module basic_500_3000_500_40_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_309,In_449);
nor U1 (N_1,In_281,In_157);
nor U2 (N_2,In_391,In_463);
and U3 (N_3,In_326,In_52);
nand U4 (N_4,In_422,In_261);
and U5 (N_5,In_153,In_464);
nor U6 (N_6,In_99,In_476);
or U7 (N_7,In_176,In_138);
and U8 (N_8,In_260,In_252);
nand U9 (N_9,In_368,In_336);
and U10 (N_10,In_384,In_226);
and U11 (N_11,In_251,In_298);
nand U12 (N_12,In_358,In_144);
nor U13 (N_13,In_338,In_125);
nand U14 (N_14,In_340,In_42);
and U15 (N_15,In_345,In_308);
nor U16 (N_16,In_161,In_342);
or U17 (N_17,In_407,In_201);
nor U18 (N_18,In_3,In_271);
and U19 (N_19,In_137,In_12);
or U20 (N_20,In_243,In_447);
and U21 (N_21,In_155,In_113);
and U22 (N_22,In_423,In_275);
nand U23 (N_23,In_96,In_36);
nand U24 (N_24,In_34,In_288);
and U25 (N_25,In_499,In_300);
and U26 (N_26,In_483,In_87);
xor U27 (N_27,In_428,In_418);
nor U28 (N_28,In_285,In_445);
nor U29 (N_29,In_453,In_146);
nand U30 (N_30,In_236,In_71);
nor U31 (N_31,In_2,In_51);
or U32 (N_32,In_235,In_13);
nor U33 (N_33,In_98,In_208);
and U34 (N_34,In_493,In_439);
and U35 (N_35,In_192,In_92);
and U36 (N_36,In_492,In_101);
nor U37 (N_37,In_451,In_294);
or U38 (N_38,In_389,In_16);
and U39 (N_39,In_323,In_297);
nand U40 (N_40,In_459,In_435);
nand U41 (N_41,In_373,In_434);
nor U42 (N_42,In_387,In_145);
nand U43 (N_43,In_234,In_420);
nand U44 (N_44,In_202,In_331);
and U45 (N_45,In_303,In_238);
nand U46 (N_46,In_468,In_398);
or U47 (N_47,In_307,In_286);
nand U48 (N_48,In_410,In_403);
and U49 (N_49,In_170,In_258);
or U50 (N_50,In_211,In_344);
nor U51 (N_51,In_124,In_86);
and U52 (N_52,In_458,In_262);
nand U53 (N_53,In_195,In_363);
nor U54 (N_54,In_355,In_390);
nor U55 (N_55,In_200,In_315);
and U56 (N_56,In_26,In_94);
or U57 (N_57,In_359,In_205);
and U58 (N_58,In_7,In_247);
nand U59 (N_59,In_479,In_40);
or U60 (N_60,In_77,In_379);
nor U61 (N_61,In_119,In_53);
nor U62 (N_62,In_54,In_227);
or U63 (N_63,In_18,In_218);
or U64 (N_64,In_497,In_282);
and U65 (N_65,In_267,In_107);
xor U66 (N_66,In_454,In_478);
and U67 (N_67,In_246,In_5);
and U68 (N_68,In_450,In_470);
and U69 (N_69,In_278,In_240);
and U70 (N_70,In_184,In_9);
or U71 (N_71,In_109,In_217);
or U72 (N_72,In_498,In_20);
nor U73 (N_73,In_381,In_215);
and U74 (N_74,In_228,In_102);
and U75 (N_75,N_34,In_47);
or U76 (N_76,N_47,In_474);
and U77 (N_77,In_22,In_78);
nand U78 (N_78,N_52,In_393);
and U79 (N_79,In_296,In_123);
or U80 (N_80,In_335,In_382);
or U81 (N_81,In_305,In_438);
nor U82 (N_82,In_62,N_60);
or U83 (N_83,In_84,In_370);
and U84 (N_84,In_245,In_491);
or U85 (N_85,In_82,In_224);
nand U86 (N_86,In_333,In_142);
and U87 (N_87,In_120,N_41);
nand U88 (N_88,In_477,In_490);
nand U89 (N_89,In_166,In_306);
nand U90 (N_90,In_116,In_0);
or U91 (N_91,In_241,In_291);
nor U92 (N_92,In_229,In_356);
and U93 (N_93,In_143,In_399);
nand U94 (N_94,In_104,N_5);
nand U95 (N_95,In_473,In_462);
or U96 (N_96,In_214,In_11);
and U97 (N_97,In_110,In_437);
nand U98 (N_98,In_495,N_38);
xnor U99 (N_99,In_83,In_351);
nand U100 (N_100,In_253,In_225);
nor U101 (N_101,In_48,In_386);
or U102 (N_102,N_3,In_349);
and U103 (N_103,In_179,In_374);
or U104 (N_104,In_429,In_206);
nand U105 (N_105,In_219,In_128);
and U106 (N_106,In_369,In_264);
and U107 (N_107,In_310,N_66);
nand U108 (N_108,N_10,In_209);
nor U109 (N_109,In_117,In_321);
or U110 (N_110,N_18,In_45);
and U111 (N_111,N_58,In_289);
nand U112 (N_112,In_317,In_149);
nor U113 (N_113,In_89,In_172);
or U114 (N_114,In_38,In_159);
or U115 (N_115,In_322,N_62);
nor U116 (N_116,In_332,In_133);
and U117 (N_117,In_160,In_352);
nand U118 (N_118,In_55,In_85);
and U119 (N_119,N_49,In_314);
nand U120 (N_120,N_67,N_53);
or U121 (N_121,In_233,In_348);
nand U122 (N_122,N_2,In_480);
nand U123 (N_123,N_14,In_402);
or U124 (N_124,In_248,In_199);
nor U125 (N_125,In_396,In_198);
or U126 (N_126,In_57,In_266);
nor U127 (N_127,In_293,In_140);
xnor U128 (N_128,In_24,In_421);
nand U129 (N_129,In_457,In_88);
nand U130 (N_130,N_63,In_4);
xnor U131 (N_131,In_136,In_268);
or U132 (N_132,In_416,In_183);
or U133 (N_133,In_482,N_72);
or U134 (N_134,In_371,N_17);
or U135 (N_135,In_397,In_460);
nor U136 (N_136,N_36,In_162);
or U137 (N_137,In_156,In_486);
nor U138 (N_138,In_61,N_64);
and U139 (N_139,In_360,N_69);
and U140 (N_140,In_412,In_175);
nand U141 (N_141,In_442,In_93);
nor U142 (N_142,In_181,N_59);
and U143 (N_143,In_173,In_167);
or U144 (N_144,In_485,In_191);
nand U145 (N_145,In_446,In_272);
or U146 (N_146,N_23,N_68);
or U147 (N_147,In_90,In_400);
nor U148 (N_148,In_150,In_452);
or U149 (N_149,In_204,In_406);
nand U150 (N_150,In_425,In_32);
nor U151 (N_151,N_120,N_142);
nor U152 (N_152,N_105,In_171);
nor U153 (N_153,In_121,In_318);
and U154 (N_154,N_108,In_432);
nor U155 (N_155,N_1,In_430);
nand U156 (N_156,In_91,In_250);
nand U157 (N_157,In_372,In_50);
nor U158 (N_158,N_99,In_312);
or U159 (N_159,In_64,In_455);
and U160 (N_160,In_196,N_54);
or U161 (N_161,In_216,In_465);
nand U162 (N_162,N_121,In_223);
and U163 (N_163,N_82,In_44);
nor U164 (N_164,In_14,N_75);
nor U165 (N_165,In_466,In_259);
or U166 (N_166,In_174,In_254);
and U167 (N_167,In_395,In_106);
and U168 (N_168,N_141,In_31);
nor U169 (N_169,N_28,N_21);
and U170 (N_170,In_456,In_30);
nor U171 (N_171,N_127,In_320);
and U172 (N_172,N_70,In_154);
nor U173 (N_173,In_194,In_164);
or U174 (N_174,In_231,N_100);
or U175 (N_175,In_213,N_115);
and U176 (N_176,In_496,In_242);
nor U177 (N_177,In_58,N_143);
nor U178 (N_178,In_239,N_39);
nand U179 (N_179,N_81,In_188);
or U180 (N_180,N_16,In_68);
and U181 (N_181,In_256,N_125);
nor U182 (N_182,In_427,In_367);
nor U183 (N_183,In_378,In_168);
or U184 (N_184,N_84,In_301);
nor U185 (N_185,N_122,In_377);
xor U186 (N_186,In_302,N_24);
nor U187 (N_187,In_112,In_385);
and U188 (N_188,In_280,In_424);
and U189 (N_189,In_19,In_75);
and U190 (N_190,In_221,N_114);
and U191 (N_191,N_19,N_22);
and U192 (N_192,In_292,N_149);
nor U193 (N_193,N_78,N_111);
and U194 (N_194,In_97,In_274);
nor U195 (N_195,In_290,In_265);
or U196 (N_196,N_98,In_489);
or U197 (N_197,In_132,In_66);
and U198 (N_198,N_136,In_383);
and U199 (N_199,In_152,In_433);
and U200 (N_200,In_79,In_43);
and U201 (N_201,In_187,N_80);
nand U202 (N_202,In_27,In_1);
or U203 (N_203,N_29,In_277);
xor U204 (N_204,In_376,In_494);
nand U205 (N_205,In_313,In_444);
nand U206 (N_206,In_108,In_413);
nand U207 (N_207,In_284,In_366);
nor U208 (N_208,In_65,N_85);
nand U209 (N_209,In_73,In_401);
or U210 (N_210,In_273,In_461);
nor U211 (N_211,In_111,In_255);
and U212 (N_212,N_133,In_165);
nor U213 (N_213,In_375,In_114);
or U214 (N_214,N_119,N_117);
and U215 (N_215,In_67,N_131);
nand U216 (N_216,In_270,N_20);
or U217 (N_217,In_60,In_276);
nand U218 (N_218,N_86,N_33);
and U219 (N_219,N_124,In_10);
or U220 (N_220,N_4,In_394);
nor U221 (N_221,N_103,In_139);
or U222 (N_222,In_441,N_106);
nor U223 (N_223,In_190,In_177);
nand U224 (N_224,In_304,N_96);
nand U225 (N_225,In_207,In_388);
and U226 (N_226,In_417,N_224);
or U227 (N_227,In_431,N_31);
nor U228 (N_228,In_80,N_116);
nand U229 (N_229,N_154,N_89);
and U230 (N_230,In_122,In_100);
or U231 (N_231,N_93,N_197);
and U232 (N_232,In_127,N_43);
and U233 (N_233,N_137,N_8);
and U234 (N_234,In_354,In_203);
nor U235 (N_235,In_118,In_448);
or U236 (N_236,In_295,N_175);
or U237 (N_237,N_40,In_440);
or U238 (N_238,In_63,N_91);
and U239 (N_239,N_210,In_443);
nor U240 (N_240,In_279,N_88);
and U241 (N_241,In_404,In_212);
xnor U242 (N_242,In_23,N_205);
nand U243 (N_243,N_13,N_152);
or U244 (N_244,In_134,In_249);
or U245 (N_245,N_139,N_61);
nor U246 (N_246,In_411,In_319);
and U247 (N_247,N_76,In_299);
and U248 (N_248,In_182,In_76);
or U249 (N_249,N_161,In_28);
or U250 (N_250,N_0,N_219);
nand U251 (N_251,N_158,N_55);
or U252 (N_252,N_192,In_141);
nand U253 (N_253,N_213,N_184);
nand U254 (N_254,N_6,N_190);
and U255 (N_255,In_8,N_128);
and U256 (N_256,N_207,N_144);
nand U257 (N_257,N_153,In_6);
nor U258 (N_258,In_37,N_50);
or U259 (N_259,In_469,N_7);
xnor U260 (N_260,In_35,N_57);
or U261 (N_261,In_180,N_37);
and U262 (N_262,In_316,In_15);
or U263 (N_263,N_25,N_138);
nor U264 (N_264,N_107,In_475);
and U265 (N_265,In_364,N_156);
nand U266 (N_266,In_409,In_263);
or U267 (N_267,N_186,N_45);
and U268 (N_268,N_223,In_237);
nand U269 (N_269,N_162,In_337);
or U270 (N_270,In_69,N_216);
and U271 (N_271,In_327,N_217);
nand U272 (N_272,N_65,N_44);
nand U273 (N_273,In_419,In_471);
nand U274 (N_274,N_179,In_21);
nand U275 (N_275,N_159,N_206);
and U276 (N_276,In_472,N_180);
or U277 (N_277,In_484,In_56);
or U278 (N_278,N_71,In_41);
nor U279 (N_279,N_170,In_357);
nor U280 (N_280,N_87,N_178);
nor U281 (N_281,N_211,N_166);
or U282 (N_282,N_167,In_230);
nand U283 (N_283,N_164,In_467);
nor U284 (N_284,In_59,In_380);
xor U285 (N_285,In_329,N_203);
or U286 (N_286,In_426,In_186);
nand U287 (N_287,N_73,N_208);
nand U288 (N_288,N_126,In_33);
and U289 (N_289,N_15,In_330);
nand U290 (N_290,N_30,N_12);
or U291 (N_291,N_157,N_168);
and U292 (N_292,N_11,N_176);
nor U293 (N_293,In_126,N_209);
nor U294 (N_294,N_182,In_135);
nor U295 (N_295,In_287,N_174);
and U296 (N_296,N_160,N_9);
or U297 (N_297,N_200,N_169);
nand U298 (N_298,In_488,N_222);
and U299 (N_299,In_324,In_341);
or U300 (N_300,N_291,In_115);
nand U301 (N_301,In_405,In_362);
and U302 (N_302,In_189,N_140);
or U303 (N_303,In_95,N_248);
nor U304 (N_304,N_294,N_283);
nor U305 (N_305,N_260,N_256);
nor U306 (N_306,N_193,N_173);
and U307 (N_307,N_79,In_343);
nor U308 (N_308,In_129,N_237);
nand U309 (N_309,In_487,In_169);
nor U310 (N_310,N_46,N_282);
and U311 (N_311,In_72,N_266);
or U312 (N_312,In_70,N_239);
nor U313 (N_313,N_97,N_241);
or U314 (N_314,N_236,In_151);
nand U315 (N_315,In_415,N_92);
nor U316 (N_316,In_283,N_238);
or U317 (N_317,N_253,N_129);
or U318 (N_318,N_181,In_350);
nor U319 (N_319,N_146,N_280);
or U320 (N_320,N_250,N_276);
and U321 (N_321,N_271,N_287);
nor U322 (N_322,In_147,N_102);
nor U323 (N_323,In_436,In_29);
nor U324 (N_324,N_195,In_414);
xnor U325 (N_325,In_103,N_185);
nor U326 (N_326,N_56,N_90);
or U327 (N_327,N_163,In_148);
nor U328 (N_328,N_296,N_252);
and U329 (N_329,N_279,N_135);
and U330 (N_330,N_274,N_225);
or U331 (N_331,N_147,N_242);
or U332 (N_332,N_187,N_220);
or U333 (N_333,N_151,In_178);
and U334 (N_334,In_105,In_220);
and U335 (N_335,In_257,N_234);
or U336 (N_336,In_334,In_347);
nor U337 (N_337,In_131,N_299);
nand U338 (N_338,N_148,In_361);
nand U339 (N_339,In_197,N_229);
nor U340 (N_340,N_255,In_25);
nand U341 (N_341,In_325,N_261);
nand U342 (N_342,N_113,N_215);
nand U343 (N_343,N_257,In_269);
xor U344 (N_344,N_110,N_251);
or U345 (N_345,N_214,N_204);
nand U346 (N_346,N_228,N_145);
and U347 (N_347,In_346,N_221);
and U348 (N_348,In_210,In_232);
nand U349 (N_349,N_83,N_189);
nor U350 (N_350,N_244,In_81);
nor U351 (N_351,N_290,N_285);
and U352 (N_352,N_273,N_281);
nand U353 (N_353,In_39,N_284);
nor U354 (N_354,In_74,In_46);
or U355 (N_355,N_230,N_202);
and U356 (N_356,In_222,N_235);
nand U357 (N_357,N_191,N_288);
and U358 (N_358,N_123,N_245);
or U359 (N_359,In_193,N_246);
or U360 (N_360,N_101,N_165);
or U361 (N_361,N_94,N_172);
nand U362 (N_362,N_268,N_95);
and U363 (N_363,In_49,N_249);
nor U364 (N_364,N_275,N_212);
nand U365 (N_365,N_263,N_289);
nand U366 (N_366,N_262,N_232);
nand U367 (N_367,N_254,N_278);
nand U368 (N_368,In_353,N_231);
nor U369 (N_369,N_196,In_328);
nand U370 (N_370,N_32,N_295);
and U371 (N_371,N_109,N_177);
nor U372 (N_372,In_244,N_243);
nor U373 (N_373,In_185,N_297);
and U374 (N_374,N_150,In_311);
nand U375 (N_375,N_130,N_310);
or U376 (N_376,N_306,N_338);
nand U377 (N_377,N_334,N_331);
nor U378 (N_378,N_360,N_26);
and U379 (N_379,N_201,N_363);
and U380 (N_380,N_155,N_312);
nor U381 (N_381,N_339,N_301);
and U382 (N_382,In_408,In_17);
and U383 (N_383,N_335,N_258);
nand U384 (N_384,N_233,N_315);
xnor U385 (N_385,N_303,N_362);
or U386 (N_386,N_272,N_330);
and U387 (N_387,N_328,N_345);
and U388 (N_388,N_286,N_227);
nand U389 (N_389,N_118,N_341);
and U390 (N_390,N_259,N_307);
nor U391 (N_391,N_359,N_269);
and U392 (N_392,In_130,N_368);
nand U393 (N_393,N_198,N_74);
or U394 (N_394,N_264,N_51);
nand U395 (N_395,N_270,N_293);
nand U396 (N_396,N_320,In_163);
nor U397 (N_397,N_370,N_322);
nor U398 (N_398,N_374,N_298);
and U399 (N_399,N_48,N_240);
or U400 (N_400,N_352,N_369);
xnor U401 (N_401,N_361,N_325);
nand U402 (N_402,N_357,In_392);
and U403 (N_403,N_42,N_188);
xor U404 (N_404,N_302,N_171);
and U405 (N_405,N_323,N_354);
nor U406 (N_406,N_27,N_311);
and U407 (N_407,N_277,N_358);
or U408 (N_408,In_365,N_218);
and U409 (N_409,N_247,N_366);
and U410 (N_410,N_308,N_342);
xor U411 (N_411,N_104,N_355);
nor U412 (N_412,N_321,In_339);
and U413 (N_413,N_356,N_313);
nand U414 (N_414,N_183,N_132);
or U415 (N_415,N_347,N_327);
or U416 (N_416,N_292,N_314);
nor U417 (N_417,N_351,N_346);
and U418 (N_418,N_324,N_317);
nor U419 (N_419,N_77,N_367);
and U420 (N_420,N_112,N_336);
or U421 (N_421,In_158,N_305);
nor U422 (N_422,N_365,N_329);
or U423 (N_423,N_340,N_343);
nor U424 (N_424,N_316,N_353);
nand U425 (N_425,N_319,N_309);
or U426 (N_426,N_348,N_134);
nor U427 (N_427,N_332,N_300);
nor U428 (N_428,N_373,N_337);
and U429 (N_429,N_371,N_265);
nor U430 (N_430,N_344,N_267);
and U431 (N_431,In_481,N_326);
nand U432 (N_432,N_226,N_35);
nor U433 (N_433,N_333,N_304);
and U434 (N_434,N_199,N_194);
or U435 (N_435,N_350,N_364);
nand U436 (N_436,N_318,N_349);
nand U437 (N_437,N_372,N_331);
nand U438 (N_438,N_338,N_344);
and U439 (N_439,In_408,N_272);
nand U440 (N_440,N_240,N_302);
nor U441 (N_441,N_316,N_198);
and U442 (N_442,N_314,N_233);
nand U443 (N_443,N_312,N_345);
nand U444 (N_444,In_365,N_369);
nand U445 (N_445,N_272,N_48);
or U446 (N_446,N_306,N_363);
and U447 (N_447,N_218,N_343);
or U448 (N_448,N_337,N_365);
and U449 (N_449,N_322,N_48);
and U450 (N_450,N_443,N_393);
nand U451 (N_451,N_417,N_399);
and U452 (N_452,N_375,N_397);
and U453 (N_453,N_413,N_447);
or U454 (N_454,N_438,N_446);
or U455 (N_455,N_392,N_376);
nand U456 (N_456,N_379,N_418);
and U457 (N_457,N_406,N_440);
nand U458 (N_458,N_423,N_433);
nand U459 (N_459,N_429,N_449);
nand U460 (N_460,N_431,N_437);
nor U461 (N_461,N_408,N_420);
xor U462 (N_462,N_395,N_445);
nor U463 (N_463,N_402,N_394);
nand U464 (N_464,N_386,N_409);
nor U465 (N_465,N_427,N_400);
nor U466 (N_466,N_382,N_434);
nor U467 (N_467,N_390,N_380);
and U468 (N_468,N_435,N_412);
and U469 (N_469,N_416,N_442);
nor U470 (N_470,N_405,N_385);
nand U471 (N_471,N_401,N_388);
xnor U472 (N_472,N_387,N_398);
nor U473 (N_473,N_448,N_384);
or U474 (N_474,N_389,N_404);
nand U475 (N_475,N_407,N_428);
nand U476 (N_476,N_425,N_424);
and U477 (N_477,N_391,N_439);
nor U478 (N_478,N_414,N_410);
nor U479 (N_479,N_436,N_378);
nand U480 (N_480,N_430,N_415);
nand U481 (N_481,N_381,N_444);
or U482 (N_482,N_383,N_419);
or U483 (N_483,N_421,N_403);
or U484 (N_484,N_422,N_377);
and U485 (N_485,N_426,N_441);
and U486 (N_486,N_396,N_432);
nand U487 (N_487,N_411,N_443);
nor U488 (N_488,N_425,N_403);
and U489 (N_489,N_436,N_380);
and U490 (N_490,N_383,N_421);
nor U491 (N_491,N_385,N_433);
nor U492 (N_492,N_391,N_382);
nor U493 (N_493,N_380,N_388);
and U494 (N_494,N_392,N_398);
xor U495 (N_495,N_428,N_400);
nand U496 (N_496,N_378,N_379);
xnor U497 (N_497,N_390,N_446);
nand U498 (N_498,N_406,N_444);
and U499 (N_499,N_419,N_436);
and U500 (N_500,N_435,N_391);
and U501 (N_501,N_402,N_377);
or U502 (N_502,N_415,N_425);
nand U503 (N_503,N_434,N_403);
and U504 (N_504,N_404,N_431);
and U505 (N_505,N_437,N_432);
nand U506 (N_506,N_387,N_429);
nand U507 (N_507,N_395,N_394);
nand U508 (N_508,N_378,N_415);
and U509 (N_509,N_433,N_400);
or U510 (N_510,N_418,N_440);
or U511 (N_511,N_407,N_394);
nor U512 (N_512,N_403,N_385);
and U513 (N_513,N_378,N_419);
nor U514 (N_514,N_413,N_436);
nor U515 (N_515,N_383,N_388);
and U516 (N_516,N_388,N_430);
and U517 (N_517,N_406,N_432);
and U518 (N_518,N_406,N_413);
nor U519 (N_519,N_377,N_449);
and U520 (N_520,N_433,N_375);
and U521 (N_521,N_427,N_423);
and U522 (N_522,N_380,N_431);
and U523 (N_523,N_426,N_391);
and U524 (N_524,N_442,N_404);
and U525 (N_525,N_465,N_506);
nor U526 (N_526,N_492,N_521);
or U527 (N_527,N_457,N_516);
or U528 (N_528,N_470,N_487);
nand U529 (N_529,N_501,N_514);
or U530 (N_530,N_518,N_494);
nand U531 (N_531,N_462,N_504);
nand U532 (N_532,N_508,N_469);
and U533 (N_533,N_451,N_483);
and U534 (N_534,N_478,N_524);
xnor U535 (N_535,N_497,N_455);
xnor U536 (N_536,N_519,N_517);
nor U537 (N_537,N_458,N_523);
nand U538 (N_538,N_480,N_481);
nor U539 (N_539,N_498,N_475);
xor U540 (N_540,N_491,N_471);
nand U541 (N_541,N_513,N_489);
nor U542 (N_542,N_520,N_450);
and U543 (N_543,N_474,N_459);
or U544 (N_544,N_496,N_482);
nor U545 (N_545,N_502,N_468);
and U546 (N_546,N_493,N_522);
and U547 (N_547,N_511,N_453);
or U548 (N_548,N_499,N_456);
and U549 (N_549,N_509,N_473);
nor U550 (N_550,N_510,N_512);
nand U551 (N_551,N_515,N_460);
and U552 (N_552,N_479,N_486);
nor U553 (N_553,N_476,N_477);
or U554 (N_554,N_467,N_485);
nand U555 (N_555,N_505,N_500);
nor U556 (N_556,N_490,N_488);
or U557 (N_557,N_472,N_466);
or U558 (N_558,N_484,N_463);
and U559 (N_559,N_503,N_507);
and U560 (N_560,N_495,N_454);
or U561 (N_561,N_464,N_461);
and U562 (N_562,N_452,N_450);
nand U563 (N_563,N_492,N_491);
nand U564 (N_564,N_470,N_490);
nor U565 (N_565,N_471,N_494);
nand U566 (N_566,N_454,N_492);
xor U567 (N_567,N_494,N_462);
nor U568 (N_568,N_523,N_521);
nand U569 (N_569,N_498,N_472);
xor U570 (N_570,N_495,N_476);
and U571 (N_571,N_450,N_497);
nand U572 (N_572,N_493,N_465);
and U573 (N_573,N_495,N_475);
and U574 (N_574,N_513,N_485);
xnor U575 (N_575,N_500,N_466);
or U576 (N_576,N_494,N_473);
nor U577 (N_577,N_474,N_509);
and U578 (N_578,N_489,N_465);
and U579 (N_579,N_462,N_510);
nor U580 (N_580,N_504,N_498);
and U581 (N_581,N_485,N_454);
and U582 (N_582,N_505,N_470);
nor U583 (N_583,N_472,N_492);
or U584 (N_584,N_451,N_477);
or U585 (N_585,N_520,N_453);
and U586 (N_586,N_471,N_500);
or U587 (N_587,N_510,N_513);
or U588 (N_588,N_523,N_495);
or U589 (N_589,N_468,N_486);
nor U590 (N_590,N_511,N_501);
nand U591 (N_591,N_515,N_498);
and U592 (N_592,N_462,N_480);
or U593 (N_593,N_458,N_486);
and U594 (N_594,N_507,N_502);
nor U595 (N_595,N_473,N_454);
and U596 (N_596,N_474,N_499);
nand U597 (N_597,N_486,N_466);
nand U598 (N_598,N_459,N_473);
nand U599 (N_599,N_512,N_450);
or U600 (N_600,N_543,N_579);
nand U601 (N_601,N_564,N_554);
and U602 (N_602,N_532,N_562);
nand U603 (N_603,N_567,N_549);
nor U604 (N_604,N_528,N_575);
nor U605 (N_605,N_584,N_566);
or U606 (N_606,N_590,N_547);
or U607 (N_607,N_538,N_537);
nor U608 (N_608,N_586,N_560);
xnor U609 (N_609,N_536,N_594);
nand U610 (N_610,N_550,N_571);
nor U611 (N_611,N_548,N_599);
nand U612 (N_612,N_572,N_525);
nand U613 (N_613,N_540,N_527);
nand U614 (N_614,N_568,N_577);
and U615 (N_615,N_593,N_592);
nand U616 (N_616,N_574,N_555);
and U617 (N_617,N_541,N_529);
and U618 (N_618,N_576,N_556);
nor U619 (N_619,N_563,N_573);
nor U620 (N_620,N_581,N_558);
and U621 (N_621,N_539,N_552);
nand U622 (N_622,N_580,N_561);
or U623 (N_623,N_589,N_565);
and U624 (N_624,N_591,N_533);
or U625 (N_625,N_582,N_557);
nand U626 (N_626,N_526,N_534);
and U627 (N_627,N_551,N_569);
nor U628 (N_628,N_535,N_531);
and U629 (N_629,N_545,N_587);
and U630 (N_630,N_578,N_546);
and U631 (N_631,N_597,N_598);
nand U632 (N_632,N_559,N_553);
and U633 (N_633,N_596,N_544);
or U634 (N_634,N_542,N_570);
nand U635 (N_635,N_585,N_588);
and U636 (N_636,N_583,N_530);
or U637 (N_637,N_595,N_581);
nor U638 (N_638,N_534,N_555);
nor U639 (N_639,N_553,N_571);
nor U640 (N_640,N_578,N_543);
nor U641 (N_641,N_526,N_597);
nand U642 (N_642,N_546,N_528);
and U643 (N_643,N_584,N_583);
or U644 (N_644,N_555,N_558);
nand U645 (N_645,N_557,N_579);
nor U646 (N_646,N_588,N_536);
or U647 (N_647,N_576,N_540);
and U648 (N_648,N_568,N_530);
nor U649 (N_649,N_578,N_551);
or U650 (N_650,N_554,N_571);
and U651 (N_651,N_592,N_576);
and U652 (N_652,N_585,N_590);
nand U653 (N_653,N_546,N_581);
or U654 (N_654,N_589,N_550);
nor U655 (N_655,N_570,N_553);
nor U656 (N_656,N_548,N_558);
and U657 (N_657,N_535,N_559);
or U658 (N_658,N_546,N_570);
or U659 (N_659,N_532,N_527);
nor U660 (N_660,N_567,N_565);
and U661 (N_661,N_566,N_539);
or U662 (N_662,N_535,N_565);
or U663 (N_663,N_570,N_535);
and U664 (N_664,N_541,N_558);
nand U665 (N_665,N_557,N_536);
nand U666 (N_666,N_586,N_553);
nor U667 (N_667,N_557,N_597);
and U668 (N_668,N_570,N_528);
or U669 (N_669,N_557,N_573);
nor U670 (N_670,N_552,N_561);
or U671 (N_671,N_596,N_551);
xor U672 (N_672,N_579,N_592);
nor U673 (N_673,N_571,N_585);
and U674 (N_674,N_546,N_591);
nand U675 (N_675,N_626,N_664);
xnor U676 (N_676,N_611,N_660);
or U677 (N_677,N_651,N_638);
nor U678 (N_678,N_603,N_605);
nand U679 (N_679,N_645,N_640);
nor U680 (N_680,N_606,N_641);
xnor U681 (N_681,N_653,N_629);
and U682 (N_682,N_618,N_615);
and U683 (N_683,N_636,N_637);
nand U684 (N_684,N_617,N_642);
and U685 (N_685,N_608,N_609);
or U686 (N_686,N_639,N_625);
nand U687 (N_687,N_600,N_658);
nand U688 (N_688,N_654,N_632);
and U689 (N_689,N_610,N_635);
nand U690 (N_690,N_647,N_627);
and U691 (N_691,N_649,N_604);
nor U692 (N_692,N_631,N_646);
nor U693 (N_693,N_624,N_663);
or U694 (N_694,N_622,N_628);
or U695 (N_695,N_665,N_620);
and U696 (N_696,N_671,N_672);
nor U697 (N_697,N_657,N_633);
nor U698 (N_698,N_602,N_655);
nand U699 (N_699,N_612,N_607);
nor U700 (N_700,N_601,N_644);
nor U701 (N_701,N_648,N_630);
nor U702 (N_702,N_652,N_668);
nor U703 (N_703,N_656,N_661);
nor U704 (N_704,N_670,N_643);
nand U705 (N_705,N_673,N_623);
and U706 (N_706,N_619,N_613);
nand U707 (N_707,N_666,N_659);
or U708 (N_708,N_614,N_634);
nor U709 (N_709,N_662,N_667);
and U710 (N_710,N_674,N_669);
or U711 (N_711,N_650,N_616);
nor U712 (N_712,N_621,N_634);
nor U713 (N_713,N_621,N_653);
xor U714 (N_714,N_634,N_603);
nand U715 (N_715,N_661,N_659);
nor U716 (N_716,N_603,N_630);
and U717 (N_717,N_602,N_648);
or U718 (N_718,N_612,N_631);
and U719 (N_719,N_606,N_661);
or U720 (N_720,N_663,N_659);
nor U721 (N_721,N_644,N_658);
nor U722 (N_722,N_653,N_610);
nand U723 (N_723,N_669,N_618);
and U724 (N_724,N_662,N_601);
and U725 (N_725,N_641,N_616);
nand U726 (N_726,N_637,N_613);
nor U727 (N_727,N_644,N_632);
or U728 (N_728,N_656,N_648);
and U729 (N_729,N_610,N_629);
or U730 (N_730,N_612,N_639);
nor U731 (N_731,N_653,N_674);
or U732 (N_732,N_630,N_671);
and U733 (N_733,N_611,N_671);
xnor U734 (N_734,N_620,N_650);
and U735 (N_735,N_661,N_657);
and U736 (N_736,N_620,N_627);
nor U737 (N_737,N_655,N_653);
and U738 (N_738,N_653,N_601);
or U739 (N_739,N_642,N_619);
and U740 (N_740,N_637,N_641);
and U741 (N_741,N_627,N_614);
nor U742 (N_742,N_658,N_619);
nand U743 (N_743,N_640,N_607);
nand U744 (N_744,N_600,N_619);
and U745 (N_745,N_660,N_639);
nor U746 (N_746,N_662,N_672);
and U747 (N_747,N_665,N_667);
or U748 (N_748,N_660,N_601);
nand U749 (N_749,N_662,N_614);
nand U750 (N_750,N_735,N_709);
and U751 (N_751,N_677,N_679);
and U752 (N_752,N_703,N_739);
nor U753 (N_753,N_733,N_742);
or U754 (N_754,N_696,N_746);
or U755 (N_755,N_734,N_744);
and U756 (N_756,N_705,N_690);
nor U757 (N_757,N_687,N_730);
or U758 (N_758,N_745,N_678);
and U759 (N_759,N_694,N_743);
nor U760 (N_760,N_736,N_700);
or U761 (N_761,N_741,N_718);
nor U762 (N_762,N_714,N_721);
or U763 (N_763,N_698,N_686);
or U764 (N_764,N_747,N_702);
nand U765 (N_765,N_717,N_737);
and U766 (N_766,N_681,N_684);
nor U767 (N_767,N_712,N_728);
or U768 (N_768,N_689,N_722);
and U769 (N_769,N_693,N_716);
nand U770 (N_770,N_692,N_699);
nand U771 (N_771,N_729,N_740);
and U772 (N_772,N_688,N_710);
or U773 (N_773,N_706,N_707);
nand U774 (N_774,N_738,N_723);
nand U775 (N_775,N_697,N_704);
and U776 (N_776,N_748,N_724);
and U777 (N_777,N_675,N_680);
or U778 (N_778,N_713,N_682);
and U779 (N_779,N_727,N_749);
nor U780 (N_780,N_726,N_711);
and U781 (N_781,N_695,N_720);
and U782 (N_782,N_685,N_676);
nor U783 (N_783,N_708,N_725);
nand U784 (N_784,N_691,N_719);
or U785 (N_785,N_731,N_683);
xor U786 (N_786,N_715,N_701);
and U787 (N_787,N_732,N_747);
nand U788 (N_788,N_746,N_737);
nand U789 (N_789,N_734,N_702);
or U790 (N_790,N_744,N_735);
or U791 (N_791,N_734,N_696);
nor U792 (N_792,N_746,N_723);
xor U793 (N_793,N_691,N_709);
and U794 (N_794,N_692,N_730);
nand U795 (N_795,N_730,N_744);
nor U796 (N_796,N_719,N_707);
or U797 (N_797,N_720,N_707);
nand U798 (N_798,N_707,N_687);
and U799 (N_799,N_740,N_747);
or U800 (N_800,N_739,N_682);
nand U801 (N_801,N_741,N_703);
nor U802 (N_802,N_684,N_719);
nand U803 (N_803,N_721,N_697);
nor U804 (N_804,N_725,N_687);
nand U805 (N_805,N_688,N_678);
and U806 (N_806,N_710,N_743);
nand U807 (N_807,N_745,N_719);
nand U808 (N_808,N_685,N_698);
nor U809 (N_809,N_695,N_712);
and U810 (N_810,N_719,N_739);
nand U811 (N_811,N_746,N_713);
or U812 (N_812,N_702,N_723);
or U813 (N_813,N_728,N_746);
and U814 (N_814,N_713,N_678);
nand U815 (N_815,N_738,N_745);
and U816 (N_816,N_701,N_722);
xnor U817 (N_817,N_694,N_691);
nor U818 (N_818,N_680,N_692);
xnor U819 (N_819,N_709,N_718);
nand U820 (N_820,N_748,N_723);
or U821 (N_821,N_729,N_747);
and U822 (N_822,N_740,N_713);
nand U823 (N_823,N_695,N_728);
nand U824 (N_824,N_740,N_745);
and U825 (N_825,N_768,N_762);
nand U826 (N_826,N_800,N_815);
xor U827 (N_827,N_752,N_787);
and U828 (N_828,N_773,N_781);
and U829 (N_829,N_769,N_804);
nand U830 (N_830,N_816,N_779);
or U831 (N_831,N_756,N_788);
nor U832 (N_832,N_765,N_820);
nor U833 (N_833,N_817,N_780);
or U834 (N_834,N_822,N_758);
and U835 (N_835,N_754,N_801);
or U836 (N_836,N_782,N_819);
nand U837 (N_837,N_814,N_807);
and U838 (N_838,N_750,N_789);
nand U839 (N_839,N_823,N_778);
nor U840 (N_840,N_790,N_795);
nand U841 (N_841,N_767,N_810);
nor U842 (N_842,N_776,N_813);
nor U843 (N_843,N_757,N_783);
nor U844 (N_844,N_811,N_802);
nor U845 (N_845,N_803,N_821);
or U846 (N_846,N_785,N_808);
or U847 (N_847,N_784,N_755);
or U848 (N_848,N_792,N_775);
nand U849 (N_849,N_774,N_824);
nor U850 (N_850,N_753,N_771);
nand U851 (N_851,N_798,N_772);
and U852 (N_852,N_794,N_760);
nand U853 (N_853,N_796,N_786);
or U854 (N_854,N_770,N_791);
and U855 (N_855,N_799,N_777);
and U856 (N_856,N_763,N_809);
or U857 (N_857,N_764,N_805);
or U858 (N_858,N_797,N_806);
and U859 (N_859,N_818,N_751);
or U860 (N_860,N_766,N_761);
nand U861 (N_861,N_812,N_793);
nand U862 (N_862,N_759,N_760);
nand U863 (N_863,N_813,N_756);
and U864 (N_864,N_785,N_816);
and U865 (N_865,N_799,N_758);
nor U866 (N_866,N_788,N_766);
nand U867 (N_867,N_807,N_753);
nor U868 (N_868,N_772,N_752);
nand U869 (N_869,N_816,N_799);
nand U870 (N_870,N_755,N_760);
nand U871 (N_871,N_812,N_795);
nand U872 (N_872,N_811,N_805);
and U873 (N_873,N_751,N_790);
or U874 (N_874,N_812,N_765);
or U875 (N_875,N_790,N_775);
nor U876 (N_876,N_819,N_759);
nor U877 (N_877,N_810,N_755);
nor U878 (N_878,N_769,N_816);
nor U879 (N_879,N_811,N_798);
nand U880 (N_880,N_753,N_797);
or U881 (N_881,N_761,N_770);
nor U882 (N_882,N_769,N_809);
nor U883 (N_883,N_807,N_799);
nand U884 (N_884,N_814,N_803);
or U885 (N_885,N_762,N_821);
or U886 (N_886,N_774,N_802);
and U887 (N_887,N_776,N_772);
nor U888 (N_888,N_761,N_769);
or U889 (N_889,N_779,N_753);
nand U890 (N_890,N_785,N_778);
nor U891 (N_891,N_796,N_804);
and U892 (N_892,N_791,N_789);
nor U893 (N_893,N_752,N_799);
or U894 (N_894,N_789,N_799);
nand U895 (N_895,N_811,N_820);
and U896 (N_896,N_797,N_792);
xnor U897 (N_897,N_751,N_783);
nor U898 (N_898,N_755,N_807);
and U899 (N_899,N_789,N_773);
nor U900 (N_900,N_842,N_846);
nor U901 (N_901,N_835,N_897);
nor U902 (N_902,N_879,N_873);
nor U903 (N_903,N_874,N_868);
nand U904 (N_904,N_862,N_839);
and U905 (N_905,N_825,N_898);
or U906 (N_906,N_895,N_899);
and U907 (N_907,N_861,N_875);
nor U908 (N_908,N_888,N_885);
or U909 (N_909,N_856,N_827);
nand U910 (N_910,N_890,N_841);
or U911 (N_911,N_860,N_864);
nor U912 (N_912,N_896,N_889);
and U913 (N_913,N_848,N_853);
and U914 (N_914,N_894,N_887);
and U915 (N_915,N_884,N_866);
xnor U916 (N_916,N_865,N_850);
nand U917 (N_917,N_833,N_859);
nand U918 (N_918,N_840,N_867);
or U919 (N_919,N_836,N_882);
and U920 (N_920,N_830,N_847);
nand U921 (N_921,N_828,N_880);
and U922 (N_922,N_832,N_886);
nor U923 (N_923,N_844,N_851);
nand U924 (N_924,N_852,N_855);
and U925 (N_925,N_857,N_831);
and U926 (N_926,N_829,N_843);
nor U927 (N_927,N_849,N_858);
and U928 (N_928,N_863,N_870);
and U929 (N_929,N_869,N_872);
and U930 (N_930,N_834,N_871);
nand U931 (N_931,N_826,N_845);
nand U932 (N_932,N_878,N_893);
and U933 (N_933,N_892,N_854);
or U934 (N_934,N_838,N_883);
nand U935 (N_935,N_881,N_891);
nor U936 (N_936,N_877,N_876);
and U937 (N_937,N_837,N_850);
and U938 (N_938,N_888,N_868);
or U939 (N_939,N_853,N_867);
or U940 (N_940,N_883,N_833);
or U941 (N_941,N_869,N_892);
or U942 (N_942,N_847,N_834);
nand U943 (N_943,N_827,N_832);
nand U944 (N_944,N_826,N_841);
nor U945 (N_945,N_864,N_859);
and U946 (N_946,N_870,N_860);
nor U947 (N_947,N_899,N_859);
nand U948 (N_948,N_854,N_842);
and U949 (N_949,N_832,N_849);
and U950 (N_950,N_850,N_855);
or U951 (N_951,N_865,N_863);
and U952 (N_952,N_847,N_836);
nand U953 (N_953,N_864,N_899);
nand U954 (N_954,N_868,N_842);
and U955 (N_955,N_855,N_874);
or U956 (N_956,N_854,N_835);
and U957 (N_957,N_842,N_896);
or U958 (N_958,N_878,N_868);
and U959 (N_959,N_882,N_826);
nor U960 (N_960,N_845,N_832);
and U961 (N_961,N_863,N_839);
nor U962 (N_962,N_880,N_839);
or U963 (N_963,N_872,N_890);
and U964 (N_964,N_834,N_885);
and U965 (N_965,N_873,N_872);
nand U966 (N_966,N_860,N_830);
and U967 (N_967,N_869,N_866);
nor U968 (N_968,N_857,N_853);
or U969 (N_969,N_852,N_891);
or U970 (N_970,N_894,N_843);
nand U971 (N_971,N_881,N_844);
xor U972 (N_972,N_827,N_854);
nand U973 (N_973,N_851,N_841);
nand U974 (N_974,N_884,N_870);
nand U975 (N_975,N_953,N_957);
or U976 (N_976,N_930,N_929);
nor U977 (N_977,N_956,N_974);
or U978 (N_978,N_964,N_907);
nand U979 (N_979,N_960,N_910);
or U980 (N_980,N_928,N_939);
or U981 (N_981,N_926,N_951);
or U982 (N_982,N_922,N_933);
nor U983 (N_983,N_940,N_943);
xor U984 (N_984,N_925,N_902);
nor U985 (N_985,N_935,N_918);
nor U986 (N_986,N_941,N_962);
and U987 (N_987,N_919,N_924);
xnor U988 (N_988,N_909,N_917);
nand U989 (N_989,N_911,N_969);
nand U990 (N_990,N_908,N_920);
or U991 (N_991,N_931,N_901);
or U992 (N_992,N_959,N_968);
nand U993 (N_993,N_949,N_973);
nand U994 (N_994,N_963,N_954);
or U995 (N_995,N_948,N_958);
nand U996 (N_996,N_904,N_937);
or U997 (N_997,N_952,N_916);
or U998 (N_998,N_936,N_938);
and U999 (N_999,N_966,N_944);
nor U1000 (N_1000,N_913,N_972);
nand U1001 (N_1001,N_945,N_946);
and U1002 (N_1002,N_923,N_900);
nor U1003 (N_1003,N_905,N_965);
nor U1004 (N_1004,N_934,N_942);
or U1005 (N_1005,N_927,N_947);
nand U1006 (N_1006,N_967,N_971);
nand U1007 (N_1007,N_903,N_955);
and U1008 (N_1008,N_932,N_970);
nor U1009 (N_1009,N_961,N_950);
nor U1010 (N_1010,N_915,N_906);
nand U1011 (N_1011,N_912,N_921);
or U1012 (N_1012,N_914,N_953);
or U1013 (N_1013,N_935,N_970);
or U1014 (N_1014,N_911,N_930);
or U1015 (N_1015,N_968,N_908);
or U1016 (N_1016,N_901,N_922);
nand U1017 (N_1017,N_922,N_904);
or U1018 (N_1018,N_958,N_935);
nand U1019 (N_1019,N_921,N_900);
or U1020 (N_1020,N_961,N_906);
and U1021 (N_1021,N_946,N_936);
and U1022 (N_1022,N_920,N_915);
or U1023 (N_1023,N_910,N_962);
or U1024 (N_1024,N_910,N_911);
nor U1025 (N_1025,N_916,N_946);
or U1026 (N_1026,N_970,N_941);
nor U1027 (N_1027,N_939,N_927);
and U1028 (N_1028,N_956,N_935);
nor U1029 (N_1029,N_962,N_920);
nand U1030 (N_1030,N_902,N_963);
and U1031 (N_1031,N_926,N_923);
or U1032 (N_1032,N_903,N_905);
and U1033 (N_1033,N_961,N_957);
or U1034 (N_1034,N_913,N_957);
and U1035 (N_1035,N_905,N_956);
nand U1036 (N_1036,N_974,N_911);
and U1037 (N_1037,N_906,N_944);
and U1038 (N_1038,N_950,N_914);
nor U1039 (N_1039,N_966,N_937);
and U1040 (N_1040,N_900,N_960);
and U1041 (N_1041,N_968,N_930);
nand U1042 (N_1042,N_961,N_943);
nand U1043 (N_1043,N_960,N_903);
and U1044 (N_1044,N_940,N_972);
nor U1045 (N_1045,N_913,N_903);
nor U1046 (N_1046,N_971,N_957);
nand U1047 (N_1047,N_973,N_970);
nand U1048 (N_1048,N_930,N_900);
nand U1049 (N_1049,N_966,N_973);
and U1050 (N_1050,N_1040,N_993);
or U1051 (N_1051,N_1017,N_1036);
nor U1052 (N_1052,N_1028,N_998);
nand U1053 (N_1053,N_1043,N_1002);
nand U1054 (N_1054,N_983,N_1039);
and U1055 (N_1055,N_988,N_1048);
nor U1056 (N_1056,N_1049,N_1023);
or U1057 (N_1057,N_994,N_984);
xor U1058 (N_1058,N_1031,N_999);
or U1059 (N_1059,N_990,N_989);
xnor U1060 (N_1060,N_1041,N_1022);
nor U1061 (N_1061,N_1046,N_1010);
nor U1062 (N_1062,N_1009,N_1025);
nand U1063 (N_1063,N_1020,N_1006);
nor U1064 (N_1064,N_981,N_1011);
nand U1065 (N_1065,N_1045,N_997);
nand U1066 (N_1066,N_1003,N_975);
or U1067 (N_1067,N_1034,N_992);
nor U1068 (N_1068,N_996,N_977);
and U1069 (N_1069,N_1016,N_995);
xnor U1070 (N_1070,N_1024,N_980);
nand U1071 (N_1071,N_986,N_1018);
nor U1072 (N_1072,N_982,N_1012);
nor U1073 (N_1073,N_1038,N_1019);
xor U1074 (N_1074,N_1027,N_1032);
and U1075 (N_1075,N_1004,N_976);
nand U1076 (N_1076,N_1013,N_1037);
nor U1077 (N_1077,N_1007,N_991);
or U1078 (N_1078,N_987,N_1035);
nor U1079 (N_1079,N_979,N_1015);
or U1080 (N_1080,N_1021,N_1014);
or U1081 (N_1081,N_1005,N_1044);
nor U1082 (N_1082,N_1001,N_1047);
or U1083 (N_1083,N_1042,N_1029);
and U1084 (N_1084,N_978,N_1008);
nand U1085 (N_1085,N_1026,N_1030);
nand U1086 (N_1086,N_985,N_1000);
and U1087 (N_1087,N_1033,N_983);
or U1088 (N_1088,N_1042,N_989);
nor U1089 (N_1089,N_985,N_998);
and U1090 (N_1090,N_1029,N_975);
and U1091 (N_1091,N_993,N_1037);
nor U1092 (N_1092,N_992,N_1015);
and U1093 (N_1093,N_992,N_1002);
and U1094 (N_1094,N_999,N_995);
or U1095 (N_1095,N_997,N_1034);
or U1096 (N_1096,N_1033,N_1011);
nor U1097 (N_1097,N_1028,N_975);
or U1098 (N_1098,N_1019,N_976);
nor U1099 (N_1099,N_1021,N_1030);
and U1100 (N_1100,N_1013,N_981);
and U1101 (N_1101,N_1034,N_1037);
nor U1102 (N_1102,N_990,N_1008);
nor U1103 (N_1103,N_1012,N_1047);
or U1104 (N_1104,N_1033,N_1029);
nand U1105 (N_1105,N_1001,N_1036);
nor U1106 (N_1106,N_1009,N_1031);
and U1107 (N_1107,N_1010,N_1043);
nor U1108 (N_1108,N_1022,N_976);
nand U1109 (N_1109,N_994,N_1041);
or U1110 (N_1110,N_1030,N_1019);
nand U1111 (N_1111,N_1036,N_1048);
and U1112 (N_1112,N_987,N_1038);
or U1113 (N_1113,N_984,N_1013);
nand U1114 (N_1114,N_978,N_1016);
nor U1115 (N_1115,N_988,N_1002);
nand U1116 (N_1116,N_1032,N_978);
and U1117 (N_1117,N_983,N_996);
and U1118 (N_1118,N_1019,N_1039);
and U1119 (N_1119,N_1027,N_1010);
nor U1120 (N_1120,N_1040,N_1001);
or U1121 (N_1121,N_1004,N_1041);
and U1122 (N_1122,N_1023,N_1048);
and U1123 (N_1123,N_1014,N_1038);
nor U1124 (N_1124,N_1010,N_982);
or U1125 (N_1125,N_1051,N_1110);
and U1126 (N_1126,N_1058,N_1066);
nand U1127 (N_1127,N_1061,N_1095);
and U1128 (N_1128,N_1121,N_1106);
nor U1129 (N_1129,N_1077,N_1074);
and U1130 (N_1130,N_1099,N_1072);
or U1131 (N_1131,N_1113,N_1069);
nor U1132 (N_1132,N_1089,N_1083);
nand U1133 (N_1133,N_1091,N_1096);
or U1134 (N_1134,N_1092,N_1067);
nand U1135 (N_1135,N_1122,N_1116);
nand U1136 (N_1136,N_1050,N_1123);
and U1137 (N_1137,N_1117,N_1101);
and U1138 (N_1138,N_1068,N_1087);
nand U1139 (N_1139,N_1107,N_1120);
or U1140 (N_1140,N_1098,N_1063);
nand U1141 (N_1141,N_1052,N_1119);
nand U1142 (N_1142,N_1103,N_1080);
nor U1143 (N_1143,N_1108,N_1111);
nand U1144 (N_1144,N_1073,N_1093);
and U1145 (N_1145,N_1124,N_1082);
and U1146 (N_1146,N_1088,N_1085);
nand U1147 (N_1147,N_1059,N_1097);
nand U1148 (N_1148,N_1109,N_1064);
nor U1149 (N_1149,N_1081,N_1086);
nor U1150 (N_1150,N_1054,N_1078);
nand U1151 (N_1151,N_1065,N_1115);
or U1152 (N_1152,N_1084,N_1094);
nand U1153 (N_1153,N_1076,N_1060);
nor U1154 (N_1154,N_1102,N_1112);
and U1155 (N_1155,N_1079,N_1062);
and U1156 (N_1156,N_1057,N_1075);
nor U1157 (N_1157,N_1056,N_1104);
nor U1158 (N_1158,N_1100,N_1118);
nand U1159 (N_1159,N_1114,N_1055);
nand U1160 (N_1160,N_1071,N_1070);
or U1161 (N_1161,N_1090,N_1053);
nor U1162 (N_1162,N_1105,N_1113);
nor U1163 (N_1163,N_1061,N_1057);
and U1164 (N_1164,N_1096,N_1123);
nand U1165 (N_1165,N_1063,N_1124);
and U1166 (N_1166,N_1115,N_1110);
xor U1167 (N_1167,N_1107,N_1105);
nor U1168 (N_1168,N_1071,N_1107);
and U1169 (N_1169,N_1102,N_1110);
nor U1170 (N_1170,N_1075,N_1067);
or U1171 (N_1171,N_1055,N_1092);
or U1172 (N_1172,N_1093,N_1090);
and U1173 (N_1173,N_1116,N_1057);
or U1174 (N_1174,N_1089,N_1061);
nand U1175 (N_1175,N_1119,N_1108);
nand U1176 (N_1176,N_1071,N_1093);
nor U1177 (N_1177,N_1121,N_1061);
nand U1178 (N_1178,N_1066,N_1104);
or U1179 (N_1179,N_1070,N_1083);
nor U1180 (N_1180,N_1115,N_1108);
nand U1181 (N_1181,N_1070,N_1102);
or U1182 (N_1182,N_1070,N_1062);
nor U1183 (N_1183,N_1066,N_1080);
or U1184 (N_1184,N_1065,N_1068);
nand U1185 (N_1185,N_1117,N_1116);
and U1186 (N_1186,N_1108,N_1086);
or U1187 (N_1187,N_1105,N_1078);
nor U1188 (N_1188,N_1115,N_1070);
or U1189 (N_1189,N_1061,N_1100);
nor U1190 (N_1190,N_1073,N_1086);
or U1191 (N_1191,N_1106,N_1122);
or U1192 (N_1192,N_1069,N_1117);
nand U1193 (N_1193,N_1069,N_1092);
nor U1194 (N_1194,N_1058,N_1102);
nand U1195 (N_1195,N_1102,N_1081);
or U1196 (N_1196,N_1070,N_1080);
and U1197 (N_1197,N_1119,N_1053);
or U1198 (N_1198,N_1086,N_1075);
xor U1199 (N_1199,N_1084,N_1112);
and U1200 (N_1200,N_1142,N_1172);
nor U1201 (N_1201,N_1189,N_1145);
nand U1202 (N_1202,N_1182,N_1132);
nand U1203 (N_1203,N_1148,N_1152);
nor U1204 (N_1204,N_1141,N_1192);
xnor U1205 (N_1205,N_1193,N_1157);
nor U1206 (N_1206,N_1188,N_1197);
nor U1207 (N_1207,N_1147,N_1128);
and U1208 (N_1208,N_1176,N_1175);
and U1209 (N_1209,N_1156,N_1130);
nor U1210 (N_1210,N_1137,N_1166);
nand U1211 (N_1211,N_1131,N_1127);
nor U1212 (N_1212,N_1174,N_1150);
nand U1213 (N_1213,N_1134,N_1160);
or U1214 (N_1214,N_1144,N_1164);
nor U1215 (N_1215,N_1183,N_1143);
or U1216 (N_1216,N_1159,N_1195);
nor U1217 (N_1217,N_1185,N_1161);
or U1218 (N_1218,N_1139,N_1154);
nor U1219 (N_1219,N_1129,N_1177);
nand U1220 (N_1220,N_1196,N_1151);
xor U1221 (N_1221,N_1199,N_1167);
nor U1222 (N_1222,N_1126,N_1179);
and U1223 (N_1223,N_1125,N_1135);
nand U1224 (N_1224,N_1186,N_1165);
and U1225 (N_1225,N_1173,N_1158);
nor U1226 (N_1226,N_1184,N_1168);
or U1227 (N_1227,N_1171,N_1198);
or U1228 (N_1228,N_1191,N_1149);
or U1229 (N_1229,N_1140,N_1153);
nor U1230 (N_1230,N_1178,N_1138);
nor U1231 (N_1231,N_1180,N_1136);
nand U1232 (N_1232,N_1169,N_1155);
nand U1233 (N_1233,N_1133,N_1163);
or U1234 (N_1234,N_1181,N_1170);
and U1235 (N_1235,N_1162,N_1187);
nor U1236 (N_1236,N_1146,N_1194);
and U1237 (N_1237,N_1190,N_1163);
nor U1238 (N_1238,N_1145,N_1180);
or U1239 (N_1239,N_1188,N_1148);
or U1240 (N_1240,N_1169,N_1189);
nand U1241 (N_1241,N_1153,N_1170);
nand U1242 (N_1242,N_1176,N_1162);
and U1243 (N_1243,N_1175,N_1156);
nand U1244 (N_1244,N_1194,N_1142);
and U1245 (N_1245,N_1176,N_1166);
or U1246 (N_1246,N_1163,N_1146);
nand U1247 (N_1247,N_1139,N_1189);
nor U1248 (N_1248,N_1198,N_1156);
and U1249 (N_1249,N_1132,N_1130);
nand U1250 (N_1250,N_1125,N_1158);
nand U1251 (N_1251,N_1127,N_1135);
or U1252 (N_1252,N_1187,N_1197);
nor U1253 (N_1253,N_1189,N_1131);
and U1254 (N_1254,N_1149,N_1180);
nor U1255 (N_1255,N_1153,N_1172);
and U1256 (N_1256,N_1167,N_1188);
nor U1257 (N_1257,N_1149,N_1179);
nand U1258 (N_1258,N_1133,N_1187);
nor U1259 (N_1259,N_1159,N_1146);
nor U1260 (N_1260,N_1177,N_1152);
and U1261 (N_1261,N_1196,N_1187);
nor U1262 (N_1262,N_1158,N_1156);
nor U1263 (N_1263,N_1185,N_1168);
nand U1264 (N_1264,N_1140,N_1166);
and U1265 (N_1265,N_1176,N_1141);
or U1266 (N_1266,N_1179,N_1164);
nand U1267 (N_1267,N_1128,N_1185);
or U1268 (N_1268,N_1183,N_1139);
and U1269 (N_1269,N_1186,N_1177);
nand U1270 (N_1270,N_1180,N_1133);
and U1271 (N_1271,N_1166,N_1199);
and U1272 (N_1272,N_1159,N_1175);
nand U1273 (N_1273,N_1183,N_1194);
nor U1274 (N_1274,N_1176,N_1179);
or U1275 (N_1275,N_1243,N_1200);
nand U1276 (N_1276,N_1231,N_1260);
or U1277 (N_1277,N_1255,N_1238);
or U1278 (N_1278,N_1268,N_1215);
nor U1279 (N_1279,N_1206,N_1240);
nor U1280 (N_1280,N_1258,N_1235);
nand U1281 (N_1281,N_1214,N_1265);
or U1282 (N_1282,N_1213,N_1241);
nand U1283 (N_1283,N_1236,N_1229);
and U1284 (N_1284,N_1226,N_1266);
nand U1285 (N_1285,N_1228,N_1224);
nor U1286 (N_1286,N_1273,N_1251);
or U1287 (N_1287,N_1217,N_1267);
nor U1288 (N_1288,N_1244,N_1252);
or U1289 (N_1289,N_1203,N_1254);
and U1290 (N_1290,N_1239,N_1256);
nand U1291 (N_1291,N_1233,N_1219);
nor U1292 (N_1292,N_1234,N_1253);
and U1293 (N_1293,N_1250,N_1246);
or U1294 (N_1294,N_1222,N_1225);
nand U1295 (N_1295,N_1216,N_1212);
nand U1296 (N_1296,N_1259,N_1209);
nand U1297 (N_1297,N_1271,N_1261);
nor U1298 (N_1298,N_1272,N_1274);
nor U1299 (N_1299,N_1264,N_1202);
nand U1300 (N_1300,N_1221,N_1257);
nand U1301 (N_1301,N_1249,N_1205);
and U1302 (N_1302,N_1227,N_1248);
or U1303 (N_1303,N_1230,N_1262);
nor U1304 (N_1304,N_1245,N_1208);
nand U1305 (N_1305,N_1201,N_1210);
nand U1306 (N_1306,N_1232,N_1218);
or U1307 (N_1307,N_1207,N_1270);
nand U1308 (N_1308,N_1242,N_1269);
nor U1309 (N_1309,N_1211,N_1220);
nor U1310 (N_1310,N_1263,N_1237);
or U1311 (N_1311,N_1204,N_1247);
nor U1312 (N_1312,N_1223,N_1204);
nor U1313 (N_1313,N_1253,N_1225);
nand U1314 (N_1314,N_1230,N_1222);
nor U1315 (N_1315,N_1256,N_1242);
and U1316 (N_1316,N_1217,N_1262);
nor U1317 (N_1317,N_1268,N_1208);
and U1318 (N_1318,N_1227,N_1214);
or U1319 (N_1319,N_1257,N_1247);
and U1320 (N_1320,N_1265,N_1241);
nor U1321 (N_1321,N_1260,N_1218);
nand U1322 (N_1322,N_1242,N_1270);
nand U1323 (N_1323,N_1244,N_1210);
or U1324 (N_1324,N_1241,N_1260);
or U1325 (N_1325,N_1229,N_1224);
and U1326 (N_1326,N_1273,N_1205);
and U1327 (N_1327,N_1202,N_1224);
and U1328 (N_1328,N_1242,N_1218);
or U1329 (N_1329,N_1210,N_1234);
nand U1330 (N_1330,N_1236,N_1201);
xor U1331 (N_1331,N_1222,N_1266);
and U1332 (N_1332,N_1226,N_1263);
nand U1333 (N_1333,N_1234,N_1211);
and U1334 (N_1334,N_1237,N_1262);
or U1335 (N_1335,N_1237,N_1214);
nand U1336 (N_1336,N_1204,N_1267);
nor U1337 (N_1337,N_1271,N_1238);
nor U1338 (N_1338,N_1220,N_1274);
nand U1339 (N_1339,N_1272,N_1256);
or U1340 (N_1340,N_1227,N_1225);
nor U1341 (N_1341,N_1227,N_1250);
and U1342 (N_1342,N_1248,N_1212);
nand U1343 (N_1343,N_1250,N_1262);
or U1344 (N_1344,N_1268,N_1245);
and U1345 (N_1345,N_1208,N_1234);
nand U1346 (N_1346,N_1204,N_1225);
nor U1347 (N_1347,N_1241,N_1263);
or U1348 (N_1348,N_1241,N_1259);
and U1349 (N_1349,N_1224,N_1246);
nand U1350 (N_1350,N_1333,N_1345);
nand U1351 (N_1351,N_1294,N_1306);
nor U1352 (N_1352,N_1296,N_1338);
nor U1353 (N_1353,N_1320,N_1291);
nor U1354 (N_1354,N_1322,N_1290);
nor U1355 (N_1355,N_1330,N_1295);
nand U1356 (N_1356,N_1276,N_1334);
nand U1357 (N_1357,N_1340,N_1308);
and U1358 (N_1358,N_1283,N_1310);
xor U1359 (N_1359,N_1277,N_1280);
and U1360 (N_1360,N_1282,N_1325);
and U1361 (N_1361,N_1285,N_1304);
nor U1362 (N_1362,N_1300,N_1297);
and U1363 (N_1363,N_1286,N_1289);
nand U1364 (N_1364,N_1301,N_1298);
nand U1365 (N_1365,N_1323,N_1341);
nand U1366 (N_1366,N_1312,N_1339);
and U1367 (N_1367,N_1321,N_1302);
nor U1368 (N_1368,N_1342,N_1311);
nor U1369 (N_1369,N_1349,N_1305);
nand U1370 (N_1370,N_1299,N_1292);
and U1371 (N_1371,N_1288,N_1337);
and U1372 (N_1372,N_1275,N_1328);
or U1373 (N_1373,N_1324,N_1316);
nor U1374 (N_1374,N_1348,N_1278);
and U1375 (N_1375,N_1293,N_1326);
nand U1376 (N_1376,N_1346,N_1307);
nor U1377 (N_1377,N_1303,N_1347);
nor U1378 (N_1378,N_1318,N_1313);
or U1379 (N_1379,N_1287,N_1343);
and U1380 (N_1380,N_1331,N_1336);
or U1381 (N_1381,N_1281,N_1314);
or U1382 (N_1382,N_1344,N_1315);
or U1383 (N_1383,N_1327,N_1317);
nor U1384 (N_1384,N_1319,N_1329);
or U1385 (N_1385,N_1284,N_1335);
and U1386 (N_1386,N_1309,N_1332);
nand U1387 (N_1387,N_1279,N_1343);
nor U1388 (N_1388,N_1285,N_1322);
nor U1389 (N_1389,N_1300,N_1284);
and U1390 (N_1390,N_1299,N_1284);
xnor U1391 (N_1391,N_1342,N_1285);
or U1392 (N_1392,N_1278,N_1283);
nand U1393 (N_1393,N_1344,N_1296);
and U1394 (N_1394,N_1325,N_1291);
and U1395 (N_1395,N_1321,N_1292);
nand U1396 (N_1396,N_1313,N_1317);
or U1397 (N_1397,N_1293,N_1328);
or U1398 (N_1398,N_1291,N_1345);
and U1399 (N_1399,N_1325,N_1324);
and U1400 (N_1400,N_1300,N_1295);
nor U1401 (N_1401,N_1280,N_1279);
or U1402 (N_1402,N_1322,N_1333);
nand U1403 (N_1403,N_1282,N_1308);
nor U1404 (N_1404,N_1292,N_1328);
and U1405 (N_1405,N_1281,N_1300);
nand U1406 (N_1406,N_1298,N_1338);
nand U1407 (N_1407,N_1299,N_1311);
and U1408 (N_1408,N_1336,N_1322);
xor U1409 (N_1409,N_1302,N_1326);
or U1410 (N_1410,N_1321,N_1285);
and U1411 (N_1411,N_1339,N_1307);
or U1412 (N_1412,N_1295,N_1340);
and U1413 (N_1413,N_1279,N_1292);
nand U1414 (N_1414,N_1288,N_1344);
and U1415 (N_1415,N_1341,N_1284);
nor U1416 (N_1416,N_1341,N_1292);
or U1417 (N_1417,N_1319,N_1322);
nor U1418 (N_1418,N_1304,N_1283);
and U1419 (N_1419,N_1283,N_1333);
nor U1420 (N_1420,N_1290,N_1282);
or U1421 (N_1421,N_1282,N_1275);
or U1422 (N_1422,N_1296,N_1341);
or U1423 (N_1423,N_1308,N_1304);
and U1424 (N_1424,N_1332,N_1334);
and U1425 (N_1425,N_1400,N_1416);
nand U1426 (N_1426,N_1410,N_1378);
nor U1427 (N_1427,N_1395,N_1380);
nor U1428 (N_1428,N_1379,N_1352);
nor U1429 (N_1429,N_1375,N_1356);
or U1430 (N_1430,N_1364,N_1363);
nor U1431 (N_1431,N_1376,N_1422);
nand U1432 (N_1432,N_1412,N_1411);
and U1433 (N_1433,N_1396,N_1360);
nor U1434 (N_1434,N_1406,N_1358);
and U1435 (N_1435,N_1385,N_1369);
or U1436 (N_1436,N_1414,N_1405);
or U1437 (N_1437,N_1393,N_1382);
nor U1438 (N_1438,N_1417,N_1354);
or U1439 (N_1439,N_1399,N_1387);
and U1440 (N_1440,N_1374,N_1370);
and U1441 (N_1441,N_1418,N_1389);
nand U1442 (N_1442,N_1361,N_1359);
nand U1443 (N_1443,N_1423,N_1408);
and U1444 (N_1444,N_1386,N_1365);
and U1445 (N_1445,N_1401,N_1353);
and U1446 (N_1446,N_1397,N_1413);
nand U1447 (N_1447,N_1381,N_1351);
or U1448 (N_1448,N_1350,N_1372);
nor U1449 (N_1449,N_1366,N_1420);
and U1450 (N_1450,N_1415,N_1394);
nand U1451 (N_1451,N_1419,N_1404);
nand U1452 (N_1452,N_1362,N_1371);
nand U1453 (N_1453,N_1390,N_1355);
or U1454 (N_1454,N_1398,N_1368);
or U1455 (N_1455,N_1383,N_1409);
and U1456 (N_1456,N_1421,N_1373);
nor U1457 (N_1457,N_1424,N_1392);
nor U1458 (N_1458,N_1384,N_1407);
or U1459 (N_1459,N_1388,N_1391);
and U1460 (N_1460,N_1377,N_1403);
and U1461 (N_1461,N_1402,N_1357);
nand U1462 (N_1462,N_1367,N_1374);
nand U1463 (N_1463,N_1363,N_1389);
and U1464 (N_1464,N_1383,N_1398);
nor U1465 (N_1465,N_1404,N_1360);
and U1466 (N_1466,N_1411,N_1354);
nand U1467 (N_1467,N_1423,N_1359);
nand U1468 (N_1468,N_1359,N_1365);
nand U1469 (N_1469,N_1369,N_1381);
nor U1470 (N_1470,N_1383,N_1394);
or U1471 (N_1471,N_1377,N_1416);
nor U1472 (N_1472,N_1416,N_1405);
and U1473 (N_1473,N_1360,N_1381);
nand U1474 (N_1474,N_1380,N_1412);
or U1475 (N_1475,N_1414,N_1424);
or U1476 (N_1476,N_1372,N_1412);
and U1477 (N_1477,N_1381,N_1392);
nor U1478 (N_1478,N_1422,N_1407);
nand U1479 (N_1479,N_1420,N_1362);
nand U1480 (N_1480,N_1370,N_1378);
or U1481 (N_1481,N_1389,N_1424);
nor U1482 (N_1482,N_1397,N_1420);
nor U1483 (N_1483,N_1404,N_1374);
or U1484 (N_1484,N_1385,N_1371);
or U1485 (N_1485,N_1357,N_1415);
nor U1486 (N_1486,N_1413,N_1374);
or U1487 (N_1487,N_1396,N_1401);
nor U1488 (N_1488,N_1361,N_1362);
nor U1489 (N_1489,N_1405,N_1413);
nor U1490 (N_1490,N_1353,N_1402);
nand U1491 (N_1491,N_1357,N_1384);
and U1492 (N_1492,N_1356,N_1365);
nand U1493 (N_1493,N_1401,N_1366);
nor U1494 (N_1494,N_1422,N_1409);
nor U1495 (N_1495,N_1377,N_1396);
and U1496 (N_1496,N_1404,N_1351);
or U1497 (N_1497,N_1363,N_1422);
nand U1498 (N_1498,N_1390,N_1405);
and U1499 (N_1499,N_1408,N_1417);
and U1500 (N_1500,N_1478,N_1495);
nand U1501 (N_1501,N_1477,N_1483);
or U1502 (N_1502,N_1429,N_1468);
nor U1503 (N_1503,N_1428,N_1498);
nor U1504 (N_1504,N_1458,N_1455);
nand U1505 (N_1505,N_1472,N_1432);
nor U1506 (N_1506,N_1492,N_1475);
nand U1507 (N_1507,N_1491,N_1447);
nand U1508 (N_1508,N_1466,N_1481);
and U1509 (N_1509,N_1449,N_1462);
or U1510 (N_1510,N_1437,N_1494);
and U1511 (N_1511,N_1488,N_1427);
nor U1512 (N_1512,N_1496,N_1460);
and U1513 (N_1513,N_1434,N_1470);
nand U1514 (N_1514,N_1440,N_1441);
or U1515 (N_1515,N_1451,N_1474);
xnor U1516 (N_1516,N_1499,N_1467);
and U1517 (N_1517,N_1425,N_1497);
nand U1518 (N_1518,N_1476,N_1464);
or U1519 (N_1519,N_1446,N_1487);
nand U1520 (N_1520,N_1473,N_1431);
nand U1521 (N_1521,N_1484,N_1426);
nor U1522 (N_1522,N_1435,N_1438);
or U1523 (N_1523,N_1448,N_1457);
and U1524 (N_1524,N_1450,N_1456);
or U1525 (N_1525,N_1444,N_1442);
nand U1526 (N_1526,N_1454,N_1461);
and U1527 (N_1527,N_1443,N_1433);
nand U1528 (N_1528,N_1493,N_1482);
or U1529 (N_1529,N_1480,N_1489);
nor U1530 (N_1530,N_1439,N_1490);
nand U1531 (N_1531,N_1445,N_1452);
nand U1532 (N_1532,N_1430,N_1469);
nand U1533 (N_1533,N_1453,N_1459);
nor U1534 (N_1534,N_1436,N_1463);
nor U1535 (N_1535,N_1479,N_1465);
or U1536 (N_1536,N_1486,N_1471);
nand U1537 (N_1537,N_1485,N_1469);
nand U1538 (N_1538,N_1498,N_1487);
xor U1539 (N_1539,N_1483,N_1488);
nand U1540 (N_1540,N_1476,N_1478);
or U1541 (N_1541,N_1495,N_1490);
nand U1542 (N_1542,N_1432,N_1431);
or U1543 (N_1543,N_1466,N_1472);
nand U1544 (N_1544,N_1462,N_1479);
nor U1545 (N_1545,N_1435,N_1460);
xor U1546 (N_1546,N_1453,N_1475);
or U1547 (N_1547,N_1476,N_1456);
and U1548 (N_1548,N_1428,N_1427);
nand U1549 (N_1549,N_1436,N_1484);
nor U1550 (N_1550,N_1488,N_1490);
or U1551 (N_1551,N_1463,N_1484);
nor U1552 (N_1552,N_1469,N_1470);
nand U1553 (N_1553,N_1453,N_1434);
nor U1554 (N_1554,N_1428,N_1442);
nor U1555 (N_1555,N_1474,N_1489);
or U1556 (N_1556,N_1498,N_1488);
nand U1557 (N_1557,N_1480,N_1450);
or U1558 (N_1558,N_1467,N_1498);
and U1559 (N_1559,N_1429,N_1434);
xor U1560 (N_1560,N_1427,N_1498);
xnor U1561 (N_1561,N_1464,N_1463);
nor U1562 (N_1562,N_1489,N_1488);
and U1563 (N_1563,N_1443,N_1489);
xor U1564 (N_1564,N_1469,N_1461);
nand U1565 (N_1565,N_1475,N_1497);
xor U1566 (N_1566,N_1446,N_1475);
nand U1567 (N_1567,N_1465,N_1489);
nor U1568 (N_1568,N_1478,N_1488);
nor U1569 (N_1569,N_1468,N_1460);
or U1570 (N_1570,N_1448,N_1481);
nand U1571 (N_1571,N_1433,N_1446);
and U1572 (N_1572,N_1448,N_1434);
or U1573 (N_1573,N_1437,N_1454);
nor U1574 (N_1574,N_1470,N_1438);
and U1575 (N_1575,N_1546,N_1565);
nand U1576 (N_1576,N_1545,N_1503);
nand U1577 (N_1577,N_1517,N_1547);
or U1578 (N_1578,N_1534,N_1539);
nor U1579 (N_1579,N_1552,N_1523);
nor U1580 (N_1580,N_1569,N_1532);
nand U1581 (N_1581,N_1518,N_1562);
or U1582 (N_1582,N_1504,N_1537);
nand U1583 (N_1583,N_1556,N_1522);
or U1584 (N_1584,N_1528,N_1543);
nand U1585 (N_1585,N_1527,N_1501);
nor U1586 (N_1586,N_1554,N_1553);
or U1587 (N_1587,N_1510,N_1561);
nand U1588 (N_1588,N_1519,N_1557);
or U1589 (N_1589,N_1516,N_1506);
and U1590 (N_1590,N_1511,N_1540);
or U1591 (N_1591,N_1558,N_1533);
and U1592 (N_1592,N_1573,N_1568);
xor U1593 (N_1593,N_1515,N_1574);
nor U1594 (N_1594,N_1551,N_1529);
nor U1595 (N_1595,N_1542,N_1500);
or U1596 (N_1596,N_1513,N_1567);
or U1597 (N_1597,N_1555,N_1536);
nor U1598 (N_1598,N_1525,N_1559);
and U1599 (N_1599,N_1566,N_1524);
nand U1600 (N_1600,N_1549,N_1544);
and U1601 (N_1601,N_1571,N_1531);
nor U1602 (N_1602,N_1538,N_1563);
xor U1603 (N_1603,N_1530,N_1560);
nor U1604 (N_1604,N_1502,N_1564);
nor U1605 (N_1605,N_1508,N_1521);
nand U1606 (N_1606,N_1541,N_1509);
nand U1607 (N_1607,N_1572,N_1514);
nor U1608 (N_1608,N_1570,N_1548);
or U1609 (N_1609,N_1507,N_1512);
or U1610 (N_1610,N_1535,N_1520);
or U1611 (N_1611,N_1505,N_1550);
nor U1612 (N_1612,N_1526,N_1513);
nand U1613 (N_1613,N_1566,N_1565);
or U1614 (N_1614,N_1505,N_1525);
and U1615 (N_1615,N_1523,N_1505);
or U1616 (N_1616,N_1501,N_1522);
or U1617 (N_1617,N_1503,N_1565);
and U1618 (N_1618,N_1560,N_1526);
nor U1619 (N_1619,N_1520,N_1573);
and U1620 (N_1620,N_1548,N_1542);
nor U1621 (N_1621,N_1527,N_1512);
and U1622 (N_1622,N_1525,N_1551);
nor U1623 (N_1623,N_1530,N_1564);
nand U1624 (N_1624,N_1560,N_1502);
nor U1625 (N_1625,N_1573,N_1560);
or U1626 (N_1626,N_1508,N_1529);
nor U1627 (N_1627,N_1508,N_1545);
or U1628 (N_1628,N_1531,N_1570);
xor U1629 (N_1629,N_1570,N_1555);
nand U1630 (N_1630,N_1503,N_1548);
nor U1631 (N_1631,N_1500,N_1515);
nor U1632 (N_1632,N_1508,N_1503);
nor U1633 (N_1633,N_1509,N_1531);
nor U1634 (N_1634,N_1560,N_1554);
nor U1635 (N_1635,N_1565,N_1548);
nand U1636 (N_1636,N_1569,N_1528);
nor U1637 (N_1637,N_1505,N_1503);
or U1638 (N_1638,N_1572,N_1506);
or U1639 (N_1639,N_1538,N_1546);
or U1640 (N_1640,N_1511,N_1568);
nand U1641 (N_1641,N_1519,N_1559);
or U1642 (N_1642,N_1523,N_1509);
nand U1643 (N_1643,N_1525,N_1508);
nand U1644 (N_1644,N_1564,N_1528);
or U1645 (N_1645,N_1528,N_1538);
or U1646 (N_1646,N_1544,N_1536);
nand U1647 (N_1647,N_1547,N_1527);
nor U1648 (N_1648,N_1536,N_1552);
and U1649 (N_1649,N_1572,N_1543);
nand U1650 (N_1650,N_1630,N_1639);
nor U1651 (N_1651,N_1599,N_1601);
and U1652 (N_1652,N_1642,N_1605);
or U1653 (N_1653,N_1583,N_1640);
nand U1654 (N_1654,N_1612,N_1575);
nor U1655 (N_1655,N_1609,N_1577);
or U1656 (N_1656,N_1649,N_1603);
nor U1657 (N_1657,N_1607,N_1625);
nand U1658 (N_1658,N_1615,N_1611);
nor U1659 (N_1659,N_1624,N_1602);
and U1660 (N_1660,N_1618,N_1638);
and U1661 (N_1661,N_1629,N_1585);
nand U1662 (N_1662,N_1597,N_1644);
or U1663 (N_1663,N_1645,N_1576);
or U1664 (N_1664,N_1634,N_1584);
nand U1665 (N_1665,N_1620,N_1579);
and U1666 (N_1666,N_1635,N_1595);
nor U1667 (N_1667,N_1580,N_1633);
and U1668 (N_1668,N_1582,N_1592);
nor U1669 (N_1669,N_1621,N_1648);
xor U1670 (N_1670,N_1610,N_1578);
xor U1671 (N_1671,N_1628,N_1591);
and U1672 (N_1672,N_1623,N_1619);
and U1673 (N_1673,N_1616,N_1608);
or U1674 (N_1674,N_1631,N_1594);
or U1675 (N_1675,N_1636,N_1598);
and U1676 (N_1676,N_1600,N_1588);
and U1677 (N_1677,N_1626,N_1614);
nor U1678 (N_1678,N_1637,N_1646);
nor U1679 (N_1679,N_1617,N_1593);
nand U1680 (N_1680,N_1643,N_1632);
and U1681 (N_1681,N_1622,N_1613);
nor U1682 (N_1682,N_1641,N_1586);
and U1683 (N_1683,N_1596,N_1606);
nand U1684 (N_1684,N_1581,N_1590);
nor U1685 (N_1685,N_1647,N_1587);
nand U1686 (N_1686,N_1589,N_1604);
or U1687 (N_1687,N_1627,N_1590);
or U1688 (N_1688,N_1618,N_1593);
nand U1689 (N_1689,N_1620,N_1632);
and U1690 (N_1690,N_1597,N_1583);
and U1691 (N_1691,N_1615,N_1605);
nand U1692 (N_1692,N_1613,N_1641);
and U1693 (N_1693,N_1648,N_1624);
nand U1694 (N_1694,N_1629,N_1604);
or U1695 (N_1695,N_1585,N_1622);
and U1696 (N_1696,N_1584,N_1616);
nor U1697 (N_1697,N_1622,N_1628);
and U1698 (N_1698,N_1649,N_1582);
and U1699 (N_1699,N_1625,N_1602);
or U1700 (N_1700,N_1638,N_1617);
nand U1701 (N_1701,N_1613,N_1603);
and U1702 (N_1702,N_1608,N_1612);
or U1703 (N_1703,N_1579,N_1637);
nor U1704 (N_1704,N_1584,N_1612);
and U1705 (N_1705,N_1584,N_1635);
nor U1706 (N_1706,N_1643,N_1596);
nor U1707 (N_1707,N_1610,N_1616);
or U1708 (N_1708,N_1609,N_1627);
nor U1709 (N_1709,N_1628,N_1583);
nand U1710 (N_1710,N_1595,N_1649);
and U1711 (N_1711,N_1604,N_1645);
xor U1712 (N_1712,N_1589,N_1625);
or U1713 (N_1713,N_1585,N_1597);
and U1714 (N_1714,N_1597,N_1582);
or U1715 (N_1715,N_1588,N_1609);
and U1716 (N_1716,N_1614,N_1589);
nand U1717 (N_1717,N_1600,N_1613);
or U1718 (N_1718,N_1633,N_1643);
and U1719 (N_1719,N_1643,N_1644);
or U1720 (N_1720,N_1606,N_1639);
nor U1721 (N_1721,N_1585,N_1615);
or U1722 (N_1722,N_1606,N_1611);
and U1723 (N_1723,N_1604,N_1623);
and U1724 (N_1724,N_1595,N_1627);
or U1725 (N_1725,N_1673,N_1654);
nor U1726 (N_1726,N_1686,N_1666);
nor U1727 (N_1727,N_1714,N_1667);
nand U1728 (N_1728,N_1695,N_1652);
and U1729 (N_1729,N_1669,N_1684);
nand U1730 (N_1730,N_1718,N_1671);
and U1731 (N_1731,N_1685,N_1700);
or U1732 (N_1732,N_1721,N_1705);
nand U1733 (N_1733,N_1678,N_1663);
and U1734 (N_1734,N_1687,N_1655);
nor U1735 (N_1735,N_1699,N_1690);
nand U1736 (N_1736,N_1722,N_1676);
or U1737 (N_1737,N_1697,N_1650);
and U1738 (N_1738,N_1657,N_1717);
nor U1739 (N_1739,N_1683,N_1694);
and U1740 (N_1740,N_1706,N_1720);
or U1741 (N_1741,N_1689,N_1653);
nor U1742 (N_1742,N_1716,N_1675);
or U1743 (N_1743,N_1682,N_1713);
and U1744 (N_1744,N_1708,N_1668);
nand U1745 (N_1745,N_1692,N_1707);
nor U1746 (N_1746,N_1701,N_1672);
nand U1747 (N_1747,N_1711,N_1680);
nand U1748 (N_1748,N_1677,N_1661);
and U1749 (N_1749,N_1664,N_1709);
nor U1750 (N_1750,N_1704,N_1693);
and U1751 (N_1751,N_1703,N_1719);
or U1752 (N_1752,N_1665,N_1715);
and U1753 (N_1753,N_1712,N_1656);
or U1754 (N_1754,N_1681,N_1688);
nand U1755 (N_1755,N_1696,N_1710);
and U1756 (N_1756,N_1724,N_1662);
nand U1757 (N_1757,N_1659,N_1698);
nand U1758 (N_1758,N_1658,N_1674);
nor U1759 (N_1759,N_1670,N_1723);
nor U1760 (N_1760,N_1660,N_1702);
or U1761 (N_1761,N_1691,N_1651);
and U1762 (N_1762,N_1679,N_1661);
or U1763 (N_1763,N_1657,N_1718);
and U1764 (N_1764,N_1685,N_1683);
and U1765 (N_1765,N_1724,N_1715);
and U1766 (N_1766,N_1650,N_1719);
nand U1767 (N_1767,N_1713,N_1691);
nand U1768 (N_1768,N_1657,N_1719);
and U1769 (N_1769,N_1686,N_1716);
nor U1770 (N_1770,N_1717,N_1703);
nand U1771 (N_1771,N_1664,N_1670);
and U1772 (N_1772,N_1702,N_1681);
and U1773 (N_1773,N_1691,N_1701);
and U1774 (N_1774,N_1713,N_1683);
and U1775 (N_1775,N_1671,N_1691);
nand U1776 (N_1776,N_1650,N_1720);
or U1777 (N_1777,N_1689,N_1664);
or U1778 (N_1778,N_1669,N_1661);
and U1779 (N_1779,N_1724,N_1679);
nor U1780 (N_1780,N_1659,N_1662);
or U1781 (N_1781,N_1668,N_1698);
nand U1782 (N_1782,N_1662,N_1702);
and U1783 (N_1783,N_1703,N_1673);
and U1784 (N_1784,N_1689,N_1685);
nor U1785 (N_1785,N_1653,N_1698);
or U1786 (N_1786,N_1710,N_1700);
and U1787 (N_1787,N_1677,N_1719);
nor U1788 (N_1788,N_1655,N_1659);
and U1789 (N_1789,N_1686,N_1652);
nor U1790 (N_1790,N_1711,N_1703);
nand U1791 (N_1791,N_1651,N_1710);
nor U1792 (N_1792,N_1705,N_1672);
nand U1793 (N_1793,N_1723,N_1671);
nand U1794 (N_1794,N_1654,N_1704);
nand U1795 (N_1795,N_1656,N_1709);
and U1796 (N_1796,N_1715,N_1666);
or U1797 (N_1797,N_1716,N_1723);
and U1798 (N_1798,N_1663,N_1691);
nand U1799 (N_1799,N_1713,N_1653);
nand U1800 (N_1800,N_1759,N_1788);
and U1801 (N_1801,N_1779,N_1781);
nand U1802 (N_1802,N_1732,N_1742);
or U1803 (N_1803,N_1750,N_1763);
and U1804 (N_1804,N_1741,N_1725);
or U1805 (N_1805,N_1765,N_1733);
or U1806 (N_1806,N_1757,N_1787);
nand U1807 (N_1807,N_1775,N_1736);
nor U1808 (N_1808,N_1768,N_1743);
nor U1809 (N_1809,N_1762,N_1761);
or U1810 (N_1810,N_1778,N_1734);
nand U1811 (N_1811,N_1752,N_1758);
nor U1812 (N_1812,N_1793,N_1740);
xor U1813 (N_1813,N_1731,N_1749);
and U1814 (N_1814,N_1794,N_1789);
nand U1815 (N_1815,N_1767,N_1770);
or U1816 (N_1816,N_1774,N_1756);
nor U1817 (N_1817,N_1782,N_1769);
nor U1818 (N_1818,N_1755,N_1783);
nor U1819 (N_1819,N_1760,N_1790);
or U1820 (N_1820,N_1748,N_1791);
and U1821 (N_1821,N_1729,N_1766);
nand U1822 (N_1822,N_1728,N_1726);
xnor U1823 (N_1823,N_1746,N_1727);
and U1824 (N_1824,N_1777,N_1796);
or U1825 (N_1825,N_1730,N_1797);
nor U1826 (N_1826,N_1776,N_1771);
nor U1827 (N_1827,N_1780,N_1798);
or U1828 (N_1828,N_1744,N_1772);
nand U1829 (N_1829,N_1751,N_1735);
and U1830 (N_1830,N_1792,N_1799);
nor U1831 (N_1831,N_1764,N_1786);
nor U1832 (N_1832,N_1739,N_1747);
nand U1833 (N_1833,N_1737,N_1753);
nor U1834 (N_1834,N_1784,N_1745);
or U1835 (N_1835,N_1785,N_1754);
xnor U1836 (N_1836,N_1773,N_1738);
nor U1837 (N_1837,N_1795,N_1729);
nand U1838 (N_1838,N_1727,N_1748);
or U1839 (N_1839,N_1794,N_1758);
nor U1840 (N_1840,N_1733,N_1767);
and U1841 (N_1841,N_1778,N_1792);
and U1842 (N_1842,N_1795,N_1733);
or U1843 (N_1843,N_1796,N_1742);
nand U1844 (N_1844,N_1738,N_1734);
and U1845 (N_1845,N_1788,N_1740);
or U1846 (N_1846,N_1733,N_1735);
or U1847 (N_1847,N_1792,N_1755);
nand U1848 (N_1848,N_1754,N_1769);
nor U1849 (N_1849,N_1733,N_1797);
nor U1850 (N_1850,N_1734,N_1768);
or U1851 (N_1851,N_1776,N_1766);
and U1852 (N_1852,N_1774,N_1788);
nand U1853 (N_1853,N_1757,N_1772);
nand U1854 (N_1854,N_1789,N_1799);
nor U1855 (N_1855,N_1732,N_1791);
and U1856 (N_1856,N_1759,N_1777);
xor U1857 (N_1857,N_1742,N_1740);
and U1858 (N_1858,N_1736,N_1798);
nand U1859 (N_1859,N_1725,N_1786);
nand U1860 (N_1860,N_1779,N_1756);
nand U1861 (N_1861,N_1783,N_1764);
or U1862 (N_1862,N_1779,N_1767);
nor U1863 (N_1863,N_1787,N_1776);
or U1864 (N_1864,N_1748,N_1758);
or U1865 (N_1865,N_1771,N_1787);
and U1866 (N_1866,N_1786,N_1777);
or U1867 (N_1867,N_1745,N_1762);
nor U1868 (N_1868,N_1751,N_1781);
and U1869 (N_1869,N_1761,N_1735);
nand U1870 (N_1870,N_1733,N_1761);
nor U1871 (N_1871,N_1792,N_1727);
nor U1872 (N_1872,N_1753,N_1743);
nor U1873 (N_1873,N_1789,N_1739);
nor U1874 (N_1874,N_1799,N_1761);
and U1875 (N_1875,N_1859,N_1829);
nor U1876 (N_1876,N_1844,N_1851);
or U1877 (N_1877,N_1871,N_1848);
xnor U1878 (N_1878,N_1822,N_1856);
and U1879 (N_1879,N_1837,N_1864);
nand U1880 (N_1880,N_1839,N_1835);
nand U1881 (N_1881,N_1803,N_1872);
nand U1882 (N_1882,N_1868,N_1857);
and U1883 (N_1883,N_1849,N_1815);
and U1884 (N_1884,N_1841,N_1833);
or U1885 (N_1885,N_1805,N_1874);
nor U1886 (N_1886,N_1850,N_1823);
nor U1887 (N_1887,N_1870,N_1812);
nand U1888 (N_1888,N_1855,N_1828);
and U1889 (N_1889,N_1852,N_1846);
and U1890 (N_1890,N_1873,N_1827);
nand U1891 (N_1891,N_1824,N_1819);
nor U1892 (N_1892,N_1831,N_1863);
or U1893 (N_1893,N_1807,N_1826);
or U1894 (N_1894,N_1820,N_1858);
and U1895 (N_1895,N_1802,N_1806);
or U1896 (N_1896,N_1810,N_1853);
nor U1897 (N_1897,N_1845,N_1847);
nor U1898 (N_1898,N_1865,N_1811);
or U1899 (N_1899,N_1860,N_1862);
nand U1900 (N_1900,N_1842,N_1854);
nor U1901 (N_1901,N_1866,N_1836);
nand U1902 (N_1902,N_1840,N_1818);
and U1903 (N_1903,N_1834,N_1804);
and U1904 (N_1904,N_1867,N_1817);
nor U1905 (N_1905,N_1825,N_1814);
nand U1906 (N_1906,N_1832,N_1843);
and U1907 (N_1907,N_1800,N_1809);
nand U1908 (N_1908,N_1838,N_1816);
or U1909 (N_1909,N_1830,N_1861);
and U1910 (N_1910,N_1808,N_1813);
or U1911 (N_1911,N_1821,N_1801);
and U1912 (N_1912,N_1869,N_1825);
nor U1913 (N_1913,N_1801,N_1828);
or U1914 (N_1914,N_1844,N_1828);
nor U1915 (N_1915,N_1870,N_1854);
or U1916 (N_1916,N_1802,N_1811);
nor U1917 (N_1917,N_1858,N_1836);
or U1918 (N_1918,N_1833,N_1862);
and U1919 (N_1919,N_1865,N_1803);
nand U1920 (N_1920,N_1845,N_1805);
or U1921 (N_1921,N_1868,N_1821);
or U1922 (N_1922,N_1806,N_1819);
and U1923 (N_1923,N_1801,N_1873);
nor U1924 (N_1924,N_1853,N_1862);
and U1925 (N_1925,N_1841,N_1809);
or U1926 (N_1926,N_1819,N_1831);
and U1927 (N_1927,N_1828,N_1808);
and U1928 (N_1928,N_1856,N_1807);
nand U1929 (N_1929,N_1872,N_1825);
or U1930 (N_1930,N_1868,N_1869);
and U1931 (N_1931,N_1846,N_1853);
or U1932 (N_1932,N_1814,N_1850);
or U1933 (N_1933,N_1819,N_1873);
nand U1934 (N_1934,N_1826,N_1827);
and U1935 (N_1935,N_1840,N_1852);
and U1936 (N_1936,N_1850,N_1800);
or U1937 (N_1937,N_1811,N_1858);
and U1938 (N_1938,N_1862,N_1814);
and U1939 (N_1939,N_1854,N_1816);
nand U1940 (N_1940,N_1829,N_1840);
nand U1941 (N_1941,N_1834,N_1823);
and U1942 (N_1942,N_1855,N_1839);
or U1943 (N_1943,N_1826,N_1845);
or U1944 (N_1944,N_1803,N_1856);
xor U1945 (N_1945,N_1873,N_1842);
nor U1946 (N_1946,N_1824,N_1810);
and U1947 (N_1947,N_1812,N_1811);
nor U1948 (N_1948,N_1816,N_1864);
nor U1949 (N_1949,N_1811,N_1856);
or U1950 (N_1950,N_1885,N_1895);
or U1951 (N_1951,N_1892,N_1893);
nand U1952 (N_1952,N_1916,N_1937);
nor U1953 (N_1953,N_1942,N_1940);
nand U1954 (N_1954,N_1906,N_1930);
and U1955 (N_1955,N_1917,N_1941);
or U1956 (N_1956,N_1887,N_1878);
or U1957 (N_1957,N_1896,N_1905);
nand U1958 (N_1958,N_1919,N_1901);
or U1959 (N_1959,N_1909,N_1934);
and U1960 (N_1960,N_1932,N_1914);
nand U1961 (N_1961,N_1927,N_1943);
or U1962 (N_1962,N_1904,N_1888);
nor U1963 (N_1963,N_1881,N_1924);
and U1964 (N_1964,N_1931,N_1898);
nand U1965 (N_1965,N_1939,N_1913);
nor U1966 (N_1966,N_1938,N_1947);
xor U1967 (N_1967,N_1907,N_1876);
xor U1968 (N_1968,N_1889,N_1910);
and U1969 (N_1969,N_1882,N_1899);
and U1970 (N_1970,N_1875,N_1925);
or U1971 (N_1971,N_1922,N_1923);
and U1972 (N_1972,N_1890,N_1935);
nor U1973 (N_1973,N_1894,N_1884);
and U1974 (N_1974,N_1897,N_1886);
and U1975 (N_1975,N_1929,N_1891);
xor U1976 (N_1976,N_1877,N_1928);
nand U1977 (N_1977,N_1926,N_1946);
and U1978 (N_1978,N_1908,N_1883);
or U1979 (N_1979,N_1903,N_1949);
nand U1980 (N_1980,N_1945,N_1918);
nor U1981 (N_1981,N_1879,N_1911);
nand U1982 (N_1982,N_1902,N_1936);
nand U1983 (N_1983,N_1915,N_1933);
nand U1984 (N_1984,N_1880,N_1920);
nor U1985 (N_1985,N_1912,N_1900);
nand U1986 (N_1986,N_1921,N_1944);
or U1987 (N_1987,N_1948,N_1926);
nand U1988 (N_1988,N_1879,N_1918);
nor U1989 (N_1989,N_1948,N_1897);
nor U1990 (N_1990,N_1905,N_1941);
and U1991 (N_1991,N_1907,N_1898);
and U1992 (N_1992,N_1934,N_1887);
or U1993 (N_1993,N_1933,N_1947);
xor U1994 (N_1994,N_1918,N_1921);
nor U1995 (N_1995,N_1876,N_1919);
nor U1996 (N_1996,N_1946,N_1937);
xnor U1997 (N_1997,N_1914,N_1879);
or U1998 (N_1998,N_1917,N_1899);
nor U1999 (N_1999,N_1924,N_1892);
nand U2000 (N_2000,N_1937,N_1920);
xnor U2001 (N_2001,N_1937,N_1914);
nand U2002 (N_2002,N_1916,N_1878);
and U2003 (N_2003,N_1888,N_1949);
or U2004 (N_2004,N_1926,N_1937);
nor U2005 (N_2005,N_1899,N_1909);
nand U2006 (N_2006,N_1921,N_1920);
nand U2007 (N_2007,N_1912,N_1896);
or U2008 (N_2008,N_1877,N_1934);
nand U2009 (N_2009,N_1946,N_1901);
nor U2010 (N_2010,N_1917,N_1907);
nor U2011 (N_2011,N_1878,N_1888);
nor U2012 (N_2012,N_1883,N_1920);
nand U2013 (N_2013,N_1938,N_1914);
nor U2014 (N_2014,N_1890,N_1932);
nor U2015 (N_2015,N_1884,N_1877);
xnor U2016 (N_2016,N_1921,N_1883);
or U2017 (N_2017,N_1932,N_1944);
or U2018 (N_2018,N_1946,N_1888);
nand U2019 (N_2019,N_1918,N_1911);
or U2020 (N_2020,N_1876,N_1901);
nand U2021 (N_2021,N_1908,N_1902);
nor U2022 (N_2022,N_1888,N_1939);
nand U2023 (N_2023,N_1919,N_1896);
nand U2024 (N_2024,N_1930,N_1945);
or U2025 (N_2025,N_1982,N_1974);
or U2026 (N_2026,N_2013,N_1967);
and U2027 (N_2027,N_1977,N_1998);
and U2028 (N_2028,N_2003,N_1963);
nor U2029 (N_2029,N_1979,N_2018);
nor U2030 (N_2030,N_2007,N_1980);
nor U2031 (N_2031,N_1970,N_2009);
and U2032 (N_2032,N_2024,N_1973);
or U2033 (N_2033,N_1984,N_1965);
nor U2034 (N_2034,N_2022,N_1995);
nand U2035 (N_2035,N_1990,N_1952);
nand U2036 (N_2036,N_1962,N_2015);
nor U2037 (N_2037,N_1964,N_1993);
or U2038 (N_2038,N_1985,N_1950);
and U2039 (N_2039,N_1961,N_1981);
nand U2040 (N_2040,N_2002,N_1954);
nand U2041 (N_2041,N_1986,N_1960);
nand U2042 (N_2042,N_2004,N_1966);
and U2043 (N_2043,N_2008,N_1953);
nor U2044 (N_2044,N_1957,N_1972);
and U2045 (N_2045,N_2021,N_1996);
or U2046 (N_2046,N_1992,N_1956);
nor U2047 (N_2047,N_1959,N_2005);
nor U2048 (N_2048,N_1969,N_1955);
nand U2049 (N_2049,N_1999,N_2011);
and U2050 (N_2050,N_1989,N_1971);
nor U2051 (N_2051,N_2017,N_2000);
nand U2052 (N_2052,N_2014,N_2016);
or U2053 (N_2053,N_1988,N_2010);
and U2054 (N_2054,N_1968,N_1994);
or U2055 (N_2055,N_2019,N_1958);
nor U2056 (N_2056,N_2001,N_1997);
and U2057 (N_2057,N_1991,N_2006);
nor U2058 (N_2058,N_1951,N_1975);
and U2059 (N_2059,N_1983,N_2012);
nand U2060 (N_2060,N_2023,N_1987);
or U2061 (N_2061,N_1976,N_2020);
nor U2062 (N_2062,N_1978,N_2007);
or U2063 (N_2063,N_1975,N_2004);
nor U2064 (N_2064,N_1964,N_1971);
and U2065 (N_2065,N_1953,N_1985);
and U2066 (N_2066,N_1952,N_1999);
nor U2067 (N_2067,N_1953,N_2021);
nor U2068 (N_2068,N_1981,N_1951);
nand U2069 (N_2069,N_1996,N_1958);
and U2070 (N_2070,N_1954,N_2003);
or U2071 (N_2071,N_1965,N_1961);
nor U2072 (N_2072,N_1998,N_1968);
and U2073 (N_2073,N_2014,N_1961);
and U2074 (N_2074,N_1988,N_1961);
nand U2075 (N_2075,N_1969,N_1962);
or U2076 (N_2076,N_2015,N_2014);
nand U2077 (N_2077,N_1962,N_1950);
or U2078 (N_2078,N_2018,N_1970);
nand U2079 (N_2079,N_1959,N_1958);
and U2080 (N_2080,N_1979,N_1985);
nor U2081 (N_2081,N_1987,N_1952);
nor U2082 (N_2082,N_1987,N_2000);
nand U2083 (N_2083,N_1959,N_1953);
and U2084 (N_2084,N_1988,N_2022);
nor U2085 (N_2085,N_1952,N_1975);
nand U2086 (N_2086,N_1981,N_1977);
or U2087 (N_2087,N_2022,N_1967);
nor U2088 (N_2088,N_2023,N_1964);
and U2089 (N_2089,N_1994,N_1969);
nor U2090 (N_2090,N_1986,N_2001);
nor U2091 (N_2091,N_1957,N_2010);
nand U2092 (N_2092,N_1987,N_1999);
and U2093 (N_2093,N_1993,N_1991);
nand U2094 (N_2094,N_1957,N_1958);
and U2095 (N_2095,N_1972,N_2005);
nor U2096 (N_2096,N_1959,N_2017);
nand U2097 (N_2097,N_1965,N_1979);
nor U2098 (N_2098,N_1971,N_1983);
and U2099 (N_2099,N_1984,N_1987);
or U2100 (N_2100,N_2078,N_2076);
or U2101 (N_2101,N_2073,N_2079);
and U2102 (N_2102,N_2033,N_2056);
nand U2103 (N_2103,N_2055,N_2094);
nor U2104 (N_2104,N_2068,N_2038);
and U2105 (N_2105,N_2044,N_2083);
nand U2106 (N_2106,N_2090,N_2046);
and U2107 (N_2107,N_2095,N_2035);
nand U2108 (N_2108,N_2036,N_2045);
and U2109 (N_2109,N_2075,N_2074);
nor U2110 (N_2110,N_2039,N_2071);
and U2111 (N_2111,N_2086,N_2061);
nor U2112 (N_2112,N_2058,N_2081);
or U2113 (N_2113,N_2072,N_2064);
and U2114 (N_2114,N_2047,N_2091);
nor U2115 (N_2115,N_2085,N_2030);
nor U2116 (N_2116,N_2054,N_2084);
or U2117 (N_2117,N_2026,N_2087);
or U2118 (N_2118,N_2028,N_2067);
or U2119 (N_2119,N_2093,N_2089);
nor U2120 (N_2120,N_2041,N_2037);
or U2121 (N_2121,N_2066,N_2042);
and U2122 (N_2122,N_2057,N_2040);
nor U2123 (N_2123,N_2059,N_2098);
nand U2124 (N_2124,N_2096,N_2048);
or U2125 (N_2125,N_2077,N_2099);
nor U2126 (N_2126,N_2088,N_2032);
nand U2127 (N_2127,N_2049,N_2027);
nand U2128 (N_2128,N_2062,N_2034);
or U2129 (N_2129,N_2092,N_2070);
nor U2130 (N_2130,N_2051,N_2082);
and U2131 (N_2131,N_2069,N_2097);
nand U2132 (N_2132,N_2031,N_2053);
or U2133 (N_2133,N_2029,N_2052);
or U2134 (N_2134,N_2065,N_2043);
or U2135 (N_2135,N_2063,N_2080);
or U2136 (N_2136,N_2025,N_2060);
or U2137 (N_2137,N_2050,N_2088);
nor U2138 (N_2138,N_2075,N_2045);
and U2139 (N_2139,N_2098,N_2043);
or U2140 (N_2140,N_2084,N_2032);
nand U2141 (N_2141,N_2090,N_2025);
or U2142 (N_2142,N_2092,N_2049);
and U2143 (N_2143,N_2066,N_2039);
or U2144 (N_2144,N_2072,N_2059);
nand U2145 (N_2145,N_2065,N_2091);
nor U2146 (N_2146,N_2083,N_2064);
nor U2147 (N_2147,N_2045,N_2092);
and U2148 (N_2148,N_2080,N_2090);
nand U2149 (N_2149,N_2062,N_2029);
nor U2150 (N_2150,N_2089,N_2071);
or U2151 (N_2151,N_2054,N_2074);
nand U2152 (N_2152,N_2072,N_2094);
nor U2153 (N_2153,N_2073,N_2093);
nor U2154 (N_2154,N_2026,N_2080);
or U2155 (N_2155,N_2032,N_2034);
or U2156 (N_2156,N_2074,N_2029);
nand U2157 (N_2157,N_2054,N_2088);
or U2158 (N_2158,N_2068,N_2042);
xor U2159 (N_2159,N_2066,N_2084);
and U2160 (N_2160,N_2051,N_2075);
nor U2161 (N_2161,N_2051,N_2065);
nand U2162 (N_2162,N_2049,N_2035);
and U2163 (N_2163,N_2042,N_2078);
or U2164 (N_2164,N_2093,N_2082);
nand U2165 (N_2165,N_2029,N_2030);
nor U2166 (N_2166,N_2041,N_2085);
nand U2167 (N_2167,N_2082,N_2097);
and U2168 (N_2168,N_2076,N_2049);
nor U2169 (N_2169,N_2075,N_2065);
or U2170 (N_2170,N_2058,N_2051);
and U2171 (N_2171,N_2072,N_2028);
nand U2172 (N_2172,N_2097,N_2038);
nand U2173 (N_2173,N_2055,N_2079);
nand U2174 (N_2174,N_2075,N_2025);
or U2175 (N_2175,N_2104,N_2106);
nand U2176 (N_2176,N_2152,N_2121);
nand U2177 (N_2177,N_2164,N_2102);
and U2178 (N_2178,N_2171,N_2107);
nor U2179 (N_2179,N_2150,N_2147);
and U2180 (N_2180,N_2163,N_2112);
xor U2181 (N_2181,N_2105,N_2137);
nor U2182 (N_2182,N_2125,N_2143);
and U2183 (N_2183,N_2158,N_2127);
or U2184 (N_2184,N_2154,N_2135);
and U2185 (N_2185,N_2169,N_2146);
and U2186 (N_2186,N_2172,N_2166);
and U2187 (N_2187,N_2110,N_2123);
and U2188 (N_2188,N_2140,N_2159);
and U2189 (N_2189,N_2124,N_2145);
xor U2190 (N_2190,N_2162,N_2132);
xnor U2191 (N_2191,N_2100,N_2113);
nand U2192 (N_2192,N_2153,N_2130);
nor U2193 (N_2193,N_2148,N_2156);
or U2194 (N_2194,N_2151,N_2138);
and U2195 (N_2195,N_2133,N_2170);
and U2196 (N_2196,N_2111,N_2157);
nor U2197 (N_2197,N_2141,N_2115);
or U2198 (N_2198,N_2128,N_2165);
or U2199 (N_2199,N_2101,N_2109);
nor U2200 (N_2200,N_2119,N_2167);
or U2201 (N_2201,N_2173,N_2134);
nor U2202 (N_2202,N_2139,N_2144);
or U2203 (N_2203,N_2108,N_2103);
xnor U2204 (N_2204,N_2120,N_2161);
nor U2205 (N_2205,N_2168,N_2155);
or U2206 (N_2206,N_2116,N_2114);
nand U2207 (N_2207,N_2122,N_2160);
or U2208 (N_2208,N_2136,N_2126);
nand U2209 (N_2209,N_2117,N_2149);
nand U2210 (N_2210,N_2142,N_2129);
or U2211 (N_2211,N_2174,N_2131);
and U2212 (N_2212,N_2118,N_2116);
or U2213 (N_2213,N_2165,N_2155);
nand U2214 (N_2214,N_2107,N_2167);
and U2215 (N_2215,N_2156,N_2107);
nor U2216 (N_2216,N_2130,N_2129);
nand U2217 (N_2217,N_2137,N_2107);
nand U2218 (N_2218,N_2106,N_2151);
and U2219 (N_2219,N_2114,N_2107);
xnor U2220 (N_2220,N_2123,N_2151);
or U2221 (N_2221,N_2152,N_2132);
and U2222 (N_2222,N_2101,N_2149);
xnor U2223 (N_2223,N_2154,N_2125);
nor U2224 (N_2224,N_2147,N_2105);
or U2225 (N_2225,N_2133,N_2151);
or U2226 (N_2226,N_2154,N_2152);
nor U2227 (N_2227,N_2130,N_2173);
nand U2228 (N_2228,N_2138,N_2112);
and U2229 (N_2229,N_2154,N_2139);
and U2230 (N_2230,N_2145,N_2108);
nor U2231 (N_2231,N_2144,N_2163);
and U2232 (N_2232,N_2152,N_2124);
nor U2233 (N_2233,N_2117,N_2162);
nand U2234 (N_2234,N_2161,N_2172);
xnor U2235 (N_2235,N_2133,N_2113);
nand U2236 (N_2236,N_2115,N_2108);
nand U2237 (N_2237,N_2140,N_2100);
and U2238 (N_2238,N_2163,N_2126);
nand U2239 (N_2239,N_2145,N_2101);
or U2240 (N_2240,N_2100,N_2155);
or U2241 (N_2241,N_2104,N_2139);
nor U2242 (N_2242,N_2173,N_2123);
nand U2243 (N_2243,N_2161,N_2158);
nor U2244 (N_2244,N_2139,N_2130);
nand U2245 (N_2245,N_2109,N_2119);
or U2246 (N_2246,N_2100,N_2105);
or U2247 (N_2247,N_2114,N_2174);
nor U2248 (N_2248,N_2109,N_2165);
nand U2249 (N_2249,N_2172,N_2135);
nor U2250 (N_2250,N_2227,N_2194);
and U2251 (N_2251,N_2238,N_2244);
nand U2252 (N_2252,N_2178,N_2230);
nor U2253 (N_2253,N_2240,N_2243);
and U2254 (N_2254,N_2217,N_2212);
or U2255 (N_2255,N_2228,N_2234);
and U2256 (N_2256,N_2193,N_2204);
nor U2257 (N_2257,N_2209,N_2220);
nand U2258 (N_2258,N_2199,N_2233);
nand U2259 (N_2259,N_2248,N_2241);
or U2260 (N_2260,N_2218,N_2231);
nor U2261 (N_2261,N_2188,N_2210);
xnor U2262 (N_2262,N_2191,N_2207);
and U2263 (N_2263,N_2179,N_2232);
or U2264 (N_2264,N_2206,N_2180);
nand U2265 (N_2265,N_2195,N_2176);
nor U2266 (N_2266,N_2181,N_2200);
or U2267 (N_2267,N_2236,N_2183);
and U2268 (N_2268,N_2196,N_2214);
nor U2269 (N_2269,N_2201,N_2242);
nor U2270 (N_2270,N_2246,N_2237);
nor U2271 (N_2271,N_2216,N_2205);
nor U2272 (N_2272,N_2239,N_2247);
or U2273 (N_2273,N_2202,N_2229);
or U2274 (N_2274,N_2215,N_2185);
nand U2275 (N_2275,N_2186,N_2190);
nand U2276 (N_2276,N_2175,N_2184);
or U2277 (N_2277,N_2223,N_2189);
and U2278 (N_2278,N_2187,N_2226);
and U2279 (N_2279,N_2222,N_2235);
and U2280 (N_2280,N_2177,N_2224);
nor U2281 (N_2281,N_2192,N_2182);
nor U2282 (N_2282,N_2213,N_2245);
xor U2283 (N_2283,N_2197,N_2221);
and U2284 (N_2284,N_2225,N_2249);
nor U2285 (N_2285,N_2198,N_2211);
xor U2286 (N_2286,N_2203,N_2208);
and U2287 (N_2287,N_2219,N_2225);
nand U2288 (N_2288,N_2193,N_2231);
and U2289 (N_2289,N_2228,N_2240);
nor U2290 (N_2290,N_2240,N_2192);
and U2291 (N_2291,N_2177,N_2239);
nor U2292 (N_2292,N_2200,N_2238);
nand U2293 (N_2293,N_2180,N_2244);
or U2294 (N_2294,N_2192,N_2183);
nor U2295 (N_2295,N_2194,N_2221);
or U2296 (N_2296,N_2224,N_2235);
or U2297 (N_2297,N_2208,N_2240);
or U2298 (N_2298,N_2243,N_2193);
and U2299 (N_2299,N_2249,N_2234);
nor U2300 (N_2300,N_2225,N_2242);
nand U2301 (N_2301,N_2222,N_2238);
or U2302 (N_2302,N_2244,N_2218);
or U2303 (N_2303,N_2180,N_2179);
nor U2304 (N_2304,N_2228,N_2211);
and U2305 (N_2305,N_2247,N_2202);
nor U2306 (N_2306,N_2183,N_2246);
or U2307 (N_2307,N_2241,N_2191);
or U2308 (N_2308,N_2197,N_2208);
or U2309 (N_2309,N_2244,N_2245);
nor U2310 (N_2310,N_2249,N_2224);
and U2311 (N_2311,N_2190,N_2228);
nand U2312 (N_2312,N_2231,N_2217);
nand U2313 (N_2313,N_2201,N_2241);
or U2314 (N_2314,N_2244,N_2239);
or U2315 (N_2315,N_2246,N_2245);
nand U2316 (N_2316,N_2212,N_2209);
or U2317 (N_2317,N_2249,N_2181);
nor U2318 (N_2318,N_2236,N_2242);
and U2319 (N_2319,N_2233,N_2180);
and U2320 (N_2320,N_2177,N_2176);
xnor U2321 (N_2321,N_2234,N_2243);
nor U2322 (N_2322,N_2201,N_2237);
nand U2323 (N_2323,N_2233,N_2238);
nor U2324 (N_2324,N_2233,N_2201);
nand U2325 (N_2325,N_2282,N_2260);
nand U2326 (N_2326,N_2261,N_2311);
nor U2327 (N_2327,N_2285,N_2317);
and U2328 (N_2328,N_2316,N_2280);
or U2329 (N_2329,N_2255,N_2269);
nor U2330 (N_2330,N_2304,N_2296);
nand U2331 (N_2331,N_2262,N_2273);
nand U2332 (N_2332,N_2319,N_2297);
nand U2333 (N_2333,N_2310,N_2251);
or U2334 (N_2334,N_2307,N_2279);
and U2335 (N_2335,N_2266,N_2277);
nor U2336 (N_2336,N_2299,N_2284);
or U2337 (N_2337,N_2286,N_2292);
or U2338 (N_2338,N_2287,N_2265);
and U2339 (N_2339,N_2303,N_2256);
nand U2340 (N_2340,N_2301,N_2278);
nor U2341 (N_2341,N_2270,N_2276);
nor U2342 (N_2342,N_2298,N_2254);
nand U2343 (N_2343,N_2259,N_2290);
or U2344 (N_2344,N_2318,N_2283);
nor U2345 (N_2345,N_2313,N_2288);
nor U2346 (N_2346,N_2323,N_2321);
and U2347 (N_2347,N_2264,N_2306);
and U2348 (N_2348,N_2294,N_2268);
or U2349 (N_2349,N_2312,N_2305);
or U2350 (N_2350,N_2253,N_2308);
nor U2351 (N_2351,N_2272,N_2250);
nor U2352 (N_2352,N_2324,N_2293);
and U2353 (N_2353,N_2252,N_2302);
nor U2354 (N_2354,N_2271,N_2309);
nand U2355 (N_2355,N_2257,N_2274);
nand U2356 (N_2356,N_2320,N_2291);
nand U2357 (N_2357,N_2263,N_2281);
or U2358 (N_2358,N_2275,N_2300);
or U2359 (N_2359,N_2314,N_2267);
nor U2360 (N_2360,N_2258,N_2295);
and U2361 (N_2361,N_2322,N_2315);
nand U2362 (N_2362,N_2289,N_2281);
or U2363 (N_2363,N_2299,N_2313);
nor U2364 (N_2364,N_2310,N_2295);
nand U2365 (N_2365,N_2288,N_2260);
nor U2366 (N_2366,N_2303,N_2278);
xor U2367 (N_2367,N_2305,N_2322);
nor U2368 (N_2368,N_2260,N_2259);
nand U2369 (N_2369,N_2321,N_2289);
or U2370 (N_2370,N_2316,N_2295);
nand U2371 (N_2371,N_2306,N_2273);
nor U2372 (N_2372,N_2280,N_2267);
or U2373 (N_2373,N_2252,N_2272);
nand U2374 (N_2374,N_2294,N_2295);
and U2375 (N_2375,N_2294,N_2313);
nor U2376 (N_2376,N_2297,N_2318);
and U2377 (N_2377,N_2251,N_2259);
or U2378 (N_2378,N_2260,N_2305);
xnor U2379 (N_2379,N_2270,N_2305);
nand U2380 (N_2380,N_2323,N_2281);
nor U2381 (N_2381,N_2270,N_2314);
nand U2382 (N_2382,N_2279,N_2278);
nand U2383 (N_2383,N_2316,N_2252);
nor U2384 (N_2384,N_2299,N_2251);
and U2385 (N_2385,N_2294,N_2303);
nor U2386 (N_2386,N_2307,N_2259);
nand U2387 (N_2387,N_2311,N_2283);
or U2388 (N_2388,N_2263,N_2270);
and U2389 (N_2389,N_2302,N_2268);
nand U2390 (N_2390,N_2312,N_2322);
or U2391 (N_2391,N_2252,N_2250);
nand U2392 (N_2392,N_2317,N_2288);
xnor U2393 (N_2393,N_2275,N_2256);
nand U2394 (N_2394,N_2282,N_2266);
and U2395 (N_2395,N_2295,N_2299);
nor U2396 (N_2396,N_2306,N_2254);
nand U2397 (N_2397,N_2253,N_2312);
or U2398 (N_2398,N_2270,N_2273);
nand U2399 (N_2399,N_2261,N_2291);
or U2400 (N_2400,N_2339,N_2377);
nor U2401 (N_2401,N_2380,N_2344);
nor U2402 (N_2402,N_2326,N_2395);
or U2403 (N_2403,N_2362,N_2361);
or U2404 (N_2404,N_2349,N_2371);
or U2405 (N_2405,N_2375,N_2368);
and U2406 (N_2406,N_2378,N_2381);
or U2407 (N_2407,N_2336,N_2342);
nand U2408 (N_2408,N_2391,N_2338);
nand U2409 (N_2409,N_2348,N_2389);
and U2410 (N_2410,N_2383,N_2356);
nor U2411 (N_2411,N_2385,N_2372);
xor U2412 (N_2412,N_2328,N_2343);
nand U2413 (N_2413,N_2366,N_2393);
or U2414 (N_2414,N_2330,N_2327);
nor U2415 (N_2415,N_2350,N_2352);
nor U2416 (N_2416,N_2384,N_2390);
or U2417 (N_2417,N_2386,N_2382);
xnor U2418 (N_2418,N_2388,N_2329);
nor U2419 (N_2419,N_2359,N_2370);
nand U2420 (N_2420,N_2379,N_2351);
or U2421 (N_2421,N_2396,N_2394);
nor U2422 (N_2422,N_2364,N_2399);
or U2423 (N_2423,N_2358,N_2376);
or U2424 (N_2424,N_2397,N_2354);
nand U2425 (N_2425,N_2363,N_2341);
or U2426 (N_2426,N_2346,N_2355);
or U2427 (N_2427,N_2369,N_2340);
or U2428 (N_2428,N_2345,N_2373);
nor U2429 (N_2429,N_2325,N_2360);
nand U2430 (N_2430,N_2357,N_2333);
nor U2431 (N_2431,N_2392,N_2337);
nand U2432 (N_2432,N_2353,N_2367);
nand U2433 (N_2433,N_2332,N_2334);
nor U2434 (N_2434,N_2387,N_2331);
nor U2435 (N_2435,N_2335,N_2365);
nor U2436 (N_2436,N_2398,N_2374);
xnor U2437 (N_2437,N_2347,N_2340);
and U2438 (N_2438,N_2353,N_2347);
nand U2439 (N_2439,N_2329,N_2335);
nand U2440 (N_2440,N_2382,N_2349);
nand U2441 (N_2441,N_2349,N_2334);
nand U2442 (N_2442,N_2385,N_2393);
or U2443 (N_2443,N_2378,N_2343);
or U2444 (N_2444,N_2353,N_2383);
and U2445 (N_2445,N_2348,N_2336);
nand U2446 (N_2446,N_2335,N_2368);
or U2447 (N_2447,N_2390,N_2362);
and U2448 (N_2448,N_2381,N_2336);
or U2449 (N_2449,N_2391,N_2382);
nor U2450 (N_2450,N_2387,N_2367);
or U2451 (N_2451,N_2343,N_2399);
nand U2452 (N_2452,N_2358,N_2331);
and U2453 (N_2453,N_2387,N_2397);
and U2454 (N_2454,N_2380,N_2362);
nand U2455 (N_2455,N_2380,N_2359);
nor U2456 (N_2456,N_2361,N_2339);
or U2457 (N_2457,N_2333,N_2351);
nor U2458 (N_2458,N_2396,N_2328);
and U2459 (N_2459,N_2337,N_2343);
nand U2460 (N_2460,N_2388,N_2359);
nor U2461 (N_2461,N_2380,N_2393);
or U2462 (N_2462,N_2332,N_2353);
nor U2463 (N_2463,N_2392,N_2399);
and U2464 (N_2464,N_2385,N_2356);
and U2465 (N_2465,N_2376,N_2349);
and U2466 (N_2466,N_2394,N_2341);
and U2467 (N_2467,N_2371,N_2355);
nor U2468 (N_2468,N_2383,N_2360);
and U2469 (N_2469,N_2369,N_2362);
and U2470 (N_2470,N_2329,N_2340);
nor U2471 (N_2471,N_2333,N_2371);
nand U2472 (N_2472,N_2397,N_2371);
or U2473 (N_2473,N_2392,N_2369);
nand U2474 (N_2474,N_2385,N_2340);
or U2475 (N_2475,N_2460,N_2429);
nand U2476 (N_2476,N_2423,N_2440);
xor U2477 (N_2477,N_2431,N_2467);
nor U2478 (N_2478,N_2404,N_2471);
or U2479 (N_2479,N_2448,N_2470);
and U2480 (N_2480,N_2434,N_2441);
nand U2481 (N_2481,N_2419,N_2453);
nor U2482 (N_2482,N_2407,N_2462);
nor U2483 (N_2483,N_2401,N_2450);
xor U2484 (N_2484,N_2474,N_2417);
or U2485 (N_2485,N_2415,N_2436);
nand U2486 (N_2486,N_2459,N_2439);
and U2487 (N_2487,N_2402,N_2438);
nor U2488 (N_2488,N_2444,N_2428);
or U2489 (N_2489,N_2463,N_2425);
nand U2490 (N_2490,N_2451,N_2447);
or U2491 (N_2491,N_2426,N_2424);
nor U2492 (N_2492,N_2435,N_2400);
or U2493 (N_2493,N_2442,N_2464);
nand U2494 (N_2494,N_2445,N_2437);
and U2495 (N_2495,N_2432,N_2430);
and U2496 (N_2496,N_2458,N_2456);
or U2497 (N_2497,N_2472,N_2413);
or U2498 (N_2498,N_2433,N_2461);
nor U2499 (N_2499,N_2454,N_2457);
or U2500 (N_2500,N_2416,N_2422);
or U2501 (N_2501,N_2449,N_2411);
and U2502 (N_2502,N_2455,N_2465);
nor U2503 (N_2503,N_2412,N_2443);
nand U2504 (N_2504,N_2408,N_2421);
and U2505 (N_2505,N_2427,N_2406);
nand U2506 (N_2506,N_2414,N_2468);
nand U2507 (N_2507,N_2466,N_2405);
or U2508 (N_2508,N_2420,N_2452);
and U2509 (N_2509,N_2418,N_2473);
nand U2510 (N_2510,N_2403,N_2469);
or U2511 (N_2511,N_2409,N_2410);
nand U2512 (N_2512,N_2446,N_2441);
or U2513 (N_2513,N_2427,N_2472);
and U2514 (N_2514,N_2448,N_2450);
nor U2515 (N_2515,N_2415,N_2429);
and U2516 (N_2516,N_2414,N_2466);
and U2517 (N_2517,N_2464,N_2450);
nand U2518 (N_2518,N_2427,N_2417);
nand U2519 (N_2519,N_2447,N_2426);
or U2520 (N_2520,N_2455,N_2444);
or U2521 (N_2521,N_2425,N_2410);
nor U2522 (N_2522,N_2402,N_2459);
and U2523 (N_2523,N_2409,N_2425);
nor U2524 (N_2524,N_2411,N_2432);
or U2525 (N_2525,N_2458,N_2462);
nand U2526 (N_2526,N_2472,N_2464);
nand U2527 (N_2527,N_2432,N_2416);
and U2528 (N_2528,N_2406,N_2469);
nand U2529 (N_2529,N_2415,N_2432);
nor U2530 (N_2530,N_2474,N_2412);
or U2531 (N_2531,N_2448,N_2422);
or U2532 (N_2532,N_2403,N_2468);
nor U2533 (N_2533,N_2473,N_2441);
and U2534 (N_2534,N_2462,N_2438);
and U2535 (N_2535,N_2412,N_2430);
or U2536 (N_2536,N_2419,N_2454);
nor U2537 (N_2537,N_2409,N_2437);
nor U2538 (N_2538,N_2435,N_2440);
nor U2539 (N_2539,N_2417,N_2471);
and U2540 (N_2540,N_2467,N_2404);
and U2541 (N_2541,N_2415,N_2440);
or U2542 (N_2542,N_2439,N_2430);
or U2543 (N_2543,N_2423,N_2458);
nand U2544 (N_2544,N_2424,N_2438);
nor U2545 (N_2545,N_2401,N_2467);
or U2546 (N_2546,N_2466,N_2425);
and U2547 (N_2547,N_2441,N_2472);
or U2548 (N_2548,N_2430,N_2429);
nand U2549 (N_2549,N_2453,N_2432);
and U2550 (N_2550,N_2542,N_2534);
or U2551 (N_2551,N_2527,N_2544);
and U2552 (N_2552,N_2539,N_2512);
or U2553 (N_2553,N_2519,N_2496);
nand U2554 (N_2554,N_2511,N_2510);
xnor U2555 (N_2555,N_2517,N_2509);
nand U2556 (N_2556,N_2481,N_2532);
or U2557 (N_2557,N_2545,N_2480);
nor U2558 (N_2558,N_2522,N_2475);
or U2559 (N_2559,N_2503,N_2515);
xor U2560 (N_2560,N_2484,N_2485);
xnor U2561 (N_2561,N_2477,N_2516);
or U2562 (N_2562,N_2483,N_2488);
nand U2563 (N_2563,N_2548,N_2502);
and U2564 (N_2564,N_2526,N_2518);
nand U2565 (N_2565,N_2500,N_2478);
nor U2566 (N_2566,N_2529,N_2541);
xor U2567 (N_2567,N_2501,N_2547);
and U2568 (N_2568,N_2530,N_2535);
and U2569 (N_2569,N_2524,N_2537);
nand U2570 (N_2570,N_2513,N_2505);
nor U2571 (N_2571,N_2495,N_2492);
and U2572 (N_2572,N_2494,N_2476);
and U2573 (N_2573,N_2546,N_2514);
and U2574 (N_2574,N_2493,N_2531);
nand U2575 (N_2575,N_2540,N_2486);
nand U2576 (N_2576,N_2533,N_2489);
or U2577 (N_2577,N_2543,N_2490);
nor U2578 (N_2578,N_2523,N_2508);
or U2579 (N_2579,N_2507,N_2506);
nand U2580 (N_2580,N_2491,N_2549);
and U2581 (N_2581,N_2521,N_2520);
nor U2582 (N_2582,N_2499,N_2482);
nand U2583 (N_2583,N_2525,N_2498);
nand U2584 (N_2584,N_2538,N_2487);
nand U2585 (N_2585,N_2504,N_2479);
or U2586 (N_2586,N_2528,N_2536);
nor U2587 (N_2587,N_2497,N_2500);
nand U2588 (N_2588,N_2503,N_2487);
and U2589 (N_2589,N_2523,N_2496);
nand U2590 (N_2590,N_2504,N_2480);
nor U2591 (N_2591,N_2513,N_2532);
and U2592 (N_2592,N_2487,N_2531);
or U2593 (N_2593,N_2508,N_2496);
or U2594 (N_2594,N_2529,N_2493);
nor U2595 (N_2595,N_2521,N_2519);
or U2596 (N_2596,N_2532,N_2498);
nand U2597 (N_2597,N_2531,N_2532);
and U2598 (N_2598,N_2488,N_2501);
nand U2599 (N_2599,N_2520,N_2548);
or U2600 (N_2600,N_2491,N_2506);
nand U2601 (N_2601,N_2529,N_2536);
nor U2602 (N_2602,N_2516,N_2492);
and U2603 (N_2603,N_2476,N_2520);
xnor U2604 (N_2604,N_2477,N_2475);
and U2605 (N_2605,N_2523,N_2485);
nand U2606 (N_2606,N_2522,N_2516);
and U2607 (N_2607,N_2503,N_2533);
nor U2608 (N_2608,N_2479,N_2511);
nand U2609 (N_2609,N_2527,N_2524);
xor U2610 (N_2610,N_2481,N_2549);
and U2611 (N_2611,N_2494,N_2533);
or U2612 (N_2612,N_2499,N_2525);
and U2613 (N_2613,N_2479,N_2501);
nor U2614 (N_2614,N_2482,N_2496);
and U2615 (N_2615,N_2486,N_2495);
nand U2616 (N_2616,N_2499,N_2508);
nor U2617 (N_2617,N_2532,N_2534);
and U2618 (N_2618,N_2534,N_2522);
and U2619 (N_2619,N_2498,N_2546);
or U2620 (N_2620,N_2493,N_2526);
nand U2621 (N_2621,N_2517,N_2525);
or U2622 (N_2622,N_2512,N_2531);
and U2623 (N_2623,N_2499,N_2494);
nor U2624 (N_2624,N_2499,N_2535);
nand U2625 (N_2625,N_2552,N_2592);
and U2626 (N_2626,N_2585,N_2586);
nor U2627 (N_2627,N_2596,N_2624);
nor U2628 (N_2628,N_2604,N_2594);
or U2629 (N_2629,N_2555,N_2583);
and U2630 (N_2630,N_2589,N_2581);
and U2631 (N_2631,N_2565,N_2558);
and U2632 (N_2632,N_2614,N_2600);
and U2633 (N_2633,N_2557,N_2587);
and U2634 (N_2634,N_2597,N_2578);
and U2635 (N_2635,N_2606,N_2562);
nor U2636 (N_2636,N_2553,N_2599);
xor U2637 (N_2637,N_2593,N_2556);
nor U2638 (N_2638,N_2619,N_2595);
nor U2639 (N_2639,N_2601,N_2571);
nor U2640 (N_2640,N_2603,N_2613);
nor U2641 (N_2641,N_2584,N_2563);
and U2642 (N_2642,N_2573,N_2611);
nor U2643 (N_2643,N_2550,N_2574);
nand U2644 (N_2644,N_2605,N_2590);
or U2645 (N_2645,N_2618,N_2576);
nor U2646 (N_2646,N_2580,N_2570);
nand U2647 (N_2647,N_2598,N_2551);
and U2648 (N_2648,N_2579,N_2567);
nor U2649 (N_2649,N_2566,N_2622);
nand U2650 (N_2650,N_2559,N_2616);
or U2651 (N_2651,N_2554,N_2620);
and U2652 (N_2652,N_2588,N_2572);
or U2653 (N_2653,N_2607,N_2568);
nor U2654 (N_2654,N_2617,N_2564);
or U2655 (N_2655,N_2577,N_2610);
nand U2656 (N_2656,N_2609,N_2615);
nor U2657 (N_2657,N_2561,N_2612);
nor U2658 (N_2658,N_2621,N_2623);
nand U2659 (N_2659,N_2602,N_2575);
or U2660 (N_2660,N_2608,N_2569);
nand U2661 (N_2661,N_2582,N_2591);
nand U2662 (N_2662,N_2560,N_2615);
or U2663 (N_2663,N_2557,N_2565);
nor U2664 (N_2664,N_2605,N_2570);
and U2665 (N_2665,N_2562,N_2623);
nand U2666 (N_2666,N_2586,N_2610);
or U2667 (N_2667,N_2563,N_2591);
or U2668 (N_2668,N_2594,N_2552);
and U2669 (N_2669,N_2616,N_2613);
nor U2670 (N_2670,N_2582,N_2550);
or U2671 (N_2671,N_2577,N_2595);
nand U2672 (N_2672,N_2597,N_2551);
and U2673 (N_2673,N_2550,N_2593);
and U2674 (N_2674,N_2566,N_2574);
and U2675 (N_2675,N_2611,N_2577);
nand U2676 (N_2676,N_2567,N_2609);
nand U2677 (N_2677,N_2585,N_2591);
nand U2678 (N_2678,N_2596,N_2620);
or U2679 (N_2679,N_2613,N_2624);
nand U2680 (N_2680,N_2565,N_2598);
nand U2681 (N_2681,N_2597,N_2618);
nor U2682 (N_2682,N_2608,N_2554);
nand U2683 (N_2683,N_2577,N_2568);
or U2684 (N_2684,N_2552,N_2589);
or U2685 (N_2685,N_2560,N_2550);
nand U2686 (N_2686,N_2594,N_2597);
nor U2687 (N_2687,N_2624,N_2580);
nor U2688 (N_2688,N_2621,N_2613);
nand U2689 (N_2689,N_2604,N_2606);
or U2690 (N_2690,N_2583,N_2620);
or U2691 (N_2691,N_2612,N_2582);
and U2692 (N_2692,N_2558,N_2556);
nand U2693 (N_2693,N_2580,N_2619);
nor U2694 (N_2694,N_2593,N_2620);
and U2695 (N_2695,N_2566,N_2552);
and U2696 (N_2696,N_2570,N_2556);
and U2697 (N_2697,N_2576,N_2588);
and U2698 (N_2698,N_2580,N_2614);
or U2699 (N_2699,N_2573,N_2592);
nand U2700 (N_2700,N_2697,N_2679);
or U2701 (N_2701,N_2660,N_2670);
and U2702 (N_2702,N_2661,N_2692);
nand U2703 (N_2703,N_2695,N_2686);
nand U2704 (N_2704,N_2635,N_2641);
xnor U2705 (N_2705,N_2676,N_2645);
nand U2706 (N_2706,N_2689,N_2637);
and U2707 (N_2707,N_2634,N_2656);
nand U2708 (N_2708,N_2651,N_2655);
nor U2709 (N_2709,N_2636,N_2663);
or U2710 (N_2710,N_2698,N_2646);
or U2711 (N_2711,N_2630,N_2629);
nand U2712 (N_2712,N_2625,N_2644);
or U2713 (N_2713,N_2628,N_2666);
nor U2714 (N_2714,N_2654,N_2684);
nor U2715 (N_2715,N_2649,N_2627);
nor U2716 (N_2716,N_2626,N_2642);
or U2717 (N_2717,N_2662,N_2677);
or U2718 (N_2718,N_2687,N_2690);
nor U2719 (N_2719,N_2675,N_2640);
or U2720 (N_2720,N_2632,N_2674);
nand U2721 (N_2721,N_2671,N_2678);
xor U2722 (N_2722,N_2631,N_2650);
and U2723 (N_2723,N_2685,N_2657);
or U2724 (N_2724,N_2682,N_2638);
nand U2725 (N_2725,N_2647,N_2639);
nand U2726 (N_2726,N_2643,N_2652);
nor U2727 (N_2727,N_2673,N_2633);
nand U2728 (N_2728,N_2664,N_2653);
and U2729 (N_2729,N_2694,N_2667);
nand U2730 (N_2730,N_2658,N_2688);
nand U2731 (N_2731,N_2699,N_2691);
or U2732 (N_2732,N_2672,N_2669);
and U2733 (N_2733,N_2693,N_2668);
nor U2734 (N_2734,N_2648,N_2683);
nand U2735 (N_2735,N_2696,N_2659);
nor U2736 (N_2736,N_2680,N_2681);
nand U2737 (N_2737,N_2665,N_2671);
nand U2738 (N_2738,N_2669,N_2679);
and U2739 (N_2739,N_2647,N_2668);
or U2740 (N_2740,N_2675,N_2630);
nand U2741 (N_2741,N_2625,N_2670);
and U2742 (N_2742,N_2639,N_2686);
nor U2743 (N_2743,N_2659,N_2699);
or U2744 (N_2744,N_2640,N_2627);
and U2745 (N_2745,N_2674,N_2633);
nand U2746 (N_2746,N_2636,N_2687);
nor U2747 (N_2747,N_2634,N_2659);
and U2748 (N_2748,N_2646,N_2658);
and U2749 (N_2749,N_2678,N_2677);
or U2750 (N_2750,N_2654,N_2634);
nand U2751 (N_2751,N_2627,N_2687);
nand U2752 (N_2752,N_2659,N_2663);
nand U2753 (N_2753,N_2646,N_2672);
or U2754 (N_2754,N_2630,N_2656);
and U2755 (N_2755,N_2697,N_2629);
or U2756 (N_2756,N_2641,N_2667);
nand U2757 (N_2757,N_2641,N_2697);
or U2758 (N_2758,N_2650,N_2643);
and U2759 (N_2759,N_2653,N_2651);
nor U2760 (N_2760,N_2653,N_2688);
xnor U2761 (N_2761,N_2682,N_2699);
and U2762 (N_2762,N_2658,N_2645);
and U2763 (N_2763,N_2631,N_2687);
or U2764 (N_2764,N_2688,N_2667);
or U2765 (N_2765,N_2663,N_2686);
or U2766 (N_2766,N_2671,N_2699);
nor U2767 (N_2767,N_2699,N_2626);
or U2768 (N_2768,N_2650,N_2639);
nor U2769 (N_2769,N_2693,N_2635);
and U2770 (N_2770,N_2698,N_2699);
nor U2771 (N_2771,N_2630,N_2683);
nor U2772 (N_2772,N_2661,N_2699);
nand U2773 (N_2773,N_2669,N_2664);
or U2774 (N_2774,N_2671,N_2698);
or U2775 (N_2775,N_2711,N_2739);
or U2776 (N_2776,N_2755,N_2762);
nand U2777 (N_2777,N_2717,N_2727);
and U2778 (N_2778,N_2761,N_2771);
nor U2779 (N_2779,N_2700,N_2760);
nand U2780 (N_2780,N_2730,N_2733);
nor U2781 (N_2781,N_2713,N_2742);
or U2782 (N_2782,N_2712,N_2704);
nor U2783 (N_2783,N_2701,N_2763);
nor U2784 (N_2784,N_2767,N_2745);
or U2785 (N_2785,N_2766,N_2752);
and U2786 (N_2786,N_2715,N_2746);
nor U2787 (N_2787,N_2722,N_2721);
and U2788 (N_2788,N_2707,N_2747);
nor U2789 (N_2789,N_2719,N_2728);
or U2790 (N_2790,N_2726,N_2718);
or U2791 (N_2791,N_2765,N_2773);
nand U2792 (N_2792,N_2738,N_2736);
or U2793 (N_2793,N_2743,N_2768);
and U2794 (N_2794,N_2714,N_2729);
and U2795 (N_2795,N_2709,N_2725);
and U2796 (N_2796,N_2731,N_2750);
nor U2797 (N_2797,N_2757,N_2723);
or U2798 (N_2798,N_2749,N_2705);
nor U2799 (N_2799,N_2720,N_2748);
and U2800 (N_2800,N_2740,N_2758);
or U2801 (N_2801,N_2764,N_2741);
and U2802 (N_2802,N_2769,N_2702);
nand U2803 (N_2803,N_2732,N_2710);
or U2804 (N_2804,N_2756,N_2744);
nor U2805 (N_2805,N_2754,N_2770);
and U2806 (N_2806,N_2751,N_2774);
nand U2807 (N_2807,N_2703,N_2716);
and U2808 (N_2808,N_2759,N_2772);
or U2809 (N_2809,N_2735,N_2724);
and U2810 (N_2810,N_2706,N_2708);
xnor U2811 (N_2811,N_2737,N_2753);
or U2812 (N_2812,N_2734,N_2753);
and U2813 (N_2813,N_2748,N_2751);
nand U2814 (N_2814,N_2721,N_2745);
and U2815 (N_2815,N_2728,N_2716);
nand U2816 (N_2816,N_2762,N_2721);
nand U2817 (N_2817,N_2732,N_2702);
nand U2818 (N_2818,N_2746,N_2774);
or U2819 (N_2819,N_2754,N_2752);
nor U2820 (N_2820,N_2730,N_2749);
and U2821 (N_2821,N_2702,N_2707);
nor U2822 (N_2822,N_2770,N_2738);
and U2823 (N_2823,N_2710,N_2742);
and U2824 (N_2824,N_2735,N_2730);
and U2825 (N_2825,N_2734,N_2710);
and U2826 (N_2826,N_2707,N_2754);
nor U2827 (N_2827,N_2725,N_2739);
nand U2828 (N_2828,N_2756,N_2720);
nor U2829 (N_2829,N_2732,N_2773);
nor U2830 (N_2830,N_2731,N_2747);
and U2831 (N_2831,N_2735,N_2743);
and U2832 (N_2832,N_2732,N_2765);
nor U2833 (N_2833,N_2737,N_2707);
or U2834 (N_2834,N_2710,N_2721);
nor U2835 (N_2835,N_2773,N_2701);
and U2836 (N_2836,N_2770,N_2745);
nand U2837 (N_2837,N_2748,N_2736);
nor U2838 (N_2838,N_2769,N_2753);
and U2839 (N_2839,N_2762,N_2770);
nand U2840 (N_2840,N_2743,N_2745);
and U2841 (N_2841,N_2770,N_2729);
and U2842 (N_2842,N_2747,N_2758);
nand U2843 (N_2843,N_2760,N_2716);
nand U2844 (N_2844,N_2741,N_2737);
nor U2845 (N_2845,N_2720,N_2744);
nand U2846 (N_2846,N_2756,N_2755);
and U2847 (N_2847,N_2735,N_2701);
nor U2848 (N_2848,N_2755,N_2707);
nor U2849 (N_2849,N_2723,N_2744);
or U2850 (N_2850,N_2823,N_2829);
or U2851 (N_2851,N_2803,N_2791);
nand U2852 (N_2852,N_2783,N_2817);
nor U2853 (N_2853,N_2824,N_2849);
nand U2854 (N_2854,N_2848,N_2793);
or U2855 (N_2855,N_2790,N_2835);
and U2856 (N_2856,N_2812,N_2810);
or U2857 (N_2857,N_2775,N_2780);
or U2858 (N_2858,N_2779,N_2837);
nand U2859 (N_2859,N_2805,N_2834);
nor U2860 (N_2860,N_2797,N_2843);
nor U2861 (N_2861,N_2796,N_2832);
nand U2862 (N_2862,N_2836,N_2785);
nor U2863 (N_2863,N_2802,N_2815);
nor U2864 (N_2864,N_2818,N_2777);
nand U2865 (N_2865,N_2807,N_2813);
nand U2866 (N_2866,N_2821,N_2847);
nand U2867 (N_2867,N_2786,N_2830);
nor U2868 (N_2868,N_2822,N_2787);
and U2869 (N_2869,N_2789,N_2827);
or U2870 (N_2870,N_2808,N_2798);
or U2871 (N_2871,N_2811,N_2840);
nor U2872 (N_2872,N_2782,N_2831);
and U2873 (N_2873,N_2776,N_2804);
and U2874 (N_2874,N_2799,N_2795);
or U2875 (N_2875,N_2826,N_2844);
and U2876 (N_2876,N_2788,N_2838);
nor U2877 (N_2877,N_2839,N_2781);
xnor U2878 (N_2878,N_2828,N_2801);
nand U2879 (N_2879,N_2794,N_2806);
nand U2880 (N_2880,N_2841,N_2809);
and U2881 (N_2881,N_2825,N_2820);
xor U2882 (N_2882,N_2842,N_2833);
or U2883 (N_2883,N_2784,N_2800);
nand U2884 (N_2884,N_2819,N_2792);
nand U2885 (N_2885,N_2778,N_2816);
nor U2886 (N_2886,N_2814,N_2846);
nand U2887 (N_2887,N_2845,N_2776);
or U2888 (N_2888,N_2819,N_2782);
nor U2889 (N_2889,N_2788,N_2841);
and U2890 (N_2890,N_2796,N_2791);
nand U2891 (N_2891,N_2819,N_2848);
nand U2892 (N_2892,N_2779,N_2825);
nor U2893 (N_2893,N_2791,N_2809);
and U2894 (N_2894,N_2843,N_2824);
nor U2895 (N_2895,N_2805,N_2790);
and U2896 (N_2896,N_2816,N_2779);
and U2897 (N_2897,N_2815,N_2780);
nor U2898 (N_2898,N_2789,N_2793);
xnor U2899 (N_2899,N_2842,N_2810);
and U2900 (N_2900,N_2811,N_2814);
and U2901 (N_2901,N_2848,N_2828);
and U2902 (N_2902,N_2841,N_2816);
nor U2903 (N_2903,N_2807,N_2847);
and U2904 (N_2904,N_2788,N_2815);
nor U2905 (N_2905,N_2831,N_2816);
and U2906 (N_2906,N_2799,N_2828);
and U2907 (N_2907,N_2802,N_2784);
nand U2908 (N_2908,N_2828,N_2811);
nor U2909 (N_2909,N_2786,N_2825);
nor U2910 (N_2910,N_2819,N_2820);
nand U2911 (N_2911,N_2846,N_2796);
nand U2912 (N_2912,N_2805,N_2817);
nand U2913 (N_2913,N_2841,N_2823);
and U2914 (N_2914,N_2796,N_2783);
or U2915 (N_2915,N_2780,N_2806);
nor U2916 (N_2916,N_2822,N_2835);
or U2917 (N_2917,N_2841,N_2811);
or U2918 (N_2918,N_2812,N_2804);
nor U2919 (N_2919,N_2822,N_2826);
nand U2920 (N_2920,N_2797,N_2819);
or U2921 (N_2921,N_2801,N_2783);
nor U2922 (N_2922,N_2810,N_2776);
and U2923 (N_2923,N_2818,N_2785);
nand U2924 (N_2924,N_2776,N_2799);
nor U2925 (N_2925,N_2897,N_2853);
or U2926 (N_2926,N_2906,N_2864);
or U2927 (N_2927,N_2889,N_2901);
nand U2928 (N_2928,N_2871,N_2892);
nor U2929 (N_2929,N_2911,N_2865);
nand U2930 (N_2930,N_2859,N_2873);
and U2931 (N_2931,N_2887,N_2854);
nand U2932 (N_2932,N_2884,N_2880);
or U2933 (N_2933,N_2905,N_2885);
and U2934 (N_2934,N_2862,N_2891);
and U2935 (N_2935,N_2908,N_2850);
and U2936 (N_2936,N_2886,N_2895);
and U2937 (N_2937,N_2878,N_2876);
or U2938 (N_2938,N_2902,N_2910);
or U2939 (N_2939,N_2879,N_2867);
nor U2940 (N_2940,N_2909,N_2920);
nor U2941 (N_2941,N_2923,N_2877);
nor U2942 (N_2942,N_2907,N_2918);
or U2943 (N_2943,N_2851,N_2883);
nand U2944 (N_2944,N_2881,N_2852);
or U2945 (N_2945,N_2915,N_2916);
or U2946 (N_2946,N_2898,N_2857);
nand U2947 (N_2947,N_2890,N_2912);
or U2948 (N_2948,N_2888,N_2882);
nand U2949 (N_2949,N_2924,N_2913);
or U2950 (N_2950,N_2899,N_2858);
nand U2951 (N_2951,N_2903,N_2866);
nor U2952 (N_2952,N_2914,N_2863);
and U2953 (N_2953,N_2874,N_2872);
or U2954 (N_2954,N_2855,N_2875);
and U2955 (N_2955,N_2860,N_2900);
nor U2956 (N_2956,N_2917,N_2896);
nor U2957 (N_2957,N_2868,N_2922);
nor U2958 (N_2958,N_2921,N_2904);
and U2959 (N_2959,N_2893,N_2919);
and U2960 (N_2960,N_2869,N_2894);
and U2961 (N_2961,N_2870,N_2856);
or U2962 (N_2962,N_2861,N_2891);
nor U2963 (N_2963,N_2916,N_2880);
xor U2964 (N_2964,N_2910,N_2877);
and U2965 (N_2965,N_2865,N_2920);
or U2966 (N_2966,N_2909,N_2915);
nor U2967 (N_2967,N_2921,N_2882);
nor U2968 (N_2968,N_2902,N_2911);
and U2969 (N_2969,N_2863,N_2871);
or U2970 (N_2970,N_2861,N_2851);
nand U2971 (N_2971,N_2924,N_2917);
or U2972 (N_2972,N_2896,N_2903);
and U2973 (N_2973,N_2916,N_2920);
and U2974 (N_2974,N_2877,N_2874);
and U2975 (N_2975,N_2901,N_2912);
and U2976 (N_2976,N_2901,N_2856);
nor U2977 (N_2977,N_2853,N_2913);
xor U2978 (N_2978,N_2907,N_2908);
nor U2979 (N_2979,N_2870,N_2852);
and U2980 (N_2980,N_2924,N_2902);
or U2981 (N_2981,N_2860,N_2887);
or U2982 (N_2982,N_2923,N_2865);
or U2983 (N_2983,N_2885,N_2878);
and U2984 (N_2984,N_2906,N_2866);
nand U2985 (N_2985,N_2856,N_2894);
and U2986 (N_2986,N_2901,N_2892);
nand U2987 (N_2987,N_2898,N_2893);
nand U2988 (N_2988,N_2853,N_2886);
nor U2989 (N_2989,N_2882,N_2891);
nor U2990 (N_2990,N_2857,N_2854);
nor U2991 (N_2991,N_2889,N_2898);
nand U2992 (N_2992,N_2852,N_2867);
nand U2993 (N_2993,N_2861,N_2864);
nand U2994 (N_2994,N_2900,N_2912);
and U2995 (N_2995,N_2914,N_2852);
nand U2996 (N_2996,N_2854,N_2903);
or U2997 (N_2997,N_2862,N_2919);
nand U2998 (N_2998,N_2923,N_2893);
nand U2999 (N_2999,N_2904,N_2868);
nor UO_0 (O_0,N_2973,N_2949);
nor UO_1 (O_1,N_2976,N_2984);
and UO_2 (O_2,N_2946,N_2951);
nand UO_3 (O_3,N_2939,N_2966);
nand UO_4 (O_4,N_2947,N_2987);
or UO_5 (O_5,N_2959,N_2942);
and UO_6 (O_6,N_2982,N_2950);
nand UO_7 (O_7,N_2981,N_2992);
or UO_8 (O_8,N_2932,N_2979);
nor UO_9 (O_9,N_2988,N_2963);
and UO_10 (O_10,N_2971,N_2999);
nand UO_11 (O_11,N_2929,N_2926);
nor UO_12 (O_12,N_2927,N_2957);
or UO_13 (O_13,N_2980,N_2948);
or UO_14 (O_14,N_2965,N_2972);
or UO_15 (O_15,N_2993,N_2955);
nor UO_16 (O_16,N_2956,N_2938);
or UO_17 (O_17,N_2925,N_2936);
nor UO_18 (O_18,N_2995,N_2997);
nand UO_19 (O_19,N_2977,N_2934);
nand UO_20 (O_20,N_2969,N_2945);
nor UO_21 (O_21,N_2967,N_2935);
and UO_22 (O_22,N_2943,N_2989);
nor UO_23 (O_23,N_2928,N_2961);
and UO_24 (O_24,N_2937,N_2998);
or UO_25 (O_25,N_2964,N_2983);
or UO_26 (O_26,N_2931,N_2974);
nand UO_27 (O_27,N_2962,N_2953);
and UO_28 (O_28,N_2933,N_2960);
and UO_29 (O_29,N_2975,N_2991);
xnor UO_30 (O_30,N_2968,N_2958);
and UO_31 (O_31,N_2996,N_2954);
or UO_32 (O_32,N_2986,N_2970);
or UO_33 (O_33,N_2941,N_2985);
or UO_34 (O_34,N_2990,N_2940);
nor UO_35 (O_35,N_2978,N_2994);
nor UO_36 (O_36,N_2930,N_2952);
and UO_37 (O_37,N_2944,N_2993);
nor UO_38 (O_38,N_2992,N_2984);
nor UO_39 (O_39,N_2988,N_2937);
nand UO_40 (O_40,N_2964,N_2938);
and UO_41 (O_41,N_2974,N_2937);
or UO_42 (O_42,N_2988,N_2973);
and UO_43 (O_43,N_2994,N_2966);
or UO_44 (O_44,N_2971,N_2983);
nor UO_45 (O_45,N_2986,N_2953);
or UO_46 (O_46,N_2949,N_2964);
nor UO_47 (O_47,N_2979,N_2973);
nand UO_48 (O_48,N_2931,N_2959);
nand UO_49 (O_49,N_2980,N_2961);
nor UO_50 (O_50,N_2991,N_2962);
nand UO_51 (O_51,N_2955,N_2990);
and UO_52 (O_52,N_2973,N_2964);
and UO_53 (O_53,N_2947,N_2994);
nand UO_54 (O_54,N_2940,N_2998);
and UO_55 (O_55,N_2999,N_2977);
or UO_56 (O_56,N_2960,N_2945);
nor UO_57 (O_57,N_2949,N_2996);
and UO_58 (O_58,N_2947,N_2942);
and UO_59 (O_59,N_2947,N_2968);
and UO_60 (O_60,N_2964,N_2998);
or UO_61 (O_61,N_2991,N_2955);
nand UO_62 (O_62,N_2968,N_2960);
nor UO_63 (O_63,N_2927,N_2983);
nor UO_64 (O_64,N_2927,N_2950);
nor UO_65 (O_65,N_2981,N_2993);
nand UO_66 (O_66,N_2998,N_2992);
and UO_67 (O_67,N_2988,N_2943);
or UO_68 (O_68,N_2989,N_2971);
nor UO_69 (O_69,N_2955,N_2992);
nand UO_70 (O_70,N_2939,N_2983);
or UO_71 (O_71,N_2933,N_2982);
or UO_72 (O_72,N_2925,N_2976);
nor UO_73 (O_73,N_2962,N_2956);
and UO_74 (O_74,N_2956,N_2989);
nor UO_75 (O_75,N_2929,N_2943);
nand UO_76 (O_76,N_2930,N_2981);
nor UO_77 (O_77,N_2970,N_2985);
or UO_78 (O_78,N_2943,N_2946);
xor UO_79 (O_79,N_2992,N_2934);
or UO_80 (O_80,N_2948,N_2950);
nor UO_81 (O_81,N_2977,N_2986);
nand UO_82 (O_82,N_2945,N_2943);
nor UO_83 (O_83,N_2985,N_2975);
nor UO_84 (O_84,N_2989,N_2949);
or UO_85 (O_85,N_2969,N_2949);
or UO_86 (O_86,N_2989,N_2974);
nor UO_87 (O_87,N_2977,N_2961);
nand UO_88 (O_88,N_2931,N_2942);
nor UO_89 (O_89,N_2952,N_2936);
nor UO_90 (O_90,N_2940,N_2993);
nand UO_91 (O_91,N_2966,N_2968);
and UO_92 (O_92,N_2948,N_2984);
and UO_93 (O_93,N_2931,N_2984);
xor UO_94 (O_94,N_2981,N_2935);
nand UO_95 (O_95,N_2990,N_2985);
or UO_96 (O_96,N_2928,N_2985);
nor UO_97 (O_97,N_2973,N_2939);
nand UO_98 (O_98,N_2925,N_2989);
nand UO_99 (O_99,N_2963,N_2933);
and UO_100 (O_100,N_2989,N_2983);
or UO_101 (O_101,N_2948,N_2952);
nor UO_102 (O_102,N_2931,N_2977);
nand UO_103 (O_103,N_2961,N_2927);
nor UO_104 (O_104,N_2958,N_2983);
or UO_105 (O_105,N_2940,N_2930);
nor UO_106 (O_106,N_2976,N_2931);
nand UO_107 (O_107,N_2991,N_2945);
or UO_108 (O_108,N_2976,N_2944);
or UO_109 (O_109,N_2994,N_2931);
or UO_110 (O_110,N_2965,N_2994);
nand UO_111 (O_111,N_2937,N_2979);
nor UO_112 (O_112,N_2996,N_2974);
nand UO_113 (O_113,N_2983,N_2955);
or UO_114 (O_114,N_2995,N_2943);
nand UO_115 (O_115,N_2934,N_2989);
or UO_116 (O_116,N_2958,N_2981);
nor UO_117 (O_117,N_2981,N_2975);
and UO_118 (O_118,N_2930,N_2964);
nand UO_119 (O_119,N_2942,N_2985);
or UO_120 (O_120,N_2952,N_2977);
nand UO_121 (O_121,N_2939,N_2943);
nor UO_122 (O_122,N_2980,N_2947);
or UO_123 (O_123,N_2961,N_2949);
nor UO_124 (O_124,N_2927,N_2952);
nand UO_125 (O_125,N_2938,N_2928);
nor UO_126 (O_126,N_2927,N_2953);
nor UO_127 (O_127,N_2951,N_2939);
or UO_128 (O_128,N_2935,N_2947);
and UO_129 (O_129,N_2957,N_2951);
and UO_130 (O_130,N_2955,N_2926);
nor UO_131 (O_131,N_2965,N_2941);
nand UO_132 (O_132,N_2990,N_2966);
and UO_133 (O_133,N_2926,N_2940);
nand UO_134 (O_134,N_2965,N_2967);
or UO_135 (O_135,N_2959,N_2949);
or UO_136 (O_136,N_2965,N_2982);
or UO_137 (O_137,N_2956,N_2926);
and UO_138 (O_138,N_2999,N_2940);
nand UO_139 (O_139,N_2937,N_2961);
nand UO_140 (O_140,N_2957,N_2947);
or UO_141 (O_141,N_2948,N_2995);
or UO_142 (O_142,N_2952,N_2925);
and UO_143 (O_143,N_2960,N_2928);
nor UO_144 (O_144,N_2951,N_2963);
or UO_145 (O_145,N_2933,N_2949);
and UO_146 (O_146,N_2970,N_2954);
nor UO_147 (O_147,N_2999,N_2950);
nor UO_148 (O_148,N_2965,N_2958);
nor UO_149 (O_149,N_2982,N_2926);
nor UO_150 (O_150,N_2967,N_2977);
nand UO_151 (O_151,N_2970,N_2943);
nand UO_152 (O_152,N_2932,N_2994);
and UO_153 (O_153,N_2931,N_2964);
or UO_154 (O_154,N_2944,N_2966);
nor UO_155 (O_155,N_2948,N_2972);
and UO_156 (O_156,N_2940,N_2959);
or UO_157 (O_157,N_2995,N_2932);
nand UO_158 (O_158,N_2997,N_2960);
and UO_159 (O_159,N_2944,N_2967);
nor UO_160 (O_160,N_2997,N_2927);
nand UO_161 (O_161,N_2930,N_2995);
and UO_162 (O_162,N_2969,N_2950);
or UO_163 (O_163,N_2947,N_2938);
nand UO_164 (O_164,N_2994,N_2939);
nand UO_165 (O_165,N_2969,N_2937);
nand UO_166 (O_166,N_2994,N_2945);
nor UO_167 (O_167,N_2946,N_2995);
and UO_168 (O_168,N_2975,N_2994);
nor UO_169 (O_169,N_2936,N_2957);
nor UO_170 (O_170,N_2934,N_2959);
nand UO_171 (O_171,N_2995,N_2937);
nor UO_172 (O_172,N_2971,N_2985);
or UO_173 (O_173,N_2959,N_2943);
nand UO_174 (O_174,N_2978,N_2996);
nor UO_175 (O_175,N_2964,N_2952);
and UO_176 (O_176,N_2998,N_2941);
or UO_177 (O_177,N_2938,N_2941);
and UO_178 (O_178,N_2969,N_2948);
or UO_179 (O_179,N_2925,N_2962);
nand UO_180 (O_180,N_2957,N_2934);
nor UO_181 (O_181,N_2973,N_2938);
nor UO_182 (O_182,N_2973,N_2959);
nor UO_183 (O_183,N_2938,N_2983);
nand UO_184 (O_184,N_2928,N_2998);
or UO_185 (O_185,N_2952,N_2968);
or UO_186 (O_186,N_2944,N_2952);
or UO_187 (O_187,N_2962,N_2977);
nand UO_188 (O_188,N_2958,N_2978);
xor UO_189 (O_189,N_2953,N_2971);
or UO_190 (O_190,N_2978,N_2933);
nand UO_191 (O_191,N_2954,N_2957);
and UO_192 (O_192,N_2964,N_2956);
or UO_193 (O_193,N_2942,N_2999);
nor UO_194 (O_194,N_2952,N_2989);
nand UO_195 (O_195,N_2953,N_2980);
and UO_196 (O_196,N_2970,N_2988);
and UO_197 (O_197,N_2966,N_2963);
and UO_198 (O_198,N_2938,N_2988);
and UO_199 (O_199,N_2925,N_2998);
or UO_200 (O_200,N_2952,N_2960);
nor UO_201 (O_201,N_2961,N_2967);
and UO_202 (O_202,N_2928,N_2955);
and UO_203 (O_203,N_2975,N_2953);
or UO_204 (O_204,N_2974,N_2962);
nor UO_205 (O_205,N_2996,N_2927);
nand UO_206 (O_206,N_2969,N_2991);
nand UO_207 (O_207,N_2953,N_2958);
nor UO_208 (O_208,N_2987,N_2975);
nor UO_209 (O_209,N_2927,N_2977);
and UO_210 (O_210,N_2932,N_2933);
nand UO_211 (O_211,N_2932,N_2953);
nand UO_212 (O_212,N_2947,N_2970);
or UO_213 (O_213,N_2996,N_2960);
and UO_214 (O_214,N_2965,N_2962);
nor UO_215 (O_215,N_2961,N_2956);
or UO_216 (O_216,N_2966,N_2969);
nand UO_217 (O_217,N_2938,N_2966);
xnor UO_218 (O_218,N_2982,N_2927);
and UO_219 (O_219,N_2972,N_2997);
nor UO_220 (O_220,N_2980,N_2984);
or UO_221 (O_221,N_2941,N_2953);
nand UO_222 (O_222,N_2996,N_2975);
nor UO_223 (O_223,N_2971,N_2997);
nand UO_224 (O_224,N_2957,N_2949);
or UO_225 (O_225,N_2963,N_2952);
or UO_226 (O_226,N_2958,N_2962);
nand UO_227 (O_227,N_2950,N_2979);
or UO_228 (O_228,N_2930,N_2944);
nand UO_229 (O_229,N_2951,N_2992);
nor UO_230 (O_230,N_2927,N_2973);
and UO_231 (O_231,N_2951,N_2983);
or UO_232 (O_232,N_2940,N_2991);
nand UO_233 (O_233,N_2961,N_2990);
and UO_234 (O_234,N_2926,N_2952);
xor UO_235 (O_235,N_2925,N_2968);
or UO_236 (O_236,N_2957,N_2988);
nand UO_237 (O_237,N_2961,N_2983);
nand UO_238 (O_238,N_2939,N_2931);
nor UO_239 (O_239,N_2928,N_2999);
nor UO_240 (O_240,N_2997,N_2981);
nand UO_241 (O_241,N_2976,N_2981);
nor UO_242 (O_242,N_2933,N_2994);
nor UO_243 (O_243,N_2970,N_2951);
nor UO_244 (O_244,N_2972,N_2925);
and UO_245 (O_245,N_2964,N_2945);
and UO_246 (O_246,N_2963,N_2928);
nand UO_247 (O_247,N_2936,N_2965);
or UO_248 (O_248,N_2993,N_2973);
and UO_249 (O_249,N_2974,N_2927);
and UO_250 (O_250,N_2987,N_2968);
nor UO_251 (O_251,N_2955,N_2929);
nand UO_252 (O_252,N_2993,N_2988);
or UO_253 (O_253,N_2995,N_2962);
or UO_254 (O_254,N_2961,N_2992);
and UO_255 (O_255,N_2928,N_2967);
nor UO_256 (O_256,N_2936,N_2972);
and UO_257 (O_257,N_2942,N_2938);
nand UO_258 (O_258,N_2950,N_2932);
and UO_259 (O_259,N_2962,N_2997);
or UO_260 (O_260,N_2939,N_2934);
and UO_261 (O_261,N_2969,N_2982);
nor UO_262 (O_262,N_2958,N_2932);
and UO_263 (O_263,N_2949,N_2956);
or UO_264 (O_264,N_2993,N_2971);
and UO_265 (O_265,N_2972,N_2939);
or UO_266 (O_266,N_2977,N_2933);
or UO_267 (O_267,N_2983,N_2982);
nor UO_268 (O_268,N_2936,N_2976);
or UO_269 (O_269,N_2969,N_2984);
nor UO_270 (O_270,N_2981,N_2956);
or UO_271 (O_271,N_2979,N_2938);
nor UO_272 (O_272,N_2948,N_2979);
or UO_273 (O_273,N_2949,N_2941);
or UO_274 (O_274,N_2986,N_2969);
nor UO_275 (O_275,N_2954,N_2949);
or UO_276 (O_276,N_2927,N_2946);
nor UO_277 (O_277,N_2955,N_2975);
or UO_278 (O_278,N_2978,N_2951);
and UO_279 (O_279,N_2938,N_2950);
and UO_280 (O_280,N_2925,N_2940);
and UO_281 (O_281,N_2995,N_2941);
nor UO_282 (O_282,N_2980,N_2974);
nand UO_283 (O_283,N_2952,N_2950);
or UO_284 (O_284,N_2963,N_2950);
nor UO_285 (O_285,N_2939,N_2958);
or UO_286 (O_286,N_2976,N_2979);
nor UO_287 (O_287,N_2997,N_2937);
nor UO_288 (O_288,N_2976,N_2977);
or UO_289 (O_289,N_2975,N_2963);
nor UO_290 (O_290,N_2968,N_2943);
or UO_291 (O_291,N_2983,N_2975);
or UO_292 (O_292,N_2965,N_2979);
and UO_293 (O_293,N_2931,N_2993);
and UO_294 (O_294,N_2943,N_2951);
nor UO_295 (O_295,N_2965,N_2957);
nand UO_296 (O_296,N_2982,N_2937);
or UO_297 (O_297,N_2995,N_2935);
nor UO_298 (O_298,N_2986,N_2937);
nor UO_299 (O_299,N_2968,N_2944);
nor UO_300 (O_300,N_2935,N_2962);
nand UO_301 (O_301,N_2932,N_2997);
and UO_302 (O_302,N_2961,N_2968);
and UO_303 (O_303,N_2929,N_2991);
nand UO_304 (O_304,N_2996,N_2952);
nor UO_305 (O_305,N_2964,N_2968);
or UO_306 (O_306,N_2999,N_2927);
and UO_307 (O_307,N_2990,N_2975);
nand UO_308 (O_308,N_2933,N_2984);
or UO_309 (O_309,N_2970,N_2968);
or UO_310 (O_310,N_2931,N_2951);
or UO_311 (O_311,N_2991,N_2932);
nand UO_312 (O_312,N_2974,N_2987);
nor UO_313 (O_313,N_2931,N_2981);
or UO_314 (O_314,N_2985,N_2967);
nor UO_315 (O_315,N_2998,N_2950);
or UO_316 (O_316,N_2972,N_2969);
or UO_317 (O_317,N_2976,N_2935);
nand UO_318 (O_318,N_2989,N_2969);
or UO_319 (O_319,N_2976,N_2968);
nor UO_320 (O_320,N_2985,N_2962);
or UO_321 (O_321,N_2943,N_2971);
nand UO_322 (O_322,N_2996,N_2935);
nor UO_323 (O_323,N_2970,N_2926);
or UO_324 (O_324,N_2980,N_2986);
or UO_325 (O_325,N_2997,N_2948);
and UO_326 (O_326,N_2999,N_2947);
and UO_327 (O_327,N_2947,N_2974);
nor UO_328 (O_328,N_2982,N_2941);
and UO_329 (O_329,N_2927,N_2968);
or UO_330 (O_330,N_2966,N_2970);
nor UO_331 (O_331,N_2927,N_2992);
nor UO_332 (O_332,N_2948,N_2946);
nor UO_333 (O_333,N_2961,N_2955);
and UO_334 (O_334,N_2980,N_2997);
or UO_335 (O_335,N_2979,N_2994);
and UO_336 (O_336,N_2932,N_2976);
or UO_337 (O_337,N_2937,N_2996);
or UO_338 (O_338,N_2967,N_2953);
and UO_339 (O_339,N_2988,N_2979);
xnor UO_340 (O_340,N_2943,N_2991);
or UO_341 (O_341,N_2942,N_2955);
nand UO_342 (O_342,N_2958,N_2975);
or UO_343 (O_343,N_2972,N_2982);
or UO_344 (O_344,N_2939,N_2956);
nand UO_345 (O_345,N_2955,N_2979);
nand UO_346 (O_346,N_2993,N_2938);
xnor UO_347 (O_347,N_2951,N_2956);
nand UO_348 (O_348,N_2938,N_2929);
nand UO_349 (O_349,N_2948,N_2982);
nor UO_350 (O_350,N_2979,N_2991);
nor UO_351 (O_351,N_2929,N_2994);
or UO_352 (O_352,N_2926,N_2935);
nor UO_353 (O_353,N_2988,N_2969);
nor UO_354 (O_354,N_2982,N_2954);
nand UO_355 (O_355,N_2967,N_2955);
nor UO_356 (O_356,N_2968,N_2926);
nor UO_357 (O_357,N_2981,N_2929);
and UO_358 (O_358,N_2944,N_2991);
and UO_359 (O_359,N_2995,N_2988);
nor UO_360 (O_360,N_2929,N_2977);
or UO_361 (O_361,N_2976,N_2954);
nand UO_362 (O_362,N_2927,N_2981);
or UO_363 (O_363,N_2945,N_2961);
or UO_364 (O_364,N_2926,N_2986);
nor UO_365 (O_365,N_2982,N_2947);
nor UO_366 (O_366,N_2975,N_2967);
nor UO_367 (O_367,N_2965,N_2960);
and UO_368 (O_368,N_2995,N_2949);
nand UO_369 (O_369,N_2933,N_2954);
and UO_370 (O_370,N_2995,N_2973);
nand UO_371 (O_371,N_2948,N_2965);
nand UO_372 (O_372,N_2942,N_2925);
or UO_373 (O_373,N_2928,N_2952);
nand UO_374 (O_374,N_2947,N_2984);
nor UO_375 (O_375,N_2938,N_2951);
or UO_376 (O_376,N_2985,N_2957);
nor UO_377 (O_377,N_2963,N_2938);
nor UO_378 (O_378,N_2976,N_2973);
nor UO_379 (O_379,N_2988,N_2935);
nor UO_380 (O_380,N_2945,N_2993);
nor UO_381 (O_381,N_2972,N_2955);
or UO_382 (O_382,N_2947,N_2995);
or UO_383 (O_383,N_2992,N_2958);
nand UO_384 (O_384,N_2962,N_2946);
nand UO_385 (O_385,N_2995,N_2970);
or UO_386 (O_386,N_2987,N_2945);
nand UO_387 (O_387,N_2966,N_2945);
and UO_388 (O_388,N_2940,N_2948);
or UO_389 (O_389,N_2964,N_2937);
nor UO_390 (O_390,N_2991,N_2933);
or UO_391 (O_391,N_2991,N_2967);
xnor UO_392 (O_392,N_2961,N_2998);
nor UO_393 (O_393,N_2941,N_2935);
or UO_394 (O_394,N_2994,N_2983);
and UO_395 (O_395,N_2975,N_2970);
nor UO_396 (O_396,N_2977,N_2928);
nand UO_397 (O_397,N_2968,N_2951);
or UO_398 (O_398,N_2939,N_2993);
and UO_399 (O_399,N_2984,N_2953);
nand UO_400 (O_400,N_2961,N_2995);
and UO_401 (O_401,N_2929,N_2985);
or UO_402 (O_402,N_2973,N_2956);
or UO_403 (O_403,N_2985,N_2995);
or UO_404 (O_404,N_2999,N_2936);
and UO_405 (O_405,N_2985,N_2961);
and UO_406 (O_406,N_2949,N_2953);
or UO_407 (O_407,N_2934,N_2967);
or UO_408 (O_408,N_2974,N_2958);
nand UO_409 (O_409,N_2931,N_2943);
nand UO_410 (O_410,N_2954,N_2950);
nand UO_411 (O_411,N_2998,N_2932);
or UO_412 (O_412,N_2927,N_2972);
and UO_413 (O_413,N_2985,N_2969);
nor UO_414 (O_414,N_2950,N_2990);
or UO_415 (O_415,N_2949,N_2978);
and UO_416 (O_416,N_2966,N_2962);
or UO_417 (O_417,N_2998,N_2977);
nand UO_418 (O_418,N_2937,N_2976);
or UO_419 (O_419,N_2925,N_2985);
or UO_420 (O_420,N_2966,N_2947);
or UO_421 (O_421,N_2956,N_2942);
or UO_422 (O_422,N_2950,N_2926);
and UO_423 (O_423,N_2942,N_2954);
and UO_424 (O_424,N_2979,N_2978);
or UO_425 (O_425,N_2981,N_2950);
or UO_426 (O_426,N_2930,N_2951);
nor UO_427 (O_427,N_2947,N_2962);
nor UO_428 (O_428,N_2934,N_2930);
and UO_429 (O_429,N_2976,N_2963);
and UO_430 (O_430,N_2937,N_2941);
nor UO_431 (O_431,N_2967,N_2945);
xnor UO_432 (O_432,N_2951,N_2971);
and UO_433 (O_433,N_2961,N_2973);
nor UO_434 (O_434,N_2974,N_2956);
xnor UO_435 (O_435,N_2955,N_2982);
or UO_436 (O_436,N_2951,N_2993);
nand UO_437 (O_437,N_2962,N_2964);
nand UO_438 (O_438,N_2970,N_2939);
and UO_439 (O_439,N_2998,N_2962);
nand UO_440 (O_440,N_2939,N_2945);
nor UO_441 (O_441,N_2992,N_2935);
and UO_442 (O_442,N_2972,N_2996);
and UO_443 (O_443,N_2994,N_2969);
or UO_444 (O_444,N_2958,N_2951);
and UO_445 (O_445,N_2982,N_2968);
nand UO_446 (O_446,N_2980,N_2995);
and UO_447 (O_447,N_2977,N_2964);
nor UO_448 (O_448,N_2963,N_2936);
or UO_449 (O_449,N_2950,N_2940);
nand UO_450 (O_450,N_2934,N_2991);
nand UO_451 (O_451,N_2929,N_2975);
and UO_452 (O_452,N_2972,N_2929);
nand UO_453 (O_453,N_2980,N_2965);
nand UO_454 (O_454,N_2947,N_2934);
or UO_455 (O_455,N_2970,N_2932);
and UO_456 (O_456,N_2944,N_2961);
nor UO_457 (O_457,N_2941,N_2928);
or UO_458 (O_458,N_2934,N_2929);
or UO_459 (O_459,N_2997,N_2938);
or UO_460 (O_460,N_2954,N_2981);
nand UO_461 (O_461,N_2948,N_2941);
and UO_462 (O_462,N_2967,N_2997);
and UO_463 (O_463,N_2972,N_2954);
or UO_464 (O_464,N_2992,N_2964);
nor UO_465 (O_465,N_2967,N_2999);
nand UO_466 (O_466,N_2960,N_2964);
nand UO_467 (O_467,N_2989,N_2950);
nor UO_468 (O_468,N_2991,N_2972);
nand UO_469 (O_469,N_2941,N_2934);
nand UO_470 (O_470,N_2929,N_2939);
nand UO_471 (O_471,N_2937,N_2952);
or UO_472 (O_472,N_2959,N_2925);
nor UO_473 (O_473,N_2957,N_2945);
nor UO_474 (O_474,N_2929,N_2999);
nor UO_475 (O_475,N_2970,N_2967);
or UO_476 (O_476,N_2958,N_2957);
or UO_477 (O_477,N_2949,N_2976);
xnor UO_478 (O_478,N_2996,N_2925);
or UO_479 (O_479,N_2985,N_2996);
nor UO_480 (O_480,N_2973,N_2980);
or UO_481 (O_481,N_2930,N_2987);
nor UO_482 (O_482,N_2949,N_2993);
or UO_483 (O_483,N_2981,N_2946);
and UO_484 (O_484,N_2999,N_2965);
and UO_485 (O_485,N_2952,N_2957);
nand UO_486 (O_486,N_2981,N_2942);
and UO_487 (O_487,N_2990,N_2982);
nand UO_488 (O_488,N_2926,N_2965);
and UO_489 (O_489,N_2964,N_2957);
and UO_490 (O_490,N_2934,N_2943);
or UO_491 (O_491,N_2955,N_2927);
and UO_492 (O_492,N_2970,N_2955);
nand UO_493 (O_493,N_2969,N_2981);
and UO_494 (O_494,N_2979,N_2939);
or UO_495 (O_495,N_2931,N_2985);
nor UO_496 (O_496,N_2995,N_2945);
nand UO_497 (O_497,N_2936,N_2954);
or UO_498 (O_498,N_2973,N_2942);
nand UO_499 (O_499,N_2929,N_2947);
endmodule