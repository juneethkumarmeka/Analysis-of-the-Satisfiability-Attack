module basic_1500_15000_2000_15_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_1407,In_1017);
or U1 (N_1,In_685,In_601);
xor U2 (N_2,In_737,In_1287);
and U3 (N_3,In_542,In_223);
and U4 (N_4,In_185,In_1128);
xnor U5 (N_5,In_956,In_1162);
xor U6 (N_6,In_1003,In_1144);
nand U7 (N_7,In_929,In_372);
and U8 (N_8,In_350,In_919);
nor U9 (N_9,In_1153,In_1220);
nand U10 (N_10,In_404,In_139);
nor U11 (N_11,In_1120,In_460);
nand U12 (N_12,In_876,In_409);
nor U13 (N_13,In_67,In_498);
and U14 (N_14,In_782,In_1458);
and U15 (N_15,In_529,In_671);
nor U16 (N_16,In_1160,In_1404);
nor U17 (N_17,In_68,In_1078);
nor U18 (N_18,In_1256,In_94);
or U19 (N_19,In_1300,In_444);
xor U20 (N_20,In_699,In_805);
nand U21 (N_21,In_1035,In_286);
and U22 (N_22,In_377,In_1400);
and U23 (N_23,In_518,In_809);
and U24 (N_24,In_622,In_183);
and U25 (N_25,In_423,In_279);
nor U26 (N_26,In_694,In_1413);
nand U27 (N_27,In_134,In_207);
or U28 (N_28,In_989,In_1224);
nand U29 (N_29,In_927,In_1206);
or U30 (N_30,In_554,In_90);
xor U31 (N_31,In_142,In_1124);
and U32 (N_32,In_1317,In_294);
nand U33 (N_33,In_274,In_254);
or U34 (N_34,In_718,In_1350);
nor U35 (N_35,In_1323,In_722);
or U36 (N_36,In_1345,In_552);
nand U37 (N_37,In_890,In_1043);
xor U38 (N_38,In_878,In_625);
xnor U39 (N_39,In_315,In_1092);
nand U40 (N_40,In_468,In_517);
and U41 (N_41,In_131,In_482);
nand U42 (N_42,In_193,In_1408);
xor U43 (N_43,In_1422,In_874);
nand U44 (N_44,In_644,In_893);
or U45 (N_45,In_1490,In_609);
or U46 (N_46,In_222,In_786);
xnor U47 (N_47,In_287,In_435);
or U48 (N_48,In_1339,In_1188);
xnor U49 (N_49,In_1100,In_985);
and U50 (N_50,In_769,In_150);
nor U51 (N_51,In_706,In_758);
xor U52 (N_52,In_0,In_633);
nand U53 (N_53,In_60,In_1429);
or U54 (N_54,In_302,In_1455);
and U55 (N_55,In_485,In_1045);
or U56 (N_56,In_1143,In_1320);
and U57 (N_57,In_353,In_797);
and U58 (N_58,In_1231,In_1298);
or U59 (N_59,In_472,In_865);
or U60 (N_60,In_474,In_702);
xor U61 (N_61,In_708,In_417);
and U62 (N_62,In_1204,In_1151);
nor U63 (N_63,In_1122,In_1000);
and U64 (N_64,In_749,In_750);
nand U65 (N_65,In_261,In_78);
nor U66 (N_66,In_584,In_1068);
and U67 (N_67,In_1084,In_31);
nor U68 (N_68,In_788,In_1251);
xor U69 (N_69,In_1411,In_692);
and U70 (N_70,In_1216,In_469);
nand U71 (N_71,In_546,In_301);
and U72 (N_72,In_1129,In_1386);
or U73 (N_73,In_1001,In_1343);
nand U74 (N_74,In_103,In_1174);
xnor U75 (N_75,In_1460,In_130);
or U76 (N_76,In_647,In_457);
xor U77 (N_77,In_1240,In_292);
xnor U78 (N_78,In_607,In_320);
nand U79 (N_79,In_276,In_716);
and U80 (N_80,In_351,In_1493);
nand U81 (N_81,In_1178,In_1089);
nor U82 (N_82,In_1452,In_132);
nor U83 (N_83,In_145,In_58);
nor U84 (N_84,In_566,In_977);
or U85 (N_85,In_1448,In_511);
nand U86 (N_86,In_1098,In_871);
nor U87 (N_87,In_1402,In_1192);
nor U88 (N_88,In_1182,In_323);
or U89 (N_89,In_401,In_1197);
or U90 (N_90,In_75,In_1239);
xnor U91 (N_91,In_211,In_1180);
xnor U92 (N_92,In_1468,In_925);
xnor U93 (N_93,In_1279,In_955);
nor U94 (N_94,In_523,In_1465);
and U95 (N_95,In_376,In_663);
nor U96 (N_96,In_459,In_1449);
xor U97 (N_97,In_793,In_338);
xnor U98 (N_98,In_214,In_1042);
nand U99 (N_99,In_932,In_1288);
or U100 (N_100,In_105,In_611);
nor U101 (N_101,In_1166,In_1241);
nand U102 (N_102,In_819,In_1269);
xor U103 (N_103,In_1119,In_1027);
nor U104 (N_104,In_1156,In_1070);
nand U105 (N_105,In_966,In_1275);
nor U106 (N_106,In_82,In_504);
or U107 (N_107,In_220,In_668);
nand U108 (N_108,In_466,In_532);
nor U109 (N_109,In_486,In_964);
nand U110 (N_110,In_670,In_1387);
nor U111 (N_111,In_698,In_1041);
xnor U112 (N_112,In_133,In_1342);
nand U113 (N_113,In_38,In_244);
nor U114 (N_114,In_569,In_135);
nor U115 (N_115,In_76,In_767);
and U116 (N_116,In_1095,In_202);
xor U117 (N_117,In_186,In_1196);
xor U118 (N_118,In_648,In_125);
nand U119 (N_119,In_1135,In_352);
and U120 (N_120,In_791,In_1483);
nand U121 (N_121,In_218,In_1372);
nor U122 (N_122,In_641,In_73);
and U123 (N_123,In_495,In_1218);
nand U124 (N_124,In_386,In_55);
nor U125 (N_125,In_728,In_715);
and U126 (N_126,In_796,In_1481);
or U127 (N_127,In_157,In_575);
or U128 (N_128,In_1217,In_1243);
and U129 (N_129,In_201,In_1295);
or U130 (N_130,In_934,In_208);
nor U131 (N_131,In_226,In_93);
nand U132 (N_132,In_683,In_762);
nand U133 (N_133,In_121,In_70);
nand U134 (N_134,In_826,In_424);
and U135 (N_135,In_790,In_59);
nor U136 (N_136,In_574,In_210);
nand U137 (N_137,In_148,In_399);
xnor U138 (N_138,In_1333,In_3);
and U139 (N_139,In_727,In_988);
xnor U140 (N_140,In_316,In_608);
or U141 (N_141,In_561,In_996);
nor U142 (N_142,In_820,In_421);
and U143 (N_143,In_992,In_751);
or U144 (N_144,In_428,In_1139);
nand U145 (N_145,In_1112,In_658);
nand U146 (N_146,In_1430,In_258);
and U147 (N_147,In_1497,In_322);
and U148 (N_148,In_1071,In_490);
or U149 (N_149,In_414,In_475);
nor U150 (N_150,In_1055,In_1207);
nor U151 (N_151,In_115,In_1393);
and U152 (N_152,In_308,In_1008);
nor U153 (N_153,In_438,In_593);
and U154 (N_154,In_736,In_1346);
nor U155 (N_155,In_288,In_898);
xnor U156 (N_156,In_242,In_605);
xor U157 (N_157,In_571,In_524);
nand U158 (N_158,In_373,In_233);
or U159 (N_159,In_84,In_311);
and U160 (N_160,In_74,In_666);
nor U161 (N_161,In_408,In_1443);
nor U162 (N_162,In_448,In_1337);
nor U163 (N_163,In_1155,In_1395);
xnor U164 (N_164,In_332,In_1439);
and U165 (N_165,In_206,In_61);
xnor U166 (N_166,In_418,In_1470);
nor U167 (N_167,In_1210,In_422);
and U168 (N_168,In_953,In_682);
xnor U169 (N_169,In_230,In_381);
or U170 (N_170,In_531,In_99);
and U171 (N_171,In_429,In_1396);
nand U172 (N_172,In_167,In_1421);
or U173 (N_173,In_975,In_931);
or U174 (N_174,In_978,In_283);
or U175 (N_175,In_328,In_33);
or U176 (N_176,In_689,In_369);
nor U177 (N_177,In_23,In_392);
or U178 (N_178,In_873,In_1399);
and U179 (N_179,In_540,In_164);
or U180 (N_180,In_492,In_817);
and U181 (N_181,In_774,In_655);
nand U182 (N_182,In_808,In_1423);
and U183 (N_183,In_861,In_825);
nor U184 (N_184,In_544,In_360);
or U185 (N_185,In_1260,In_1356);
and U186 (N_186,In_57,In_535);
xnor U187 (N_187,In_949,In_366);
nor U188 (N_188,In_1134,In_772);
and U189 (N_189,In_519,In_251);
or U190 (N_190,In_789,In_1115);
or U191 (N_191,In_897,In_397);
and U192 (N_192,In_1307,In_645);
nand U193 (N_193,In_1173,In_522);
nor U194 (N_194,In_631,In_7);
or U195 (N_195,In_1037,In_509);
nor U196 (N_196,In_1132,In_1082);
and U197 (N_197,In_1103,In_1185);
or U198 (N_198,In_1164,In_1097);
xnor U199 (N_199,In_1163,In_488);
xor U200 (N_200,In_91,In_1059);
and U201 (N_201,In_1363,In_229);
or U202 (N_202,In_180,In_738);
nor U203 (N_203,In_792,In_604);
and U204 (N_204,In_1004,In_613);
and U205 (N_205,In_1187,In_1499);
xnor U206 (N_206,In_1314,In_795);
xor U207 (N_207,In_358,In_1085);
nor U208 (N_208,In_650,In_143);
nor U209 (N_209,In_52,In_500);
and U210 (N_210,In_962,In_1427);
nor U211 (N_211,In_231,In_415);
and U212 (N_212,In_553,In_541);
and U213 (N_213,In_36,In_635);
or U214 (N_214,In_732,In_506);
nand U215 (N_215,In_14,In_69);
xor U216 (N_216,In_963,In_1259);
nand U217 (N_217,In_1347,In_1158);
or U218 (N_218,In_907,In_467);
or U219 (N_219,In_43,In_269);
nor U220 (N_220,In_1226,In_773);
nand U221 (N_221,In_307,In_759);
and U222 (N_222,In_119,In_1113);
and U223 (N_223,In_860,In_654);
nor U224 (N_224,In_113,In_990);
or U225 (N_225,In_854,In_1102);
nand U226 (N_226,In_83,In_866);
nor U227 (N_227,In_1437,In_1147);
nor U228 (N_228,In_1238,In_238);
and U229 (N_229,In_1385,In_859);
or U230 (N_230,In_562,In_551);
and U231 (N_231,In_305,In_1273);
nor U232 (N_232,In_1294,In_1235);
xnor U233 (N_233,In_1203,In_98);
and U234 (N_234,In_623,In_1077);
xor U235 (N_235,In_304,In_799);
nor U236 (N_236,In_361,In_1332);
or U237 (N_237,In_1368,In_205);
nand U238 (N_238,In_1149,In_179);
and U239 (N_239,In_638,In_109);
or U240 (N_240,In_20,In_754);
and U241 (N_241,In_1029,In_255);
nand U242 (N_242,In_363,In_282);
nor U243 (N_243,In_944,In_124);
or U244 (N_244,In_1334,In_80);
nor U245 (N_245,In_1378,In_291);
and U246 (N_246,In_1123,In_1431);
xnor U247 (N_247,In_537,In_162);
nor U248 (N_248,In_382,In_1398);
nor U249 (N_249,In_15,In_1244);
nand U250 (N_250,In_849,In_266);
xnor U251 (N_251,In_107,In_602);
nand U252 (N_252,In_434,In_200);
or U253 (N_253,In_168,In_1117);
and U254 (N_254,In_97,In_51);
and U255 (N_255,In_169,In_171);
nor U256 (N_256,In_921,In_1140);
or U257 (N_257,In_875,In_1108);
and U258 (N_258,In_526,In_431);
xnor U259 (N_259,In_595,In_812);
nand U260 (N_260,In_550,In_1401);
and U261 (N_261,In_1321,In_123);
nand U262 (N_262,In_1436,In_1303);
nor U263 (N_263,In_1280,In_111);
or U264 (N_264,In_165,In_1488);
nand U265 (N_265,In_273,In_775);
or U266 (N_266,In_995,In_646);
xor U267 (N_267,In_1127,In_649);
and U268 (N_268,In_1405,In_126);
xor U269 (N_269,In_748,In_1195);
nor U270 (N_270,In_661,In_471);
and U271 (N_271,In_1109,In_400);
nor U272 (N_272,In_1193,In_112);
or U273 (N_273,In_462,In_1199);
nor U274 (N_274,In_1383,In_1270);
nor U275 (N_275,In_1019,In_629);
nand U276 (N_276,In_798,In_1489);
or U277 (N_277,In_359,In_979);
nand U278 (N_278,In_1394,In_1425);
nor U279 (N_279,In_880,In_1258);
xor U280 (N_280,In_600,In_1130);
and U281 (N_281,In_513,In_343);
nor U282 (N_282,In_810,In_712);
nand U283 (N_283,In_704,In_711);
nor U284 (N_284,In_879,In_1491);
or U285 (N_285,In_1271,In_855);
or U286 (N_286,In_686,In_505);
nand U287 (N_287,In_1311,In_79);
or U288 (N_288,In_981,In_733);
xor U289 (N_289,In_1286,In_140);
and U290 (N_290,In_437,In_888);
nor U291 (N_291,In_263,In_1110);
nand U292 (N_292,In_306,In_297);
nor U293 (N_293,In_664,In_656);
xor U294 (N_294,In_1444,In_657);
nand U295 (N_295,In_16,In_1340);
or U296 (N_296,In_1229,In_912);
nor U297 (N_297,In_224,In_724);
xnor U298 (N_298,In_1415,In_512);
nand U299 (N_299,In_936,In_533);
nor U300 (N_300,In_1292,In_585);
xnor U301 (N_301,In_1291,In_195);
nor U302 (N_302,In_289,In_354);
xnor U303 (N_303,In_807,In_1200);
and U304 (N_304,In_507,In_998);
nor U305 (N_305,In_10,In_449);
or U306 (N_306,In_259,In_1360);
nand U307 (N_307,In_1322,In_25);
or U308 (N_308,In_1018,In_1324);
xor U309 (N_309,In_1107,In_1028);
nand U310 (N_310,In_1086,In_327);
and U311 (N_311,In_440,In_939);
or U312 (N_312,In_906,In_675);
nor U313 (N_313,In_345,In_917);
and U314 (N_314,In_29,In_1299);
nand U315 (N_315,In_760,In_1066);
nand U316 (N_316,In_563,In_892);
nor U317 (N_317,In_872,In_252);
nand U318 (N_318,In_539,In_735);
and U319 (N_319,In_521,In_1484);
or U320 (N_320,In_86,In_740);
or U321 (N_321,In_1148,In_101);
nand U322 (N_322,In_624,In_1305);
xnor U323 (N_323,In_869,In_267);
xnor U324 (N_324,In_862,In_1276);
or U325 (N_325,In_1169,In_1450);
nand U326 (N_326,In_1114,In_24);
xor U327 (N_327,In_146,In_1362);
nand U328 (N_328,In_298,In_783);
nand U329 (N_329,In_309,In_1464);
and U330 (N_330,In_175,In_1354);
or U331 (N_331,In_480,In_1426);
nor U332 (N_332,In_12,In_1096);
nand U333 (N_333,In_1225,In_1289);
nand U334 (N_334,In_1494,In_705);
and U335 (N_335,In_1278,In_946);
xor U336 (N_336,In_347,In_1133);
xor U337 (N_337,In_1482,In_284);
xor U338 (N_338,In_821,In_940);
nand U339 (N_339,In_6,In_779);
nand U340 (N_340,In_451,In_1016);
nand U341 (N_341,In_314,In_831);
and U342 (N_342,In_824,In_1104);
or U343 (N_343,In_761,In_1403);
nand U344 (N_344,In_1463,In_1351);
xor U345 (N_345,In_1414,In_497);
and U346 (N_346,In_272,In_1061);
nor U347 (N_347,In_1283,In_555);
and U348 (N_348,In_547,In_194);
and U349 (N_349,In_1369,In_384);
nor U350 (N_350,In_768,In_110);
and U351 (N_351,In_695,In_643);
and U352 (N_352,In_225,In_234);
xor U353 (N_353,In_1296,In_356);
nand U354 (N_354,In_548,In_954);
nand U355 (N_355,In_221,In_752);
nand U356 (N_356,In_590,In_281);
or U357 (N_357,In_494,In_703);
and U358 (N_358,In_1285,In_1247);
and U359 (N_359,In_127,In_1492);
xnor U360 (N_360,In_22,In_395);
nor U361 (N_361,In_719,In_501);
and U362 (N_362,In_994,In_1433);
or U363 (N_363,In_1047,In_577);
nor U364 (N_364,In_161,In_586);
or U365 (N_365,In_318,In_1485);
xnor U366 (N_366,In_958,In_867);
or U367 (N_367,In_1230,In_1141);
or U368 (N_368,In_1032,In_1391);
or U369 (N_369,In_673,In_388);
nand U370 (N_370,In_1462,In_581);
xnor U371 (N_371,In_1063,In_49);
or U372 (N_372,In_803,In_1126);
or U373 (N_373,In_1222,In_340);
nor U374 (N_374,In_1376,In_1441);
or U375 (N_375,In_357,In_355);
and U376 (N_376,In_972,In_1076);
or U377 (N_377,In_784,In_178);
xnor U378 (N_378,In_745,In_1219);
or U379 (N_379,In_1212,In_443);
or U380 (N_380,In_730,In_834);
and U381 (N_381,In_1025,In_1268);
or U382 (N_382,In_1424,In_822);
and U383 (N_383,In_326,In_1262);
xor U384 (N_384,In_312,In_572);
nand U385 (N_385,In_1390,In_1355);
nor U386 (N_386,In_374,In_1293);
and U387 (N_387,In_957,In_1125);
or U388 (N_388,In_1131,In_811);
or U389 (N_389,In_344,In_842);
nor U390 (N_390,In_528,In_910);
and U391 (N_391,In_741,In_235);
and U392 (N_392,In_589,In_1384);
nor U393 (N_393,In_1075,In_886);
or U394 (N_394,In_260,In_1062);
and U395 (N_395,In_746,In_228);
nand U396 (N_396,In_56,In_739);
or U397 (N_397,In_837,In_249);
xor U398 (N_398,In_534,In_198);
or U399 (N_399,In_915,In_1495);
nand U400 (N_400,In_1228,In_688);
nand U401 (N_401,In_938,In_396);
xnor U402 (N_402,In_293,In_1121);
nor U403 (N_403,In_1091,In_691);
nand U404 (N_404,In_814,In_1194);
xnor U405 (N_405,In_1146,In_1020);
nand U406 (N_406,In_1272,In_174);
nand U407 (N_407,In_766,In_427);
and U408 (N_408,In_380,In_385);
nand U409 (N_409,In_446,In_652);
and U410 (N_410,In_450,In_970);
nand U411 (N_411,In_780,In_952);
xnor U412 (N_412,In_147,In_514);
and U413 (N_413,In_1033,In_348);
xnor U414 (N_414,In_679,In_549);
and U415 (N_415,In_525,In_213);
and U416 (N_416,In_197,In_209);
or U417 (N_417,In_904,In_203);
nor U418 (N_418,In_1467,In_1056);
xnor U419 (N_419,In_634,In_394);
nand U420 (N_420,In_72,In_1221);
xnor U421 (N_421,In_37,In_250);
nor U422 (N_422,In_65,In_684);
nand U423 (N_423,In_239,In_1412);
xor U424 (N_424,In_403,In_857);
and U425 (N_425,In_1,In_1245);
or U426 (N_426,In_1046,In_568);
and U427 (N_427,In_1406,In_1049);
nand U428 (N_428,In_909,In_905);
or U429 (N_429,In_1060,In_144);
and U430 (N_430,In_1159,In_829);
nand U431 (N_431,In_1052,In_630);
nand U432 (N_432,In_478,In_390);
nor U433 (N_433,In_1417,In_1208);
nand U434 (N_434,In_280,In_1418);
or U435 (N_435,In_116,In_453);
nand U436 (N_436,In_710,In_1081);
or U437 (N_437,In_1446,In_599);
xnor U438 (N_438,In_1142,In_1252);
or U439 (N_439,In_236,In_617);
nor U440 (N_440,In_1456,In_1435);
or U441 (N_441,In_199,In_1316);
or U442 (N_442,In_785,In_844);
nor U443 (N_443,In_1344,In_1254);
and U444 (N_444,In_1152,In_456);
nand U445 (N_445,In_639,In_247);
or U446 (N_446,In_1451,In_412);
nor U447 (N_447,In_845,In_828);
and U448 (N_448,In_128,In_1447);
nand U449 (N_449,In_1030,In_1161);
or U450 (N_450,In_614,In_1261);
and U451 (N_451,In_499,In_1013);
xor U452 (N_452,In_1318,In_846);
and U453 (N_453,In_676,In_425);
xor U454 (N_454,In_187,In_1352);
nand U455 (N_455,In_982,In_442);
nand U456 (N_456,In_900,In_756);
or U457 (N_457,In_40,In_945);
nand U458 (N_458,In_1181,In_227);
and U459 (N_459,In_868,In_1358);
and U460 (N_460,In_913,In_916);
and U461 (N_461,In_1179,In_971);
nor U462 (N_462,In_721,In_219);
and U463 (N_463,In_942,In_836);
or U464 (N_464,In_926,In_1338);
or U465 (N_465,In_1263,In_303);
xnor U466 (N_466,In_1330,In_290);
or U467 (N_467,In_947,In_151);
or U468 (N_468,In_102,In_1459);
xor U469 (N_469,In_87,In_1306);
nor U470 (N_470,In_1348,In_764);
nor U471 (N_471,In_943,In_1410);
xnor U472 (N_472,In_700,In_182);
and U473 (N_473,In_1073,In_4);
nor U474 (N_474,In_217,In_95);
nand U475 (N_475,In_838,In_1010);
or U476 (N_476,In_974,In_190);
xor U477 (N_477,In_1116,In_687);
and U478 (N_478,In_833,In_1453);
and U479 (N_479,In_13,In_85);
nor U480 (N_480,In_1064,In_1442);
and U481 (N_481,In_479,In_757);
or U482 (N_482,In_268,In_53);
or U483 (N_483,In_454,In_1198);
or U484 (N_484,In_317,In_800);
nor U485 (N_485,In_66,In_1248);
nand U486 (N_486,In_129,In_18);
and U487 (N_487,In_181,In_1175);
nand U488 (N_488,In_1301,In_296);
and U489 (N_489,In_1172,In_778);
nor U490 (N_490,In_889,In_166);
and U491 (N_491,In_1496,In_463);
nand U492 (N_492,In_1065,In_1349);
xor U493 (N_493,In_63,In_248);
xor U494 (N_494,In_1101,In_44);
xor U495 (N_495,In_743,In_720);
or U496 (N_496,In_612,In_1072);
or U497 (N_497,In_153,In_173);
xor U498 (N_498,In_794,In_851);
or U499 (N_499,In_1266,In_1454);
xor U500 (N_500,In_582,In_299);
and U501 (N_501,In_271,In_576);
nor U502 (N_502,In_701,In_196);
xnor U503 (N_503,In_122,In_30);
xnor U504 (N_504,In_92,In_1093);
nor U505 (N_505,In_747,In_680);
and U506 (N_506,In_321,In_830);
xor U507 (N_507,In_1267,In_914);
or U508 (N_508,In_1021,In_1234);
xor U509 (N_509,In_580,In_1040);
xnor U510 (N_510,In_1328,In_362);
or U511 (N_511,In_591,In_136);
nor U512 (N_512,In_1297,In_96);
and U513 (N_513,In_596,In_407);
and U514 (N_514,In_336,In_1428);
nor U515 (N_515,In_765,In_1011);
xor U516 (N_516,In_678,In_806);
xor U517 (N_517,In_364,In_564);
and U518 (N_518,In_669,In_379);
xnor U519 (N_519,In_781,In_465);
nor U520 (N_520,In_367,In_1392);
xor U521 (N_521,In_951,In_787);
nor U522 (N_522,In_725,In_461);
or U523 (N_523,In_510,In_1389);
nor U524 (N_524,In_430,In_991);
xnor U525 (N_525,In_346,In_11);
and U526 (N_526,In_1005,In_245);
nand U527 (N_527,In_1325,In_158);
nand U528 (N_528,In_753,In_45);
nand U529 (N_529,In_1186,In_967);
nor U530 (N_530,In_39,In_1367);
nand U531 (N_531,In_545,In_216);
nand U532 (N_532,In_163,In_667);
or U533 (N_533,In_681,In_28);
or U534 (N_534,In_895,In_378);
and U535 (N_535,In_54,In_1308);
or U536 (N_536,In_389,In_1312);
nand U537 (N_537,In_1475,In_1457);
and U538 (N_538,In_1053,In_1026);
and U539 (N_539,In_232,In_1237);
nor U540 (N_540,In_1250,In_1054);
nand U541 (N_541,In_411,In_243);
and U542 (N_542,In_637,In_331);
nor U543 (N_543,In_300,In_455);
nand U544 (N_544,In_398,In_565);
and U545 (N_545,In_870,In_965);
xnor U546 (N_546,In_1138,In_579);
nor U547 (N_547,In_827,In_1177);
xor U548 (N_548,In_1336,In_987);
or U549 (N_549,In_21,In_1335);
or U550 (N_550,In_559,In_1373);
and U551 (N_551,In_81,In_1067);
xnor U552 (N_552,In_17,In_726);
nor U553 (N_553,In_391,In_744);
nor U554 (N_554,In_1034,In_1015);
or U555 (N_555,In_104,In_843);
and U556 (N_556,In_1167,In_405);
and U557 (N_557,In_923,In_1253);
nand U558 (N_558,In_192,In_1074);
and U559 (N_559,In_1099,In_961);
xor U560 (N_560,In_1419,In_1111);
xor U561 (N_561,In_334,In_1150);
nor U562 (N_562,In_333,In_41);
xor U563 (N_563,In_864,In_473);
or U564 (N_564,In_1157,In_714);
or U565 (N_565,In_933,In_918);
xor U566 (N_566,In_1284,In_1105);
and U567 (N_567,In_160,In_1341);
and U568 (N_568,In_137,In_557);
nand U569 (N_569,In_335,In_1050);
nand U570 (N_570,In_980,In_1265);
nor U571 (N_571,In_606,In_212);
xnor U572 (N_572,In_1039,In_1031);
nor U573 (N_573,In_516,In_922);
and U574 (N_574,In_42,In_592);
nand U575 (N_575,In_941,In_152);
nand U576 (N_576,In_1051,In_818);
nor U577 (N_577,In_481,In_295);
nor U578 (N_578,In_48,In_1486);
nor U579 (N_579,In_402,In_1473);
and U580 (N_580,In_1009,In_1190);
nand U581 (N_581,In_960,In_406);
xnor U582 (N_582,In_863,In_620);
nor U583 (N_583,In_986,In_1365);
nor U584 (N_584,In_177,In_1191);
nand U585 (N_585,In_341,In_1223);
nor U586 (N_586,In_1282,In_191);
and U587 (N_587,In_968,In_1006);
or U588 (N_588,In_1136,In_587);
nand U589 (N_589,In_902,In_1487);
or U590 (N_590,In_717,In_853);
and U591 (N_591,In_1176,In_1184);
or U592 (N_592,In_877,In_410);
nor U593 (N_593,In_984,In_368);
xor U594 (N_594,In_285,In_159);
and U595 (N_595,In_1478,In_1168);
xnor U596 (N_596,In_1498,In_447);
nor U597 (N_597,In_729,In_1371);
xor U598 (N_598,In_46,In_742);
or U599 (N_599,In_628,In_1476);
and U600 (N_600,In_1058,In_891);
nand U601 (N_601,In_616,In_1069);
nand U602 (N_602,In_588,In_804);
or U603 (N_603,In_636,In_515);
or U604 (N_604,In_755,In_632);
xnor U605 (N_605,In_771,In_27);
or U606 (N_606,In_660,In_1302);
or U607 (N_607,In_594,In_155);
or U608 (N_608,In_256,In_615);
or U609 (N_609,In_840,In_1434);
and U610 (N_610,In_1137,In_973);
nand U611 (N_611,In_839,In_677);
or U612 (N_612,In_930,In_1012);
xnor U613 (N_613,In_1474,In_1479);
xnor U614 (N_614,In_329,In_342);
or U615 (N_615,In_887,In_1106);
or U616 (N_616,In_610,In_324);
and U617 (N_617,In_924,In_1313);
or U618 (N_618,In_1036,In_393);
nand U619 (N_619,In_1057,In_1381);
nor U620 (N_620,In_1094,In_100);
and U621 (N_621,In_1118,In_433);
or U622 (N_622,In_470,In_603);
or U623 (N_623,In_375,In_997);
xor U624 (N_624,In_264,In_50);
xnor U625 (N_625,In_1331,In_1304);
nand U626 (N_626,In_117,In_1090);
nand U627 (N_627,In_278,In_856);
and U628 (N_628,In_776,In_1357);
xor U629 (N_629,In_215,In_520);
xnor U630 (N_630,In_858,In_154);
nor U631 (N_631,In_763,In_441);
xnor U632 (N_632,In_1370,In_483);
or U633 (N_633,In_88,In_172);
xnor U634 (N_634,In_583,In_1480);
nor U635 (N_635,In_34,In_120);
xnor U636 (N_636,In_908,In_313);
nand U637 (N_637,In_1397,In_1409);
xnor U638 (N_638,In_270,In_257);
or U639 (N_639,In_662,In_1319);
nor U640 (N_640,In_1189,In_118);
or U641 (N_641,In_439,In_1274);
and U642 (N_642,In_330,In_493);
or U643 (N_643,In_1290,In_149);
nor U644 (N_644,In_1361,In_1087);
xnor U645 (N_645,In_1375,In_693);
and U646 (N_646,In_426,In_189);
nor U647 (N_647,In_503,In_310);
or U648 (N_648,In_1154,In_1183);
nor U649 (N_649,In_852,In_976);
or U650 (N_650,In_1083,In_458);
nor U651 (N_651,In_530,In_883);
xnor U652 (N_652,In_1327,In_240);
xnor U653 (N_653,In_464,In_419);
xor U654 (N_654,In_896,In_106);
nor U655 (N_655,In_325,In_665);
nand U656 (N_656,In_1227,In_1215);
or U657 (N_657,In_1353,In_1170);
nor U658 (N_658,In_696,In_1214);
and U659 (N_659,In_1359,In_598);
or U660 (N_660,In_432,In_1461);
and U661 (N_661,In_275,In_1079);
xnor U662 (N_662,In_835,In_476);
nand U663 (N_663,In_47,In_138);
nor U664 (N_664,In_881,In_1038);
and U665 (N_665,In_1211,In_1432);
and U666 (N_666,In_935,In_64);
and U667 (N_667,In_1445,In_937);
xnor U668 (N_668,In_1209,In_241);
or U669 (N_669,In_188,In_911);
nand U670 (N_670,In_597,In_1471);
xnor U671 (N_671,In_627,In_948);
and U672 (N_672,In_1281,In_1242);
or U673 (N_673,In_950,In_141);
and U674 (N_674,In_567,In_894);
nor U675 (N_675,In_1379,In_556);
nor U676 (N_676,In_651,In_999);
or U677 (N_677,In_265,In_823);
xnor U678 (N_678,In_1388,In_445);
or U679 (N_679,In_156,In_484);
nor U680 (N_680,In_262,In_489);
nor U681 (N_681,In_1233,In_108);
xor U682 (N_682,In_1326,In_801);
nand U683 (N_683,In_1236,In_1257);
xnor U684 (N_684,In_1023,In_349);
nor U685 (N_685,In_1438,In_642);
nand U686 (N_686,In_496,In_558);
nand U687 (N_687,In_536,In_1366);
xor U688 (N_688,In_1469,In_697);
xnor U689 (N_689,In_1165,In_487);
nor U690 (N_690,In_32,In_370);
nor U691 (N_691,In_184,In_640);
nor U692 (N_692,In_1277,In_1232);
xnor U693 (N_693,In_365,In_653);
nor U694 (N_694,In_920,In_1202);
nand U695 (N_695,In_477,In_1477);
nor U696 (N_696,In_713,In_1014);
and U697 (N_697,In_71,In_452);
nor U698 (N_698,In_723,In_1044);
nand U699 (N_699,In_1420,In_1201);
nand U700 (N_700,In_969,In_816);
xor U701 (N_701,In_1382,In_959);
nor U702 (N_702,In_1264,In_371);
nor U703 (N_703,In_626,In_901);
xnor U704 (N_704,In_387,In_850);
and U705 (N_705,In_1255,In_770);
xnor U706 (N_706,In_1205,In_993);
nand U707 (N_707,In_35,In_1249);
and U708 (N_708,In_416,In_813);
or U709 (N_709,In_659,In_413);
nor U710 (N_710,In_543,In_903);
nor U711 (N_711,In_1246,In_848);
or U712 (N_712,In_436,In_802);
or U713 (N_713,In_1145,In_538);
or U714 (N_714,In_882,In_1309);
or U715 (N_715,In_1022,In_77);
nor U716 (N_716,In_707,In_204);
xnor U717 (N_717,In_841,In_578);
or U718 (N_718,In_1213,In_114);
nand U719 (N_719,In_1048,In_928);
nand U720 (N_720,In_1466,In_237);
nor U721 (N_721,In_277,In_8);
and U722 (N_722,In_885,In_337);
xor U723 (N_723,In_621,In_383);
and U724 (N_724,In_1380,In_1024);
nor U725 (N_725,In_1377,In_339);
nor U726 (N_726,In_253,In_1007);
nand U727 (N_727,In_672,In_5);
nor U728 (N_728,In_570,In_1364);
nor U729 (N_729,In_884,In_618);
or U730 (N_730,In_1088,In_1374);
xor U731 (N_731,In_815,In_619);
or U732 (N_732,In_502,In_89);
or U733 (N_733,In_527,In_674);
nor U734 (N_734,In_176,In_508);
nand U735 (N_735,In_9,In_420);
nor U736 (N_736,In_560,In_2);
or U737 (N_737,In_1310,In_777);
nand U738 (N_738,In_734,In_899);
or U739 (N_739,In_1329,In_1472);
and U740 (N_740,In_170,In_1315);
xor U741 (N_741,In_847,In_1002);
or U742 (N_742,In_1171,In_573);
nor U743 (N_743,In_690,In_19);
or U744 (N_744,In_983,In_1416);
nor U745 (N_745,In_709,In_319);
nand U746 (N_746,In_1080,In_246);
and U747 (N_747,In_62,In_491);
xnor U748 (N_748,In_731,In_26);
or U749 (N_749,In_832,In_1440);
xnor U750 (N_750,In_66,In_1275);
nand U751 (N_751,In_54,In_499);
or U752 (N_752,In_1486,In_320);
xnor U753 (N_753,In_122,In_270);
and U754 (N_754,In_203,In_1081);
or U755 (N_755,In_408,In_650);
nor U756 (N_756,In_1218,In_263);
nand U757 (N_757,In_1356,In_1183);
and U758 (N_758,In_811,In_671);
nand U759 (N_759,In_879,In_1259);
nand U760 (N_760,In_808,In_930);
xnor U761 (N_761,In_368,In_1049);
or U762 (N_762,In_1269,In_184);
nor U763 (N_763,In_1135,In_929);
nor U764 (N_764,In_45,In_437);
nor U765 (N_765,In_357,In_854);
or U766 (N_766,In_1131,In_1428);
nor U767 (N_767,In_1217,In_1209);
nand U768 (N_768,In_782,In_431);
and U769 (N_769,In_1427,In_1131);
nor U770 (N_770,In_678,In_481);
nor U771 (N_771,In_1045,In_1104);
xor U772 (N_772,In_555,In_1398);
or U773 (N_773,In_209,In_1107);
nor U774 (N_774,In_841,In_151);
nand U775 (N_775,In_1344,In_588);
nor U776 (N_776,In_1240,In_274);
xnor U777 (N_777,In_1356,In_960);
and U778 (N_778,In_436,In_394);
or U779 (N_779,In_901,In_539);
xnor U780 (N_780,In_573,In_1323);
and U781 (N_781,In_748,In_738);
xnor U782 (N_782,In_1203,In_837);
xnor U783 (N_783,In_73,In_811);
xor U784 (N_784,In_1249,In_146);
nor U785 (N_785,In_1277,In_1217);
and U786 (N_786,In_926,In_1214);
nand U787 (N_787,In_1200,In_1319);
nand U788 (N_788,In_998,In_929);
xor U789 (N_789,In_381,In_75);
nor U790 (N_790,In_932,In_357);
and U791 (N_791,In_1402,In_825);
xnor U792 (N_792,In_1106,In_28);
nand U793 (N_793,In_756,In_30);
or U794 (N_794,In_1171,In_306);
nand U795 (N_795,In_1396,In_1419);
nand U796 (N_796,In_940,In_116);
or U797 (N_797,In_521,In_1335);
nand U798 (N_798,In_450,In_1440);
nand U799 (N_799,In_331,In_1157);
nor U800 (N_800,In_807,In_1394);
nor U801 (N_801,In_1139,In_254);
nor U802 (N_802,In_373,In_193);
or U803 (N_803,In_14,In_536);
nor U804 (N_804,In_1198,In_264);
nor U805 (N_805,In_1238,In_834);
nand U806 (N_806,In_238,In_1410);
or U807 (N_807,In_833,In_513);
nor U808 (N_808,In_6,In_1432);
or U809 (N_809,In_1189,In_749);
xor U810 (N_810,In_714,In_1403);
nand U811 (N_811,In_89,In_436);
nand U812 (N_812,In_420,In_1408);
xnor U813 (N_813,In_812,In_44);
and U814 (N_814,In_1321,In_1489);
or U815 (N_815,In_679,In_405);
or U816 (N_816,In_292,In_902);
nor U817 (N_817,In_39,In_1089);
or U818 (N_818,In_243,In_652);
and U819 (N_819,In_1144,In_1347);
nor U820 (N_820,In_295,In_237);
and U821 (N_821,In_1373,In_777);
nor U822 (N_822,In_485,In_704);
and U823 (N_823,In_1175,In_185);
or U824 (N_824,In_1057,In_889);
nand U825 (N_825,In_1290,In_524);
nor U826 (N_826,In_685,In_1023);
nand U827 (N_827,In_1173,In_1489);
nand U828 (N_828,In_1325,In_705);
and U829 (N_829,In_645,In_138);
or U830 (N_830,In_201,In_195);
xnor U831 (N_831,In_1406,In_548);
xor U832 (N_832,In_254,In_1296);
xnor U833 (N_833,In_660,In_586);
or U834 (N_834,In_1353,In_52);
xnor U835 (N_835,In_1263,In_99);
or U836 (N_836,In_1034,In_1196);
nand U837 (N_837,In_1223,In_675);
nand U838 (N_838,In_431,In_1034);
or U839 (N_839,In_962,In_776);
and U840 (N_840,In_1494,In_1369);
and U841 (N_841,In_579,In_244);
nor U842 (N_842,In_1027,In_839);
xor U843 (N_843,In_1024,In_622);
and U844 (N_844,In_1491,In_36);
or U845 (N_845,In_1434,In_592);
nor U846 (N_846,In_1380,In_431);
xnor U847 (N_847,In_534,In_564);
or U848 (N_848,In_17,In_839);
xor U849 (N_849,In_800,In_1351);
nor U850 (N_850,In_441,In_1225);
or U851 (N_851,In_662,In_629);
nand U852 (N_852,In_811,In_495);
xor U853 (N_853,In_138,In_495);
or U854 (N_854,In_15,In_826);
nand U855 (N_855,In_664,In_1424);
or U856 (N_856,In_381,In_705);
nor U857 (N_857,In_959,In_869);
or U858 (N_858,In_1010,In_176);
xnor U859 (N_859,In_279,In_335);
xor U860 (N_860,In_543,In_1162);
or U861 (N_861,In_1202,In_656);
nand U862 (N_862,In_585,In_955);
nand U863 (N_863,In_916,In_165);
nand U864 (N_864,In_1404,In_163);
xnor U865 (N_865,In_82,In_833);
and U866 (N_866,In_122,In_12);
xnor U867 (N_867,In_1235,In_810);
nor U868 (N_868,In_654,In_727);
nand U869 (N_869,In_368,In_23);
and U870 (N_870,In_1122,In_298);
nor U871 (N_871,In_1303,In_847);
and U872 (N_872,In_48,In_1359);
and U873 (N_873,In_1413,In_1162);
xnor U874 (N_874,In_438,In_1015);
nor U875 (N_875,In_1440,In_427);
and U876 (N_876,In_72,In_452);
nor U877 (N_877,In_1397,In_1342);
nor U878 (N_878,In_923,In_954);
nor U879 (N_879,In_593,In_257);
or U880 (N_880,In_135,In_486);
nand U881 (N_881,In_945,In_1452);
xnor U882 (N_882,In_1012,In_1495);
xnor U883 (N_883,In_505,In_997);
nor U884 (N_884,In_1226,In_1242);
xor U885 (N_885,In_536,In_855);
and U886 (N_886,In_1190,In_331);
nor U887 (N_887,In_972,In_1381);
nand U888 (N_888,In_0,In_1418);
nor U889 (N_889,In_995,In_922);
or U890 (N_890,In_1382,In_403);
nand U891 (N_891,In_877,In_322);
or U892 (N_892,In_1145,In_578);
nand U893 (N_893,In_16,In_539);
and U894 (N_894,In_34,In_627);
and U895 (N_895,In_622,In_538);
nand U896 (N_896,In_1079,In_816);
nand U897 (N_897,In_1389,In_105);
nand U898 (N_898,In_1353,In_79);
or U899 (N_899,In_229,In_68);
and U900 (N_900,In_423,In_731);
nor U901 (N_901,In_675,In_175);
nor U902 (N_902,In_832,In_394);
and U903 (N_903,In_788,In_1177);
or U904 (N_904,In_566,In_137);
xor U905 (N_905,In_746,In_720);
nand U906 (N_906,In_892,In_954);
or U907 (N_907,In_642,In_1076);
or U908 (N_908,In_1408,In_423);
nor U909 (N_909,In_1394,In_1486);
nor U910 (N_910,In_1261,In_1346);
nor U911 (N_911,In_428,In_1110);
nor U912 (N_912,In_1201,In_501);
xnor U913 (N_913,In_938,In_1456);
nor U914 (N_914,In_1073,In_1473);
and U915 (N_915,In_1210,In_972);
xor U916 (N_916,In_351,In_507);
or U917 (N_917,In_685,In_28);
or U918 (N_918,In_764,In_1430);
and U919 (N_919,In_1310,In_911);
xor U920 (N_920,In_90,In_1459);
nor U921 (N_921,In_357,In_974);
nor U922 (N_922,In_559,In_85);
or U923 (N_923,In_1066,In_773);
or U924 (N_924,In_1437,In_1342);
xor U925 (N_925,In_1445,In_1381);
nor U926 (N_926,In_53,In_175);
or U927 (N_927,In_121,In_165);
nand U928 (N_928,In_770,In_1036);
and U929 (N_929,In_1072,In_318);
or U930 (N_930,In_1006,In_1174);
xor U931 (N_931,In_1276,In_236);
or U932 (N_932,In_822,In_791);
or U933 (N_933,In_1072,In_655);
nand U934 (N_934,In_18,In_715);
or U935 (N_935,In_1474,In_945);
nand U936 (N_936,In_1205,In_750);
and U937 (N_937,In_1257,In_1357);
nand U938 (N_938,In_91,In_1415);
xor U939 (N_939,In_1299,In_404);
xnor U940 (N_940,In_15,In_1171);
nand U941 (N_941,In_65,In_649);
and U942 (N_942,In_1398,In_1015);
nor U943 (N_943,In_1295,In_1055);
nor U944 (N_944,In_1116,In_1184);
nor U945 (N_945,In_1370,In_999);
nand U946 (N_946,In_528,In_562);
or U947 (N_947,In_1228,In_62);
nor U948 (N_948,In_443,In_1140);
nand U949 (N_949,In_1135,In_164);
nor U950 (N_950,In_384,In_196);
or U951 (N_951,In_1065,In_1495);
nand U952 (N_952,In_950,In_786);
nand U953 (N_953,In_1097,In_48);
nand U954 (N_954,In_1199,In_1334);
nor U955 (N_955,In_141,In_1046);
xnor U956 (N_956,In_1461,In_1228);
nor U957 (N_957,In_827,In_395);
nor U958 (N_958,In_1215,In_1156);
or U959 (N_959,In_1242,In_55);
nand U960 (N_960,In_1325,In_1144);
xnor U961 (N_961,In_1488,In_907);
or U962 (N_962,In_837,In_652);
nand U963 (N_963,In_344,In_133);
or U964 (N_964,In_1443,In_1194);
nand U965 (N_965,In_1370,In_326);
and U966 (N_966,In_600,In_1372);
and U967 (N_967,In_982,In_147);
and U968 (N_968,In_1387,In_232);
or U969 (N_969,In_1055,In_1375);
and U970 (N_970,In_1087,In_517);
nor U971 (N_971,In_698,In_1470);
nand U972 (N_972,In_573,In_958);
or U973 (N_973,In_427,In_343);
or U974 (N_974,In_1183,In_858);
or U975 (N_975,In_86,In_165);
and U976 (N_976,In_717,In_191);
or U977 (N_977,In_304,In_815);
or U978 (N_978,In_1491,In_1112);
or U979 (N_979,In_262,In_1188);
xnor U980 (N_980,In_834,In_242);
nand U981 (N_981,In_186,In_131);
or U982 (N_982,In_942,In_1368);
and U983 (N_983,In_1070,In_672);
nor U984 (N_984,In_835,In_143);
xor U985 (N_985,In_195,In_235);
and U986 (N_986,In_623,In_1351);
and U987 (N_987,In_576,In_412);
xor U988 (N_988,In_61,In_1360);
nand U989 (N_989,In_814,In_1277);
nor U990 (N_990,In_681,In_916);
or U991 (N_991,In_826,In_277);
nand U992 (N_992,In_589,In_898);
xor U993 (N_993,In_1008,In_169);
or U994 (N_994,In_918,In_516);
and U995 (N_995,In_1327,In_832);
nor U996 (N_996,In_484,In_300);
and U997 (N_997,In_9,In_259);
nand U998 (N_998,In_1096,In_803);
and U999 (N_999,In_912,In_1094);
or U1000 (N_1000,N_843,N_778);
nor U1001 (N_1001,N_922,N_55);
nand U1002 (N_1002,N_511,N_22);
nor U1003 (N_1003,N_373,N_720);
and U1004 (N_1004,N_305,N_752);
nand U1005 (N_1005,N_649,N_19);
xnor U1006 (N_1006,N_17,N_127);
or U1007 (N_1007,N_495,N_998);
nor U1008 (N_1008,N_247,N_601);
and U1009 (N_1009,N_958,N_287);
and U1010 (N_1010,N_555,N_957);
xnor U1011 (N_1011,N_900,N_662);
and U1012 (N_1012,N_997,N_806);
nand U1013 (N_1013,N_297,N_242);
and U1014 (N_1014,N_238,N_407);
nor U1015 (N_1015,N_603,N_79);
xor U1016 (N_1016,N_303,N_481);
xnor U1017 (N_1017,N_702,N_751);
nor U1018 (N_1018,N_626,N_479);
nand U1019 (N_1019,N_231,N_943);
xor U1020 (N_1020,N_356,N_188);
and U1021 (N_1021,N_24,N_875);
and U1022 (N_1022,N_872,N_400);
nor U1023 (N_1023,N_657,N_936);
and U1024 (N_1024,N_325,N_978);
and U1025 (N_1025,N_250,N_146);
nor U1026 (N_1026,N_651,N_731);
nand U1027 (N_1027,N_929,N_696);
xor U1028 (N_1028,N_976,N_49);
or U1029 (N_1029,N_189,N_505);
nand U1030 (N_1030,N_629,N_15);
or U1031 (N_1031,N_834,N_638);
and U1032 (N_1032,N_541,N_719);
and U1033 (N_1033,N_167,N_40);
xnor U1034 (N_1034,N_46,N_658);
nor U1035 (N_1035,N_882,N_97);
xor U1036 (N_1036,N_164,N_502);
nand U1037 (N_1037,N_472,N_320);
nand U1038 (N_1038,N_95,N_573);
and U1039 (N_1039,N_367,N_483);
and U1040 (N_1040,N_873,N_123);
nand U1041 (N_1041,N_909,N_119);
nor U1042 (N_1042,N_235,N_216);
nand U1043 (N_1043,N_947,N_299);
nand U1044 (N_1044,N_920,N_624);
nand U1045 (N_1045,N_608,N_493);
nor U1046 (N_1046,N_270,N_286);
and U1047 (N_1047,N_448,N_469);
and U1048 (N_1048,N_265,N_730);
or U1049 (N_1049,N_0,N_849);
and U1050 (N_1050,N_380,N_881);
xor U1051 (N_1051,N_723,N_918);
and U1052 (N_1052,N_864,N_755);
or U1053 (N_1053,N_600,N_888);
nand U1054 (N_1054,N_961,N_521);
xnor U1055 (N_1055,N_399,N_422);
xor U1056 (N_1056,N_342,N_398);
or U1057 (N_1057,N_53,N_903);
and U1058 (N_1058,N_508,N_532);
or U1059 (N_1059,N_642,N_948);
xnor U1060 (N_1060,N_425,N_243);
or U1061 (N_1061,N_239,N_648);
xnor U1062 (N_1062,N_294,N_574);
or U1063 (N_1063,N_126,N_896);
nand U1064 (N_1064,N_383,N_768);
or U1065 (N_1065,N_366,N_312);
xor U1066 (N_1066,N_518,N_546);
nand U1067 (N_1067,N_656,N_331);
nand U1068 (N_1068,N_543,N_132);
xnor U1069 (N_1069,N_722,N_817);
nand U1070 (N_1070,N_330,N_458);
nand U1071 (N_1071,N_438,N_424);
xor U1072 (N_1072,N_455,N_606);
nand U1073 (N_1073,N_646,N_758);
nand U1074 (N_1074,N_637,N_522);
nand U1075 (N_1075,N_906,N_309);
nand U1076 (N_1076,N_28,N_290);
and U1077 (N_1077,N_482,N_799);
and U1078 (N_1078,N_104,N_426);
nand U1079 (N_1079,N_59,N_214);
xor U1080 (N_1080,N_322,N_847);
and U1081 (N_1081,N_45,N_468);
and U1082 (N_1082,N_332,N_939);
nor U1083 (N_1083,N_489,N_402);
nand U1084 (N_1084,N_803,N_134);
xnor U1085 (N_1085,N_108,N_484);
or U1086 (N_1086,N_578,N_435);
nor U1087 (N_1087,N_317,N_116);
nor U1088 (N_1088,N_158,N_473);
and U1089 (N_1089,N_210,N_636);
nand U1090 (N_1090,N_615,N_259);
or U1091 (N_1091,N_418,N_512);
nor U1092 (N_1092,N_839,N_343);
xnor U1093 (N_1093,N_419,N_241);
and U1094 (N_1094,N_694,N_691);
or U1095 (N_1095,N_395,N_644);
nor U1096 (N_1096,N_571,N_995);
or U1097 (N_1097,N_740,N_826);
nand U1098 (N_1098,N_491,N_496);
nor U1099 (N_1099,N_340,N_570);
or U1100 (N_1100,N_897,N_2);
nor U1101 (N_1101,N_678,N_80);
xor U1102 (N_1102,N_612,N_335);
nor U1103 (N_1103,N_82,N_683);
and U1104 (N_1104,N_57,N_863);
or U1105 (N_1105,N_219,N_413);
nand U1106 (N_1106,N_128,N_403);
nand U1107 (N_1107,N_627,N_833);
or U1108 (N_1108,N_766,N_793);
nor U1109 (N_1109,N_810,N_439);
and U1110 (N_1110,N_237,N_314);
and U1111 (N_1111,N_739,N_862);
or U1112 (N_1112,N_783,N_699);
xnor U1113 (N_1113,N_263,N_351);
nor U1114 (N_1114,N_60,N_355);
and U1115 (N_1115,N_4,N_973);
and U1116 (N_1116,N_951,N_474);
nor U1117 (N_1117,N_20,N_647);
and U1118 (N_1118,N_218,N_911);
or U1119 (N_1119,N_92,N_728);
nor U1120 (N_1120,N_744,N_892);
and U1121 (N_1121,N_180,N_273);
xnor U1122 (N_1122,N_851,N_971);
or U1123 (N_1123,N_490,N_292);
nand U1124 (N_1124,N_724,N_359);
nand U1125 (N_1125,N_791,N_234);
xnor U1126 (N_1126,N_344,N_765);
or U1127 (N_1127,N_676,N_618);
nand U1128 (N_1128,N_148,N_328);
nand U1129 (N_1129,N_954,N_827);
xnor U1130 (N_1130,N_446,N_232);
nand U1131 (N_1131,N_829,N_860);
and U1132 (N_1132,N_634,N_200);
nand U1133 (N_1133,N_753,N_240);
nor U1134 (N_1134,N_423,N_650);
nand U1135 (N_1135,N_197,N_185);
nand U1136 (N_1136,N_462,N_575);
xor U1137 (N_1137,N_371,N_831);
and U1138 (N_1138,N_786,N_252);
nor U1139 (N_1139,N_224,N_712);
nor U1140 (N_1140,N_497,N_725);
and U1141 (N_1141,N_244,N_280);
nand U1142 (N_1142,N_893,N_401);
and U1143 (N_1143,N_196,N_856);
nor U1144 (N_1144,N_152,N_602);
and U1145 (N_1145,N_414,N_926);
nor U1146 (N_1146,N_186,N_825);
nand U1147 (N_1147,N_865,N_75);
nand U1148 (N_1148,N_348,N_397);
and U1149 (N_1149,N_572,N_952);
xnor U1150 (N_1150,N_486,N_143);
nor U1151 (N_1151,N_433,N_52);
nor U1152 (N_1152,N_178,N_985);
xnor U1153 (N_1153,N_176,N_51);
or U1154 (N_1154,N_391,N_930);
nor U1155 (N_1155,N_376,N_655);
nand U1156 (N_1156,N_925,N_223);
or U1157 (N_1157,N_96,N_315);
xnor U1158 (N_1158,N_544,N_44);
or U1159 (N_1159,N_111,N_733);
or U1160 (N_1160,N_538,N_558);
xor U1161 (N_1161,N_855,N_254);
xnor U1162 (N_1162,N_110,N_345);
or U1163 (N_1163,N_107,N_278);
nor U1164 (N_1164,N_449,N_289);
nor U1165 (N_1165,N_537,N_557);
xor U1166 (N_1166,N_592,N_747);
nand U1167 (N_1167,N_692,N_807);
nand U1168 (N_1168,N_828,N_979);
nor U1169 (N_1169,N_498,N_378);
nor U1170 (N_1170,N_434,N_142);
and U1171 (N_1171,N_883,N_736);
and U1172 (N_1172,N_494,N_835);
and U1173 (N_1173,N_70,N_809);
nand U1174 (N_1174,N_771,N_23);
xor U1175 (N_1175,N_184,N_800);
nand U1176 (N_1176,N_745,N_100);
xor U1177 (N_1177,N_307,N_727);
nand U1178 (N_1178,N_777,N_302);
or U1179 (N_1179,N_837,N_967);
nand U1180 (N_1180,N_689,N_974);
xor U1181 (N_1181,N_861,N_179);
or U1182 (N_1182,N_715,N_296);
or U1183 (N_1183,N_229,N_977);
xnor U1184 (N_1184,N_871,N_531);
nand U1185 (N_1185,N_716,N_598);
or U1186 (N_1186,N_63,N_452);
nor U1187 (N_1187,N_569,N_151);
nand U1188 (N_1188,N_159,N_282);
nand U1189 (N_1189,N_90,N_412);
nand U1190 (N_1190,N_787,N_106);
nor U1191 (N_1191,N_198,N_118);
nand U1192 (N_1192,N_905,N_515);
and U1193 (N_1193,N_748,N_10);
nand U1194 (N_1194,N_684,N_870);
and U1195 (N_1195,N_761,N_352);
and U1196 (N_1196,N_545,N_620);
nor U1197 (N_1197,N_705,N_587);
or U1198 (N_1198,N_346,N_659);
or U1199 (N_1199,N_155,N_276);
xor U1200 (N_1200,N_21,N_671);
xnor U1201 (N_1201,N_962,N_854);
and U1202 (N_1202,N_451,N_157);
or U1203 (N_1203,N_945,N_131);
nor U1204 (N_1204,N_842,N_277);
or U1205 (N_1205,N_972,N_135);
nand U1206 (N_1206,N_37,N_996);
nor U1207 (N_1207,N_792,N_361);
xor U1208 (N_1208,N_919,N_554);
nand U1209 (N_1209,N_408,N_710);
nand U1210 (N_1210,N_393,N_898);
xor U1211 (N_1211,N_421,N_295);
nor U1212 (N_1212,N_640,N_960);
xnor U1213 (N_1213,N_595,N_822);
xor U1214 (N_1214,N_830,N_653);
and U1215 (N_1215,N_480,N_641);
nor U1216 (N_1216,N_666,N_221);
and U1217 (N_1217,N_983,N_841);
nor U1218 (N_1218,N_306,N_713);
xnor U1219 (N_1219,N_275,N_12);
or U1220 (N_1220,N_818,N_389);
nor U1221 (N_1221,N_341,N_639);
and U1222 (N_1222,N_9,N_409);
nor U1223 (N_1223,N_30,N_160);
nand U1224 (N_1224,N_514,N_526);
and U1225 (N_1225,N_222,N_124);
xnor U1226 (N_1226,N_144,N_946);
nand U1227 (N_1227,N_623,N_886);
or U1228 (N_1228,N_567,N_547);
nor U1229 (N_1229,N_625,N_779);
or U1230 (N_1230,N_99,N_884);
or U1231 (N_1231,N_520,N_927);
or U1232 (N_1232,N_770,N_704);
nand U1233 (N_1233,N_207,N_316);
nand U1234 (N_1234,N_838,N_813);
xor U1235 (N_1235,N_551,N_323);
nand U1236 (N_1236,N_660,N_867);
nand U1237 (N_1237,N_227,N_665);
and U1238 (N_1238,N_271,N_597);
nand U1239 (N_1239,N_932,N_68);
xor U1240 (N_1240,N_467,N_668);
and U1241 (N_1241,N_251,N_992);
xnor U1242 (N_1242,N_533,N_141);
and U1243 (N_1243,N_27,N_153);
nand U1244 (N_1244,N_16,N_56);
nand U1245 (N_1245,N_476,N_729);
nor U1246 (N_1246,N_129,N_616);
nor U1247 (N_1247,N_794,N_388);
or U1248 (N_1248,N_894,N_941);
nand U1249 (N_1249,N_324,N_174);
or U1250 (N_1250,N_39,N_910);
or U1251 (N_1251,N_584,N_591);
and U1252 (N_1252,N_246,N_695);
and U1253 (N_1253,N_445,N_274);
nor U1254 (N_1254,N_610,N_86);
xnor U1255 (N_1255,N_844,N_81);
or U1256 (N_1256,N_669,N_528);
or U1257 (N_1257,N_621,N_802);
xnor U1258 (N_1258,N_553,N_857);
nor U1259 (N_1259,N_74,N_327);
and U1260 (N_1260,N_887,N_969);
and U1261 (N_1261,N_673,N_364);
xor U1262 (N_1262,N_970,N_233);
nor U1263 (N_1263,N_256,N_607);
xor U1264 (N_1264,N_891,N_944);
nand U1265 (N_1265,N_195,N_172);
nor U1266 (N_1266,N_921,N_199);
nor U1267 (N_1267,N_581,N_840);
and U1268 (N_1268,N_226,N_949);
nand U1269 (N_1269,N_411,N_585);
nor U1270 (N_1270,N_536,N_980);
xnor U1271 (N_1271,N_850,N_769);
or U1272 (N_1272,N_688,N_812);
nor U1273 (N_1273,N_13,N_816);
nor U1274 (N_1274,N_773,N_808);
nand U1275 (N_1275,N_801,N_248);
and U1276 (N_1276,N_261,N_71);
nor U1277 (N_1277,N_923,N_443);
xnor U1278 (N_1278,N_133,N_154);
and U1279 (N_1279,N_614,N_741);
nand U1280 (N_1280,N_820,N_166);
nand U1281 (N_1281,N_47,N_776);
or U1282 (N_1282,N_953,N_717);
or U1283 (N_1283,N_427,N_162);
xor U1284 (N_1284,N_566,N_631);
nor U1285 (N_1285,N_457,N_645);
or U1286 (N_1286,N_58,N_788);
nor U1287 (N_1287,N_742,N_268);
xnor U1288 (N_1288,N_115,N_304);
nand U1289 (N_1289,N_635,N_83);
and U1290 (N_1290,N_228,N_54);
nand U1291 (N_1291,N_853,N_982);
nor U1292 (N_1292,N_815,N_145);
and U1293 (N_1293,N_895,N_698);
and U1294 (N_1294,N_913,N_150);
nor U1295 (N_1295,N_103,N_501);
nand U1296 (N_1296,N_846,N_91);
nand U1297 (N_1297,N_619,N_375);
nor U1298 (N_1298,N_137,N_685);
xnor U1299 (N_1299,N_372,N_249);
xor U1300 (N_1300,N_301,N_697);
or U1301 (N_1301,N_1,N_789);
and U1302 (N_1302,N_576,N_459);
and U1303 (N_1303,N_681,N_6);
or U1304 (N_1304,N_77,N_734);
and U1305 (N_1305,N_169,N_140);
or U1306 (N_1306,N_101,N_805);
xor U1307 (N_1307,N_738,N_743);
and U1308 (N_1308,N_213,N_622);
or U1309 (N_1309,N_475,N_994);
and U1310 (N_1310,N_524,N_611);
and U1311 (N_1311,N_950,N_726);
xnor U1312 (N_1312,N_350,N_506);
nor U1313 (N_1313,N_318,N_487);
xor U1314 (N_1314,N_202,N_109);
nor U1315 (N_1315,N_663,N_488);
and U1316 (N_1316,N_105,N_852);
xnor U1317 (N_1317,N_313,N_879);
nand U1318 (N_1318,N_362,N_548);
and U1319 (N_1319,N_711,N_321);
xor U1320 (N_1320,N_173,N_390);
xor U1321 (N_1321,N_530,N_599);
or U1322 (N_1322,N_191,N_319);
or U1323 (N_1323,N_347,N_379);
nor U1324 (N_1324,N_763,N_561);
xor U1325 (N_1325,N_590,N_593);
or U1326 (N_1326,N_464,N_682);
nor U1327 (N_1327,N_18,N_670);
nor U1328 (N_1328,N_262,N_7);
xor U1329 (N_1329,N_14,N_78);
xor U1330 (N_1330,N_876,N_337);
nor U1331 (N_1331,N_163,N_194);
nor U1332 (N_1332,N_440,N_507);
nand U1333 (N_1333,N_284,N_975);
nor U1334 (N_1334,N_529,N_499);
nor U1335 (N_1335,N_613,N_394);
xnor U1336 (N_1336,N_504,N_796);
xnor U1337 (N_1337,N_293,N_374);
nor U1338 (N_1338,N_429,N_121);
and U1339 (N_1339,N_667,N_415);
nor U1340 (N_1340,N_260,N_845);
nor U1341 (N_1341,N_935,N_230);
xnor U1342 (N_1342,N_764,N_336);
nor U1343 (N_1343,N_353,N_357);
xnor U1344 (N_1344,N_182,N_756);
xnor U1345 (N_1345,N_754,N_999);
and U1346 (N_1346,N_48,N_981);
or U1347 (N_1347,N_125,N_774);
or U1348 (N_1348,N_29,N_69);
nand U1349 (N_1349,N_33,N_370);
nand U1350 (N_1350,N_382,N_255);
nor U1351 (N_1351,N_643,N_525);
nor U1352 (N_1352,N_664,N_986);
or U1353 (N_1353,N_938,N_594);
or U1354 (N_1354,N_334,N_785);
and U1355 (N_1355,N_706,N_329);
nor U1356 (N_1356,N_279,N_757);
nor U1357 (N_1357,N_914,N_338);
nor U1358 (N_1358,N_183,N_510);
nor U1359 (N_1359,N_385,N_604);
nor U1360 (N_1360,N_212,N_444);
xnor U1361 (N_1361,N_565,N_61);
and U1362 (N_1362,N_675,N_396);
nor U1363 (N_1363,N_354,N_72);
or U1364 (N_1364,N_384,N_288);
nor U1365 (N_1365,N_477,N_453);
nor U1366 (N_1366,N_31,N_269);
nand U1367 (N_1367,N_762,N_775);
or U1368 (N_1368,N_955,N_441);
nor U1369 (N_1369,N_114,N_782);
nand U1370 (N_1370,N_877,N_549);
or U1371 (N_1371,N_93,N_386);
nor U1372 (N_1372,N_406,N_804);
and U1373 (N_1373,N_492,N_596);
or U1374 (N_1374,N_693,N_456);
nand U1375 (N_1375,N_880,N_750);
nor U1376 (N_1376,N_956,N_392);
xor U1377 (N_1377,N_560,N_707);
or U1378 (N_1378,N_283,N_217);
and U1379 (N_1379,N_326,N_257);
and U1380 (N_1380,N_89,N_517);
nand U1381 (N_1381,N_737,N_236);
and U1382 (N_1382,N_211,N_85);
and U1383 (N_1383,N_908,N_98);
nand U1384 (N_1384,N_417,N_966);
xor U1385 (N_1385,N_513,N_5);
or U1386 (N_1386,N_703,N_933);
nor U1387 (N_1387,N_192,N_963);
xor U1388 (N_1388,N_404,N_201);
and U1389 (N_1389,N_405,N_586);
nand U1390 (N_1390,N_11,N_25);
nand U1391 (N_1391,N_66,N_869);
or U1392 (N_1392,N_187,N_899);
xnor U1393 (N_1393,N_358,N_215);
and U1394 (N_1394,N_432,N_130);
xnor U1395 (N_1395,N_266,N_718);
or U1396 (N_1396,N_442,N_917);
xor U1397 (N_1397,N_912,N_363);
nor U1398 (N_1398,N_661,N_87);
or U1399 (N_1399,N_206,N_577);
xnor U1400 (N_1400,N_420,N_959);
nor U1401 (N_1401,N_915,N_814);
and U1402 (N_1402,N_220,N_527);
xnor U1403 (N_1403,N_258,N_466);
xnor U1404 (N_1404,N_50,N_746);
xnor U1405 (N_1405,N_62,N_858);
nor U1406 (N_1406,N_36,N_461);
and U1407 (N_1407,N_94,N_32);
nor U1408 (N_1408,N_253,N_868);
or U1409 (N_1409,N_550,N_781);
nand U1410 (N_1410,N_387,N_580);
and U1411 (N_1411,N_878,N_583);
and U1412 (N_1412,N_700,N_721);
and U1413 (N_1413,N_790,N_8);
nand U1414 (N_1414,N_931,N_735);
and U1415 (N_1415,N_463,N_848);
or U1416 (N_1416,N_795,N_500);
nor U1417 (N_1417,N_937,N_410);
and U1418 (N_1418,N_122,N_890);
xnor U1419 (N_1419,N_245,N_64);
or U1420 (N_1420,N_759,N_523);
nor U1421 (N_1421,N_349,N_934);
or U1422 (N_1422,N_563,N_360);
or U1423 (N_1423,N_171,N_907);
nor U1424 (N_1424,N_630,N_964);
xnor U1425 (N_1425,N_714,N_381);
xor U1426 (N_1426,N_628,N_709);
nand U1427 (N_1427,N_3,N_987);
or U1428 (N_1428,N_165,N_552);
and U1429 (N_1429,N_365,N_672);
xor U1430 (N_1430,N_35,N_798);
or U1431 (N_1431,N_609,N_377);
nand U1432 (N_1432,N_701,N_225);
nor U1433 (N_1433,N_450,N_485);
nor U1434 (N_1434,N_928,N_333);
and U1435 (N_1435,N_113,N_968);
nor U1436 (N_1436,N_120,N_836);
xnor U1437 (N_1437,N_267,N_885);
nand U1438 (N_1438,N_519,N_821);
nand U1439 (N_1439,N_991,N_285);
nand U1440 (N_1440,N_677,N_589);
nand U1441 (N_1441,N_904,N_298);
and U1442 (N_1442,N_147,N_708);
or U1443 (N_1443,N_824,N_139);
or U1444 (N_1444,N_264,N_168);
nor U1445 (N_1445,N_43,N_732);
and U1446 (N_1446,N_416,N_208);
or U1447 (N_1447,N_564,N_509);
xor U1448 (N_1448,N_540,N_562);
or U1449 (N_1449,N_680,N_65);
nand U1450 (N_1450,N_535,N_633);
nand U1451 (N_1451,N_652,N_161);
nand U1452 (N_1452,N_272,N_26);
nand U1453 (N_1453,N_582,N_42);
nor U1454 (N_1454,N_874,N_436);
nand U1455 (N_1455,N_654,N_989);
and U1456 (N_1456,N_889,N_539);
nand U1457 (N_1457,N_942,N_674);
nor U1458 (N_1458,N_556,N_209);
or U1459 (N_1459,N_428,N_503);
nand U1460 (N_1460,N_310,N_916);
or U1461 (N_1461,N_993,N_568);
or U1462 (N_1462,N_308,N_454);
nand U1463 (N_1463,N_823,N_859);
nor U1464 (N_1464,N_460,N_749);
nand U1465 (N_1465,N_117,N_149);
or U1466 (N_1466,N_772,N_311);
xor U1467 (N_1467,N_478,N_339);
and U1468 (N_1468,N_203,N_465);
nor U1469 (N_1469,N_534,N_368);
or U1470 (N_1470,N_369,N_204);
nand U1471 (N_1471,N_588,N_797);
xnor U1472 (N_1472,N_431,N_76);
nand U1473 (N_1473,N_516,N_832);
and U1474 (N_1474,N_679,N_866);
and U1475 (N_1475,N_901,N_579);
xor U1476 (N_1476,N_88,N_156);
nand U1477 (N_1477,N_175,N_924);
and U1478 (N_1478,N_984,N_965);
xor U1479 (N_1479,N_84,N_811);
and U1480 (N_1480,N_38,N_138);
or U1481 (N_1481,N_112,N_617);
or U1482 (N_1482,N_605,N_205);
nor U1483 (N_1483,N_990,N_686);
nor U1484 (N_1484,N_760,N_193);
xor U1485 (N_1485,N_470,N_34);
and U1486 (N_1486,N_136,N_559);
nand U1487 (N_1487,N_41,N_632);
nor U1488 (N_1488,N_940,N_300);
nand U1489 (N_1489,N_181,N_447);
or U1490 (N_1490,N_767,N_430);
and U1491 (N_1491,N_471,N_819);
nand U1492 (N_1492,N_780,N_687);
nand U1493 (N_1493,N_690,N_291);
and U1494 (N_1494,N_281,N_902);
xnor U1495 (N_1495,N_784,N_177);
nor U1496 (N_1496,N_170,N_437);
and U1497 (N_1497,N_67,N_190);
and U1498 (N_1498,N_988,N_102);
xnor U1499 (N_1499,N_542,N_73);
or U1500 (N_1500,N_531,N_509);
and U1501 (N_1501,N_841,N_52);
or U1502 (N_1502,N_679,N_220);
nand U1503 (N_1503,N_881,N_829);
xor U1504 (N_1504,N_469,N_623);
or U1505 (N_1505,N_207,N_603);
xor U1506 (N_1506,N_662,N_573);
or U1507 (N_1507,N_315,N_68);
nand U1508 (N_1508,N_2,N_586);
nor U1509 (N_1509,N_762,N_788);
nand U1510 (N_1510,N_702,N_173);
nand U1511 (N_1511,N_216,N_946);
nor U1512 (N_1512,N_164,N_699);
nor U1513 (N_1513,N_655,N_47);
xnor U1514 (N_1514,N_299,N_515);
xnor U1515 (N_1515,N_216,N_874);
xnor U1516 (N_1516,N_139,N_246);
and U1517 (N_1517,N_181,N_766);
xnor U1518 (N_1518,N_415,N_691);
nand U1519 (N_1519,N_2,N_440);
or U1520 (N_1520,N_455,N_712);
nor U1521 (N_1521,N_613,N_158);
nand U1522 (N_1522,N_71,N_949);
nand U1523 (N_1523,N_813,N_65);
xnor U1524 (N_1524,N_701,N_99);
or U1525 (N_1525,N_948,N_557);
xnor U1526 (N_1526,N_115,N_17);
nand U1527 (N_1527,N_2,N_900);
or U1528 (N_1528,N_741,N_309);
and U1529 (N_1529,N_456,N_50);
and U1530 (N_1530,N_161,N_346);
and U1531 (N_1531,N_256,N_231);
or U1532 (N_1532,N_817,N_45);
nor U1533 (N_1533,N_760,N_976);
and U1534 (N_1534,N_268,N_828);
xor U1535 (N_1535,N_451,N_10);
nand U1536 (N_1536,N_228,N_489);
or U1537 (N_1537,N_593,N_317);
or U1538 (N_1538,N_612,N_285);
nand U1539 (N_1539,N_661,N_672);
and U1540 (N_1540,N_41,N_348);
xnor U1541 (N_1541,N_639,N_399);
nor U1542 (N_1542,N_809,N_459);
nor U1543 (N_1543,N_377,N_983);
and U1544 (N_1544,N_217,N_414);
and U1545 (N_1545,N_222,N_325);
xor U1546 (N_1546,N_788,N_754);
or U1547 (N_1547,N_708,N_649);
or U1548 (N_1548,N_165,N_336);
nand U1549 (N_1549,N_199,N_638);
nor U1550 (N_1550,N_462,N_385);
xnor U1551 (N_1551,N_360,N_171);
nand U1552 (N_1552,N_694,N_882);
xnor U1553 (N_1553,N_999,N_606);
xor U1554 (N_1554,N_555,N_219);
or U1555 (N_1555,N_200,N_982);
and U1556 (N_1556,N_845,N_504);
and U1557 (N_1557,N_99,N_642);
nand U1558 (N_1558,N_801,N_914);
or U1559 (N_1559,N_148,N_851);
or U1560 (N_1560,N_724,N_83);
xnor U1561 (N_1561,N_910,N_226);
xnor U1562 (N_1562,N_552,N_949);
xnor U1563 (N_1563,N_766,N_532);
xnor U1564 (N_1564,N_482,N_147);
nand U1565 (N_1565,N_141,N_326);
nand U1566 (N_1566,N_693,N_722);
or U1567 (N_1567,N_221,N_983);
and U1568 (N_1568,N_432,N_59);
xnor U1569 (N_1569,N_460,N_455);
xnor U1570 (N_1570,N_915,N_688);
and U1571 (N_1571,N_727,N_500);
xor U1572 (N_1572,N_719,N_966);
xnor U1573 (N_1573,N_164,N_628);
or U1574 (N_1574,N_85,N_874);
and U1575 (N_1575,N_479,N_378);
xnor U1576 (N_1576,N_851,N_900);
xnor U1577 (N_1577,N_547,N_920);
nor U1578 (N_1578,N_90,N_137);
nand U1579 (N_1579,N_678,N_133);
nand U1580 (N_1580,N_852,N_32);
nor U1581 (N_1581,N_734,N_331);
nor U1582 (N_1582,N_714,N_311);
and U1583 (N_1583,N_266,N_526);
nand U1584 (N_1584,N_911,N_746);
nor U1585 (N_1585,N_888,N_97);
xor U1586 (N_1586,N_248,N_676);
and U1587 (N_1587,N_46,N_259);
or U1588 (N_1588,N_529,N_267);
xor U1589 (N_1589,N_315,N_44);
or U1590 (N_1590,N_583,N_470);
xnor U1591 (N_1591,N_423,N_195);
xor U1592 (N_1592,N_766,N_716);
or U1593 (N_1593,N_194,N_92);
and U1594 (N_1594,N_808,N_539);
nor U1595 (N_1595,N_761,N_178);
or U1596 (N_1596,N_780,N_810);
xor U1597 (N_1597,N_884,N_815);
xor U1598 (N_1598,N_888,N_720);
and U1599 (N_1599,N_295,N_731);
nor U1600 (N_1600,N_107,N_512);
or U1601 (N_1601,N_909,N_992);
nand U1602 (N_1602,N_27,N_151);
nor U1603 (N_1603,N_180,N_403);
and U1604 (N_1604,N_385,N_503);
nor U1605 (N_1605,N_402,N_248);
nand U1606 (N_1606,N_227,N_64);
xnor U1607 (N_1607,N_399,N_92);
nor U1608 (N_1608,N_454,N_964);
nand U1609 (N_1609,N_192,N_42);
nor U1610 (N_1610,N_852,N_139);
or U1611 (N_1611,N_350,N_114);
or U1612 (N_1612,N_958,N_864);
nor U1613 (N_1613,N_891,N_706);
nor U1614 (N_1614,N_926,N_626);
nor U1615 (N_1615,N_739,N_660);
or U1616 (N_1616,N_66,N_454);
xor U1617 (N_1617,N_605,N_641);
nand U1618 (N_1618,N_749,N_513);
and U1619 (N_1619,N_691,N_339);
and U1620 (N_1620,N_694,N_19);
and U1621 (N_1621,N_327,N_248);
nand U1622 (N_1622,N_453,N_883);
xor U1623 (N_1623,N_598,N_419);
nand U1624 (N_1624,N_322,N_357);
or U1625 (N_1625,N_755,N_748);
nor U1626 (N_1626,N_134,N_875);
nor U1627 (N_1627,N_624,N_220);
or U1628 (N_1628,N_9,N_921);
or U1629 (N_1629,N_435,N_14);
and U1630 (N_1630,N_249,N_919);
and U1631 (N_1631,N_444,N_843);
or U1632 (N_1632,N_248,N_76);
or U1633 (N_1633,N_292,N_946);
or U1634 (N_1634,N_909,N_849);
and U1635 (N_1635,N_887,N_74);
nand U1636 (N_1636,N_424,N_463);
nor U1637 (N_1637,N_287,N_365);
or U1638 (N_1638,N_811,N_857);
nand U1639 (N_1639,N_809,N_950);
nand U1640 (N_1640,N_248,N_424);
xor U1641 (N_1641,N_180,N_150);
or U1642 (N_1642,N_522,N_246);
nor U1643 (N_1643,N_370,N_626);
nand U1644 (N_1644,N_557,N_813);
and U1645 (N_1645,N_204,N_873);
nor U1646 (N_1646,N_95,N_758);
and U1647 (N_1647,N_887,N_918);
nor U1648 (N_1648,N_966,N_666);
and U1649 (N_1649,N_211,N_693);
nand U1650 (N_1650,N_296,N_624);
xor U1651 (N_1651,N_268,N_704);
xnor U1652 (N_1652,N_681,N_256);
or U1653 (N_1653,N_321,N_387);
or U1654 (N_1654,N_16,N_311);
nand U1655 (N_1655,N_58,N_330);
nor U1656 (N_1656,N_580,N_897);
xor U1657 (N_1657,N_522,N_63);
nor U1658 (N_1658,N_227,N_872);
nor U1659 (N_1659,N_519,N_804);
and U1660 (N_1660,N_230,N_293);
xor U1661 (N_1661,N_637,N_85);
xnor U1662 (N_1662,N_726,N_359);
nor U1663 (N_1663,N_545,N_826);
nand U1664 (N_1664,N_101,N_570);
nand U1665 (N_1665,N_22,N_509);
nand U1666 (N_1666,N_683,N_655);
or U1667 (N_1667,N_91,N_179);
or U1668 (N_1668,N_429,N_825);
and U1669 (N_1669,N_458,N_217);
xor U1670 (N_1670,N_957,N_486);
nand U1671 (N_1671,N_286,N_963);
xor U1672 (N_1672,N_268,N_591);
and U1673 (N_1673,N_734,N_459);
xnor U1674 (N_1674,N_478,N_634);
xor U1675 (N_1675,N_196,N_575);
or U1676 (N_1676,N_45,N_920);
or U1677 (N_1677,N_397,N_641);
xnor U1678 (N_1678,N_828,N_377);
and U1679 (N_1679,N_661,N_401);
nor U1680 (N_1680,N_600,N_598);
or U1681 (N_1681,N_560,N_817);
xor U1682 (N_1682,N_749,N_579);
nand U1683 (N_1683,N_757,N_258);
nor U1684 (N_1684,N_269,N_112);
or U1685 (N_1685,N_130,N_284);
xnor U1686 (N_1686,N_20,N_961);
or U1687 (N_1687,N_942,N_235);
or U1688 (N_1688,N_976,N_25);
and U1689 (N_1689,N_820,N_188);
and U1690 (N_1690,N_358,N_652);
nand U1691 (N_1691,N_657,N_231);
and U1692 (N_1692,N_465,N_806);
xnor U1693 (N_1693,N_53,N_996);
or U1694 (N_1694,N_572,N_139);
or U1695 (N_1695,N_186,N_274);
nand U1696 (N_1696,N_706,N_963);
and U1697 (N_1697,N_486,N_702);
and U1698 (N_1698,N_604,N_43);
nand U1699 (N_1699,N_849,N_853);
nand U1700 (N_1700,N_299,N_982);
nand U1701 (N_1701,N_237,N_257);
and U1702 (N_1702,N_727,N_722);
and U1703 (N_1703,N_560,N_946);
nor U1704 (N_1704,N_995,N_373);
xor U1705 (N_1705,N_942,N_99);
xnor U1706 (N_1706,N_227,N_905);
and U1707 (N_1707,N_334,N_469);
xnor U1708 (N_1708,N_949,N_118);
xor U1709 (N_1709,N_209,N_18);
xnor U1710 (N_1710,N_408,N_14);
and U1711 (N_1711,N_249,N_332);
or U1712 (N_1712,N_626,N_294);
and U1713 (N_1713,N_393,N_331);
and U1714 (N_1714,N_35,N_549);
nand U1715 (N_1715,N_58,N_857);
nand U1716 (N_1716,N_812,N_729);
nor U1717 (N_1717,N_51,N_61);
xor U1718 (N_1718,N_150,N_326);
xor U1719 (N_1719,N_33,N_774);
xnor U1720 (N_1720,N_263,N_177);
and U1721 (N_1721,N_807,N_51);
and U1722 (N_1722,N_570,N_275);
or U1723 (N_1723,N_200,N_66);
and U1724 (N_1724,N_337,N_450);
nor U1725 (N_1725,N_990,N_659);
nand U1726 (N_1726,N_193,N_373);
and U1727 (N_1727,N_598,N_579);
or U1728 (N_1728,N_25,N_318);
and U1729 (N_1729,N_730,N_258);
or U1730 (N_1730,N_944,N_82);
xnor U1731 (N_1731,N_354,N_189);
nand U1732 (N_1732,N_88,N_396);
or U1733 (N_1733,N_869,N_163);
and U1734 (N_1734,N_738,N_497);
nor U1735 (N_1735,N_586,N_608);
nor U1736 (N_1736,N_334,N_315);
nor U1737 (N_1737,N_869,N_985);
nor U1738 (N_1738,N_46,N_652);
xor U1739 (N_1739,N_212,N_534);
nand U1740 (N_1740,N_506,N_136);
nor U1741 (N_1741,N_999,N_960);
or U1742 (N_1742,N_699,N_445);
nand U1743 (N_1743,N_470,N_500);
or U1744 (N_1744,N_895,N_879);
nor U1745 (N_1745,N_0,N_114);
and U1746 (N_1746,N_809,N_250);
nand U1747 (N_1747,N_769,N_49);
xor U1748 (N_1748,N_502,N_275);
xnor U1749 (N_1749,N_693,N_479);
xnor U1750 (N_1750,N_768,N_699);
xor U1751 (N_1751,N_561,N_494);
and U1752 (N_1752,N_733,N_951);
xor U1753 (N_1753,N_685,N_159);
and U1754 (N_1754,N_383,N_891);
nand U1755 (N_1755,N_624,N_161);
or U1756 (N_1756,N_959,N_226);
and U1757 (N_1757,N_326,N_972);
and U1758 (N_1758,N_203,N_9);
nor U1759 (N_1759,N_695,N_292);
nor U1760 (N_1760,N_810,N_637);
nor U1761 (N_1761,N_125,N_643);
nor U1762 (N_1762,N_824,N_207);
or U1763 (N_1763,N_814,N_278);
or U1764 (N_1764,N_389,N_375);
nor U1765 (N_1765,N_281,N_383);
xnor U1766 (N_1766,N_254,N_51);
or U1767 (N_1767,N_139,N_611);
nand U1768 (N_1768,N_454,N_243);
and U1769 (N_1769,N_333,N_289);
and U1770 (N_1770,N_166,N_154);
nand U1771 (N_1771,N_511,N_362);
or U1772 (N_1772,N_200,N_383);
or U1773 (N_1773,N_32,N_248);
or U1774 (N_1774,N_797,N_494);
nor U1775 (N_1775,N_185,N_395);
nor U1776 (N_1776,N_993,N_555);
nand U1777 (N_1777,N_243,N_702);
or U1778 (N_1778,N_954,N_684);
nor U1779 (N_1779,N_720,N_664);
and U1780 (N_1780,N_486,N_714);
nand U1781 (N_1781,N_275,N_699);
and U1782 (N_1782,N_88,N_691);
nand U1783 (N_1783,N_67,N_477);
nor U1784 (N_1784,N_492,N_349);
and U1785 (N_1785,N_77,N_915);
and U1786 (N_1786,N_39,N_528);
nor U1787 (N_1787,N_208,N_707);
or U1788 (N_1788,N_452,N_457);
and U1789 (N_1789,N_924,N_787);
nor U1790 (N_1790,N_874,N_218);
and U1791 (N_1791,N_951,N_563);
nor U1792 (N_1792,N_974,N_792);
nor U1793 (N_1793,N_771,N_211);
xor U1794 (N_1794,N_927,N_148);
nor U1795 (N_1795,N_976,N_800);
xnor U1796 (N_1796,N_617,N_526);
xnor U1797 (N_1797,N_628,N_734);
nand U1798 (N_1798,N_959,N_316);
and U1799 (N_1799,N_909,N_393);
nor U1800 (N_1800,N_709,N_428);
nand U1801 (N_1801,N_794,N_903);
or U1802 (N_1802,N_641,N_504);
nand U1803 (N_1803,N_585,N_591);
xor U1804 (N_1804,N_889,N_390);
and U1805 (N_1805,N_67,N_249);
xor U1806 (N_1806,N_507,N_473);
nand U1807 (N_1807,N_842,N_647);
and U1808 (N_1808,N_799,N_159);
or U1809 (N_1809,N_918,N_799);
nor U1810 (N_1810,N_735,N_399);
nor U1811 (N_1811,N_25,N_814);
or U1812 (N_1812,N_404,N_416);
xnor U1813 (N_1813,N_366,N_35);
nor U1814 (N_1814,N_677,N_272);
nand U1815 (N_1815,N_738,N_552);
and U1816 (N_1816,N_116,N_596);
xor U1817 (N_1817,N_349,N_329);
xor U1818 (N_1818,N_949,N_244);
nand U1819 (N_1819,N_726,N_138);
or U1820 (N_1820,N_428,N_257);
and U1821 (N_1821,N_449,N_915);
xnor U1822 (N_1822,N_326,N_189);
and U1823 (N_1823,N_468,N_39);
nor U1824 (N_1824,N_870,N_974);
and U1825 (N_1825,N_131,N_990);
and U1826 (N_1826,N_614,N_219);
nand U1827 (N_1827,N_513,N_517);
xnor U1828 (N_1828,N_112,N_11);
and U1829 (N_1829,N_703,N_940);
nor U1830 (N_1830,N_897,N_348);
xnor U1831 (N_1831,N_702,N_784);
xor U1832 (N_1832,N_946,N_56);
or U1833 (N_1833,N_128,N_244);
and U1834 (N_1834,N_48,N_18);
xnor U1835 (N_1835,N_987,N_748);
nand U1836 (N_1836,N_36,N_379);
xor U1837 (N_1837,N_793,N_226);
and U1838 (N_1838,N_270,N_289);
nand U1839 (N_1839,N_366,N_99);
and U1840 (N_1840,N_172,N_327);
and U1841 (N_1841,N_664,N_7);
or U1842 (N_1842,N_79,N_902);
or U1843 (N_1843,N_877,N_529);
nand U1844 (N_1844,N_383,N_298);
nor U1845 (N_1845,N_944,N_781);
nand U1846 (N_1846,N_681,N_199);
and U1847 (N_1847,N_194,N_506);
nor U1848 (N_1848,N_638,N_324);
nor U1849 (N_1849,N_441,N_945);
xor U1850 (N_1850,N_857,N_931);
xnor U1851 (N_1851,N_554,N_738);
xnor U1852 (N_1852,N_870,N_96);
xor U1853 (N_1853,N_194,N_207);
nand U1854 (N_1854,N_626,N_446);
nand U1855 (N_1855,N_607,N_819);
or U1856 (N_1856,N_444,N_708);
xnor U1857 (N_1857,N_484,N_46);
nand U1858 (N_1858,N_197,N_626);
nand U1859 (N_1859,N_535,N_441);
nor U1860 (N_1860,N_775,N_17);
and U1861 (N_1861,N_753,N_907);
or U1862 (N_1862,N_35,N_446);
nand U1863 (N_1863,N_5,N_100);
nand U1864 (N_1864,N_409,N_317);
xor U1865 (N_1865,N_621,N_660);
and U1866 (N_1866,N_680,N_985);
or U1867 (N_1867,N_642,N_390);
and U1868 (N_1868,N_462,N_370);
and U1869 (N_1869,N_446,N_348);
and U1870 (N_1870,N_463,N_204);
nor U1871 (N_1871,N_148,N_326);
nor U1872 (N_1872,N_41,N_60);
and U1873 (N_1873,N_455,N_599);
or U1874 (N_1874,N_828,N_697);
nand U1875 (N_1875,N_544,N_782);
nand U1876 (N_1876,N_339,N_29);
nand U1877 (N_1877,N_517,N_693);
xor U1878 (N_1878,N_859,N_578);
nand U1879 (N_1879,N_151,N_921);
nor U1880 (N_1880,N_793,N_455);
nand U1881 (N_1881,N_137,N_969);
nor U1882 (N_1882,N_29,N_438);
nor U1883 (N_1883,N_566,N_974);
and U1884 (N_1884,N_84,N_341);
or U1885 (N_1885,N_323,N_468);
nor U1886 (N_1886,N_981,N_794);
nand U1887 (N_1887,N_246,N_861);
nand U1888 (N_1888,N_831,N_505);
or U1889 (N_1889,N_107,N_303);
or U1890 (N_1890,N_810,N_686);
and U1891 (N_1891,N_758,N_622);
nand U1892 (N_1892,N_183,N_755);
nand U1893 (N_1893,N_875,N_379);
xor U1894 (N_1894,N_898,N_912);
or U1895 (N_1895,N_318,N_697);
nand U1896 (N_1896,N_791,N_254);
or U1897 (N_1897,N_143,N_541);
nor U1898 (N_1898,N_832,N_20);
and U1899 (N_1899,N_832,N_620);
and U1900 (N_1900,N_493,N_477);
nand U1901 (N_1901,N_895,N_2);
nand U1902 (N_1902,N_465,N_967);
and U1903 (N_1903,N_567,N_958);
or U1904 (N_1904,N_94,N_619);
and U1905 (N_1905,N_774,N_607);
nand U1906 (N_1906,N_236,N_146);
or U1907 (N_1907,N_804,N_682);
xnor U1908 (N_1908,N_780,N_90);
nor U1909 (N_1909,N_840,N_756);
and U1910 (N_1910,N_576,N_238);
and U1911 (N_1911,N_585,N_266);
nor U1912 (N_1912,N_243,N_200);
nor U1913 (N_1913,N_28,N_649);
nand U1914 (N_1914,N_739,N_424);
nand U1915 (N_1915,N_644,N_173);
or U1916 (N_1916,N_86,N_962);
nor U1917 (N_1917,N_307,N_428);
or U1918 (N_1918,N_3,N_683);
and U1919 (N_1919,N_223,N_84);
nor U1920 (N_1920,N_149,N_519);
or U1921 (N_1921,N_534,N_949);
and U1922 (N_1922,N_259,N_788);
or U1923 (N_1923,N_18,N_88);
nor U1924 (N_1924,N_229,N_822);
and U1925 (N_1925,N_459,N_830);
xor U1926 (N_1926,N_298,N_414);
xor U1927 (N_1927,N_229,N_839);
nor U1928 (N_1928,N_159,N_795);
xor U1929 (N_1929,N_777,N_664);
nor U1930 (N_1930,N_471,N_562);
nor U1931 (N_1931,N_144,N_235);
or U1932 (N_1932,N_979,N_483);
xor U1933 (N_1933,N_50,N_408);
or U1934 (N_1934,N_691,N_329);
nor U1935 (N_1935,N_110,N_824);
nand U1936 (N_1936,N_898,N_46);
or U1937 (N_1937,N_569,N_859);
xor U1938 (N_1938,N_64,N_147);
nand U1939 (N_1939,N_641,N_15);
nor U1940 (N_1940,N_841,N_248);
or U1941 (N_1941,N_327,N_932);
and U1942 (N_1942,N_765,N_274);
nor U1943 (N_1943,N_832,N_416);
nor U1944 (N_1944,N_896,N_55);
or U1945 (N_1945,N_30,N_434);
nand U1946 (N_1946,N_415,N_558);
nand U1947 (N_1947,N_366,N_235);
nor U1948 (N_1948,N_820,N_130);
and U1949 (N_1949,N_476,N_596);
or U1950 (N_1950,N_734,N_228);
or U1951 (N_1951,N_753,N_293);
nand U1952 (N_1952,N_713,N_213);
xnor U1953 (N_1953,N_238,N_43);
nand U1954 (N_1954,N_803,N_644);
nor U1955 (N_1955,N_726,N_408);
or U1956 (N_1956,N_975,N_367);
xnor U1957 (N_1957,N_909,N_37);
xor U1958 (N_1958,N_777,N_563);
xor U1959 (N_1959,N_994,N_209);
and U1960 (N_1960,N_494,N_654);
and U1961 (N_1961,N_483,N_808);
or U1962 (N_1962,N_787,N_508);
or U1963 (N_1963,N_279,N_935);
or U1964 (N_1964,N_88,N_31);
and U1965 (N_1965,N_619,N_557);
xnor U1966 (N_1966,N_435,N_171);
or U1967 (N_1967,N_578,N_877);
nor U1968 (N_1968,N_87,N_890);
xor U1969 (N_1969,N_12,N_564);
and U1970 (N_1970,N_359,N_141);
and U1971 (N_1971,N_351,N_73);
or U1972 (N_1972,N_757,N_49);
xor U1973 (N_1973,N_5,N_567);
or U1974 (N_1974,N_838,N_550);
and U1975 (N_1975,N_1,N_163);
xor U1976 (N_1976,N_109,N_967);
or U1977 (N_1977,N_352,N_370);
xnor U1978 (N_1978,N_532,N_185);
and U1979 (N_1979,N_828,N_482);
nand U1980 (N_1980,N_167,N_675);
and U1981 (N_1981,N_541,N_83);
nand U1982 (N_1982,N_830,N_942);
xor U1983 (N_1983,N_629,N_797);
xnor U1984 (N_1984,N_294,N_14);
xnor U1985 (N_1985,N_234,N_313);
and U1986 (N_1986,N_851,N_137);
and U1987 (N_1987,N_408,N_914);
and U1988 (N_1988,N_42,N_720);
and U1989 (N_1989,N_301,N_445);
or U1990 (N_1990,N_674,N_61);
nor U1991 (N_1991,N_677,N_471);
and U1992 (N_1992,N_113,N_372);
xnor U1993 (N_1993,N_161,N_296);
nor U1994 (N_1994,N_879,N_34);
and U1995 (N_1995,N_988,N_171);
xor U1996 (N_1996,N_800,N_541);
or U1997 (N_1997,N_124,N_567);
xnor U1998 (N_1998,N_143,N_488);
and U1999 (N_1999,N_999,N_676);
xnor U2000 (N_2000,N_1900,N_1876);
nand U2001 (N_2001,N_1787,N_1622);
nor U2002 (N_2002,N_1326,N_1884);
xnor U2003 (N_2003,N_1068,N_1005);
or U2004 (N_2004,N_1138,N_1383);
or U2005 (N_2005,N_1828,N_1352);
and U2006 (N_2006,N_1476,N_1936);
and U2007 (N_2007,N_1516,N_1151);
and U2008 (N_2008,N_1901,N_1971);
xnor U2009 (N_2009,N_1805,N_1701);
nor U2010 (N_2010,N_1466,N_1974);
nand U2011 (N_2011,N_1188,N_1109);
xor U2012 (N_2012,N_1888,N_1010);
and U2013 (N_2013,N_1248,N_1461);
nor U2014 (N_2014,N_1205,N_1446);
nor U2015 (N_2015,N_1897,N_1186);
nor U2016 (N_2016,N_1289,N_1447);
nand U2017 (N_2017,N_1645,N_1176);
xnor U2018 (N_2018,N_1565,N_1750);
or U2019 (N_2019,N_1296,N_1267);
or U2020 (N_2020,N_1742,N_1274);
nand U2021 (N_2021,N_1564,N_1295);
xnor U2022 (N_2022,N_1611,N_1252);
nand U2023 (N_2023,N_1146,N_1591);
and U2024 (N_2024,N_1480,N_1862);
nand U2025 (N_2025,N_1525,N_1669);
nand U2026 (N_2026,N_1962,N_1991);
or U2027 (N_2027,N_1297,N_1871);
xnor U2028 (N_2028,N_1505,N_1899);
xnor U2029 (N_2029,N_1756,N_1945);
xnor U2030 (N_2030,N_1639,N_1330);
and U2031 (N_2031,N_1287,N_1154);
and U2032 (N_2032,N_1391,N_1533);
and U2033 (N_2033,N_1382,N_1618);
nor U2034 (N_2034,N_1174,N_1209);
nand U2035 (N_2035,N_1780,N_1975);
nand U2036 (N_2036,N_1934,N_1989);
xnor U2037 (N_2037,N_1674,N_1958);
xnor U2038 (N_2038,N_1996,N_1143);
xor U2039 (N_2039,N_1272,N_1061);
or U2040 (N_2040,N_1924,N_1182);
or U2041 (N_2041,N_1173,N_1395);
nor U2042 (N_2042,N_1834,N_1025);
nor U2043 (N_2043,N_1967,N_1230);
or U2044 (N_2044,N_1624,N_1632);
xnor U2045 (N_2045,N_1221,N_1549);
xor U2046 (N_2046,N_1728,N_1022);
and U2047 (N_2047,N_1367,N_1265);
and U2048 (N_2048,N_1609,N_1983);
and U2049 (N_2049,N_1465,N_1096);
and U2050 (N_2050,N_1441,N_1054);
and U2051 (N_2051,N_1570,N_1518);
xnor U2052 (N_2052,N_1148,N_1698);
and U2053 (N_2053,N_1191,N_1699);
xor U2054 (N_2054,N_1359,N_1830);
and U2055 (N_2055,N_1571,N_1732);
and U2056 (N_2056,N_1088,N_1941);
nor U2057 (N_2057,N_1052,N_1215);
nand U2058 (N_2058,N_1016,N_1459);
and U2059 (N_2059,N_1140,N_1377);
nand U2060 (N_2060,N_1986,N_1372);
xnor U2061 (N_2061,N_1966,N_1492);
xnor U2062 (N_2062,N_1489,N_1360);
and U2063 (N_2063,N_1916,N_1069);
or U2064 (N_2064,N_1860,N_1740);
nor U2065 (N_2065,N_1385,N_1692);
xor U2066 (N_2066,N_1712,N_1262);
and U2067 (N_2067,N_1921,N_1895);
or U2068 (N_2068,N_1579,N_1055);
xor U2069 (N_2069,N_1613,N_1169);
nand U2070 (N_2070,N_1021,N_1908);
and U2071 (N_2071,N_1536,N_1988);
nor U2072 (N_2072,N_1535,N_1636);
nor U2073 (N_2073,N_1883,N_1702);
and U2074 (N_2074,N_1841,N_1387);
nand U2075 (N_2075,N_1523,N_1723);
or U2076 (N_2076,N_1027,N_1625);
xnor U2077 (N_2077,N_1757,N_1922);
or U2078 (N_2078,N_1208,N_1693);
and U2079 (N_2079,N_1759,N_1013);
nor U2080 (N_2080,N_1919,N_1784);
nor U2081 (N_2081,N_1233,N_1575);
nand U2082 (N_2082,N_1322,N_1709);
nor U2083 (N_2083,N_1543,N_1070);
nand U2084 (N_2084,N_1158,N_1846);
xnor U2085 (N_2085,N_1848,N_1339);
nand U2086 (N_2086,N_1494,N_1445);
xor U2087 (N_2087,N_1199,N_1724);
or U2088 (N_2088,N_1126,N_1519);
or U2089 (N_2089,N_1105,N_1462);
xnor U2090 (N_2090,N_1124,N_1413);
and U2091 (N_2091,N_1464,N_1521);
nor U2092 (N_2092,N_1635,N_1559);
nor U2093 (N_2093,N_1059,N_1039);
and U2094 (N_2094,N_1909,N_1280);
nand U2095 (N_2095,N_1878,N_1134);
nor U2096 (N_2096,N_1077,N_1179);
nor U2097 (N_2097,N_1074,N_1081);
nor U2098 (N_2098,N_1682,N_1875);
nor U2099 (N_2099,N_1153,N_1665);
nor U2100 (N_2100,N_1165,N_1951);
xor U2101 (N_2101,N_1578,N_1408);
and U2102 (N_2102,N_1977,N_1623);
or U2103 (N_2103,N_1576,N_1247);
nand U2104 (N_2104,N_1269,N_1911);
nand U2105 (N_2105,N_1325,N_1063);
nand U2106 (N_2106,N_1691,N_1243);
and U2107 (N_2107,N_1361,N_1453);
xor U2108 (N_2108,N_1356,N_1393);
or U2109 (N_2109,N_1402,N_1075);
nor U2110 (N_2110,N_1303,N_1946);
nor U2111 (N_2111,N_1586,N_1286);
nor U2112 (N_2112,N_1440,N_1117);
and U2113 (N_2113,N_1341,N_1019);
nand U2114 (N_2114,N_1515,N_1261);
and U2115 (N_2115,N_1204,N_1398);
or U2116 (N_2116,N_1870,N_1972);
nand U2117 (N_2117,N_1201,N_1171);
nand U2118 (N_2118,N_1420,N_1947);
or U2119 (N_2119,N_1646,N_1679);
and U2120 (N_2120,N_1668,N_1128);
nor U2121 (N_2121,N_1690,N_1125);
xnor U2122 (N_2122,N_1006,N_1782);
nor U2123 (N_2123,N_1345,N_1984);
nor U2124 (N_2124,N_1202,N_1599);
and U2125 (N_2125,N_1566,N_1244);
nor U2126 (N_2126,N_1416,N_1089);
and U2127 (N_2127,N_1431,N_1907);
or U2128 (N_2128,N_1813,N_1706);
nand U2129 (N_2129,N_1127,N_1593);
nor U2130 (N_2130,N_1455,N_1002);
nor U2131 (N_2131,N_1263,N_1275);
and U2132 (N_2132,N_1654,N_1042);
xor U2133 (N_2133,N_1568,N_1863);
and U2134 (N_2134,N_1386,N_1111);
xor U2135 (N_2135,N_1615,N_1601);
xnor U2136 (N_2136,N_1850,N_1219);
nor U2137 (N_2137,N_1246,N_1826);
xnor U2138 (N_2138,N_1452,N_1251);
and U2139 (N_2139,N_1700,N_1789);
and U2140 (N_2140,N_1545,N_1527);
nand U2141 (N_2141,N_1843,N_1094);
and U2142 (N_2142,N_1853,N_1852);
xor U2143 (N_2143,N_1491,N_1486);
nor U2144 (N_2144,N_1032,N_1896);
and U2145 (N_2145,N_1987,N_1558);
nor U2146 (N_2146,N_1587,N_1800);
and U2147 (N_2147,N_1546,N_1836);
nand U2148 (N_2148,N_1115,N_1648);
and U2149 (N_2149,N_1595,N_1304);
xnor U2150 (N_2150,N_1087,N_1879);
and U2151 (N_2151,N_1882,N_1011);
xor U2152 (N_2152,N_1891,N_1467);
nor U2153 (N_2153,N_1137,N_1887);
nand U2154 (N_2154,N_1057,N_1554);
xor U2155 (N_2155,N_1849,N_1633);
or U2156 (N_2156,N_1985,N_1172);
or U2157 (N_2157,N_1167,N_1241);
nand U2158 (N_2158,N_1827,N_1569);
or U2159 (N_2159,N_1004,N_1815);
nor U2160 (N_2160,N_1050,N_1744);
or U2161 (N_2161,N_1048,N_1638);
and U2162 (N_2162,N_1616,N_1239);
xor U2163 (N_2163,N_1630,N_1617);
or U2164 (N_2164,N_1493,N_1735);
nand U2165 (N_2165,N_1964,N_1769);
xor U2166 (N_2166,N_1661,N_1316);
nand U2167 (N_2167,N_1764,N_1023);
nor U2168 (N_2168,N_1537,N_1671);
nor U2169 (N_2169,N_1886,N_1574);
nand U2170 (N_2170,N_1307,N_1428);
nand U2171 (N_2171,N_1979,N_1028);
and U2172 (N_2172,N_1334,N_1676);
or U2173 (N_2173,N_1475,N_1538);
nand U2174 (N_2174,N_1955,N_1046);
nand U2175 (N_2175,N_1995,N_1064);
and U2176 (N_2176,N_1379,N_1583);
nand U2177 (N_2177,N_1510,N_1880);
nand U2178 (N_2178,N_1066,N_1018);
xnor U2179 (N_2179,N_1426,N_1652);
or U2180 (N_2180,N_1009,N_1684);
nor U2181 (N_2181,N_1403,N_1741);
or U2182 (N_2182,N_1157,N_1647);
nand U2183 (N_2183,N_1956,N_1155);
nor U2184 (N_2184,N_1412,N_1708);
nor U2185 (N_2185,N_1754,N_1328);
nand U2186 (N_2186,N_1765,N_1133);
nor U2187 (N_2187,N_1073,N_1300);
nor U2188 (N_2188,N_1422,N_1193);
xor U2189 (N_2189,N_1346,N_1181);
xnor U2190 (N_2190,N_1534,N_1722);
or U2191 (N_2191,N_1969,N_1953);
nand U2192 (N_2192,N_1184,N_1187);
or U2193 (N_2193,N_1981,N_1619);
or U2194 (N_2194,N_1563,N_1145);
and U2195 (N_2195,N_1450,N_1315);
xnor U2196 (N_2196,N_1855,N_1488);
or U2197 (N_2197,N_1771,N_1605);
nand U2198 (N_2198,N_1890,N_1331);
or U2199 (N_2199,N_1550,N_1823);
xnor U2200 (N_2200,N_1806,N_1673);
or U2201 (N_2201,N_1271,N_1542);
nand U2202 (N_2202,N_1954,N_1746);
or U2203 (N_2203,N_1670,N_1490);
or U2204 (N_2204,N_1344,N_1675);
nand U2205 (N_2205,N_1118,N_1399);
and U2206 (N_2206,N_1437,N_1266);
or U2207 (N_2207,N_1851,N_1802);
xnor U2208 (N_2208,N_1062,N_1284);
or U2209 (N_2209,N_1577,N_1795);
xnor U2210 (N_2210,N_1842,N_1093);
xor U2211 (N_2211,N_1317,N_1240);
nor U2212 (N_2212,N_1822,N_1640);
or U2213 (N_2213,N_1857,N_1938);
nor U2214 (N_2214,N_1293,N_1185);
xor U2215 (N_2215,N_1767,N_1161);
or U2216 (N_2216,N_1968,N_1007);
xor U2217 (N_2217,N_1818,N_1479);
xnor U2218 (N_2218,N_1819,N_1003);
or U2219 (N_2219,N_1726,N_1444);
xnor U2220 (N_2220,N_1727,N_1596);
and U2221 (N_2221,N_1643,N_1268);
or U2222 (N_2222,N_1725,N_1045);
and U2223 (N_2223,N_1644,N_1034);
xor U2224 (N_2224,N_1792,N_1793);
nor U2225 (N_2225,N_1373,N_1253);
or U2226 (N_2226,N_1439,N_1481);
and U2227 (N_2227,N_1350,N_1781);
and U2228 (N_2228,N_1365,N_1291);
xor U2229 (N_2229,N_1306,N_1456);
nor U2230 (N_2230,N_1509,N_1392);
xnor U2231 (N_2231,N_1547,N_1443);
xnor U2232 (N_2232,N_1614,N_1310);
or U2233 (N_2233,N_1960,N_1083);
and U2234 (N_2234,N_1001,N_1498);
nor U2235 (N_2235,N_1423,N_1703);
and U2236 (N_2236,N_1507,N_1324);
and U2237 (N_2237,N_1948,N_1332);
xnor U2238 (N_2238,N_1904,N_1747);
nand U2239 (N_2239,N_1257,N_1106);
and U2240 (N_2240,N_1748,N_1950);
and U2241 (N_2241,N_1033,N_1312);
and U2242 (N_2242,N_1734,N_1417);
and U2243 (N_2243,N_1905,N_1680);
nor U2244 (N_2244,N_1225,N_1943);
nand U2245 (N_2245,N_1942,N_1910);
or U2246 (N_2246,N_1687,N_1840);
and U2247 (N_2247,N_1915,N_1602);
nor U2248 (N_2248,N_1845,N_1928);
xor U2249 (N_2249,N_1785,N_1292);
nand U2250 (N_2250,N_1917,N_1362);
xor U2251 (N_2251,N_1353,N_1065);
xor U2252 (N_2252,N_1336,N_1949);
nand U2253 (N_2253,N_1368,N_1142);
nand U2254 (N_2254,N_1606,N_1520);
nor U2255 (N_2255,N_1604,N_1804);
nand U2256 (N_2256,N_1715,N_1457);
and U2257 (N_2257,N_1047,N_1528);
or U2258 (N_2258,N_1937,N_1342);
or U2259 (N_2259,N_1079,N_1831);
nor U2260 (N_2260,N_1594,N_1433);
and U2261 (N_2261,N_1110,N_1760);
and U2262 (N_2262,N_1603,N_1207);
nand U2263 (N_2263,N_1541,N_1530);
xor U2264 (N_2264,N_1551,N_1477);
or U2265 (N_2265,N_1471,N_1686);
nand U2266 (N_2266,N_1348,N_1349);
or U2267 (N_2267,N_1689,N_1540);
nor U2268 (N_2268,N_1084,N_1309);
nand U2269 (N_2269,N_1276,N_1056);
xnor U2270 (N_2270,N_1961,N_1130);
or U2271 (N_2271,N_1474,N_1980);
nand U2272 (N_2272,N_1031,N_1432);
and U2273 (N_2273,N_1641,N_1600);
nand U2274 (N_2274,N_1695,N_1076);
or U2275 (N_2275,N_1288,N_1610);
xnor U2276 (N_2276,N_1885,N_1147);
xnor U2277 (N_2277,N_1278,N_1721);
or U2278 (N_2278,N_1258,N_1730);
and U2279 (N_2279,N_1683,N_1347);
nand U2280 (N_2280,N_1195,N_1211);
nor U2281 (N_2281,N_1000,N_1302);
xnor U2282 (N_2282,N_1957,N_1539);
nor U2283 (N_2283,N_1688,N_1801);
and U2284 (N_2284,N_1404,N_1067);
or U2285 (N_2285,N_1249,N_1672);
nand U2286 (N_2286,N_1327,N_1598);
nand U2287 (N_2287,N_1053,N_1872);
nor U2288 (N_2288,N_1397,N_1357);
nand U2289 (N_2289,N_1448,N_1768);
xnor U2290 (N_2290,N_1729,N_1178);
nor U2291 (N_2291,N_1926,N_1763);
and U2292 (N_2292,N_1008,N_1844);
xnor U2293 (N_2293,N_1370,N_1217);
and U2294 (N_2294,N_1035,N_1743);
nand U2295 (N_2295,N_1835,N_1892);
and U2296 (N_2296,N_1524,N_1838);
nand U2297 (N_2297,N_1657,N_1235);
nor U2298 (N_2298,N_1029,N_1484);
and U2299 (N_2299,N_1553,N_1485);
nor U2300 (N_2300,N_1659,N_1790);
xor U2301 (N_2301,N_1982,N_1501);
or U2302 (N_2302,N_1993,N_1931);
and U2303 (N_2303,N_1496,N_1214);
or U2304 (N_2304,N_1552,N_1152);
xnor U2305 (N_2305,N_1058,N_1135);
nor U2306 (N_2306,N_1237,N_1573);
nand U2307 (N_2307,N_1799,N_1914);
and U2308 (N_2308,N_1320,N_1183);
or U2309 (N_2309,N_1514,N_1994);
or U2310 (N_2310,N_1086,N_1584);
and U2311 (N_2311,N_1608,N_1620);
xnor U2312 (N_2312,N_1168,N_1920);
nand U2313 (N_2313,N_1343,N_1737);
xnor U2314 (N_2314,N_1959,N_1856);
nor U2315 (N_2315,N_1582,N_1777);
or U2316 (N_2316,N_1612,N_1889);
and U2317 (N_2317,N_1704,N_1893);
nor U2318 (N_2318,N_1364,N_1999);
and U2319 (N_2319,N_1816,N_1470);
and U2320 (N_2320,N_1371,N_1642);
or U2321 (N_2321,N_1797,N_1811);
nand U2322 (N_2322,N_1585,N_1129);
nor U2323 (N_2323,N_1311,N_1529);
xnor U2324 (N_2324,N_1044,N_1508);
nor U2325 (N_2325,N_1697,N_1259);
nor U2326 (N_2326,N_1281,N_1144);
and U2327 (N_2327,N_1716,N_1132);
nand U2328 (N_2328,N_1913,N_1020);
and U2329 (N_2329,N_1794,N_1588);
and U2330 (N_2330,N_1085,N_1101);
xor U2331 (N_2331,N_1482,N_1203);
xor U2332 (N_2332,N_1429,N_1839);
nor U2333 (N_2333,N_1772,N_1363);
nor U2334 (N_2334,N_1299,N_1629);
xnor U2335 (N_2335,N_1572,N_1504);
nand U2336 (N_2336,N_1305,N_1779);
or U2337 (N_2337,N_1024,N_1798);
nor U2338 (N_2338,N_1378,N_1273);
nand U2339 (N_2339,N_1092,N_1663);
nand U2340 (N_2340,N_1166,N_1978);
nor U2341 (N_2341,N_1512,N_1098);
and U2342 (N_2342,N_1338,N_1414);
nor U2343 (N_2343,N_1944,N_1164);
nor U2344 (N_2344,N_1631,N_1912);
nor U2345 (N_2345,N_1817,N_1998);
xor U2346 (N_2346,N_1104,N_1100);
nand U2347 (N_2347,N_1270,N_1532);
nand U2348 (N_2348,N_1150,N_1285);
or U2349 (N_2349,N_1375,N_1229);
and U2350 (N_2350,N_1522,N_1634);
nor U2351 (N_2351,N_1731,N_1454);
and U2352 (N_2352,N_1333,N_1369);
nand U2353 (N_2353,N_1072,N_1869);
or U2354 (N_2354,N_1037,N_1078);
or U2355 (N_2355,N_1194,N_1681);
or U2356 (N_2356,N_1678,N_1255);
and U2357 (N_2357,N_1156,N_1436);
xnor U2358 (N_2358,N_1992,N_1866);
or U2359 (N_2359,N_1277,N_1177);
or U2360 (N_2360,N_1390,N_1854);
or U2361 (N_2361,N_1607,N_1796);
nor U2362 (N_2362,N_1038,N_1548);
nand U2363 (N_2363,N_1298,N_1405);
xor U2364 (N_2364,N_1116,N_1873);
or U2365 (N_2365,N_1355,N_1506);
nand U2366 (N_2366,N_1766,N_1366);
or U2367 (N_2367,N_1015,N_1718);
nand U2368 (N_2368,N_1090,N_1113);
nand U2369 (N_2369,N_1775,N_1242);
or U2370 (N_2370,N_1282,N_1502);
or U2371 (N_2371,N_1930,N_1581);
or U2372 (N_2372,N_1517,N_1858);
nor U2373 (N_2373,N_1122,N_1120);
and U2374 (N_2374,N_1231,N_1354);
nand U2375 (N_2375,N_1590,N_1929);
xor U2376 (N_2376,N_1495,N_1927);
or U2377 (N_2377,N_1807,N_1017);
nand U2378 (N_2378,N_1649,N_1463);
and U2379 (N_2379,N_1175,N_1099);
nor U2380 (N_2380,N_1112,N_1778);
xnor U2381 (N_2381,N_1705,N_1932);
xnor U2382 (N_2382,N_1419,N_1589);
xor U2383 (N_2383,N_1865,N_1389);
and U2384 (N_2384,N_1425,N_1163);
nand U2385 (N_2385,N_1323,N_1560);
xor U2386 (N_2386,N_1562,N_1753);
or U2387 (N_2387,N_1898,N_1511);
or U2388 (N_2388,N_1561,N_1216);
nor U2389 (N_2389,N_1224,N_1256);
nand U2390 (N_2390,N_1103,N_1903);
or U2391 (N_2391,N_1318,N_1427);
or U2392 (N_2392,N_1192,N_1160);
xor U2393 (N_2393,N_1597,N_1503);
nand U2394 (N_2394,N_1881,N_1745);
nor U2395 (N_2395,N_1051,N_1837);
or U2396 (N_2396,N_1874,N_1400);
or U2397 (N_2397,N_1902,N_1200);
nor U2398 (N_2398,N_1736,N_1990);
xor U2399 (N_2399,N_1119,N_1335);
nand U2400 (N_2400,N_1279,N_1867);
xnor U2401 (N_2401,N_1213,N_1685);
xor U2402 (N_2402,N_1963,N_1821);
and U2403 (N_2403,N_1526,N_1340);
nor U2404 (N_2404,N_1245,N_1933);
nor U2405 (N_2405,N_1555,N_1234);
nor U2406 (N_2406,N_1713,N_1809);
or U2407 (N_2407,N_1786,N_1918);
or U2408 (N_2408,N_1131,N_1222);
or U2409 (N_2409,N_1468,N_1808);
nor U2410 (N_2410,N_1762,N_1656);
nor U2411 (N_2411,N_1733,N_1650);
nand U2412 (N_2412,N_1483,N_1415);
or U2413 (N_2413,N_1162,N_1232);
or U2414 (N_2414,N_1449,N_1592);
or U2415 (N_2415,N_1319,N_1513);
and U2416 (N_2416,N_1254,N_1940);
nor U2417 (N_2417,N_1651,N_1424);
and U2418 (N_2418,N_1189,N_1627);
or U2419 (N_2419,N_1301,N_1337);
or U2420 (N_2420,N_1859,N_1236);
and U2421 (N_2421,N_1710,N_1626);
nand U2422 (N_2422,N_1043,N_1351);
nor U2423 (N_2423,N_1190,N_1170);
nor U2424 (N_2424,N_1030,N_1923);
and U2425 (N_2425,N_1720,N_1653);
or U2426 (N_2426,N_1012,N_1877);
and U2427 (N_2427,N_1556,N_1198);
and U2428 (N_2428,N_1861,N_1711);
nand U2429 (N_2429,N_1283,N_1696);
nor U2430 (N_2430,N_1976,N_1250);
or U2431 (N_2431,N_1773,N_1409);
xor U2432 (N_2432,N_1141,N_1438);
nand U2433 (N_2433,N_1107,N_1557);
and U2434 (N_2434,N_1783,N_1410);
nor U2435 (N_2435,N_1060,N_1814);
and U2436 (N_2436,N_1567,N_1394);
nor U2437 (N_2437,N_1666,N_1761);
nand U2438 (N_2438,N_1040,N_1210);
nand U2439 (N_2439,N_1314,N_1091);
nor U2440 (N_2440,N_1717,N_1384);
nand U2441 (N_2441,N_1406,N_1041);
nand U2442 (N_2442,N_1223,N_1123);
and U2443 (N_2443,N_1082,N_1473);
or U2444 (N_2444,N_1628,N_1290);
xnor U2445 (N_2445,N_1707,N_1965);
or U2446 (N_2446,N_1868,N_1212);
nor U2447 (N_2447,N_1791,N_1694);
nor U2448 (N_2448,N_1531,N_1758);
and U2449 (N_2449,N_1776,N_1460);
or U2450 (N_2450,N_1939,N_1894);
nor U2451 (N_2451,N_1071,N_1036);
or U2452 (N_2452,N_1997,N_1755);
and U2453 (N_2453,N_1294,N_1226);
nor U2454 (N_2454,N_1829,N_1820);
or U2455 (N_2455,N_1376,N_1442);
and U2456 (N_2456,N_1396,N_1500);
and U2457 (N_2457,N_1313,N_1227);
or U2458 (N_2458,N_1803,N_1637);
or U2459 (N_2459,N_1114,N_1925);
and U2460 (N_2460,N_1421,N_1434);
xnor U2461 (N_2461,N_1411,N_1487);
xnor U2462 (N_2462,N_1264,N_1220);
xnor U2463 (N_2463,N_1660,N_1833);
nor U2464 (N_2464,N_1739,N_1864);
and U2465 (N_2465,N_1499,N_1149);
and U2466 (N_2466,N_1770,N_1952);
or U2467 (N_2467,N_1136,N_1810);
nand U2468 (N_2468,N_1497,N_1451);
nor U2469 (N_2469,N_1664,N_1380);
xnor U2470 (N_2470,N_1121,N_1662);
nand U2471 (N_2471,N_1472,N_1469);
nand U2472 (N_2472,N_1049,N_1321);
or U2473 (N_2473,N_1102,N_1935);
nor U2474 (N_2474,N_1719,N_1430);
nor U2475 (N_2475,N_1159,N_1658);
or U2476 (N_2476,N_1108,N_1655);
xor U2477 (N_2477,N_1260,N_1218);
nor U2478 (N_2478,N_1667,N_1774);
nor U2479 (N_2479,N_1407,N_1812);
xnor U2480 (N_2480,N_1832,N_1014);
and U2481 (N_2481,N_1228,N_1906);
xor U2482 (N_2482,N_1080,N_1677);
nand U2483 (N_2483,N_1435,N_1970);
nor U2484 (N_2484,N_1418,N_1329);
nand U2485 (N_2485,N_1374,N_1749);
nand U2486 (N_2486,N_1458,N_1097);
or U2487 (N_2487,N_1238,N_1973);
nor U2488 (N_2488,N_1139,N_1788);
nand U2489 (N_2489,N_1358,N_1180);
xor U2490 (N_2490,N_1751,N_1752);
or U2491 (N_2491,N_1824,N_1388);
nor U2492 (N_2492,N_1825,N_1544);
xnor U2493 (N_2493,N_1206,N_1308);
xnor U2494 (N_2494,N_1401,N_1621);
nand U2495 (N_2495,N_1381,N_1478);
nand U2496 (N_2496,N_1714,N_1196);
xnor U2497 (N_2497,N_1095,N_1738);
nand U2498 (N_2498,N_1847,N_1580);
or U2499 (N_2499,N_1026,N_1197);
nor U2500 (N_2500,N_1319,N_1942);
and U2501 (N_2501,N_1751,N_1375);
xor U2502 (N_2502,N_1095,N_1250);
and U2503 (N_2503,N_1445,N_1683);
or U2504 (N_2504,N_1044,N_1926);
nor U2505 (N_2505,N_1720,N_1184);
and U2506 (N_2506,N_1092,N_1591);
nand U2507 (N_2507,N_1837,N_1348);
and U2508 (N_2508,N_1727,N_1601);
xnor U2509 (N_2509,N_1385,N_1435);
and U2510 (N_2510,N_1449,N_1361);
or U2511 (N_2511,N_1059,N_1364);
or U2512 (N_2512,N_1555,N_1685);
or U2513 (N_2513,N_1003,N_1326);
nor U2514 (N_2514,N_1605,N_1392);
xor U2515 (N_2515,N_1535,N_1021);
nor U2516 (N_2516,N_1447,N_1685);
and U2517 (N_2517,N_1868,N_1265);
or U2518 (N_2518,N_1646,N_1314);
or U2519 (N_2519,N_1095,N_1105);
or U2520 (N_2520,N_1928,N_1544);
or U2521 (N_2521,N_1276,N_1546);
nand U2522 (N_2522,N_1840,N_1288);
nand U2523 (N_2523,N_1520,N_1481);
xor U2524 (N_2524,N_1503,N_1212);
nand U2525 (N_2525,N_1469,N_1075);
nor U2526 (N_2526,N_1689,N_1330);
and U2527 (N_2527,N_1686,N_1651);
nand U2528 (N_2528,N_1870,N_1076);
nand U2529 (N_2529,N_1191,N_1405);
or U2530 (N_2530,N_1545,N_1319);
nor U2531 (N_2531,N_1499,N_1363);
nor U2532 (N_2532,N_1422,N_1150);
nand U2533 (N_2533,N_1817,N_1154);
nand U2534 (N_2534,N_1999,N_1214);
nand U2535 (N_2535,N_1340,N_1856);
xnor U2536 (N_2536,N_1804,N_1493);
nor U2537 (N_2537,N_1726,N_1571);
and U2538 (N_2538,N_1630,N_1023);
nand U2539 (N_2539,N_1207,N_1172);
nand U2540 (N_2540,N_1511,N_1922);
xor U2541 (N_2541,N_1439,N_1333);
and U2542 (N_2542,N_1189,N_1886);
and U2543 (N_2543,N_1132,N_1113);
or U2544 (N_2544,N_1344,N_1009);
nor U2545 (N_2545,N_1949,N_1148);
nand U2546 (N_2546,N_1526,N_1671);
nand U2547 (N_2547,N_1525,N_1295);
nand U2548 (N_2548,N_1796,N_1689);
nand U2549 (N_2549,N_1389,N_1971);
or U2550 (N_2550,N_1668,N_1117);
nor U2551 (N_2551,N_1653,N_1462);
or U2552 (N_2552,N_1976,N_1209);
nand U2553 (N_2553,N_1634,N_1439);
and U2554 (N_2554,N_1617,N_1257);
or U2555 (N_2555,N_1957,N_1900);
or U2556 (N_2556,N_1248,N_1647);
or U2557 (N_2557,N_1617,N_1354);
or U2558 (N_2558,N_1399,N_1854);
nand U2559 (N_2559,N_1454,N_1986);
nor U2560 (N_2560,N_1778,N_1053);
nor U2561 (N_2561,N_1211,N_1053);
and U2562 (N_2562,N_1010,N_1319);
nor U2563 (N_2563,N_1007,N_1793);
or U2564 (N_2564,N_1881,N_1642);
xnor U2565 (N_2565,N_1462,N_1833);
or U2566 (N_2566,N_1020,N_1485);
or U2567 (N_2567,N_1264,N_1389);
or U2568 (N_2568,N_1297,N_1153);
or U2569 (N_2569,N_1851,N_1746);
and U2570 (N_2570,N_1066,N_1999);
and U2571 (N_2571,N_1612,N_1179);
and U2572 (N_2572,N_1065,N_1981);
nor U2573 (N_2573,N_1729,N_1476);
or U2574 (N_2574,N_1417,N_1888);
xor U2575 (N_2575,N_1462,N_1233);
nand U2576 (N_2576,N_1031,N_1194);
and U2577 (N_2577,N_1818,N_1812);
or U2578 (N_2578,N_1326,N_1002);
nor U2579 (N_2579,N_1622,N_1107);
or U2580 (N_2580,N_1365,N_1222);
xor U2581 (N_2581,N_1949,N_1790);
xor U2582 (N_2582,N_1262,N_1442);
xor U2583 (N_2583,N_1675,N_1825);
and U2584 (N_2584,N_1989,N_1764);
nand U2585 (N_2585,N_1997,N_1576);
nor U2586 (N_2586,N_1563,N_1632);
and U2587 (N_2587,N_1275,N_1123);
xnor U2588 (N_2588,N_1952,N_1731);
nor U2589 (N_2589,N_1959,N_1330);
nor U2590 (N_2590,N_1453,N_1004);
nand U2591 (N_2591,N_1309,N_1187);
nand U2592 (N_2592,N_1686,N_1222);
nand U2593 (N_2593,N_1133,N_1399);
and U2594 (N_2594,N_1794,N_1416);
and U2595 (N_2595,N_1311,N_1042);
and U2596 (N_2596,N_1280,N_1049);
xnor U2597 (N_2597,N_1111,N_1083);
or U2598 (N_2598,N_1100,N_1377);
xnor U2599 (N_2599,N_1408,N_1026);
and U2600 (N_2600,N_1575,N_1548);
nor U2601 (N_2601,N_1682,N_1260);
nand U2602 (N_2602,N_1611,N_1550);
and U2603 (N_2603,N_1683,N_1127);
xnor U2604 (N_2604,N_1812,N_1384);
nor U2605 (N_2605,N_1286,N_1243);
nor U2606 (N_2606,N_1297,N_1653);
nor U2607 (N_2607,N_1584,N_1960);
or U2608 (N_2608,N_1402,N_1351);
nand U2609 (N_2609,N_1929,N_1577);
xor U2610 (N_2610,N_1490,N_1978);
nor U2611 (N_2611,N_1749,N_1751);
nand U2612 (N_2612,N_1778,N_1939);
nand U2613 (N_2613,N_1646,N_1424);
xor U2614 (N_2614,N_1298,N_1500);
nor U2615 (N_2615,N_1448,N_1609);
nand U2616 (N_2616,N_1483,N_1815);
and U2617 (N_2617,N_1376,N_1900);
nor U2618 (N_2618,N_1451,N_1042);
and U2619 (N_2619,N_1569,N_1108);
or U2620 (N_2620,N_1555,N_1504);
and U2621 (N_2621,N_1486,N_1264);
nor U2622 (N_2622,N_1415,N_1368);
or U2623 (N_2623,N_1784,N_1813);
nand U2624 (N_2624,N_1672,N_1998);
or U2625 (N_2625,N_1970,N_1045);
xor U2626 (N_2626,N_1743,N_1903);
or U2627 (N_2627,N_1694,N_1527);
nor U2628 (N_2628,N_1586,N_1972);
and U2629 (N_2629,N_1677,N_1189);
xnor U2630 (N_2630,N_1764,N_1715);
and U2631 (N_2631,N_1862,N_1351);
or U2632 (N_2632,N_1975,N_1476);
nor U2633 (N_2633,N_1135,N_1138);
or U2634 (N_2634,N_1956,N_1949);
nor U2635 (N_2635,N_1120,N_1797);
nor U2636 (N_2636,N_1167,N_1501);
or U2637 (N_2637,N_1317,N_1377);
nor U2638 (N_2638,N_1632,N_1054);
and U2639 (N_2639,N_1480,N_1697);
xor U2640 (N_2640,N_1372,N_1854);
nand U2641 (N_2641,N_1099,N_1420);
and U2642 (N_2642,N_1658,N_1090);
and U2643 (N_2643,N_1485,N_1848);
nor U2644 (N_2644,N_1032,N_1415);
or U2645 (N_2645,N_1085,N_1526);
or U2646 (N_2646,N_1881,N_1330);
nor U2647 (N_2647,N_1122,N_1204);
and U2648 (N_2648,N_1500,N_1921);
nor U2649 (N_2649,N_1063,N_1368);
nor U2650 (N_2650,N_1565,N_1294);
and U2651 (N_2651,N_1106,N_1275);
nand U2652 (N_2652,N_1834,N_1923);
and U2653 (N_2653,N_1720,N_1778);
xor U2654 (N_2654,N_1199,N_1419);
or U2655 (N_2655,N_1565,N_1677);
nor U2656 (N_2656,N_1248,N_1773);
or U2657 (N_2657,N_1138,N_1580);
or U2658 (N_2658,N_1658,N_1491);
nor U2659 (N_2659,N_1058,N_1714);
xnor U2660 (N_2660,N_1310,N_1553);
nand U2661 (N_2661,N_1610,N_1765);
nand U2662 (N_2662,N_1086,N_1953);
and U2663 (N_2663,N_1457,N_1742);
nand U2664 (N_2664,N_1349,N_1021);
and U2665 (N_2665,N_1799,N_1868);
xnor U2666 (N_2666,N_1169,N_1234);
nand U2667 (N_2667,N_1963,N_1105);
xnor U2668 (N_2668,N_1243,N_1320);
or U2669 (N_2669,N_1190,N_1009);
or U2670 (N_2670,N_1661,N_1752);
or U2671 (N_2671,N_1529,N_1030);
nand U2672 (N_2672,N_1300,N_1601);
or U2673 (N_2673,N_1862,N_1559);
or U2674 (N_2674,N_1128,N_1662);
nor U2675 (N_2675,N_1930,N_1061);
nor U2676 (N_2676,N_1167,N_1872);
nor U2677 (N_2677,N_1033,N_1335);
nand U2678 (N_2678,N_1746,N_1646);
xor U2679 (N_2679,N_1348,N_1286);
nand U2680 (N_2680,N_1944,N_1705);
and U2681 (N_2681,N_1219,N_1052);
nor U2682 (N_2682,N_1331,N_1302);
or U2683 (N_2683,N_1655,N_1352);
nor U2684 (N_2684,N_1650,N_1073);
or U2685 (N_2685,N_1945,N_1839);
xor U2686 (N_2686,N_1861,N_1886);
nor U2687 (N_2687,N_1752,N_1302);
nand U2688 (N_2688,N_1681,N_1927);
or U2689 (N_2689,N_1078,N_1809);
nor U2690 (N_2690,N_1675,N_1171);
and U2691 (N_2691,N_1952,N_1092);
and U2692 (N_2692,N_1531,N_1274);
xor U2693 (N_2693,N_1665,N_1040);
or U2694 (N_2694,N_1989,N_1081);
nand U2695 (N_2695,N_1615,N_1268);
or U2696 (N_2696,N_1947,N_1087);
and U2697 (N_2697,N_1910,N_1607);
and U2698 (N_2698,N_1641,N_1325);
and U2699 (N_2699,N_1995,N_1163);
or U2700 (N_2700,N_1935,N_1719);
nand U2701 (N_2701,N_1754,N_1427);
or U2702 (N_2702,N_1333,N_1198);
or U2703 (N_2703,N_1730,N_1386);
or U2704 (N_2704,N_1934,N_1532);
nor U2705 (N_2705,N_1548,N_1790);
and U2706 (N_2706,N_1418,N_1723);
xnor U2707 (N_2707,N_1890,N_1797);
nand U2708 (N_2708,N_1936,N_1483);
and U2709 (N_2709,N_1999,N_1463);
nor U2710 (N_2710,N_1649,N_1146);
nor U2711 (N_2711,N_1784,N_1311);
or U2712 (N_2712,N_1757,N_1952);
xor U2713 (N_2713,N_1028,N_1504);
nor U2714 (N_2714,N_1976,N_1740);
nand U2715 (N_2715,N_1530,N_1761);
and U2716 (N_2716,N_1924,N_1185);
and U2717 (N_2717,N_1101,N_1296);
nand U2718 (N_2718,N_1221,N_1803);
or U2719 (N_2719,N_1340,N_1549);
and U2720 (N_2720,N_1511,N_1643);
and U2721 (N_2721,N_1760,N_1145);
and U2722 (N_2722,N_1583,N_1838);
or U2723 (N_2723,N_1336,N_1947);
nand U2724 (N_2724,N_1666,N_1937);
nand U2725 (N_2725,N_1718,N_1621);
or U2726 (N_2726,N_1306,N_1643);
nor U2727 (N_2727,N_1218,N_1287);
and U2728 (N_2728,N_1185,N_1710);
xnor U2729 (N_2729,N_1482,N_1014);
nor U2730 (N_2730,N_1326,N_1738);
xnor U2731 (N_2731,N_1160,N_1503);
nand U2732 (N_2732,N_1317,N_1445);
nor U2733 (N_2733,N_1139,N_1217);
and U2734 (N_2734,N_1092,N_1344);
and U2735 (N_2735,N_1387,N_1013);
nor U2736 (N_2736,N_1785,N_1263);
nand U2737 (N_2737,N_1311,N_1438);
or U2738 (N_2738,N_1708,N_1068);
and U2739 (N_2739,N_1397,N_1844);
nor U2740 (N_2740,N_1885,N_1460);
or U2741 (N_2741,N_1226,N_1908);
xor U2742 (N_2742,N_1313,N_1878);
or U2743 (N_2743,N_1110,N_1115);
xor U2744 (N_2744,N_1861,N_1007);
nor U2745 (N_2745,N_1106,N_1129);
and U2746 (N_2746,N_1295,N_1679);
and U2747 (N_2747,N_1820,N_1684);
xor U2748 (N_2748,N_1739,N_1317);
and U2749 (N_2749,N_1228,N_1501);
nand U2750 (N_2750,N_1674,N_1268);
nand U2751 (N_2751,N_1090,N_1373);
nor U2752 (N_2752,N_1582,N_1616);
nor U2753 (N_2753,N_1206,N_1546);
or U2754 (N_2754,N_1856,N_1464);
and U2755 (N_2755,N_1071,N_1239);
and U2756 (N_2756,N_1267,N_1951);
xnor U2757 (N_2757,N_1252,N_1972);
or U2758 (N_2758,N_1919,N_1627);
or U2759 (N_2759,N_1232,N_1003);
nor U2760 (N_2760,N_1334,N_1628);
and U2761 (N_2761,N_1883,N_1848);
or U2762 (N_2762,N_1205,N_1696);
xnor U2763 (N_2763,N_1608,N_1673);
xor U2764 (N_2764,N_1840,N_1503);
nand U2765 (N_2765,N_1636,N_1248);
xnor U2766 (N_2766,N_1895,N_1802);
xnor U2767 (N_2767,N_1418,N_1122);
or U2768 (N_2768,N_1166,N_1078);
nor U2769 (N_2769,N_1316,N_1581);
nand U2770 (N_2770,N_1480,N_1032);
nor U2771 (N_2771,N_1803,N_1207);
or U2772 (N_2772,N_1539,N_1285);
and U2773 (N_2773,N_1613,N_1208);
xnor U2774 (N_2774,N_1498,N_1106);
xor U2775 (N_2775,N_1732,N_1484);
nor U2776 (N_2776,N_1788,N_1624);
and U2777 (N_2777,N_1984,N_1371);
and U2778 (N_2778,N_1454,N_1870);
and U2779 (N_2779,N_1927,N_1582);
or U2780 (N_2780,N_1213,N_1128);
nand U2781 (N_2781,N_1557,N_1572);
and U2782 (N_2782,N_1734,N_1181);
and U2783 (N_2783,N_1328,N_1037);
nand U2784 (N_2784,N_1677,N_1771);
nand U2785 (N_2785,N_1785,N_1807);
or U2786 (N_2786,N_1679,N_1344);
and U2787 (N_2787,N_1705,N_1893);
xnor U2788 (N_2788,N_1602,N_1175);
nor U2789 (N_2789,N_1836,N_1093);
or U2790 (N_2790,N_1800,N_1742);
nand U2791 (N_2791,N_1581,N_1943);
and U2792 (N_2792,N_1217,N_1967);
and U2793 (N_2793,N_1605,N_1584);
nor U2794 (N_2794,N_1871,N_1402);
nor U2795 (N_2795,N_1122,N_1821);
nor U2796 (N_2796,N_1659,N_1030);
and U2797 (N_2797,N_1908,N_1832);
nor U2798 (N_2798,N_1663,N_1909);
or U2799 (N_2799,N_1467,N_1150);
xor U2800 (N_2800,N_1342,N_1847);
nand U2801 (N_2801,N_1242,N_1005);
xnor U2802 (N_2802,N_1408,N_1165);
nor U2803 (N_2803,N_1893,N_1708);
xnor U2804 (N_2804,N_1745,N_1243);
xnor U2805 (N_2805,N_1887,N_1207);
xor U2806 (N_2806,N_1801,N_1297);
nor U2807 (N_2807,N_1457,N_1877);
xnor U2808 (N_2808,N_1584,N_1326);
or U2809 (N_2809,N_1328,N_1257);
nor U2810 (N_2810,N_1676,N_1579);
xor U2811 (N_2811,N_1730,N_1328);
nor U2812 (N_2812,N_1549,N_1032);
or U2813 (N_2813,N_1309,N_1229);
and U2814 (N_2814,N_1002,N_1234);
nor U2815 (N_2815,N_1433,N_1036);
xnor U2816 (N_2816,N_1884,N_1216);
nor U2817 (N_2817,N_1779,N_1091);
xor U2818 (N_2818,N_1913,N_1667);
and U2819 (N_2819,N_1909,N_1169);
nand U2820 (N_2820,N_1233,N_1290);
nand U2821 (N_2821,N_1333,N_1306);
nand U2822 (N_2822,N_1455,N_1162);
nor U2823 (N_2823,N_1414,N_1086);
xor U2824 (N_2824,N_1561,N_1223);
nor U2825 (N_2825,N_1343,N_1240);
and U2826 (N_2826,N_1945,N_1624);
and U2827 (N_2827,N_1626,N_1965);
or U2828 (N_2828,N_1623,N_1079);
or U2829 (N_2829,N_1288,N_1487);
xnor U2830 (N_2830,N_1733,N_1740);
nand U2831 (N_2831,N_1929,N_1436);
and U2832 (N_2832,N_1505,N_1501);
nor U2833 (N_2833,N_1097,N_1727);
nor U2834 (N_2834,N_1094,N_1385);
and U2835 (N_2835,N_1292,N_1067);
nor U2836 (N_2836,N_1101,N_1199);
nand U2837 (N_2837,N_1024,N_1182);
xnor U2838 (N_2838,N_1250,N_1254);
nand U2839 (N_2839,N_1738,N_1247);
and U2840 (N_2840,N_1257,N_1299);
xnor U2841 (N_2841,N_1876,N_1307);
xor U2842 (N_2842,N_1482,N_1933);
nor U2843 (N_2843,N_1537,N_1316);
nand U2844 (N_2844,N_1242,N_1346);
nand U2845 (N_2845,N_1885,N_1980);
or U2846 (N_2846,N_1611,N_1233);
nand U2847 (N_2847,N_1846,N_1586);
and U2848 (N_2848,N_1578,N_1373);
and U2849 (N_2849,N_1215,N_1085);
nand U2850 (N_2850,N_1365,N_1165);
xor U2851 (N_2851,N_1967,N_1139);
nor U2852 (N_2852,N_1535,N_1903);
nor U2853 (N_2853,N_1411,N_1062);
or U2854 (N_2854,N_1280,N_1072);
nor U2855 (N_2855,N_1279,N_1050);
nand U2856 (N_2856,N_1998,N_1226);
or U2857 (N_2857,N_1924,N_1225);
nand U2858 (N_2858,N_1369,N_1013);
nor U2859 (N_2859,N_1358,N_1094);
and U2860 (N_2860,N_1448,N_1118);
or U2861 (N_2861,N_1608,N_1987);
nand U2862 (N_2862,N_1005,N_1654);
nand U2863 (N_2863,N_1032,N_1323);
nor U2864 (N_2864,N_1823,N_1300);
nor U2865 (N_2865,N_1888,N_1833);
or U2866 (N_2866,N_1699,N_1950);
and U2867 (N_2867,N_1316,N_1355);
nor U2868 (N_2868,N_1374,N_1402);
or U2869 (N_2869,N_1835,N_1829);
nand U2870 (N_2870,N_1675,N_1823);
xnor U2871 (N_2871,N_1427,N_1209);
nor U2872 (N_2872,N_1080,N_1819);
and U2873 (N_2873,N_1636,N_1770);
xor U2874 (N_2874,N_1929,N_1130);
and U2875 (N_2875,N_1817,N_1052);
nand U2876 (N_2876,N_1736,N_1937);
and U2877 (N_2877,N_1522,N_1611);
nor U2878 (N_2878,N_1580,N_1713);
nor U2879 (N_2879,N_1737,N_1892);
nor U2880 (N_2880,N_1268,N_1445);
nand U2881 (N_2881,N_1943,N_1130);
nand U2882 (N_2882,N_1111,N_1185);
nor U2883 (N_2883,N_1671,N_1513);
xor U2884 (N_2884,N_1819,N_1651);
or U2885 (N_2885,N_1841,N_1904);
nand U2886 (N_2886,N_1479,N_1916);
xnor U2887 (N_2887,N_1852,N_1960);
nor U2888 (N_2888,N_1014,N_1751);
nand U2889 (N_2889,N_1201,N_1053);
nand U2890 (N_2890,N_1332,N_1777);
nor U2891 (N_2891,N_1276,N_1094);
nor U2892 (N_2892,N_1842,N_1969);
nand U2893 (N_2893,N_1404,N_1008);
or U2894 (N_2894,N_1873,N_1639);
and U2895 (N_2895,N_1522,N_1711);
xnor U2896 (N_2896,N_1453,N_1023);
or U2897 (N_2897,N_1026,N_1132);
nand U2898 (N_2898,N_1529,N_1367);
or U2899 (N_2899,N_1976,N_1653);
or U2900 (N_2900,N_1542,N_1913);
nand U2901 (N_2901,N_1406,N_1352);
and U2902 (N_2902,N_1261,N_1434);
xor U2903 (N_2903,N_1541,N_1501);
and U2904 (N_2904,N_1684,N_1218);
nor U2905 (N_2905,N_1612,N_1724);
and U2906 (N_2906,N_1896,N_1625);
nor U2907 (N_2907,N_1533,N_1648);
or U2908 (N_2908,N_1670,N_1306);
nor U2909 (N_2909,N_1675,N_1128);
nor U2910 (N_2910,N_1906,N_1445);
nand U2911 (N_2911,N_1028,N_1425);
nor U2912 (N_2912,N_1261,N_1489);
xor U2913 (N_2913,N_1693,N_1662);
nand U2914 (N_2914,N_1827,N_1205);
or U2915 (N_2915,N_1795,N_1303);
nand U2916 (N_2916,N_1923,N_1727);
or U2917 (N_2917,N_1523,N_1316);
nor U2918 (N_2918,N_1565,N_1644);
nand U2919 (N_2919,N_1211,N_1581);
xnor U2920 (N_2920,N_1063,N_1516);
nand U2921 (N_2921,N_1078,N_1686);
and U2922 (N_2922,N_1556,N_1831);
and U2923 (N_2923,N_1943,N_1527);
nand U2924 (N_2924,N_1589,N_1813);
nor U2925 (N_2925,N_1393,N_1778);
xor U2926 (N_2926,N_1005,N_1442);
and U2927 (N_2927,N_1111,N_1261);
xor U2928 (N_2928,N_1712,N_1401);
xor U2929 (N_2929,N_1810,N_1490);
and U2930 (N_2930,N_1404,N_1004);
xor U2931 (N_2931,N_1962,N_1345);
nor U2932 (N_2932,N_1945,N_1715);
xor U2933 (N_2933,N_1693,N_1998);
nor U2934 (N_2934,N_1948,N_1304);
or U2935 (N_2935,N_1606,N_1235);
or U2936 (N_2936,N_1517,N_1980);
xor U2937 (N_2937,N_1869,N_1745);
and U2938 (N_2938,N_1247,N_1604);
and U2939 (N_2939,N_1755,N_1885);
xor U2940 (N_2940,N_1599,N_1124);
nand U2941 (N_2941,N_1111,N_1836);
xor U2942 (N_2942,N_1323,N_1759);
nor U2943 (N_2943,N_1572,N_1531);
xnor U2944 (N_2944,N_1801,N_1935);
or U2945 (N_2945,N_1656,N_1458);
nand U2946 (N_2946,N_1964,N_1330);
and U2947 (N_2947,N_1095,N_1544);
nand U2948 (N_2948,N_1326,N_1518);
nor U2949 (N_2949,N_1149,N_1298);
and U2950 (N_2950,N_1206,N_1228);
and U2951 (N_2951,N_1009,N_1027);
nand U2952 (N_2952,N_1474,N_1731);
nor U2953 (N_2953,N_1309,N_1616);
xor U2954 (N_2954,N_1011,N_1776);
and U2955 (N_2955,N_1342,N_1501);
or U2956 (N_2956,N_1930,N_1626);
xor U2957 (N_2957,N_1684,N_1855);
or U2958 (N_2958,N_1276,N_1538);
nor U2959 (N_2959,N_1334,N_1585);
nand U2960 (N_2960,N_1973,N_1867);
and U2961 (N_2961,N_1634,N_1677);
nand U2962 (N_2962,N_1843,N_1326);
xnor U2963 (N_2963,N_1072,N_1396);
nor U2964 (N_2964,N_1878,N_1269);
nand U2965 (N_2965,N_1534,N_1238);
nand U2966 (N_2966,N_1364,N_1486);
and U2967 (N_2967,N_1911,N_1135);
and U2968 (N_2968,N_1374,N_1797);
nor U2969 (N_2969,N_1172,N_1496);
or U2970 (N_2970,N_1438,N_1325);
xnor U2971 (N_2971,N_1975,N_1438);
or U2972 (N_2972,N_1110,N_1965);
or U2973 (N_2973,N_1490,N_1000);
or U2974 (N_2974,N_1477,N_1181);
nand U2975 (N_2975,N_1100,N_1590);
and U2976 (N_2976,N_1570,N_1503);
xor U2977 (N_2977,N_1324,N_1697);
nand U2978 (N_2978,N_1576,N_1312);
or U2979 (N_2979,N_1946,N_1456);
nand U2980 (N_2980,N_1682,N_1101);
or U2981 (N_2981,N_1373,N_1006);
and U2982 (N_2982,N_1421,N_1752);
and U2983 (N_2983,N_1506,N_1950);
nor U2984 (N_2984,N_1470,N_1915);
xor U2985 (N_2985,N_1556,N_1143);
or U2986 (N_2986,N_1312,N_1765);
nand U2987 (N_2987,N_1850,N_1912);
xnor U2988 (N_2988,N_1009,N_1253);
or U2989 (N_2989,N_1598,N_1058);
nor U2990 (N_2990,N_1641,N_1119);
xnor U2991 (N_2991,N_1350,N_1877);
and U2992 (N_2992,N_1894,N_1241);
xnor U2993 (N_2993,N_1669,N_1839);
and U2994 (N_2994,N_1843,N_1428);
and U2995 (N_2995,N_1933,N_1587);
xnor U2996 (N_2996,N_1617,N_1051);
xor U2997 (N_2997,N_1360,N_1437);
and U2998 (N_2998,N_1067,N_1886);
xnor U2999 (N_2999,N_1559,N_1484);
nor U3000 (N_3000,N_2587,N_2900);
nor U3001 (N_3001,N_2064,N_2202);
xnor U3002 (N_3002,N_2463,N_2426);
xnor U3003 (N_3003,N_2005,N_2114);
or U3004 (N_3004,N_2142,N_2875);
nor U3005 (N_3005,N_2550,N_2646);
nand U3006 (N_3006,N_2304,N_2641);
nor U3007 (N_3007,N_2205,N_2155);
or U3008 (N_3008,N_2312,N_2097);
nor U3009 (N_3009,N_2422,N_2280);
or U3010 (N_3010,N_2532,N_2291);
xor U3011 (N_3011,N_2621,N_2166);
nor U3012 (N_3012,N_2605,N_2937);
nor U3013 (N_3013,N_2040,N_2909);
nor U3014 (N_3014,N_2810,N_2228);
and U3015 (N_3015,N_2065,N_2079);
xnor U3016 (N_3016,N_2635,N_2598);
nand U3017 (N_3017,N_2666,N_2823);
xor U3018 (N_3018,N_2632,N_2735);
xor U3019 (N_3019,N_2583,N_2405);
nand U3020 (N_3020,N_2989,N_2962);
or U3021 (N_3021,N_2767,N_2969);
nand U3022 (N_3022,N_2763,N_2894);
xnor U3023 (N_3023,N_2792,N_2683);
nand U3024 (N_3024,N_2068,N_2663);
nor U3025 (N_3025,N_2163,N_2596);
xor U3026 (N_3026,N_2362,N_2251);
or U3027 (N_3027,N_2082,N_2331);
and U3028 (N_3028,N_2401,N_2180);
nor U3029 (N_3029,N_2599,N_2776);
or U3030 (N_3030,N_2582,N_2730);
nor U3031 (N_3031,N_2600,N_2073);
or U3032 (N_3032,N_2066,N_2519);
nor U3033 (N_3033,N_2870,N_2328);
nor U3034 (N_3034,N_2393,N_2160);
xor U3035 (N_3035,N_2963,N_2015);
nand U3036 (N_3036,N_2334,N_2866);
and U3037 (N_3037,N_2498,N_2306);
xor U3038 (N_3038,N_2300,N_2522);
xnor U3039 (N_3039,N_2565,N_2702);
nor U3040 (N_3040,N_2281,N_2619);
or U3041 (N_3041,N_2764,N_2929);
xor U3042 (N_3042,N_2211,N_2754);
xnor U3043 (N_3043,N_2640,N_2800);
xor U3044 (N_3044,N_2938,N_2338);
nor U3045 (N_3045,N_2671,N_2784);
nor U3046 (N_3046,N_2111,N_2419);
and U3047 (N_3047,N_2499,N_2928);
and U3048 (N_3048,N_2289,N_2464);
xor U3049 (N_3049,N_2225,N_2597);
or U3050 (N_3050,N_2379,N_2690);
xor U3051 (N_3051,N_2112,N_2162);
xor U3052 (N_3052,N_2684,N_2503);
xor U3053 (N_3053,N_2442,N_2271);
nand U3054 (N_3054,N_2734,N_2543);
nand U3055 (N_3055,N_2124,N_2725);
nand U3056 (N_3056,N_2382,N_2974);
nor U3057 (N_3057,N_2330,N_2260);
nor U3058 (N_3058,N_2631,N_2778);
xor U3059 (N_3059,N_2395,N_2006);
and U3060 (N_3060,N_2210,N_2383);
or U3061 (N_3061,N_2060,N_2854);
xnor U3062 (N_3062,N_2757,N_2022);
nor U3063 (N_3063,N_2692,N_2761);
nand U3064 (N_3064,N_2732,N_2973);
nor U3065 (N_3065,N_2525,N_2452);
xnor U3066 (N_3066,N_2749,N_2988);
nand U3067 (N_3067,N_2174,N_2448);
nand U3068 (N_3068,N_2831,N_2562);
or U3069 (N_3069,N_2195,N_2775);
nor U3070 (N_3070,N_2638,N_2373);
or U3071 (N_3071,N_2737,N_2558);
nand U3072 (N_3072,N_2615,N_2071);
nand U3073 (N_3073,N_2341,N_2453);
xor U3074 (N_3074,N_2359,N_2361);
or U3075 (N_3075,N_2356,N_2964);
nand U3076 (N_3076,N_2493,N_2482);
xnor U3077 (N_3077,N_2956,N_2440);
and U3078 (N_3078,N_2648,N_2552);
or U3079 (N_3079,N_2380,N_2283);
nand U3080 (N_3080,N_2669,N_2461);
and U3081 (N_3081,N_2850,N_2184);
nand U3082 (N_3082,N_2220,N_2152);
nor U3083 (N_3083,N_2096,N_2591);
or U3084 (N_3084,N_2141,N_2892);
nor U3085 (N_3085,N_2520,N_2122);
or U3086 (N_3086,N_2949,N_2206);
or U3087 (N_3087,N_2898,N_2910);
or U3088 (N_3088,N_2150,N_2798);
or U3089 (N_3089,N_2420,N_2433);
nand U3090 (N_3090,N_2069,N_2901);
or U3091 (N_3091,N_2710,N_2010);
nor U3092 (N_3092,N_2801,N_2149);
or U3093 (N_3093,N_2247,N_2078);
nor U3094 (N_3094,N_2233,N_2610);
nand U3095 (N_3095,N_2877,N_2335);
nor U3096 (N_3096,N_2604,N_2906);
nor U3097 (N_3097,N_2527,N_2945);
xnor U3098 (N_3098,N_2513,N_2665);
nand U3099 (N_3099,N_2930,N_2835);
or U3100 (N_3100,N_2363,N_2743);
and U3101 (N_3101,N_2042,N_2480);
nor U3102 (N_3102,N_2360,N_2645);
nor U3103 (N_3103,N_2662,N_2000);
xnor U3104 (N_3104,N_2779,N_2344);
or U3105 (N_3105,N_2614,N_2712);
nor U3106 (N_3106,N_2869,N_2209);
or U3107 (N_3107,N_2644,N_2018);
xnor U3108 (N_3108,N_2534,N_2146);
and U3109 (N_3109,N_2127,N_2014);
and U3110 (N_3110,N_2218,N_2549);
xor U3111 (N_3111,N_2790,N_2516);
and U3112 (N_3112,N_2178,N_2102);
xor U3113 (N_3113,N_2609,N_2001);
or U3114 (N_3114,N_2287,N_2862);
nor U3115 (N_3115,N_2240,N_2385);
xor U3116 (N_3116,N_2595,N_2884);
and U3117 (N_3117,N_2853,N_2704);
and U3118 (N_3118,N_2315,N_2540);
nand U3119 (N_3119,N_2512,N_2313);
nor U3120 (N_3120,N_2242,N_2417);
or U3121 (N_3121,N_2826,N_2657);
xor U3122 (N_3122,N_2758,N_2517);
xor U3123 (N_3123,N_2264,N_2714);
and U3124 (N_3124,N_2837,N_2849);
and U3125 (N_3125,N_2311,N_2818);
or U3126 (N_3126,N_2366,N_2027);
nand U3127 (N_3127,N_2469,N_2394);
nor U3128 (N_3128,N_2840,N_2972);
xor U3129 (N_3129,N_2941,N_2308);
and U3130 (N_3130,N_2353,N_2979);
xor U3131 (N_3131,N_2090,N_2059);
or U3132 (N_3132,N_2694,N_2556);
and U3133 (N_3133,N_2670,N_2724);
nor U3134 (N_3134,N_2773,N_2617);
and U3135 (N_3135,N_2667,N_2489);
xor U3136 (N_3136,N_2542,N_2098);
and U3137 (N_3137,N_2867,N_2926);
or U3138 (N_3138,N_2302,N_2076);
nand U3139 (N_3139,N_2968,N_2893);
xnor U3140 (N_3140,N_2895,N_2736);
xnor U3141 (N_3141,N_2033,N_2113);
xor U3142 (N_3142,N_2653,N_2285);
xnor U3143 (N_3143,N_2744,N_2584);
xnor U3144 (N_3144,N_2301,N_2045);
xor U3145 (N_3145,N_2157,N_2212);
nor U3146 (N_3146,N_2838,N_2351);
xnor U3147 (N_3147,N_2423,N_2728);
and U3148 (N_3148,N_2381,N_2117);
nand U3149 (N_3149,N_2686,N_2899);
or U3150 (N_3150,N_2942,N_2204);
or U3151 (N_3151,N_2004,N_2881);
xnor U3152 (N_3152,N_2269,N_2797);
xnor U3153 (N_3153,N_2093,N_2820);
nor U3154 (N_3154,N_2507,N_2459);
xor U3155 (N_3155,N_2267,N_2530);
nand U3156 (N_3156,N_2878,N_2274);
and U3157 (N_3157,N_2265,N_2496);
and U3158 (N_3158,N_2024,N_2538);
and U3159 (N_3159,N_2606,N_2780);
and U3160 (N_3160,N_2647,N_2032);
and U3161 (N_3161,N_2414,N_2103);
nor U3162 (N_3162,N_2276,N_2343);
or U3163 (N_3163,N_2055,N_2321);
xor U3164 (N_3164,N_2703,N_2116);
and U3165 (N_3165,N_2721,N_2664);
and U3166 (N_3166,N_2486,N_2882);
nor U3167 (N_3167,N_2782,N_2412);
nand U3168 (N_3168,N_2954,N_2025);
xnor U3169 (N_3169,N_2396,N_2947);
or U3170 (N_3170,N_2056,N_2087);
or U3171 (N_3171,N_2063,N_2234);
and U3172 (N_3172,N_2544,N_2563);
or U3173 (N_3173,N_2475,N_2326);
or U3174 (N_3174,N_2258,N_2151);
xor U3175 (N_3175,N_2526,N_2914);
nor U3176 (N_3176,N_2781,N_2250);
nor U3177 (N_3177,N_2659,N_2249);
and U3178 (N_3178,N_2227,N_2660);
nand U3179 (N_3179,N_2633,N_2768);
nor U3180 (N_3180,N_2975,N_2727);
xor U3181 (N_3181,N_2329,N_2462);
and U3182 (N_3182,N_2788,N_2237);
xnor U3183 (N_3183,N_2245,N_2483);
nand U3184 (N_3184,N_2751,N_2812);
or U3185 (N_3185,N_2514,N_2698);
and U3186 (N_3186,N_2934,N_2841);
or U3187 (N_3187,N_2791,N_2913);
nand U3188 (N_3188,N_2369,N_2197);
nand U3189 (N_3189,N_2348,N_2083);
xor U3190 (N_3190,N_2454,N_2924);
xnor U3191 (N_3191,N_2700,N_2794);
nand U3192 (N_3192,N_2357,N_2580);
and U3193 (N_3193,N_2750,N_2084);
nor U3194 (N_3194,N_2572,N_2175);
nand U3195 (N_3195,N_2203,N_2611);
or U3196 (N_3196,N_2575,N_2322);
xnor U3197 (N_3197,N_2731,N_2559);
nor U3198 (N_3198,N_2777,N_2846);
nor U3199 (N_3199,N_2325,N_2783);
and U3200 (N_3200,N_2697,N_2089);
nand U3201 (N_3201,N_2997,N_2957);
nand U3202 (N_3202,N_2772,N_2188);
and U3203 (N_3203,N_2137,N_2923);
and U3204 (N_3204,N_2257,N_2613);
or U3205 (N_3205,N_2072,N_2115);
nor U3206 (N_3206,N_2432,N_2983);
and U3207 (N_3207,N_2502,N_2239);
or U3208 (N_3208,N_2477,N_2421);
or U3209 (N_3209,N_2649,N_2017);
nand U3210 (N_3210,N_2876,N_2009);
or U3211 (N_3211,N_2711,N_2392);
nor U3212 (N_3212,N_2349,N_2872);
and U3213 (N_3213,N_2156,N_2282);
nor U3214 (N_3214,N_2323,N_2446);
or U3215 (N_3215,N_2140,N_2588);
and U3216 (N_3216,N_2165,N_2101);
or U3217 (N_3217,N_2198,N_2658);
nand U3218 (N_3218,N_2678,N_2745);
or U3219 (N_3219,N_2216,N_2139);
nand U3220 (N_3220,N_2656,N_2438);
or U3221 (N_3221,N_2147,N_2034);
xnor U3222 (N_3222,N_2377,N_2965);
and U3223 (N_3223,N_2427,N_2762);
nor U3224 (N_3224,N_2629,N_2011);
xnor U3225 (N_3225,N_2707,N_2418);
and U3226 (N_3226,N_2295,N_2691);
and U3227 (N_3227,N_2521,N_2386);
and U3228 (N_3228,N_2852,N_2564);
nor U3229 (N_3229,N_2317,N_2278);
nor U3230 (N_3230,N_2290,N_2766);
xnor U3231 (N_3231,N_2046,N_2708);
nand U3232 (N_3232,N_2129,N_2879);
or U3233 (N_3233,N_2814,N_2201);
nand U3234 (N_3234,N_2793,N_2890);
xnor U3235 (N_3235,N_2316,N_2029);
nand U3236 (N_3236,N_2693,N_2885);
nand U3237 (N_3237,N_2471,N_2307);
xnor U3238 (N_3238,N_2171,N_2808);
xor U3239 (N_3239,N_2019,N_2787);
nor U3240 (N_3240,N_2048,N_2026);
nand U3241 (N_3241,N_2752,N_2504);
and U3242 (N_3242,N_2581,N_2539);
nand U3243 (N_3243,N_2943,N_2829);
xor U3244 (N_3244,N_2603,N_2524);
and U3245 (N_3245,N_2235,N_2608);
nand U3246 (N_3246,N_2528,N_2679);
nand U3247 (N_3247,N_2976,N_2618);
nor U3248 (N_3248,N_2789,N_2476);
and U3249 (N_3249,N_2230,N_2570);
nand U3250 (N_3250,N_2490,N_2813);
or U3251 (N_3251,N_2346,N_2560);
nor U3252 (N_3252,N_2626,N_2992);
and U3253 (N_3253,N_2991,N_2863);
xor U3254 (N_3254,N_2465,N_2181);
nor U3255 (N_3255,N_2713,N_2927);
xnor U3256 (N_3256,N_2824,N_2051);
and U3257 (N_3257,N_2441,N_2460);
nor U3258 (N_3258,N_2410,N_2008);
nor U3259 (N_3259,N_2428,N_2436);
nand U3260 (N_3260,N_2158,N_2053);
xnor U3261 (N_3261,N_2320,N_2121);
xor U3262 (N_3262,N_2594,N_2905);
or U3263 (N_3263,N_2642,N_2990);
and U3264 (N_3264,N_2057,N_2447);
nand U3265 (N_3265,N_2263,N_2261);
or U3266 (N_3266,N_2718,N_2795);
xor U3267 (N_3267,N_2858,N_2554);
xnor U3268 (N_3268,N_2485,N_2845);
nor U3269 (N_3269,N_2848,N_2553);
and U3270 (N_3270,N_2709,N_2856);
nor U3271 (N_3271,N_2297,N_2571);
xnor U3272 (N_3272,N_2303,N_2996);
nand U3273 (N_3273,N_2016,N_2630);
and U3274 (N_3274,N_2473,N_2830);
nor U3275 (N_3275,N_2479,N_2925);
nor U3276 (N_3276,N_2387,N_2628);
and U3277 (N_3277,N_2370,N_2807);
nand U3278 (N_3278,N_2319,N_2193);
nand U3279 (N_3279,N_2739,N_2953);
and U3280 (N_3280,N_2434,N_2847);
xnor U3281 (N_3281,N_2756,N_2529);
nand U3282 (N_3282,N_2173,N_2602);
xor U3283 (N_3283,N_2148,N_2196);
or U3284 (N_3284,N_2951,N_2105);
nand U3285 (N_3285,N_2980,N_2574);
and U3286 (N_3286,N_2268,N_2318);
nor U3287 (N_3287,N_2921,N_2468);
nand U3288 (N_3288,N_2213,N_2050);
nor U3289 (N_3289,N_2855,N_2183);
or U3290 (N_3290,N_2589,N_2946);
nor U3291 (N_3291,N_2217,N_2955);
nor U3292 (N_3292,N_2091,N_2031);
nand U3293 (N_3293,N_2952,N_2624);
nand U3294 (N_3294,N_2309,N_2058);
xnor U3295 (N_3295,N_2857,N_2508);
xor U3296 (N_3296,N_2456,N_2437);
and U3297 (N_3297,N_2836,N_2043);
nand U3298 (N_3298,N_2548,N_2842);
nor U3299 (N_3299,N_2748,N_2967);
or U3300 (N_3300,N_2922,N_2491);
nor U3301 (N_3301,N_2337,N_2747);
nand U3302 (N_3302,N_2903,N_2138);
or U3303 (N_3303,N_2993,N_2809);
and U3304 (N_3304,N_2593,N_2451);
xnor U3305 (N_3305,N_2803,N_2135);
xor U3306 (N_3306,N_2350,N_2144);
nor U3307 (N_3307,N_2932,N_2176);
and U3308 (N_3308,N_2995,N_2785);
or U3309 (N_3309,N_2959,N_2774);
xnor U3310 (N_3310,N_2917,N_2236);
nor U3311 (N_3311,N_2668,N_2277);
and U3312 (N_3312,N_2865,N_2273);
xor U3313 (N_3313,N_2871,N_2896);
nand U3314 (N_3314,N_2241,N_2687);
nand U3315 (N_3315,N_2106,N_2719);
nand U3316 (N_3316,N_2936,N_2391);
xor U3317 (N_3317,N_2622,N_2682);
nand U3318 (N_3318,N_2052,N_2874);
or U3319 (N_3319,N_2811,N_2288);
nand U3320 (N_3320,N_2695,N_2219);
nand U3321 (N_3321,N_2035,N_2760);
nor U3322 (N_3322,N_2286,N_2472);
or U3323 (N_3323,N_2190,N_2915);
nand U3324 (N_3324,N_2492,N_2481);
xor U3325 (N_3325,N_2279,N_2799);
nand U3326 (N_3326,N_2833,N_2753);
xor U3327 (N_3327,N_2187,N_2561);
nand U3328 (N_3328,N_2651,N_2998);
xor U3329 (N_3329,N_2497,N_2095);
xnor U3330 (N_3330,N_2720,N_2742);
and U3331 (N_3331,N_2255,N_2689);
xnor U3332 (N_3332,N_2966,N_2672);
nand U3333 (N_3333,N_2047,N_2569);
nand U3334 (N_3334,N_2390,N_2179);
nand U3335 (N_3335,N_2224,N_2021);
xor U3336 (N_3336,N_2637,N_2505);
or U3337 (N_3337,N_2576,N_2038);
xor U3338 (N_3338,N_2537,N_2981);
nor U3339 (N_3339,N_2100,N_2612);
xnor U3340 (N_3340,N_2207,N_2616);
nor U3341 (N_3341,N_2822,N_2248);
and U3342 (N_3342,N_2868,N_2229);
xor U3343 (N_3343,N_2802,N_2435);
nand U3344 (N_3344,N_2891,N_2916);
nor U3345 (N_3345,N_2408,N_2404);
or U3346 (N_3346,N_2827,N_2406);
nor U3347 (N_3347,N_2425,N_2738);
nor U3348 (N_3348,N_2132,N_2467);
nand U3349 (N_3349,N_2221,N_2950);
and U3350 (N_3350,N_2887,N_2399);
nand U3351 (N_3351,N_2685,N_2123);
xor U3352 (N_3352,N_2030,N_2192);
nand U3353 (N_3353,N_2256,N_2706);
or U3354 (N_3354,N_2298,N_2832);
nor U3355 (N_3355,N_2275,N_2167);
or U3356 (N_3356,N_2495,N_2643);
nand U3357 (N_3357,N_2450,N_2086);
or U3358 (N_3358,N_2908,N_2523);
xnor U3359 (N_3359,N_2397,N_2092);
nand U3360 (N_3360,N_2620,N_2374);
xnor U3361 (N_3361,N_2259,N_2960);
nand U3362 (N_3362,N_2864,N_2458);
and U3363 (N_3363,N_2935,N_2185);
nor U3364 (N_3364,N_2880,N_2449);
and U3365 (N_3365,N_2354,N_2500);
nand U3366 (N_3366,N_2765,N_2510);
or U3367 (N_3367,N_2296,N_2246);
nand U3368 (N_3368,N_2367,N_2545);
nor U3369 (N_3369,N_2159,N_2886);
nand U3370 (N_3370,N_2586,N_2371);
and U3371 (N_3371,N_2054,N_2919);
and U3372 (N_3372,N_2920,N_2796);
or U3373 (N_3373,N_2070,N_2639);
nor U3374 (N_3374,N_2324,N_2978);
nand U3375 (N_3375,N_2931,N_2501);
nand U3376 (N_3376,N_2701,N_2200);
nand U3377 (N_3377,N_2120,N_2168);
nor U3378 (N_3378,N_2262,N_2531);
nor U3379 (N_3379,N_2722,N_2478);
nor U3380 (N_3380,N_2424,N_2839);
xnor U3381 (N_3381,N_2819,N_2627);
xnor U3382 (N_3382,N_2085,N_2339);
nor U3383 (N_3383,N_2049,N_2948);
and U3384 (N_3384,N_2457,N_2169);
nand U3385 (N_3385,N_2515,N_2843);
or U3386 (N_3386,N_2970,N_2161);
and U3387 (N_3387,N_2654,N_2012);
xnor U3388 (N_3388,N_2145,N_2266);
xnor U3389 (N_3389,N_2585,N_2696);
or U3390 (N_3390,N_2770,N_2681);
xnor U3391 (N_3391,N_2509,N_2579);
or U3392 (N_3392,N_2873,N_2416);
or U3393 (N_3393,N_2314,N_2834);
and U3394 (N_3394,N_2336,N_2555);
xnor U3395 (N_3395,N_2455,N_2533);
xnor U3396 (N_3396,N_2292,N_2828);
and U3397 (N_3397,N_2413,N_2741);
nand U3398 (N_3398,N_2445,N_2494);
and U3399 (N_3399,N_2705,N_2094);
xnor U3400 (N_3400,N_2506,N_2443);
nor U3401 (N_3401,N_2729,N_2655);
nand U3402 (N_3402,N_2985,N_2804);
nor U3403 (N_3403,N_2067,N_2182);
nand U3404 (N_3404,N_2439,N_2153);
nand U3405 (N_3405,N_2134,N_2634);
or U3406 (N_3406,N_2013,N_2474);
nor U3407 (N_3407,N_2716,N_2238);
nand U3408 (N_3408,N_2805,N_2118);
or U3409 (N_3409,N_2075,N_2222);
and U3410 (N_3410,N_2566,N_2546);
nand U3411 (N_3411,N_2844,N_2347);
xnor U3412 (N_3412,N_2940,N_2194);
xnor U3413 (N_3413,N_2039,N_2535);
and U3414 (N_3414,N_2077,N_2723);
and U3415 (N_3415,N_2340,N_2674);
nand U3416 (N_3416,N_2825,N_2568);
and U3417 (N_3417,N_2104,N_2243);
nor U3418 (N_3418,N_2310,N_2272);
nor U3419 (N_3419,N_2164,N_2415);
and U3420 (N_3420,N_2215,N_2889);
xnor U3421 (N_3421,N_2108,N_2902);
nor U3422 (N_3422,N_2208,N_2590);
nor U3423 (N_3423,N_2677,N_2430);
xor U3424 (N_3424,N_2675,N_2551);
xor U3425 (N_3425,N_2400,N_2699);
nand U3426 (N_3426,N_2567,N_2821);
nand U3427 (N_3427,N_2364,N_2933);
nand U3428 (N_3428,N_2939,N_2688);
or U3429 (N_3429,N_2110,N_2003);
xor U3430 (N_3430,N_2470,N_2578);
and U3431 (N_3431,N_2170,N_2109);
nor U3432 (N_3432,N_2177,N_2897);
nand U3433 (N_3433,N_2020,N_2623);
nor U3434 (N_3434,N_2352,N_2368);
nand U3435 (N_3435,N_2409,N_2883);
and U3436 (N_3436,N_2511,N_2816);
xor U3437 (N_3437,N_2986,N_2547);
nand U3438 (N_3438,N_2125,N_2223);
and U3439 (N_3439,N_2002,N_2061);
nor U3440 (N_3440,N_2817,N_2918);
nor U3441 (N_3441,N_2403,N_2484);
xnor U3442 (N_3442,N_2411,N_2081);
and U3443 (N_3443,N_2244,N_2518);
xnor U3444 (N_3444,N_2759,N_2607);
nand U3445 (N_3445,N_2214,N_2636);
and U3446 (N_3446,N_2541,N_2293);
nand U3447 (N_3447,N_2342,N_2859);
and U3448 (N_3448,N_2284,N_2186);
nor U3449 (N_3449,N_2378,N_2365);
or U3450 (N_3450,N_2007,N_2536);
nor U3451 (N_3451,N_2088,N_2305);
xnor U3452 (N_3452,N_2402,N_2199);
xnor U3453 (N_3453,N_2376,N_2806);
and U3454 (N_3454,N_2673,N_2154);
and U3455 (N_3455,N_2252,N_2971);
and U3456 (N_3456,N_2389,N_2044);
xnor U3457 (N_3457,N_2851,N_2143);
or U3458 (N_3458,N_2388,N_2912);
xnor U3459 (N_3459,N_2861,N_2191);
nor U3460 (N_3460,N_2680,N_2487);
or U3461 (N_3461,N_2601,N_2786);
xnor U3462 (N_3462,N_2128,N_2041);
or U3463 (N_3463,N_2333,N_2755);
xnor U3464 (N_3464,N_2904,N_2036);
and U3465 (N_3465,N_2984,N_2189);
or U3466 (N_3466,N_2652,N_2133);
and U3467 (N_3467,N_2136,N_2726);
nor U3468 (N_3468,N_2232,N_2270);
nand U3469 (N_3469,N_2625,N_2592);
xor U3470 (N_3470,N_2345,N_2130);
and U3471 (N_3471,N_2231,N_2062);
or U3472 (N_3472,N_2907,N_2717);
xnor U3473 (N_3473,N_2226,N_2384);
nand U3474 (N_3474,N_2488,N_2994);
and U3475 (N_3475,N_2661,N_2982);
or U3476 (N_3476,N_2126,N_2557);
and U3477 (N_3477,N_2746,N_2769);
xnor U3478 (N_3478,N_2961,N_2080);
nand U3479 (N_3479,N_2299,N_2860);
xnor U3480 (N_3480,N_2358,N_2740);
nand U3481 (N_3481,N_2573,N_2888);
nand U3482 (N_3482,N_2431,N_2099);
nor U3483 (N_3483,N_2676,N_2327);
or U3484 (N_3484,N_2944,N_2028);
nand U3485 (N_3485,N_2023,N_2398);
nor U3486 (N_3486,N_2466,N_2131);
and U3487 (N_3487,N_2429,N_2815);
nor U3488 (N_3488,N_2254,N_2355);
nor U3489 (N_3489,N_2253,N_2733);
nor U3490 (N_3490,N_2294,N_2999);
or U3491 (N_3491,N_2577,N_2119);
nand U3492 (N_3492,N_2650,N_2107);
nand U3493 (N_3493,N_2987,N_2407);
and U3494 (N_3494,N_2444,N_2977);
xnor U3495 (N_3495,N_2372,N_2037);
nand U3496 (N_3496,N_2332,N_2172);
nor U3497 (N_3497,N_2911,N_2958);
nand U3498 (N_3498,N_2375,N_2715);
nor U3499 (N_3499,N_2771,N_2074);
xnor U3500 (N_3500,N_2791,N_2083);
and U3501 (N_3501,N_2302,N_2675);
nand U3502 (N_3502,N_2964,N_2436);
nor U3503 (N_3503,N_2878,N_2017);
nand U3504 (N_3504,N_2302,N_2284);
nor U3505 (N_3505,N_2469,N_2747);
nand U3506 (N_3506,N_2537,N_2041);
and U3507 (N_3507,N_2664,N_2822);
nand U3508 (N_3508,N_2854,N_2297);
nor U3509 (N_3509,N_2956,N_2950);
xnor U3510 (N_3510,N_2728,N_2944);
xor U3511 (N_3511,N_2472,N_2372);
nand U3512 (N_3512,N_2126,N_2259);
nand U3513 (N_3513,N_2788,N_2002);
or U3514 (N_3514,N_2995,N_2129);
and U3515 (N_3515,N_2855,N_2070);
and U3516 (N_3516,N_2466,N_2615);
nand U3517 (N_3517,N_2689,N_2259);
and U3518 (N_3518,N_2093,N_2512);
nand U3519 (N_3519,N_2217,N_2672);
nand U3520 (N_3520,N_2034,N_2185);
and U3521 (N_3521,N_2948,N_2100);
xnor U3522 (N_3522,N_2210,N_2589);
nor U3523 (N_3523,N_2256,N_2879);
xor U3524 (N_3524,N_2205,N_2695);
xor U3525 (N_3525,N_2170,N_2600);
or U3526 (N_3526,N_2761,N_2190);
or U3527 (N_3527,N_2281,N_2488);
or U3528 (N_3528,N_2929,N_2522);
nor U3529 (N_3529,N_2924,N_2899);
nand U3530 (N_3530,N_2014,N_2887);
nor U3531 (N_3531,N_2754,N_2534);
xor U3532 (N_3532,N_2336,N_2859);
xnor U3533 (N_3533,N_2905,N_2019);
or U3534 (N_3534,N_2793,N_2903);
and U3535 (N_3535,N_2256,N_2057);
nor U3536 (N_3536,N_2884,N_2601);
xnor U3537 (N_3537,N_2403,N_2947);
and U3538 (N_3538,N_2186,N_2002);
xor U3539 (N_3539,N_2800,N_2725);
and U3540 (N_3540,N_2652,N_2756);
or U3541 (N_3541,N_2049,N_2582);
or U3542 (N_3542,N_2722,N_2867);
or U3543 (N_3543,N_2383,N_2269);
nor U3544 (N_3544,N_2250,N_2747);
and U3545 (N_3545,N_2877,N_2234);
and U3546 (N_3546,N_2481,N_2275);
nand U3547 (N_3547,N_2471,N_2743);
nor U3548 (N_3548,N_2506,N_2342);
nor U3549 (N_3549,N_2288,N_2465);
and U3550 (N_3550,N_2641,N_2665);
xor U3551 (N_3551,N_2466,N_2092);
and U3552 (N_3552,N_2109,N_2905);
nor U3553 (N_3553,N_2236,N_2576);
or U3554 (N_3554,N_2706,N_2330);
and U3555 (N_3555,N_2763,N_2213);
or U3556 (N_3556,N_2335,N_2652);
nor U3557 (N_3557,N_2697,N_2791);
and U3558 (N_3558,N_2335,N_2545);
or U3559 (N_3559,N_2181,N_2208);
nand U3560 (N_3560,N_2845,N_2089);
and U3561 (N_3561,N_2009,N_2983);
nor U3562 (N_3562,N_2308,N_2399);
xor U3563 (N_3563,N_2822,N_2486);
and U3564 (N_3564,N_2009,N_2743);
or U3565 (N_3565,N_2171,N_2647);
nand U3566 (N_3566,N_2890,N_2202);
nand U3567 (N_3567,N_2141,N_2681);
nor U3568 (N_3568,N_2225,N_2705);
xnor U3569 (N_3569,N_2652,N_2796);
nand U3570 (N_3570,N_2581,N_2731);
and U3571 (N_3571,N_2838,N_2293);
and U3572 (N_3572,N_2008,N_2017);
nor U3573 (N_3573,N_2565,N_2910);
nor U3574 (N_3574,N_2836,N_2624);
nand U3575 (N_3575,N_2621,N_2664);
xor U3576 (N_3576,N_2632,N_2354);
xor U3577 (N_3577,N_2342,N_2173);
nor U3578 (N_3578,N_2161,N_2006);
xor U3579 (N_3579,N_2676,N_2160);
and U3580 (N_3580,N_2586,N_2368);
nand U3581 (N_3581,N_2437,N_2240);
or U3582 (N_3582,N_2964,N_2272);
nand U3583 (N_3583,N_2571,N_2343);
or U3584 (N_3584,N_2223,N_2368);
and U3585 (N_3585,N_2806,N_2164);
nor U3586 (N_3586,N_2293,N_2859);
xnor U3587 (N_3587,N_2590,N_2213);
nor U3588 (N_3588,N_2211,N_2088);
or U3589 (N_3589,N_2974,N_2863);
or U3590 (N_3590,N_2491,N_2364);
xnor U3591 (N_3591,N_2463,N_2527);
or U3592 (N_3592,N_2325,N_2819);
or U3593 (N_3593,N_2515,N_2280);
and U3594 (N_3594,N_2493,N_2895);
nand U3595 (N_3595,N_2134,N_2589);
nand U3596 (N_3596,N_2533,N_2435);
nand U3597 (N_3597,N_2380,N_2143);
or U3598 (N_3598,N_2749,N_2622);
nor U3599 (N_3599,N_2617,N_2325);
nor U3600 (N_3600,N_2983,N_2116);
and U3601 (N_3601,N_2825,N_2424);
xor U3602 (N_3602,N_2560,N_2977);
nand U3603 (N_3603,N_2422,N_2590);
or U3604 (N_3604,N_2845,N_2651);
and U3605 (N_3605,N_2629,N_2583);
xnor U3606 (N_3606,N_2408,N_2202);
or U3607 (N_3607,N_2623,N_2395);
xnor U3608 (N_3608,N_2843,N_2045);
nand U3609 (N_3609,N_2355,N_2687);
nor U3610 (N_3610,N_2290,N_2919);
or U3611 (N_3611,N_2256,N_2315);
and U3612 (N_3612,N_2596,N_2868);
nor U3613 (N_3613,N_2917,N_2647);
nand U3614 (N_3614,N_2554,N_2530);
nor U3615 (N_3615,N_2196,N_2034);
xor U3616 (N_3616,N_2410,N_2731);
and U3617 (N_3617,N_2599,N_2263);
or U3618 (N_3618,N_2191,N_2366);
nor U3619 (N_3619,N_2818,N_2458);
or U3620 (N_3620,N_2604,N_2898);
or U3621 (N_3621,N_2341,N_2209);
nand U3622 (N_3622,N_2144,N_2573);
nand U3623 (N_3623,N_2972,N_2867);
nor U3624 (N_3624,N_2858,N_2786);
nor U3625 (N_3625,N_2348,N_2611);
nor U3626 (N_3626,N_2109,N_2804);
or U3627 (N_3627,N_2126,N_2286);
nand U3628 (N_3628,N_2617,N_2377);
nor U3629 (N_3629,N_2512,N_2128);
xnor U3630 (N_3630,N_2986,N_2612);
nand U3631 (N_3631,N_2149,N_2578);
nor U3632 (N_3632,N_2807,N_2859);
and U3633 (N_3633,N_2585,N_2667);
and U3634 (N_3634,N_2367,N_2028);
and U3635 (N_3635,N_2325,N_2584);
nand U3636 (N_3636,N_2394,N_2926);
xnor U3637 (N_3637,N_2291,N_2095);
xnor U3638 (N_3638,N_2925,N_2167);
or U3639 (N_3639,N_2469,N_2293);
nand U3640 (N_3640,N_2785,N_2197);
nand U3641 (N_3641,N_2097,N_2779);
xor U3642 (N_3642,N_2712,N_2972);
nand U3643 (N_3643,N_2641,N_2458);
xor U3644 (N_3644,N_2061,N_2858);
nand U3645 (N_3645,N_2012,N_2078);
or U3646 (N_3646,N_2372,N_2670);
or U3647 (N_3647,N_2531,N_2309);
nor U3648 (N_3648,N_2668,N_2820);
nor U3649 (N_3649,N_2999,N_2071);
nor U3650 (N_3650,N_2049,N_2795);
and U3651 (N_3651,N_2985,N_2599);
nand U3652 (N_3652,N_2680,N_2823);
nor U3653 (N_3653,N_2772,N_2294);
or U3654 (N_3654,N_2625,N_2944);
xor U3655 (N_3655,N_2795,N_2731);
nand U3656 (N_3656,N_2705,N_2440);
xnor U3657 (N_3657,N_2550,N_2288);
nand U3658 (N_3658,N_2074,N_2121);
and U3659 (N_3659,N_2386,N_2424);
xor U3660 (N_3660,N_2680,N_2887);
nand U3661 (N_3661,N_2607,N_2103);
xor U3662 (N_3662,N_2592,N_2087);
nand U3663 (N_3663,N_2695,N_2096);
nor U3664 (N_3664,N_2144,N_2375);
or U3665 (N_3665,N_2610,N_2892);
xor U3666 (N_3666,N_2077,N_2608);
xnor U3667 (N_3667,N_2725,N_2681);
nor U3668 (N_3668,N_2464,N_2568);
or U3669 (N_3669,N_2975,N_2728);
xor U3670 (N_3670,N_2869,N_2804);
nor U3671 (N_3671,N_2765,N_2598);
nand U3672 (N_3672,N_2307,N_2961);
and U3673 (N_3673,N_2664,N_2688);
and U3674 (N_3674,N_2723,N_2689);
nand U3675 (N_3675,N_2913,N_2628);
xor U3676 (N_3676,N_2999,N_2448);
and U3677 (N_3677,N_2887,N_2432);
or U3678 (N_3678,N_2368,N_2767);
and U3679 (N_3679,N_2396,N_2487);
nand U3680 (N_3680,N_2518,N_2530);
and U3681 (N_3681,N_2058,N_2908);
nand U3682 (N_3682,N_2463,N_2037);
nand U3683 (N_3683,N_2395,N_2946);
xor U3684 (N_3684,N_2728,N_2881);
xor U3685 (N_3685,N_2866,N_2533);
and U3686 (N_3686,N_2358,N_2460);
nor U3687 (N_3687,N_2135,N_2670);
nor U3688 (N_3688,N_2806,N_2191);
nand U3689 (N_3689,N_2096,N_2842);
or U3690 (N_3690,N_2193,N_2626);
nor U3691 (N_3691,N_2839,N_2317);
nor U3692 (N_3692,N_2550,N_2019);
xor U3693 (N_3693,N_2542,N_2432);
and U3694 (N_3694,N_2935,N_2751);
and U3695 (N_3695,N_2623,N_2996);
nand U3696 (N_3696,N_2402,N_2399);
xnor U3697 (N_3697,N_2353,N_2847);
xor U3698 (N_3698,N_2438,N_2273);
or U3699 (N_3699,N_2949,N_2381);
nand U3700 (N_3700,N_2941,N_2557);
nor U3701 (N_3701,N_2777,N_2017);
or U3702 (N_3702,N_2817,N_2504);
and U3703 (N_3703,N_2744,N_2572);
nand U3704 (N_3704,N_2620,N_2353);
nor U3705 (N_3705,N_2207,N_2092);
and U3706 (N_3706,N_2622,N_2891);
nor U3707 (N_3707,N_2321,N_2459);
and U3708 (N_3708,N_2839,N_2006);
and U3709 (N_3709,N_2674,N_2093);
xor U3710 (N_3710,N_2878,N_2148);
xor U3711 (N_3711,N_2376,N_2843);
and U3712 (N_3712,N_2362,N_2796);
and U3713 (N_3713,N_2268,N_2964);
xnor U3714 (N_3714,N_2954,N_2282);
nand U3715 (N_3715,N_2415,N_2834);
nor U3716 (N_3716,N_2744,N_2496);
or U3717 (N_3717,N_2364,N_2560);
or U3718 (N_3718,N_2164,N_2768);
or U3719 (N_3719,N_2934,N_2075);
and U3720 (N_3720,N_2618,N_2503);
nor U3721 (N_3721,N_2829,N_2838);
or U3722 (N_3722,N_2172,N_2490);
and U3723 (N_3723,N_2456,N_2716);
nand U3724 (N_3724,N_2757,N_2695);
or U3725 (N_3725,N_2610,N_2241);
nand U3726 (N_3726,N_2127,N_2467);
xor U3727 (N_3727,N_2993,N_2205);
xor U3728 (N_3728,N_2625,N_2363);
and U3729 (N_3729,N_2477,N_2484);
xor U3730 (N_3730,N_2353,N_2975);
nor U3731 (N_3731,N_2280,N_2802);
nor U3732 (N_3732,N_2690,N_2781);
nor U3733 (N_3733,N_2267,N_2946);
and U3734 (N_3734,N_2999,N_2200);
nor U3735 (N_3735,N_2696,N_2237);
nand U3736 (N_3736,N_2747,N_2779);
and U3737 (N_3737,N_2764,N_2669);
xnor U3738 (N_3738,N_2278,N_2827);
xor U3739 (N_3739,N_2897,N_2157);
and U3740 (N_3740,N_2642,N_2245);
nor U3741 (N_3741,N_2809,N_2863);
or U3742 (N_3742,N_2149,N_2785);
nand U3743 (N_3743,N_2052,N_2179);
xnor U3744 (N_3744,N_2251,N_2230);
or U3745 (N_3745,N_2332,N_2072);
or U3746 (N_3746,N_2760,N_2019);
nand U3747 (N_3747,N_2397,N_2306);
xnor U3748 (N_3748,N_2618,N_2967);
nand U3749 (N_3749,N_2463,N_2182);
or U3750 (N_3750,N_2506,N_2056);
and U3751 (N_3751,N_2495,N_2031);
and U3752 (N_3752,N_2302,N_2485);
and U3753 (N_3753,N_2368,N_2534);
nor U3754 (N_3754,N_2728,N_2865);
nand U3755 (N_3755,N_2369,N_2203);
xnor U3756 (N_3756,N_2603,N_2442);
nor U3757 (N_3757,N_2283,N_2859);
and U3758 (N_3758,N_2072,N_2194);
xnor U3759 (N_3759,N_2388,N_2358);
or U3760 (N_3760,N_2203,N_2950);
nor U3761 (N_3761,N_2879,N_2131);
nand U3762 (N_3762,N_2934,N_2229);
and U3763 (N_3763,N_2225,N_2540);
nand U3764 (N_3764,N_2226,N_2197);
xnor U3765 (N_3765,N_2871,N_2236);
nor U3766 (N_3766,N_2800,N_2449);
nor U3767 (N_3767,N_2361,N_2179);
or U3768 (N_3768,N_2912,N_2779);
xor U3769 (N_3769,N_2652,N_2892);
or U3770 (N_3770,N_2273,N_2455);
nand U3771 (N_3771,N_2091,N_2051);
or U3772 (N_3772,N_2184,N_2221);
and U3773 (N_3773,N_2700,N_2740);
and U3774 (N_3774,N_2652,N_2945);
nor U3775 (N_3775,N_2302,N_2940);
or U3776 (N_3776,N_2910,N_2277);
or U3777 (N_3777,N_2372,N_2874);
nor U3778 (N_3778,N_2946,N_2707);
nand U3779 (N_3779,N_2989,N_2345);
xor U3780 (N_3780,N_2512,N_2375);
xor U3781 (N_3781,N_2592,N_2010);
nor U3782 (N_3782,N_2100,N_2178);
and U3783 (N_3783,N_2710,N_2362);
nor U3784 (N_3784,N_2911,N_2345);
nor U3785 (N_3785,N_2724,N_2069);
nor U3786 (N_3786,N_2414,N_2686);
xor U3787 (N_3787,N_2221,N_2394);
nand U3788 (N_3788,N_2712,N_2287);
or U3789 (N_3789,N_2792,N_2316);
xnor U3790 (N_3790,N_2627,N_2007);
xnor U3791 (N_3791,N_2108,N_2882);
nor U3792 (N_3792,N_2566,N_2473);
nand U3793 (N_3793,N_2720,N_2689);
nor U3794 (N_3794,N_2091,N_2518);
nand U3795 (N_3795,N_2477,N_2974);
nor U3796 (N_3796,N_2310,N_2936);
and U3797 (N_3797,N_2284,N_2518);
or U3798 (N_3798,N_2065,N_2653);
or U3799 (N_3799,N_2557,N_2204);
nand U3800 (N_3800,N_2157,N_2222);
xor U3801 (N_3801,N_2235,N_2048);
or U3802 (N_3802,N_2944,N_2702);
and U3803 (N_3803,N_2580,N_2973);
nor U3804 (N_3804,N_2274,N_2267);
xnor U3805 (N_3805,N_2767,N_2825);
and U3806 (N_3806,N_2862,N_2271);
xnor U3807 (N_3807,N_2889,N_2185);
xnor U3808 (N_3808,N_2693,N_2627);
nor U3809 (N_3809,N_2102,N_2598);
or U3810 (N_3810,N_2592,N_2704);
or U3811 (N_3811,N_2489,N_2837);
and U3812 (N_3812,N_2337,N_2957);
and U3813 (N_3813,N_2791,N_2674);
and U3814 (N_3814,N_2156,N_2068);
nand U3815 (N_3815,N_2484,N_2616);
xor U3816 (N_3816,N_2678,N_2873);
nand U3817 (N_3817,N_2795,N_2086);
and U3818 (N_3818,N_2336,N_2471);
nand U3819 (N_3819,N_2681,N_2841);
nor U3820 (N_3820,N_2500,N_2192);
nor U3821 (N_3821,N_2136,N_2513);
nor U3822 (N_3822,N_2192,N_2989);
nand U3823 (N_3823,N_2213,N_2328);
nor U3824 (N_3824,N_2045,N_2071);
nand U3825 (N_3825,N_2488,N_2341);
nor U3826 (N_3826,N_2417,N_2948);
nand U3827 (N_3827,N_2954,N_2654);
nand U3828 (N_3828,N_2215,N_2673);
or U3829 (N_3829,N_2505,N_2063);
nand U3830 (N_3830,N_2638,N_2859);
or U3831 (N_3831,N_2347,N_2621);
and U3832 (N_3832,N_2681,N_2927);
or U3833 (N_3833,N_2025,N_2594);
or U3834 (N_3834,N_2458,N_2215);
xnor U3835 (N_3835,N_2077,N_2746);
and U3836 (N_3836,N_2065,N_2779);
nor U3837 (N_3837,N_2553,N_2576);
xnor U3838 (N_3838,N_2779,N_2791);
and U3839 (N_3839,N_2819,N_2137);
nand U3840 (N_3840,N_2110,N_2673);
nor U3841 (N_3841,N_2219,N_2870);
and U3842 (N_3842,N_2379,N_2953);
and U3843 (N_3843,N_2153,N_2829);
xor U3844 (N_3844,N_2285,N_2405);
xor U3845 (N_3845,N_2369,N_2911);
or U3846 (N_3846,N_2694,N_2612);
nor U3847 (N_3847,N_2224,N_2125);
nor U3848 (N_3848,N_2615,N_2745);
nor U3849 (N_3849,N_2648,N_2406);
xor U3850 (N_3850,N_2470,N_2949);
and U3851 (N_3851,N_2660,N_2606);
xor U3852 (N_3852,N_2056,N_2519);
nor U3853 (N_3853,N_2188,N_2823);
nor U3854 (N_3854,N_2430,N_2871);
or U3855 (N_3855,N_2349,N_2839);
and U3856 (N_3856,N_2261,N_2189);
or U3857 (N_3857,N_2792,N_2382);
nand U3858 (N_3858,N_2565,N_2389);
or U3859 (N_3859,N_2961,N_2411);
xnor U3860 (N_3860,N_2014,N_2080);
xor U3861 (N_3861,N_2398,N_2504);
nand U3862 (N_3862,N_2465,N_2400);
or U3863 (N_3863,N_2906,N_2017);
xnor U3864 (N_3864,N_2798,N_2718);
nand U3865 (N_3865,N_2779,N_2557);
nor U3866 (N_3866,N_2934,N_2041);
and U3867 (N_3867,N_2744,N_2023);
xor U3868 (N_3868,N_2474,N_2215);
or U3869 (N_3869,N_2858,N_2307);
nand U3870 (N_3870,N_2222,N_2345);
nor U3871 (N_3871,N_2246,N_2719);
nor U3872 (N_3872,N_2144,N_2295);
nand U3873 (N_3873,N_2760,N_2259);
nand U3874 (N_3874,N_2785,N_2033);
or U3875 (N_3875,N_2323,N_2848);
xor U3876 (N_3876,N_2416,N_2367);
or U3877 (N_3877,N_2772,N_2565);
nand U3878 (N_3878,N_2102,N_2322);
nand U3879 (N_3879,N_2971,N_2284);
and U3880 (N_3880,N_2669,N_2078);
nand U3881 (N_3881,N_2122,N_2962);
xnor U3882 (N_3882,N_2581,N_2371);
and U3883 (N_3883,N_2037,N_2170);
or U3884 (N_3884,N_2959,N_2255);
xnor U3885 (N_3885,N_2379,N_2178);
and U3886 (N_3886,N_2642,N_2964);
nand U3887 (N_3887,N_2181,N_2901);
nand U3888 (N_3888,N_2857,N_2585);
and U3889 (N_3889,N_2665,N_2937);
or U3890 (N_3890,N_2035,N_2238);
or U3891 (N_3891,N_2851,N_2433);
nor U3892 (N_3892,N_2100,N_2412);
nand U3893 (N_3893,N_2948,N_2515);
and U3894 (N_3894,N_2312,N_2940);
or U3895 (N_3895,N_2065,N_2777);
nor U3896 (N_3896,N_2331,N_2241);
or U3897 (N_3897,N_2500,N_2061);
and U3898 (N_3898,N_2372,N_2739);
and U3899 (N_3899,N_2444,N_2338);
or U3900 (N_3900,N_2013,N_2677);
xnor U3901 (N_3901,N_2514,N_2218);
nor U3902 (N_3902,N_2592,N_2705);
nand U3903 (N_3903,N_2673,N_2775);
xor U3904 (N_3904,N_2773,N_2715);
xor U3905 (N_3905,N_2711,N_2811);
or U3906 (N_3906,N_2054,N_2982);
nand U3907 (N_3907,N_2550,N_2491);
nand U3908 (N_3908,N_2280,N_2253);
nor U3909 (N_3909,N_2634,N_2145);
nand U3910 (N_3910,N_2130,N_2069);
xnor U3911 (N_3911,N_2607,N_2018);
xor U3912 (N_3912,N_2162,N_2283);
xnor U3913 (N_3913,N_2174,N_2292);
nor U3914 (N_3914,N_2881,N_2776);
nand U3915 (N_3915,N_2230,N_2557);
or U3916 (N_3916,N_2845,N_2226);
nor U3917 (N_3917,N_2591,N_2633);
or U3918 (N_3918,N_2114,N_2107);
and U3919 (N_3919,N_2078,N_2549);
and U3920 (N_3920,N_2404,N_2546);
or U3921 (N_3921,N_2340,N_2513);
and U3922 (N_3922,N_2805,N_2995);
or U3923 (N_3923,N_2064,N_2591);
nor U3924 (N_3924,N_2427,N_2428);
nor U3925 (N_3925,N_2868,N_2080);
nor U3926 (N_3926,N_2399,N_2114);
or U3927 (N_3927,N_2757,N_2487);
nor U3928 (N_3928,N_2020,N_2690);
nand U3929 (N_3929,N_2495,N_2110);
nand U3930 (N_3930,N_2781,N_2744);
and U3931 (N_3931,N_2592,N_2486);
nor U3932 (N_3932,N_2952,N_2071);
or U3933 (N_3933,N_2166,N_2658);
or U3934 (N_3934,N_2675,N_2501);
nor U3935 (N_3935,N_2011,N_2708);
and U3936 (N_3936,N_2837,N_2311);
xor U3937 (N_3937,N_2449,N_2465);
nand U3938 (N_3938,N_2020,N_2129);
xor U3939 (N_3939,N_2555,N_2804);
nand U3940 (N_3940,N_2890,N_2314);
nor U3941 (N_3941,N_2640,N_2436);
xor U3942 (N_3942,N_2298,N_2715);
and U3943 (N_3943,N_2715,N_2733);
or U3944 (N_3944,N_2120,N_2302);
or U3945 (N_3945,N_2322,N_2451);
nor U3946 (N_3946,N_2893,N_2231);
or U3947 (N_3947,N_2984,N_2750);
or U3948 (N_3948,N_2920,N_2668);
or U3949 (N_3949,N_2581,N_2132);
xnor U3950 (N_3950,N_2946,N_2086);
or U3951 (N_3951,N_2186,N_2115);
nand U3952 (N_3952,N_2893,N_2894);
nand U3953 (N_3953,N_2246,N_2465);
or U3954 (N_3954,N_2959,N_2743);
xnor U3955 (N_3955,N_2125,N_2495);
nand U3956 (N_3956,N_2770,N_2925);
nand U3957 (N_3957,N_2953,N_2197);
nand U3958 (N_3958,N_2937,N_2584);
or U3959 (N_3959,N_2140,N_2530);
xor U3960 (N_3960,N_2727,N_2722);
xor U3961 (N_3961,N_2080,N_2949);
nand U3962 (N_3962,N_2798,N_2848);
nor U3963 (N_3963,N_2267,N_2952);
nand U3964 (N_3964,N_2693,N_2849);
or U3965 (N_3965,N_2144,N_2164);
nand U3966 (N_3966,N_2203,N_2175);
and U3967 (N_3967,N_2210,N_2826);
nor U3968 (N_3968,N_2250,N_2009);
and U3969 (N_3969,N_2529,N_2438);
xnor U3970 (N_3970,N_2439,N_2203);
xnor U3971 (N_3971,N_2932,N_2615);
nor U3972 (N_3972,N_2593,N_2603);
xnor U3973 (N_3973,N_2043,N_2881);
xnor U3974 (N_3974,N_2662,N_2578);
and U3975 (N_3975,N_2847,N_2365);
and U3976 (N_3976,N_2656,N_2712);
and U3977 (N_3977,N_2314,N_2042);
or U3978 (N_3978,N_2920,N_2064);
xor U3979 (N_3979,N_2426,N_2778);
or U3980 (N_3980,N_2922,N_2403);
and U3981 (N_3981,N_2856,N_2930);
xnor U3982 (N_3982,N_2786,N_2092);
xnor U3983 (N_3983,N_2219,N_2109);
nand U3984 (N_3984,N_2983,N_2689);
xnor U3985 (N_3985,N_2949,N_2861);
nand U3986 (N_3986,N_2564,N_2873);
and U3987 (N_3987,N_2813,N_2388);
nand U3988 (N_3988,N_2582,N_2212);
nor U3989 (N_3989,N_2460,N_2668);
nand U3990 (N_3990,N_2546,N_2832);
nand U3991 (N_3991,N_2517,N_2309);
nand U3992 (N_3992,N_2738,N_2769);
and U3993 (N_3993,N_2060,N_2349);
nor U3994 (N_3994,N_2423,N_2883);
and U3995 (N_3995,N_2685,N_2112);
nand U3996 (N_3996,N_2731,N_2694);
nand U3997 (N_3997,N_2642,N_2547);
nand U3998 (N_3998,N_2142,N_2574);
or U3999 (N_3999,N_2312,N_2208);
or U4000 (N_4000,N_3922,N_3705);
or U4001 (N_4001,N_3386,N_3070);
and U4002 (N_4002,N_3385,N_3455);
nor U4003 (N_4003,N_3409,N_3194);
or U4004 (N_4004,N_3485,N_3394);
xor U4005 (N_4005,N_3104,N_3663);
and U4006 (N_4006,N_3546,N_3000);
nand U4007 (N_4007,N_3549,N_3665);
or U4008 (N_4008,N_3303,N_3220);
nor U4009 (N_4009,N_3206,N_3298);
nand U4010 (N_4010,N_3135,N_3519);
nand U4011 (N_4011,N_3933,N_3333);
nor U4012 (N_4012,N_3481,N_3741);
and U4013 (N_4013,N_3789,N_3670);
and U4014 (N_4014,N_3863,N_3696);
or U4015 (N_4015,N_3074,N_3141);
xnor U4016 (N_4016,N_3996,N_3138);
xor U4017 (N_4017,N_3974,N_3879);
nand U4018 (N_4018,N_3729,N_3860);
xnor U4019 (N_4019,N_3189,N_3157);
and U4020 (N_4020,N_3521,N_3427);
nand U4021 (N_4021,N_3545,N_3906);
nor U4022 (N_4022,N_3589,N_3039);
nand U4023 (N_4023,N_3660,N_3606);
nor U4024 (N_4024,N_3825,N_3739);
xor U4025 (N_4025,N_3105,N_3969);
xor U4026 (N_4026,N_3083,N_3833);
and U4027 (N_4027,N_3057,N_3384);
xnor U4028 (N_4028,N_3793,N_3668);
and U4029 (N_4029,N_3136,N_3732);
nand U4030 (N_4030,N_3012,N_3588);
and U4031 (N_4031,N_3006,N_3004);
or U4032 (N_4032,N_3803,N_3015);
and U4033 (N_4033,N_3197,N_3888);
and U4034 (N_4034,N_3475,N_3140);
nor U4035 (N_4035,N_3877,N_3401);
nor U4036 (N_4036,N_3112,N_3227);
nor U4037 (N_4037,N_3210,N_3581);
or U4038 (N_4038,N_3465,N_3760);
or U4039 (N_4039,N_3402,N_3518);
nand U4040 (N_4040,N_3076,N_3239);
and U4041 (N_4041,N_3734,N_3586);
nor U4042 (N_4042,N_3348,N_3535);
nor U4043 (N_4043,N_3516,N_3850);
or U4044 (N_4044,N_3139,N_3980);
or U4045 (N_4045,N_3576,N_3802);
or U4046 (N_4046,N_3332,N_3926);
and U4047 (N_4047,N_3615,N_3899);
and U4048 (N_4048,N_3867,N_3600);
xnor U4049 (N_4049,N_3150,N_3986);
and U4050 (N_4050,N_3875,N_3654);
or U4051 (N_4051,N_3495,N_3752);
or U4052 (N_4052,N_3810,N_3678);
nor U4053 (N_4053,N_3073,N_3154);
and U4054 (N_4054,N_3770,N_3274);
nor U4055 (N_4055,N_3471,N_3257);
nor U4056 (N_4056,N_3349,N_3417);
xor U4057 (N_4057,N_3859,N_3077);
or U4058 (N_4058,N_3450,N_3594);
or U4059 (N_4059,N_3451,N_3474);
or U4060 (N_4060,N_3331,N_3709);
and U4061 (N_4061,N_3469,N_3609);
nor U4062 (N_4062,N_3362,N_3746);
and U4063 (N_4063,N_3261,N_3292);
nor U4064 (N_4064,N_3021,N_3673);
or U4065 (N_4065,N_3484,N_3540);
xor U4066 (N_4066,N_3617,N_3132);
nor U4067 (N_4067,N_3737,N_3256);
or U4068 (N_4068,N_3264,N_3610);
xnor U4069 (N_4069,N_3997,N_3568);
xnor U4070 (N_4070,N_3873,N_3943);
and U4071 (N_4071,N_3932,N_3815);
nand U4072 (N_4072,N_3062,N_3965);
nand U4073 (N_4073,N_3477,N_3635);
nor U4074 (N_4074,N_3953,N_3740);
nor U4075 (N_4075,N_3082,N_3319);
or U4076 (N_4076,N_3107,N_3356);
xnor U4077 (N_4077,N_3499,N_3856);
nor U4078 (N_4078,N_3351,N_3822);
or U4079 (N_4079,N_3228,N_3501);
or U4080 (N_4080,N_3056,N_3109);
nand U4081 (N_4081,N_3857,N_3837);
nand U4082 (N_4082,N_3761,N_3149);
and U4083 (N_4083,N_3410,N_3466);
or U4084 (N_4084,N_3940,N_3018);
nor U4085 (N_4085,N_3942,N_3171);
and U4086 (N_4086,N_3643,N_3988);
xnor U4087 (N_4087,N_3065,N_3921);
xor U4088 (N_4088,N_3565,N_3037);
nor U4089 (N_4089,N_3676,N_3829);
nand U4090 (N_4090,N_3278,N_3975);
xnor U4091 (N_4091,N_3184,N_3438);
xnor U4092 (N_4092,N_3376,N_3086);
nand U4093 (N_4093,N_3551,N_3176);
or U4094 (N_4094,N_3767,N_3631);
and U4095 (N_4095,N_3914,N_3880);
and U4096 (N_4096,N_3005,N_3266);
nand U4097 (N_4097,N_3907,N_3453);
and U4098 (N_4098,N_3909,N_3207);
and U4099 (N_4099,N_3329,N_3145);
nor U4100 (N_4100,N_3142,N_3308);
or U4101 (N_4101,N_3075,N_3778);
and U4102 (N_4102,N_3839,N_3273);
and U4103 (N_4103,N_3851,N_3637);
xor U4104 (N_4104,N_3188,N_3026);
or U4105 (N_4105,N_3337,N_3447);
nand U4106 (N_4106,N_3350,N_3180);
and U4107 (N_4107,N_3702,N_3464);
xor U4108 (N_4108,N_3796,N_3869);
nand U4109 (N_4109,N_3569,N_3375);
or U4110 (N_4110,N_3153,N_3653);
nor U4111 (N_4111,N_3934,N_3232);
xor U4112 (N_4112,N_3299,N_3941);
and U4113 (N_4113,N_3088,N_3787);
xnor U4114 (N_4114,N_3068,N_3395);
xnor U4115 (N_4115,N_3945,N_3230);
nor U4116 (N_4116,N_3658,N_3539);
xor U4117 (N_4117,N_3397,N_3411);
xnor U4118 (N_4118,N_3698,N_3585);
nand U4119 (N_4119,N_3764,N_3215);
nor U4120 (N_4120,N_3182,N_3035);
nor U4121 (N_4121,N_3664,N_3960);
nor U4122 (N_4122,N_3775,N_3573);
or U4123 (N_4123,N_3727,N_3683);
xor U4124 (N_4124,N_3710,N_3510);
or U4125 (N_4125,N_3255,N_3725);
and U4126 (N_4126,N_3419,N_3728);
nor U4127 (N_4127,N_3458,N_3853);
or U4128 (N_4128,N_3025,N_3396);
nand U4129 (N_4129,N_3642,N_3842);
xnor U4130 (N_4130,N_3721,N_3054);
xnor U4131 (N_4131,N_3618,N_3029);
xnor U4132 (N_4132,N_3774,N_3849);
nor U4133 (N_4133,N_3201,N_3317);
and U4134 (N_4134,N_3315,N_3553);
nor U4135 (N_4135,N_3249,N_3406);
nand U4136 (N_4136,N_3523,N_3017);
nor U4137 (N_4137,N_3442,N_3806);
nor U4138 (N_4138,N_3126,N_3704);
xor U4139 (N_4139,N_3420,N_3488);
and U4140 (N_4140,N_3325,N_3982);
xnor U4141 (N_4141,N_3008,N_3958);
xnor U4142 (N_4142,N_3616,N_3038);
or U4143 (N_4143,N_3408,N_3911);
nor U4144 (N_4144,N_3354,N_3338);
xor U4145 (N_4145,N_3625,N_3099);
xnor U4146 (N_4146,N_3042,N_3280);
xor U4147 (N_4147,N_3509,N_3582);
nand U4148 (N_4148,N_3460,N_3003);
nand U4149 (N_4149,N_3199,N_3883);
xnor U4150 (N_4150,N_3454,N_3759);
or U4151 (N_4151,N_3555,N_3282);
xnor U4152 (N_4152,N_3393,N_3925);
xnor U4153 (N_4153,N_3707,N_3514);
or U4154 (N_4154,N_3213,N_3797);
xor U4155 (N_4155,N_3301,N_3445);
xnor U4156 (N_4156,N_3370,N_3684);
or U4157 (N_4157,N_3231,N_3889);
and U4158 (N_4158,N_3391,N_3459);
nor U4159 (N_4159,N_3659,N_3052);
nand U4160 (N_4160,N_3198,N_3685);
nand U4161 (N_4161,N_3884,N_3253);
nor U4162 (N_4162,N_3304,N_3924);
or U4163 (N_4163,N_3515,N_3529);
xnor U4164 (N_4164,N_3089,N_3367);
nor U4165 (N_4165,N_3712,N_3542);
nor U4166 (N_4166,N_3532,N_3520);
nor U4167 (N_4167,N_3238,N_3195);
nand U4168 (N_4168,N_3938,N_3972);
and U4169 (N_4169,N_3808,N_3049);
and U4170 (N_4170,N_3413,N_3738);
nor U4171 (N_4171,N_3998,N_3689);
or U4172 (N_4172,N_3841,N_3896);
nor U4173 (N_4173,N_3389,N_3601);
and U4174 (N_4174,N_3047,N_3269);
nand U4175 (N_4175,N_3840,N_3719);
nor U4176 (N_4176,N_3784,N_3493);
nor U4177 (N_4177,N_3577,N_3927);
or U4178 (N_4178,N_3602,N_3782);
nor U4179 (N_4179,N_3828,N_3224);
nor U4180 (N_4180,N_3591,N_3050);
nor U4181 (N_4181,N_3405,N_3826);
xnor U4182 (N_4182,N_3124,N_3805);
nand U4183 (N_4183,N_3548,N_3671);
xnor U4184 (N_4184,N_3064,N_3834);
nor U4185 (N_4185,N_3811,N_3010);
nand U4186 (N_4186,N_3644,N_3930);
or U4187 (N_4187,N_3779,N_3095);
or U4188 (N_4188,N_3800,N_3439);
nand U4189 (N_4189,N_3378,N_3868);
xor U4190 (N_4190,N_3700,N_3128);
nand U4191 (N_4191,N_3745,N_3587);
nor U4192 (N_4192,N_3844,N_3881);
nor U4193 (N_4193,N_3456,N_3984);
nor U4194 (N_4194,N_3248,N_3426);
or U4195 (N_4195,N_3750,N_3111);
or U4196 (N_4196,N_3123,N_3776);
nor U4197 (N_4197,N_3084,N_3715);
and U4198 (N_4198,N_3309,N_3757);
or U4199 (N_4199,N_3032,N_3030);
xor U4200 (N_4200,N_3165,N_3716);
and U4201 (N_4201,N_3612,N_3358);
nor U4202 (N_4202,N_3987,N_3870);
and U4203 (N_4203,N_3887,N_3125);
nand U4204 (N_4204,N_3843,N_3167);
nor U4205 (N_4205,N_3814,N_3148);
nor U4206 (N_4206,N_3432,N_3836);
or U4207 (N_4207,N_3913,N_3936);
or U4208 (N_4208,N_3033,N_3462);
xor U4209 (N_4209,N_3636,N_3619);
xnor U4210 (N_4210,N_3871,N_3178);
xnor U4211 (N_4211,N_3743,N_3392);
xor U4212 (N_4212,N_3687,N_3983);
and U4213 (N_4213,N_3046,N_3059);
nand U4214 (N_4214,N_3892,N_3311);
xor U4215 (N_4215,N_3119,N_3865);
nor U4216 (N_4216,N_3657,N_3202);
and U4217 (N_4217,N_3762,N_3809);
nor U4218 (N_4218,N_3517,N_3507);
and U4219 (N_4219,N_3819,N_3622);
xor U4220 (N_4220,N_3723,N_3316);
nor U4221 (N_4221,N_3430,N_3302);
xor U4222 (N_4222,N_3288,N_3058);
xnor U4223 (N_4223,N_3160,N_3724);
and U4224 (N_4224,N_3570,N_3788);
or U4225 (N_4225,N_3277,N_3259);
nor U4226 (N_4226,N_3832,N_3603);
nand U4227 (N_4227,N_3599,N_3749);
or U4228 (N_4228,N_3666,N_3371);
and U4229 (N_4229,N_3677,N_3106);
nor U4230 (N_4230,N_3152,N_3571);
xor U4231 (N_4231,N_3262,N_3024);
or U4232 (N_4232,N_3818,N_3265);
and U4233 (N_4233,N_3116,N_3071);
and U4234 (N_4234,N_3977,N_3090);
or U4235 (N_4235,N_3085,N_3744);
nand U4236 (N_4236,N_3798,N_3443);
or U4237 (N_4237,N_3342,N_3699);
xor U4238 (N_4238,N_3604,N_3956);
or U4239 (N_4239,N_3830,N_3374);
or U4240 (N_4240,N_3159,N_3009);
and U4241 (N_4241,N_3931,N_3363);
and U4242 (N_4242,N_3204,N_3639);
xor U4243 (N_4243,N_3632,N_3785);
and U4244 (N_4244,N_3929,N_3377);
xnor U4245 (N_4245,N_3640,N_3334);
nand U4246 (N_4246,N_3023,N_3667);
nand U4247 (N_4247,N_3034,N_3944);
nor U4248 (N_4248,N_3897,N_3433);
xor U4249 (N_4249,N_3366,N_3271);
xor U4250 (N_4250,N_3713,N_3578);
and U4251 (N_4251,N_3703,N_3381);
or U4252 (N_4252,N_3444,N_3326);
and U4253 (N_4253,N_3904,N_3966);
xor U4254 (N_4254,N_3669,N_3313);
nor U4255 (N_4255,N_3322,N_3827);
nand U4256 (N_4256,N_3686,N_3066);
nor U4257 (N_4257,N_3694,N_3891);
nand U4258 (N_4258,N_3177,N_3866);
or U4259 (N_4259,N_3359,N_3369);
xnor U4260 (N_4260,N_3649,N_3087);
nor U4261 (N_4261,N_3629,N_3218);
nand U4262 (N_4262,N_3478,N_3792);
or U4263 (N_4263,N_3043,N_3560);
or U4264 (N_4264,N_3211,N_3959);
and U4265 (N_4265,N_3848,N_3648);
nand U4266 (N_4266,N_3284,N_3838);
and U4267 (N_4267,N_3820,N_3613);
nand U4268 (N_4268,N_3550,N_3002);
and U4269 (N_4269,N_3735,N_3534);
nand U4270 (N_4270,N_3388,N_3324);
or U4271 (N_4271,N_3435,N_3108);
xor U4272 (N_4272,N_3981,N_3415);
nor U4273 (N_4273,N_3185,N_3258);
nand U4274 (N_4274,N_3855,N_3915);
nand U4275 (N_4275,N_3053,N_3060);
and U4276 (N_4276,N_3225,N_3561);
or U4277 (N_4277,N_3970,N_3607);
and U4278 (N_4278,N_3424,N_3028);
nor U4279 (N_4279,N_3656,N_3339);
nor U4280 (N_4280,N_3387,N_3200);
or U4281 (N_4281,N_3916,N_3268);
or U4282 (N_4282,N_3222,N_3276);
nor U4283 (N_4283,N_3252,N_3731);
xor U4284 (N_4284,N_3511,N_3494);
xnor U4285 (N_4285,N_3559,N_3063);
and U4286 (N_4286,N_3067,N_3237);
or U4287 (N_4287,N_3482,N_3080);
and U4288 (N_4288,N_3964,N_3022);
nand U4289 (N_4289,N_3726,N_3151);
and U4290 (N_4290,N_3158,N_3242);
and U4291 (N_4291,N_3163,N_3250);
or U4292 (N_4292,N_3722,N_3681);
nand U4293 (N_4293,N_3835,N_3496);
xor U4294 (N_4294,N_3908,N_3270);
nand U4295 (N_4295,N_3885,N_3720);
nor U4296 (N_4296,N_3245,N_3437);
or U4297 (N_4297,N_3596,N_3852);
and U4298 (N_4298,N_3372,N_3293);
xnor U4299 (N_4299,N_3212,N_3431);
nand U4300 (N_4300,N_3260,N_3628);
or U4301 (N_4301,N_3783,N_3679);
xnor U4302 (N_4302,N_3187,N_3414);
nor U4303 (N_4303,N_3620,N_3706);
or U4304 (N_4304,N_3320,N_3407);
nand U4305 (N_4305,N_3161,N_3147);
xor U4306 (N_4306,N_3630,N_3799);
nand U4307 (N_4307,N_3920,N_3463);
nor U4308 (N_4308,N_3113,N_3114);
and U4309 (N_4309,N_3364,N_3742);
nand U4310 (N_4310,N_3524,N_3020);
nor U4311 (N_4311,N_3680,N_3504);
or U4312 (N_4312,N_3917,N_3583);
and U4313 (N_4313,N_3991,N_3697);
or U4314 (N_4314,N_3072,N_3078);
nand U4315 (N_4315,N_3590,N_3263);
nand U4316 (N_4316,N_3564,N_3655);
nand U4317 (N_4317,N_3247,N_3747);
nand U4318 (N_4318,N_3169,N_3234);
and U4319 (N_4319,N_3291,N_3756);
nand U4320 (N_4320,N_3821,N_3491);
or U4321 (N_4321,N_3131,N_3283);
and U4322 (N_4322,N_3110,N_3963);
or U4323 (N_4323,N_3978,N_3428);
nand U4324 (N_4324,N_3209,N_3682);
xnor U4325 (N_4325,N_3876,N_3452);
and U4326 (N_4326,N_3556,N_3390);
nor U4327 (N_4327,N_3769,N_3097);
or U4328 (N_4328,N_3893,N_3748);
and U4329 (N_4329,N_3971,N_3117);
nand U4330 (N_4330,N_3214,N_3330);
or U4331 (N_4331,N_3016,N_3403);
nand U4332 (N_4332,N_3595,N_3134);
nand U4333 (N_4333,N_3882,N_3773);
or U4334 (N_4334,N_3638,N_3497);
nor U4335 (N_4335,N_3900,N_3382);
or U4336 (N_4336,N_3467,N_3305);
or U4337 (N_4337,N_3918,N_3421);
and U4338 (N_4338,N_3133,N_3624);
or U4339 (N_4339,N_3285,N_3845);
nor U4340 (N_4340,N_3634,N_3973);
nor U4341 (N_4341,N_3281,N_3777);
nor U4342 (N_4342,N_3203,N_3544);
nand U4343 (N_4343,N_3902,N_3300);
nand U4344 (N_4344,N_3120,N_3768);
xor U4345 (N_4345,N_3692,N_3208);
and U4346 (N_4346,N_3036,N_3353);
nand U4347 (N_4347,N_3254,N_3318);
and U4348 (N_4348,N_3878,N_3446);
nand U4349 (N_4349,N_3967,N_3340);
xor U4350 (N_4350,N_3217,N_3098);
or U4351 (N_4351,N_3480,N_3506);
or U4352 (N_4352,N_3192,N_3823);
xnor U4353 (N_4353,N_3781,N_3448);
xor U4354 (N_4354,N_3297,N_3347);
or U4355 (N_4355,N_3647,N_3306);
and U4356 (N_4356,N_3976,N_3874);
or U4357 (N_4357,N_3817,N_3235);
xnor U4358 (N_4358,N_3275,N_3766);
or U4359 (N_4359,N_3525,N_3733);
xor U4360 (N_4360,N_3379,N_3557);
and U4361 (N_4361,N_3041,N_3989);
or U4362 (N_4362,N_3804,N_3813);
nor U4363 (N_4363,N_3079,N_3627);
or U4364 (N_4364,N_3193,N_3864);
xnor U4365 (N_4365,N_3919,N_3013);
nand U4366 (N_4366,N_3674,N_3051);
nand U4367 (N_4367,N_3717,N_3190);
xor U4368 (N_4368,N_3541,N_3383);
xnor U4369 (N_4369,N_3341,N_3861);
or U4370 (N_4370,N_3957,N_3490);
xor U4371 (N_4371,N_3122,N_3816);
nor U4372 (N_4372,N_3572,N_3675);
nand U4373 (N_4373,N_3412,N_3693);
and U4374 (N_4374,N_3574,N_3999);
xnor U4375 (N_4375,N_3172,N_3538);
nand U4376 (N_4376,N_3910,N_3531);
and U4377 (N_4377,N_3711,N_3449);
nor U4378 (N_4378,N_3102,N_3343);
nand U4379 (N_4379,N_3310,N_3502);
and U4380 (N_4380,N_3240,N_3399);
nand U4381 (N_4381,N_3441,N_3854);
or U4382 (N_4382,N_3295,N_3708);
and U4383 (N_4383,N_3498,N_3547);
nand U4384 (N_4384,N_3751,N_3241);
xor U4385 (N_4385,N_3730,N_3527);
nor U4386 (N_4386,N_3626,N_3069);
nand U4387 (N_4387,N_3948,N_3672);
nand U4388 (N_4388,N_3791,N_3790);
or U4389 (N_4389,N_3352,N_3890);
nand U4390 (N_4390,N_3346,N_3552);
xnor U4391 (N_4391,N_3422,N_3166);
nand U4392 (N_4392,N_3380,N_3968);
or U4393 (N_4393,N_3164,N_3952);
nor U4394 (N_4394,N_3690,N_3307);
nand U4395 (N_4395,N_3226,N_3605);
xor U4396 (N_4396,N_3592,N_3831);
nand U4397 (N_4397,N_3758,N_3429);
nand U4398 (N_4398,N_3183,N_3650);
and U4399 (N_4399,N_3061,N_3287);
nand U4400 (N_4400,N_3505,N_3794);
nand U4401 (N_4401,N_3895,N_3144);
xnor U4402 (N_4402,N_3186,N_3526);
nor U4403 (N_4403,N_3905,N_3489);
nand U4404 (N_4404,N_3344,N_3321);
nand U4405 (N_4405,N_3898,N_3961);
and U4406 (N_4406,N_3652,N_3962);
nand U4407 (N_4407,N_3470,N_3537);
and U4408 (N_4408,N_3623,N_3236);
or U4409 (N_4409,N_3040,N_3862);
and U4410 (N_4410,N_3646,N_3812);
or U4411 (N_4411,N_3503,N_3995);
xnor U4412 (N_4412,N_3121,N_3229);
nand U4413 (N_4413,N_3558,N_3081);
and U4414 (N_4414,N_3162,N_3701);
and U4415 (N_4415,N_3404,N_3048);
or U4416 (N_4416,N_3223,N_3949);
or U4417 (N_4417,N_3328,N_3714);
or U4418 (N_4418,N_3175,N_3912);
nand U4419 (N_4419,N_3323,N_3267);
nand U4420 (N_4420,N_3279,N_3174);
xor U4421 (N_4421,N_3368,N_3947);
nand U4422 (N_4422,N_3566,N_3513);
nand U4423 (N_4423,N_3651,N_3027);
and U4424 (N_4424,N_3345,N_3314);
nand U4425 (N_4425,N_3951,N_3901);
or U4426 (N_4426,N_3221,N_3508);
xor U4427 (N_4427,N_3954,N_3327);
xor U4428 (N_4428,N_3562,N_3473);
xor U4429 (N_4429,N_3872,N_3423);
xor U4430 (N_4430,N_3436,N_3661);
or U4431 (N_4431,N_3094,N_3718);
nand U4432 (N_4432,N_3251,N_3894);
nand U4433 (N_4433,N_3858,N_3786);
nand U4434 (N_4434,N_3014,N_3824);
nor U4435 (N_4435,N_3492,N_3522);
nor U4436 (N_4436,N_3479,N_3695);
and U4437 (N_4437,N_3091,N_3554);
xor U4438 (N_4438,N_3688,N_3156);
xor U4439 (N_4439,N_3979,N_3641);
nor U4440 (N_4440,N_3755,N_3290);
nand U4441 (N_4441,N_3946,N_3373);
and U4442 (N_4442,N_3584,N_3416);
xnor U4443 (N_4443,N_3533,N_3168);
nand U4444 (N_4444,N_3939,N_3272);
xnor U4445 (N_4445,N_3146,N_3512);
or U4446 (N_4446,N_3611,N_3530);
nor U4447 (N_4447,N_3101,N_3130);
and U4448 (N_4448,N_3486,N_3886);
nand U4449 (N_4449,N_3476,N_3001);
or U4450 (N_4450,N_3468,N_3801);
and U4451 (N_4451,N_3289,N_3336);
nand U4452 (N_4452,N_3312,N_3461);
xnor U4453 (N_4453,N_3127,N_3137);
or U4454 (N_4454,N_3246,N_3662);
xor U4455 (N_4455,N_3847,N_3903);
and U4456 (N_4456,N_3045,N_3621);
nor U4457 (N_4457,N_3418,N_3181);
nor U4458 (N_4458,N_3179,N_3771);
nand U4459 (N_4459,N_3115,N_3994);
nor U4460 (N_4460,N_3093,N_3092);
nand U4461 (N_4461,N_3440,N_3244);
or U4462 (N_4462,N_3807,N_3219);
or U4463 (N_4463,N_3103,N_3923);
nand U4464 (N_4464,N_3335,N_3575);
and U4465 (N_4465,N_3955,N_3780);
nand U4466 (N_4466,N_3011,N_3129);
or U4467 (N_4467,N_3935,N_3173);
xor U4468 (N_4468,N_3763,N_3563);
nand U4469 (N_4469,N_3096,N_3753);
or U4470 (N_4470,N_3155,N_3434);
nor U4471 (N_4471,N_3360,N_3355);
xor U4472 (N_4472,N_3736,N_3992);
nor U4473 (N_4473,N_3993,N_3500);
nand U4474 (N_4474,N_3216,N_3598);
or U4475 (N_4475,N_3985,N_3143);
xor U4476 (N_4476,N_3170,N_3286);
nand U4477 (N_4477,N_3191,N_3365);
nor U4478 (N_4478,N_3007,N_3044);
or U4479 (N_4479,N_3400,N_3928);
nor U4480 (N_4480,N_3100,N_3633);
or U4481 (N_4481,N_3597,N_3567);
nand U4482 (N_4482,N_3205,N_3196);
xnor U4483 (N_4483,N_3608,N_3055);
and U4484 (N_4484,N_3937,N_3528);
nor U4485 (N_4485,N_3457,N_3243);
nand U4486 (N_4486,N_3579,N_3614);
xor U4487 (N_4487,N_3019,N_3483);
xor U4488 (N_4488,N_3846,N_3691);
xor U4489 (N_4489,N_3772,N_3950);
or U4490 (N_4490,N_3357,N_3487);
xnor U4491 (N_4491,N_3536,N_3425);
nor U4492 (N_4492,N_3754,N_3118);
xnor U4493 (N_4493,N_3031,N_3472);
or U4494 (N_4494,N_3593,N_3296);
nand U4495 (N_4495,N_3233,N_3398);
or U4496 (N_4496,N_3580,N_3765);
and U4497 (N_4497,N_3645,N_3990);
nand U4498 (N_4498,N_3795,N_3361);
and U4499 (N_4499,N_3543,N_3294);
or U4500 (N_4500,N_3461,N_3128);
nand U4501 (N_4501,N_3453,N_3430);
and U4502 (N_4502,N_3214,N_3419);
and U4503 (N_4503,N_3959,N_3406);
xor U4504 (N_4504,N_3679,N_3949);
or U4505 (N_4505,N_3977,N_3900);
and U4506 (N_4506,N_3268,N_3034);
or U4507 (N_4507,N_3690,N_3167);
xnor U4508 (N_4508,N_3694,N_3426);
nor U4509 (N_4509,N_3922,N_3338);
xnor U4510 (N_4510,N_3973,N_3615);
nor U4511 (N_4511,N_3340,N_3565);
nand U4512 (N_4512,N_3635,N_3915);
xor U4513 (N_4513,N_3115,N_3516);
and U4514 (N_4514,N_3025,N_3991);
or U4515 (N_4515,N_3804,N_3997);
nor U4516 (N_4516,N_3927,N_3965);
nor U4517 (N_4517,N_3353,N_3092);
and U4518 (N_4518,N_3157,N_3834);
nor U4519 (N_4519,N_3014,N_3462);
nor U4520 (N_4520,N_3330,N_3898);
and U4521 (N_4521,N_3489,N_3148);
nand U4522 (N_4522,N_3554,N_3302);
nand U4523 (N_4523,N_3612,N_3083);
or U4524 (N_4524,N_3990,N_3704);
or U4525 (N_4525,N_3306,N_3303);
xnor U4526 (N_4526,N_3893,N_3328);
nand U4527 (N_4527,N_3868,N_3311);
xnor U4528 (N_4528,N_3080,N_3459);
or U4529 (N_4529,N_3443,N_3210);
or U4530 (N_4530,N_3231,N_3477);
xnor U4531 (N_4531,N_3309,N_3410);
nor U4532 (N_4532,N_3152,N_3844);
xnor U4533 (N_4533,N_3064,N_3234);
xnor U4534 (N_4534,N_3692,N_3184);
nor U4535 (N_4535,N_3852,N_3964);
or U4536 (N_4536,N_3677,N_3119);
and U4537 (N_4537,N_3810,N_3987);
nand U4538 (N_4538,N_3630,N_3355);
and U4539 (N_4539,N_3520,N_3892);
and U4540 (N_4540,N_3349,N_3763);
nor U4541 (N_4541,N_3706,N_3747);
xor U4542 (N_4542,N_3352,N_3784);
xor U4543 (N_4543,N_3123,N_3231);
and U4544 (N_4544,N_3180,N_3951);
nor U4545 (N_4545,N_3627,N_3896);
and U4546 (N_4546,N_3859,N_3403);
nand U4547 (N_4547,N_3494,N_3430);
xor U4548 (N_4548,N_3423,N_3755);
and U4549 (N_4549,N_3496,N_3269);
and U4550 (N_4550,N_3828,N_3963);
and U4551 (N_4551,N_3607,N_3126);
nor U4552 (N_4552,N_3285,N_3943);
nand U4553 (N_4553,N_3055,N_3056);
or U4554 (N_4554,N_3195,N_3525);
nand U4555 (N_4555,N_3488,N_3280);
nor U4556 (N_4556,N_3637,N_3998);
xnor U4557 (N_4557,N_3841,N_3706);
nor U4558 (N_4558,N_3892,N_3809);
nand U4559 (N_4559,N_3382,N_3605);
nor U4560 (N_4560,N_3914,N_3320);
or U4561 (N_4561,N_3728,N_3730);
or U4562 (N_4562,N_3418,N_3363);
nor U4563 (N_4563,N_3849,N_3860);
and U4564 (N_4564,N_3213,N_3809);
xnor U4565 (N_4565,N_3187,N_3397);
and U4566 (N_4566,N_3374,N_3224);
and U4567 (N_4567,N_3548,N_3164);
and U4568 (N_4568,N_3033,N_3536);
nand U4569 (N_4569,N_3983,N_3042);
xnor U4570 (N_4570,N_3032,N_3519);
and U4571 (N_4571,N_3415,N_3949);
and U4572 (N_4572,N_3669,N_3117);
nor U4573 (N_4573,N_3113,N_3442);
nand U4574 (N_4574,N_3210,N_3674);
nand U4575 (N_4575,N_3005,N_3172);
nor U4576 (N_4576,N_3555,N_3700);
nand U4577 (N_4577,N_3469,N_3321);
and U4578 (N_4578,N_3659,N_3129);
nor U4579 (N_4579,N_3166,N_3244);
nand U4580 (N_4580,N_3814,N_3908);
and U4581 (N_4581,N_3576,N_3463);
and U4582 (N_4582,N_3525,N_3565);
and U4583 (N_4583,N_3597,N_3454);
nand U4584 (N_4584,N_3826,N_3047);
or U4585 (N_4585,N_3041,N_3405);
and U4586 (N_4586,N_3564,N_3263);
nand U4587 (N_4587,N_3607,N_3804);
xnor U4588 (N_4588,N_3264,N_3630);
and U4589 (N_4589,N_3396,N_3732);
nor U4590 (N_4590,N_3011,N_3853);
or U4591 (N_4591,N_3978,N_3858);
nor U4592 (N_4592,N_3829,N_3159);
nor U4593 (N_4593,N_3948,N_3677);
nor U4594 (N_4594,N_3830,N_3725);
and U4595 (N_4595,N_3978,N_3713);
and U4596 (N_4596,N_3403,N_3219);
or U4597 (N_4597,N_3447,N_3456);
nor U4598 (N_4598,N_3865,N_3355);
or U4599 (N_4599,N_3033,N_3655);
and U4600 (N_4600,N_3221,N_3387);
nand U4601 (N_4601,N_3279,N_3993);
xor U4602 (N_4602,N_3619,N_3094);
nand U4603 (N_4603,N_3551,N_3466);
nor U4604 (N_4604,N_3405,N_3228);
nand U4605 (N_4605,N_3737,N_3513);
and U4606 (N_4606,N_3940,N_3200);
xor U4607 (N_4607,N_3838,N_3672);
or U4608 (N_4608,N_3178,N_3530);
or U4609 (N_4609,N_3460,N_3312);
and U4610 (N_4610,N_3898,N_3806);
xnor U4611 (N_4611,N_3982,N_3848);
or U4612 (N_4612,N_3572,N_3583);
xnor U4613 (N_4613,N_3856,N_3918);
or U4614 (N_4614,N_3554,N_3060);
nor U4615 (N_4615,N_3868,N_3184);
or U4616 (N_4616,N_3025,N_3833);
xor U4617 (N_4617,N_3713,N_3624);
xor U4618 (N_4618,N_3984,N_3471);
and U4619 (N_4619,N_3186,N_3930);
and U4620 (N_4620,N_3954,N_3541);
nor U4621 (N_4621,N_3802,N_3156);
nand U4622 (N_4622,N_3432,N_3916);
nor U4623 (N_4623,N_3384,N_3358);
xor U4624 (N_4624,N_3348,N_3358);
xor U4625 (N_4625,N_3675,N_3235);
or U4626 (N_4626,N_3296,N_3747);
nand U4627 (N_4627,N_3102,N_3553);
xor U4628 (N_4628,N_3803,N_3383);
or U4629 (N_4629,N_3232,N_3062);
and U4630 (N_4630,N_3060,N_3551);
nand U4631 (N_4631,N_3194,N_3101);
nand U4632 (N_4632,N_3466,N_3335);
xor U4633 (N_4633,N_3638,N_3287);
xor U4634 (N_4634,N_3783,N_3411);
nand U4635 (N_4635,N_3011,N_3441);
nand U4636 (N_4636,N_3186,N_3672);
xor U4637 (N_4637,N_3472,N_3358);
xnor U4638 (N_4638,N_3534,N_3020);
and U4639 (N_4639,N_3837,N_3372);
nand U4640 (N_4640,N_3347,N_3365);
nand U4641 (N_4641,N_3994,N_3716);
or U4642 (N_4642,N_3384,N_3399);
and U4643 (N_4643,N_3519,N_3601);
and U4644 (N_4644,N_3518,N_3882);
nand U4645 (N_4645,N_3585,N_3792);
xor U4646 (N_4646,N_3044,N_3022);
xor U4647 (N_4647,N_3808,N_3688);
xor U4648 (N_4648,N_3007,N_3812);
nor U4649 (N_4649,N_3250,N_3159);
and U4650 (N_4650,N_3335,N_3817);
and U4651 (N_4651,N_3202,N_3675);
xnor U4652 (N_4652,N_3146,N_3844);
nor U4653 (N_4653,N_3832,N_3367);
nor U4654 (N_4654,N_3535,N_3181);
nand U4655 (N_4655,N_3012,N_3060);
nand U4656 (N_4656,N_3086,N_3939);
xnor U4657 (N_4657,N_3839,N_3237);
and U4658 (N_4658,N_3434,N_3248);
or U4659 (N_4659,N_3833,N_3436);
nand U4660 (N_4660,N_3777,N_3741);
nand U4661 (N_4661,N_3205,N_3477);
and U4662 (N_4662,N_3396,N_3904);
and U4663 (N_4663,N_3542,N_3870);
or U4664 (N_4664,N_3845,N_3078);
and U4665 (N_4665,N_3821,N_3199);
nor U4666 (N_4666,N_3773,N_3299);
or U4667 (N_4667,N_3585,N_3290);
nor U4668 (N_4668,N_3528,N_3344);
nor U4669 (N_4669,N_3748,N_3333);
and U4670 (N_4670,N_3917,N_3846);
nand U4671 (N_4671,N_3476,N_3893);
or U4672 (N_4672,N_3199,N_3991);
or U4673 (N_4673,N_3011,N_3902);
nand U4674 (N_4674,N_3497,N_3204);
or U4675 (N_4675,N_3122,N_3253);
nand U4676 (N_4676,N_3208,N_3836);
or U4677 (N_4677,N_3008,N_3682);
nor U4678 (N_4678,N_3857,N_3542);
nor U4679 (N_4679,N_3286,N_3855);
nor U4680 (N_4680,N_3980,N_3457);
xor U4681 (N_4681,N_3355,N_3223);
nand U4682 (N_4682,N_3938,N_3551);
and U4683 (N_4683,N_3598,N_3912);
nand U4684 (N_4684,N_3837,N_3561);
and U4685 (N_4685,N_3687,N_3905);
and U4686 (N_4686,N_3493,N_3187);
nor U4687 (N_4687,N_3339,N_3032);
xor U4688 (N_4688,N_3819,N_3057);
or U4689 (N_4689,N_3560,N_3162);
nor U4690 (N_4690,N_3454,N_3144);
and U4691 (N_4691,N_3071,N_3284);
xor U4692 (N_4692,N_3234,N_3595);
or U4693 (N_4693,N_3652,N_3211);
xnor U4694 (N_4694,N_3364,N_3370);
and U4695 (N_4695,N_3071,N_3897);
nand U4696 (N_4696,N_3084,N_3406);
nor U4697 (N_4697,N_3957,N_3257);
xor U4698 (N_4698,N_3526,N_3871);
nand U4699 (N_4699,N_3404,N_3119);
nand U4700 (N_4700,N_3379,N_3548);
xor U4701 (N_4701,N_3660,N_3132);
and U4702 (N_4702,N_3688,N_3656);
or U4703 (N_4703,N_3025,N_3441);
or U4704 (N_4704,N_3420,N_3917);
xor U4705 (N_4705,N_3174,N_3761);
or U4706 (N_4706,N_3616,N_3465);
nand U4707 (N_4707,N_3004,N_3095);
nor U4708 (N_4708,N_3719,N_3128);
nand U4709 (N_4709,N_3257,N_3853);
or U4710 (N_4710,N_3316,N_3925);
nand U4711 (N_4711,N_3713,N_3268);
nand U4712 (N_4712,N_3850,N_3839);
nand U4713 (N_4713,N_3827,N_3141);
nor U4714 (N_4714,N_3562,N_3527);
or U4715 (N_4715,N_3433,N_3752);
or U4716 (N_4716,N_3733,N_3421);
xnor U4717 (N_4717,N_3223,N_3518);
or U4718 (N_4718,N_3051,N_3400);
and U4719 (N_4719,N_3590,N_3421);
nor U4720 (N_4720,N_3847,N_3443);
or U4721 (N_4721,N_3408,N_3971);
and U4722 (N_4722,N_3850,N_3600);
and U4723 (N_4723,N_3291,N_3323);
and U4724 (N_4724,N_3310,N_3092);
nor U4725 (N_4725,N_3869,N_3346);
nor U4726 (N_4726,N_3772,N_3640);
and U4727 (N_4727,N_3437,N_3930);
nor U4728 (N_4728,N_3971,N_3551);
nor U4729 (N_4729,N_3890,N_3276);
nand U4730 (N_4730,N_3342,N_3009);
nor U4731 (N_4731,N_3110,N_3916);
or U4732 (N_4732,N_3707,N_3918);
and U4733 (N_4733,N_3077,N_3928);
or U4734 (N_4734,N_3150,N_3440);
nor U4735 (N_4735,N_3863,N_3745);
nor U4736 (N_4736,N_3988,N_3105);
xnor U4737 (N_4737,N_3150,N_3428);
and U4738 (N_4738,N_3955,N_3992);
and U4739 (N_4739,N_3178,N_3952);
or U4740 (N_4740,N_3872,N_3241);
nand U4741 (N_4741,N_3293,N_3842);
or U4742 (N_4742,N_3069,N_3454);
and U4743 (N_4743,N_3028,N_3208);
nor U4744 (N_4744,N_3169,N_3119);
and U4745 (N_4745,N_3580,N_3641);
or U4746 (N_4746,N_3869,N_3538);
nand U4747 (N_4747,N_3011,N_3852);
and U4748 (N_4748,N_3030,N_3932);
xnor U4749 (N_4749,N_3036,N_3076);
or U4750 (N_4750,N_3287,N_3206);
nand U4751 (N_4751,N_3869,N_3331);
nand U4752 (N_4752,N_3655,N_3239);
nand U4753 (N_4753,N_3606,N_3013);
nand U4754 (N_4754,N_3350,N_3137);
nor U4755 (N_4755,N_3648,N_3728);
and U4756 (N_4756,N_3416,N_3601);
and U4757 (N_4757,N_3335,N_3420);
nor U4758 (N_4758,N_3427,N_3484);
xnor U4759 (N_4759,N_3688,N_3834);
and U4760 (N_4760,N_3154,N_3856);
or U4761 (N_4761,N_3296,N_3370);
and U4762 (N_4762,N_3793,N_3118);
nand U4763 (N_4763,N_3215,N_3583);
nor U4764 (N_4764,N_3905,N_3018);
nand U4765 (N_4765,N_3059,N_3146);
and U4766 (N_4766,N_3991,N_3226);
and U4767 (N_4767,N_3101,N_3454);
and U4768 (N_4768,N_3095,N_3841);
or U4769 (N_4769,N_3683,N_3026);
nor U4770 (N_4770,N_3162,N_3614);
and U4771 (N_4771,N_3168,N_3494);
and U4772 (N_4772,N_3238,N_3227);
nand U4773 (N_4773,N_3941,N_3667);
or U4774 (N_4774,N_3314,N_3357);
or U4775 (N_4775,N_3171,N_3610);
xor U4776 (N_4776,N_3783,N_3222);
and U4777 (N_4777,N_3133,N_3817);
nand U4778 (N_4778,N_3378,N_3965);
nor U4779 (N_4779,N_3830,N_3069);
nor U4780 (N_4780,N_3217,N_3944);
or U4781 (N_4781,N_3677,N_3842);
xnor U4782 (N_4782,N_3126,N_3916);
or U4783 (N_4783,N_3313,N_3960);
xor U4784 (N_4784,N_3995,N_3564);
xnor U4785 (N_4785,N_3841,N_3001);
nand U4786 (N_4786,N_3248,N_3505);
or U4787 (N_4787,N_3540,N_3322);
and U4788 (N_4788,N_3622,N_3072);
nand U4789 (N_4789,N_3767,N_3982);
or U4790 (N_4790,N_3712,N_3786);
nand U4791 (N_4791,N_3747,N_3895);
xor U4792 (N_4792,N_3137,N_3080);
or U4793 (N_4793,N_3341,N_3600);
nor U4794 (N_4794,N_3321,N_3856);
nor U4795 (N_4795,N_3530,N_3681);
or U4796 (N_4796,N_3229,N_3835);
or U4797 (N_4797,N_3385,N_3420);
or U4798 (N_4798,N_3018,N_3949);
xor U4799 (N_4799,N_3557,N_3282);
nand U4800 (N_4800,N_3836,N_3841);
xnor U4801 (N_4801,N_3736,N_3488);
xor U4802 (N_4802,N_3059,N_3150);
nand U4803 (N_4803,N_3968,N_3971);
xor U4804 (N_4804,N_3360,N_3988);
nor U4805 (N_4805,N_3697,N_3402);
nor U4806 (N_4806,N_3847,N_3373);
xnor U4807 (N_4807,N_3301,N_3420);
nor U4808 (N_4808,N_3112,N_3516);
and U4809 (N_4809,N_3892,N_3614);
xnor U4810 (N_4810,N_3452,N_3891);
or U4811 (N_4811,N_3017,N_3742);
and U4812 (N_4812,N_3692,N_3031);
nor U4813 (N_4813,N_3491,N_3954);
nand U4814 (N_4814,N_3130,N_3855);
nor U4815 (N_4815,N_3866,N_3750);
or U4816 (N_4816,N_3871,N_3585);
nand U4817 (N_4817,N_3470,N_3312);
xnor U4818 (N_4818,N_3051,N_3594);
nor U4819 (N_4819,N_3095,N_3225);
nand U4820 (N_4820,N_3044,N_3767);
xor U4821 (N_4821,N_3494,N_3057);
xor U4822 (N_4822,N_3415,N_3167);
nor U4823 (N_4823,N_3544,N_3859);
or U4824 (N_4824,N_3265,N_3082);
nor U4825 (N_4825,N_3052,N_3797);
or U4826 (N_4826,N_3522,N_3831);
nor U4827 (N_4827,N_3406,N_3618);
or U4828 (N_4828,N_3192,N_3305);
and U4829 (N_4829,N_3069,N_3288);
xnor U4830 (N_4830,N_3422,N_3394);
nor U4831 (N_4831,N_3351,N_3786);
and U4832 (N_4832,N_3474,N_3620);
and U4833 (N_4833,N_3589,N_3577);
xnor U4834 (N_4834,N_3294,N_3302);
xor U4835 (N_4835,N_3862,N_3831);
and U4836 (N_4836,N_3559,N_3980);
or U4837 (N_4837,N_3875,N_3825);
xor U4838 (N_4838,N_3014,N_3603);
nand U4839 (N_4839,N_3985,N_3349);
or U4840 (N_4840,N_3766,N_3652);
nor U4841 (N_4841,N_3509,N_3495);
xor U4842 (N_4842,N_3293,N_3226);
xor U4843 (N_4843,N_3383,N_3216);
xor U4844 (N_4844,N_3400,N_3577);
and U4845 (N_4845,N_3934,N_3926);
xnor U4846 (N_4846,N_3930,N_3989);
or U4847 (N_4847,N_3579,N_3499);
xnor U4848 (N_4848,N_3250,N_3342);
and U4849 (N_4849,N_3837,N_3804);
nor U4850 (N_4850,N_3712,N_3406);
xor U4851 (N_4851,N_3592,N_3850);
or U4852 (N_4852,N_3534,N_3543);
nand U4853 (N_4853,N_3828,N_3281);
xnor U4854 (N_4854,N_3440,N_3962);
nor U4855 (N_4855,N_3058,N_3757);
and U4856 (N_4856,N_3507,N_3435);
and U4857 (N_4857,N_3212,N_3971);
nor U4858 (N_4858,N_3086,N_3850);
nor U4859 (N_4859,N_3644,N_3371);
xnor U4860 (N_4860,N_3337,N_3668);
or U4861 (N_4861,N_3292,N_3397);
or U4862 (N_4862,N_3446,N_3043);
nor U4863 (N_4863,N_3091,N_3506);
xor U4864 (N_4864,N_3848,N_3389);
nor U4865 (N_4865,N_3168,N_3728);
nand U4866 (N_4866,N_3224,N_3557);
or U4867 (N_4867,N_3728,N_3312);
nand U4868 (N_4868,N_3185,N_3122);
nor U4869 (N_4869,N_3030,N_3451);
xor U4870 (N_4870,N_3569,N_3194);
xor U4871 (N_4871,N_3868,N_3292);
xnor U4872 (N_4872,N_3001,N_3136);
and U4873 (N_4873,N_3136,N_3721);
nor U4874 (N_4874,N_3497,N_3683);
or U4875 (N_4875,N_3081,N_3811);
xnor U4876 (N_4876,N_3097,N_3861);
nor U4877 (N_4877,N_3305,N_3314);
and U4878 (N_4878,N_3035,N_3396);
and U4879 (N_4879,N_3333,N_3530);
or U4880 (N_4880,N_3392,N_3381);
and U4881 (N_4881,N_3780,N_3724);
nor U4882 (N_4882,N_3631,N_3246);
xnor U4883 (N_4883,N_3113,N_3307);
or U4884 (N_4884,N_3629,N_3715);
nand U4885 (N_4885,N_3340,N_3676);
nand U4886 (N_4886,N_3327,N_3510);
nand U4887 (N_4887,N_3098,N_3976);
xnor U4888 (N_4888,N_3723,N_3437);
and U4889 (N_4889,N_3206,N_3593);
xnor U4890 (N_4890,N_3235,N_3113);
nor U4891 (N_4891,N_3154,N_3021);
or U4892 (N_4892,N_3934,N_3052);
nand U4893 (N_4893,N_3722,N_3021);
or U4894 (N_4894,N_3126,N_3882);
xor U4895 (N_4895,N_3455,N_3629);
xnor U4896 (N_4896,N_3106,N_3370);
nor U4897 (N_4897,N_3644,N_3075);
or U4898 (N_4898,N_3432,N_3106);
and U4899 (N_4899,N_3972,N_3267);
and U4900 (N_4900,N_3057,N_3220);
nand U4901 (N_4901,N_3309,N_3829);
nor U4902 (N_4902,N_3458,N_3494);
nor U4903 (N_4903,N_3128,N_3539);
nand U4904 (N_4904,N_3980,N_3903);
xnor U4905 (N_4905,N_3517,N_3716);
nor U4906 (N_4906,N_3054,N_3475);
xor U4907 (N_4907,N_3309,N_3824);
nand U4908 (N_4908,N_3425,N_3603);
nor U4909 (N_4909,N_3582,N_3872);
xnor U4910 (N_4910,N_3857,N_3198);
or U4911 (N_4911,N_3723,N_3234);
and U4912 (N_4912,N_3690,N_3370);
or U4913 (N_4913,N_3082,N_3902);
nor U4914 (N_4914,N_3264,N_3013);
and U4915 (N_4915,N_3415,N_3475);
nand U4916 (N_4916,N_3589,N_3915);
or U4917 (N_4917,N_3755,N_3272);
and U4918 (N_4918,N_3886,N_3313);
xor U4919 (N_4919,N_3149,N_3216);
nand U4920 (N_4920,N_3354,N_3310);
xor U4921 (N_4921,N_3492,N_3215);
nand U4922 (N_4922,N_3956,N_3948);
or U4923 (N_4923,N_3448,N_3938);
nand U4924 (N_4924,N_3522,N_3816);
nand U4925 (N_4925,N_3831,N_3704);
nor U4926 (N_4926,N_3556,N_3566);
nand U4927 (N_4927,N_3464,N_3186);
and U4928 (N_4928,N_3617,N_3416);
xor U4929 (N_4929,N_3279,N_3140);
and U4930 (N_4930,N_3759,N_3310);
nor U4931 (N_4931,N_3171,N_3631);
nor U4932 (N_4932,N_3304,N_3473);
xor U4933 (N_4933,N_3006,N_3057);
nand U4934 (N_4934,N_3873,N_3267);
or U4935 (N_4935,N_3981,N_3899);
and U4936 (N_4936,N_3150,N_3291);
and U4937 (N_4937,N_3342,N_3192);
and U4938 (N_4938,N_3795,N_3331);
or U4939 (N_4939,N_3691,N_3323);
or U4940 (N_4940,N_3326,N_3492);
and U4941 (N_4941,N_3842,N_3611);
or U4942 (N_4942,N_3462,N_3552);
nor U4943 (N_4943,N_3278,N_3675);
or U4944 (N_4944,N_3218,N_3286);
and U4945 (N_4945,N_3204,N_3623);
xnor U4946 (N_4946,N_3703,N_3383);
nand U4947 (N_4947,N_3727,N_3406);
nor U4948 (N_4948,N_3335,N_3375);
xor U4949 (N_4949,N_3440,N_3663);
and U4950 (N_4950,N_3569,N_3311);
or U4951 (N_4951,N_3617,N_3500);
and U4952 (N_4952,N_3669,N_3139);
nor U4953 (N_4953,N_3310,N_3724);
or U4954 (N_4954,N_3891,N_3651);
and U4955 (N_4955,N_3568,N_3144);
and U4956 (N_4956,N_3502,N_3397);
or U4957 (N_4957,N_3129,N_3867);
or U4958 (N_4958,N_3793,N_3447);
and U4959 (N_4959,N_3936,N_3772);
or U4960 (N_4960,N_3548,N_3735);
or U4961 (N_4961,N_3399,N_3564);
nand U4962 (N_4962,N_3140,N_3259);
nor U4963 (N_4963,N_3550,N_3380);
xor U4964 (N_4964,N_3044,N_3037);
nand U4965 (N_4965,N_3933,N_3695);
and U4966 (N_4966,N_3661,N_3893);
xnor U4967 (N_4967,N_3518,N_3477);
or U4968 (N_4968,N_3596,N_3196);
nor U4969 (N_4969,N_3088,N_3028);
or U4970 (N_4970,N_3843,N_3670);
and U4971 (N_4971,N_3196,N_3779);
xnor U4972 (N_4972,N_3205,N_3734);
nor U4973 (N_4973,N_3045,N_3166);
and U4974 (N_4974,N_3291,N_3361);
nand U4975 (N_4975,N_3422,N_3295);
and U4976 (N_4976,N_3092,N_3003);
or U4977 (N_4977,N_3576,N_3854);
nand U4978 (N_4978,N_3083,N_3971);
or U4979 (N_4979,N_3486,N_3998);
and U4980 (N_4980,N_3241,N_3449);
nor U4981 (N_4981,N_3131,N_3207);
xor U4982 (N_4982,N_3791,N_3475);
and U4983 (N_4983,N_3419,N_3132);
and U4984 (N_4984,N_3823,N_3808);
or U4985 (N_4985,N_3559,N_3254);
and U4986 (N_4986,N_3684,N_3476);
xor U4987 (N_4987,N_3791,N_3554);
or U4988 (N_4988,N_3723,N_3328);
nand U4989 (N_4989,N_3399,N_3933);
or U4990 (N_4990,N_3715,N_3198);
or U4991 (N_4991,N_3386,N_3273);
and U4992 (N_4992,N_3641,N_3284);
or U4993 (N_4993,N_3081,N_3276);
or U4994 (N_4994,N_3796,N_3239);
and U4995 (N_4995,N_3367,N_3661);
or U4996 (N_4996,N_3278,N_3616);
or U4997 (N_4997,N_3384,N_3897);
xnor U4998 (N_4998,N_3436,N_3030);
nor U4999 (N_4999,N_3396,N_3322);
or U5000 (N_5000,N_4864,N_4951);
and U5001 (N_5001,N_4046,N_4200);
and U5002 (N_5002,N_4796,N_4909);
nor U5003 (N_5003,N_4869,N_4925);
nand U5004 (N_5004,N_4654,N_4936);
or U5005 (N_5005,N_4192,N_4375);
and U5006 (N_5006,N_4014,N_4761);
nand U5007 (N_5007,N_4444,N_4636);
or U5008 (N_5008,N_4231,N_4672);
nor U5009 (N_5009,N_4013,N_4763);
xnor U5010 (N_5010,N_4197,N_4342);
xor U5011 (N_5011,N_4582,N_4183);
nor U5012 (N_5012,N_4798,N_4259);
and U5013 (N_5013,N_4256,N_4136);
nor U5014 (N_5014,N_4392,N_4324);
xnor U5015 (N_5015,N_4993,N_4077);
nor U5016 (N_5016,N_4190,N_4076);
and U5017 (N_5017,N_4308,N_4310);
xnor U5018 (N_5018,N_4056,N_4641);
and U5019 (N_5019,N_4495,N_4617);
nand U5020 (N_5020,N_4009,N_4890);
nor U5021 (N_5021,N_4861,N_4750);
or U5022 (N_5022,N_4346,N_4002);
xor U5023 (N_5023,N_4174,N_4773);
and U5024 (N_5024,N_4915,N_4648);
nand U5025 (N_5025,N_4599,N_4221);
xnor U5026 (N_5026,N_4363,N_4880);
and U5027 (N_5027,N_4838,N_4911);
and U5028 (N_5028,N_4998,N_4003);
or U5029 (N_5029,N_4224,N_4433);
nor U5030 (N_5030,N_4906,N_4974);
or U5031 (N_5031,N_4952,N_4932);
xnor U5032 (N_5032,N_4338,N_4788);
nand U5033 (N_5033,N_4534,N_4218);
xor U5034 (N_5034,N_4461,N_4341);
and U5035 (N_5035,N_4419,N_4188);
and U5036 (N_5036,N_4910,N_4859);
or U5037 (N_5037,N_4947,N_4748);
nor U5038 (N_5038,N_4185,N_4724);
xnor U5039 (N_5039,N_4178,N_4128);
xor U5040 (N_5040,N_4460,N_4887);
xnor U5041 (N_5041,N_4250,N_4849);
or U5042 (N_5042,N_4867,N_4557);
and U5043 (N_5043,N_4704,N_4559);
and U5044 (N_5044,N_4543,N_4402);
nand U5045 (N_5045,N_4105,N_4085);
nand U5046 (N_5046,N_4209,N_4030);
and U5047 (N_5047,N_4248,N_4094);
nand U5048 (N_5048,N_4561,N_4758);
xnor U5049 (N_5049,N_4370,N_4286);
or U5050 (N_5050,N_4583,N_4605);
or U5051 (N_5051,N_4022,N_4143);
nor U5052 (N_5052,N_4431,N_4067);
xor U5053 (N_5053,N_4207,N_4088);
nand U5054 (N_5054,N_4538,N_4327);
or U5055 (N_5055,N_4558,N_4570);
or U5056 (N_5056,N_4113,N_4501);
nor U5057 (N_5057,N_4752,N_4836);
xor U5058 (N_5058,N_4108,N_4294);
and U5059 (N_5059,N_4670,N_4420);
and U5060 (N_5060,N_4114,N_4851);
and U5061 (N_5061,N_4302,N_4789);
or U5062 (N_5062,N_4516,N_4845);
or U5063 (N_5063,N_4186,N_4973);
nand U5064 (N_5064,N_4611,N_4142);
xnor U5065 (N_5065,N_4512,N_4098);
nand U5066 (N_5066,N_4903,N_4151);
or U5067 (N_5067,N_4463,N_4615);
or U5068 (N_5068,N_4918,N_4580);
nor U5069 (N_5069,N_4667,N_4691);
nand U5070 (N_5070,N_4596,N_4959);
nor U5071 (N_5071,N_4817,N_4235);
nand U5072 (N_5072,N_4391,N_4692);
and U5073 (N_5073,N_4297,N_4874);
or U5074 (N_5074,N_4282,N_4535);
and U5075 (N_5075,N_4233,N_4548);
nor U5076 (N_5076,N_4709,N_4336);
xnor U5077 (N_5077,N_4124,N_4782);
nor U5078 (N_5078,N_4530,N_4048);
or U5079 (N_5079,N_4746,N_4627);
and U5080 (N_5080,N_4793,N_4162);
nor U5081 (N_5081,N_4245,N_4977);
nor U5082 (N_5082,N_4766,N_4774);
nor U5083 (N_5083,N_4533,N_4117);
and U5084 (N_5084,N_4157,N_4702);
nor U5085 (N_5085,N_4191,N_4304);
or U5086 (N_5086,N_4340,N_4787);
nand U5087 (N_5087,N_4007,N_4799);
nor U5088 (N_5088,N_4892,N_4870);
nand U5089 (N_5089,N_4837,N_4924);
and U5090 (N_5090,N_4521,N_4155);
nor U5091 (N_5091,N_4883,N_4412);
and U5092 (N_5092,N_4919,N_4115);
nand U5093 (N_5093,N_4161,N_4531);
nor U5094 (N_5094,N_4179,N_4971);
nor U5095 (N_5095,N_4265,N_4352);
nor U5096 (N_5096,N_4290,N_4868);
and U5097 (N_5097,N_4445,N_4622);
nor U5098 (N_5098,N_4283,N_4006);
and U5099 (N_5099,N_4413,N_4442);
or U5100 (N_5100,N_4242,N_4180);
nor U5101 (N_5101,N_4705,N_4372);
and U5102 (N_5102,N_4339,N_4464);
nor U5103 (N_5103,N_4872,N_4497);
and U5104 (N_5104,N_4134,N_4866);
and U5105 (N_5105,N_4285,N_4549);
and U5106 (N_5106,N_4454,N_4011);
nand U5107 (N_5107,N_4061,N_4216);
and U5108 (N_5108,N_4386,N_4726);
nand U5109 (N_5109,N_4620,N_4275);
nand U5110 (N_5110,N_4163,N_4542);
nor U5111 (N_5111,N_4312,N_4417);
nor U5112 (N_5112,N_4194,N_4945);
or U5113 (N_5113,N_4689,N_4853);
xnor U5114 (N_5114,N_4358,N_4320);
and U5115 (N_5115,N_4368,N_4537);
or U5116 (N_5116,N_4121,N_4978);
or U5117 (N_5117,N_4095,N_4371);
nand U5118 (N_5118,N_4650,N_4768);
nor U5119 (N_5119,N_4057,N_4070);
and U5120 (N_5120,N_4100,N_4741);
nand U5121 (N_5121,N_4377,N_4955);
or U5122 (N_5122,N_4626,N_4008);
nor U5123 (N_5123,N_4567,N_4465);
and U5124 (N_5124,N_4860,N_4062);
and U5125 (N_5125,N_4840,N_4471);
nor U5126 (N_5126,N_4828,N_4019);
or U5127 (N_5127,N_4529,N_4571);
xnor U5128 (N_5128,N_4226,N_4393);
xor U5129 (N_5129,N_4292,N_4314);
nor U5130 (N_5130,N_4991,N_4655);
xor U5131 (N_5131,N_4408,N_4806);
and U5132 (N_5132,N_4450,N_4624);
and U5133 (N_5133,N_4982,N_4629);
nor U5134 (N_5134,N_4976,N_4271);
nand U5135 (N_5135,N_4418,N_4676);
and U5136 (N_5136,N_4159,N_4749);
nor U5137 (N_5137,N_4387,N_4255);
or U5138 (N_5138,N_4988,N_4589);
nor U5139 (N_5139,N_4457,N_4089);
or U5140 (N_5140,N_4263,N_4050);
xnor U5141 (N_5141,N_4715,N_4810);
or U5142 (N_5142,N_4335,N_4281);
or U5143 (N_5143,N_4274,N_4997);
or U5144 (N_5144,N_4225,N_4720);
nor U5145 (N_5145,N_4894,N_4922);
or U5146 (N_5146,N_4833,N_4045);
nand U5147 (N_5147,N_4034,N_4760);
or U5148 (N_5148,N_4477,N_4244);
nand U5149 (N_5149,N_4764,N_4829);
and U5150 (N_5150,N_4176,N_4299);
nor U5151 (N_5151,N_4972,N_4239);
nor U5152 (N_5152,N_4928,N_4917);
nand U5153 (N_5153,N_4528,N_4814);
and U5154 (N_5154,N_4981,N_4276);
nand U5155 (N_5155,N_4807,N_4104);
xor U5156 (N_5156,N_4133,N_4850);
nor U5157 (N_5157,N_4153,N_4222);
and U5158 (N_5158,N_4364,N_4958);
nor U5159 (N_5159,N_4323,N_4278);
nand U5160 (N_5160,N_4141,N_4343);
xnor U5161 (N_5161,N_4588,N_4914);
and U5162 (N_5162,N_4688,N_4926);
nor U5163 (N_5163,N_4303,N_4205);
or U5164 (N_5164,N_4356,N_4171);
nand U5165 (N_5165,N_4632,N_4354);
nor U5166 (N_5166,N_4819,N_4434);
xor U5167 (N_5167,N_4122,N_4373);
xor U5168 (N_5168,N_4662,N_4421);
nand U5169 (N_5169,N_4081,N_4489);
xnor U5170 (N_5170,N_4016,N_4490);
nand U5171 (N_5171,N_4778,N_4734);
or U5172 (N_5172,N_4266,N_4904);
nor U5173 (N_5173,N_4269,N_4069);
or U5174 (N_5174,N_4964,N_4772);
or U5175 (N_5175,N_4996,N_4573);
and U5176 (N_5176,N_4227,N_4249);
or U5177 (N_5177,N_4131,N_4443);
nor U5178 (N_5178,N_4992,N_4468);
nor U5179 (N_5179,N_4287,N_4895);
xnor U5180 (N_5180,N_4051,N_4683);
xnor U5181 (N_5181,N_4252,N_4695);
nand U5182 (N_5182,N_4084,N_4639);
nor U5183 (N_5183,N_4873,N_4505);
and U5184 (N_5184,N_4172,N_4148);
nand U5185 (N_5185,N_4506,N_4601);
and U5186 (N_5186,N_4321,N_4270);
nor U5187 (N_5187,N_4110,N_4515);
nand U5188 (N_5188,N_4762,N_4732);
nor U5189 (N_5189,N_4469,N_4129);
nand U5190 (N_5190,N_4968,N_4811);
and U5191 (N_5191,N_4722,N_4839);
nand U5192 (N_5192,N_4033,N_4415);
nand U5193 (N_5193,N_4842,N_4488);
nand U5194 (N_5194,N_4899,N_4927);
or U5195 (N_5195,N_4078,N_4306);
xnor U5196 (N_5196,N_4618,N_4594);
xor U5197 (N_5197,N_4169,N_4995);
nand U5198 (N_5198,N_4504,N_4254);
nor U5199 (N_5199,N_4448,N_4714);
and U5200 (N_5200,N_4429,N_4809);
and U5201 (N_5201,N_4877,N_4541);
nand U5202 (N_5202,N_4210,N_4332);
xor U5203 (N_5203,N_4073,N_4160);
nor U5204 (N_5204,N_4446,N_4625);
nand U5205 (N_5205,N_4884,N_4074);
and U5206 (N_5206,N_4289,N_4147);
nor U5207 (N_5207,N_4735,N_4491);
xor U5208 (N_5208,N_4930,N_4536);
nor U5209 (N_5209,N_4264,N_4103);
nand U5210 (N_5210,N_4856,N_4039);
xor U5211 (N_5211,N_4712,N_4195);
xnor U5212 (N_5212,N_4272,N_4765);
and U5213 (N_5213,N_4309,N_4954);
or U5214 (N_5214,N_4507,N_4158);
nor U5215 (N_5215,N_4994,N_4027);
nand U5216 (N_5216,N_4745,N_4687);
nand U5217 (N_5217,N_4711,N_4637);
or U5218 (N_5218,N_4487,N_4767);
nand U5219 (N_5219,N_4154,N_4660);
nor U5220 (N_5220,N_4219,N_4140);
or U5221 (N_5221,N_4719,N_4815);
xor U5222 (N_5222,N_4923,N_4032);
nor U5223 (N_5223,N_4737,N_4018);
nor U5224 (N_5224,N_4168,N_4485);
nand U5225 (N_5225,N_4424,N_4293);
and U5226 (N_5226,N_4781,N_4345);
and U5227 (N_5227,N_4990,N_4025);
and U5228 (N_5228,N_4579,N_4822);
nor U5229 (N_5229,N_4355,N_4730);
nor U5230 (N_5230,N_4987,N_4747);
nand U5231 (N_5231,N_4005,N_4437);
or U5232 (N_5232,N_4079,N_4891);
nand U5233 (N_5233,N_4937,N_4674);
nand U5234 (N_5234,N_4623,N_4328);
and U5235 (N_5235,N_4483,N_4847);
and U5236 (N_5236,N_4280,N_4344);
nand U5237 (N_5237,N_4820,N_4396);
nor U5238 (N_5238,N_4566,N_4843);
or U5239 (N_5239,N_4524,N_4590);
nor U5240 (N_5240,N_4832,N_4610);
xnor U5241 (N_5241,N_4347,N_4826);
nand U5242 (N_5242,N_4948,N_4825);
and U5243 (N_5243,N_4112,N_4152);
nor U5244 (N_5244,N_4333,N_4539);
xnor U5245 (N_5245,N_4021,N_4956);
xor U5246 (N_5246,N_4325,N_4931);
nand U5247 (N_5247,N_4241,N_4585);
nand U5248 (N_5248,N_4587,N_4693);
xor U5249 (N_5249,N_4379,N_4776);
xor U5250 (N_5250,N_4196,N_4770);
or U5251 (N_5251,N_4812,N_4149);
and U5252 (N_5252,N_4970,N_4686);
and U5253 (N_5253,N_4779,N_4311);
xor U5254 (N_5254,N_4775,N_4545);
or U5255 (N_5255,N_4075,N_4498);
xnor U5256 (N_5256,N_4633,N_4564);
and U5257 (N_5257,N_4438,N_4664);
and U5258 (N_5258,N_4756,N_4889);
xor U5259 (N_5259,N_4823,N_4784);
nand U5260 (N_5260,N_4298,N_4026);
and U5261 (N_5261,N_4012,N_4404);
and U5262 (N_5262,N_4044,N_4351);
xnor U5263 (N_5263,N_4795,N_4661);
or U5264 (N_5264,N_4532,N_4929);
nand U5265 (N_5265,N_4150,N_4120);
nand U5266 (N_5266,N_4246,N_4020);
or U5267 (N_5267,N_4059,N_4651);
xor U5268 (N_5268,N_4606,N_4879);
or U5269 (N_5269,N_4232,N_4472);
nor U5270 (N_5270,N_4902,N_4729);
nor U5271 (N_5271,N_4844,N_4983);
xor U5272 (N_5272,N_4634,N_4436);
and U5273 (N_5273,N_4106,N_4223);
nand U5274 (N_5274,N_4499,N_4562);
and U5275 (N_5275,N_4156,N_4273);
nand U5276 (N_5276,N_4757,N_4547);
or U5277 (N_5277,N_4102,N_4854);
or U5278 (N_5278,N_4514,N_4360);
nor U5279 (N_5279,N_4934,N_4804);
xor U5280 (N_5280,N_4721,N_4522);
or U5281 (N_5281,N_4646,N_4382);
and U5282 (N_5282,N_4574,N_4049);
nand U5283 (N_5283,N_4199,N_4119);
nor U5284 (N_5284,N_4551,N_4953);
nor U5285 (N_5285,N_4440,N_4912);
nand U5286 (N_5286,N_4685,N_4941);
xor U5287 (N_5287,N_4619,N_4790);
nand U5288 (N_5288,N_4572,N_4432);
and U5289 (N_5289,N_4410,N_4068);
nor U5290 (N_5290,N_4201,N_4656);
or U5291 (N_5291,N_4097,N_4944);
xnor U5292 (N_5292,N_4550,N_4659);
and U5293 (N_5293,N_4001,N_4093);
xnor U5294 (N_5294,N_4486,N_4791);
xor U5295 (N_5295,N_4603,N_4349);
or U5296 (N_5296,N_4666,N_4565);
nand U5297 (N_5297,N_4510,N_4898);
xor U5298 (N_5298,N_4901,N_4214);
or U5299 (N_5299,N_4337,N_4933);
nor U5300 (N_5300,N_4015,N_4665);
nand U5301 (N_5301,N_4043,N_4058);
and U5302 (N_5302,N_4613,N_4206);
or U5303 (N_5303,N_4690,N_4525);
and U5304 (N_5304,N_4479,N_4876);
xor U5305 (N_5305,N_4247,N_4397);
and U5306 (N_5306,N_4608,N_4401);
nor U5307 (N_5307,N_4717,N_4780);
nor U5308 (N_5308,N_4319,N_4376);
nor U5309 (N_5309,N_4458,N_4064);
or U5310 (N_5310,N_4852,N_4643);
xnor U5311 (N_5311,N_4649,N_4288);
nand U5312 (N_5312,N_4638,N_4706);
nand U5313 (N_5313,N_4130,N_4389);
xor U5314 (N_5314,N_4359,N_4082);
or U5315 (N_5315,N_4985,N_4885);
and U5316 (N_5316,N_4546,N_4586);
nor U5317 (N_5317,N_4848,N_4494);
xnor U5318 (N_5318,N_4357,N_4694);
nand U5319 (N_5319,N_4165,N_4967);
nor U5320 (N_5320,N_4957,N_4307);
nand U5321 (N_5321,N_4897,N_4071);
and U5322 (N_5322,N_4331,N_4380);
or U5323 (N_5323,N_4063,N_4592);
or U5324 (N_5324,N_4710,N_4353);
or U5325 (N_5325,N_4581,N_4520);
or U5326 (N_5326,N_4220,N_4803);
nor U5327 (N_5327,N_4399,N_4184);
and U5328 (N_5328,N_4805,N_4965);
xor U5329 (N_5329,N_4125,N_4801);
nand U5330 (N_5330,N_4708,N_4631);
xor U5331 (N_5331,N_4447,N_4426);
or U5332 (N_5332,N_4427,N_4042);
and U5333 (N_5333,N_4028,N_4913);
and U5334 (N_5334,N_4701,N_4198);
nor U5335 (N_5335,N_4086,N_4466);
xor U5336 (N_5336,N_4630,N_4480);
nand U5337 (N_5337,N_4317,N_4657);
nor U5338 (N_5338,N_4699,N_4474);
nor U5339 (N_5339,N_4475,N_4846);
and U5340 (N_5340,N_4313,N_4509);
xnor U5341 (N_5341,N_4260,N_4553);
or U5342 (N_5342,N_4166,N_4663);
or U5343 (N_5343,N_4578,N_4361);
nand U5344 (N_5344,N_4523,N_4065);
or U5345 (N_5345,N_4350,N_4743);
nand U5346 (N_5346,N_4144,N_4544);
xor U5347 (N_5347,N_4609,N_4821);
xnor U5348 (N_5348,N_4511,N_4430);
and U5349 (N_5349,N_4786,N_4326);
nand U5350 (N_5350,N_4939,N_4723);
and U5351 (N_5351,N_4644,N_4900);
and U5352 (N_5352,N_4137,N_4513);
nand U5353 (N_5353,N_4476,N_4671);
xor U5354 (N_5354,N_4301,N_4769);
nor U5355 (N_5355,N_4023,N_4211);
nor U5356 (N_5356,N_4496,N_4940);
or U5357 (N_5357,N_4481,N_4212);
and U5358 (N_5358,N_4568,N_4060);
or U5359 (N_5359,N_4946,N_4645);
and U5360 (N_5360,N_4236,N_4208);
nor U5361 (N_5361,N_4237,N_4405);
nand U5362 (N_5362,N_4083,N_4334);
xor U5363 (N_5363,N_4193,N_4000);
nand U5364 (N_5364,N_4595,N_4484);
xor U5365 (N_5365,N_4593,N_4938);
or U5366 (N_5366,N_4673,N_4950);
xor U5367 (N_5367,N_4855,N_4680);
nand U5368 (N_5368,N_4284,N_4575);
xnor U5369 (N_5369,N_4871,N_4203);
xnor U5370 (N_5370,N_4441,N_4451);
or U5371 (N_5371,N_4600,N_4920);
or U5372 (N_5372,N_4228,N_4777);
or U5373 (N_5373,N_4123,N_4696);
nand U5374 (N_5374,N_4697,N_4725);
xnor U5375 (N_5375,N_4099,N_4738);
and U5376 (N_5376,N_4213,N_4234);
nand U5377 (N_5377,N_4090,N_4107);
nor U5378 (N_5378,N_4942,N_4116);
and U5379 (N_5379,N_4508,N_4759);
xor U5380 (N_5380,N_4614,N_4467);
nor U5381 (N_5381,N_4830,N_4949);
nand U5382 (N_5382,N_4818,N_4388);
xor U5383 (N_5383,N_4217,N_4604);
and U5384 (N_5384,N_4591,N_4518);
and U5385 (N_5385,N_4986,N_4727);
nor U5386 (N_5386,N_4669,N_4792);
and U5387 (N_5387,N_4554,N_4841);
or U5388 (N_5388,N_4398,N_4439);
nor U5389 (N_5389,N_4091,N_4167);
and U5390 (N_5390,N_4362,N_4975);
nor U5391 (N_5391,N_4041,N_4517);
nor U5392 (N_5392,N_4602,N_4989);
and U5393 (N_5393,N_4492,N_4204);
nor U5394 (N_5394,N_4348,N_4962);
nand U5395 (N_5395,N_4452,N_4751);
xnor U5396 (N_5396,N_4177,N_4395);
or U5397 (N_5397,N_4598,N_4146);
xnor U5398 (N_5398,N_4744,N_4238);
nand U5399 (N_5399,N_4733,N_4597);
nand U5400 (N_5400,N_4881,N_4040);
nor U5401 (N_5401,N_4893,N_4035);
xor U5402 (N_5402,N_4173,N_4963);
xnor U5403 (N_5403,N_4300,N_4916);
xor U5404 (N_5404,N_4834,N_4718);
or U5405 (N_5405,N_4857,N_4563);
and U5406 (N_5406,N_4980,N_4315);
and U5407 (N_5407,N_4616,N_4369);
xnor U5408 (N_5408,N_4066,N_4414);
xor U5409 (N_5409,N_4560,N_4257);
nor U5410 (N_5410,N_4652,N_4678);
and U5411 (N_5411,N_4935,N_4943);
and U5412 (N_5412,N_4875,N_4653);
nand U5413 (N_5413,N_4808,N_4305);
xor U5414 (N_5414,N_4296,N_4010);
or U5415 (N_5415,N_4886,N_4366);
and U5416 (N_5416,N_4576,N_4527);
or U5417 (N_5417,N_4268,N_4961);
or U5418 (N_5418,N_4316,N_4642);
and U5419 (N_5419,N_4607,N_4004);
and U5420 (N_5420,N_4882,N_4908);
nand U5421 (N_5421,N_4230,N_4921);
nand U5422 (N_5422,N_4365,N_4087);
and U5423 (N_5423,N_4979,N_4519);
and U5424 (N_5424,N_4394,N_4029);
nor U5425 (N_5425,N_4707,N_4384);
or U5426 (N_5426,N_4731,N_4175);
nand U5427 (N_5427,N_4640,N_4835);
nor U5428 (N_5428,N_4827,N_4716);
and U5429 (N_5429,N_4552,N_4456);
xnor U5430 (N_5430,N_4682,N_4999);
or U5431 (N_5431,N_4047,N_4482);
or U5432 (N_5432,N_4739,N_4367);
and U5433 (N_5433,N_4540,N_4984);
nor U5434 (N_5434,N_4318,N_4658);
xnor U5435 (N_5435,N_4684,N_4677);
nand U5436 (N_5436,N_4502,N_4253);
or U5437 (N_5437,N_4858,N_4813);
nor U5438 (N_5438,N_4403,N_4700);
or U5439 (N_5439,N_4428,N_4753);
nand U5440 (N_5440,N_4736,N_4031);
and U5441 (N_5441,N_4824,N_4036);
nor U5442 (N_5442,N_4017,N_4681);
xor U5443 (N_5443,N_4831,N_4295);
nand U5444 (N_5444,N_4785,N_4390);
nor U5445 (N_5445,N_4267,N_4621);
xor U5446 (N_5446,N_4187,N_4569);
xor U5447 (N_5447,N_4182,N_4406);
nor U5448 (N_5448,N_4101,N_4960);
nand U5449 (N_5449,N_4409,N_4478);
xor U5450 (N_5450,N_4279,N_4385);
nor U5451 (N_5451,N_4905,N_4584);
nor U5452 (N_5452,N_4577,N_4742);
and U5453 (N_5453,N_4797,N_4966);
nor U5454 (N_5454,N_4455,N_4189);
nor U5455 (N_5455,N_4635,N_4072);
nand U5456 (N_5456,N_4181,N_4802);
nor U5457 (N_5457,N_4038,N_4668);
xor U5458 (N_5458,N_4383,N_4423);
nor U5459 (N_5459,N_4794,N_4111);
and U5460 (N_5460,N_4816,N_4728);
or U5461 (N_5461,N_4096,N_4612);
xor U5462 (N_5462,N_4215,N_4526);
or U5463 (N_5463,N_4500,N_4698);
nand U5464 (N_5464,N_4138,N_4896);
nor U5465 (N_5465,N_4453,N_4258);
nand U5466 (N_5466,N_4322,N_4054);
xor U5467 (N_5467,N_4783,N_4164);
xnor U5468 (N_5468,N_4555,N_4679);
nand U5469 (N_5469,N_4243,N_4109);
nor U5470 (N_5470,N_4771,N_4628);
nand U5471 (N_5471,N_4400,N_4878);
and U5472 (N_5472,N_4381,N_4865);
nand U5473 (N_5473,N_4229,N_4800);
nand U5474 (N_5474,N_4053,N_4037);
and U5475 (N_5475,N_4556,N_4740);
nand U5476 (N_5476,N_4675,N_4459);
xor U5477 (N_5477,N_4462,N_4713);
or U5478 (N_5478,N_4378,N_4127);
nor U5479 (N_5479,N_4449,N_4969);
and U5480 (N_5480,N_4240,N_4473);
or U5481 (N_5481,N_4329,N_4416);
or U5482 (N_5482,N_4407,N_4863);
xor U5483 (N_5483,N_4503,N_4862);
and U5484 (N_5484,N_4755,N_4888);
and U5485 (N_5485,N_4703,N_4470);
or U5486 (N_5486,N_4261,N_4330);
or U5487 (N_5487,N_4754,N_4907);
and U5488 (N_5488,N_4291,N_4493);
and U5489 (N_5489,N_4425,N_4251);
and U5490 (N_5490,N_4202,N_4435);
or U5491 (N_5491,N_4170,N_4647);
nor U5492 (N_5492,N_4055,N_4139);
and U5493 (N_5493,N_4422,N_4080);
nand U5494 (N_5494,N_4374,N_4132);
nor U5495 (N_5495,N_4092,N_4411);
xnor U5496 (N_5496,N_4126,N_4052);
or U5497 (N_5497,N_4118,N_4277);
xor U5498 (N_5498,N_4024,N_4145);
xnor U5499 (N_5499,N_4135,N_4262);
nand U5500 (N_5500,N_4447,N_4972);
nor U5501 (N_5501,N_4683,N_4294);
xor U5502 (N_5502,N_4127,N_4284);
and U5503 (N_5503,N_4898,N_4695);
nand U5504 (N_5504,N_4710,N_4298);
nor U5505 (N_5505,N_4906,N_4690);
and U5506 (N_5506,N_4442,N_4718);
or U5507 (N_5507,N_4367,N_4149);
and U5508 (N_5508,N_4677,N_4853);
xor U5509 (N_5509,N_4100,N_4405);
or U5510 (N_5510,N_4230,N_4975);
xnor U5511 (N_5511,N_4796,N_4797);
nand U5512 (N_5512,N_4962,N_4357);
or U5513 (N_5513,N_4375,N_4086);
and U5514 (N_5514,N_4649,N_4485);
or U5515 (N_5515,N_4348,N_4312);
nor U5516 (N_5516,N_4366,N_4789);
xnor U5517 (N_5517,N_4551,N_4342);
nand U5518 (N_5518,N_4303,N_4427);
and U5519 (N_5519,N_4802,N_4063);
and U5520 (N_5520,N_4230,N_4139);
nor U5521 (N_5521,N_4073,N_4464);
nor U5522 (N_5522,N_4880,N_4767);
and U5523 (N_5523,N_4321,N_4304);
nand U5524 (N_5524,N_4724,N_4651);
and U5525 (N_5525,N_4111,N_4941);
or U5526 (N_5526,N_4533,N_4092);
nand U5527 (N_5527,N_4900,N_4866);
nand U5528 (N_5528,N_4562,N_4633);
nor U5529 (N_5529,N_4623,N_4278);
nand U5530 (N_5530,N_4914,N_4373);
nand U5531 (N_5531,N_4475,N_4012);
nor U5532 (N_5532,N_4963,N_4162);
nor U5533 (N_5533,N_4289,N_4907);
nor U5534 (N_5534,N_4672,N_4765);
nor U5535 (N_5535,N_4826,N_4941);
xnor U5536 (N_5536,N_4054,N_4588);
nor U5537 (N_5537,N_4276,N_4379);
and U5538 (N_5538,N_4266,N_4220);
nand U5539 (N_5539,N_4905,N_4966);
nand U5540 (N_5540,N_4573,N_4614);
nor U5541 (N_5541,N_4093,N_4858);
or U5542 (N_5542,N_4828,N_4870);
xor U5543 (N_5543,N_4125,N_4771);
nor U5544 (N_5544,N_4980,N_4510);
or U5545 (N_5545,N_4920,N_4839);
xnor U5546 (N_5546,N_4595,N_4753);
xnor U5547 (N_5547,N_4555,N_4254);
and U5548 (N_5548,N_4634,N_4849);
nor U5549 (N_5549,N_4115,N_4003);
xnor U5550 (N_5550,N_4571,N_4453);
nand U5551 (N_5551,N_4339,N_4566);
or U5552 (N_5552,N_4459,N_4749);
or U5553 (N_5553,N_4482,N_4511);
or U5554 (N_5554,N_4682,N_4146);
nand U5555 (N_5555,N_4377,N_4357);
and U5556 (N_5556,N_4449,N_4207);
nand U5557 (N_5557,N_4502,N_4079);
xor U5558 (N_5558,N_4154,N_4572);
nand U5559 (N_5559,N_4477,N_4614);
and U5560 (N_5560,N_4467,N_4023);
xnor U5561 (N_5561,N_4160,N_4054);
nand U5562 (N_5562,N_4415,N_4487);
nor U5563 (N_5563,N_4992,N_4545);
nor U5564 (N_5564,N_4593,N_4320);
or U5565 (N_5565,N_4898,N_4837);
nand U5566 (N_5566,N_4740,N_4728);
nand U5567 (N_5567,N_4967,N_4452);
nand U5568 (N_5568,N_4512,N_4317);
nand U5569 (N_5569,N_4287,N_4546);
and U5570 (N_5570,N_4970,N_4499);
nand U5571 (N_5571,N_4574,N_4729);
and U5572 (N_5572,N_4927,N_4348);
or U5573 (N_5573,N_4185,N_4446);
xor U5574 (N_5574,N_4329,N_4498);
nand U5575 (N_5575,N_4869,N_4238);
xor U5576 (N_5576,N_4019,N_4198);
and U5577 (N_5577,N_4671,N_4307);
nand U5578 (N_5578,N_4481,N_4546);
and U5579 (N_5579,N_4765,N_4307);
and U5580 (N_5580,N_4124,N_4083);
or U5581 (N_5581,N_4475,N_4960);
xor U5582 (N_5582,N_4388,N_4835);
and U5583 (N_5583,N_4041,N_4668);
and U5584 (N_5584,N_4526,N_4033);
nor U5585 (N_5585,N_4322,N_4101);
xor U5586 (N_5586,N_4759,N_4870);
nand U5587 (N_5587,N_4549,N_4884);
nand U5588 (N_5588,N_4387,N_4549);
nand U5589 (N_5589,N_4948,N_4028);
or U5590 (N_5590,N_4871,N_4642);
nor U5591 (N_5591,N_4212,N_4948);
nor U5592 (N_5592,N_4966,N_4027);
nor U5593 (N_5593,N_4977,N_4752);
xnor U5594 (N_5594,N_4868,N_4680);
or U5595 (N_5595,N_4861,N_4375);
or U5596 (N_5596,N_4576,N_4423);
xor U5597 (N_5597,N_4957,N_4671);
nor U5598 (N_5598,N_4756,N_4280);
nand U5599 (N_5599,N_4154,N_4071);
nand U5600 (N_5600,N_4906,N_4904);
and U5601 (N_5601,N_4615,N_4484);
or U5602 (N_5602,N_4764,N_4487);
or U5603 (N_5603,N_4829,N_4320);
or U5604 (N_5604,N_4368,N_4453);
xnor U5605 (N_5605,N_4768,N_4825);
and U5606 (N_5606,N_4305,N_4228);
and U5607 (N_5607,N_4719,N_4854);
and U5608 (N_5608,N_4341,N_4008);
or U5609 (N_5609,N_4262,N_4355);
nand U5610 (N_5610,N_4235,N_4556);
nor U5611 (N_5611,N_4171,N_4393);
xor U5612 (N_5612,N_4214,N_4476);
or U5613 (N_5613,N_4731,N_4375);
nor U5614 (N_5614,N_4835,N_4367);
xor U5615 (N_5615,N_4912,N_4103);
or U5616 (N_5616,N_4434,N_4762);
nor U5617 (N_5617,N_4483,N_4928);
or U5618 (N_5618,N_4733,N_4809);
and U5619 (N_5619,N_4038,N_4343);
and U5620 (N_5620,N_4775,N_4123);
nand U5621 (N_5621,N_4083,N_4610);
nor U5622 (N_5622,N_4727,N_4234);
and U5623 (N_5623,N_4275,N_4624);
and U5624 (N_5624,N_4643,N_4085);
nor U5625 (N_5625,N_4633,N_4354);
xor U5626 (N_5626,N_4148,N_4512);
or U5627 (N_5627,N_4366,N_4807);
xor U5628 (N_5628,N_4072,N_4100);
and U5629 (N_5629,N_4476,N_4165);
and U5630 (N_5630,N_4607,N_4615);
xor U5631 (N_5631,N_4890,N_4972);
xor U5632 (N_5632,N_4219,N_4263);
nor U5633 (N_5633,N_4108,N_4365);
xnor U5634 (N_5634,N_4067,N_4651);
nand U5635 (N_5635,N_4373,N_4295);
nand U5636 (N_5636,N_4237,N_4610);
nor U5637 (N_5637,N_4071,N_4963);
nor U5638 (N_5638,N_4029,N_4812);
or U5639 (N_5639,N_4847,N_4863);
xor U5640 (N_5640,N_4864,N_4253);
and U5641 (N_5641,N_4607,N_4651);
xor U5642 (N_5642,N_4968,N_4376);
and U5643 (N_5643,N_4715,N_4660);
nor U5644 (N_5644,N_4361,N_4120);
nand U5645 (N_5645,N_4304,N_4223);
and U5646 (N_5646,N_4914,N_4100);
xnor U5647 (N_5647,N_4670,N_4204);
xor U5648 (N_5648,N_4465,N_4790);
and U5649 (N_5649,N_4359,N_4155);
nor U5650 (N_5650,N_4609,N_4773);
nand U5651 (N_5651,N_4074,N_4066);
nor U5652 (N_5652,N_4844,N_4065);
or U5653 (N_5653,N_4505,N_4629);
nand U5654 (N_5654,N_4312,N_4462);
and U5655 (N_5655,N_4846,N_4571);
or U5656 (N_5656,N_4890,N_4929);
xnor U5657 (N_5657,N_4957,N_4539);
nor U5658 (N_5658,N_4514,N_4259);
nor U5659 (N_5659,N_4584,N_4598);
nor U5660 (N_5660,N_4877,N_4479);
xor U5661 (N_5661,N_4170,N_4840);
or U5662 (N_5662,N_4963,N_4606);
nand U5663 (N_5663,N_4093,N_4961);
nor U5664 (N_5664,N_4615,N_4529);
and U5665 (N_5665,N_4901,N_4743);
nor U5666 (N_5666,N_4466,N_4856);
nand U5667 (N_5667,N_4159,N_4708);
or U5668 (N_5668,N_4720,N_4945);
xnor U5669 (N_5669,N_4891,N_4651);
and U5670 (N_5670,N_4259,N_4318);
or U5671 (N_5671,N_4622,N_4258);
or U5672 (N_5672,N_4017,N_4224);
or U5673 (N_5673,N_4591,N_4430);
nand U5674 (N_5674,N_4431,N_4594);
or U5675 (N_5675,N_4583,N_4837);
nor U5676 (N_5676,N_4071,N_4852);
nor U5677 (N_5677,N_4441,N_4516);
and U5678 (N_5678,N_4504,N_4449);
nand U5679 (N_5679,N_4158,N_4149);
xor U5680 (N_5680,N_4925,N_4783);
nor U5681 (N_5681,N_4127,N_4717);
nand U5682 (N_5682,N_4973,N_4816);
xor U5683 (N_5683,N_4098,N_4763);
nand U5684 (N_5684,N_4546,N_4730);
and U5685 (N_5685,N_4374,N_4378);
and U5686 (N_5686,N_4787,N_4215);
nor U5687 (N_5687,N_4655,N_4454);
nand U5688 (N_5688,N_4657,N_4231);
nand U5689 (N_5689,N_4624,N_4773);
xnor U5690 (N_5690,N_4316,N_4345);
nor U5691 (N_5691,N_4707,N_4277);
or U5692 (N_5692,N_4153,N_4728);
or U5693 (N_5693,N_4656,N_4455);
and U5694 (N_5694,N_4733,N_4532);
and U5695 (N_5695,N_4005,N_4321);
xnor U5696 (N_5696,N_4761,N_4092);
nor U5697 (N_5697,N_4924,N_4370);
and U5698 (N_5698,N_4469,N_4350);
and U5699 (N_5699,N_4047,N_4261);
or U5700 (N_5700,N_4985,N_4685);
and U5701 (N_5701,N_4753,N_4742);
nand U5702 (N_5702,N_4853,N_4666);
xnor U5703 (N_5703,N_4732,N_4998);
xor U5704 (N_5704,N_4969,N_4745);
and U5705 (N_5705,N_4420,N_4257);
or U5706 (N_5706,N_4130,N_4605);
nor U5707 (N_5707,N_4314,N_4979);
nand U5708 (N_5708,N_4600,N_4768);
and U5709 (N_5709,N_4024,N_4079);
or U5710 (N_5710,N_4422,N_4301);
and U5711 (N_5711,N_4419,N_4815);
or U5712 (N_5712,N_4203,N_4812);
xnor U5713 (N_5713,N_4484,N_4945);
nor U5714 (N_5714,N_4593,N_4718);
or U5715 (N_5715,N_4409,N_4018);
nand U5716 (N_5716,N_4110,N_4475);
nand U5717 (N_5717,N_4690,N_4633);
nand U5718 (N_5718,N_4154,N_4374);
xor U5719 (N_5719,N_4956,N_4451);
and U5720 (N_5720,N_4344,N_4543);
and U5721 (N_5721,N_4262,N_4580);
or U5722 (N_5722,N_4013,N_4864);
or U5723 (N_5723,N_4273,N_4861);
xnor U5724 (N_5724,N_4615,N_4710);
nor U5725 (N_5725,N_4179,N_4124);
and U5726 (N_5726,N_4791,N_4360);
nand U5727 (N_5727,N_4105,N_4230);
or U5728 (N_5728,N_4224,N_4100);
nor U5729 (N_5729,N_4927,N_4694);
or U5730 (N_5730,N_4979,N_4044);
nor U5731 (N_5731,N_4808,N_4408);
nor U5732 (N_5732,N_4996,N_4934);
nand U5733 (N_5733,N_4855,N_4394);
or U5734 (N_5734,N_4207,N_4342);
or U5735 (N_5735,N_4355,N_4231);
nor U5736 (N_5736,N_4280,N_4022);
or U5737 (N_5737,N_4660,N_4397);
or U5738 (N_5738,N_4862,N_4878);
and U5739 (N_5739,N_4884,N_4936);
and U5740 (N_5740,N_4117,N_4023);
nand U5741 (N_5741,N_4216,N_4903);
or U5742 (N_5742,N_4481,N_4537);
and U5743 (N_5743,N_4358,N_4810);
nor U5744 (N_5744,N_4404,N_4324);
nor U5745 (N_5745,N_4013,N_4862);
or U5746 (N_5746,N_4462,N_4489);
xnor U5747 (N_5747,N_4244,N_4275);
nor U5748 (N_5748,N_4791,N_4180);
and U5749 (N_5749,N_4230,N_4074);
and U5750 (N_5750,N_4363,N_4302);
and U5751 (N_5751,N_4838,N_4154);
or U5752 (N_5752,N_4931,N_4529);
nand U5753 (N_5753,N_4494,N_4865);
and U5754 (N_5754,N_4620,N_4493);
nor U5755 (N_5755,N_4766,N_4143);
nand U5756 (N_5756,N_4969,N_4886);
nor U5757 (N_5757,N_4646,N_4906);
nor U5758 (N_5758,N_4885,N_4679);
or U5759 (N_5759,N_4574,N_4091);
nor U5760 (N_5760,N_4966,N_4798);
or U5761 (N_5761,N_4083,N_4931);
nand U5762 (N_5762,N_4372,N_4344);
and U5763 (N_5763,N_4291,N_4043);
nor U5764 (N_5764,N_4809,N_4121);
and U5765 (N_5765,N_4955,N_4146);
or U5766 (N_5766,N_4927,N_4325);
and U5767 (N_5767,N_4685,N_4214);
nor U5768 (N_5768,N_4050,N_4485);
xnor U5769 (N_5769,N_4284,N_4412);
and U5770 (N_5770,N_4717,N_4227);
nand U5771 (N_5771,N_4398,N_4910);
xnor U5772 (N_5772,N_4951,N_4671);
xnor U5773 (N_5773,N_4773,N_4170);
nor U5774 (N_5774,N_4401,N_4879);
or U5775 (N_5775,N_4734,N_4554);
xnor U5776 (N_5776,N_4001,N_4955);
nor U5777 (N_5777,N_4290,N_4836);
xor U5778 (N_5778,N_4739,N_4692);
and U5779 (N_5779,N_4775,N_4604);
nand U5780 (N_5780,N_4446,N_4019);
nor U5781 (N_5781,N_4458,N_4474);
nor U5782 (N_5782,N_4767,N_4966);
or U5783 (N_5783,N_4708,N_4682);
nand U5784 (N_5784,N_4320,N_4739);
xor U5785 (N_5785,N_4144,N_4150);
or U5786 (N_5786,N_4470,N_4214);
xnor U5787 (N_5787,N_4437,N_4133);
xnor U5788 (N_5788,N_4462,N_4997);
nand U5789 (N_5789,N_4152,N_4399);
or U5790 (N_5790,N_4087,N_4456);
nor U5791 (N_5791,N_4939,N_4372);
xnor U5792 (N_5792,N_4744,N_4615);
nor U5793 (N_5793,N_4173,N_4311);
or U5794 (N_5794,N_4279,N_4817);
nor U5795 (N_5795,N_4331,N_4150);
and U5796 (N_5796,N_4893,N_4415);
nand U5797 (N_5797,N_4055,N_4622);
xnor U5798 (N_5798,N_4152,N_4180);
nand U5799 (N_5799,N_4561,N_4736);
nand U5800 (N_5800,N_4687,N_4150);
and U5801 (N_5801,N_4204,N_4329);
or U5802 (N_5802,N_4712,N_4025);
or U5803 (N_5803,N_4389,N_4545);
nand U5804 (N_5804,N_4791,N_4022);
and U5805 (N_5805,N_4439,N_4729);
and U5806 (N_5806,N_4996,N_4225);
or U5807 (N_5807,N_4143,N_4884);
nand U5808 (N_5808,N_4397,N_4568);
xnor U5809 (N_5809,N_4390,N_4541);
and U5810 (N_5810,N_4241,N_4966);
nor U5811 (N_5811,N_4526,N_4179);
xnor U5812 (N_5812,N_4880,N_4637);
and U5813 (N_5813,N_4645,N_4578);
xnor U5814 (N_5814,N_4461,N_4382);
nor U5815 (N_5815,N_4002,N_4629);
nor U5816 (N_5816,N_4388,N_4579);
or U5817 (N_5817,N_4412,N_4061);
xnor U5818 (N_5818,N_4108,N_4637);
and U5819 (N_5819,N_4178,N_4542);
nand U5820 (N_5820,N_4355,N_4994);
or U5821 (N_5821,N_4697,N_4400);
xnor U5822 (N_5822,N_4128,N_4676);
nand U5823 (N_5823,N_4853,N_4250);
nand U5824 (N_5824,N_4874,N_4557);
nand U5825 (N_5825,N_4992,N_4516);
nor U5826 (N_5826,N_4133,N_4743);
nor U5827 (N_5827,N_4912,N_4033);
and U5828 (N_5828,N_4139,N_4069);
or U5829 (N_5829,N_4678,N_4664);
xor U5830 (N_5830,N_4443,N_4961);
nand U5831 (N_5831,N_4362,N_4466);
or U5832 (N_5832,N_4452,N_4697);
or U5833 (N_5833,N_4514,N_4606);
and U5834 (N_5834,N_4956,N_4861);
nand U5835 (N_5835,N_4892,N_4272);
nor U5836 (N_5836,N_4518,N_4194);
and U5837 (N_5837,N_4787,N_4119);
and U5838 (N_5838,N_4415,N_4889);
xnor U5839 (N_5839,N_4022,N_4478);
and U5840 (N_5840,N_4450,N_4875);
nand U5841 (N_5841,N_4281,N_4674);
nand U5842 (N_5842,N_4789,N_4146);
and U5843 (N_5843,N_4960,N_4829);
xnor U5844 (N_5844,N_4355,N_4945);
and U5845 (N_5845,N_4793,N_4198);
nor U5846 (N_5846,N_4122,N_4232);
and U5847 (N_5847,N_4873,N_4439);
xor U5848 (N_5848,N_4493,N_4361);
and U5849 (N_5849,N_4518,N_4763);
xnor U5850 (N_5850,N_4443,N_4279);
xor U5851 (N_5851,N_4169,N_4761);
xnor U5852 (N_5852,N_4117,N_4391);
xor U5853 (N_5853,N_4248,N_4829);
or U5854 (N_5854,N_4767,N_4459);
or U5855 (N_5855,N_4529,N_4135);
or U5856 (N_5856,N_4906,N_4870);
and U5857 (N_5857,N_4714,N_4831);
xnor U5858 (N_5858,N_4036,N_4198);
nor U5859 (N_5859,N_4960,N_4590);
or U5860 (N_5860,N_4323,N_4301);
nor U5861 (N_5861,N_4568,N_4025);
nand U5862 (N_5862,N_4620,N_4051);
nand U5863 (N_5863,N_4654,N_4940);
nor U5864 (N_5864,N_4535,N_4381);
and U5865 (N_5865,N_4811,N_4788);
or U5866 (N_5866,N_4970,N_4117);
or U5867 (N_5867,N_4039,N_4634);
and U5868 (N_5868,N_4438,N_4903);
xor U5869 (N_5869,N_4319,N_4115);
and U5870 (N_5870,N_4681,N_4542);
or U5871 (N_5871,N_4495,N_4240);
xor U5872 (N_5872,N_4228,N_4366);
nor U5873 (N_5873,N_4580,N_4215);
or U5874 (N_5874,N_4557,N_4961);
or U5875 (N_5875,N_4193,N_4841);
xor U5876 (N_5876,N_4411,N_4864);
nor U5877 (N_5877,N_4558,N_4704);
or U5878 (N_5878,N_4866,N_4822);
nor U5879 (N_5879,N_4203,N_4590);
nand U5880 (N_5880,N_4782,N_4495);
nor U5881 (N_5881,N_4884,N_4359);
xor U5882 (N_5882,N_4412,N_4358);
nor U5883 (N_5883,N_4958,N_4943);
or U5884 (N_5884,N_4174,N_4989);
and U5885 (N_5885,N_4611,N_4404);
nand U5886 (N_5886,N_4859,N_4080);
xor U5887 (N_5887,N_4410,N_4626);
nor U5888 (N_5888,N_4359,N_4041);
or U5889 (N_5889,N_4550,N_4345);
xnor U5890 (N_5890,N_4235,N_4566);
xnor U5891 (N_5891,N_4706,N_4087);
or U5892 (N_5892,N_4048,N_4459);
and U5893 (N_5893,N_4750,N_4222);
xor U5894 (N_5894,N_4014,N_4944);
nand U5895 (N_5895,N_4218,N_4939);
xnor U5896 (N_5896,N_4551,N_4169);
nor U5897 (N_5897,N_4143,N_4987);
nand U5898 (N_5898,N_4359,N_4181);
xor U5899 (N_5899,N_4694,N_4349);
or U5900 (N_5900,N_4186,N_4348);
or U5901 (N_5901,N_4306,N_4668);
xor U5902 (N_5902,N_4086,N_4461);
xnor U5903 (N_5903,N_4033,N_4916);
and U5904 (N_5904,N_4008,N_4989);
nand U5905 (N_5905,N_4679,N_4084);
nor U5906 (N_5906,N_4502,N_4561);
nand U5907 (N_5907,N_4558,N_4038);
xor U5908 (N_5908,N_4423,N_4732);
xnor U5909 (N_5909,N_4495,N_4009);
or U5910 (N_5910,N_4233,N_4237);
or U5911 (N_5911,N_4767,N_4406);
nand U5912 (N_5912,N_4449,N_4188);
xnor U5913 (N_5913,N_4872,N_4336);
or U5914 (N_5914,N_4185,N_4030);
and U5915 (N_5915,N_4267,N_4504);
nand U5916 (N_5916,N_4931,N_4162);
and U5917 (N_5917,N_4441,N_4675);
or U5918 (N_5918,N_4927,N_4188);
xnor U5919 (N_5919,N_4001,N_4770);
or U5920 (N_5920,N_4356,N_4200);
nand U5921 (N_5921,N_4487,N_4167);
or U5922 (N_5922,N_4239,N_4885);
and U5923 (N_5923,N_4738,N_4838);
nor U5924 (N_5924,N_4966,N_4984);
and U5925 (N_5925,N_4186,N_4388);
xor U5926 (N_5926,N_4840,N_4414);
xnor U5927 (N_5927,N_4014,N_4980);
nor U5928 (N_5928,N_4018,N_4474);
nor U5929 (N_5929,N_4240,N_4823);
xor U5930 (N_5930,N_4587,N_4554);
and U5931 (N_5931,N_4790,N_4536);
or U5932 (N_5932,N_4580,N_4826);
xor U5933 (N_5933,N_4148,N_4333);
and U5934 (N_5934,N_4138,N_4934);
nand U5935 (N_5935,N_4239,N_4904);
and U5936 (N_5936,N_4667,N_4192);
and U5937 (N_5937,N_4790,N_4312);
xnor U5938 (N_5938,N_4528,N_4984);
nor U5939 (N_5939,N_4390,N_4537);
or U5940 (N_5940,N_4973,N_4964);
or U5941 (N_5941,N_4056,N_4069);
nand U5942 (N_5942,N_4202,N_4077);
xor U5943 (N_5943,N_4629,N_4023);
xnor U5944 (N_5944,N_4077,N_4568);
and U5945 (N_5945,N_4661,N_4174);
nand U5946 (N_5946,N_4039,N_4917);
or U5947 (N_5947,N_4313,N_4309);
xnor U5948 (N_5948,N_4062,N_4506);
or U5949 (N_5949,N_4683,N_4896);
nand U5950 (N_5950,N_4674,N_4442);
or U5951 (N_5951,N_4100,N_4713);
nand U5952 (N_5952,N_4396,N_4871);
nand U5953 (N_5953,N_4528,N_4841);
or U5954 (N_5954,N_4016,N_4806);
xor U5955 (N_5955,N_4866,N_4196);
nor U5956 (N_5956,N_4186,N_4743);
xnor U5957 (N_5957,N_4599,N_4520);
nand U5958 (N_5958,N_4552,N_4492);
nor U5959 (N_5959,N_4257,N_4553);
nand U5960 (N_5960,N_4682,N_4961);
and U5961 (N_5961,N_4489,N_4728);
nand U5962 (N_5962,N_4123,N_4481);
or U5963 (N_5963,N_4102,N_4144);
xor U5964 (N_5964,N_4795,N_4886);
nand U5965 (N_5965,N_4612,N_4033);
nand U5966 (N_5966,N_4423,N_4901);
and U5967 (N_5967,N_4936,N_4477);
or U5968 (N_5968,N_4100,N_4729);
or U5969 (N_5969,N_4258,N_4176);
and U5970 (N_5970,N_4095,N_4818);
or U5971 (N_5971,N_4104,N_4515);
nand U5972 (N_5972,N_4568,N_4772);
nor U5973 (N_5973,N_4977,N_4201);
and U5974 (N_5974,N_4281,N_4015);
xor U5975 (N_5975,N_4469,N_4942);
nand U5976 (N_5976,N_4902,N_4631);
xnor U5977 (N_5977,N_4913,N_4576);
nand U5978 (N_5978,N_4698,N_4003);
nor U5979 (N_5979,N_4907,N_4958);
nor U5980 (N_5980,N_4087,N_4280);
xor U5981 (N_5981,N_4219,N_4972);
nand U5982 (N_5982,N_4710,N_4224);
or U5983 (N_5983,N_4129,N_4658);
nor U5984 (N_5984,N_4244,N_4320);
and U5985 (N_5985,N_4290,N_4663);
xor U5986 (N_5986,N_4602,N_4320);
nor U5987 (N_5987,N_4292,N_4286);
nor U5988 (N_5988,N_4368,N_4747);
nand U5989 (N_5989,N_4860,N_4536);
and U5990 (N_5990,N_4559,N_4860);
xnor U5991 (N_5991,N_4369,N_4249);
xor U5992 (N_5992,N_4257,N_4648);
and U5993 (N_5993,N_4143,N_4900);
nor U5994 (N_5994,N_4192,N_4002);
or U5995 (N_5995,N_4080,N_4160);
or U5996 (N_5996,N_4182,N_4135);
and U5997 (N_5997,N_4312,N_4051);
nor U5998 (N_5998,N_4859,N_4781);
or U5999 (N_5999,N_4966,N_4265);
or U6000 (N_6000,N_5874,N_5750);
and U6001 (N_6001,N_5703,N_5018);
nor U6002 (N_6002,N_5841,N_5479);
nand U6003 (N_6003,N_5572,N_5986);
or U6004 (N_6004,N_5324,N_5711);
xor U6005 (N_6005,N_5641,N_5893);
or U6006 (N_6006,N_5152,N_5632);
and U6007 (N_6007,N_5737,N_5700);
nand U6008 (N_6008,N_5755,N_5735);
and U6009 (N_6009,N_5752,N_5513);
or U6010 (N_6010,N_5283,N_5395);
or U6011 (N_6011,N_5399,N_5655);
nor U6012 (N_6012,N_5690,N_5445);
nor U6013 (N_6013,N_5944,N_5681);
or U6014 (N_6014,N_5454,N_5758);
or U6015 (N_6015,N_5771,N_5914);
nor U6016 (N_6016,N_5719,N_5340);
or U6017 (N_6017,N_5618,N_5665);
nor U6018 (N_6018,N_5895,N_5963);
xnor U6019 (N_6019,N_5877,N_5140);
and U6020 (N_6020,N_5002,N_5535);
nand U6021 (N_6021,N_5346,N_5834);
or U6022 (N_6022,N_5991,N_5166);
xor U6023 (N_6023,N_5011,N_5226);
nor U6024 (N_6024,N_5858,N_5325);
and U6025 (N_6025,N_5113,N_5886);
and U6026 (N_6026,N_5006,N_5142);
xnor U6027 (N_6027,N_5805,N_5542);
and U6028 (N_6028,N_5687,N_5987);
and U6029 (N_6029,N_5724,N_5713);
and U6030 (N_6030,N_5281,N_5407);
and U6031 (N_6031,N_5129,N_5249);
nor U6032 (N_6032,N_5382,N_5459);
xnor U6033 (N_6033,N_5205,N_5613);
xnor U6034 (N_6034,N_5231,N_5876);
and U6035 (N_6035,N_5087,N_5617);
and U6036 (N_6036,N_5585,N_5107);
nor U6037 (N_6037,N_5736,N_5322);
nand U6038 (N_6038,N_5334,N_5278);
and U6039 (N_6039,N_5526,N_5929);
or U6040 (N_6040,N_5518,N_5562);
and U6041 (N_6041,N_5491,N_5507);
nor U6042 (N_6042,N_5162,N_5483);
or U6043 (N_6043,N_5500,N_5159);
xor U6044 (N_6044,N_5994,N_5754);
or U6045 (N_6045,N_5300,N_5235);
xnor U6046 (N_6046,N_5461,N_5345);
or U6047 (N_6047,N_5765,N_5280);
or U6048 (N_6048,N_5000,N_5748);
nor U6049 (N_6049,N_5026,N_5447);
xnor U6050 (N_6050,N_5998,N_5635);
and U6051 (N_6051,N_5849,N_5309);
or U6052 (N_6052,N_5191,N_5381);
and U6053 (N_6053,N_5882,N_5509);
nor U6054 (N_6054,N_5552,N_5151);
xnor U6055 (N_6055,N_5145,N_5534);
xor U6056 (N_6056,N_5287,N_5845);
nor U6057 (N_6057,N_5361,N_5153);
nor U6058 (N_6058,N_5359,N_5085);
nor U6059 (N_6059,N_5127,N_5707);
nor U6060 (N_6060,N_5599,N_5606);
xor U6061 (N_6061,N_5063,N_5715);
or U6062 (N_6062,N_5316,N_5331);
nor U6063 (N_6063,N_5260,N_5842);
nand U6064 (N_6064,N_5699,N_5517);
xnor U6065 (N_6065,N_5462,N_5385);
xnor U6066 (N_6066,N_5695,N_5326);
or U6067 (N_6067,N_5293,N_5716);
nand U6068 (N_6068,N_5939,N_5012);
nor U6069 (N_6069,N_5588,N_5933);
nand U6070 (N_6070,N_5993,N_5243);
xnor U6071 (N_6071,N_5527,N_5441);
and U6072 (N_6072,N_5015,N_5852);
or U6073 (N_6073,N_5157,N_5123);
and U6074 (N_6074,N_5496,N_5712);
xnor U6075 (N_6075,N_5003,N_5192);
or U6076 (N_6076,N_5060,N_5439);
or U6077 (N_6077,N_5682,N_5451);
nand U6078 (N_6078,N_5823,N_5136);
nand U6079 (N_6079,N_5443,N_5938);
and U6080 (N_6080,N_5753,N_5953);
xnor U6081 (N_6081,N_5756,N_5387);
xnor U6082 (N_6082,N_5955,N_5071);
and U6083 (N_6083,N_5729,N_5868);
nand U6084 (N_6084,N_5614,N_5415);
or U6085 (N_6085,N_5220,N_5821);
or U6086 (N_6086,N_5409,N_5052);
or U6087 (N_6087,N_5918,N_5551);
nor U6088 (N_6088,N_5651,N_5775);
or U6089 (N_6089,N_5110,N_5265);
xor U6090 (N_6090,N_5652,N_5024);
nor U6091 (N_6091,N_5592,N_5802);
and U6092 (N_6092,N_5383,N_5266);
xor U6093 (N_6093,N_5034,N_5025);
or U6094 (N_6094,N_5314,N_5400);
nand U6095 (N_6095,N_5117,N_5471);
nand U6096 (N_6096,N_5571,N_5298);
and U6097 (N_6097,N_5574,N_5485);
and U6098 (N_6098,N_5568,N_5165);
or U6099 (N_6099,N_5369,N_5610);
and U6100 (N_6100,N_5899,N_5785);
nand U6101 (N_6101,N_5384,N_5807);
nand U6102 (N_6102,N_5320,N_5596);
and U6103 (N_6103,N_5290,N_5550);
nand U6104 (N_6104,N_5629,N_5777);
nand U6105 (N_6105,N_5636,N_5639);
or U6106 (N_6106,N_5952,N_5591);
nand U6107 (N_6107,N_5154,N_5965);
nor U6108 (N_6108,N_5187,N_5795);
or U6109 (N_6109,N_5520,N_5839);
and U6110 (N_6110,N_5229,N_5351);
nor U6111 (N_6111,N_5814,N_5161);
and U6112 (N_6112,N_5059,N_5313);
nand U6113 (N_6113,N_5945,N_5554);
and U6114 (N_6114,N_5648,N_5553);
and U6115 (N_6115,N_5227,N_5837);
or U6116 (N_6116,N_5259,N_5956);
and U6117 (N_6117,N_5124,N_5198);
or U6118 (N_6118,N_5630,N_5913);
or U6119 (N_6119,N_5078,N_5565);
nand U6120 (N_6120,N_5048,N_5444);
xor U6121 (N_6121,N_5075,N_5718);
nor U6122 (N_6122,N_5657,N_5464);
or U6123 (N_6123,N_5446,N_5722);
or U6124 (N_6124,N_5150,N_5267);
nor U6125 (N_6125,N_5867,N_5790);
nor U6126 (N_6126,N_5363,N_5809);
nand U6127 (N_6127,N_5989,N_5423);
nor U6128 (N_6128,N_5883,N_5065);
xnor U6129 (N_6129,N_5905,N_5533);
and U6130 (N_6130,N_5578,N_5970);
xnor U6131 (N_6131,N_5607,N_5625);
nor U6132 (N_6132,N_5547,N_5094);
xnor U6133 (N_6133,N_5277,N_5402);
or U6134 (N_6134,N_5672,N_5693);
and U6135 (N_6135,N_5698,N_5437);
or U6136 (N_6136,N_5335,N_5926);
or U6137 (N_6137,N_5723,N_5850);
and U6138 (N_6138,N_5307,N_5296);
xor U6139 (N_6139,N_5642,N_5621);
nand U6140 (N_6140,N_5431,N_5244);
nand U6141 (N_6141,N_5132,N_5812);
xnor U6142 (N_6142,N_5808,N_5274);
nor U6143 (N_6143,N_5264,N_5769);
nand U6144 (N_6144,N_5594,N_5194);
nor U6145 (N_6145,N_5028,N_5149);
nor U6146 (N_6146,N_5178,N_5356);
nand U6147 (N_6147,N_5119,N_5138);
xor U6148 (N_6148,N_5321,N_5019);
and U6149 (N_6149,N_5806,N_5438);
nand U6150 (N_6150,N_5996,N_5484);
and U6151 (N_6151,N_5257,N_5872);
nand U6152 (N_6152,N_5680,N_5469);
or U6153 (N_6153,N_5671,N_5115);
xnor U6154 (N_6154,N_5661,N_5948);
and U6155 (N_6155,N_5640,N_5694);
nor U6156 (N_6156,N_5378,N_5846);
nand U6157 (N_6157,N_5584,N_5337);
nand U6158 (N_6158,N_5401,N_5966);
or U6159 (N_6159,N_5920,N_5362);
nand U6160 (N_6160,N_5083,N_5559);
nor U6161 (N_6161,N_5389,N_5819);
or U6162 (N_6162,N_5541,N_5426);
or U6163 (N_6163,N_5549,N_5336);
xnor U6164 (N_6164,N_5961,N_5408);
xor U6165 (N_6165,N_5066,N_5794);
nand U6166 (N_6166,N_5263,N_5902);
or U6167 (N_6167,N_5077,N_5386);
or U6168 (N_6168,N_5091,N_5792);
nor U6169 (N_6169,N_5105,N_5366);
nor U6170 (N_6170,N_5580,N_5420);
nor U6171 (N_6171,N_5310,N_5367);
xor U6172 (N_6172,N_5251,N_5788);
or U6173 (N_6173,N_5312,N_5167);
nand U6174 (N_6174,N_5116,N_5885);
nor U6175 (N_6175,N_5631,N_5076);
xnor U6176 (N_6176,N_5204,N_5398);
nor U6177 (N_6177,N_5793,N_5360);
xor U6178 (N_6178,N_5619,N_5772);
nor U6179 (N_6179,N_5761,N_5583);
nand U6180 (N_6180,N_5811,N_5728);
or U6181 (N_6181,N_5530,N_5173);
or U6182 (N_6182,N_5742,N_5995);
or U6183 (N_6183,N_5637,N_5947);
or U6184 (N_6184,N_5611,N_5764);
and U6185 (N_6185,N_5044,N_5328);
nor U6186 (N_6186,N_5977,N_5181);
and U6187 (N_6187,N_5228,N_5089);
or U6188 (N_6188,N_5787,N_5416);
xnor U6189 (N_6189,N_5391,N_5412);
xor U6190 (N_6190,N_5531,N_5179);
or U6191 (N_6191,N_5211,N_5815);
nor U6192 (N_6192,N_5058,N_5714);
nor U6193 (N_6193,N_5350,N_5847);
or U6194 (N_6194,N_5813,N_5176);
nor U6195 (N_6195,N_5037,N_5759);
xor U6196 (N_6196,N_5333,N_5009);
xor U6197 (N_6197,N_5394,N_5061);
nor U6198 (N_6198,N_5158,N_5906);
or U6199 (N_6199,N_5200,N_5062);
or U6200 (N_6200,N_5799,N_5236);
and U6201 (N_6201,N_5050,N_5212);
nor U6202 (N_6202,N_5308,N_5358);
xnor U6203 (N_6203,N_5909,N_5141);
and U6204 (N_6204,N_5907,N_5352);
xor U6205 (N_6205,N_5282,N_5543);
or U6206 (N_6206,N_5894,N_5174);
or U6207 (N_6207,N_5099,N_5419);
nand U6208 (N_6208,N_5840,N_5143);
nor U6209 (N_6209,N_5064,N_5701);
and U6210 (N_6210,N_5999,N_5983);
or U6211 (N_6211,N_5988,N_5820);
nor U6212 (N_6212,N_5576,N_5673);
xor U6213 (N_6213,N_5207,N_5074);
or U6214 (N_6214,N_5563,N_5931);
nand U6215 (N_6215,N_5573,N_5798);
and U6216 (N_6216,N_5878,N_5873);
or U6217 (N_6217,N_5896,N_5021);
and U6218 (N_6218,N_5031,N_5744);
or U6219 (N_6219,N_5195,N_5271);
nor U6220 (N_6220,N_5555,N_5747);
nand U6221 (N_6221,N_5692,N_5767);
nand U6222 (N_6222,N_5467,N_5684);
and U6223 (N_6223,N_5344,N_5403);
or U6224 (N_6224,N_5008,N_5967);
xnor U6225 (N_6225,N_5460,N_5010);
and U6226 (N_6226,N_5406,N_5088);
nor U6227 (N_6227,N_5688,N_5303);
xor U6228 (N_6228,N_5486,N_5916);
nor U6229 (N_6229,N_5863,N_5968);
nand U6230 (N_6230,N_5349,N_5348);
nor U6231 (N_6231,N_5473,N_5388);
nor U6232 (N_6232,N_5442,N_5848);
and U6233 (N_6233,N_5668,N_5193);
nor U6234 (N_6234,N_5502,N_5739);
or U6235 (N_6235,N_5940,N_5217);
nand U6236 (N_6236,N_5273,N_5175);
and U6237 (N_6237,N_5586,N_5049);
xor U6238 (N_6238,N_5843,N_5557);
xnor U6239 (N_6239,N_5449,N_5978);
xor U6240 (N_6240,N_5969,N_5206);
nor U6241 (N_6241,N_5664,N_5919);
xnor U6242 (N_6242,N_5338,N_5086);
and U6243 (N_6243,N_5134,N_5111);
nor U6244 (N_6244,N_5170,N_5160);
and U6245 (N_6245,N_5120,N_5958);
xnor U6246 (N_6246,N_5475,N_5934);
xor U6247 (N_6247,N_5504,N_5949);
or U6248 (N_6248,N_5045,N_5601);
nand U6249 (N_6249,N_5686,N_5501);
and U6250 (N_6250,N_5245,N_5519);
and U6251 (N_6251,N_5577,N_5604);
and U6252 (N_6252,N_5376,N_5634);
nor U6253 (N_6253,N_5288,N_5247);
and U6254 (N_6254,N_5890,N_5633);
or U6255 (N_6255,N_5252,N_5546);
nor U6256 (N_6256,N_5219,N_5494);
nand U6257 (N_6257,N_5126,N_5817);
nor U6258 (N_6258,N_5221,N_5844);
and U6259 (N_6259,N_5935,N_5666);
and U6260 (N_6260,N_5169,N_5511);
or U6261 (N_6261,N_5295,N_5972);
and U6262 (N_6262,N_5589,N_5645);
and U6263 (N_6263,N_5499,N_5435);
nand U6264 (N_6264,N_5862,N_5239);
nor U6265 (N_6265,N_5946,N_5434);
nand U6266 (N_6266,N_5942,N_5751);
nand U6267 (N_6267,N_5608,N_5838);
xnor U6268 (N_6268,N_5733,N_5757);
nor U6269 (N_6269,N_5250,N_5825);
or U6270 (N_6270,N_5368,N_5380);
or U6271 (N_6271,N_5540,N_5581);
nand U6272 (N_6272,N_5644,N_5315);
nor U6273 (N_6273,N_5023,N_5524);
nand U6274 (N_6274,N_5605,N_5624);
nand U6275 (N_6275,N_5801,N_5458);
or U6276 (N_6276,N_5102,N_5255);
nand U6277 (N_6277,N_5210,N_5881);
or U6278 (N_6278,N_5171,N_5749);
or U6279 (N_6279,N_5332,N_5017);
or U6280 (N_6280,N_5100,N_5675);
nor U6281 (N_6281,N_5615,N_5096);
nor U6282 (N_6282,N_5297,N_5892);
and U6283 (N_6283,N_5662,N_5069);
nor U6284 (N_6284,N_5921,N_5373);
and U6285 (N_6285,N_5822,N_5778);
nand U6286 (N_6286,N_5405,N_5190);
or U6287 (N_6287,N_5616,N_5292);
nor U6288 (N_6288,N_5683,N_5397);
nand U6289 (N_6289,N_5133,N_5238);
xnor U6290 (N_6290,N_5545,N_5803);
nand U6291 (N_6291,N_5804,N_5685);
or U6292 (N_6292,N_5342,N_5139);
xnor U6293 (N_6293,N_5523,N_5185);
nor U6294 (N_6294,N_5101,N_5357);
or U6295 (N_6295,N_5029,N_5131);
or U6296 (N_6296,N_5979,N_5184);
xnor U6297 (N_6297,N_5020,N_5791);
nor U6298 (N_6298,N_5936,N_5879);
xnor U6299 (N_6299,N_5669,N_5022);
or U6300 (N_6300,N_5833,N_5598);
nor U6301 (N_6301,N_5390,N_5275);
nor U6302 (N_6302,N_5781,N_5468);
nand U6303 (N_6303,N_5436,N_5717);
and U6304 (N_6304,N_5232,N_5068);
nand U6305 (N_6305,N_5646,N_5528);
nand U6306 (N_6306,N_5284,N_5891);
xor U6307 (N_6307,N_5649,N_5304);
nand U6308 (N_6308,N_5498,N_5951);
and U6309 (N_6309,N_5448,N_5144);
nand U6310 (N_6310,N_5773,N_5566);
or U6311 (N_6311,N_5696,N_5726);
and U6312 (N_6312,N_5476,N_5474);
nor U6313 (N_6313,N_5164,N_5928);
or U6314 (N_6314,N_5109,N_5489);
or U6315 (N_6315,N_5984,N_5915);
or U6316 (N_6316,N_5053,N_5593);
or U6317 (N_6317,N_5561,N_5595);
nor U6318 (N_6318,N_5763,N_5130);
nor U6319 (N_6319,N_5741,N_5323);
or U6320 (N_6320,N_5343,N_5377);
xor U6321 (N_6321,N_5600,N_5835);
or U6322 (N_6322,N_5663,N_5081);
xor U6323 (N_6323,N_5702,N_5208);
or U6324 (N_6324,N_5432,N_5466);
xor U6325 (N_6325,N_5962,N_5537);
nand U6326 (N_6326,N_5904,N_5371);
nor U6327 (N_6327,N_5364,N_5897);
nor U6328 (N_6328,N_5587,N_5470);
nor U6329 (N_6329,N_5354,N_5828);
nor U6330 (N_6330,N_5253,N_5971);
xor U6331 (N_6331,N_5121,N_5903);
and U6332 (N_6332,N_5421,N_5268);
xnor U6333 (N_6333,N_5954,N_5532);
and U6334 (N_6334,N_5225,N_5455);
xnor U6335 (N_6335,N_5341,N_5112);
xor U6336 (N_6336,N_5318,N_5302);
xnor U6337 (N_6337,N_5704,N_5079);
and U6338 (N_6338,N_5035,N_5997);
nor U6339 (N_6339,N_5853,N_5317);
or U6340 (N_6340,N_5481,N_5118);
xnor U6341 (N_6341,N_5456,N_5135);
nand U6342 (N_6342,N_5708,N_5103);
xnor U6343 (N_6343,N_5197,N_5261);
and U6344 (N_6344,N_5305,N_5720);
nand U6345 (N_6345,N_5379,N_5981);
xor U6346 (N_6346,N_5647,N_5670);
or U6347 (N_6347,N_5213,N_5864);
nor U6348 (N_6348,N_5612,N_5774);
xor U6349 (N_6349,N_5521,N_5242);
and U6350 (N_6350,N_5538,N_5347);
nor U6351 (N_6351,N_5230,N_5570);
or U6352 (N_6352,N_5544,N_5870);
xnor U6353 (N_6353,N_5871,N_5480);
and U6354 (N_6354,N_5365,N_5452);
xnor U6355 (N_6355,N_5067,N_5556);
nor U6356 (N_6356,N_5051,N_5046);
nor U6357 (N_6357,N_5472,N_5797);
and U6358 (N_6358,N_5924,N_5440);
nor U6359 (N_6359,N_5168,N_5855);
or U6360 (N_6360,N_5285,N_5286);
xor U6361 (N_6361,N_5901,N_5810);
nand U6362 (N_6362,N_5214,N_5766);
nor U6363 (N_6363,N_5218,N_5038);
nor U6364 (N_6364,N_5860,N_5569);
and U6365 (N_6365,N_5564,N_5005);
xor U6366 (N_6366,N_5910,N_5740);
or U6367 (N_6367,N_5567,N_5660);
nor U6368 (N_6368,N_5016,N_5422);
nor U6369 (N_6369,N_5628,N_5900);
nand U6370 (N_6370,N_5536,N_5146);
and U6371 (N_6371,N_5982,N_5301);
nand U6372 (N_6372,N_5240,N_5027);
nor U6373 (N_6373,N_5033,N_5887);
xor U6374 (N_6374,N_5927,N_5784);
xnor U6375 (N_6375,N_5678,N_5638);
nor U6376 (N_6376,N_5223,N_5047);
and U6377 (N_6377,N_5603,N_5224);
or U6378 (N_6378,N_5912,N_5976);
nand U6379 (N_6379,N_5950,N_5959);
and U6380 (N_6380,N_5677,N_5548);
nor U6381 (N_6381,N_5495,N_5830);
or U6382 (N_6382,N_5055,N_5216);
nand U6383 (N_6383,N_5490,N_5258);
and U6384 (N_6384,N_5254,N_5869);
nor U6385 (N_6385,N_5450,N_5505);
and U6386 (N_6386,N_5911,N_5857);
nor U6387 (N_6387,N_5932,N_5183);
nand U6388 (N_6388,N_5861,N_5917);
nor U6389 (N_6389,N_5789,N_5137);
nor U6390 (N_6390,N_5721,N_5732);
nand U6391 (N_6391,N_5404,N_5339);
nand U6392 (N_6392,N_5925,N_5311);
xor U6393 (N_6393,N_5525,N_5768);
and U6394 (N_6394,N_5880,N_5180);
nand U6395 (N_6395,N_5597,N_5674);
xor U6396 (N_6396,N_5488,N_5941);
or U6397 (N_6397,N_5609,N_5043);
nand U6398 (N_6398,N_5656,N_5514);
or U6399 (N_6399,N_5482,N_5056);
nor U6400 (N_6400,N_5209,N_5054);
or U6401 (N_6401,N_5582,N_5057);
and U6402 (N_6402,N_5372,N_5202);
xor U6403 (N_6403,N_5627,N_5330);
nand U6404 (N_6404,N_5508,N_5072);
xor U6405 (N_6405,N_5626,N_5114);
xor U6406 (N_6406,N_5734,N_5128);
nor U6407 (N_6407,N_5800,N_5155);
or U6408 (N_6408,N_5497,N_5780);
or U6409 (N_6409,N_5430,N_5477);
and U6410 (N_6410,N_5215,N_5510);
and U6411 (N_6411,N_5410,N_5199);
nand U6412 (N_6412,N_5092,N_5427);
xor U6413 (N_6413,N_5859,N_5516);
and U6414 (N_6414,N_5706,N_5299);
xor U6415 (N_6415,N_5992,N_5623);
nand U6416 (N_6416,N_5854,N_5659);
or U6417 (N_6417,N_5590,N_5201);
nor U6418 (N_6418,N_5004,N_5975);
nor U6419 (N_6419,N_5964,N_5014);
and U6420 (N_6420,N_5487,N_5007);
and U6421 (N_6421,N_5827,N_5602);
and U6422 (N_6422,N_5319,N_5279);
nand U6423 (N_6423,N_5163,N_5492);
and U6424 (N_6424,N_5457,N_5943);
or U6425 (N_6425,N_5375,N_5013);
xnor U6426 (N_6426,N_5622,N_5889);
nor U6427 (N_6427,N_5782,N_5189);
nor U6428 (N_6428,N_5465,N_5353);
nand U6429 (N_6429,N_5957,N_5186);
or U6430 (N_6430,N_5433,N_5743);
xnor U6431 (N_6431,N_5425,N_5990);
or U6432 (N_6432,N_5973,N_5515);
nor U6433 (N_6433,N_5705,N_5985);
or U6434 (N_6434,N_5270,N_5503);
nand U6435 (N_6435,N_5233,N_5746);
xor U6436 (N_6436,N_5147,N_5030);
xor U6437 (N_6437,N_5414,N_5930);
xor U6438 (N_6438,N_5262,N_5084);
and U6439 (N_6439,N_5779,N_5041);
nand U6440 (N_6440,N_5898,N_5203);
or U6441 (N_6441,N_5831,N_5709);
and U6442 (N_6442,N_5738,N_5522);
xnor U6443 (N_6443,N_5539,N_5796);
nand U6444 (N_6444,N_5392,N_5710);
or U6445 (N_6445,N_5818,N_5095);
or U6446 (N_6446,N_5922,N_5417);
nor U6447 (N_6447,N_5776,N_5851);
and U6448 (N_6448,N_5816,N_5836);
nor U6449 (N_6449,N_5658,N_5248);
and U6450 (N_6450,N_5276,N_5125);
and U6451 (N_6451,N_5036,N_5960);
xor U6452 (N_6452,N_5923,N_5865);
xor U6453 (N_6453,N_5272,N_5691);
nor U6454 (N_6454,N_5182,N_5222);
or U6455 (N_6455,N_5884,N_5730);
xor U6456 (N_6456,N_5256,N_5620);
and U6457 (N_6457,N_5080,N_5098);
xnor U6458 (N_6458,N_5393,N_5453);
nand U6459 (N_6459,N_5246,N_5396);
or U6460 (N_6460,N_5786,N_5697);
xnor U6461 (N_6461,N_5643,N_5042);
nand U6462 (N_6462,N_5725,N_5888);
and U6463 (N_6463,N_5579,N_5374);
xor U6464 (N_6464,N_5172,N_5234);
and U6465 (N_6465,N_5097,N_5676);
or U6466 (N_6466,N_5196,N_5760);
or U6467 (N_6467,N_5493,N_5770);
xnor U6468 (N_6468,N_5040,N_5575);
xor U6469 (N_6469,N_5032,N_5429);
nand U6470 (N_6470,N_5291,N_5148);
and U6471 (N_6471,N_5073,N_5875);
or U6472 (N_6472,N_5506,N_5650);
and U6473 (N_6473,N_5856,N_5106);
or U6474 (N_6474,N_5824,N_5731);
nor U6475 (N_6475,N_5306,N_5355);
nor U6476 (N_6476,N_5418,N_5269);
nand U6477 (N_6477,N_5070,N_5329);
nor U6478 (N_6478,N_5327,N_5826);
nand U6479 (N_6479,N_5241,N_5294);
and U6480 (N_6480,N_5177,N_5478);
xnor U6481 (N_6481,N_5411,N_5529);
nor U6482 (N_6482,N_5679,N_5689);
xnor U6483 (N_6483,N_5653,N_5001);
and U6484 (N_6484,N_5866,N_5654);
and U6485 (N_6485,N_5108,N_5104);
nor U6486 (N_6486,N_5039,N_5980);
nor U6487 (N_6487,N_5937,N_5090);
or U6488 (N_6488,N_5762,N_5560);
nand U6489 (N_6489,N_5082,N_5413);
nand U6490 (N_6490,N_5832,N_5745);
nand U6491 (N_6491,N_5829,N_5188);
nand U6492 (N_6492,N_5908,N_5156);
nand U6493 (N_6493,N_5428,N_5463);
xnor U6494 (N_6494,N_5727,N_5512);
or U6495 (N_6495,N_5558,N_5093);
xnor U6496 (N_6496,N_5289,N_5237);
xor U6497 (N_6497,N_5424,N_5667);
nand U6498 (N_6498,N_5783,N_5974);
or U6499 (N_6499,N_5122,N_5370);
nand U6500 (N_6500,N_5087,N_5161);
and U6501 (N_6501,N_5330,N_5227);
and U6502 (N_6502,N_5883,N_5549);
and U6503 (N_6503,N_5270,N_5987);
nor U6504 (N_6504,N_5623,N_5515);
and U6505 (N_6505,N_5153,N_5002);
and U6506 (N_6506,N_5767,N_5680);
and U6507 (N_6507,N_5266,N_5028);
nand U6508 (N_6508,N_5427,N_5860);
nand U6509 (N_6509,N_5206,N_5160);
and U6510 (N_6510,N_5467,N_5595);
and U6511 (N_6511,N_5217,N_5560);
and U6512 (N_6512,N_5701,N_5668);
xor U6513 (N_6513,N_5897,N_5391);
and U6514 (N_6514,N_5359,N_5404);
nand U6515 (N_6515,N_5990,N_5119);
nor U6516 (N_6516,N_5720,N_5971);
and U6517 (N_6517,N_5110,N_5656);
nor U6518 (N_6518,N_5552,N_5494);
and U6519 (N_6519,N_5072,N_5254);
nand U6520 (N_6520,N_5572,N_5289);
nand U6521 (N_6521,N_5306,N_5254);
nor U6522 (N_6522,N_5938,N_5264);
or U6523 (N_6523,N_5045,N_5683);
or U6524 (N_6524,N_5053,N_5518);
nand U6525 (N_6525,N_5425,N_5377);
xnor U6526 (N_6526,N_5866,N_5969);
nand U6527 (N_6527,N_5589,N_5624);
and U6528 (N_6528,N_5719,N_5771);
and U6529 (N_6529,N_5163,N_5335);
and U6530 (N_6530,N_5938,N_5056);
nor U6531 (N_6531,N_5046,N_5369);
xor U6532 (N_6532,N_5852,N_5150);
xor U6533 (N_6533,N_5195,N_5871);
and U6534 (N_6534,N_5793,N_5022);
or U6535 (N_6535,N_5072,N_5467);
nor U6536 (N_6536,N_5893,N_5117);
nor U6537 (N_6537,N_5882,N_5411);
or U6538 (N_6538,N_5930,N_5192);
or U6539 (N_6539,N_5556,N_5868);
xnor U6540 (N_6540,N_5730,N_5318);
or U6541 (N_6541,N_5528,N_5250);
or U6542 (N_6542,N_5066,N_5923);
nor U6543 (N_6543,N_5660,N_5424);
nand U6544 (N_6544,N_5180,N_5228);
nand U6545 (N_6545,N_5303,N_5155);
nand U6546 (N_6546,N_5157,N_5004);
xor U6547 (N_6547,N_5602,N_5267);
xor U6548 (N_6548,N_5066,N_5097);
and U6549 (N_6549,N_5733,N_5205);
and U6550 (N_6550,N_5795,N_5987);
or U6551 (N_6551,N_5618,N_5782);
nor U6552 (N_6552,N_5728,N_5179);
nor U6553 (N_6553,N_5957,N_5738);
xor U6554 (N_6554,N_5253,N_5323);
and U6555 (N_6555,N_5672,N_5133);
nand U6556 (N_6556,N_5273,N_5926);
nand U6557 (N_6557,N_5729,N_5299);
and U6558 (N_6558,N_5822,N_5061);
or U6559 (N_6559,N_5657,N_5593);
xnor U6560 (N_6560,N_5318,N_5064);
and U6561 (N_6561,N_5275,N_5104);
or U6562 (N_6562,N_5432,N_5160);
nor U6563 (N_6563,N_5587,N_5240);
nor U6564 (N_6564,N_5733,N_5979);
or U6565 (N_6565,N_5505,N_5570);
or U6566 (N_6566,N_5027,N_5958);
xor U6567 (N_6567,N_5596,N_5929);
nor U6568 (N_6568,N_5677,N_5517);
xnor U6569 (N_6569,N_5425,N_5665);
or U6570 (N_6570,N_5826,N_5614);
or U6571 (N_6571,N_5314,N_5891);
nor U6572 (N_6572,N_5721,N_5746);
and U6573 (N_6573,N_5606,N_5700);
nor U6574 (N_6574,N_5299,N_5882);
xnor U6575 (N_6575,N_5899,N_5244);
or U6576 (N_6576,N_5417,N_5088);
and U6577 (N_6577,N_5871,N_5453);
nand U6578 (N_6578,N_5867,N_5166);
xnor U6579 (N_6579,N_5318,N_5375);
nand U6580 (N_6580,N_5690,N_5739);
and U6581 (N_6581,N_5942,N_5351);
or U6582 (N_6582,N_5990,N_5003);
or U6583 (N_6583,N_5604,N_5597);
nor U6584 (N_6584,N_5588,N_5650);
nor U6585 (N_6585,N_5690,N_5352);
xnor U6586 (N_6586,N_5748,N_5872);
nand U6587 (N_6587,N_5495,N_5712);
nor U6588 (N_6588,N_5596,N_5248);
nand U6589 (N_6589,N_5614,N_5842);
or U6590 (N_6590,N_5755,N_5234);
or U6591 (N_6591,N_5496,N_5780);
xnor U6592 (N_6592,N_5965,N_5693);
or U6593 (N_6593,N_5091,N_5625);
or U6594 (N_6594,N_5559,N_5785);
nor U6595 (N_6595,N_5296,N_5236);
xnor U6596 (N_6596,N_5027,N_5072);
nand U6597 (N_6597,N_5529,N_5853);
nand U6598 (N_6598,N_5579,N_5136);
xnor U6599 (N_6599,N_5999,N_5281);
nand U6600 (N_6600,N_5074,N_5890);
nor U6601 (N_6601,N_5078,N_5008);
nand U6602 (N_6602,N_5166,N_5870);
or U6603 (N_6603,N_5537,N_5102);
xor U6604 (N_6604,N_5049,N_5754);
or U6605 (N_6605,N_5919,N_5472);
xor U6606 (N_6606,N_5155,N_5153);
xor U6607 (N_6607,N_5999,N_5870);
nor U6608 (N_6608,N_5840,N_5144);
xnor U6609 (N_6609,N_5835,N_5277);
or U6610 (N_6610,N_5771,N_5699);
and U6611 (N_6611,N_5112,N_5208);
xnor U6612 (N_6612,N_5409,N_5791);
nor U6613 (N_6613,N_5864,N_5712);
nand U6614 (N_6614,N_5249,N_5577);
nor U6615 (N_6615,N_5461,N_5847);
nand U6616 (N_6616,N_5444,N_5747);
nand U6617 (N_6617,N_5222,N_5781);
nor U6618 (N_6618,N_5038,N_5986);
and U6619 (N_6619,N_5546,N_5350);
or U6620 (N_6620,N_5125,N_5234);
nor U6621 (N_6621,N_5288,N_5437);
xnor U6622 (N_6622,N_5269,N_5037);
or U6623 (N_6623,N_5344,N_5583);
or U6624 (N_6624,N_5173,N_5271);
nand U6625 (N_6625,N_5839,N_5788);
and U6626 (N_6626,N_5739,N_5899);
or U6627 (N_6627,N_5366,N_5657);
nor U6628 (N_6628,N_5133,N_5784);
and U6629 (N_6629,N_5569,N_5812);
or U6630 (N_6630,N_5753,N_5132);
or U6631 (N_6631,N_5834,N_5142);
nand U6632 (N_6632,N_5956,N_5388);
xnor U6633 (N_6633,N_5517,N_5409);
nor U6634 (N_6634,N_5132,N_5631);
xor U6635 (N_6635,N_5037,N_5949);
and U6636 (N_6636,N_5989,N_5121);
and U6637 (N_6637,N_5177,N_5550);
xor U6638 (N_6638,N_5719,N_5510);
nor U6639 (N_6639,N_5377,N_5280);
and U6640 (N_6640,N_5558,N_5055);
nor U6641 (N_6641,N_5561,N_5986);
nand U6642 (N_6642,N_5513,N_5267);
xor U6643 (N_6643,N_5371,N_5456);
nor U6644 (N_6644,N_5436,N_5124);
and U6645 (N_6645,N_5512,N_5136);
nor U6646 (N_6646,N_5707,N_5606);
xnor U6647 (N_6647,N_5548,N_5417);
and U6648 (N_6648,N_5140,N_5972);
and U6649 (N_6649,N_5893,N_5229);
xnor U6650 (N_6650,N_5407,N_5104);
nor U6651 (N_6651,N_5909,N_5936);
nor U6652 (N_6652,N_5563,N_5449);
nand U6653 (N_6653,N_5869,N_5038);
and U6654 (N_6654,N_5185,N_5016);
and U6655 (N_6655,N_5925,N_5183);
and U6656 (N_6656,N_5352,N_5622);
and U6657 (N_6657,N_5446,N_5782);
nor U6658 (N_6658,N_5536,N_5918);
and U6659 (N_6659,N_5453,N_5142);
nor U6660 (N_6660,N_5508,N_5265);
nand U6661 (N_6661,N_5806,N_5197);
and U6662 (N_6662,N_5866,N_5976);
or U6663 (N_6663,N_5549,N_5864);
xnor U6664 (N_6664,N_5232,N_5055);
nor U6665 (N_6665,N_5381,N_5240);
and U6666 (N_6666,N_5299,N_5157);
nand U6667 (N_6667,N_5624,N_5082);
and U6668 (N_6668,N_5569,N_5017);
or U6669 (N_6669,N_5027,N_5405);
nor U6670 (N_6670,N_5057,N_5816);
nor U6671 (N_6671,N_5074,N_5211);
nand U6672 (N_6672,N_5819,N_5200);
nand U6673 (N_6673,N_5699,N_5217);
and U6674 (N_6674,N_5080,N_5020);
or U6675 (N_6675,N_5289,N_5859);
xnor U6676 (N_6676,N_5174,N_5941);
nor U6677 (N_6677,N_5263,N_5157);
or U6678 (N_6678,N_5940,N_5692);
or U6679 (N_6679,N_5446,N_5563);
nor U6680 (N_6680,N_5861,N_5930);
nor U6681 (N_6681,N_5868,N_5237);
and U6682 (N_6682,N_5534,N_5837);
nor U6683 (N_6683,N_5199,N_5746);
and U6684 (N_6684,N_5980,N_5332);
and U6685 (N_6685,N_5546,N_5206);
xnor U6686 (N_6686,N_5354,N_5662);
or U6687 (N_6687,N_5920,N_5116);
and U6688 (N_6688,N_5340,N_5488);
nor U6689 (N_6689,N_5631,N_5615);
nand U6690 (N_6690,N_5939,N_5605);
and U6691 (N_6691,N_5206,N_5636);
xnor U6692 (N_6692,N_5007,N_5873);
nor U6693 (N_6693,N_5331,N_5343);
or U6694 (N_6694,N_5932,N_5873);
xnor U6695 (N_6695,N_5572,N_5773);
nand U6696 (N_6696,N_5482,N_5759);
or U6697 (N_6697,N_5074,N_5592);
nand U6698 (N_6698,N_5838,N_5100);
nand U6699 (N_6699,N_5016,N_5926);
or U6700 (N_6700,N_5864,N_5426);
or U6701 (N_6701,N_5675,N_5884);
xor U6702 (N_6702,N_5000,N_5208);
nand U6703 (N_6703,N_5411,N_5809);
or U6704 (N_6704,N_5027,N_5156);
and U6705 (N_6705,N_5084,N_5649);
nor U6706 (N_6706,N_5814,N_5007);
nand U6707 (N_6707,N_5134,N_5519);
and U6708 (N_6708,N_5538,N_5551);
or U6709 (N_6709,N_5428,N_5162);
nand U6710 (N_6710,N_5737,N_5094);
nand U6711 (N_6711,N_5176,N_5677);
nand U6712 (N_6712,N_5495,N_5406);
xor U6713 (N_6713,N_5374,N_5751);
xor U6714 (N_6714,N_5201,N_5606);
nand U6715 (N_6715,N_5541,N_5857);
nand U6716 (N_6716,N_5621,N_5608);
xnor U6717 (N_6717,N_5486,N_5110);
xor U6718 (N_6718,N_5901,N_5714);
and U6719 (N_6719,N_5380,N_5825);
nand U6720 (N_6720,N_5357,N_5023);
or U6721 (N_6721,N_5985,N_5661);
xor U6722 (N_6722,N_5582,N_5709);
xnor U6723 (N_6723,N_5119,N_5154);
or U6724 (N_6724,N_5559,N_5113);
and U6725 (N_6725,N_5965,N_5445);
nor U6726 (N_6726,N_5378,N_5929);
or U6727 (N_6727,N_5534,N_5091);
nand U6728 (N_6728,N_5208,N_5597);
xor U6729 (N_6729,N_5057,N_5501);
and U6730 (N_6730,N_5201,N_5808);
or U6731 (N_6731,N_5858,N_5363);
and U6732 (N_6732,N_5465,N_5420);
and U6733 (N_6733,N_5721,N_5227);
xor U6734 (N_6734,N_5155,N_5256);
nand U6735 (N_6735,N_5500,N_5181);
or U6736 (N_6736,N_5463,N_5880);
xor U6737 (N_6737,N_5371,N_5967);
nand U6738 (N_6738,N_5474,N_5213);
xnor U6739 (N_6739,N_5980,N_5422);
nand U6740 (N_6740,N_5699,N_5893);
and U6741 (N_6741,N_5308,N_5691);
nand U6742 (N_6742,N_5134,N_5576);
nand U6743 (N_6743,N_5139,N_5379);
xor U6744 (N_6744,N_5526,N_5836);
or U6745 (N_6745,N_5713,N_5016);
xor U6746 (N_6746,N_5410,N_5308);
or U6747 (N_6747,N_5651,N_5236);
or U6748 (N_6748,N_5464,N_5375);
xor U6749 (N_6749,N_5411,N_5650);
nand U6750 (N_6750,N_5024,N_5118);
xnor U6751 (N_6751,N_5502,N_5162);
nor U6752 (N_6752,N_5817,N_5487);
or U6753 (N_6753,N_5672,N_5933);
and U6754 (N_6754,N_5055,N_5758);
nand U6755 (N_6755,N_5358,N_5963);
nor U6756 (N_6756,N_5948,N_5815);
nand U6757 (N_6757,N_5939,N_5210);
xor U6758 (N_6758,N_5430,N_5388);
nor U6759 (N_6759,N_5706,N_5132);
nand U6760 (N_6760,N_5609,N_5781);
and U6761 (N_6761,N_5621,N_5885);
and U6762 (N_6762,N_5594,N_5091);
or U6763 (N_6763,N_5140,N_5174);
or U6764 (N_6764,N_5880,N_5150);
or U6765 (N_6765,N_5089,N_5937);
xnor U6766 (N_6766,N_5864,N_5339);
nor U6767 (N_6767,N_5732,N_5971);
xnor U6768 (N_6768,N_5640,N_5545);
nor U6769 (N_6769,N_5797,N_5277);
nor U6770 (N_6770,N_5458,N_5792);
nand U6771 (N_6771,N_5976,N_5391);
and U6772 (N_6772,N_5744,N_5140);
or U6773 (N_6773,N_5230,N_5382);
xor U6774 (N_6774,N_5603,N_5119);
nor U6775 (N_6775,N_5185,N_5171);
xor U6776 (N_6776,N_5506,N_5608);
xor U6777 (N_6777,N_5610,N_5618);
and U6778 (N_6778,N_5431,N_5172);
nand U6779 (N_6779,N_5235,N_5470);
and U6780 (N_6780,N_5598,N_5448);
nand U6781 (N_6781,N_5145,N_5851);
or U6782 (N_6782,N_5428,N_5727);
or U6783 (N_6783,N_5829,N_5240);
and U6784 (N_6784,N_5659,N_5972);
xnor U6785 (N_6785,N_5567,N_5436);
nor U6786 (N_6786,N_5893,N_5642);
or U6787 (N_6787,N_5972,N_5882);
and U6788 (N_6788,N_5145,N_5560);
and U6789 (N_6789,N_5451,N_5472);
and U6790 (N_6790,N_5556,N_5123);
xor U6791 (N_6791,N_5078,N_5304);
xor U6792 (N_6792,N_5452,N_5728);
nand U6793 (N_6793,N_5995,N_5501);
nand U6794 (N_6794,N_5771,N_5842);
or U6795 (N_6795,N_5691,N_5358);
xnor U6796 (N_6796,N_5507,N_5973);
xor U6797 (N_6797,N_5697,N_5969);
xor U6798 (N_6798,N_5247,N_5666);
nor U6799 (N_6799,N_5642,N_5840);
nand U6800 (N_6800,N_5709,N_5636);
nand U6801 (N_6801,N_5271,N_5842);
and U6802 (N_6802,N_5090,N_5478);
or U6803 (N_6803,N_5309,N_5986);
nand U6804 (N_6804,N_5407,N_5470);
nand U6805 (N_6805,N_5161,N_5166);
nand U6806 (N_6806,N_5383,N_5871);
or U6807 (N_6807,N_5144,N_5439);
nor U6808 (N_6808,N_5212,N_5315);
or U6809 (N_6809,N_5237,N_5136);
xnor U6810 (N_6810,N_5213,N_5469);
nand U6811 (N_6811,N_5830,N_5052);
or U6812 (N_6812,N_5525,N_5897);
or U6813 (N_6813,N_5930,N_5183);
nor U6814 (N_6814,N_5080,N_5841);
nor U6815 (N_6815,N_5577,N_5451);
xor U6816 (N_6816,N_5002,N_5372);
nor U6817 (N_6817,N_5536,N_5993);
and U6818 (N_6818,N_5684,N_5757);
nor U6819 (N_6819,N_5495,N_5859);
xor U6820 (N_6820,N_5707,N_5451);
nand U6821 (N_6821,N_5077,N_5689);
and U6822 (N_6822,N_5048,N_5622);
or U6823 (N_6823,N_5759,N_5812);
nand U6824 (N_6824,N_5073,N_5250);
nor U6825 (N_6825,N_5140,N_5853);
or U6826 (N_6826,N_5422,N_5283);
nand U6827 (N_6827,N_5535,N_5498);
nor U6828 (N_6828,N_5264,N_5127);
and U6829 (N_6829,N_5507,N_5498);
xnor U6830 (N_6830,N_5375,N_5591);
and U6831 (N_6831,N_5488,N_5355);
nand U6832 (N_6832,N_5770,N_5725);
and U6833 (N_6833,N_5465,N_5044);
or U6834 (N_6834,N_5388,N_5180);
or U6835 (N_6835,N_5119,N_5033);
nand U6836 (N_6836,N_5746,N_5024);
xnor U6837 (N_6837,N_5306,N_5924);
xor U6838 (N_6838,N_5442,N_5752);
xnor U6839 (N_6839,N_5580,N_5250);
nand U6840 (N_6840,N_5282,N_5799);
nand U6841 (N_6841,N_5336,N_5743);
and U6842 (N_6842,N_5981,N_5895);
and U6843 (N_6843,N_5134,N_5266);
nand U6844 (N_6844,N_5764,N_5183);
nand U6845 (N_6845,N_5018,N_5746);
nand U6846 (N_6846,N_5918,N_5761);
or U6847 (N_6847,N_5727,N_5216);
and U6848 (N_6848,N_5314,N_5730);
nor U6849 (N_6849,N_5075,N_5801);
xor U6850 (N_6850,N_5618,N_5041);
and U6851 (N_6851,N_5957,N_5020);
nand U6852 (N_6852,N_5526,N_5897);
xor U6853 (N_6853,N_5480,N_5587);
or U6854 (N_6854,N_5430,N_5894);
and U6855 (N_6855,N_5509,N_5867);
nand U6856 (N_6856,N_5234,N_5103);
or U6857 (N_6857,N_5032,N_5912);
nor U6858 (N_6858,N_5376,N_5369);
or U6859 (N_6859,N_5774,N_5335);
and U6860 (N_6860,N_5931,N_5394);
and U6861 (N_6861,N_5521,N_5790);
nor U6862 (N_6862,N_5241,N_5588);
and U6863 (N_6863,N_5794,N_5373);
xnor U6864 (N_6864,N_5161,N_5335);
xor U6865 (N_6865,N_5225,N_5894);
xor U6866 (N_6866,N_5237,N_5809);
xor U6867 (N_6867,N_5429,N_5458);
or U6868 (N_6868,N_5014,N_5205);
nand U6869 (N_6869,N_5390,N_5761);
or U6870 (N_6870,N_5237,N_5324);
xor U6871 (N_6871,N_5780,N_5035);
or U6872 (N_6872,N_5799,N_5273);
and U6873 (N_6873,N_5380,N_5301);
nor U6874 (N_6874,N_5790,N_5263);
xor U6875 (N_6875,N_5827,N_5970);
or U6876 (N_6876,N_5683,N_5374);
or U6877 (N_6877,N_5188,N_5761);
xor U6878 (N_6878,N_5230,N_5083);
nand U6879 (N_6879,N_5114,N_5424);
nand U6880 (N_6880,N_5997,N_5914);
and U6881 (N_6881,N_5680,N_5751);
or U6882 (N_6882,N_5931,N_5233);
nor U6883 (N_6883,N_5849,N_5446);
nor U6884 (N_6884,N_5760,N_5441);
nand U6885 (N_6885,N_5284,N_5454);
or U6886 (N_6886,N_5365,N_5700);
or U6887 (N_6887,N_5491,N_5531);
xor U6888 (N_6888,N_5311,N_5190);
and U6889 (N_6889,N_5422,N_5391);
or U6890 (N_6890,N_5102,N_5202);
or U6891 (N_6891,N_5741,N_5880);
and U6892 (N_6892,N_5550,N_5097);
or U6893 (N_6893,N_5228,N_5223);
nor U6894 (N_6894,N_5984,N_5711);
nor U6895 (N_6895,N_5221,N_5568);
and U6896 (N_6896,N_5915,N_5649);
nor U6897 (N_6897,N_5220,N_5243);
nor U6898 (N_6898,N_5971,N_5965);
or U6899 (N_6899,N_5016,N_5655);
and U6900 (N_6900,N_5215,N_5030);
nor U6901 (N_6901,N_5339,N_5048);
nor U6902 (N_6902,N_5309,N_5037);
nor U6903 (N_6903,N_5213,N_5504);
xor U6904 (N_6904,N_5746,N_5925);
or U6905 (N_6905,N_5558,N_5767);
nor U6906 (N_6906,N_5326,N_5774);
or U6907 (N_6907,N_5450,N_5855);
nand U6908 (N_6908,N_5386,N_5197);
xnor U6909 (N_6909,N_5802,N_5812);
and U6910 (N_6910,N_5564,N_5543);
and U6911 (N_6911,N_5074,N_5104);
or U6912 (N_6912,N_5018,N_5152);
xor U6913 (N_6913,N_5611,N_5454);
nand U6914 (N_6914,N_5877,N_5026);
xnor U6915 (N_6915,N_5248,N_5464);
or U6916 (N_6916,N_5360,N_5270);
and U6917 (N_6917,N_5671,N_5696);
nand U6918 (N_6918,N_5170,N_5931);
or U6919 (N_6919,N_5231,N_5952);
or U6920 (N_6920,N_5798,N_5369);
nand U6921 (N_6921,N_5463,N_5649);
or U6922 (N_6922,N_5090,N_5164);
or U6923 (N_6923,N_5527,N_5143);
nor U6924 (N_6924,N_5515,N_5745);
nand U6925 (N_6925,N_5097,N_5224);
nand U6926 (N_6926,N_5511,N_5782);
or U6927 (N_6927,N_5532,N_5268);
xnor U6928 (N_6928,N_5815,N_5568);
nor U6929 (N_6929,N_5100,N_5448);
nand U6930 (N_6930,N_5134,N_5805);
or U6931 (N_6931,N_5186,N_5256);
or U6932 (N_6932,N_5132,N_5951);
nand U6933 (N_6933,N_5489,N_5414);
or U6934 (N_6934,N_5967,N_5585);
nand U6935 (N_6935,N_5582,N_5006);
nor U6936 (N_6936,N_5399,N_5729);
nor U6937 (N_6937,N_5587,N_5498);
or U6938 (N_6938,N_5466,N_5668);
and U6939 (N_6939,N_5571,N_5792);
nand U6940 (N_6940,N_5769,N_5517);
nor U6941 (N_6941,N_5778,N_5836);
nand U6942 (N_6942,N_5244,N_5586);
or U6943 (N_6943,N_5710,N_5247);
and U6944 (N_6944,N_5325,N_5983);
or U6945 (N_6945,N_5876,N_5936);
xnor U6946 (N_6946,N_5814,N_5873);
and U6947 (N_6947,N_5116,N_5665);
nand U6948 (N_6948,N_5657,N_5889);
xnor U6949 (N_6949,N_5736,N_5954);
xnor U6950 (N_6950,N_5363,N_5492);
or U6951 (N_6951,N_5702,N_5947);
nand U6952 (N_6952,N_5866,N_5547);
xor U6953 (N_6953,N_5917,N_5674);
nand U6954 (N_6954,N_5535,N_5257);
and U6955 (N_6955,N_5294,N_5511);
and U6956 (N_6956,N_5918,N_5711);
xor U6957 (N_6957,N_5207,N_5702);
or U6958 (N_6958,N_5005,N_5887);
and U6959 (N_6959,N_5577,N_5946);
and U6960 (N_6960,N_5445,N_5488);
xor U6961 (N_6961,N_5228,N_5871);
or U6962 (N_6962,N_5915,N_5711);
nor U6963 (N_6963,N_5851,N_5300);
nor U6964 (N_6964,N_5450,N_5319);
nor U6965 (N_6965,N_5898,N_5723);
nor U6966 (N_6966,N_5418,N_5385);
nand U6967 (N_6967,N_5788,N_5948);
nand U6968 (N_6968,N_5871,N_5303);
nor U6969 (N_6969,N_5510,N_5779);
and U6970 (N_6970,N_5423,N_5614);
nand U6971 (N_6971,N_5781,N_5516);
and U6972 (N_6972,N_5429,N_5096);
nand U6973 (N_6973,N_5485,N_5106);
or U6974 (N_6974,N_5560,N_5946);
nand U6975 (N_6975,N_5420,N_5158);
nand U6976 (N_6976,N_5255,N_5989);
nand U6977 (N_6977,N_5853,N_5358);
and U6978 (N_6978,N_5369,N_5422);
or U6979 (N_6979,N_5156,N_5036);
xor U6980 (N_6980,N_5453,N_5335);
nor U6981 (N_6981,N_5124,N_5423);
nand U6982 (N_6982,N_5465,N_5199);
or U6983 (N_6983,N_5551,N_5586);
and U6984 (N_6984,N_5817,N_5374);
nor U6985 (N_6985,N_5509,N_5576);
nand U6986 (N_6986,N_5384,N_5095);
and U6987 (N_6987,N_5231,N_5761);
nor U6988 (N_6988,N_5020,N_5087);
and U6989 (N_6989,N_5376,N_5397);
nand U6990 (N_6990,N_5255,N_5548);
nand U6991 (N_6991,N_5126,N_5443);
and U6992 (N_6992,N_5698,N_5087);
xor U6993 (N_6993,N_5291,N_5517);
or U6994 (N_6994,N_5095,N_5576);
or U6995 (N_6995,N_5027,N_5540);
xnor U6996 (N_6996,N_5572,N_5831);
and U6997 (N_6997,N_5150,N_5903);
or U6998 (N_6998,N_5055,N_5677);
and U6999 (N_6999,N_5739,N_5432);
nand U7000 (N_7000,N_6018,N_6202);
and U7001 (N_7001,N_6218,N_6711);
or U7002 (N_7002,N_6979,N_6215);
or U7003 (N_7003,N_6751,N_6161);
or U7004 (N_7004,N_6994,N_6805);
and U7005 (N_7005,N_6432,N_6718);
nor U7006 (N_7006,N_6801,N_6935);
nand U7007 (N_7007,N_6581,N_6545);
nand U7008 (N_7008,N_6458,N_6316);
nand U7009 (N_7009,N_6537,N_6734);
xnor U7010 (N_7010,N_6883,N_6904);
nor U7011 (N_7011,N_6291,N_6926);
and U7012 (N_7012,N_6838,N_6111);
xnor U7013 (N_7013,N_6040,N_6305);
nand U7014 (N_7014,N_6747,N_6995);
nor U7015 (N_7015,N_6705,N_6236);
nor U7016 (N_7016,N_6564,N_6219);
nor U7017 (N_7017,N_6532,N_6478);
or U7018 (N_7018,N_6619,N_6501);
xnor U7019 (N_7019,N_6508,N_6128);
nand U7020 (N_7020,N_6041,N_6333);
and U7021 (N_7021,N_6870,N_6715);
nor U7022 (N_7022,N_6209,N_6496);
nand U7023 (N_7023,N_6541,N_6140);
xnor U7024 (N_7024,N_6690,N_6370);
or U7025 (N_7025,N_6756,N_6712);
and U7026 (N_7026,N_6286,N_6616);
nand U7027 (N_7027,N_6518,N_6383);
nor U7028 (N_7028,N_6396,N_6073);
nand U7029 (N_7029,N_6210,N_6526);
nand U7030 (N_7030,N_6039,N_6669);
or U7031 (N_7031,N_6860,N_6068);
nor U7032 (N_7032,N_6583,N_6334);
nor U7033 (N_7033,N_6632,N_6266);
nand U7034 (N_7034,N_6562,N_6164);
nand U7035 (N_7035,N_6137,N_6951);
and U7036 (N_7036,N_6788,N_6520);
or U7037 (N_7037,N_6819,N_6782);
and U7038 (N_7038,N_6445,N_6058);
nor U7039 (N_7039,N_6067,N_6512);
xor U7040 (N_7040,N_6416,N_6276);
xor U7041 (N_7041,N_6138,N_6909);
or U7042 (N_7042,N_6798,N_6470);
or U7043 (N_7043,N_6672,N_6303);
nand U7044 (N_7044,N_6835,N_6611);
nand U7045 (N_7045,N_6373,N_6101);
nor U7046 (N_7046,N_6027,N_6548);
nor U7047 (N_7047,N_6425,N_6659);
nor U7048 (N_7048,N_6515,N_6451);
xnor U7049 (N_7049,N_6066,N_6230);
or U7050 (N_7050,N_6634,N_6667);
or U7051 (N_7051,N_6604,N_6369);
and U7052 (N_7052,N_6254,N_6925);
or U7053 (N_7053,N_6643,N_6016);
xnor U7054 (N_7054,N_6129,N_6142);
nor U7055 (N_7055,N_6580,N_6124);
and U7056 (N_7056,N_6681,N_6586);
nand U7057 (N_7057,N_6899,N_6504);
nor U7058 (N_7058,N_6623,N_6354);
or U7059 (N_7059,N_6176,N_6412);
and U7060 (N_7060,N_6948,N_6130);
nand U7061 (N_7061,N_6259,N_6280);
nor U7062 (N_7062,N_6543,N_6069);
nor U7063 (N_7063,N_6131,N_6208);
xor U7064 (N_7064,N_6574,N_6197);
nand U7065 (N_7065,N_6689,N_6404);
xor U7066 (N_7066,N_6653,N_6555);
nor U7067 (N_7067,N_6088,N_6189);
and U7068 (N_7068,N_6930,N_6043);
xor U7069 (N_7069,N_6380,N_6895);
and U7070 (N_7070,N_6503,N_6031);
nand U7071 (N_7071,N_6488,N_6491);
xnor U7072 (N_7072,N_6597,N_6765);
and U7073 (N_7073,N_6434,N_6549);
nand U7074 (N_7074,N_6566,N_6076);
or U7075 (N_7075,N_6652,N_6729);
and U7076 (N_7076,N_6850,N_6704);
nor U7077 (N_7077,N_6882,N_6047);
or U7078 (N_7078,N_6135,N_6575);
and U7079 (N_7079,N_6993,N_6072);
xor U7080 (N_7080,N_6185,N_6063);
or U7081 (N_7081,N_6519,N_6531);
nand U7082 (N_7082,N_6061,N_6961);
or U7083 (N_7083,N_6989,N_6848);
xnor U7084 (N_7084,N_6954,N_6405);
nor U7085 (N_7085,N_6193,N_6045);
and U7086 (N_7086,N_6213,N_6893);
nor U7087 (N_7087,N_6177,N_6028);
xnor U7088 (N_7088,N_6803,N_6625);
and U7089 (N_7089,N_6695,N_6326);
nor U7090 (N_7090,N_6113,N_6457);
nand U7091 (N_7091,N_6945,N_6618);
and U7092 (N_7092,N_6645,N_6139);
nor U7093 (N_7093,N_6024,N_6107);
nor U7094 (N_7094,N_6637,N_6627);
and U7095 (N_7095,N_6570,N_6206);
nor U7096 (N_7096,N_6832,N_6677);
and U7097 (N_7097,N_6292,N_6184);
nand U7098 (N_7098,N_6336,N_6448);
or U7099 (N_7099,N_6296,N_6557);
or U7100 (N_7100,N_6114,N_6340);
xnor U7101 (N_7101,N_6441,N_6392);
nor U7102 (N_7102,N_6235,N_6513);
xor U7103 (N_7103,N_6271,N_6071);
nor U7104 (N_7104,N_6269,N_6790);
xor U7105 (N_7105,N_6482,N_6023);
nor U7106 (N_7106,N_6005,N_6984);
xnor U7107 (N_7107,N_6430,N_6987);
nor U7108 (N_7108,N_6998,N_6845);
and U7109 (N_7109,N_6399,N_6789);
nor U7110 (N_7110,N_6827,N_6858);
xnor U7111 (N_7111,N_6602,N_6844);
nor U7112 (N_7112,N_6939,N_6004);
and U7113 (N_7113,N_6914,N_6795);
or U7114 (N_7114,N_6661,N_6676);
xor U7115 (N_7115,N_6364,N_6620);
xnor U7116 (N_7116,N_6194,N_6603);
nand U7117 (N_7117,N_6679,N_6720);
or U7118 (N_7118,N_6757,N_6356);
or U7119 (N_7119,N_6062,N_6477);
nor U7120 (N_7120,N_6083,N_6861);
nand U7121 (N_7121,N_6431,N_6360);
or U7122 (N_7122,N_6455,N_6959);
and U7123 (N_7123,N_6009,N_6320);
or U7124 (N_7124,N_6622,N_6484);
nor U7125 (N_7125,N_6818,N_6560);
nand U7126 (N_7126,N_6792,N_6258);
nand U7127 (N_7127,N_6947,N_6927);
nor U7128 (N_7128,N_6724,N_6701);
and U7129 (N_7129,N_6226,N_6162);
and U7130 (N_7130,N_6997,N_6579);
or U7131 (N_7131,N_6578,N_6825);
and U7132 (N_7132,N_6272,N_6243);
nor U7133 (N_7133,N_6942,N_6558);
nand U7134 (N_7134,N_6968,N_6294);
or U7135 (N_7135,N_6099,N_6890);
xnor U7136 (N_7136,N_6443,N_6025);
nand U7137 (N_7137,N_6651,N_6401);
nor U7138 (N_7138,N_6234,N_6332);
and U7139 (N_7139,N_6536,N_6078);
nand U7140 (N_7140,N_6466,N_6932);
xnor U7141 (N_7141,N_6461,N_6808);
and U7142 (N_7142,N_6937,N_6389);
and U7143 (N_7143,N_6148,N_6529);
nor U7144 (N_7144,N_6395,N_6530);
or U7145 (N_7145,N_6826,N_6863);
xnor U7146 (N_7146,N_6797,N_6688);
and U7147 (N_7147,N_6507,N_6535);
or U7148 (N_7148,N_6666,N_6875);
or U7149 (N_7149,N_6281,N_6517);
xor U7150 (N_7150,N_6884,N_6500);
and U7151 (N_7151,N_6468,N_6398);
nor U7152 (N_7152,N_6232,N_6778);
xor U7153 (N_7153,N_6382,N_6582);
nand U7154 (N_7154,N_6594,N_6924);
and U7155 (N_7155,N_6640,N_6471);
and U7156 (N_7156,N_6136,N_6736);
xor U7157 (N_7157,N_6685,N_6901);
and U7158 (N_7158,N_6132,N_6384);
and U7159 (N_7159,N_6601,N_6878);
nor U7160 (N_7160,N_6919,N_6033);
nand U7161 (N_7161,N_6522,N_6203);
xor U7162 (N_7162,N_6587,N_6742);
and U7163 (N_7163,N_6183,N_6344);
or U7164 (N_7164,N_6605,N_6973);
and U7165 (N_7165,N_6388,N_6319);
or U7166 (N_7166,N_6999,N_6056);
and U7167 (N_7167,N_6565,N_6426);
or U7168 (N_7168,N_6318,N_6506);
and U7169 (N_7169,N_6338,N_6008);
nand U7170 (N_7170,N_6190,N_6525);
or U7171 (N_7171,N_6248,N_6938);
xor U7172 (N_7172,N_6160,N_6436);
and U7173 (N_7173,N_6020,N_6417);
xnor U7174 (N_7174,N_6096,N_6894);
xnor U7175 (N_7175,N_6196,N_6379);
nand U7176 (N_7176,N_6728,N_6082);
nand U7177 (N_7177,N_6842,N_6420);
xnor U7178 (N_7178,N_6264,N_6793);
and U7179 (N_7179,N_6149,N_6084);
nand U7180 (N_7180,N_6171,N_6889);
and U7181 (N_7181,N_6493,N_6684);
and U7182 (N_7182,N_6915,N_6192);
xor U7183 (N_7183,N_6245,N_6527);
and U7184 (N_7184,N_6547,N_6607);
or U7185 (N_7185,N_6125,N_6996);
xor U7186 (N_7186,N_6559,N_6642);
or U7187 (N_7187,N_6635,N_6969);
nor U7188 (N_7188,N_6911,N_6780);
nand U7189 (N_7189,N_6165,N_6026);
or U7190 (N_7190,N_6181,N_6038);
or U7191 (N_7191,N_6774,N_6377);
or U7192 (N_7192,N_6204,N_6776);
nand U7193 (N_7193,N_6662,N_6873);
and U7194 (N_7194,N_6936,N_6567);
xor U7195 (N_7195,N_6748,N_6308);
or U7196 (N_7196,N_6049,N_6182);
nor U7197 (N_7197,N_6740,N_6497);
nand U7198 (N_7198,N_6775,N_6849);
nand U7199 (N_7199,N_6853,N_6002);
xnor U7200 (N_7200,N_6864,N_6631);
xnor U7201 (N_7201,N_6116,N_6486);
nor U7202 (N_7202,N_6505,N_6670);
nor U7203 (N_7203,N_6376,N_6606);
xor U7204 (N_7204,N_6714,N_6741);
and U7205 (N_7205,N_6381,N_6359);
nor U7206 (N_7206,N_6521,N_6810);
nor U7207 (N_7207,N_6962,N_6134);
nor U7208 (N_7208,N_6654,N_6386);
xor U7209 (N_7209,N_6820,N_6761);
or U7210 (N_7210,N_6828,N_6166);
nor U7211 (N_7211,N_6299,N_6674);
xor U7212 (N_7212,N_6551,N_6897);
xor U7213 (N_7213,N_6900,N_6422);
nor U7214 (N_7214,N_6610,N_6106);
nor U7215 (N_7215,N_6673,N_6785);
and U7216 (N_7216,N_6922,N_6593);
nand U7217 (N_7217,N_6881,N_6053);
xor U7218 (N_7218,N_6485,N_6591);
nand U7219 (N_7219,N_6006,N_6141);
and U7220 (N_7220,N_6198,N_6145);
xor U7221 (N_7221,N_6779,N_6042);
and U7222 (N_7222,N_6238,N_6007);
nor U7223 (N_7223,N_6524,N_6152);
and U7224 (N_7224,N_6304,N_6614);
and U7225 (N_7225,N_6424,N_6201);
or U7226 (N_7226,N_6867,N_6990);
xor U7227 (N_7227,N_6086,N_6239);
xnor U7228 (N_7228,N_6419,N_6624);
xnor U7229 (N_7229,N_6366,N_6514);
and U7230 (N_7230,N_6242,N_6978);
or U7231 (N_7231,N_6353,N_6017);
nor U7232 (N_7232,N_6663,N_6312);
nor U7233 (N_7233,N_6730,N_6691);
or U7234 (N_7234,N_6260,N_6064);
nor U7235 (N_7235,N_6928,N_6568);
and U7236 (N_7236,N_6091,N_6306);
and U7237 (N_7237,N_6363,N_6563);
or U7238 (N_7238,N_6977,N_6953);
nor U7239 (N_7239,N_6097,N_6214);
nand U7240 (N_7240,N_6133,N_6469);
xor U7241 (N_7241,N_6075,N_6777);
and U7242 (N_7242,N_6186,N_6121);
nand U7243 (N_7243,N_6358,N_6717);
and U7244 (N_7244,N_6081,N_6302);
or U7245 (N_7245,N_6284,N_6946);
nor U7246 (N_7246,N_6065,N_6290);
nor U7247 (N_7247,N_6408,N_6330);
nor U7248 (N_7248,N_6608,N_6112);
nand U7249 (N_7249,N_6630,N_6029);
and U7250 (N_7250,N_6743,N_6885);
or U7251 (N_7251,N_6722,N_6768);
nor U7252 (N_7252,N_6289,N_6092);
nand U7253 (N_7253,N_6371,N_6888);
or U7254 (N_7254,N_6589,N_6626);
or U7255 (N_7255,N_6975,N_6080);
and U7256 (N_7256,N_6079,N_6000);
and U7257 (N_7257,N_6511,N_6014);
and U7258 (N_7258,N_6686,N_6841);
and U7259 (N_7259,N_6944,N_6200);
nand U7260 (N_7260,N_6613,N_6971);
or U7261 (N_7261,N_6843,N_6721);
or U7262 (N_7262,N_6698,N_6172);
or U7263 (N_7263,N_6755,N_6647);
or U7264 (N_7264,N_6804,N_6749);
nand U7265 (N_7265,N_6710,N_6700);
nand U7266 (N_7266,N_6322,N_6949);
xnor U7267 (N_7267,N_6912,N_6746);
and U7268 (N_7268,N_6809,N_6313);
and U7269 (N_7269,N_6343,N_6905);
xnor U7270 (N_7270,N_6732,N_6950);
nand U7271 (N_7271,N_6829,N_6224);
and U7272 (N_7272,N_6699,N_6766);
nand U7273 (N_7273,N_6444,N_6475);
nor U7274 (N_7274,N_6090,N_6435);
and U7275 (N_7275,N_6816,N_6963);
and U7276 (N_7276,N_6246,N_6918);
nor U7277 (N_7277,N_6054,N_6599);
nand U7278 (N_7278,N_6982,N_6745);
nor U7279 (N_7279,N_6415,N_6429);
or U7280 (N_7280,N_6077,N_6314);
nand U7281 (N_7281,N_6929,N_6211);
and U7282 (N_7282,N_6390,N_6750);
nand U7283 (N_7283,N_6830,N_6146);
and U7284 (N_7284,N_6648,N_6921);
and U7285 (N_7285,N_6941,N_6753);
or U7286 (N_7286,N_6480,N_6010);
and U7287 (N_7287,N_6621,N_6463);
or U7288 (N_7288,N_6671,N_6220);
and U7289 (N_7289,N_6167,N_6854);
or U7290 (N_7290,N_6811,N_6095);
nor U7291 (N_7291,N_6769,N_6773);
or U7292 (N_7292,N_6288,N_6495);
or U7293 (N_7293,N_6481,N_6244);
and U7294 (N_7294,N_6903,N_6241);
xor U7295 (N_7295,N_6813,N_6298);
and U7296 (N_7296,N_6976,N_6833);
nor U7297 (N_7297,N_6655,N_6034);
and U7298 (N_7298,N_6931,N_6709);
and U7299 (N_7299,N_6231,N_6473);
nand U7300 (N_7300,N_6365,N_6301);
xnor U7301 (N_7301,N_6683,N_6986);
nor U7302 (N_7302,N_6315,N_6839);
xor U7303 (N_7303,N_6806,N_6019);
xnor U7304 (N_7304,N_6263,N_6085);
or U7305 (N_7305,N_6852,N_6433);
nor U7306 (N_7306,N_6955,N_6791);
nand U7307 (N_7307,N_6898,N_6665);
or U7308 (N_7308,N_6158,N_6913);
and U7309 (N_7309,N_6629,N_6752);
nand U7310 (N_7310,N_6030,N_6658);
or U7311 (N_7311,N_6649,N_6173);
nor U7312 (N_7312,N_6237,N_6474);
xnor U7313 (N_7313,N_6044,N_6644);
or U7314 (N_7314,N_6680,N_6050);
nand U7315 (N_7315,N_6784,N_6891);
nor U7316 (N_7316,N_6467,N_6588);
nor U7317 (N_7317,N_6759,N_6571);
xor U7318 (N_7318,N_6542,N_6253);
and U7319 (N_7319,N_6822,N_6059);
and U7320 (N_7320,N_6459,N_6410);
and U7321 (N_7321,N_6708,N_6847);
or U7322 (N_7322,N_6980,N_6221);
nor U7323 (N_7323,N_6692,N_6540);
xnor U7324 (N_7324,N_6857,N_6225);
nand U7325 (N_7325,N_6411,N_6550);
and U7326 (N_7326,N_6851,N_6702);
nand U7327 (N_7327,N_6011,N_6887);
nor U7328 (N_7328,N_6917,N_6546);
xor U7329 (N_7329,N_6787,N_6617);
xor U7330 (N_7330,N_6102,N_6351);
and U7331 (N_7331,N_6187,N_6533);
nor U7332 (N_7332,N_6057,N_6636);
nand U7333 (N_7333,N_6122,N_6807);
nor U7334 (N_7334,N_6483,N_6275);
nand U7335 (N_7335,N_6727,N_6633);
or U7336 (N_7336,N_6179,N_6494);
or U7337 (N_7337,N_6821,N_6638);
nand U7338 (N_7338,N_6277,N_6772);
and U7339 (N_7339,N_6438,N_6022);
xnor U7340 (N_7340,N_6409,N_6199);
nand U7341 (N_7341,N_6966,N_6297);
nand U7342 (N_7342,N_6222,N_6916);
nand U7343 (N_7343,N_6118,N_6960);
or U7344 (N_7344,N_6817,N_6476);
nand U7345 (N_7345,N_6440,N_6229);
or U7346 (N_7346,N_6534,N_6256);
nand U7347 (N_7347,N_6378,N_6402);
and U7348 (N_7348,N_6735,N_6910);
nand U7349 (N_7349,N_6802,N_6988);
and U7350 (N_7350,N_6492,N_6628);
xnor U7351 (N_7351,N_6595,N_6178);
xnor U7352 (N_7352,N_6325,N_6285);
nor U7353 (N_7353,N_6339,N_6584);
and U7354 (N_7354,N_6877,N_6035);
and U7355 (N_7355,N_6323,N_6418);
xor U7356 (N_7356,N_6697,N_6762);
nor U7357 (N_7357,N_6552,N_6207);
nor U7358 (N_7358,N_6874,N_6970);
nor U7359 (N_7359,N_6449,N_6021);
or U7360 (N_7360,N_6170,N_6127);
nand U7361 (N_7361,N_6573,N_6933);
nand U7362 (N_7362,N_6725,N_6413);
nand U7363 (N_7363,N_6771,N_6341);
nand U7364 (N_7364,N_6087,N_6329);
and U7365 (N_7365,N_6646,N_6823);
nand U7366 (N_7366,N_6965,N_6217);
or U7367 (N_7367,N_6387,N_6309);
nand U7368 (N_7368,N_6974,N_6615);
or U7369 (N_7369,N_6110,N_6153);
nor U7370 (N_7370,N_6331,N_6126);
xor U7371 (N_7371,N_6760,N_6716);
or U7372 (N_7372,N_6682,N_6585);
xnor U7373 (N_7373,N_6400,N_6923);
xor U7374 (N_7374,N_6865,N_6479);
nor U7375 (N_7375,N_6556,N_6046);
nand U7376 (N_7376,N_6675,N_6279);
xnor U7377 (N_7377,N_6855,N_6347);
or U7378 (N_7378,N_6880,N_6060);
or U7379 (N_7379,N_6036,N_6846);
xor U7380 (N_7380,N_6738,N_6561);
and U7381 (N_7381,N_6427,N_6233);
nand U7382 (N_7382,N_6733,N_6052);
and U7383 (N_7383,N_6109,N_6143);
and U7384 (N_7384,N_6490,N_6967);
or U7385 (N_7385,N_6337,N_6770);
xnor U7386 (N_7386,N_6499,N_6876);
and U7387 (N_7387,N_6287,N_6311);
or U7388 (N_7388,N_6981,N_6423);
and U7389 (N_7389,N_6015,N_6093);
nor U7390 (N_7390,N_6834,N_6032);
nor U7391 (N_7391,N_6355,N_6767);
and U7392 (N_7392,N_6321,N_6972);
nor U7393 (N_7393,N_6706,N_6367);
nor U7394 (N_7394,N_6055,N_6991);
nor U7395 (N_7395,N_6799,N_6660);
xnor U7396 (N_7396,N_6155,N_6569);
nor U7397 (N_7397,N_6836,N_6108);
nand U7398 (N_7398,N_6454,N_6456);
nor U7399 (N_7399,N_6668,N_6447);
and U7400 (N_7400,N_6783,N_6327);
xor U7401 (N_7401,N_6596,N_6528);
nand U7402 (N_7402,N_6012,N_6100);
xnor U7403 (N_7403,N_6592,N_6255);
xnor U7404 (N_7404,N_6437,N_6862);
xor U7405 (N_7405,N_6726,N_6737);
nand U7406 (N_7406,N_6048,N_6074);
or U7407 (N_7407,N_6103,N_6013);
nor U7408 (N_7408,N_6641,N_6147);
nand U7409 (N_7409,N_6159,N_6707);
nand U7410 (N_7410,N_6502,N_6693);
xor U7411 (N_7411,N_6442,N_6317);
and U7412 (N_7412,N_6781,N_6509);
nand U7413 (N_7413,N_6163,N_6452);
xor U7414 (N_7414,N_6157,N_6345);
xnor U7415 (N_7415,N_6453,N_6538);
nand U7416 (N_7416,N_6003,N_6815);
xor U7417 (N_7417,N_6267,N_6964);
nand U7418 (N_7418,N_6554,N_6920);
nand U7419 (N_7419,N_6576,N_6572);
nand U7420 (N_7420,N_6349,N_6465);
or U7421 (N_7421,N_6872,N_6421);
xnor U7422 (N_7422,N_6639,N_6800);
nor U7423 (N_7423,N_6374,N_6227);
and U7424 (N_7424,N_6144,N_6886);
xnor U7425 (N_7425,N_6168,N_6270);
nand U7426 (N_7426,N_6739,N_6723);
or U7427 (N_7427,N_6278,N_6151);
nor U7428 (N_7428,N_6544,N_6983);
and U7429 (N_7429,N_6385,N_6464);
xor U7430 (N_7430,N_6731,N_6051);
xnor U7431 (N_7431,N_6696,N_6089);
and U7432 (N_7432,N_6868,N_6119);
and U7433 (N_7433,N_6216,N_6758);
xor U7434 (N_7434,N_6307,N_6664);
or U7435 (N_7435,N_6462,N_6394);
and U7436 (N_7436,N_6117,N_6273);
nand U7437 (N_7437,N_6188,N_6115);
or U7438 (N_7438,N_6812,N_6169);
nor U7439 (N_7439,N_6678,N_6251);
nand U7440 (N_7440,N_6744,N_6391);
xnor U7441 (N_7441,N_6856,N_6037);
or U7442 (N_7442,N_6283,N_6361);
xnor U7443 (N_7443,N_6837,N_6257);
xor U7444 (N_7444,N_6539,N_6902);
nand U7445 (N_7445,N_6352,N_6335);
xnor U7446 (N_7446,N_6407,N_6205);
nand U7447 (N_7447,N_6450,N_6598);
nand U7448 (N_7448,N_6840,N_6871);
nand U7449 (N_7449,N_6105,N_6397);
or U7450 (N_7450,N_6191,N_6348);
or U7451 (N_7451,N_6156,N_6446);
and U7452 (N_7452,N_6265,N_6958);
nor U7453 (N_7453,N_6150,N_6814);
nand U7454 (N_7454,N_6590,N_6859);
and U7455 (N_7455,N_6368,N_6328);
nand U7456 (N_7456,N_6489,N_6510);
xnor U7457 (N_7457,N_6250,N_6357);
nand U7458 (N_7458,N_6869,N_6472);
or U7459 (N_7459,N_6293,N_6375);
and U7460 (N_7460,N_6553,N_6174);
xor U7461 (N_7461,N_6249,N_6831);
and U7462 (N_7462,N_6094,N_6439);
xnor U7463 (N_7463,N_6350,N_6906);
and U7464 (N_7464,N_6247,N_6713);
nor U7465 (N_7465,N_6703,N_6764);
nor U7466 (N_7466,N_6952,N_6403);
and U7467 (N_7467,N_6180,N_6957);
nor U7468 (N_7468,N_6896,N_6120);
nor U7469 (N_7469,N_6934,N_6212);
nor U7470 (N_7470,N_6282,N_6892);
or U7471 (N_7471,N_6516,N_6223);
nand U7472 (N_7472,N_6295,N_6650);
or U7473 (N_7473,N_6940,N_6070);
and U7474 (N_7474,N_6175,N_6612);
nor U7475 (N_7475,N_6796,N_6600);
nor U7476 (N_7476,N_6719,N_6123);
xor U7477 (N_7477,N_6261,N_6985);
nor U7478 (N_7478,N_6414,N_6794);
or U7479 (N_7479,N_6908,N_6346);
and U7480 (N_7480,N_6310,N_6609);
and U7481 (N_7481,N_6252,N_6406);
xor U7482 (N_7482,N_6342,N_6324);
nor U7483 (N_7483,N_6228,N_6428);
nand U7484 (N_7484,N_6098,N_6907);
or U7485 (N_7485,N_6001,N_6657);
nand U7486 (N_7486,N_6943,N_6754);
or U7487 (N_7487,N_6362,N_6879);
nor U7488 (N_7488,N_6656,N_6240);
nor U7489 (N_7489,N_6460,N_6487);
and U7490 (N_7490,N_6195,N_6154);
xor U7491 (N_7491,N_6393,N_6694);
xor U7492 (N_7492,N_6300,N_6498);
nor U7493 (N_7493,N_6268,N_6372);
nor U7494 (N_7494,N_6577,N_6763);
xnor U7495 (N_7495,N_6104,N_6523);
and U7496 (N_7496,N_6262,N_6992);
or U7497 (N_7497,N_6956,N_6824);
or U7498 (N_7498,N_6687,N_6274);
nand U7499 (N_7499,N_6786,N_6866);
or U7500 (N_7500,N_6318,N_6762);
nor U7501 (N_7501,N_6135,N_6922);
or U7502 (N_7502,N_6820,N_6525);
and U7503 (N_7503,N_6598,N_6030);
nand U7504 (N_7504,N_6849,N_6053);
nand U7505 (N_7505,N_6535,N_6869);
or U7506 (N_7506,N_6819,N_6425);
nor U7507 (N_7507,N_6361,N_6088);
xor U7508 (N_7508,N_6584,N_6902);
nand U7509 (N_7509,N_6733,N_6620);
xor U7510 (N_7510,N_6981,N_6029);
xor U7511 (N_7511,N_6056,N_6816);
and U7512 (N_7512,N_6840,N_6392);
and U7513 (N_7513,N_6482,N_6262);
or U7514 (N_7514,N_6106,N_6402);
and U7515 (N_7515,N_6878,N_6850);
nor U7516 (N_7516,N_6349,N_6576);
nor U7517 (N_7517,N_6219,N_6536);
nor U7518 (N_7518,N_6434,N_6709);
xor U7519 (N_7519,N_6548,N_6975);
and U7520 (N_7520,N_6904,N_6621);
nor U7521 (N_7521,N_6346,N_6318);
nand U7522 (N_7522,N_6845,N_6483);
nor U7523 (N_7523,N_6676,N_6578);
nand U7524 (N_7524,N_6827,N_6310);
and U7525 (N_7525,N_6078,N_6696);
or U7526 (N_7526,N_6437,N_6860);
xnor U7527 (N_7527,N_6046,N_6514);
and U7528 (N_7528,N_6958,N_6188);
xnor U7529 (N_7529,N_6720,N_6865);
and U7530 (N_7530,N_6403,N_6440);
nand U7531 (N_7531,N_6394,N_6712);
or U7532 (N_7532,N_6946,N_6210);
and U7533 (N_7533,N_6069,N_6220);
xor U7534 (N_7534,N_6227,N_6932);
nor U7535 (N_7535,N_6842,N_6418);
or U7536 (N_7536,N_6964,N_6516);
nand U7537 (N_7537,N_6791,N_6468);
nor U7538 (N_7538,N_6330,N_6000);
or U7539 (N_7539,N_6972,N_6306);
xor U7540 (N_7540,N_6485,N_6660);
or U7541 (N_7541,N_6875,N_6189);
nand U7542 (N_7542,N_6648,N_6933);
nor U7543 (N_7543,N_6280,N_6319);
and U7544 (N_7544,N_6415,N_6901);
and U7545 (N_7545,N_6697,N_6699);
xor U7546 (N_7546,N_6759,N_6150);
nand U7547 (N_7547,N_6707,N_6878);
xor U7548 (N_7548,N_6944,N_6113);
or U7549 (N_7549,N_6556,N_6841);
nor U7550 (N_7550,N_6599,N_6772);
xor U7551 (N_7551,N_6469,N_6532);
xor U7552 (N_7552,N_6198,N_6027);
nand U7553 (N_7553,N_6364,N_6312);
and U7554 (N_7554,N_6547,N_6512);
nand U7555 (N_7555,N_6974,N_6212);
nand U7556 (N_7556,N_6933,N_6441);
or U7557 (N_7557,N_6194,N_6521);
or U7558 (N_7558,N_6889,N_6159);
or U7559 (N_7559,N_6271,N_6955);
and U7560 (N_7560,N_6867,N_6589);
and U7561 (N_7561,N_6859,N_6494);
and U7562 (N_7562,N_6852,N_6157);
or U7563 (N_7563,N_6904,N_6388);
and U7564 (N_7564,N_6912,N_6481);
nor U7565 (N_7565,N_6670,N_6530);
nand U7566 (N_7566,N_6995,N_6933);
and U7567 (N_7567,N_6400,N_6559);
or U7568 (N_7568,N_6201,N_6518);
nor U7569 (N_7569,N_6180,N_6751);
and U7570 (N_7570,N_6839,N_6513);
nor U7571 (N_7571,N_6228,N_6274);
xor U7572 (N_7572,N_6002,N_6203);
nand U7573 (N_7573,N_6848,N_6156);
nand U7574 (N_7574,N_6277,N_6948);
nor U7575 (N_7575,N_6146,N_6719);
or U7576 (N_7576,N_6788,N_6253);
nor U7577 (N_7577,N_6139,N_6007);
or U7578 (N_7578,N_6728,N_6660);
and U7579 (N_7579,N_6493,N_6998);
nand U7580 (N_7580,N_6411,N_6848);
and U7581 (N_7581,N_6021,N_6890);
xnor U7582 (N_7582,N_6355,N_6975);
and U7583 (N_7583,N_6634,N_6295);
and U7584 (N_7584,N_6703,N_6469);
nand U7585 (N_7585,N_6410,N_6561);
or U7586 (N_7586,N_6351,N_6283);
or U7587 (N_7587,N_6725,N_6013);
nand U7588 (N_7588,N_6256,N_6713);
nor U7589 (N_7589,N_6271,N_6874);
or U7590 (N_7590,N_6533,N_6590);
xnor U7591 (N_7591,N_6123,N_6000);
or U7592 (N_7592,N_6934,N_6460);
and U7593 (N_7593,N_6465,N_6937);
or U7594 (N_7594,N_6564,N_6539);
nor U7595 (N_7595,N_6036,N_6772);
or U7596 (N_7596,N_6321,N_6749);
and U7597 (N_7597,N_6705,N_6588);
nor U7598 (N_7598,N_6160,N_6348);
and U7599 (N_7599,N_6289,N_6660);
nand U7600 (N_7600,N_6821,N_6274);
xor U7601 (N_7601,N_6287,N_6592);
or U7602 (N_7602,N_6285,N_6655);
nand U7603 (N_7603,N_6905,N_6034);
xnor U7604 (N_7604,N_6629,N_6134);
or U7605 (N_7605,N_6275,N_6998);
and U7606 (N_7606,N_6079,N_6041);
nand U7607 (N_7607,N_6475,N_6522);
or U7608 (N_7608,N_6028,N_6980);
and U7609 (N_7609,N_6947,N_6780);
nor U7610 (N_7610,N_6908,N_6774);
nor U7611 (N_7611,N_6292,N_6434);
xor U7612 (N_7612,N_6431,N_6998);
nand U7613 (N_7613,N_6790,N_6852);
nand U7614 (N_7614,N_6593,N_6943);
or U7615 (N_7615,N_6976,N_6387);
or U7616 (N_7616,N_6947,N_6724);
and U7617 (N_7617,N_6195,N_6680);
nor U7618 (N_7618,N_6666,N_6788);
xnor U7619 (N_7619,N_6926,N_6183);
xnor U7620 (N_7620,N_6868,N_6497);
or U7621 (N_7621,N_6829,N_6685);
and U7622 (N_7622,N_6684,N_6946);
or U7623 (N_7623,N_6765,N_6206);
nand U7624 (N_7624,N_6584,N_6017);
nor U7625 (N_7625,N_6829,N_6411);
xnor U7626 (N_7626,N_6266,N_6243);
or U7627 (N_7627,N_6579,N_6182);
and U7628 (N_7628,N_6657,N_6305);
or U7629 (N_7629,N_6883,N_6501);
xnor U7630 (N_7630,N_6401,N_6710);
and U7631 (N_7631,N_6655,N_6619);
nor U7632 (N_7632,N_6712,N_6660);
nand U7633 (N_7633,N_6127,N_6621);
or U7634 (N_7634,N_6725,N_6374);
and U7635 (N_7635,N_6171,N_6926);
xor U7636 (N_7636,N_6329,N_6620);
or U7637 (N_7637,N_6240,N_6988);
nor U7638 (N_7638,N_6415,N_6181);
or U7639 (N_7639,N_6617,N_6142);
or U7640 (N_7640,N_6639,N_6273);
or U7641 (N_7641,N_6206,N_6334);
and U7642 (N_7642,N_6498,N_6781);
nand U7643 (N_7643,N_6020,N_6090);
nand U7644 (N_7644,N_6786,N_6210);
nor U7645 (N_7645,N_6832,N_6890);
and U7646 (N_7646,N_6723,N_6495);
and U7647 (N_7647,N_6530,N_6264);
and U7648 (N_7648,N_6517,N_6525);
or U7649 (N_7649,N_6771,N_6912);
or U7650 (N_7650,N_6494,N_6834);
nor U7651 (N_7651,N_6177,N_6859);
and U7652 (N_7652,N_6849,N_6988);
or U7653 (N_7653,N_6340,N_6382);
nor U7654 (N_7654,N_6647,N_6542);
and U7655 (N_7655,N_6306,N_6930);
nor U7656 (N_7656,N_6369,N_6190);
nor U7657 (N_7657,N_6804,N_6242);
and U7658 (N_7658,N_6721,N_6765);
nand U7659 (N_7659,N_6152,N_6258);
and U7660 (N_7660,N_6455,N_6872);
or U7661 (N_7661,N_6691,N_6230);
xnor U7662 (N_7662,N_6374,N_6164);
or U7663 (N_7663,N_6505,N_6077);
or U7664 (N_7664,N_6029,N_6366);
xor U7665 (N_7665,N_6636,N_6845);
nor U7666 (N_7666,N_6877,N_6967);
or U7667 (N_7667,N_6475,N_6566);
or U7668 (N_7668,N_6512,N_6180);
nand U7669 (N_7669,N_6906,N_6635);
or U7670 (N_7670,N_6704,N_6942);
nand U7671 (N_7671,N_6289,N_6986);
and U7672 (N_7672,N_6845,N_6361);
or U7673 (N_7673,N_6567,N_6805);
nor U7674 (N_7674,N_6429,N_6046);
and U7675 (N_7675,N_6929,N_6796);
nand U7676 (N_7676,N_6219,N_6880);
xnor U7677 (N_7677,N_6544,N_6369);
or U7678 (N_7678,N_6853,N_6225);
xnor U7679 (N_7679,N_6136,N_6714);
nor U7680 (N_7680,N_6751,N_6801);
nand U7681 (N_7681,N_6424,N_6256);
nor U7682 (N_7682,N_6840,N_6035);
nor U7683 (N_7683,N_6990,N_6791);
nor U7684 (N_7684,N_6018,N_6580);
nor U7685 (N_7685,N_6825,N_6348);
nand U7686 (N_7686,N_6684,N_6165);
or U7687 (N_7687,N_6659,N_6338);
xor U7688 (N_7688,N_6330,N_6813);
nand U7689 (N_7689,N_6289,N_6178);
or U7690 (N_7690,N_6232,N_6751);
xor U7691 (N_7691,N_6198,N_6550);
nor U7692 (N_7692,N_6675,N_6346);
nand U7693 (N_7693,N_6532,N_6103);
nor U7694 (N_7694,N_6354,N_6427);
nor U7695 (N_7695,N_6285,N_6668);
nand U7696 (N_7696,N_6177,N_6705);
nor U7697 (N_7697,N_6747,N_6042);
nand U7698 (N_7698,N_6620,N_6904);
nor U7699 (N_7699,N_6564,N_6341);
or U7700 (N_7700,N_6842,N_6140);
and U7701 (N_7701,N_6507,N_6809);
and U7702 (N_7702,N_6773,N_6757);
or U7703 (N_7703,N_6627,N_6089);
or U7704 (N_7704,N_6042,N_6332);
and U7705 (N_7705,N_6349,N_6474);
nand U7706 (N_7706,N_6232,N_6809);
nor U7707 (N_7707,N_6339,N_6689);
nand U7708 (N_7708,N_6993,N_6110);
nor U7709 (N_7709,N_6509,N_6090);
nand U7710 (N_7710,N_6105,N_6345);
and U7711 (N_7711,N_6173,N_6653);
nand U7712 (N_7712,N_6862,N_6436);
and U7713 (N_7713,N_6959,N_6474);
nand U7714 (N_7714,N_6642,N_6111);
nand U7715 (N_7715,N_6875,N_6396);
nor U7716 (N_7716,N_6628,N_6065);
or U7717 (N_7717,N_6419,N_6083);
and U7718 (N_7718,N_6496,N_6598);
nand U7719 (N_7719,N_6538,N_6636);
and U7720 (N_7720,N_6416,N_6802);
and U7721 (N_7721,N_6565,N_6402);
nor U7722 (N_7722,N_6073,N_6435);
or U7723 (N_7723,N_6997,N_6534);
xnor U7724 (N_7724,N_6907,N_6747);
xnor U7725 (N_7725,N_6211,N_6010);
nor U7726 (N_7726,N_6288,N_6109);
xor U7727 (N_7727,N_6210,N_6374);
nor U7728 (N_7728,N_6034,N_6421);
or U7729 (N_7729,N_6435,N_6119);
or U7730 (N_7730,N_6203,N_6470);
nor U7731 (N_7731,N_6918,N_6178);
nand U7732 (N_7732,N_6150,N_6194);
nor U7733 (N_7733,N_6799,N_6396);
xnor U7734 (N_7734,N_6081,N_6232);
nand U7735 (N_7735,N_6353,N_6377);
nor U7736 (N_7736,N_6742,N_6404);
and U7737 (N_7737,N_6976,N_6006);
nand U7738 (N_7738,N_6214,N_6995);
and U7739 (N_7739,N_6856,N_6473);
xor U7740 (N_7740,N_6389,N_6125);
nor U7741 (N_7741,N_6272,N_6415);
xnor U7742 (N_7742,N_6228,N_6709);
and U7743 (N_7743,N_6952,N_6313);
or U7744 (N_7744,N_6132,N_6280);
and U7745 (N_7745,N_6463,N_6529);
or U7746 (N_7746,N_6741,N_6516);
or U7747 (N_7747,N_6693,N_6113);
nor U7748 (N_7748,N_6451,N_6107);
or U7749 (N_7749,N_6729,N_6131);
nand U7750 (N_7750,N_6907,N_6861);
xnor U7751 (N_7751,N_6936,N_6919);
nor U7752 (N_7752,N_6492,N_6207);
nand U7753 (N_7753,N_6444,N_6172);
nor U7754 (N_7754,N_6940,N_6899);
nand U7755 (N_7755,N_6547,N_6539);
nor U7756 (N_7756,N_6045,N_6653);
nand U7757 (N_7757,N_6315,N_6565);
xor U7758 (N_7758,N_6816,N_6775);
and U7759 (N_7759,N_6702,N_6113);
xor U7760 (N_7760,N_6325,N_6562);
or U7761 (N_7761,N_6751,N_6184);
xnor U7762 (N_7762,N_6170,N_6555);
nor U7763 (N_7763,N_6895,N_6624);
xnor U7764 (N_7764,N_6452,N_6404);
xor U7765 (N_7765,N_6384,N_6801);
and U7766 (N_7766,N_6551,N_6996);
xnor U7767 (N_7767,N_6830,N_6153);
or U7768 (N_7768,N_6766,N_6209);
or U7769 (N_7769,N_6089,N_6154);
or U7770 (N_7770,N_6286,N_6161);
xnor U7771 (N_7771,N_6421,N_6663);
nor U7772 (N_7772,N_6971,N_6828);
and U7773 (N_7773,N_6828,N_6682);
and U7774 (N_7774,N_6349,N_6003);
nand U7775 (N_7775,N_6234,N_6874);
or U7776 (N_7776,N_6167,N_6784);
and U7777 (N_7777,N_6707,N_6821);
and U7778 (N_7778,N_6062,N_6611);
nand U7779 (N_7779,N_6335,N_6071);
or U7780 (N_7780,N_6734,N_6479);
or U7781 (N_7781,N_6422,N_6868);
nand U7782 (N_7782,N_6809,N_6265);
nand U7783 (N_7783,N_6181,N_6920);
and U7784 (N_7784,N_6188,N_6696);
and U7785 (N_7785,N_6474,N_6822);
nor U7786 (N_7786,N_6801,N_6549);
nor U7787 (N_7787,N_6623,N_6173);
nand U7788 (N_7788,N_6632,N_6042);
and U7789 (N_7789,N_6555,N_6339);
and U7790 (N_7790,N_6587,N_6323);
xor U7791 (N_7791,N_6245,N_6148);
xor U7792 (N_7792,N_6233,N_6119);
nor U7793 (N_7793,N_6714,N_6423);
or U7794 (N_7794,N_6163,N_6089);
nor U7795 (N_7795,N_6613,N_6752);
or U7796 (N_7796,N_6799,N_6247);
nand U7797 (N_7797,N_6287,N_6368);
nor U7798 (N_7798,N_6967,N_6227);
nand U7799 (N_7799,N_6688,N_6675);
or U7800 (N_7800,N_6707,N_6493);
xnor U7801 (N_7801,N_6678,N_6541);
nand U7802 (N_7802,N_6073,N_6119);
and U7803 (N_7803,N_6207,N_6823);
xnor U7804 (N_7804,N_6778,N_6259);
or U7805 (N_7805,N_6787,N_6139);
nor U7806 (N_7806,N_6019,N_6613);
nand U7807 (N_7807,N_6524,N_6410);
nand U7808 (N_7808,N_6705,N_6079);
nand U7809 (N_7809,N_6052,N_6894);
nor U7810 (N_7810,N_6473,N_6360);
nor U7811 (N_7811,N_6655,N_6106);
nor U7812 (N_7812,N_6903,N_6274);
nor U7813 (N_7813,N_6129,N_6625);
or U7814 (N_7814,N_6707,N_6374);
and U7815 (N_7815,N_6549,N_6089);
nor U7816 (N_7816,N_6974,N_6347);
and U7817 (N_7817,N_6202,N_6853);
or U7818 (N_7818,N_6356,N_6882);
nor U7819 (N_7819,N_6636,N_6128);
or U7820 (N_7820,N_6755,N_6013);
nor U7821 (N_7821,N_6443,N_6896);
and U7822 (N_7822,N_6181,N_6549);
or U7823 (N_7823,N_6578,N_6243);
xor U7824 (N_7824,N_6589,N_6216);
nor U7825 (N_7825,N_6942,N_6514);
nor U7826 (N_7826,N_6269,N_6169);
nor U7827 (N_7827,N_6556,N_6226);
or U7828 (N_7828,N_6112,N_6952);
xnor U7829 (N_7829,N_6835,N_6787);
nand U7830 (N_7830,N_6669,N_6474);
xor U7831 (N_7831,N_6815,N_6798);
nor U7832 (N_7832,N_6598,N_6889);
and U7833 (N_7833,N_6836,N_6428);
and U7834 (N_7834,N_6519,N_6606);
and U7835 (N_7835,N_6641,N_6774);
xor U7836 (N_7836,N_6752,N_6864);
and U7837 (N_7837,N_6469,N_6419);
nand U7838 (N_7838,N_6912,N_6280);
or U7839 (N_7839,N_6934,N_6966);
xor U7840 (N_7840,N_6086,N_6395);
and U7841 (N_7841,N_6397,N_6675);
xor U7842 (N_7842,N_6676,N_6757);
nor U7843 (N_7843,N_6205,N_6257);
and U7844 (N_7844,N_6379,N_6896);
and U7845 (N_7845,N_6701,N_6138);
or U7846 (N_7846,N_6842,N_6917);
nor U7847 (N_7847,N_6605,N_6343);
xor U7848 (N_7848,N_6500,N_6391);
and U7849 (N_7849,N_6356,N_6251);
and U7850 (N_7850,N_6961,N_6303);
nor U7851 (N_7851,N_6259,N_6482);
or U7852 (N_7852,N_6862,N_6340);
nand U7853 (N_7853,N_6460,N_6665);
xor U7854 (N_7854,N_6135,N_6419);
xnor U7855 (N_7855,N_6810,N_6322);
or U7856 (N_7856,N_6005,N_6130);
or U7857 (N_7857,N_6373,N_6134);
and U7858 (N_7858,N_6142,N_6063);
and U7859 (N_7859,N_6957,N_6854);
nor U7860 (N_7860,N_6691,N_6334);
nand U7861 (N_7861,N_6364,N_6511);
nand U7862 (N_7862,N_6583,N_6239);
or U7863 (N_7863,N_6289,N_6696);
nor U7864 (N_7864,N_6292,N_6299);
nand U7865 (N_7865,N_6276,N_6663);
xnor U7866 (N_7866,N_6453,N_6351);
nor U7867 (N_7867,N_6890,N_6573);
and U7868 (N_7868,N_6092,N_6695);
or U7869 (N_7869,N_6009,N_6399);
or U7870 (N_7870,N_6249,N_6228);
nand U7871 (N_7871,N_6303,N_6124);
and U7872 (N_7872,N_6790,N_6811);
or U7873 (N_7873,N_6224,N_6137);
nand U7874 (N_7874,N_6396,N_6943);
or U7875 (N_7875,N_6693,N_6467);
xnor U7876 (N_7876,N_6300,N_6172);
nand U7877 (N_7877,N_6593,N_6542);
nand U7878 (N_7878,N_6896,N_6916);
xor U7879 (N_7879,N_6676,N_6965);
nor U7880 (N_7880,N_6559,N_6590);
or U7881 (N_7881,N_6696,N_6940);
nand U7882 (N_7882,N_6299,N_6063);
nor U7883 (N_7883,N_6335,N_6785);
nor U7884 (N_7884,N_6609,N_6734);
and U7885 (N_7885,N_6822,N_6080);
and U7886 (N_7886,N_6800,N_6124);
and U7887 (N_7887,N_6336,N_6564);
and U7888 (N_7888,N_6151,N_6037);
and U7889 (N_7889,N_6772,N_6428);
nand U7890 (N_7890,N_6538,N_6393);
nand U7891 (N_7891,N_6763,N_6976);
nor U7892 (N_7892,N_6054,N_6605);
xnor U7893 (N_7893,N_6654,N_6862);
or U7894 (N_7894,N_6103,N_6838);
nor U7895 (N_7895,N_6133,N_6957);
xnor U7896 (N_7896,N_6242,N_6981);
nor U7897 (N_7897,N_6586,N_6398);
xor U7898 (N_7898,N_6766,N_6341);
xor U7899 (N_7899,N_6643,N_6319);
and U7900 (N_7900,N_6586,N_6180);
nand U7901 (N_7901,N_6592,N_6214);
or U7902 (N_7902,N_6426,N_6111);
xor U7903 (N_7903,N_6741,N_6040);
nor U7904 (N_7904,N_6378,N_6056);
nor U7905 (N_7905,N_6022,N_6095);
or U7906 (N_7906,N_6393,N_6639);
and U7907 (N_7907,N_6206,N_6047);
xnor U7908 (N_7908,N_6122,N_6228);
and U7909 (N_7909,N_6924,N_6402);
nor U7910 (N_7910,N_6106,N_6645);
and U7911 (N_7911,N_6490,N_6789);
and U7912 (N_7912,N_6092,N_6362);
and U7913 (N_7913,N_6854,N_6513);
and U7914 (N_7914,N_6958,N_6920);
nor U7915 (N_7915,N_6370,N_6185);
or U7916 (N_7916,N_6511,N_6352);
xor U7917 (N_7917,N_6077,N_6188);
xnor U7918 (N_7918,N_6760,N_6999);
and U7919 (N_7919,N_6509,N_6912);
and U7920 (N_7920,N_6786,N_6428);
nand U7921 (N_7921,N_6156,N_6391);
nor U7922 (N_7922,N_6375,N_6998);
nand U7923 (N_7923,N_6114,N_6746);
nor U7924 (N_7924,N_6003,N_6716);
or U7925 (N_7925,N_6414,N_6736);
xnor U7926 (N_7926,N_6424,N_6916);
nand U7927 (N_7927,N_6158,N_6138);
nand U7928 (N_7928,N_6967,N_6987);
or U7929 (N_7929,N_6688,N_6781);
xnor U7930 (N_7930,N_6164,N_6854);
xnor U7931 (N_7931,N_6682,N_6270);
nor U7932 (N_7932,N_6005,N_6681);
or U7933 (N_7933,N_6286,N_6229);
and U7934 (N_7934,N_6938,N_6775);
nor U7935 (N_7935,N_6754,N_6873);
xor U7936 (N_7936,N_6373,N_6189);
xnor U7937 (N_7937,N_6784,N_6014);
nand U7938 (N_7938,N_6176,N_6242);
and U7939 (N_7939,N_6039,N_6725);
or U7940 (N_7940,N_6288,N_6547);
or U7941 (N_7941,N_6040,N_6875);
nor U7942 (N_7942,N_6304,N_6528);
or U7943 (N_7943,N_6339,N_6560);
and U7944 (N_7944,N_6946,N_6786);
nand U7945 (N_7945,N_6799,N_6813);
and U7946 (N_7946,N_6066,N_6308);
nand U7947 (N_7947,N_6630,N_6154);
or U7948 (N_7948,N_6349,N_6926);
nand U7949 (N_7949,N_6312,N_6995);
nand U7950 (N_7950,N_6243,N_6359);
nor U7951 (N_7951,N_6525,N_6294);
xor U7952 (N_7952,N_6060,N_6121);
nand U7953 (N_7953,N_6110,N_6519);
or U7954 (N_7954,N_6843,N_6276);
nor U7955 (N_7955,N_6506,N_6863);
xor U7956 (N_7956,N_6102,N_6820);
and U7957 (N_7957,N_6451,N_6913);
or U7958 (N_7958,N_6183,N_6247);
xnor U7959 (N_7959,N_6328,N_6387);
or U7960 (N_7960,N_6778,N_6729);
and U7961 (N_7961,N_6952,N_6640);
xnor U7962 (N_7962,N_6101,N_6241);
or U7963 (N_7963,N_6231,N_6240);
or U7964 (N_7964,N_6557,N_6421);
nor U7965 (N_7965,N_6881,N_6873);
nand U7966 (N_7966,N_6295,N_6299);
nand U7967 (N_7967,N_6311,N_6319);
nand U7968 (N_7968,N_6644,N_6381);
nand U7969 (N_7969,N_6300,N_6730);
and U7970 (N_7970,N_6202,N_6459);
or U7971 (N_7971,N_6126,N_6721);
nand U7972 (N_7972,N_6208,N_6710);
nor U7973 (N_7973,N_6617,N_6470);
and U7974 (N_7974,N_6539,N_6931);
nand U7975 (N_7975,N_6499,N_6553);
xnor U7976 (N_7976,N_6836,N_6835);
nand U7977 (N_7977,N_6235,N_6944);
and U7978 (N_7978,N_6047,N_6562);
or U7979 (N_7979,N_6511,N_6892);
and U7980 (N_7980,N_6445,N_6365);
xor U7981 (N_7981,N_6497,N_6215);
nor U7982 (N_7982,N_6347,N_6614);
nor U7983 (N_7983,N_6650,N_6097);
and U7984 (N_7984,N_6897,N_6903);
nand U7985 (N_7985,N_6929,N_6202);
and U7986 (N_7986,N_6447,N_6504);
and U7987 (N_7987,N_6726,N_6926);
xnor U7988 (N_7988,N_6166,N_6330);
nor U7989 (N_7989,N_6753,N_6324);
nand U7990 (N_7990,N_6435,N_6406);
and U7991 (N_7991,N_6502,N_6302);
nand U7992 (N_7992,N_6929,N_6885);
xor U7993 (N_7993,N_6097,N_6951);
xor U7994 (N_7994,N_6241,N_6885);
and U7995 (N_7995,N_6762,N_6013);
nor U7996 (N_7996,N_6725,N_6985);
nand U7997 (N_7997,N_6673,N_6754);
xnor U7998 (N_7998,N_6644,N_6997);
xnor U7999 (N_7999,N_6708,N_6570);
nor U8000 (N_8000,N_7056,N_7731);
nor U8001 (N_8001,N_7106,N_7745);
xnor U8002 (N_8002,N_7808,N_7529);
or U8003 (N_8003,N_7233,N_7453);
or U8004 (N_8004,N_7115,N_7517);
or U8005 (N_8005,N_7036,N_7120);
nor U8006 (N_8006,N_7050,N_7399);
or U8007 (N_8007,N_7743,N_7630);
nor U8008 (N_8008,N_7464,N_7130);
xnor U8009 (N_8009,N_7504,N_7721);
nand U8010 (N_8010,N_7067,N_7790);
and U8011 (N_8011,N_7373,N_7977);
or U8012 (N_8012,N_7351,N_7324);
nand U8013 (N_8013,N_7970,N_7898);
and U8014 (N_8014,N_7741,N_7817);
nand U8015 (N_8015,N_7596,N_7034);
and U8016 (N_8016,N_7735,N_7648);
and U8017 (N_8017,N_7971,N_7098);
nor U8018 (N_8018,N_7575,N_7592);
nor U8019 (N_8019,N_7822,N_7550);
or U8020 (N_8020,N_7462,N_7625);
xor U8021 (N_8021,N_7707,N_7236);
xor U8022 (N_8022,N_7931,N_7651);
or U8023 (N_8023,N_7813,N_7472);
nand U8024 (N_8024,N_7820,N_7599);
xor U8025 (N_8025,N_7455,N_7230);
nand U8026 (N_8026,N_7670,N_7295);
or U8027 (N_8027,N_7000,N_7011);
or U8028 (N_8028,N_7087,N_7296);
nor U8029 (N_8029,N_7170,N_7640);
nand U8030 (N_8030,N_7254,N_7330);
and U8031 (N_8031,N_7012,N_7283);
xnor U8032 (N_8032,N_7736,N_7891);
and U8033 (N_8033,N_7752,N_7191);
or U8034 (N_8034,N_7674,N_7053);
or U8035 (N_8035,N_7620,N_7398);
and U8036 (N_8036,N_7787,N_7627);
xor U8037 (N_8037,N_7342,N_7387);
xor U8038 (N_8038,N_7865,N_7671);
and U8039 (N_8039,N_7659,N_7570);
xnor U8040 (N_8040,N_7785,N_7202);
and U8041 (N_8041,N_7357,N_7435);
or U8042 (N_8042,N_7047,N_7471);
or U8043 (N_8043,N_7122,N_7232);
and U8044 (N_8044,N_7359,N_7172);
nand U8045 (N_8045,N_7904,N_7512);
and U8046 (N_8046,N_7196,N_7700);
nand U8047 (N_8047,N_7069,N_7317);
nor U8048 (N_8048,N_7896,N_7880);
or U8049 (N_8049,N_7159,N_7754);
xnor U8050 (N_8050,N_7681,N_7769);
xnor U8051 (N_8051,N_7677,N_7402);
nor U8052 (N_8052,N_7497,N_7100);
nor U8053 (N_8053,N_7634,N_7108);
nor U8054 (N_8054,N_7714,N_7003);
nand U8055 (N_8055,N_7713,N_7621);
or U8056 (N_8056,N_7834,N_7883);
nand U8057 (N_8057,N_7569,N_7993);
xor U8058 (N_8058,N_7217,N_7502);
and U8059 (N_8059,N_7601,N_7458);
or U8060 (N_8060,N_7310,N_7264);
and U8061 (N_8061,N_7021,N_7597);
nand U8062 (N_8062,N_7116,N_7886);
xor U8063 (N_8063,N_7679,N_7385);
xnor U8064 (N_8064,N_7258,N_7641);
and U8065 (N_8065,N_7306,N_7650);
nand U8066 (N_8066,N_7661,N_7119);
nor U8067 (N_8067,N_7010,N_7256);
or U8068 (N_8068,N_7345,N_7452);
or U8069 (N_8069,N_7383,N_7633);
xor U8070 (N_8070,N_7262,N_7533);
nor U8071 (N_8071,N_7163,N_7438);
xor U8072 (N_8072,N_7204,N_7604);
xor U8073 (N_8073,N_7835,N_7969);
xor U8074 (N_8074,N_7783,N_7781);
or U8075 (N_8075,N_7925,N_7810);
xnor U8076 (N_8076,N_7906,N_7197);
xor U8077 (N_8077,N_7124,N_7673);
or U8078 (N_8078,N_7910,N_7521);
nor U8079 (N_8079,N_7784,N_7096);
or U8080 (N_8080,N_7117,N_7941);
nor U8081 (N_8081,N_7049,N_7770);
nand U8082 (N_8082,N_7479,N_7894);
nor U8083 (N_8083,N_7267,N_7839);
xnor U8084 (N_8084,N_7953,N_7846);
and U8085 (N_8085,N_7722,N_7718);
nor U8086 (N_8086,N_7377,N_7358);
nor U8087 (N_8087,N_7637,N_7980);
nor U8088 (N_8088,N_7020,N_7414);
or U8089 (N_8089,N_7508,N_7747);
or U8090 (N_8090,N_7928,N_7303);
and U8091 (N_8091,N_7991,N_7921);
nand U8092 (N_8092,N_7060,N_7956);
or U8093 (N_8093,N_7147,N_7544);
nand U8094 (N_8094,N_7023,N_7128);
xnor U8095 (N_8095,N_7160,N_7214);
or U8096 (N_8096,N_7972,N_7442);
nor U8097 (N_8097,N_7923,N_7724);
nand U8098 (N_8098,N_7336,N_7663);
nor U8099 (N_8099,N_7755,N_7188);
nand U8100 (N_8100,N_7573,N_7048);
xnor U8101 (N_8101,N_7384,N_7698);
nor U8102 (N_8102,N_7838,N_7123);
and U8103 (N_8103,N_7942,N_7551);
nand U8104 (N_8104,N_7897,N_7001);
and U8105 (N_8105,N_7720,N_7238);
xnor U8106 (N_8106,N_7506,N_7436);
xnor U8107 (N_8107,N_7815,N_7346);
nor U8108 (N_8108,N_7428,N_7949);
nand U8109 (N_8109,N_7201,N_7693);
nor U8110 (N_8110,N_7675,N_7166);
nand U8111 (N_8111,N_7697,N_7040);
and U8112 (N_8112,N_7261,N_7967);
nand U8113 (N_8113,N_7688,N_7433);
nand U8114 (N_8114,N_7902,N_7999);
or U8115 (N_8115,N_7657,N_7181);
or U8116 (N_8116,N_7609,N_7668);
and U8117 (N_8117,N_7142,N_7632);
nand U8118 (N_8118,N_7178,N_7607);
and U8119 (N_8119,N_7733,N_7761);
nor U8120 (N_8120,N_7951,N_7626);
nand U8121 (N_8121,N_7811,N_7901);
and U8122 (N_8122,N_7498,N_7070);
nor U8123 (N_8123,N_7473,N_7848);
xor U8124 (N_8124,N_7638,N_7646);
and U8125 (N_8125,N_7474,N_7664);
and U8126 (N_8126,N_7247,N_7890);
nor U8127 (N_8127,N_7602,N_7847);
or U8128 (N_8128,N_7682,N_7667);
nand U8129 (N_8129,N_7503,N_7706);
nand U8130 (N_8130,N_7912,N_7501);
or U8131 (N_8131,N_7263,N_7006);
xnor U8132 (N_8132,N_7726,N_7809);
or U8133 (N_8133,N_7918,N_7806);
or U8134 (N_8134,N_7024,N_7183);
xor U8135 (N_8135,N_7818,N_7366);
nand U8136 (N_8136,N_7520,N_7369);
and U8137 (N_8137,N_7141,N_7655);
or U8138 (N_8138,N_7376,N_7444);
nand U8139 (N_8139,N_7807,N_7480);
nor U8140 (N_8140,N_7760,N_7407);
nand U8141 (N_8141,N_7856,N_7078);
nand U8142 (N_8142,N_7867,N_7654);
nor U8143 (N_8143,N_7276,N_7091);
and U8144 (N_8144,N_7537,N_7986);
or U8145 (N_8145,N_7059,N_7507);
and U8146 (N_8146,N_7995,N_7631);
xor U8147 (N_8147,N_7907,N_7423);
nand U8148 (N_8148,N_7052,N_7545);
and U8149 (N_8149,N_7938,N_7546);
or U8150 (N_8150,N_7605,N_7339);
or U8151 (N_8151,N_7088,N_7882);
xor U8152 (N_8152,N_7887,N_7354);
or U8153 (N_8153,N_7594,N_7045);
or U8154 (N_8154,N_7684,N_7775);
and U8155 (N_8155,N_7269,N_7516);
or U8156 (N_8156,N_7614,N_7788);
or U8157 (N_8157,N_7071,N_7092);
nand U8158 (N_8158,N_7135,N_7909);
nand U8159 (N_8159,N_7628,N_7982);
and U8160 (N_8160,N_7054,N_7103);
xor U8161 (N_8161,N_7061,N_7680);
nand U8162 (N_8162,N_7792,N_7943);
and U8163 (N_8163,N_7364,N_7603);
or U8164 (N_8164,N_7467,N_7094);
xnor U8165 (N_8165,N_7318,N_7137);
and U8166 (N_8166,N_7460,N_7290);
xor U8167 (N_8167,N_7246,N_7212);
and U8168 (N_8168,N_7211,N_7321);
xnor U8169 (N_8169,N_7114,N_7878);
nor U8170 (N_8170,N_7885,N_7046);
and U8171 (N_8171,N_7076,N_7486);
nand U8172 (N_8172,N_7463,N_7702);
nand U8173 (N_8173,N_7275,N_7029);
or U8174 (N_8174,N_7658,N_7827);
and U8175 (N_8175,N_7765,N_7136);
nand U8176 (N_8176,N_7844,N_7138);
nor U8177 (N_8177,N_7395,N_7187);
nor U8178 (N_8178,N_7057,N_7701);
xnor U8179 (N_8179,N_7379,N_7610);
xor U8180 (N_8180,N_7773,N_7585);
nand U8181 (N_8181,N_7235,N_7328);
xor U8182 (N_8182,N_7362,N_7753);
nand U8183 (N_8183,N_7996,N_7789);
nand U8184 (N_8184,N_7313,N_7484);
nor U8185 (N_8185,N_7421,N_7412);
and U8186 (N_8186,N_7375,N_7192);
nand U8187 (N_8187,N_7031,N_7948);
nand U8188 (N_8188,N_7562,N_7756);
and U8189 (N_8189,N_7372,N_7992);
or U8190 (N_8190,N_7919,N_7449);
nor U8191 (N_8191,N_7104,N_7341);
and U8192 (N_8192,N_7988,N_7690);
xor U8193 (N_8193,N_7833,N_7505);
or U8194 (N_8194,N_7782,N_7194);
xnor U8195 (N_8195,N_7899,N_7983);
and U8196 (N_8196,N_7764,N_7203);
or U8197 (N_8197,N_7535,N_7616);
nor U8198 (N_8198,N_7647,N_7308);
and U8199 (N_8199,N_7411,N_7591);
or U8200 (N_8200,N_7043,N_7889);
nand U8201 (N_8201,N_7265,N_7237);
nand U8202 (N_8202,N_7837,N_7552);
and U8203 (N_8203,N_7649,N_7410);
or U8204 (N_8204,N_7450,N_7557);
xnor U8205 (N_8205,N_7771,N_7612);
nor U8206 (N_8206,N_7424,N_7348);
or U8207 (N_8207,N_7853,N_7780);
or U8208 (N_8208,N_7536,N_7140);
nand U8209 (N_8209,N_7344,N_7038);
nor U8210 (N_8210,N_7073,N_7274);
nand U8211 (N_8211,N_7590,N_7990);
and U8212 (N_8212,N_7494,N_7572);
nand U8213 (N_8213,N_7405,N_7145);
or U8214 (N_8214,N_7962,N_7509);
and U8215 (N_8215,N_7759,N_7797);
nand U8216 (N_8216,N_7089,N_7873);
nor U8217 (N_8217,N_7843,N_7583);
and U8218 (N_8218,N_7016,N_7491);
nand U8219 (N_8219,N_7798,N_7678);
nor U8220 (N_8220,N_7729,N_7042);
xor U8221 (N_8221,N_7488,N_7805);
or U8222 (N_8222,N_7032,N_7493);
and U8223 (N_8223,N_7824,N_7903);
and U8224 (N_8224,N_7794,N_7716);
xnor U8225 (N_8225,N_7271,N_7957);
xnor U8226 (N_8226,N_7727,N_7945);
or U8227 (N_8227,N_7587,N_7109);
xor U8228 (N_8228,N_7408,N_7672);
or U8229 (N_8229,N_7959,N_7564);
nor U8230 (N_8230,N_7447,N_7800);
and U8231 (N_8231,N_7090,N_7763);
nor U8232 (N_8232,N_7371,N_7842);
or U8233 (N_8233,N_7580,N_7476);
xnor U8234 (N_8234,N_7221,N_7974);
or U8235 (N_8235,N_7589,N_7490);
nand U8236 (N_8236,N_7582,N_7732);
nand U8237 (N_8237,N_7397,N_7329);
and U8238 (N_8238,N_7944,N_7768);
and U8239 (N_8239,N_7427,N_7224);
and U8240 (N_8240,N_7102,N_7097);
nand U8241 (N_8241,N_7240,N_7017);
or U8242 (N_8242,N_7814,N_7598);
xnor U8243 (N_8243,N_7356,N_7155);
or U8244 (N_8244,N_7253,N_7394);
nor U8245 (N_8245,N_7757,N_7965);
xnor U8246 (N_8246,N_7466,N_7704);
xnor U8247 (N_8247,N_7439,N_7854);
xor U8248 (N_8248,N_7558,N_7293);
or U8249 (N_8249,N_7665,N_7298);
nand U8250 (N_8250,N_7863,N_7370);
and U8251 (N_8251,N_7892,N_7426);
and U8252 (N_8252,N_7861,N_7037);
nand U8253 (N_8253,N_7691,N_7565);
nor U8254 (N_8254,N_7255,N_7746);
xnor U8255 (N_8255,N_7245,N_7239);
nor U8256 (N_8256,N_7075,N_7567);
or U8257 (N_8257,N_7418,N_7401);
nor U8258 (N_8258,N_7710,N_7549);
xor U8259 (N_8259,N_7134,N_7812);
nor U8260 (N_8260,N_7776,N_7185);
xnor U8261 (N_8261,N_7522,N_7568);
nor U8262 (N_8262,N_7019,N_7378);
nor U8263 (N_8263,N_7685,N_7347);
nor U8264 (N_8264,N_7936,N_7532);
or U8265 (N_8265,N_7349,N_7617);
or U8266 (N_8266,N_7132,N_7802);
nand U8267 (N_8267,N_7461,N_7884);
xnor U8268 (N_8268,N_7009,N_7588);
or U8269 (N_8269,N_7916,N_7380);
xnor U8270 (N_8270,N_7850,N_7004);
and U8271 (N_8271,N_7500,N_7561);
or U8272 (N_8272,N_7465,N_7243);
nor U8273 (N_8273,N_7652,N_7419);
or U8274 (N_8274,N_7365,N_7958);
nor U8275 (N_8275,N_7767,N_7989);
and U8276 (N_8276,N_7093,N_7635);
nor U8277 (N_8277,N_7553,N_7234);
nor U8278 (N_8278,N_7955,N_7683);
xor U8279 (N_8279,N_7252,N_7248);
or U8280 (N_8280,N_7795,N_7353);
nor U8281 (N_8281,N_7391,N_7220);
nand U8282 (N_8282,N_7624,N_7209);
nor U8283 (N_8283,N_7779,N_7744);
xor U8284 (N_8284,N_7386,N_7186);
nand U8285 (N_8285,N_7259,N_7750);
nand U8286 (N_8286,N_7403,N_7730);
nor U8287 (N_8287,N_7456,N_7162);
and U8288 (N_8288,N_7699,N_7554);
or U8289 (N_8289,N_7857,N_7639);
and U8290 (N_8290,N_7985,N_7530);
nand U8291 (N_8291,N_7022,N_7297);
and U8292 (N_8292,N_7165,N_7828);
nor U8293 (N_8293,N_7420,N_7015);
or U8294 (N_8294,N_7855,N_7257);
nand U8295 (N_8295,N_7579,N_7081);
nor U8296 (N_8296,N_7825,N_7606);
and U8297 (N_8297,N_7051,N_7039);
nand U8298 (N_8298,N_7524,N_7177);
nand U8299 (N_8299,N_7175,N_7241);
or U8300 (N_8300,N_7156,N_7244);
nor U8301 (N_8301,N_7816,N_7796);
nor U8302 (N_8302,N_7870,N_7696);
xor U8303 (N_8303,N_7388,N_7893);
or U8304 (N_8304,N_7044,N_7208);
xnor U8305 (N_8305,N_7845,N_7618);
nand U8306 (N_8306,N_7915,N_7595);
or U8307 (N_8307,N_7819,N_7095);
or U8308 (N_8308,N_7748,N_7068);
xnor U8309 (N_8309,N_7085,N_7940);
and U8310 (N_8310,N_7964,N_7302);
and U8311 (N_8311,N_7272,N_7422);
xor U8312 (N_8312,N_7457,N_7190);
xnor U8313 (N_8313,N_7643,N_7823);
and U8314 (N_8314,N_7288,N_7519);
nand U8315 (N_8315,N_7879,N_7327);
or U8316 (N_8316,N_7284,N_7363);
nor U8317 (N_8317,N_7431,N_7981);
xor U8318 (N_8318,N_7709,N_7007);
or U8319 (N_8319,N_7874,N_7518);
and U8320 (N_8320,N_7282,N_7774);
nand U8321 (N_8321,N_7499,N_7143);
nor U8322 (N_8322,N_7198,N_7669);
or U8323 (N_8323,N_7305,N_7309);
nand U8324 (N_8324,N_7429,N_7619);
nand U8325 (N_8325,N_7852,N_7278);
or U8326 (N_8326,N_7542,N_7793);
nand U8327 (N_8327,N_7778,N_7223);
and U8328 (N_8328,N_7540,N_7723);
and U8329 (N_8329,N_7139,N_7973);
nor U8330 (N_8330,N_7074,N_7030);
or U8331 (N_8331,N_7531,N_7273);
nand U8332 (N_8332,N_7751,N_7703);
nor U8333 (N_8333,N_7876,N_7035);
xnor U8334 (N_8334,N_7390,N_7547);
and U8335 (N_8335,N_7443,N_7352);
nor U8336 (N_8336,N_7291,N_7413);
and U8337 (N_8337,N_7121,N_7934);
or U8338 (N_8338,N_7566,N_7523);
nor U8339 (N_8339,N_7425,N_7311);
nand U8340 (N_8340,N_7285,N_7099);
and U8341 (N_8341,N_7866,N_7041);
xor U8342 (N_8342,N_7393,N_7027);
and U8343 (N_8343,N_7469,N_7184);
xor U8344 (N_8344,N_7062,N_7055);
xor U8345 (N_8345,N_7742,N_7451);
xnor U8346 (N_8346,N_7560,N_7513);
xnor U8347 (N_8347,N_7332,N_7441);
nand U8348 (N_8348,N_7440,N_7218);
or U8349 (N_8349,N_7576,N_7644);
or U8350 (N_8350,N_7994,N_7737);
nor U8351 (N_8351,N_7005,N_7112);
and U8352 (N_8352,N_7868,N_7528);
and U8353 (N_8353,N_7577,N_7301);
nand U8354 (N_8354,N_7926,N_7932);
nand U8355 (N_8355,N_7448,N_7200);
or U8356 (N_8356,N_7922,N_7222);
nor U8357 (N_8357,N_7350,N_7066);
and U8358 (N_8358,N_7695,N_7622);
xnor U8359 (N_8359,N_7072,N_7437);
xor U8360 (N_8360,N_7434,N_7600);
nand U8361 (N_8361,N_7538,N_7803);
nor U8362 (N_8362,N_7801,N_7979);
and U8363 (N_8363,N_7525,N_7251);
nand U8364 (N_8364,N_7749,N_7900);
and U8365 (N_8365,N_7924,N_7821);
xor U8366 (N_8366,N_7266,N_7875);
nor U8367 (N_8367,N_7478,N_7527);
nor U8368 (N_8368,N_7367,N_7826);
nor U8369 (N_8369,N_7382,N_7791);
or U8370 (N_8370,N_7656,N_7064);
and U8371 (N_8371,N_7127,N_7319);
xor U8372 (N_8372,N_7584,N_7334);
nor U8373 (N_8373,N_7719,N_7337);
nor U8374 (N_8374,N_7065,N_7772);
xor U8375 (N_8375,N_7152,N_7608);
or U8376 (N_8376,N_7277,N_7860);
xnor U8377 (N_8377,N_7492,N_7111);
nor U8378 (N_8378,N_7930,N_7937);
or U8379 (N_8379,N_7740,N_7534);
xnor U8380 (N_8380,N_7927,N_7762);
nand U8381 (N_8381,N_7169,N_7477);
nand U8382 (N_8382,N_7777,N_7454);
and U8383 (N_8383,N_7864,N_7315);
nor U8384 (N_8384,N_7167,N_7280);
and U8385 (N_8385,N_7445,N_7739);
xnor U8386 (N_8386,N_7392,N_7687);
nand U8387 (N_8387,N_7998,N_7164);
and U8388 (N_8388,N_7689,N_7268);
nand U8389 (N_8389,N_7556,N_7287);
or U8390 (N_8390,N_7242,N_7586);
or U8391 (N_8391,N_7717,N_7326);
or U8392 (N_8392,N_7470,N_7154);
xor U8393 (N_8393,N_7933,N_7331);
or U8394 (N_8394,N_7881,N_7686);
and U8395 (N_8395,N_7908,N_7728);
and U8396 (N_8396,N_7961,N_7151);
or U8397 (N_8397,N_7836,N_7199);
and U8398 (N_8398,N_7249,N_7316);
nor U8399 (N_8399,N_7666,N_7338);
or U8400 (N_8400,N_7495,N_7216);
nor U8401 (N_8401,N_7862,N_7279);
nor U8402 (N_8402,N_7496,N_7193);
xor U8403 (N_8403,N_7294,N_7829);
and U8404 (N_8404,N_7734,N_7929);
or U8405 (N_8405,N_7153,N_7613);
xor U8406 (N_8406,N_7799,N_7396);
nand U8407 (N_8407,N_7227,N_7939);
xnor U8408 (N_8408,N_7299,N_7629);
xnor U8409 (N_8409,N_7653,N_7182);
xnor U8410 (N_8410,N_7555,N_7446);
or U8411 (N_8411,N_7270,N_7541);
nor U8412 (N_8412,N_7131,N_7058);
nand U8413 (N_8413,N_7148,N_7307);
or U8414 (N_8414,N_7840,N_7766);
nor U8415 (N_8415,N_7514,N_7195);
or U8416 (N_8416,N_7314,N_7543);
or U8417 (N_8417,N_7917,N_7804);
or U8418 (N_8418,N_7578,N_7260);
xnor U8419 (N_8419,N_7173,N_7642);
and U8420 (N_8420,N_7711,N_7946);
xnor U8421 (N_8421,N_7851,N_7636);
or U8422 (N_8422,N_7077,N_7215);
and U8423 (N_8423,N_7333,N_7250);
xor U8424 (N_8424,N_7758,N_7101);
nor U8425 (N_8425,N_7581,N_7725);
and U8426 (N_8426,N_7611,N_7229);
and U8427 (N_8427,N_7905,N_7082);
xnor U8428 (N_8428,N_7468,N_7228);
xor U8429 (N_8429,N_7086,N_7400);
nand U8430 (N_8430,N_7830,N_7323);
and U8431 (N_8431,N_7968,N_7485);
nand U8432 (N_8432,N_7660,N_7292);
nand U8433 (N_8433,N_7281,N_7786);
nand U8434 (N_8434,N_7430,N_7888);
and U8435 (N_8435,N_7920,N_7947);
nand U8436 (N_8436,N_7841,N_7343);
nor U8437 (N_8437,N_7623,N_7409);
nand U8438 (N_8438,N_7014,N_7322);
xor U8439 (N_8439,N_7389,N_7559);
and U8440 (N_8440,N_7571,N_7954);
xor U8441 (N_8441,N_7404,N_7645);
or U8442 (N_8442,N_7459,N_7110);
nor U8443 (N_8443,N_7335,N_7161);
nor U8444 (N_8444,N_7872,N_7432);
and U8445 (N_8445,N_7963,N_7935);
nand U8446 (N_8446,N_7859,N_7415);
nand U8447 (N_8447,N_7515,N_7026);
nor U8448 (N_8448,N_7858,N_7416);
and U8449 (N_8449,N_7511,N_7708);
or U8450 (N_8450,N_7487,N_7483);
and U8451 (N_8451,N_7914,N_7950);
nor U8452 (N_8452,N_7406,N_7355);
xnor U8453 (N_8453,N_7374,N_7219);
or U8454 (N_8454,N_7574,N_7368);
or U8455 (N_8455,N_7107,N_7176);
nand U8456 (N_8456,N_7158,N_7877);
and U8457 (N_8457,N_7174,N_7126);
and U8458 (N_8458,N_7913,N_7289);
and U8459 (N_8459,N_7189,N_7952);
and U8460 (N_8460,N_7738,N_7207);
nand U8461 (N_8461,N_7025,N_7340);
xor U8462 (N_8462,N_7028,N_7180);
and U8463 (N_8463,N_7975,N_7526);
xnor U8464 (N_8464,N_7063,N_7360);
nand U8465 (N_8465,N_7361,N_7079);
nand U8466 (N_8466,N_7300,N_7692);
nor U8467 (N_8467,N_7210,N_7133);
xnor U8468 (N_8468,N_7978,N_7563);
nor U8469 (N_8469,N_7381,N_7118);
xnor U8470 (N_8470,N_7084,N_7615);
nor U8471 (N_8471,N_7849,N_7676);
and U8472 (N_8472,N_7482,N_7966);
nand U8473 (N_8473,N_7033,N_7125);
nor U8474 (N_8474,N_7593,N_7997);
nor U8475 (N_8475,N_7013,N_7320);
nand U8476 (N_8476,N_7715,N_7105);
nand U8477 (N_8477,N_7548,N_7171);
nand U8478 (N_8478,N_7144,N_7481);
and U8479 (N_8479,N_7325,N_7960);
nor U8480 (N_8480,N_7149,N_7129);
or U8481 (N_8481,N_7987,N_7008);
or U8482 (N_8482,N_7831,N_7510);
or U8483 (N_8483,N_7489,N_7157);
or U8484 (N_8484,N_7080,N_7539);
xor U8485 (N_8485,N_7083,N_7871);
nor U8486 (N_8486,N_7226,N_7213);
nand U8487 (N_8487,N_7205,N_7231);
nand U8488 (N_8488,N_7312,N_7984);
nor U8489 (N_8489,N_7895,N_7705);
nor U8490 (N_8490,N_7712,N_7150);
nor U8491 (N_8491,N_7832,N_7976);
and U8492 (N_8492,N_7869,N_7694);
nand U8493 (N_8493,N_7286,N_7168);
and U8494 (N_8494,N_7146,N_7225);
or U8495 (N_8495,N_7113,N_7002);
and U8496 (N_8496,N_7911,N_7018);
nand U8497 (N_8497,N_7475,N_7206);
nor U8498 (N_8498,N_7662,N_7417);
or U8499 (N_8499,N_7304,N_7179);
and U8500 (N_8500,N_7068,N_7154);
nor U8501 (N_8501,N_7967,N_7884);
and U8502 (N_8502,N_7298,N_7941);
nor U8503 (N_8503,N_7401,N_7110);
xor U8504 (N_8504,N_7913,N_7850);
nand U8505 (N_8505,N_7023,N_7496);
and U8506 (N_8506,N_7606,N_7162);
xor U8507 (N_8507,N_7258,N_7837);
nand U8508 (N_8508,N_7792,N_7208);
nor U8509 (N_8509,N_7407,N_7049);
nand U8510 (N_8510,N_7835,N_7886);
and U8511 (N_8511,N_7882,N_7544);
nor U8512 (N_8512,N_7386,N_7957);
nand U8513 (N_8513,N_7240,N_7029);
and U8514 (N_8514,N_7677,N_7238);
xor U8515 (N_8515,N_7479,N_7928);
nor U8516 (N_8516,N_7639,N_7765);
or U8517 (N_8517,N_7278,N_7020);
and U8518 (N_8518,N_7114,N_7915);
nand U8519 (N_8519,N_7325,N_7682);
and U8520 (N_8520,N_7104,N_7486);
xnor U8521 (N_8521,N_7659,N_7438);
and U8522 (N_8522,N_7170,N_7195);
nand U8523 (N_8523,N_7985,N_7870);
nand U8524 (N_8524,N_7610,N_7235);
or U8525 (N_8525,N_7122,N_7540);
xnor U8526 (N_8526,N_7308,N_7474);
and U8527 (N_8527,N_7619,N_7595);
or U8528 (N_8528,N_7993,N_7578);
or U8529 (N_8529,N_7600,N_7095);
or U8530 (N_8530,N_7009,N_7772);
and U8531 (N_8531,N_7878,N_7798);
nand U8532 (N_8532,N_7212,N_7941);
xnor U8533 (N_8533,N_7436,N_7546);
nor U8534 (N_8534,N_7150,N_7105);
and U8535 (N_8535,N_7351,N_7915);
nand U8536 (N_8536,N_7769,N_7560);
nor U8537 (N_8537,N_7990,N_7994);
or U8538 (N_8538,N_7428,N_7207);
nand U8539 (N_8539,N_7003,N_7119);
or U8540 (N_8540,N_7499,N_7216);
nor U8541 (N_8541,N_7245,N_7717);
xor U8542 (N_8542,N_7133,N_7741);
xor U8543 (N_8543,N_7425,N_7279);
or U8544 (N_8544,N_7990,N_7215);
xor U8545 (N_8545,N_7506,N_7756);
or U8546 (N_8546,N_7361,N_7724);
or U8547 (N_8547,N_7227,N_7379);
nor U8548 (N_8548,N_7893,N_7644);
and U8549 (N_8549,N_7972,N_7492);
or U8550 (N_8550,N_7181,N_7534);
and U8551 (N_8551,N_7476,N_7483);
xnor U8552 (N_8552,N_7576,N_7587);
and U8553 (N_8553,N_7825,N_7279);
nor U8554 (N_8554,N_7492,N_7866);
nor U8555 (N_8555,N_7009,N_7179);
nor U8556 (N_8556,N_7408,N_7495);
or U8557 (N_8557,N_7425,N_7956);
and U8558 (N_8558,N_7717,N_7848);
nor U8559 (N_8559,N_7728,N_7437);
xor U8560 (N_8560,N_7875,N_7730);
nand U8561 (N_8561,N_7814,N_7878);
xor U8562 (N_8562,N_7401,N_7377);
or U8563 (N_8563,N_7202,N_7652);
xor U8564 (N_8564,N_7287,N_7515);
and U8565 (N_8565,N_7876,N_7814);
nand U8566 (N_8566,N_7392,N_7811);
nand U8567 (N_8567,N_7897,N_7986);
nor U8568 (N_8568,N_7462,N_7488);
nand U8569 (N_8569,N_7364,N_7633);
nand U8570 (N_8570,N_7293,N_7534);
xor U8571 (N_8571,N_7508,N_7096);
nand U8572 (N_8572,N_7420,N_7830);
nor U8573 (N_8573,N_7061,N_7726);
and U8574 (N_8574,N_7683,N_7769);
nand U8575 (N_8575,N_7880,N_7141);
nor U8576 (N_8576,N_7851,N_7447);
nand U8577 (N_8577,N_7152,N_7108);
or U8578 (N_8578,N_7211,N_7878);
or U8579 (N_8579,N_7579,N_7627);
xnor U8580 (N_8580,N_7297,N_7108);
or U8581 (N_8581,N_7909,N_7927);
xor U8582 (N_8582,N_7886,N_7680);
nor U8583 (N_8583,N_7169,N_7646);
nor U8584 (N_8584,N_7404,N_7923);
xor U8585 (N_8585,N_7055,N_7147);
or U8586 (N_8586,N_7942,N_7696);
xor U8587 (N_8587,N_7503,N_7960);
or U8588 (N_8588,N_7975,N_7102);
or U8589 (N_8589,N_7793,N_7417);
and U8590 (N_8590,N_7346,N_7766);
nand U8591 (N_8591,N_7666,N_7136);
nor U8592 (N_8592,N_7282,N_7862);
nand U8593 (N_8593,N_7767,N_7491);
nand U8594 (N_8594,N_7303,N_7291);
and U8595 (N_8595,N_7285,N_7954);
and U8596 (N_8596,N_7268,N_7064);
nor U8597 (N_8597,N_7444,N_7736);
and U8598 (N_8598,N_7738,N_7729);
nand U8599 (N_8599,N_7297,N_7758);
xor U8600 (N_8600,N_7532,N_7933);
and U8601 (N_8601,N_7047,N_7879);
or U8602 (N_8602,N_7693,N_7276);
and U8603 (N_8603,N_7408,N_7161);
nor U8604 (N_8604,N_7962,N_7177);
xor U8605 (N_8605,N_7820,N_7422);
or U8606 (N_8606,N_7651,N_7182);
nand U8607 (N_8607,N_7484,N_7502);
nand U8608 (N_8608,N_7062,N_7250);
nor U8609 (N_8609,N_7852,N_7440);
nand U8610 (N_8610,N_7466,N_7340);
nor U8611 (N_8611,N_7657,N_7259);
xnor U8612 (N_8612,N_7250,N_7163);
xnor U8613 (N_8613,N_7272,N_7848);
xnor U8614 (N_8614,N_7158,N_7252);
and U8615 (N_8615,N_7765,N_7767);
nand U8616 (N_8616,N_7546,N_7688);
nor U8617 (N_8617,N_7408,N_7537);
nand U8618 (N_8618,N_7160,N_7622);
xnor U8619 (N_8619,N_7113,N_7096);
or U8620 (N_8620,N_7785,N_7820);
nor U8621 (N_8621,N_7703,N_7841);
nand U8622 (N_8622,N_7781,N_7123);
and U8623 (N_8623,N_7177,N_7779);
or U8624 (N_8624,N_7554,N_7846);
and U8625 (N_8625,N_7899,N_7339);
nand U8626 (N_8626,N_7472,N_7488);
nand U8627 (N_8627,N_7204,N_7761);
nor U8628 (N_8628,N_7603,N_7157);
xnor U8629 (N_8629,N_7055,N_7579);
and U8630 (N_8630,N_7085,N_7478);
or U8631 (N_8631,N_7388,N_7582);
xor U8632 (N_8632,N_7384,N_7228);
or U8633 (N_8633,N_7137,N_7853);
and U8634 (N_8634,N_7037,N_7800);
nand U8635 (N_8635,N_7244,N_7254);
nor U8636 (N_8636,N_7949,N_7599);
xnor U8637 (N_8637,N_7853,N_7606);
and U8638 (N_8638,N_7779,N_7188);
nor U8639 (N_8639,N_7709,N_7025);
or U8640 (N_8640,N_7313,N_7557);
and U8641 (N_8641,N_7646,N_7789);
or U8642 (N_8642,N_7573,N_7536);
xor U8643 (N_8643,N_7124,N_7512);
and U8644 (N_8644,N_7810,N_7633);
and U8645 (N_8645,N_7971,N_7873);
and U8646 (N_8646,N_7769,N_7194);
xor U8647 (N_8647,N_7735,N_7352);
and U8648 (N_8648,N_7474,N_7566);
or U8649 (N_8649,N_7042,N_7373);
nand U8650 (N_8650,N_7237,N_7054);
and U8651 (N_8651,N_7589,N_7495);
and U8652 (N_8652,N_7953,N_7975);
and U8653 (N_8653,N_7988,N_7731);
or U8654 (N_8654,N_7263,N_7223);
nand U8655 (N_8655,N_7420,N_7518);
xnor U8656 (N_8656,N_7532,N_7279);
nor U8657 (N_8657,N_7697,N_7357);
xor U8658 (N_8658,N_7565,N_7692);
nand U8659 (N_8659,N_7923,N_7462);
and U8660 (N_8660,N_7587,N_7863);
or U8661 (N_8661,N_7789,N_7745);
xnor U8662 (N_8662,N_7963,N_7526);
nor U8663 (N_8663,N_7400,N_7632);
xor U8664 (N_8664,N_7069,N_7356);
nor U8665 (N_8665,N_7670,N_7558);
nand U8666 (N_8666,N_7759,N_7000);
and U8667 (N_8667,N_7303,N_7157);
nand U8668 (N_8668,N_7254,N_7660);
nand U8669 (N_8669,N_7720,N_7235);
and U8670 (N_8670,N_7474,N_7998);
and U8671 (N_8671,N_7834,N_7940);
nand U8672 (N_8672,N_7908,N_7514);
and U8673 (N_8673,N_7061,N_7476);
xor U8674 (N_8674,N_7507,N_7079);
and U8675 (N_8675,N_7197,N_7425);
xnor U8676 (N_8676,N_7377,N_7872);
nand U8677 (N_8677,N_7428,N_7689);
xor U8678 (N_8678,N_7041,N_7913);
nor U8679 (N_8679,N_7971,N_7311);
and U8680 (N_8680,N_7755,N_7975);
or U8681 (N_8681,N_7482,N_7950);
and U8682 (N_8682,N_7373,N_7630);
nand U8683 (N_8683,N_7837,N_7079);
xor U8684 (N_8684,N_7148,N_7971);
xor U8685 (N_8685,N_7515,N_7935);
xnor U8686 (N_8686,N_7811,N_7632);
nor U8687 (N_8687,N_7114,N_7551);
nand U8688 (N_8688,N_7631,N_7294);
nor U8689 (N_8689,N_7264,N_7344);
nand U8690 (N_8690,N_7791,N_7840);
and U8691 (N_8691,N_7152,N_7117);
or U8692 (N_8692,N_7152,N_7037);
xor U8693 (N_8693,N_7248,N_7611);
or U8694 (N_8694,N_7629,N_7319);
xnor U8695 (N_8695,N_7913,N_7596);
nor U8696 (N_8696,N_7301,N_7191);
nand U8697 (N_8697,N_7261,N_7515);
or U8698 (N_8698,N_7429,N_7973);
and U8699 (N_8699,N_7580,N_7300);
or U8700 (N_8700,N_7388,N_7734);
or U8701 (N_8701,N_7443,N_7599);
and U8702 (N_8702,N_7210,N_7484);
nand U8703 (N_8703,N_7405,N_7970);
nand U8704 (N_8704,N_7927,N_7239);
and U8705 (N_8705,N_7437,N_7365);
nor U8706 (N_8706,N_7033,N_7719);
or U8707 (N_8707,N_7918,N_7297);
xor U8708 (N_8708,N_7543,N_7786);
nand U8709 (N_8709,N_7394,N_7505);
nand U8710 (N_8710,N_7491,N_7709);
xor U8711 (N_8711,N_7937,N_7250);
nor U8712 (N_8712,N_7724,N_7633);
xnor U8713 (N_8713,N_7641,N_7405);
or U8714 (N_8714,N_7760,N_7775);
xnor U8715 (N_8715,N_7031,N_7615);
xnor U8716 (N_8716,N_7808,N_7183);
xor U8717 (N_8717,N_7511,N_7465);
nor U8718 (N_8718,N_7908,N_7014);
or U8719 (N_8719,N_7207,N_7427);
or U8720 (N_8720,N_7419,N_7627);
and U8721 (N_8721,N_7805,N_7690);
xnor U8722 (N_8722,N_7645,N_7912);
nand U8723 (N_8723,N_7713,N_7051);
and U8724 (N_8724,N_7180,N_7461);
and U8725 (N_8725,N_7436,N_7392);
or U8726 (N_8726,N_7097,N_7866);
xor U8727 (N_8727,N_7705,N_7086);
xor U8728 (N_8728,N_7228,N_7235);
and U8729 (N_8729,N_7984,N_7348);
nand U8730 (N_8730,N_7192,N_7843);
nand U8731 (N_8731,N_7398,N_7488);
or U8732 (N_8732,N_7474,N_7703);
xnor U8733 (N_8733,N_7805,N_7191);
or U8734 (N_8734,N_7393,N_7655);
xnor U8735 (N_8735,N_7539,N_7100);
or U8736 (N_8736,N_7616,N_7034);
nor U8737 (N_8737,N_7622,N_7311);
and U8738 (N_8738,N_7300,N_7151);
and U8739 (N_8739,N_7124,N_7845);
xor U8740 (N_8740,N_7745,N_7493);
or U8741 (N_8741,N_7295,N_7433);
nand U8742 (N_8742,N_7873,N_7693);
nand U8743 (N_8743,N_7324,N_7977);
nor U8744 (N_8744,N_7083,N_7916);
xor U8745 (N_8745,N_7758,N_7243);
or U8746 (N_8746,N_7048,N_7440);
nor U8747 (N_8747,N_7910,N_7412);
or U8748 (N_8748,N_7775,N_7869);
nand U8749 (N_8749,N_7611,N_7047);
and U8750 (N_8750,N_7865,N_7518);
nand U8751 (N_8751,N_7772,N_7835);
and U8752 (N_8752,N_7327,N_7285);
or U8753 (N_8753,N_7537,N_7762);
or U8754 (N_8754,N_7660,N_7546);
xnor U8755 (N_8755,N_7784,N_7128);
and U8756 (N_8756,N_7867,N_7734);
xnor U8757 (N_8757,N_7091,N_7920);
xnor U8758 (N_8758,N_7516,N_7933);
and U8759 (N_8759,N_7941,N_7783);
xnor U8760 (N_8760,N_7209,N_7400);
nor U8761 (N_8761,N_7256,N_7964);
nor U8762 (N_8762,N_7399,N_7064);
xnor U8763 (N_8763,N_7844,N_7764);
nor U8764 (N_8764,N_7677,N_7756);
xnor U8765 (N_8765,N_7187,N_7579);
xor U8766 (N_8766,N_7420,N_7470);
nor U8767 (N_8767,N_7928,N_7192);
nor U8768 (N_8768,N_7609,N_7240);
or U8769 (N_8769,N_7711,N_7172);
nand U8770 (N_8770,N_7638,N_7230);
nor U8771 (N_8771,N_7224,N_7270);
and U8772 (N_8772,N_7973,N_7106);
nand U8773 (N_8773,N_7387,N_7364);
nand U8774 (N_8774,N_7268,N_7009);
and U8775 (N_8775,N_7705,N_7629);
xnor U8776 (N_8776,N_7021,N_7672);
or U8777 (N_8777,N_7151,N_7673);
xor U8778 (N_8778,N_7801,N_7817);
or U8779 (N_8779,N_7970,N_7107);
nand U8780 (N_8780,N_7392,N_7698);
and U8781 (N_8781,N_7379,N_7499);
nor U8782 (N_8782,N_7731,N_7676);
xor U8783 (N_8783,N_7529,N_7892);
nor U8784 (N_8784,N_7766,N_7554);
or U8785 (N_8785,N_7015,N_7587);
nor U8786 (N_8786,N_7350,N_7807);
nand U8787 (N_8787,N_7003,N_7399);
nand U8788 (N_8788,N_7181,N_7299);
nand U8789 (N_8789,N_7356,N_7916);
and U8790 (N_8790,N_7302,N_7527);
xor U8791 (N_8791,N_7246,N_7234);
nor U8792 (N_8792,N_7651,N_7116);
nand U8793 (N_8793,N_7179,N_7069);
and U8794 (N_8794,N_7492,N_7961);
nor U8795 (N_8795,N_7408,N_7426);
nand U8796 (N_8796,N_7141,N_7143);
or U8797 (N_8797,N_7774,N_7667);
xor U8798 (N_8798,N_7789,N_7003);
xnor U8799 (N_8799,N_7805,N_7810);
nor U8800 (N_8800,N_7648,N_7601);
xnor U8801 (N_8801,N_7042,N_7619);
nand U8802 (N_8802,N_7054,N_7627);
nand U8803 (N_8803,N_7401,N_7274);
or U8804 (N_8804,N_7262,N_7004);
nand U8805 (N_8805,N_7288,N_7873);
or U8806 (N_8806,N_7351,N_7506);
nor U8807 (N_8807,N_7038,N_7040);
nor U8808 (N_8808,N_7132,N_7841);
xnor U8809 (N_8809,N_7259,N_7664);
or U8810 (N_8810,N_7460,N_7592);
nor U8811 (N_8811,N_7377,N_7975);
and U8812 (N_8812,N_7775,N_7935);
xnor U8813 (N_8813,N_7187,N_7391);
and U8814 (N_8814,N_7912,N_7069);
and U8815 (N_8815,N_7549,N_7323);
or U8816 (N_8816,N_7620,N_7643);
or U8817 (N_8817,N_7826,N_7659);
or U8818 (N_8818,N_7796,N_7441);
or U8819 (N_8819,N_7614,N_7967);
or U8820 (N_8820,N_7478,N_7107);
nand U8821 (N_8821,N_7673,N_7847);
nor U8822 (N_8822,N_7418,N_7570);
nand U8823 (N_8823,N_7961,N_7596);
nand U8824 (N_8824,N_7063,N_7979);
and U8825 (N_8825,N_7175,N_7565);
nand U8826 (N_8826,N_7417,N_7426);
or U8827 (N_8827,N_7120,N_7789);
or U8828 (N_8828,N_7282,N_7604);
nand U8829 (N_8829,N_7913,N_7839);
xor U8830 (N_8830,N_7297,N_7455);
or U8831 (N_8831,N_7141,N_7171);
and U8832 (N_8832,N_7578,N_7081);
nor U8833 (N_8833,N_7431,N_7251);
or U8834 (N_8834,N_7971,N_7951);
nor U8835 (N_8835,N_7666,N_7331);
and U8836 (N_8836,N_7961,N_7145);
xor U8837 (N_8837,N_7767,N_7986);
xor U8838 (N_8838,N_7226,N_7415);
and U8839 (N_8839,N_7047,N_7818);
or U8840 (N_8840,N_7421,N_7782);
xor U8841 (N_8841,N_7113,N_7536);
or U8842 (N_8842,N_7698,N_7024);
and U8843 (N_8843,N_7929,N_7423);
xor U8844 (N_8844,N_7487,N_7834);
xor U8845 (N_8845,N_7350,N_7175);
nand U8846 (N_8846,N_7228,N_7977);
xor U8847 (N_8847,N_7371,N_7504);
xor U8848 (N_8848,N_7742,N_7942);
or U8849 (N_8849,N_7929,N_7034);
and U8850 (N_8850,N_7390,N_7477);
and U8851 (N_8851,N_7229,N_7187);
nand U8852 (N_8852,N_7943,N_7168);
and U8853 (N_8853,N_7377,N_7997);
xnor U8854 (N_8854,N_7303,N_7835);
nor U8855 (N_8855,N_7233,N_7587);
or U8856 (N_8856,N_7291,N_7357);
nand U8857 (N_8857,N_7430,N_7597);
nor U8858 (N_8858,N_7243,N_7885);
xor U8859 (N_8859,N_7712,N_7815);
nand U8860 (N_8860,N_7836,N_7280);
nor U8861 (N_8861,N_7024,N_7603);
nor U8862 (N_8862,N_7473,N_7713);
xor U8863 (N_8863,N_7529,N_7091);
nor U8864 (N_8864,N_7321,N_7070);
or U8865 (N_8865,N_7681,N_7606);
and U8866 (N_8866,N_7454,N_7675);
nand U8867 (N_8867,N_7521,N_7821);
and U8868 (N_8868,N_7216,N_7603);
and U8869 (N_8869,N_7061,N_7258);
nand U8870 (N_8870,N_7414,N_7136);
or U8871 (N_8871,N_7337,N_7681);
nor U8872 (N_8872,N_7561,N_7361);
nand U8873 (N_8873,N_7255,N_7628);
or U8874 (N_8874,N_7781,N_7923);
nor U8875 (N_8875,N_7083,N_7605);
nor U8876 (N_8876,N_7336,N_7563);
nor U8877 (N_8877,N_7791,N_7585);
or U8878 (N_8878,N_7657,N_7090);
xnor U8879 (N_8879,N_7790,N_7996);
and U8880 (N_8880,N_7076,N_7515);
xnor U8881 (N_8881,N_7093,N_7283);
xor U8882 (N_8882,N_7470,N_7304);
and U8883 (N_8883,N_7114,N_7610);
and U8884 (N_8884,N_7140,N_7429);
nor U8885 (N_8885,N_7362,N_7136);
and U8886 (N_8886,N_7774,N_7974);
or U8887 (N_8887,N_7578,N_7344);
nor U8888 (N_8888,N_7938,N_7023);
xnor U8889 (N_8889,N_7657,N_7221);
xnor U8890 (N_8890,N_7131,N_7319);
nand U8891 (N_8891,N_7256,N_7539);
xnor U8892 (N_8892,N_7800,N_7810);
or U8893 (N_8893,N_7252,N_7576);
nand U8894 (N_8894,N_7045,N_7625);
nor U8895 (N_8895,N_7690,N_7874);
nand U8896 (N_8896,N_7067,N_7002);
nand U8897 (N_8897,N_7998,N_7939);
or U8898 (N_8898,N_7819,N_7768);
or U8899 (N_8899,N_7976,N_7194);
or U8900 (N_8900,N_7057,N_7292);
xnor U8901 (N_8901,N_7013,N_7568);
and U8902 (N_8902,N_7393,N_7604);
or U8903 (N_8903,N_7209,N_7085);
or U8904 (N_8904,N_7125,N_7805);
or U8905 (N_8905,N_7687,N_7803);
nand U8906 (N_8906,N_7740,N_7487);
nor U8907 (N_8907,N_7334,N_7472);
xnor U8908 (N_8908,N_7851,N_7973);
nand U8909 (N_8909,N_7741,N_7771);
xor U8910 (N_8910,N_7341,N_7331);
xor U8911 (N_8911,N_7728,N_7826);
nand U8912 (N_8912,N_7479,N_7316);
xnor U8913 (N_8913,N_7515,N_7975);
xnor U8914 (N_8914,N_7820,N_7341);
or U8915 (N_8915,N_7188,N_7182);
or U8916 (N_8916,N_7132,N_7194);
nand U8917 (N_8917,N_7413,N_7709);
and U8918 (N_8918,N_7016,N_7818);
nand U8919 (N_8919,N_7033,N_7006);
or U8920 (N_8920,N_7764,N_7963);
nor U8921 (N_8921,N_7284,N_7159);
and U8922 (N_8922,N_7356,N_7983);
xor U8923 (N_8923,N_7971,N_7413);
nor U8924 (N_8924,N_7103,N_7827);
nor U8925 (N_8925,N_7007,N_7417);
nor U8926 (N_8926,N_7366,N_7975);
nand U8927 (N_8927,N_7368,N_7130);
xnor U8928 (N_8928,N_7362,N_7327);
nand U8929 (N_8929,N_7797,N_7199);
and U8930 (N_8930,N_7214,N_7655);
or U8931 (N_8931,N_7273,N_7075);
nand U8932 (N_8932,N_7312,N_7733);
xnor U8933 (N_8933,N_7140,N_7130);
and U8934 (N_8934,N_7173,N_7742);
nor U8935 (N_8935,N_7291,N_7771);
and U8936 (N_8936,N_7739,N_7622);
or U8937 (N_8937,N_7615,N_7552);
and U8938 (N_8938,N_7480,N_7749);
and U8939 (N_8939,N_7651,N_7151);
and U8940 (N_8940,N_7981,N_7693);
or U8941 (N_8941,N_7781,N_7188);
and U8942 (N_8942,N_7226,N_7977);
and U8943 (N_8943,N_7790,N_7061);
or U8944 (N_8944,N_7964,N_7825);
nand U8945 (N_8945,N_7569,N_7939);
xor U8946 (N_8946,N_7277,N_7393);
xnor U8947 (N_8947,N_7708,N_7919);
or U8948 (N_8948,N_7969,N_7709);
nand U8949 (N_8949,N_7402,N_7335);
nand U8950 (N_8950,N_7982,N_7256);
nand U8951 (N_8951,N_7714,N_7183);
xnor U8952 (N_8952,N_7332,N_7684);
and U8953 (N_8953,N_7613,N_7545);
nor U8954 (N_8954,N_7434,N_7581);
xnor U8955 (N_8955,N_7444,N_7181);
and U8956 (N_8956,N_7489,N_7958);
or U8957 (N_8957,N_7343,N_7728);
xnor U8958 (N_8958,N_7634,N_7119);
or U8959 (N_8959,N_7844,N_7299);
xor U8960 (N_8960,N_7388,N_7919);
nand U8961 (N_8961,N_7965,N_7104);
or U8962 (N_8962,N_7385,N_7889);
nand U8963 (N_8963,N_7723,N_7663);
nand U8964 (N_8964,N_7900,N_7757);
nand U8965 (N_8965,N_7587,N_7896);
and U8966 (N_8966,N_7726,N_7141);
or U8967 (N_8967,N_7882,N_7212);
xor U8968 (N_8968,N_7509,N_7545);
or U8969 (N_8969,N_7277,N_7751);
nor U8970 (N_8970,N_7869,N_7907);
nor U8971 (N_8971,N_7422,N_7211);
nand U8972 (N_8972,N_7181,N_7665);
and U8973 (N_8973,N_7153,N_7949);
nand U8974 (N_8974,N_7891,N_7920);
nand U8975 (N_8975,N_7342,N_7368);
nor U8976 (N_8976,N_7963,N_7556);
or U8977 (N_8977,N_7705,N_7664);
nand U8978 (N_8978,N_7491,N_7748);
nand U8979 (N_8979,N_7614,N_7369);
nor U8980 (N_8980,N_7546,N_7354);
nand U8981 (N_8981,N_7530,N_7774);
and U8982 (N_8982,N_7540,N_7924);
or U8983 (N_8983,N_7121,N_7896);
xnor U8984 (N_8984,N_7544,N_7967);
and U8985 (N_8985,N_7471,N_7414);
and U8986 (N_8986,N_7747,N_7946);
or U8987 (N_8987,N_7924,N_7158);
xnor U8988 (N_8988,N_7766,N_7776);
and U8989 (N_8989,N_7419,N_7915);
or U8990 (N_8990,N_7245,N_7946);
nand U8991 (N_8991,N_7608,N_7394);
nand U8992 (N_8992,N_7200,N_7144);
and U8993 (N_8993,N_7893,N_7535);
or U8994 (N_8994,N_7055,N_7026);
nand U8995 (N_8995,N_7553,N_7450);
xnor U8996 (N_8996,N_7519,N_7640);
xor U8997 (N_8997,N_7270,N_7143);
xor U8998 (N_8998,N_7943,N_7556);
nor U8999 (N_8999,N_7011,N_7215);
nand U9000 (N_9000,N_8892,N_8306);
xor U9001 (N_9001,N_8751,N_8449);
and U9002 (N_9002,N_8949,N_8832);
nor U9003 (N_9003,N_8473,N_8683);
nand U9004 (N_9004,N_8564,N_8695);
xor U9005 (N_9005,N_8617,N_8896);
xor U9006 (N_9006,N_8198,N_8092);
nand U9007 (N_9007,N_8062,N_8250);
xnor U9008 (N_9008,N_8681,N_8785);
xnor U9009 (N_9009,N_8304,N_8528);
nand U9010 (N_9010,N_8650,N_8270);
nand U9011 (N_9011,N_8706,N_8191);
nor U9012 (N_9012,N_8986,N_8041);
nand U9013 (N_9013,N_8374,N_8097);
xor U9014 (N_9014,N_8687,N_8063);
and U9015 (N_9015,N_8005,N_8997);
and U9016 (N_9016,N_8019,N_8794);
or U9017 (N_9017,N_8781,N_8939);
or U9018 (N_9018,N_8302,N_8548);
or U9019 (N_9019,N_8178,N_8396);
or U9020 (N_9020,N_8920,N_8287);
nand U9021 (N_9021,N_8932,N_8693);
nand U9022 (N_9022,N_8469,N_8973);
nor U9023 (N_9023,N_8242,N_8200);
nand U9024 (N_9024,N_8182,N_8740);
xnor U9025 (N_9025,N_8463,N_8582);
nor U9026 (N_9026,N_8749,N_8651);
nor U9027 (N_9027,N_8821,N_8587);
nand U9028 (N_9028,N_8883,N_8633);
nor U9029 (N_9029,N_8436,N_8635);
nand U9030 (N_9030,N_8642,N_8792);
nor U9031 (N_9031,N_8700,N_8671);
or U9032 (N_9032,N_8513,N_8991);
xor U9033 (N_9033,N_8666,N_8157);
nand U9034 (N_9034,N_8407,N_8456);
nand U9035 (N_9035,N_8047,N_8902);
xor U9036 (N_9036,N_8696,N_8723);
and U9037 (N_9037,N_8422,N_8112);
xor U9038 (N_9038,N_8232,N_8577);
nor U9039 (N_9039,N_8401,N_8917);
or U9040 (N_9040,N_8332,N_8544);
nor U9041 (N_9041,N_8527,N_8235);
xnor U9042 (N_9042,N_8234,N_8053);
xnor U9043 (N_9043,N_8095,N_8825);
nand U9044 (N_9044,N_8093,N_8835);
and U9045 (N_9045,N_8244,N_8017);
nor U9046 (N_9046,N_8934,N_8876);
or U9047 (N_9047,N_8299,N_8343);
and U9048 (N_9048,N_8219,N_8637);
and U9049 (N_9049,N_8614,N_8933);
and U9050 (N_9050,N_8579,N_8059);
nor U9051 (N_9051,N_8545,N_8950);
and U9052 (N_9052,N_8983,N_8073);
xor U9053 (N_9053,N_8368,N_8461);
nand U9054 (N_9054,N_8890,N_8521);
xnor U9055 (N_9055,N_8162,N_8455);
or U9056 (N_9056,N_8305,N_8793);
nor U9057 (N_9057,N_8638,N_8909);
xor U9058 (N_9058,N_8125,N_8111);
nor U9059 (N_9059,N_8546,N_8941);
xor U9060 (N_9060,N_8727,N_8013);
xor U9061 (N_9061,N_8877,N_8404);
xnor U9062 (N_9062,N_8926,N_8640);
nor U9063 (N_9063,N_8842,N_8854);
xor U9064 (N_9064,N_8836,N_8813);
or U9065 (N_9065,N_8300,N_8377);
or U9066 (N_9066,N_8493,N_8879);
and U9067 (N_9067,N_8143,N_8531);
nor U9068 (N_9068,N_8405,N_8946);
and U9069 (N_9069,N_8861,N_8598);
nand U9070 (N_9070,N_8601,N_8690);
xor U9071 (N_9071,N_8070,N_8606);
or U9072 (N_9072,N_8757,N_8057);
nor U9073 (N_9073,N_8938,N_8153);
nor U9074 (N_9074,N_8995,N_8196);
and U9075 (N_9075,N_8464,N_8336);
nand U9076 (N_9076,N_8241,N_8895);
or U9077 (N_9077,N_8290,N_8899);
xor U9078 (N_9078,N_8106,N_8963);
xnor U9079 (N_9079,N_8109,N_8312);
nand U9080 (N_9080,N_8383,N_8576);
xnor U9081 (N_9081,N_8662,N_8166);
or U9082 (N_9082,N_8308,N_8759);
and U9083 (N_9083,N_8978,N_8658);
nand U9084 (N_9084,N_8773,N_8929);
and U9085 (N_9085,N_8430,N_8453);
nor U9086 (N_9086,N_8316,N_8589);
and U9087 (N_9087,N_8348,N_8800);
nand U9088 (N_9088,N_8334,N_8071);
or U9089 (N_9089,N_8359,N_8210);
or U9090 (N_9090,N_8136,N_8209);
or U9091 (N_9091,N_8507,N_8502);
nand U9092 (N_9092,N_8037,N_8264);
and U9093 (N_9093,N_8889,N_8460);
or U9094 (N_9094,N_8903,N_8325);
nand U9095 (N_9095,N_8734,N_8815);
nor U9096 (N_9096,N_8742,N_8128);
or U9097 (N_9097,N_8568,N_8718);
nor U9098 (N_9098,N_8647,N_8271);
nor U9099 (N_9099,N_8443,N_8618);
or U9100 (N_9100,N_8959,N_8851);
or U9101 (N_9101,N_8186,N_8151);
and U9102 (N_9102,N_8323,N_8807);
and U9103 (N_9103,N_8943,N_8413);
or U9104 (N_9104,N_8195,N_8885);
or U9105 (N_9105,N_8893,N_8188);
or U9106 (N_9106,N_8697,N_8812);
nand U9107 (N_9107,N_8020,N_8014);
xnor U9108 (N_9108,N_8853,N_8044);
xnor U9109 (N_9109,N_8868,N_8620);
or U9110 (N_9110,N_8375,N_8703);
xor U9111 (N_9111,N_8680,N_8387);
or U9112 (N_9112,N_8600,N_8754);
nor U9113 (N_9113,N_8267,N_8714);
or U9114 (N_9114,N_8731,N_8272);
nand U9115 (N_9115,N_8243,N_8810);
xnor U9116 (N_9116,N_8038,N_8517);
nand U9117 (N_9117,N_8848,N_8801);
or U9118 (N_9118,N_8459,N_8849);
and U9119 (N_9119,N_8083,N_8645);
xnor U9120 (N_9120,N_8373,N_8948);
and U9121 (N_9121,N_8534,N_8841);
or U9122 (N_9122,N_8036,N_8284);
nor U9123 (N_9123,N_8427,N_8081);
or U9124 (N_9124,N_8538,N_8298);
or U9125 (N_9125,N_8656,N_8341);
or U9126 (N_9126,N_8878,N_8279);
nand U9127 (N_9127,N_8126,N_8079);
and U9128 (N_9128,N_8319,N_8864);
nor U9129 (N_9129,N_8722,N_8655);
nand U9130 (N_9130,N_8843,N_8424);
nor U9131 (N_9131,N_8385,N_8961);
nand U9132 (N_9132,N_8724,N_8953);
and U9133 (N_9133,N_8748,N_8468);
and U9134 (N_9134,N_8286,N_8314);
nand U9135 (N_9135,N_8924,N_8273);
or U9136 (N_9136,N_8212,N_8148);
xor U9137 (N_9137,N_8010,N_8355);
or U9138 (N_9138,N_8475,N_8543);
xnor U9139 (N_9139,N_8586,N_8599);
and U9140 (N_9140,N_8557,N_8756);
xor U9141 (N_9141,N_8729,N_8511);
xnor U9142 (N_9142,N_8964,N_8555);
nor U9143 (N_9143,N_8467,N_8347);
xnor U9144 (N_9144,N_8866,N_8872);
or U9145 (N_9145,N_8184,N_8985);
or U9146 (N_9146,N_8870,N_8281);
nor U9147 (N_9147,N_8803,N_8795);
nor U9148 (N_9148,N_8438,N_8124);
nand U9149 (N_9149,N_8674,N_8173);
nand U9150 (N_9150,N_8193,N_8726);
or U9151 (N_9151,N_8830,N_8445);
xnor U9152 (N_9152,N_8634,N_8448);
and U9153 (N_9153,N_8480,N_8536);
xor U9154 (N_9154,N_8139,N_8774);
xor U9155 (N_9155,N_8581,N_8412);
and U9156 (N_9156,N_8075,N_8560);
nor U9157 (N_9157,N_8747,N_8441);
or U9158 (N_9158,N_8657,N_8980);
nor U9159 (N_9159,N_8691,N_8022);
or U9160 (N_9160,N_8954,N_8979);
xor U9161 (N_9161,N_8216,N_8486);
or U9162 (N_9162,N_8055,N_8408);
nand U9163 (N_9163,N_8602,N_8146);
nor U9164 (N_9164,N_8624,N_8320);
and U9165 (N_9165,N_8942,N_8177);
or U9166 (N_9166,N_8156,N_8240);
xnor U9167 (N_9167,N_8894,N_8554);
and U9168 (N_9168,N_8023,N_8118);
nand U9169 (N_9169,N_8550,N_8931);
and U9170 (N_9170,N_8108,N_8969);
or U9171 (N_9171,N_8631,N_8252);
xor U9172 (N_9172,N_8491,N_8499);
nor U9173 (N_9173,N_8389,N_8831);
and U9174 (N_9174,N_8406,N_8575);
nand U9175 (N_9175,N_8990,N_8214);
nor U9176 (N_9176,N_8764,N_8914);
or U9177 (N_9177,N_8906,N_8551);
nor U9178 (N_9178,N_8409,N_8419);
nor U9179 (N_9179,N_8116,N_8294);
or U9180 (N_9180,N_8076,N_8838);
xnor U9181 (N_9181,N_8668,N_8477);
xnor U9182 (N_9182,N_8275,N_8457);
nand U9183 (N_9183,N_8621,N_8782);
nor U9184 (N_9184,N_8466,N_8494);
nand U9185 (N_9185,N_8113,N_8512);
and U9186 (N_9186,N_8537,N_8066);
xnor U9187 (N_9187,N_8094,N_8607);
nor U9188 (N_9188,N_8852,N_8172);
xor U9189 (N_9189,N_8552,N_8133);
nor U9190 (N_9190,N_8694,N_8261);
nand U9191 (N_9191,N_8940,N_8761);
nor U9192 (N_9192,N_8067,N_8826);
nand U9193 (N_9193,N_8102,N_8175);
nand U9194 (N_9194,N_8532,N_8205);
or U9195 (N_9195,N_8652,N_8391);
nor U9196 (N_9196,N_8002,N_8881);
nor U9197 (N_9197,N_8024,N_8622);
nand U9198 (N_9198,N_8790,N_8226);
xnor U9199 (N_9199,N_8705,N_8245);
or U9200 (N_9200,N_8603,N_8040);
or U9201 (N_9201,N_8288,N_8525);
xnor U9202 (N_9202,N_8266,N_8301);
nor U9203 (N_9203,N_8398,N_8702);
or U9204 (N_9204,N_8570,N_8123);
nand U9205 (N_9205,N_8716,N_8900);
or U9206 (N_9206,N_8916,N_8465);
xnor U9207 (N_9207,N_8356,N_8337);
xnor U9208 (N_9208,N_8256,N_8626);
xnor U9209 (N_9209,N_8488,N_8310);
and U9210 (N_9210,N_8016,N_8588);
or U9211 (N_9211,N_8721,N_8370);
and U9212 (N_9212,N_8130,N_8490);
nor U9213 (N_9213,N_8386,N_8770);
nor U9214 (N_9214,N_8686,N_8358);
xor U9215 (N_9215,N_8218,N_8414);
nor U9216 (N_9216,N_8547,N_8179);
nor U9217 (N_9217,N_8163,N_8048);
nand U9218 (N_9218,N_8679,N_8925);
and U9219 (N_9219,N_8935,N_8960);
nand U9220 (N_9220,N_8421,N_8875);
nand U9221 (N_9221,N_8354,N_8752);
or U9222 (N_9222,N_8955,N_8791);
xor U9223 (N_9223,N_8820,N_8280);
xnor U9224 (N_9224,N_8659,N_8152);
nor U9225 (N_9225,N_8766,N_8661);
and U9226 (N_9226,N_8224,N_8972);
nor U9227 (N_9227,N_8285,N_8796);
nand U9228 (N_9228,N_8771,N_8328);
nand U9229 (N_9229,N_8433,N_8390);
nor U9230 (N_9230,N_8091,N_8211);
nor U9231 (N_9231,N_8901,N_8372);
xnor U9232 (N_9232,N_8326,N_8003);
or U9233 (N_9233,N_8026,N_8236);
or U9234 (N_9234,N_8274,N_8199);
nor U9235 (N_9235,N_8594,N_8967);
nand U9236 (N_9236,N_8613,N_8886);
or U9237 (N_9237,N_8426,N_8452);
xnor U9238 (N_9238,N_8744,N_8444);
nand U9239 (N_9239,N_8431,N_8397);
nor U9240 (N_9240,N_8541,N_8789);
or U9241 (N_9241,N_8268,N_8471);
nor U9242 (N_9242,N_8450,N_8643);
and U9243 (N_9243,N_8117,N_8971);
xor U9244 (N_9244,N_8361,N_8228);
nand U9245 (N_9245,N_8104,N_8822);
and U9246 (N_9246,N_8446,N_8846);
xnor U9247 (N_9247,N_8798,N_8315);
nor U9248 (N_9248,N_8411,N_8293);
nand U9249 (N_9249,N_8107,N_8096);
or U9250 (N_9250,N_8018,N_8750);
or U9251 (N_9251,N_8768,N_8025);
or U9252 (N_9252,N_8031,N_8612);
and U9253 (N_9253,N_8987,N_8335);
and U9254 (N_9254,N_8699,N_8054);
xor U9255 (N_9255,N_8043,N_8912);
xnor U9256 (N_9256,N_8180,N_8231);
nor U9257 (N_9257,N_8833,N_8167);
and U9258 (N_9258,N_8871,N_8251);
and U9259 (N_9259,N_8585,N_8654);
or U9260 (N_9260,N_8454,N_8384);
or U9261 (N_9261,N_8636,N_8297);
nor U9262 (N_9262,N_8767,N_8844);
nor U9263 (N_9263,N_8197,N_8291);
nor U9264 (N_9264,N_8145,N_8246);
nor U9265 (N_9265,N_8573,N_8056);
nand U9266 (N_9266,N_8738,N_8530);
nand U9267 (N_9267,N_8503,N_8239);
nand U9268 (N_9268,N_8510,N_8590);
nand U9269 (N_9269,N_8762,N_8616);
nand U9270 (N_9270,N_8007,N_8410);
or U9271 (N_9271,N_8141,N_8930);
or U9272 (N_9272,N_8827,N_8262);
nand U9273 (N_9273,N_8451,N_8192);
or U9274 (N_9274,N_8887,N_8526);
nand U9275 (N_9275,N_8159,N_8313);
xor U9276 (N_9276,N_8565,N_8556);
or U9277 (N_9277,N_8364,N_8127);
xnor U9278 (N_9278,N_8730,N_8028);
nor U9279 (N_9279,N_8278,N_8665);
or U9280 (N_9280,N_8672,N_8630);
and U9281 (N_9281,N_8098,N_8580);
nor U9282 (N_9282,N_8033,N_8470);
xnor U9283 (N_9283,N_8458,N_8004);
and U9284 (N_9284,N_8728,N_8859);
or U9285 (N_9285,N_8623,N_8927);
or U9286 (N_9286,N_8149,N_8763);
and U9287 (N_9287,N_8011,N_8677);
nor U9288 (N_9288,N_8185,N_8360);
nand U9289 (N_9289,N_8506,N_8263);
xnor U9290 (N_9290,N_8296,N_8918);
nor U9291 (N_9291,N_8171,N_8514);
nor U9292 (N_9292,N_8090,N_8176);
nor U9293 (N_9293,N_8222,N_8150);
nor U9294 (N_9294,N_8984,N_8735);
xor U9295 (N_9295,N_8968,N_8524);
or U9296 (N_9296,N_8440,N_8061);
xnor U9297 (N_9297,N_8787,N_8559);
xor U9298 (N_9298,N_8709,N_8435);
xnor U9299 (N_9299,N_8114,N_8799);
or U9300 (N_9300,N_8676,N_8566);
nor U9301 (N_9301,N_8840,N_8845);
and U9302 (N_9302,N_8808,N_8476);
xnor U9303 (N_9303,N_8804,N_8688);
nand U9304 (N_9304,N_8283,N_8160);
nor U9305 (N_9305,N_8684,N_8472);
or U9306 (N_9306,N_8567,N_8847);
xor U9307 (N_9307,N_8778,N_8190);
xnor U9308 (N_9308,N_8753,N_8746);
and U9309 (N_9309,N_8223,N_8339);
or U9310 (N_9310,N_8068,N_8553);
nor U9311 (N_9311,N_8225,N_8673);
nor U9312 (N_9312,N_8535,N_8998);
nand U9313 (N_9313,N_8921,N_8788);
nor U9314 (N_9314,N_8089,N_8784);
xnor U9315 (N_9315,N_8257,N_8561);
xor U9316 (N_9316,N_8563,N_8233);
nor U9317 (N_9317,N_8518,N_8505);
and U9318 (N_9318,N_8936,N_8860);
xnor U9319 (N_9319,N_8610,N_8189);
nor U9320 (N_9320,N_8131,N_8378);
and U9321 (N_9321,N_8739,N_8873);
or U9322 (N_9322,N_8487,N_8164);
and U9323 (N_9323,N_8479,N_8649);
and U9324 (N_9324,N_8769,N_8856);
or U9325 (N_9325,N_8583,N_8380);
nand U9326 (N_9326,N_8099,N_8717);
nand U9327 (N_9327,N_8947,N_8110);
or U9328 (N_9328,N_8646,N_8229);
nor U9329 (N_9329,N_8072,N_8701);
nand U9330 (N_9330,N_8327,N_8147);
or U9331 (N_9331,N_8277,N_8819);
nor U9332 (N_9332,N_8282,N_8692);
or U9333 (N_9333,N_8032,N_8342);
nand U9334 (N_9334,N_8169,N_8140);
and U9335 (N_9335,N_8549,N_8006);
and U9336 (N_9336,N_8806,N_8663);
or U9337 (N_9337,N_8416,N_8352);
and U9338 (N_9338,N_8562,N_8289);
nand U9339 (N_9339,N_8082,N_8481);
xor U9340 (N_9340,N_8247,N_8904);
xor U9341 (N_9341,N_8857,N_8042);
nor U9342 (N_9342,N_8230,N_8138);
nand U9343 (N_9343,N_8824,N_8227);
nand U9344 (N_9344,N_8758,N_8132);
nor U9345 (N_9345,N_8818,N_8086);
nand U9346 (N_9346,N_8330,N_8639);
nor U9347 (N_9347,N_8863,N_8797);
and U9348 (N_9348,N_8064,N_8595);
xnor U9349 (N_9349,N_8371,N_8194);
nand U9350 (N_9350,N_8447,N_8707);
nor U9351 (N_9351,N_8351,N_8689);
nand U9352 (N_9352,N_8321,N_8501);
nor U9353 (N_9353,N_8989,N_8345);
nand U9354 (N_9354,N_8204,N_8392);
or U9355 (N_9355,N_8923,N_8121);
xnor U9356 (N_9356,N_8678,N_8399);
nand U9357 (N_9357,N_8829,N_8255);
nor U9358 (N_9358,N_8496,N_8988);
and U9359 (N_9359,N_8974,N_8322);
xnor U9360 (N_9360,N_8382,N_8737);
or U9361 (N_9361,N_8970,N_8779);
xor U9362 (N_9362,N_8303,N_8039);
nor U9363 (N_9363,N_8344,N_8571);
and U9364 (N_9364,N_8908,N_8533);
xnor U9365 (N_9365,N_8331,N_8509);
and U9366 (N_9366,N_8937,N_8403);
nand U9367 (N_9367,N_8596,N_8253);
and U9368 (N_9368,N_8858,N_8052);
nor U9369 (N_9369,N_8837,N_8945);
nand U9370 (N_9370,N_8708,N_8615);
nor U9371 (N_9371,N_8119,N_8009);
or U9372 (N_9372,N_8206,N_8485);
nor U9373 (N_9373,N_8393,N_8442);
and U9374 (N_9374,N_8743,N_8168);
or U9375 (N_9375,N_8736,N_8495);
xor U9376 (N_9376,N_8357,N_8627);
nor U9377 (N_9377,N_8604,N_8880);
and U9378 (N_9378,N_8249,N_8338);
or U9379 (N_9379,N_8202,N_8962);
or U9380 (N_9380,N_8597,N_8346);
and U9381 (N_9381,N_8425,N_8775);
or U9382 (N_9382,N_8994,N_8855);
or U9383 (N_9383,N_8423,N_8976);
xnor U9384 (N_9384,N_8155,N_8350);
nand U9385 (N_9385,N_8215,N_8910);
and U9386 (N_9386,N_8482,N_8725);
nand U9387 (N_9387,N_8713,N_8569);
or U9388 (N_9388,N_8664,N_8578);
and U9389 (N_9389,N_8915,N_8777);
nand U9390 (N_9390,N_8432,N_8307);
nand U9391 (N_9391,N_8258,N_8429);
or U9392 (N_9392,N_8213,N_8891);
or U9393 (N_9393,N_8698,N_8760);
xnor U9394 (N_9394,N_8591,N_8035);
nor U9395 (N_9395,N_8966,N_8237);
or U9396 (N_9396,N_8492,N_8888);
and U9397 (N_9397,N_8669,N_8520);
or U9398 (N_9398,N_8394,N_8478);
xor U9399 (N_9399,N_8958,N_8489);
xnor U9400 (N_9400,N_8366,N_8221);
and U9401 (N_9401,N_8074,N_8522);
nand U9402 (N_9402,N_8982,N_8865);
and U9403 (N_9403,N_8008,N_8077);
xor U9404 (N_9404,N_8653,N_8780);
nor U9405 (N_9405,N_8203,N_8165);
nor U9406 (N_9406,N_8000,N_8952);
and U9407 (N_9407,N_8483,N_8720);
or U9408 (N_9408,N_8080,N_8154);
nand U9409 (N_9409,N_8816,N_8572);
or U9410 (N_9410,N_8012,N_8592);
and U9411 (N_9411,N_8542,N_8474);
and U9412 (N_9412,N_8814,N_8101);
nor U9413 (N_9413,N_8437,N_8874);
and U9414 (N_9414,N_8975,N_8122);
xnor U9415 (N_9415,N_8869,N_8135);
xor U9416 (N_9416,N_8719,N_8276);
nor U9417 (N_9417,N_8120,N_8292);
or U9418 (N_9418,N_8508,N_8611);
nor U9419 (N_9419,N_8088,N_8993);
nand U9420 (N_9420,N_8540,N_8484);
and U9421 (N_9421,N_8641,N_8644);
and U9422 (N_9422,N_8772,N_8977);
nor U9423 (N_9423,N_8897,N_8755);
nand U9424 (N_9424,N_8439,N_8965);
nand U9425 (N_9425,N_8265,N_8884);
and U9426 (N_9426,N_8828,N_8428);
nand U9427 (N_9427,N_8882,N_8065);
xnor U9428 (N_9428,N_8129,N_8029);
or U9429 (N_9429,N_8158,N_8001);
and U9430 (N_9430,N_8625,N_8311);
or U9431 (N_9431,N_8103,N_8183);
or U9432 (N_9432,N_8238,N_8648);
and U9433 (N_9433,N_8682,N_8632);
nor U9434 (N_9434,N_8395,N_8504);
nand U9435 (N_9435,N_8660,N_8809);
and U9436 (N_9436,N_8021,N_8802);
nor U9437 (N_9437,N_8418,N_8161);
xor U9438 (N_9438,N_8134,N_8174);
and U9439 (N_9439,N_8850,N_8497);
xor U9440 (N_9440,N_8996,N_8862);
xnor U9441 (N_9441,N_8898,N_8957);
xor U9442 (N_9442,N_8050,N_8379);
nand U9443 (N_9443,N_8628,N_8919);
nor U9444 (N_9444,N_8115,N_8402);
xor U9445 (N_9445,N_8100,N_8907);
or U9446 (N_9446,N_8049,N_8711);
or U9447 (N_9447,N_8187,N_8034);
or U9448 (N_9448,N_8619,N_8685);
xnor U9449 (N_9449,N_8732,N_8201);
nand U9450 (N_9450,N_8295,N_8805);
xor U9451 (N_9451,N_8259,N_8367);
and U9452 (N_9452,N_8170,N_8704);
and U9453 (N_9453,N_8733,N_8523);
nor U9454 (N_9454,N_8105,N_8811);
or U9455 (N_9455,N_8329,N_8928);
or U9456 (N_9456,N_8333,N_8539);
nand U9457 (N_9457,N_8715,N_8922);
xnor U9458 (N_9458,N_8269,N_8516);
nor U9459 (N_9459,N_8519,N_8388);
nand U9460 (N_9460,N_8207,N_8051);
xor U9461 (N_9461,N_8498,N_8400);
xor U9462 (N_9462,N_8605,N_8670);
nor U9463 (N_9463,N_8058,N_8045);
nand U9464 (N_9464,N_8944,N_8363);
nor U9465 (N_9465,N_8584,N_8085);
and U9466 (N_9466,N_8667,N_8992);
nand U9467 (N_9467,N_8434,N_8783);
xnor U9468 (N_9468,N_8208,N_8069);
or U9469 (N_9469,N_8254,N_8362);
nand U9470 (N_9470,N_8309,N_8027);
nor U9471 (N_9471,N_8317,N_8248);
xor U9472 (N_9472,N_8324,N_8905);
xnor U9473 (N_9473,N_8220,N_8765);
and U9474 (N_9474,N_8381,N_8745);
or U9475 (N_9475,N_8349,N_8817);
xor U9476 (N_9476,N_8629,N_8999);
nor U9477 (N_9477,N_8675,N_8078);
nor U9478 (N_9478,N_8217,N_8913);
nor U9479 (N_9479,N_8608,N_8529);
nand U9480 (N_9480,N_8376,N_8369);
and U9481 (N_9481,N_8839,N_8318);
and U9482 (N_9482,N_8981,N_8340);
or U9483 (N_9483,N_8951,N_8181);
nor U9484 (N_9484,N_8741,N_8500);
nand U9485 (N_9485,N_8030,N_8515);
and U9486 (N_9486,N_8415,N_8574);
xor U9487 (N_9487,N_8710,N_8558);
nor U9488 (N_9488,N_8593,N_8911);
or U9489 (N_9489,N_8087,N_8365);
and U9490 (N_9490,N_8823,N_8712);
nor U9491 (N_9491,N_8015,N_8144);
and U9492 (N_9492,N_8137,N_8786);
xnor U9493 (N_9493,N_8420,N_8046);
and U9494 (N_9494,N_8084,N_8776);
nand U9495 (N_9495,N_8260,N_8609);
nand U9496 (N_9496,N_8060,N_8462);
xor U9497 (N_9497,N_8867,N_8834);
and U9498 (N_9498,N_8353,N_8142);
nor U9499 (N_9499,N_8417,N_8956);
nand U9500 (N_9500,N_8997,N_8804);
xor U9501 (N_9501,N_8774,N_8056);
or U9502 (N_9502,N_8578,N_8937);
and U9503 (N_9503,N_8798,N_8250);
or U9504 (N_9504,N_8223,N_8328);
or U9505 (N_9505,N_8227,N_8619);
xor U9506 (N_9506,N_8458,N_8154);
or U9507 (N_9507,N_8030,N_8500);
or U9508 (N_9508,N_8744,N_8165);
nand U9509 (N_9509,N_8016,N_8218);
or U9510 (N_9510,N_8647,N_8499);
xnor U9511 (N_9511,N_8149,N_8050);
nand U9512 (N_9512,N_8090,N_8991);
or U9513 (N_9513,N_8801,N_8216);
nor U9514 (N_9514,N_8457,N_8672);
and U9515 (N_9515,N_8104,N_8835);
nor U9516 (N_9516,N_8896,N_8217);
nand U9517 (N_9517,N_8596,N_8493);
nor U9518 (N_9518,N_8938,N_8145);
nand U9519 (N_9519,N_8214,N_8782);
or U9520 (N_9520,N_8627,N_8904);
nand U9521 (N_9521,N_8662,N_8400);
nor U9522 (N_9522,N_8897,N_8450);
or U9523 (N_9523,N_8569,N_8626);
nand U9524 (N_9524,N_8616,N_8401);
xnor U9525 (N_9525,N_8516,N_8189);
xor U9526 (N_9526,N_8550,N_8084);
nor U9527 (N_9527,N_8253,N_8766);
or U9528 (N_9528,N_8906,N_8752);
xor U9529 (N_9529,N_8678,N_8189);
xnor U9530 (N_9530,N_8079,N_8986);
or U9531 (N_9531,N_8874,N_8214);
nand U9532 (N_9532,N_8692,N_8054);
and U9533 (N_9533,N_8595,N_8383);
nor U9534 (N_9534,N_8936,N_8459);
nor U9535 (N_9535,N_8389,N_8197);
xnor U9536 (N_9536,N_8382,N_8485);
or U9537 (N_9537,N_8024,N_8843);
or U9538 (N_9538,N_8337,N_8008);
or U9539 (N_9539,N_8131,N_8021);
nor U9540 (N_9540,N_8798,N_8875);
or U9541 (N_9541,N_8701,N_8643);
nand U9542 (N_9542,N_8172,N_8352);
xor U9543 (N_9543,N_8109,N_8803);
xor U9544 (N_9544,N_8511,N_8346);
and U9545 (N_9545,N_8054,N_8032);
xor U9546 (N_9546,N_8128,N_8762);
nand U9547 (N_9547,N_8414,N_8108);
nand U9548 (N_9548,N_8707,N_8652);
or U9549 (N_9549,N_8021,N_8301);
and U9550 (N_9550,N_8663,N_8715);
xnor U9551 (N_9551,N_8304,N_8481);
nor U9552 (N_9552,N_8956,N_8882);
or U9553 (N_9553,N_8419,N_8806);
nand U9554 (N_9554,N_8821,N_8028);
nand U9555 (N_9555,N_8864,N_8151);
nand U9556 (N_9556,N_8862,N_8509);
nor U9557 (N_9557,N_8072,N_8394);
xnor U9558 (N_9558,N_8494,N_8170);
xnor U9559 (N_9559,N_8020,N_8873);
nor U9560 (N_9560,N_8751,N_8272);
or U9561 (N_9561,N_8470,N_8482);
nand U9562 (N_9562,N_8644,N_8774);
nor U9563 (N_9563,N_8277,N_8740);
nor U9564 (N_9564,N_8733,N_8592);
nor U9565 (N_9565,N_8119,N_8042);
nand U9566 (N_9566,N_8452,N_8759);
nor U9567 (N_9567,N_8248,N_8407);
nand U9568 (N_9568,N_8096,N_8766);
and U9569 (N_9569,N_8142,N_8998);
nand U9570 (N_9570,N_8885,N_8917);
and U9571 (N_9571,N_8792,N_8461);
nor U9572 (N_9572,N_8808,N_8431);
or U9573 (N_9573,N_8249,N_8876);
and U9574 (N_9574,N_8874,N_8326);
xor U9575 (N_9575,N_8961,N_8443);
nor U9576 (N_9576,N_8513,N_8160);
xor U9577 (N_9577,N_8065,N_8709);
nor U9578 (N_9578,N_8709,N_8329);
or U9579 (N_9579,N_8187,N_8915);
nand U9580 (N_9580,N_8174,N_8784);
xnor U9581 (N_9581,N_8203,N_8155);
xor U9582 (N_9582,N_8400,N_8996);
or U9583 (N_9583,N_8400,N_8057);
xor U9584 (N_9584,N_8362,N_8524);
nor U9585 (N_9585,N_8755,N_8708);
nand U9586 (N_9586,N_8168,N_8412);
nand U9587 (N_9587,N_8028,N_8681);
nor U9588 (N_9588,N_8731,N_8194);
xnor U9589 (N_9589,N_8674,N_8309);
nor U9590 (N_9590,N_8761,N_8251);
and U9591 (N_9591,N_8409,N_8786);
xor U9592 (N_9592,N_8319,N_8541);
or U9593 (N_9593,N_8845,N_8129);
nand U9594 (N_9594,N_8040,N_8884);
or U9595 (N_9595,N_8538,N_8632);
or U9596 (N_9596,N_8599,N_8011);
or U9597 (N_9597,N_8476,N_8676);
xor U9598 (N_9598,N_8886,N_8684);
and U9599 (N_9599,N_8139,N_8606);
xnor U9600 (N_9600,N_8970,N_8473);
xor U9601 (N_9601,N_8571,N_8040);
and U9602 (N_9602,N_8318,N_8262);
and U9603 (N_9603,N_8477,N_8399);
xnor U9604 (N_9604,N_8187,N_8425);
nor U9605 (N_9605,N_8069,N_8820);
and U9606 (N_9606,N_8660,N_8186);
and U9607 (N_9607,N_8503,N_8364);
or U9608 (N_9608,N_8505,N_8982);
nand U9609 (N_9609,N_8797,N_8216);
or U9610 (N_9610,N_8569,N_8042);
xor U9611 (N_9611,N_8641,N_8778);
or U9612 (N_9612,N_8573,N_8232);
nand U9613 (N_9613,N_8234,N_8571);
nand U9614 (N_9614,N_8741,N_8972);
nand U9615 (N_9615,N_8213,N_8845);
xnor U9616 (N_9616,N_8597,N_8184);
or U9617 (N_9617,N_8205,N_8520);
nand U9618 (N_9618,N_8375,N_8567);
and U9619 (N_9619,N_8340,N_8310);
xnor U9620 (N_9620,N_8451,N_8363);
or U9621 (N_9621,N_8498,N_8495);
nor U9622 (N_9622,N_8230,N_8845);
nor U9623 (N_9623,N_8416,N_8879);
or U9624 (N_9624,N_8868,N_8584);
and U9625 (N_9625,N_8078,N_8602);
nand U9626 (N_9626,N_8417,N_8759);
xnor U9627 (N_9627,N_8521,N_8787);
nand U9628 (N_9628,N_8715,N_8368);
or U9629 (N_9629,N_8851,N_8343);
or U9630 (N_9630,N_8882,N_8891);
nand U9631 (N_9631,N_8921,N_8138);
xor U9632 (N_9632,N_8402,N_8576);
and U9633 (N_9633,N_8597,N_8228);
or U9634 (N_9634,N_8791,N_8506);
nor U9635 (N_9635,N_8973,N_8697);
and U9636 (N_9636,N_8869,N_8550);
xnor U9637 (N_9637,N_8310,N_8040);
and U9638 (N_9638,N_8450,N_8508);
xor U9639 (N_9639,N_8891,N_8562);
xnor U9640 (N_9640,N_8894,N_8514);
nor U9641 (N_9641,N_8234,N_8082);
nor U9642 (N_9642,N_8712,N_8031);
xnor U9643 (N_9643,N_8920,N_8394);
or U9644 (N_9644,N_8440,N_8590);
or U9645 (N_9645,N_8669,N_8853);
xor U9646 (N_9646,N_8026,N_8845);
nand U9647 (N_9647,N_8372,N_8760);
nand U9648 (N_9648,N_8449,N_8536);
xnor U9649 (N_9649,N_8122,N_8558);
xor U9650 (N_9650,N_8238,N_8764);
and U9651 (N_9651,N_8211,N_8494);
nor U9652 (N_9652,N_8381,N_8014);
nand U9653 (N_9653,N_8876,N_8642);
xor U9654 (N_9654,N_8244,N_8684);
nand U9655 (N_9655,N_8159,N_8125);
and U9656 (N_9656,N_8063,N_8157);
xor U9657 (N_9657,N_8710,N_8891);
nand U9658 (N_9658,N_8610,N_8268);
nand U9659 (N_9659,N_8534,N_8701);
nor U9660 (N_9660,N_8739,N_8316);
nor U9661 (N_9661,N_8751,N_8131);
or U9662 (N_9662,N_8765,N_8659);
nand U9663 (N_9663,N_8569,N_8889);
nor U9664 (N_9664,N_8738,N_8933);
and U9665 (N_9665,N_8425,N_8022);
xor U9666 (N_9666,N_8652,N_8341);
or U9667 (N_9667,N_8849,N_8490);
nor U9668 (N_9668,N_8999,N_8107);
xor U9669 (N_9669,N_8763,N_8889);
or U9670 (N_9670,N_8057,N_8277);
xnor U9671 (N_9671,N_8233,N_8508);
xor U9672 (N_9672,N_8746,N_8064);
nor U9673 (N_9673,N_8621,N_8134);
or U9674 (N_9674,N_8203,N_8681);
xor U9675 (N_9675,N_8650,N_8368);
nor U9676 (N_9676,N_8680,N_8257);
and U9677 (N_9677,N_8256,N_8705);
nand U9678 (N_9678,N_8158,N_8086);
nand U9679 (N_9679,N_8059,N_8839);
or U9680 (N_9680,N_8387,N_8793);
and U9681 (N_9681,N_8160,N_8381);
nand U9682 (N_9682,N_8441,N_8000);
or U9683 (N_9683,N_8267,N_8936);
or U9684 (N_9684,N_8949,N_8997);
xnor U9685 (N_9685,N_8210,N_8905);
nand U9686 (N_9686,N_8334,N_8504);
and U9687 (N_9687,N_8441,N_8576);
and U9688 (N_9688,N_8898,N_8674);
and U9689 (N_9689,N_8875,N_8033);
or U9690 (N_9690,N_8648,N_8447);
and U9691 (N_9691,N_8768,N_8679);
xor U9692 (N_9692,N_8177,N_8085);
nand U9693 (N_9693,N_8941,N_8639);
or U9694 (N_9694,N_8269,N_8104);
xor U9695 (N_9695,N_8872,N_8264);
nor U9696 (N_9696,N_8606,N_8333);
xor U9697 (N_9697,N_8068,N_8256);
and U9698 (N_9698,N_8540,N_8702);
xnor U9699 (N_9699,N_8427,N_8750);
nor U9700 (N_9700,N_8039,N_8963);
xor U9701 (N_9701,N_8137,N_8469);
nand U9702 (N_9702,N_8355,N_8636);
nand U9703 (N_9703,N_8328,N_8637);
nor U9704 (N_9704,N_8120,N_8488);
and U9705 (N_9705,N_8957,N_8661);
nand U9706 (N_9706,N_8964,N_8045);
and U9707 (N_9707,N_8513,N_8654);
or U9708 (N_9708,N_8307,N_8535);
nand U9709 (N_9709,N_8437,N_8579);
and U9710 (N_9710,N_8678,N_8522);
and U9711 (N_9711,N_8963,N_8879);
or U9712 (N_9712,N_8956,N_8741);
and U9713 (N_9713,N_8082,N_8337);
or U9714 (N_9714,N_8921,N_8839);
nand U9715 (N_9715,N_8501,N_8824);
nor U9716 (N_9716,N_8050,N_8078);
nand U9717 (N_9717,N_8901,N_8025);
nand U9718 (N_9718,N_8762,N_8866);
and U9719 (N_9719,N_8151,N_8885);
xnor U9720 (N_9720,N_8377,N_8624);
nand U9721 (N_9721,N_8175,N_8525);
nor U9722 (N_9722,N_8681,N_8489);
nor U9723 (N_9723,N_8997,N_8090);
xor U9724 (N_9724,N_8119,N_8018);
nor U9725 (N_9725,N_8848,N_8283);
xor U9726 (N_9726,N_8532,N_8865);
nand U9727 (N_9727,N_8502,N_8136);
or U9728 (N_9728,N_8793,N_8719);
or U9729 (N_9729,N_8853,N_8968);
xor U9730 (N_9730,N_8705,N_8624);
and U9731 (N_9731,N_8716,N_8760);
nor U9732 (N_9732,N_8201,N_8728);
nand U9733 (N_9733,N_8133,N_8742);
nor U9734 (N_9734,N_8293,N_8235);
nor U9735 (N_9735,N_8397,N_8079);
nand U9736 (N_9736,N_8410,N_8612);
nor U9737 (N_9737,N_8037,N_8024);
nor U9738 (N_9738,N_8687,N_8796);
xnor U9739 (N_9739,N_8672,N_8287);
or U9740 (N_9740,N_8417,N_8173);
nor U9741 (N_9741,N_8281,N_8139);
xnor U9742 (N_9742,N_8003,N_8636);
nor U9743 (N_9743,N_8066,N_8471);
xor U9744 (N_9744,N_8478,N_8387);
nor U9745 (N_9745,N_8051,N_8806);
nor U9746 (N_9746,N_8890,N_8418);
xor U9747 (N_9747,N_8587,N_8658);
xnor U9748 (N_9748,N_8285,N_8765);
xnor U9749 (N_9749,N_8107,N_8193);
or U9750 (N_9750,N_8782,N_8334);
nor U9751 (N_9751,N_8174,N_8800);
xor U9752 (N_9752,N_8785,N_8277);
and U9753 (N_9753,N_8474,N_8397);
or U9754 (N_9754,N_8079,N_8478);
and U9755 (N_9755,N_8257,N_8777);
nand U9756 (N_9756,N_8233,N_8417);
xnor U9757 (N_9757,N_8594,N_8220);
nor U9758 (N_9758,N_8562,N_8107);
nor U9759 (N_9759,N_8149,N_8744);
nand U9760 (N_9760,N_8151,N_8111);
and U9761 (N_9761,N_8718,N_8225);
xnor U9762 (N_9762,N_8267,N_8734);
or U9763 (N_9763,N_8793,N_8929);
and U9764 (N_9764,N_8524,N_8913);
xnor U9765 (N_9765,N_8903,N_8691);
xnor U9766 (N_9766,N_8917,N_8566);
xnor U9767 (N_9767,N_8473,N_8078);
nor U9768 (N_9768,N_8408,N_8058);
or U9769 (N_9769,N_8806,N_8128);
or U9770 (N_9770,N_8189,N_8121);
nor U9771 (N_9771,N_8165,N_8592);
and U9772 (N_9772,N_8904,N_8579);
nand U9773 (N_9773,N_8180,N_8868);
and U9774 (N_9774,N_8074,N_8142);
xor U9775 (N_9775,N_8620,N_8534);
nand U9776 (N_9776,N_8314,N_8019);
nor U9777 (N_9777,N_8776,N_8525);
xnor U9778 (N_9778,N_8618,N_8625);
nor U9779 (N_9779,N_8149,N_8778);
nand U9780 (N_9780,N_8571,N_8282);
or U9781 (N_9781,N_8323,N_8894);
and U9782 (N_9782,N_8421,N_8474);
or U9783 (N_9783,N_8066,N_8053);
or U9784 (N_9784,N_8460,N_8823);
nor U9785 (N_9785,N_8171,N_8524);
and U9786 (N_9786,N_8526,N_8725);
and U9787 (N_9787,N_8586,N_8005);
and U9788 (N_9788,N_8623,N_8224);
xnor U9789 (N_9789,N_8900,N_8535);
xor U9790 (N_9790,N_8341,N_8022);
and U9791 (N_9791,N_8107,N_8055);
or U9792 (N_9792,N_8862,N_8089);
xor U9793 (N_9793,N_8161,N_8130);
xor U9794 (N_9794,N_8048,N_8530);
and U9795 (N_9795,N_8837,N_8666);
nand U9796 (N_9796,N_8743,N_8365);
nand U9797 (N_9797,N_8125,N_8656);
and U9798 (N_9798,N_8877,N_8932);
or U9799 (N_9799,N_8898,N_8739);
nand U9800 (N_9800,N_8042,N_8070);
and U9801 (N_9801,N_8216,N_8195);
nand U9802 (N_9802,N_8989,N_8915);
nor U9803 (N_9803,N_8938,N_8761);
xnor U9804 (N_9804,N_8261,N_8431);
or U9805 (N_9805,N_8328,N_8931);
and U9806 (N_9806,N_8685,N_8938);
nand U9807 (N_9807,N_8287,N_8909);
and U9808 (N_9808,N_8973,N_8507);
and U9809 (N_9809,N_8662,N_8900);
xor U9810 (N_9810,N_8469,N_8212);
or U9811 (N_9811,N_8440,N_8529);
nand U9812 (N_9812,N_8724,N_8001);
nand U9813 (N_9813,N_8729,N_8711);
nor U9814 (N_9814,N_8700,N_8839);
xnor U9815 (N_9815,N_8060,N_8147);
nand U9816 (N_9816,N_8266,N_8651);
nand U9817 (N_9817,N_8890,N_8493);
or U9818 (N_9818,N_8789,N_8465);
or U9819 (N_9819,N_8709,N_8152);
nand U9820 (N_9820,N_8670,N_8386);
and U9821 (N_9821,N_8447,N_8467);
nor U9822 (N_9822,N_8096,N_8618);
nor U9823 (N_9823,N_8694,N_8345);
nand U9824 (N_9824,N_8690,N_8190);
nor U9825 (N_9825,N_8909,N_8992);
nand U9826 (N_9826,N_8826,N_8137);
xor U9827 (N_9827,N_8058,N_8332);
and U9828 (N_9828,N_8634,N_8931);
xnor U9829 (N_9829,N_8628,N_8744);
and U9830 (N_9830,N_8348,N_8626);
nand U9831 (N_9831,N_8329,N_8179);
or U9832 (N_9832,N_8937,N_8365);
or U9833 (N_9833,N_8457,N_8145);
xor U9834 (N_9834,N_8735,N_8229);
nand U9835 (N_9835,N_8161,N_8169);
and U9836 (N_9836,N_8021,N_8917);
xor U9837 (N_9837,N_8373,N_8037);
nand U9838 (N_9838,N_8794,N_8833);
nor U9839 (N_9839,N_8828,N_8844);
xor U9840 (N_9840,N_8928,N_8848);
nand U9841 (N_9841,N_8000,N_8308);
or U9842 (N_9842,N_8577,N_8510);
or U9843 (N_9843,N_8020,N_8955);
or U9844 (N_9844,N_8667,N_8618);
xor U9845 (N_9845,N_8131,N_8424);
and U9846 (N_9846,N_8182,N_8355);
and U9847 (N_9847,N_8860,N_8310);
or U9848 (N_9848,N_8879,N_8298);
and U9849 (N_9849,N_8260,N_8662);
nor U9850 (N_9850,N_8379,N_8191);
and U9851 (N_9851,N_8654,N_8828);
or U9852 (N_9852,N_8231,N_8234);
xor U9853 (N_9853,N_8887,N_8320);
and U9854 (N_9854,N_8714,N_8653);
nor U9855 (N_9855,N_8961,N_8538);
nor U9856 (N_9856,N_8400,N_8834);
xnor U9857 (N_9857,N_8557,N_8056);
or U9858 (N_9858,N_8655,N_8142);
or U9859 (N_9859,N_8694,N_8691);
xnor U9860 (N_9860,N_8314,N_8352);
nor U9861 (N_9861,N_8807,N_8503);
nand U9862 (N_9862,N_8103,N_8875);
xnor U9863 (N_9863,N_8734,N_8962);
xnor U9864 (N_9864,N_8871,N_8393);
and U9865 (N_9865,N_8406,N_8907);
nand U9866 (N_9866,N_8659,N_8726);
nand U9867 (N_9867,N_8060,N_8934);
xnor U9868 (N_9868,N_8813,N_8500);
xor U9869 (N_9869,N_8444,N_8680);
nor U9870 (N_9870,N_8068,N_8657);
nor U9871 (N_9871,N_8857,N_8600);
or U9872 (N_9872,N_8827,N_8976);
or U9873 (N_9873,N_8582,N_8014);
and U9874 (N_9874,N_8287,N_8330);
and U9875 (N_9875,N_8651,N_8002);
nand U9876 (N_9876,N_8070,N_8694);
and U9877 (N_9877,N_8701,N_8438);
xor U9878 (N_9878,N_8353,N_8709);
xor U9879 (N_9879,N_8129,N_8031);
and U9880 (N_9880,N_8835,N_8377);
nor U9881 (N_9881,N_8843,N_8949);
or U9882 (N_9882,N_8409,N_8260);
xnor U9883 (N_9883,N_8088,N_8685);
and U9884 (N_9884,N_8400,N_8109);
nor U9885 (N_9885,N_8883,N_8065);
xor U9886 (N_9886,N_8648,N_8069);
and U9887 (N_9887,N_8779,N_8221);
nand U9888 (N_9888,N_8590,N_8111);
and U9889 (N_9889,N_8460,N_8893);
nor U9890 (N_9890,N_8435,N_8512);
nand U9891 (N_9891,N_8800,N_8776);
nor U9892 (N_9892,N_8914,N_8801);
nor U9893 (N_9893,N_8850,N_8657);
and U9894 (N_9894,N_8354,N_8026);
or U9895 (N_9895,N_8006,N_8379);
nand U9896 (N_9896,N_8257,N_8352);
nand U9897 (N_9897,N_8791,N_8596);
and U9898 (N_9898,N_8199,N_8561);
xor U9899 (N_9899,N_8856,N_8246);
or U9900 (N_9900,N_8285,N_8279);
or U9901 (N_9901,N_8905,N_8719);
and U9902 (N_9902,N_8046,N_8821);
and U9903 (N_9903,N_8041,N_8403);
nand U9904 (N_9904,N_8951,N_8925);
nand U9905 (N_9905,N_8102,N_8848);
nand U9906 (N_9906,N_8270,N_8369);
xnor U9907 (N_9907,N_8266,N_8557);
nor U9908 (N_9908,N_8216,N_8707);
or U9909 (N_9909,N_8149,N_8607);
and U9910 (N_9910,N_8970,N_8722);
xor U9911 (N_9911,N_8998,N_8498);
or U9912 (N_9912,N_8771,N_8979);
nor U9913 (N_9913,N_8398,N_8902);
and U9914 (N_9914,N_8470,N_8625);
nor U9915 (N_9915,N_8219,N_8334);
xnor U9916 (N_9916,N_8353,N_8322);
or U9917 (N_9917,N_8817,N_8330);
or U9918 (N_9918,N_8073,N_8407);
and U9919 (N_9919,N_8086,N_8253);
or U9920 (N_9920,N_8858,N_8195);
nor U9921 (N_9921,N_8817,N_8073);
nor U9922 (N_9922,N_8024,N_8214);
nor U9923 (N_9923,N_8698,N_8741);
and U9924 (N_9924,N_8931,N_8806);
or U9925 (N_9925,N_8609,N_8799);
nand U9926 (N_9926,N_8145,N_8037);
xnor U9927 (N_9927,N_8184,N_8337);
or U9928 (N_9928,N_8155,N_8734);
or U9929 (N_9929,N_8445,N_8286);
or U9930 (N_9930,N_8983,N_8001);
xor U9931 (N_9931,N_8649,N_8407);
xnor U9932 (N_9932,N_8723,N_8520);
or U9933 (N_9933,N_8773,N_8170);
xor U9934 (N_9934,N_8949,N_8541);
nand U9935 (N_9935,N_8962,N_8724);
nor U9936 (N_9936,N_8437,N_8490);
and U9937 (N_9937,N_8955,N_8412);
nor U9938 (N_9938,N_8973,N_8013);
or U9939 (N_9939,N_8882,N_8700);
or U9940 (N_9940,N_8153,N_8227);
or U9941 (N_9941,N_8228,N_8168);
nor U9942 (N_9942,N_8344,N_8372);
or U9943 (N_9943,N_8291,N_8923);
nor U9944 (N_9944,N_8867,N_8602);
nor U9945 (N_9945,N_8641,N_8278);
xor U9946 (N_9946,N_8158,N_8395);
xor U9947 (N_9947,N_8938,N_8681);
or U9948 (N_9948,N_8682,N_8470);
xnor U9949 (N_9949,N_8246,N_8393);
nor U9950 (N_9950,N_8994,N_8553);
nor U9951 (N_9951,N_8320,N_8101);
nand U9952 (N_9952,N_8021,N_8665);
or U9953 (N_9953,N_8600,N_8223);
and U9954 (N_9954,N_8952,N_8006);
nand U9955 (N_9955,N_8185,N_8334);
or U9956 (N_9956,N_8261,N_8049);
or U9957 (N_9957,N_8973,N_8424);
nand U9958 (N_9958,N_8995,N_8344);
and U9959 (N_9959,N_8699,N_8627);
xor U9960 (N_9960,N_8763,N_8214);
nor U9961 (N_9961,N_8209,N_8775);
nor U9962 (N_9962,N_8443,N_8825);
and U9963 (N_9963,N_8834,N_8915);
nor U9964 (N_9964,N_8863,N_8866);
nor U9965 (N_9965,N_8598,N_8741);
xor U9966 (N_9966,N_8776,N_8793);
nor U9967 (N_9967,N_8697,N_8756);
nand U9968 (N_9968,N_8243,N_8766);
nand U9969 (N_9969,N_8961,N_8042);
nor U9970 (N_9970,N_8743,N_8325);
xor U9971 (N_9971,N_8910,N_8117);
nor U9972 (N_9972,N_8691,N_8018);
or U9973 (N_9973,N_8636,N_8963);
or U9974 (N_9974,N_8220,N_8868);
xor U9975 (N_9975,N_8934,N_8179);
or U9976 (N_9976,N_8356,N_8624);
or U9977 (N_9977,N_8337,N_8922);
xnor U9978 (N_9978,N_8826,N_8533);
or U9979 (N_9979,N_8114,N_8563);
nand U9980 (N_9980,N_8789,N_8627);
and U9981 (N_9981,N_8459,N_8537);
xnor U9982 (N_9982,N_8915,N_8156);
or U9983 (N_9983,N_8423,N_8399);
or U9984 (N_9984,N_8348,N_8445);
nand U9985 (N_9985,N_8140,N_8908);
xnor U9986 (N_9986,N_8816,N_8754);
or U9987 (N_9987,N_8434,N_8115);
nor U9988 (N_9988,N_8882,N_8333);
and U9989 (N_9989,N_8338,N_8100);
and U9990 (N_9990,N_8987,N_8766);
nand U9991 (N_9991,N_8234,N_8654);
or U9992 (N_9992,N_8300,N_8768);
and U9993 (N_9993,N_8176,N_8232);
and U9994 (N_9994,N_8605,N_8840);
and U9995 (N_9995,N_8101,N_8450);
xor U9996 (N_9996,N_8064,N_8626);
and U9997 (N_9997,N_8624,N_8357);
and U9998 (N_9998,N_8583,N_8455);
nor U9999 (N_9999,N_8435,N_8468);
nor U10000 (N_10000,N_9166,N_9213);
nand U10001 (N_10001,N_9487,N_9311);
xnor U10002 (N_10002,N_9196,N_9492);
nor U10003 (N_10003,N_9807,N_9943);
and U10004 (N_10004,N_9366,N_9647);
nand U10005 (N_10005,N_9678,N_9950);
or U10006 (N_10006,N_9340,N_9371);
or U10007 (N_10007,N_9184,N_9866);
nand U10008 (N_10008,N_9860,N_9864);
or U10009 (N_10009,N_9242,N_9164);
and U10010 (N_10010,N_9175,N_9552);
nor U10011 (N_10011,N_9285,N_9100);
nor U10012 (N_10012,N_9185,N_9009);
or U10013 (N_10013,N_9791,N_9962);
or U10014 (N_10014,N_9924,N_9339);
and U10015 (N_10015,N_9952,N_9514);
xor U10016 (N_10016,N_9137,N_9097);
xor U10017 (N_10017,N_9964,N_9325);
and U10018 (N_10018,N_9300,N_9410);
or U10019 (N_10019,N_9226,N_9427);
nor U10020 (N_10020,N_9954,N_9178);
nor U10021 (N_10021,N_9521,N_9103);
and U10022 (N_10022,N_9031,N_9294);
nand U10023 (N_10023,N_9737,N_9169);
xor U10024 (N_10024,N_9619,N_9150);
or U10025 (N_10025,N_9604,N_9569);
nor U10026 (N_10026,N_9885,N_9529);
nand U10027 (N_10027,N_9775,N_9878);
nand U10028 (N_10028,N_9318,N_9803);
and U10029 (N_10029,N_9008,N_9387);
nor U10030 (N_10030,N_9188,N_9043);
nand U10031 (N_10031,N_9898,N_9687);
or U10032 (N_10032,N_9617,N_9152);
nand U10033 (N_10033,N_9180,N_9580);
and U10034 (N_10034,N_9802,N_9468);
or U10035 (N_10035,N_9120,N_9625);
and U10036 (N_10036,N_9706,N_9434);
xnor U10037 (N_10037,N_9527,N_9862);
or U10038 (N_10038,N_9795,N_9846);
and U10039 (N_10039,N_9089,N_9034);
nand U10040 (N_10040,N_9591,N_9078);
or U10041 (N_10041,N_9021,N_9545);
and U10042 (N_10042,N_9124,N_9224);
nand U10043 (N_10043,N_9312,N_9859);
or U10044 (N_10044,N_9852,N_9870);
xnor U10045 (N_10045,N_9025,N_9942);
nor U10046 (N_10046,N_9970,N_9108);
and U10047 (N_10047,N_9961,N_9946);
or U10048 (N_10048,N_9461,N_9844);
or U10049 (N_10049,N_9140,N_9252);
xnor U10050 (N_10050,N_9098,N_9289);
xnor U10051 (N_10051,N_9787,N_9744);
or U10052 (N_10052,N_9588,N_9331);
and U10053 (N_10053,N_9270,N_9448);
or U10054 (N_10054,N_9201,N_9128);
or U10055 (N_10055,N_9141,N_9705);
xor U10056 (N_10056,N_9075,N_9477);
and U10057 (N_10057,N_9364,N_9272);
nor U10058 (N_10058,N_9725,N_9794);
nor U10059 (N_10059,N_9922,N_9876);
and U10060 (N_10060,N_9000,N_9475);
xnor U10061 (N_10061,N_9996,N_9189);
and U10062 (N_10062,N_9784,N_9642);
nand U10063 (N_10063,N_9457,N_9296);
or U10064 (N_10064,N_9319,N_9643);
xnor U10065 (N_10065,N_9435,N_9253);
or U10066 (N_10066,N_9686,N_9131);
and U10067 (N_10067,N_9941,N_9388);
and U10068 (N_10068,N_9338,N_9723);
nand U10069 (N_10069,N_9576,N_9167);
and U10070 (N_10070,N_9717,N_9293);
xnor U10071 (N_10071,N_9187,N_9987);
nor U10072 (N_10072,N_9506,N_9732);
nor U10073 (N_10073,N_9033,N_9478);
or U10074 (N_10074,N_9072,N_9173);
nand U10075 (N_10075,N_9548,N_9231);
or U10076 (N_10076,N_9838,N_9491);
nand U10077 (N_10077,N_9443,N_9405);
or U10078 (N_10078,N_9244,N_9404);
xnor U10079 (N_10079,N_9394,N_9416);
xor U10080 (N_10080,N_9903,N_9986);
or U10081 (N_10081,N_9112,N_9337);
or U10082 (N_10082,N_9469,N_9958);
xor U10083 (N_10083,N_9248,N_9606);
nor U10084 (N_10084,N_9110,N_9016);
and U10085 (N_10085,N_9585,N_9225);
and U10086 (N_10086,N_9991,N_9909);
nor U10087 (N_10087,N_9317,N_9972);
and U10088 (N_10088,N_9194,N_9519);
xor U10089 (N_10089,N_9249,N_9589);
and U10090 (N_10090,N_9474,N_9010);
xnor U10091 (N_10091,N_9420,N_9740);
nor U10092 (N_10092,N_9851,N_9682);
or U10093 (N_10093,N_9526,N_9276);
xor U10094 (N_10094,N_9779,N_9967);
and U10095 (N_10095,N_9710,N_9875);
and U10096 (N_10096,N_9442,N_9910);
xnor U10097 (N_10097,N_9336,N_9676);
or U10098 (N_10098,N_9505,N_9171);
nand U10099 (N_10099,N_9210,N_9161);
nand U10100 (N_10100,N_9049,N_9216);
nor U10101 (N_10101,N_9947,N_9900);
and U10102 (N_10102,N_9990,N_9738);
and U10103 (N_10103,N_9623,N_9406);
xnor U10104 (N_10104,N_9843,N_9702);
or U10105 (N_10105,N_9824,N_9132);
nor U10106 (N_10106,N_9525,N_9592);
nor U10107 (N_10107,N_9808,N_9648);
or U10108 (N_10108,N_9309,N_9812);
xor U10109 (N_10109,N_9626,N_9805);
nor U10110 (N_10110,N_9672,N_9933);
nor U10111 (N_10111,N_9065,N_9939);
and U10112 (N_10112,N_9241,N_9284);
and U10113 (N_10113,N_9644,N_9279);
xor U10114 (N_10114,N_9684,N_9848);
and U10115 (N_10115,N_9635,N_9931);
nor U10116 (N_10116,N_9800,N_9104);
nor U10117 (N_10117,N_9256,N_9530);
xor U10118 (N_10118,N_9409,N_9666);
nor U10119 (N_10119,N_9245,N_9520);
and U10120 (N_10120,N_9282,N_9344);
nand U10121 (N_10121,N_9286,N_9446);
nor U10122 (N_10122,N_9022,N_9992);
nand U10123 (N_10123,N_9953,N_9746);
nor U10124 (N_10124,N_9380,N_9694);
or U10125 (N_10125,N_9561,N_9099);
and U10126 (N_10126,N_9810,N_9801);
nand U10127 (N_10127,N_9481,N_9865);
xnor U10128 (N_10128,N_9391,N_9759);
and U10129 (N_10129,N_9259,N_9711);
nand U10130 (N_10130,N_9517,N_9584);
and U10131 (N_10131,N_9788,N_9271);
nand U10132 (N_10132,N_9424,N_9873);
nor U10133 (N_10133,N_9915,N_9663);
or U10134 (N_10134,N_9280,N_9608);
or U10135 (N_10135,N_9618,N_9251);
or U10136 (N_10136,N_9165,N_9264);
nor U10137 (N_10137,N_9287,N_9148);
or U10138 (N_10138,N_9841,N_9060);
xnor U10139 (N_10139,N_9056,N_9834);
xor U10140 (N_10140,N_9799,N_9328);
or U10141 (N_10141,N_9265,N_9713);
nand U10142 (N_10142,N_9645,N_9707);
and U10143 (N_10143,N_9361,N_9959);
and U10144 (N_10144,N_9334,N_9908);
xnor U10145 (N_10145,N_9412,N_9290);
or U10146 (N_10146,N_9747,N_9955);
xor U10147 (N_10147,N_9353,N_9471);
or U10148 (N_10148,N_9275,N_9735);
nand U10149 (N_10149,N_9599,N_9845);
nand U10150 (N_10150,N_9899,N_9555);
or U10151 (N_10151,N_9114,N_9886);
or U10152 (N_10152,N_9751,N_9501);
nor U10153 (N_10153,N_9088,N_9607);
xnor U10154 (N_10154,N_9837,N_9414);
and U10155 (N_10155,N_9912,N_9534);
and U10156 (N_10156,N_9179,N_9062);
nor U10157 (N_10157,N_9699,N_9454);
nand U10158 (N_10158,N_9786,N_9206);
or U10159 (N_10159,N_9299,N_9028);
nor U10160 (N_10160,N_9722,N_9221);
xnor U10161 (N_10161,N_9087,N_9884);
nand U10162 (N_10162,N_9887,N_9639);
and U10163 (N_10163,N_9273,N_9960);
nand U10164 (N_10164,N_9726,N_9596);
xnor U10165 (N_10165,N_9879,N_9489);
nor U10166 (N_10166,N_9789,N_9346);
xnor U10167 (N_10167,N_9565,N_9162);
xnor U10168 (N_10168,N_9703,N_9556);
and U10169 (N_10169,N_9204,N_9754);
xor U10170 (N_10170,N_9039,N_9382);
nor U10171 (N_10171,N_9709,N_9237);
nand U10172 (N_10172,N_9350,N_9826);
nor U10173 (N_10173,N_9050,N_9059);
or U10174 (N_10174,N_9721,N_9069);
xnor U10175 (N_10175,N_9651,N_9698);
nor U10176 (N_10176,N_9988,N_9764);
xor U10177 (N_10177,N_9055,N_9882);
nor U10178 (N_10178,N_9701,N_9568);
and U10179 (N_10179,N_9504,N_9258);
or U10180 (N_10180,N_9030,N_9748);
or U10181 (N_10181,N_9869,N_9914);
xor U10182 (N_10182,N_9136,N_9133);
xor U10183 (N_10183,N_9816,N_9266);
xnor U10184 (N_10184,N_9278,N_9020);
nor U10185 (N_10185,N_9190,N_9611);
nand U10186 (N_10186,N_9785,N_9982);
xor U10187 (N_10187,N_9586,N_9086);
and U10188 (N_10188,N_9881,N_9329);
nor U10189 (N_10189,N_9111,N_9813);
xor U10190 (N_10190,N_9641,N_9154);
nor U10191 (N_10191,N_9392,N_9809);
nand U10192 (N_10192,N_9295,N_9255);
nand U10193 (N_10193,N_9855,N_9398);
xor U10194 (N_10194,N_9923,N_9904);
nor U10195 (N_10195,N_9428,N_9322);
xor U10196 (N_10196,N_9850,N_9743);
and U10197 (N_10197,N_9811,N_9142);
nand U10198 (N_10198,N_9681,N_9562);
and U10199 (N_10199,N_9037,N_9590);
xnor U10200 (N_10200,N_9609,N_9359);
xnor U10201 (N_10201,N_9828,N_9630);
and U10202 (N_10202,N_9306,N_9368);
xnor U10203 (N_10203,N_9724,N_9664);
and U10204 (N_10204,N_9806,N_9499);
xnor U10205 (N_10205,N_9024,N_9979);
nor U10206 (N_10206,N_9745,N_9292);
xor U10207 (N_10207,N_9831,N_9195);
nand U10208 (N_10208,N_9503,N_9096);
or U10209 (N_10209,N_9728,N_9938);
xnor U10210 (N_10210,N_9426,N_9934);
and U10211 (N_10211,N_9598,N_9127);
nor U10212 (N_10212,N_9401,N_9830);
nand U10213 (N_10213,N_9155,N_9734);
or U10214 (N_10214,N_9763,N_9369);
and U10215 (N_10215,N_9399,N_9080);
nand U10216 (N_10216,N_9767,N_9157);
nand U10217 (N_10217,N_9593,N_9181);
nor U10218 (N_10218,N_9151,N_9484);
or U10219 (N_10219,N_9143,N_9948);
xnor U10220 (N_10220,N_9153,N_9386);
xnor U10221 (N_10221,N_9458,N_9652);
nand U10222 (N_10222,N_9323,N_9758);
nand U10223 (N_10223,N_9537,N_9485);
nor U10224 (N_10224,N_9307,N_9999);
nand U10225 (N_10225,N_9782,N_9765);
nor U10226 (N_10226,N_9436,N_9889);
nand U10227 (N_10227,N_9857,N_9572);
xnor U10228 (N_10228,N_9822,N_9560);
or U10229 (N_10229,N_9536,N_9183);
nand U10230 (N_10230,N_9773,N_9298);
and U10231 (N_10231,N_9832,N_9389);
nor U10232 (N_10232,N_9460,N_9983);
nand U10233 (N_10233,N_9488,N_9633);
nor U10234 (N_10234,N_9662,N_9126);
or U10235 (N_10235,N_9470,N_9144);
xnor U10236 (N_10236,N_9796,N_9559);
nor U10237 (N_10237,N_9227,N_9036);
or U10238 (N_10238,N_9441,N_9139);
nand U10239 (N_10239,N_9352,N_9814);
or U10240 (N_10240,N_9170,N_9310);
nand U10241 (N_10241,N_9697,N_9197);
nor U10242 (N_10242,N_9483,N_9455);
nor U10243 (N_10243,N_9594,N_9291);
or U10244 (N_10244,N_9776,N_9603);
and U10245 (N_10245,N_9018,N_9753);
and U10246 (N_10246,N_9232,N_9281);
or U10247 (N_10247,N_9379,N_9957);
nand U10248 (N_10248,N_9397,N_9940);
or U10249 (N_10249,N_9730,N_9736);
or U10250 (N_10250,N_9675,N_9655);
or U10251 (N_10251,N_9771,N_9015);
and U10252 (N_10252,N_9911,N_9906);
xnor U10253 (N_10253,N_9212,N_9752);
and U10254 (N_10254,N_9007,N_9067);
nand U10255 (N_10255,N_9877,N_9544);
or U10256 (N_10256,N_9182,N_9493);
and U10257 (N_10257,N_9393,N_9739);
nor U10258 (N_10258,N_9411,N_9601);
or U10259 (N_10259,N_9650,N_9781);
xor U10260 (N_10260,N_9577,N_9835);
nand U10261 (N_10261,N_9396,N_9616);
nor U10262 (N_10262,N_9381,N_9349);
nor U10263 (N_10263,N_9466,N_9011);
nor U10264 (N_10264,N_9949,N_9006);
nand U10265 (N_10265,N_9083,N_9668);
xor U10266 (N_10266,N_9172,N_9692);
xor U10267 (N_10267,N_9581,N_9315);
and U10268 (N_10268,N_9313,N_9741);
xnor U10269 (N_10269,N_9825,N_9936);
and U10270 (N_10270,N_9376,N_9228);
nand U10271 (N_10271,N_9689,N_9624);
nand U10272 (N_10272,N_9357,N_9102);
nor U10273 (N_10273,N_9238,N_9774);
or U10274 (N_10274,N_9839,N_9342);
nor U10275 (N_10275,N_9354,N_9314);
or U10276 (N_10276,N_9042,N_9288);
and U10277 (N_10277,N_9973,N_9622);
nor U10278 (N_10278,N_9450,N_9250);
xor U10279 (N_10279,N_9177,N_9163);
and U10280 (N_10280,N_9613,N_9004);
nor U10281 (N_10281,N_9134,N_9130);
nand U10282 (N_10282,N_9229,N_9054);
and U10283 (N_10283,N_9595,N_9467);
xnor U10284 (N_10284,N_9550,N_9490);
xnor U10285 (N_10285,N_9755,N_9920);
or U10286 (N_10286,N_9551,N_9439);
and U10287 (N_10287,N_9963,N_9246);
and U10288 (N_10288,N_9965,N_9610);
nand U10289 (N_10289,N_9531,N_9343);
and U10290 (N_10290,N_9516,N_9612);
and U10291 (N_10291,N_9919,N_9935);
xnor U10292 (N_10292,N_9208,N_9892);
xor U10293 (N_10293,N_9355,N_9425);
xnor U10294 (N_10294,N_9944,N_9451);
and U10295 (N_10295,N_9649,N_9332);
nor U10296 (N_10296,N_9160,N_9567);
or U10297 (N_10297,N_9057,N_9433);
nor U10298 (N_10298,N_9989,N_9541);
nor U10299 (N_10299,N_9894,N_9512);
xnor U10300 (N_10300,N_9115,N_9400);
and U10301 (N_10301,N_9688,N_9040);
or U10302 (N_10302,N_9146,N_9677);
nand U10303 (N_10303,N_9463,N_9994);
or U10304 (N_10304,N_9017,N_9327);
or U10305 (N_10305,N_9997,N_9815);
nor U10306 (N_10306,N_9093,N_9254);
nor U10307 (N_10307,N_9928,N_9303);
nand U10308 (N_10308,N_9360,N_9533);
nand U10309 (N_10309,N_9792,N_9001);
nor U10310 (N_10310,N_9316,N_9502);
or U10311 (N_10311,N_9444,N_9497);
and U10312 (N_10312,N_9092,N_9749);
or U10313 (N_10313,N_9817,N_9695);
and U10314 (N_10314,N_9277,N_9575);
nand U10315 (N_10315,N_9351,N_9714);
and U10316 (N_10316,N_9003,N_9498);
nor U10317 (N_10317,N_9578,N_9856);
nor U10318 (N_10318,N_9304,N_9207);
nand U10319 (N_10319,N_9156,N_9109);
or U10320 (N_10320,N_9186,N_9459);
nor U10321 (N_10321,N_9440,N_9880);
nor U10322 (N_10322,N_9956,N_9883);
nand U10323 (N_10323,N_9966,N_9637);
xnor U10324 (N_10324,N_9408,N_9661);
nor U10325 (N_10325,N_9984,N_9081);
xnor U10326 (N_10326,N_9430,N_9968);
and U10327 (N_10327,N_9657,N_9925);
nand U10328 (N_10328,N_9191,N_9896);
nor U10329 (N_10329,N_9048,N_9704);
and U10330 (N_10330,N_9222,N_9239);
or U10331 (N_10331,N_9901,N_9119);
nand U10332 (N_10332,N_9367,N_9417);
xnor U10333 (N_10333,N_9605,N_9780);
and U10334 (N_10334,N_9496,N_9429);
nand U10335 (N_10335,N_9070,N_9472);
or U10336 (N_10336,N_9220,N_9659);
nor U10337 (N_10337,N_9107,N_9384);
or U10338 (N_10338,N_9921,N_9116);
nor U10339 (N_10339,N_9579,N_9587);
nor U10340 (N_10340,N_9902,N_9044);
xor U10341 (N_10341,N_9403,N_9729);
nor U10342 (N_10342,N_9449,N_9302);
xor U10343 (N_10343,N_9917,N_9413);
and U10344 (N_10344,N_9821,N_9341);
xnor U10345 (N_10345,N_9653,N_9854);
nor U10346 (N_10346,N_9975,N_9211);
and U10347 (N_10347,N_9365,N_9507);
or U10348 (N_10348,N_9793,N_9632);
xor U10349 (N_10349,N_9634,N_9432);
and U10350 (N_10350,N_9372,N_9438);
and U10351 (N_10351,N_9456,N_9066);
and U10352 (N_10352,N_9113,N_9669);
or U10353 (N_10353,N_9797,N_9897);
xor U10354 (N_10354,N_9482,N_9247);
and U10355 (N_10355,N_9638,N_9683);
or U10356 (N_10356,N_9085,N_9829);
or U10357 (N_10357,N_9777,N_9158);
and U10358 (N_10358,N_9918,N_9890);
or U10359 (N_10359,N_9553,N_9535);
or U10360 (N_10360,N_9762,N_9064);
or U10361 (N_10361,N_9118,N_9716);
xor U10362 (N_10362,N_9766,N_9523);
or U10363 (N_10363,N_9464,N_9508);
xor U10364 (N_10364,N_9082,N_9262);
xor U10365 (N_10365,N_9192,N_9974);
and U10366 (N_10366,N_9218,N_9301);
nand U10367 (N_10367,N_9026,N_9554);
and U10368 (N_10368,N_9176,N_9422);
xnor U10369 (N_10369,N_9691,N_9308);
and U10370 (N_10370,N_9861,N_9045);
nand U10371 (N_10371,N_9891,N_9077);
and U10372 (N_10372,N_9976,N_9515);
and U10373 (N_10373,N_9636,N_9423);
nor U10374 (N_10374,N_9462,N_9971);
nand U10375 (N_10375,N_9658,N_9756);
xor U10376 (N_10376,N_9094,N_9421);
and U10377 (N_10377,N_9511,N_9680);
and U10378 (N_10378,N_9546,N_9079);
nand U10379 (N_10379,N_9842,N_9640);
nand U10380 (N_10380,N_9932,N_9673);
nor U10381 (N_10381,N_9370,N_9564);
nor U10382 (N_10382,N_9868,N_9926);
nor U10383 (N_10383,N_9269,N_9833);
and U10384 (N_10384,N_9261,N_9768);
or U10385 (N_10385,N_9538,N_9363);
or U10386 (N_10386,N_9893,N_9674);
nand U10387 (N_10387,N_9977,N_9895);
nand U10388 (N_10388,N_9665,N_9129);
nor U10389 (N_10389,N_9863,N_9377);
or U10390 (N_10390,N_9047,N_9135);
nand U10391 (N_10391,N_9347,N_9073);
xnor U10392 (N_10392,N_9145,N_9566);
xnor U10393 (N_10393,N_9540,N_9872);
or U10394 (N_10394,N_9203,N_9847);
or U10395 (N_10395,N_9305,N_9620);
nor U10396 (N_10396,N_9234,N_9121);
and U10397 (N_10397,N_9627,N_9597);
or U10398 (N_10398,N_9867,N_9798);
or U10399 (N_10399,N_9685,N_9257);
nor U10400 (N_10400,N_9951,N_9916);
and U10401 (N_10401,N_9542,N_9263);
xor U10402 (N_10402,N_9035,N_9670);
nand U10403 (N_10403,N_9200,N_9750);
and U10404 (N_10404,N_9378,N_9236);
or U10405 (N_10405,N_9819,N_9106);
nor U10406 (N_10406,N_9091,N_9927);
xor U10407 (N_10407,N_9549,N_9820);
or U10408 (N_10408,N_9836,N_9849);
xor U10409 (N_10409,N_9528,N_9667);
and U10410 (N_10410,N_9495,N_9871);
or U10411 (N_10411,N_9582,N_9978);
or U10412 (N_10412,N_9117,N_9772);
or U10413 (N_10413,N_9760,N_9557);
xnor U10414 (N_10414,N_9076,N_9818);
and U10415 (N_10415,N_9159,N_9029);
nor U10416 (N_10416,N_9321,N_9374);
and U10417 (N_10417,N_9358,N_9452);
or U10418 (N_10418,N_9240,N_9679);
xor U10419 (N_10419,N_9696,N_9731);
xor U10420 (N_10420,N_9660,N_9543);
xor U10421 (N_10421,N_9905,N_9202);
xnor U10422 (N_10422,N_9524,N_9907);
or U10423 (N_10423,N_9715,N_9823);
nor U10424 (N_10424,N_9168,N_9061);
nor U10425 (N_10425,N_9518,N_9002);
nand U10426 (N_10426,N_9084,N_9419);
nor U10427 (N_10427,N_9437,N_9373);
or U10428 (N_10428,N_9693,N_9510);
nor U10429 (N_10429,N_9297,N_9719);
and U10430 (N_10430,N_9473,N_9356);
and U10431 (N_10431,N_9654,N_9013);
and U10432 (N_10432,N_9853,N_9205);
and U10433 (N_10433,N_9324,N_9742);
or U10434 (N_10434,N_9267,N_9012);
and U10435 (N_10435,N_9720,N_9283);
nor U10436 (N_10436,N_9320,N_9558);
or U10437 (N_10437,N_9125,N_9052);
nor U10438 (N_10438,N_9046,N_9500);
xor U10439 (N_10439,N_9671,N_9233);
or U10440 (N_10440,N_9074,N_9058);
xnor U10441 (N_10441,N_9038,N_9757);
and U10442 (N_10442,N_9929,N_9209);
and U10443 (N_10443,N_9969,N_9217);
nand U10444 (N_10444,N_9727,N_9395);
and U10445 (N_10445,N_9215,N_9274);
nand U10446 (N_10446,N_9614,N_9930);
and U10447 (N_10447,N_9600,N_9053);
and U10448 (N_10448,N_9937,N_9628);
and U10449 (N_10449,N_9700,N_9090);
nor U10450 (N_10450,N_9770,N_9032);
nand U10451 (N_10451,N_9712,N_9509);
nor U10452 (N_10452,N_9101,N_9214);
nand U10453 (N_10453,N_9385,N_9453);
or U10454 (N_10454,N_9330,N_9486);
xnor U10455 (N_10455,N_9761,N_9888);
nand U10456 (N_10456,N_9174,N_9375);
and U10457 (N_10457,N_9629,N_9573);
and U10458 (N_10458,N_9447,N_9494);
and U10459 (N_10459,N_9138,N_9945);
or U10460 (N_10460,N_9068,N_9260);
nor U10461 (N_10461,N_9230,N_9783);
xnor U10462 (N_10462,N_9563,N_9631);
or U10463 (N_10463,N_9345,N_9333);
nand U10464 (N_10464,N_9778,N_9219);
xor U10465 (N_10465,N_9445,N_9023);
nor U10466 (N_10466,N_9690,N_9105);
and U10467 (N_10467,N_9513,N_9005);
xor U10468 (N_10468,N_9383,N_9476);
or U10469 (N_10469,N_9123,N_9335);
nand U10470 (N_10470,N_9539,N_9615);
or U10471 (N_10471,N_9027,N_9063);
nor U10472 (N_10472,N_9790,N_9243);
and U10473 (N_10473,N_9014,N_9402);
nor U10474 (N_10474,N_9602,N_9708);
nand U10475 (N_10475,N_9827,N_9981);
and U10476 (N_10476,N_9198,N_9656);
nand U10477 (N_10477,N_9326,N_9522);
nor U10478 (N_10478,N_9149,N_9019);
nor U10479 (N_10479,N_9547,N_9985);
or U10480 (N_10480,N_9840,N_9071);
or U10481 (N_10481,N_9769,N_9874);
nor U10482 (N_10482,N_9532,N_9362);
xnor U10483 (N_10483,N_9415,N_9998);
or U10484 (N_10484,N_9199,N_9995);
or U10485 (N_10485,N_9571,N_9479);
and U10486 (N_10486,N_9348,N_9646);
xor U10487 (N_10487,N_9122,N_9390);
or U10488 (N_10488,N_9993,N_9407);
or U10489 (N_10489,N_9621,N_9858);
nor U10490 (N_10490,N_9583,N_9041);
nor U10491 (N_10491,N_9235,N_9193);
nor U10492 (N_10492,N_9718,N_9095);
or U10493 (N_10493,N_9804,N_9980);
and U10494 (N_10494,N_9268,N_9913);
xnor U10495 (N_10495,N_9570,N_9051);
xor U10496 (N_10496,N_9733,N_9465);
and U10497 (N_10497,N_9574,N_9147);
and U10498 (N_10498,N_9418,N_9431);
xor U10499 (N_10499,N_9480,N_9223);
xor U10500 (N_10500,N_9203,N_9338);
nand U10501 (N_10501,N_9299,N_9195);
nand U10502 (N_10502,N_9687,N_9575);
and U10503 (N_10503,N_9334,N_9919);
nor U10504 (N_10504,N_9683,N_9592);
nor U10505 (N_10505,N_9687,N_9681);
nand U10506 (N_10506,N_9501,N_9594);
nand U10507 (N_10507,N_9186,N_9492);
nand U10508 (N_10508,N_9784,N_9632);
nand U10509 (N_10509,N_9768,N_9891);
and U10510 (N_10510,N_9003,N_9788);
nand U10511 (N_10511,N_9163,N_9901);
xnor U10512 (N_10512,N_9573,N_9718);
nand U10513 (N_10513,N_9451,N_9194);
and U10514 (N_10514,N_9207,N_9776);
xnor U10515 (N_10515,N_9127,N_9109);
and U10516 (N_10516,N_9869,N_9711);
xnor U10517 (N_10517,N_9442,N_9939);
or U10518 (N_10518,N_9216,N_9797);
nor U10519 (N_10519,N_9442,N_9864);
nand U10520 (N_10520,N_9534,N_9756);
nand U10521 (N_10521,N_9038,N_9765);
nor U10522 (N_10522,N_9072,N_9810);
xnor U10523 (N_10523,N_9294,N_9539);
xnor U10524 (N_10524,N_9718,N_9141);
nor U10525 (N_10525,N_9958,N_9328);
nand U10526 (N_10526,N_9781,N_9134);
nor U10527 (N_10527,N_9773,N_9422);
and U10528 (N_10528,N_9250,N_9875);
nand U10529 (N_10529,N_9868,N_9513);
nor U10530 (N_10530,N_9715,N_9180);
nand U10531 (N_10531,N_9199,N_9634);
nor U10532 (N_10532,N_9104,N_9486);
and U10533 (N_10533,N_9164,N_9612);
and U10534 (N_10534,N_9246,N_9974);
nor U10535 (N_10535,N_9055,N_9818);
or U10536 (N_10536,N_9056,N_9609);
nor U10537 (N_10537,N_9432,N_9024);
or U10538 (N_10538,N_9126,N_9795);
nand U10539 (N_10539,N_9534,N_9031);
or U10540 (N_10540,N_9680,N_9780);
nor U10541 (N_10541,N_9567,N_9333);
xnor U10542 (N_10542,N_9690,N_9993);
and U10543 (N_10543,N_9975,N_9757);
nand U10544 (N_10544,N_9231,N_9405);
or U10545 (N_10545,N_9513,N_9623);
or U10546 (N_10546,N_9302,N_9028);
nand U10547 (N_10547,N_9171,N_9117);
nand U10548 (N_10548,N_9016,N_9342);
and U10549 (N_10549,N_9653,N_9785);
and U10550 (N_10550,N_9457,N_9461);
or U10551 (N_10551,N_9145,N_9465);
and U10552 (N_10552,N_9864,N_9434);
or U10553 (N_10553,N_9318,N_9386);
nand U10554 (N_10554,N_9995,N_9150);
and U10555 (N_10555,N_9292,N_9070);
xor U10556 (N_10556,N_9241,N_9439);
nor U10557 (N_10557,N_9794,N_9172);
nand U10558 (N_10558,N_9302,N_9430);
nor U10559 (N_10559,N_9592,N_9123);
or U10560 (N_10560,N_9855,N_9052);
and U10561 (N_10561,N_9108,N_9035);
nand U10562 (N_10562,N_9991,N_9289);
nor U10563 (N_10563,N_9571,N_9623);
and U10564 (N_10564,N_9686,N_9329);
or U10565 (N_10565,N_9364,N_9922);
or U10566 (N_10566,N_9710,N_9406);
nand U10567 (N_10567,N_9370,N_9792);
and U10568 (N_10568,N_9359,N_9601);
nand U10569 (N_10569,N_9852,N_9327);
and U10570 (N_10570,N_9029,N_9477);
nor U10571 (N_10571,N_9072,N_9771);
nand U10572 (N_10572,N_9302,N_9361);
and U10573 (N_10573,N_9227,N_9395);
nand U10574 (N_10574,N_9998,N_9958);
or U10575 (N_10575,N_9058,N_9208);
nor U10576 (N_10576,N_9479,N_9239);
nand U10577 (N_10577,N_9888,N_9146);
xnor U10578 (N_10578,N_9718,N_9315);
and U10579 (N_10579,N_9625,N_9908);
nand U10580 (N_10580,N_9486,N_9075);
and U10581 (N_10581,N_9107,N_9469);
and U10582 (N_10582,N_9486,N_9810);
or U10583 (N_10583,N_9800,N_9991);
xor U10584 (N_10584,N_9073,N_9704);
nand U10585 (N_10585,N_9571,N_9732);
xor U10586 (N_10586,N_9659,N_9910);
or U10587 (N_10587,N_9952,N_9988);
or U10588 (N_10588,N_9629,N_9831);
nor U10589 (N_10589,N_9403,N_9164);
nor U10590 (N_10590,N_9752,N_9636);
xnor U10591 (N_10591,N_9181,N_9415);
or U10592 (N_10592,N_9942,N_9090);
or U10593 (N_10593,N_9523,N_9225);
or U10594 (N_10594,N_9763,N_9824);
and U10595 (N_10595,N_9903,N_9162);
nand U10596 (N_10596,N_9768,N_9098);
nor U10597 (N_10597,N_9936,N_9207);
nor U10598 (N_10598,N_9166,N_9484);
xnor U10599 (N_10599,N_9976,N_9251);
nor U10600 (N_10600,N_9853,N_9788);
nand U10601 (N_10601,N_9781,N_9989);
xor U10602 (N_10602,N_9415,N_9674);
nand U10603 (N_10603,N_9253,N_9823);
and U10604 (N_10604,N_9527,N_9421);
and U10605 (N_10605,N_9488,N_9849);
or U10606 (N_10606,N_9156,N_9443);
nand U10607 (N_10607,N_9287,N_9309);
or U10608 (N_10608,N_9038,N_9546);
nand U10609 (N_10609,N_9629,N_9825);
xnor U10610 (N_10610,N_9703,N_9064);
or U10611 (N_10611,N_9485,N_9612);
xnor U10612 (N_10612,N_9525,N_9097);
xor U10613 (N_10613,N_9918,N_9206);
or U10614 (N_10614,N_9228,N_9017);
nor U10615 (N_10615,N_9937,N_9283);
nand U10616 (N_10616,N_9598,N_9623);
or U10617 (N_10617,N_9532,N_9977);
or U10618 (N_10618,N_9749,N_9073);
nor U10619 (N_10619,N_9966,N_9901);
and U10620 (N_10620,N_9307,N_9791);
nor U10621 (N_10621,N_9370,N_9742);
nand U10622 (N_10622,N_9427,N_9449);
nand U10623 (N_10623,N_9650,N_9194);
nand U10624 (N_10624,N_9313,N_9662);
and U10625 (N_10625,N_9195,N_9502);
and U10626 (N_10626,N_9335,N_9275);
and U10627 (N_10627,N_9580,N_9592);
xnor U10628 (N_10628,N_9984,N_9678);
xor U10629 (N_10629,N_9541,N_9720);
nor U10630 (N_10630,N_9135,N_9639);
or U10631 (N_10631,N_9511,N_9939);
nand U10632 (N_10632,N_9231,N_9699);
and U10633 (N_10633,N_9025,N_9051);
nand U10634 (N_10634,N_9132,N_9144);
nor U10635 (N_10635,N_9946,N_9695);
or U10636 (N_10636,N_9863,N_9457);
nand U10637 (N_10637,N_9184,N_9966);
and U10638 (N_10638,N_9204,N_9912);
and U10639 (N_10639,N_9713,N_9046);
xor U10640 (N_10640,N_9712,N_9524);
and U10641 (N_10641,N_9808,N_9542);
or U10642 (N_10642,N_9141,N_9192);
nor U10643 (N_10643,N_9671,N_9258);
nand U10644 (N_10644,N_9003,N_9953);
xor U10645 (N_10645,N_9244,N_9089);
nor U10646 (N_10646,N_9020,N_9356);
and U10647 (N_10647,N_9403,N_9312);
nor U10648 (N_10648,N_9310,N_9348);
nand U10649 (N_10649,N_9267,N_9907);
nand U10650 (N_10650,N_9843,N_9999);
xnor U10651 (N_10651,N_9034,N_9347);
nand U10652 (N_10652,N_9728,N_9335);
nand U10653 (N_10653,N_9619,N_9882);
nor U10654 (N_10654,N_9632,N_9177);
and U10655 (N_10655,N_9716,N_9859);
or U10656 (N_10656,N_9335,N_9783);
xnor U10657 (N_10657,N_9416,N_9752);
xor U10658 (N_10658,N_9157,N_9921);
xnor U10659 (N_10659,N_9548,N_9679);
and U10660 (N_10660,N_9506,N_9976);
nand U10661 (N_10661,N_9222,N_9018);
or U10662 (N_10662,N_9468,N_9041);
or U10663 (N_10663,N_9985,N_9341);
and U10664 (N_10664,N_9082,N_9629);
nor U10665 (N_10665,N_9007,N_9677);
nor U10666 (N_10666,N_9871,N_9147);
xnor U10667 (N_10667,N_9344,N_9121);
or U10668 (N_10668,N_9290,N_9547);
xor U10669 (N_10669,N_9455,N_9531);
nor U10670 (N_10670,N_9282,N_9247);
nor U10671 (N_10671,N_9874,N_9961);
nand U10672 (N_10672,N_9982,N_9330);
nand U10673 (N_10673,N_9750,N_9951);
and U10674 (N_10674,N_9851,N_9233);
xnor U10675 (N_10675,N_9182,N_9798);
xor U10676 (N_10676,N_9833,N_9087);
nor U10677 (N_10677,N_9198,N_9534);
nor U10678 (N_10678,N_9367,N_9631);
nand U10679 (N_10679,N_9656,N_9977);
or U10680 (N_10680,N_9267,N_9272);
and U10681 (N_10681,N_9269,N_9174);
and U10682 (N_10682,N_9395,N_9954);
nor U10683 (N_10683,N_9863,N_9762);
nor U10684 (N_10684,N_9042,N_9241);
and U10685 (N_10685,N_9734,N_9708);
and U10686 (N_10686,N_9596,N_9841);
and U10687 (N_10687,N_9784,N_9019);
nand U10688 (N_10688,N_9761,N_9110);
or U10689 (N_10689,N_9340,N_9587);
nand U10690 (N_10690,N_9235,N_9448);
nor U10691 (N_10691,N_9880,N_9140);
nor U10692 (N_10692,N_9111,N_9293);
nand U10693 (N_10693,N_9350,N_9590);
xnor U10694 (N_10694,N_9289,N_9722);
nor U10695 (N_10695,N_9084,N_9551);
nor U10696 (N_10696,N_9621,N_9934);
nand U10697 (N_10697,N_9483,N_9236);
nor U10698 (N_10698,N_9408,N_9731);
nand U10699 (N_10699,N_9174,N_9636);
nor U10700 (N_10700,N_9535,N_9628);
and U10701 (N_10701,N_9116,N_9834);
nor U10702 (N_10702,N_9657,N_9587);
and U10703 (N_10703,N_9156,N_9196);
nor U10704 (N_10704,N_9310,N_9836);
or U10705 (N_10705,N_9854,N_9810);
and U10706 (N_10706,N_9369,N_9561);
nor U10707 (N_10707,N_9292,N_9260);
xor U10708 (N_10708,N_9217,N_9922);
and U10709 (N_10709,N_9479,N_9763);
xnor U10710 (N_10710,N_9479,N_9797);
or U10711 (N_10711,N_9715,N_9758);
and U10712 (N_10712,N_9952,N_9162);
or U10713 (N_10713,N_9567,N_9478);
nand U10714 (N_10714,N_9285,N_9944);
and U10715 (N_10715,N_9032,N_9306);
nor U10716 (N_10716,N_9332,N_9015);
and U10717 (N_10717,N_9090,N_9748);
or U10718 (N_10718,N_9121,N_9049);
xor U10719 (N_10719,N_9439,N_9588);
or U10720 (N_10720,N_9002,N_9279);
xnor U10721 (N_10721,N_9314,N_9548);
nor U10722 (N_10722,N_9804,N_9758);
or U10723 (N_10723,N_9105,N_9234);
xnor U10724 (N_10724,N_9194,N_9348);
and U10725 (N_10725,N_9671,N_9739);
xnor U10726 (N_10726,N_9910,N_9724);
xnor U10727 (N_10727,N_9159,N_9294);
or U10728 (N_10728,N_9296,N_9661);
nor U10729 (N_10729,N_9748,N_9068);
or U10730 (N_10730,N_9782,N_9270);
xor U10731 (N_10731,N_9136,N_9705);
nand U10732 (N_10732,N_9268,N_9609);
nand U10733 (N_10733,N_9048,N_9281);
or U10734 (N_10734,N_9443,N_9343);
nor U10735 (N_10735,N_9647,N_9975);
nand U10736 (N_10736,N_9167,N_9507);
and U10737 (N_10737,N_9652,N_9741);
and U10738 (N_10738,N_9879,N_9362);
nor U10739 (N_10739,N_9614,N_9612);
xnor U10740 (N_10740,N_9198,N_9813);
nor U10741 (N_10741,N_9177,N_9677);
or U10742 (N_10742,N_9705,N_9375);
or U10743 (N_10743,N_9179,N_9106);
and U10744 (N_10744,N_9675,N_9056);
and U10745 (N_10745,N_9894,N_9435);
nand U10746 (N_10746,N_9121,N_9853);
xnor U10747 (N_10747,N_9238,N_9865);
and U10748 (N_10748,N_9879,N_9574);
nand U10749 (N_10749,N_9533,N_9267);
or U10750 (N_10750,N_9915,N_9521);
xor U10751 (N_10751,N_9936,N_9897);
or U10752 (N_10752,N_9670,N_9566);
nor U10753 (N_10753,N_9013,N_9833);
and U10754 (N_10754,N_9572,N_9496);
xnor U10755 (N_10755,N_9623,N_9264);
and U10756 (N_10756,N_9091,N_9932);
xnor U10757 (N_10757,N_9010,N_9514);
and U10758 (N_10758,N_9645,N_9015);
nor U10759 (N_10759,N_9992,N_9505);
xor U10760 (N_10760,N_9426,N_9468);
or U10761 (N_10761,N_9058,N_9467);
and U10762 (N_10762,N_9445,N_9096);
nor U10763 (N_10763,N_9051,N_9745);
nand U10764 (N_10764,N_9592,N_9991);
nor U10765 (N_10765,N_9542,N_9251);
nor U10766 (N_10766,N_9487,N_9698);
xor U10767 (N_10767,N_9994,N_9224);
xnor U10768 (N_10768,N_9030,N_9438);
xnor U10769 (N_10769,N_9360,N_9359);
and U10770 (N_10770,N_9832,N_9227);
or U10771 (N_10771,N_9448,N_9289);
nor U10772 (N_10772,N_9538,N_9792);
or U10773 (N_10773,N_9646,N_9814);
nor U10774 (N_10774,N_9523,N_9542);
nor U10775 (N_10775,N_9036,N_9093);
and U10776 (N_10776,N_9147,N_9651);
and U10777 (N_10777,N_9027,N_9430);
nor U10778 (N_10778,N_9451,N_9961);
nand U10779 (N_10779,N_9158,N_9270);
nand U10780 (N_10780,N_9920,N_9558);
and U10781 (N_10781,N_9139,N_9395);
nand U10782 (N_10782,N_9644,N_9789);
nand U10783 (N_10783,N_9642,N_9561);
nand U10784 (N_10784,N_9934,N_9421);
or U10785 (N_10785,N_9892,N_9493);
xor U10786 (N_10786,N_9882,N_9308);
and U10787 (N_10787,N_9980,N_9728);
nand U10788 (N_10788,N_9658,N_9437);
or U10789 (N_10789,N_9864,N_9748);
nand U10790 (N_10790,N_9155,N_9047);
xor U10791 (N_10791,N_9403,N_9001);
nor U10792 (N_10792,N_9514,N_9893);
or U10793 (N_10793,N_9607,N_9105);
xnor U10794 (N_10794,N_9382,N_9203);
or U10795 (N_10795,N_9444,N_9963);
nor U10796 (N_10796,N_9414,N_9688);
nor U10797 (N_10797,N_9655,N_9648);
nor U10798 (N_10798,N_9659,N_9746);
xor U10799 (N_10799,N_9061,N_9147);
and U10800 (N_10800,N_9932,N_9646);
nand U10801 (N_10801,N_9395,N_9052);
nor U10802 (N_10802,N_9459,N_9875);
nor U10803 (N_10803,N_9421,N_9727);
nand U10804 (N_10804,N_9511,N_9801);
xor U10805 (N_10805,N_9383,N_9247);
or U10806 (N_10806,N_9805,N_9236);
or U10807 (N_10807,N_9150,N_9115);
nor U10808 (N_10808,N_9372,N_9180);
nand U10809 (N_10809,N_9008,N_9927);
and U10810 (N_10810,N_9463,N_9383);
nand U10811 (N_10811,N_9950,N_9773);
or U10812 (N_10812,N_9696,N_9022);
nor U10813 (N_10813,N_9589,N_9530);
nand U10814 (N_10814,N_9495,N_9202);
and U10815 (N_10815,N_9854,N_9352);
nand U10816 (N_10816,N_9670,N_9855);
or U10817 (N_10817,N_9202,N_9136);
xor U10818 (N_10818,N_9117,N_9004);
and U10819 (N_10819,N_9190,N_9136);
and U10820 (N_10820,N_9356,N_9623);
or U10821 (N_10821,N_9051,N_9378);
xnor U10822 (N_10822,N_9531,N_9194);
and U10823 (N_10823,N_9536,N_9839);
nor U10824 (N_10824,N_9810,N_9638);
and U10825 (N_10825,N_9932,N_9256);
nand U10826 (N_10826,N_9058,N_9097);
xor U10827 (N_10827,N_9976,N_9270);
nor U10828 (N_10828,N_9519,N_9458);
or U10829 (N_10829,N_9826,N_9578);
nor U10830 (N_10830,N_9014,N_9378);
or U10831 (N_10831,N_9452,N_9434);
xor U10832 (N_10832,N_9080,N_9891);
nand U10833 (N_10833,N_9754,N_9821);
and U10834 (N_10834,N_9672,N_9735);
nor U10835 (N_10835,N_9357,N_9121);
or U10836 (N_10836,N_9279,N_9140);
nor U10837 (N_10837,N_9035,N_9539);
and U10838 (N_10838,N_9326,N_9982);
nand U10839 (N_10839,N_9590,N_9954);
or U10840 (N_10840,N_9915,N_9465);
and U10841 (N_10841,N_9097,N_9186);
nand U10842 (N_10842,N_9982,N_9867);
nand U10843 (N_10843,N_9826,N_9796);
nor U10844 (N_10844,N_9746,N_9928);
and U10845 (N_10845,N_9474,N_9858);
xnor U10846 (N_10846,N_9738,N_9244);
xor U10847 (N_10847,N_9030,N_9439);
or U10848 (N_10848,N_9285,N_9148);
or U10849 (N_10849,N_9440,N_9281);
nand U10850 (N_10850,N_9532,N_9086);
xor U10851 (N_10851,N_9206,N_9802);
and U10852 (N_10852,N_9612,N_9972);
nand U10853 (N_10853,N_9280,N_9776);
nor U10854 (N_10854,N_9730,N_9135);
and U10855 (N_10855,N_9386,N_9076);
nand U10856 (N_10856,N_9293,N_9445);
nor U10857 (N_10857,N_9166,N_9929);
nor U10858 (N_10858,N_9828,N_9635);
or U10859 (N_10859,N_9657,N_9121);
or U10860 (N_10860,N_9761,N_9204);
nor U10861 (N_10861,N_9262,N_9321);
or U10862 (N_10862,N_9319,N_9668);
xor U10863 (N_10863,N_9475,N_9293);
nand U10864 (N_10864,N_9502,N_9107);
nand U10865 (N_10865,N_9627,N_9955);
xnor U10866 (N_10866,N_9951,N_9402);
xnor U10867 (N_10867,N_9736,N_9192);
xnor U10868 (N_10868,N_9261,N_9981);
xor U10869 (N_10869,N_9728,N_9841);
xor U10870 (N_10870,N_9475,N_9226);
and U10871 (N_10871,N_9527,N_9398);
xnor U10872 (N_10872,N_9474,N_9251);
or U10873 (N_10873,N_9849,N_9801);
xnor U10874 (N_10874,N_9790,N_9681);
and U10875 (N_10875,N_9168,N_9096);
or U10876 (N_10876,N_9607,N_9358);
xor U10877 (N_10877,N_9248,N_9265);
nand U10878 (N_10878,N_9515,N_9696);
or U10879 (N_10879,N_9317,N_9214);
or U10880 (N_10880,N_9380,N_9662);
or U10881 (N_10881,N_9102,N_9002);
nor U10882 (N_10882,N_9862,N_9507);
nor U10883 (N_10883,N_9039,N_9064);
nor U10884 (N_10884,N_9913,N_9795);
or U10885 (N_10885,N_9627,N_9152);
and U10886 (N_10886,N_9826,N_9850);
and U10887 (N_10887,N_9761,N_9740);
nand U10888 (N_10888,N_9453,N_9529);
nor U10889 (N_10889,N_9128,N_9743);
nor U10890 (N_10890,N_9736,N_9818);
xor U10891 (N_10891,N_9266,N_9323);
nor U10892 (N_10892,N_9869,N_9602);
nand U10893 (N_10893,N_9612,N_9571);
or U10894 (N_10894,N_9290,N_9162);
and U10895 (N_10895,N_9883,N_9167);
and U10896 (N_10896,N_9387,N_9716);
or U10897 (N_10897,N_9684,N_9228);
nand U10898 (N_10898,N_9956,N_9003);
nand U10899 (N_10899,N_9763,N_9508);
xor U10900 (N_10900,N_9609,N_9957);
and U10901 (N_10901,N_9625,N_9776);
nor U10902 (N_10902,N_9100,N_9364);
or U10903 (N_10903,N_9712,N_9680);
and U10904 (N_10904,N_9806,N_9532);
nor U10905 (N_10905,N_9849,N_9252);
nand U10906 (N_10906,N_9380,N_9516);
and U10907 (N_10907,N_9212,N_9038);
and U10908 (N_10908,N_9941,N_9027);
nor U10909 (N_10909,N_9544,N_9405);
and U10910 (N_10910,N_9172,N_9809);
nor U10911 (N_10911,N_9974,N_9387);
xor U10912 (N_10912,N_9521,N_9876);
nor U10913 (N_10913,N_9054,N_9604);
xor U10914 (N_10914,N_9083,N_9832);
nor U10915 (N_10915,N_9473,N_9229);
nor U10916 (N_10916,N_9430,N_9956);
xor U10917 (N_10917,N_9482,N_9134);
or U10918 (N_10918,N_9415,N_9481);
nor U10919 (N_10919,N_9432,N_9729);
nand U10920 (N_10920,N_9832,N_9757);
nand U10921 (N_10921,N_9929,N_9626);
xor U10922 (N_10922,N_9211,N_9218);
nor U10923 (N_10923,N_9621,N_9362);
or U10924 (N_10924,N_9748,N_9008);
nand U10925 (N_10925,N_9111,N_9968);
xor U10926 (N_10926,N_9851,N_9835);
xnor U10927 (N_10927,N_9629,N_9549);
nand U10928 (N_10928,N_9443,N_9775);
nand U10929 (N_10929,N_9781,N_9656);
xnor U10930 (N_10930,N_9564,N_9894);
nor U10931 (N_10931,N_9557,N_9462);
nand U10932 (N_10932,N_9239,N_9454);
and U10933 (N_10933,N_9895,N_9225);
xor U10934 (N_10934,N_9816,N_9827);
nand U10935 (N_10935,N_9081,N_9452);
nor U10936 (N_10936,N_9022,N_9152);
xnor U10937 (N_10937,N_9572,N_9063);
xor U10938 (N_10938,N_9616,N_9053);
nor U10939 (N_10939,N_9625,N_9816);
and U10940 (N_10940,N_9656,N_9472);
or U10941 (N_10941,N_9942,N_9489);
or U10942 (N_10942,N_9257,N_9145);
nand U10943 (N_10943,N_9861,N_9776);
and U10944 (N_10944,N_9532,N_9940);
or U10945 (N_10945,N_9100,N_9432);
nand U10946 (N_10946,N_9264,N_9227);
or U10947 (N_10947,N_9146,N_9835);
xnor U10948 (N_10948,N_9239,N_9403);
and U10949 (N_10949,N_9218,N_9080);
nand U10950 (N_10950,N_9626,N_9890);
nand U10951 (N_10951,N_9465,N_9179);
nor U10952 (N_10952,N_9984,N_9680);
or U10953 (N_10953,N_9505,N_9400);
or U10954 (N_10954,N_9698,N_9126);
xor U10955 (N_10955,N_9117,N_9743);
nor U10956 (N_10956,N_9764,N_9188);
xor U10957 (N_10957,N_9970,N_9844);
nand U10958 (N_10958,N_9208,N_9250);
nor U10959 (N_10959,N_9523,N_9604);
nand U10960 (N_10960,N_9206,N_9048);
nand U10961 (N_10961,N_9414,N_9246);
or U10962 (N_10962,N_9382,N_9755);
xnor U10963 (N_10963,N_9715,N_9250);
and U10964 (N_10964,N_9289,N_9999);
xnor U10965 (N_10965,N_9314,N_9981);
or U10966 (N_10966,N_9121,N_9769);
and U10967 (N_10967,N_9370,N_9202);
and U10968 (N_10968,N_9402,N_9541);
nor U10969 (N_10969,N_9388,N_9383);
nor U10970 (N_10970,N_9996,N_9284);
or U10971 (N_10971,N_9422,N_9019);
xor U10972 (N_10972,N_9910,N_9845);
and U10973 (N_10973,N_9999,N_9632);
and U10974 (N_10974,N_9676,N_9059);
and U10975 (N_10975,N_9593,N_9876);
and U10976 (N_10976,N_9127,N_9490);
and U10977 (N_10977,N_9822,N_9910);
nor U10978 (N_10978,N_9662,N_9144);
or U10979 (N_10979,N_9928,N_9147);
nor U10980 (N_10980,N_9634,N_9893);
or U10981 (N_10981,N_9336,N_9706);
or U10982 (N_10982,N_9260,N_9114);
nor U10983 (N_10983,N_9591,N_9149);
nand U10984 (N_10984,N_9624,N_9876);
and U10985 (N_10985,N_9361,N_9097);
and U10986 (N_10986,N_9286,N_9463);
nand U10987 (N_10987,N_9716,N_9884);
or U10988 (N_10988,N_9079,N_9475);
xnor U10989 (N_10989,N_9987,N_9350);
or U10990 (N_10990,N_9761,N_9894);
nor U10991 (N_10991,N_9933,N_9882);
nand U10992 (N_10992,N_9815,N_9150);
and U10993 (N_10993,N_9710,N_9359);
nor U10994 (N_10994,N_9324,N_9741);
and U10995 (N_10995,N_9484,N_9384);
nand U10996 (N_10996,N_9193,N_9753);
and U10997 (N_10997,N_9696,N_9990);
nor U10998 (N_10998,N_9796,N_9341);
and U10999 (N_10999,N_9466,N_9682);
nor U11000 (N_11000,N_10509,N_10038);
or U11001 (N_11001,N_10653,N_10778);
nor U11002 (N_11002,N_10947,N_10388);
or U11003 (N_11003,N_10696,N_10008);
nor U11004 (N_11004,N_10296,N_10689);
nor U11005 (N_11005,N_10578,N_10548);
xnor U11006 (N_11006,N_10723,N_10224);
or U11007 (N_11007,N_10032,N_10655);
or U11008 (N_11008,N_10671,N_10113);
and U11009 (N_11009,N_10773,N_10564);
nand U11010 (N_11010,N_10363,N_10739);
or U11011 (N_11011,N_10675,N_10594);
or U11012 (N_11012,N_10808,N_10169);
or U11013 (N_11013,N_10307,N_10584);
nor U11014 (N_11014,N_10275,N_10920);
nor U11015 (N_11015,N_10462,N_10428);
and U11016 (N_11016,N_10801,N_10716);
nor U11017 (N_11017,N_10811,N_10108);
nor U11018 (N_11018,N_10768,N_10081);
nand U11019 (N_11019,N_10238,N_10846);
or U11020 (N_11020,N_10974,N_10112);
and U11021 (N_11021,N_10941,N_10193);
and U11022 (N_11022,N_10088,N_10771);
and U11023 (N_11023,N_10810,N_10484);
and U11024 (N_11024,N_10711,N_10332);
nor U11025 (N_11025,N_10178,N_10944);
nand U11026 (N_11026,N_10841,N_10018);
and U11027 (N_11027,N_10701,N_10954);
xnor U11028 (N_11028,N_10328,N_10987);
nor U11029 (N_11029,N_10119,N_10699);
nand U11030 (N_11030,N_10629,N_10159);
or U11031 (N_11031,N_10177,N_10499);
nor U11032 (N_11032,N_10391,N_10639);
and U11033 (N_11033,N_10382,N_10805);
or U11034 (N_11034,N_10134,N_10641);
nand U11035 (N_11035,N_10073,N_10375);
nand U11036 (N_11036,N_10361,N_10826);
xnor U11037 (N_11037,N_10515,N_10117);
and U11038 (N_11038,N_10116,N_10637);
and U11039 (N_11039,N_10676,N_10445);
and U11040 (N_11040,N_10403,N_10942);
xor U11041 (N_11041,N_10573,N_10853);
xor U11042 (N_11042,N_10604,N_10949);
and U11043 (N_11043,N_10836,N_10333);
xor U11044 (N_11044,N_10223,N_10734);
and U11045 (N_11045,N_10225,N_10442);
and U11046 (N_11046,N_10906,N_10353);
and U11047 (N_11047,N_10550,N_10083);
nand U11048 (N_11048,N_10383,N_10247);
and U11049 (N_11049,N_10522,N_10967);
xor U11050 (N_11050,N_10369,N_10389);
xnor U11051 (N_11051,N_10064,N_10397);
nand U11052 (N_11052,N_10819,N_10135);
or U11053 (N_11053,N_10301,N_10347);
and U11054 (N_11054,N_10783,N_10562);
or U11055 (N_11055,N_10843,N_10964);
and U11056 (N_11056,N_10276,N_10877);
nor U11057 (N_11057,N_10960,N_10386);
nor U11058 (N_11058,N_10308,N_10228);
nand U11059 (N_11059,N_10845,N_10208);
nand U11060 (N_11060,N_10343,N_10483);
nor U11061 (N_11061,N_10682,N_10700);
nand U11062 (N_11062,N_10965,N_10776);
xnor U11063 (N_11063,N_10005,N_10248);
xor U11064 (N_11064,N_10022,N_10530);
or U11065 (N_11065,N_10226,N_10645);
or U11066 (N_11066,N_10561,N_10980);
nand U11067 (N_11067,N_10172,N_10058);
xnor U11068 (N_11068,N_10235,N_10541);
and U11069 (N_11069,N_10636,N_10236);
and U11070 (N_11070,N_10385,N_10529);
nor U11071 (N_11071,N_10207,N_10340);
nor U11072 (N_11072,N_10714,N_10534);
or U11073 (N_11073,N_10638,N_10749);
nor U11074 (N_11074,N_10571,N_10926);
nand U11075 (N_11075,N_10559,N_10179);
or U11076 (N_11076,N_10455,N_10016);
xnor U11077 (N_11077,N_10762,N_10922);
or U11078 (N_11078,N_10693,N_10733);
and U11079 (N_11079,N_10062,N_10485);
and U11080 (N_11080,N_10697,N_10684);
nand U11081 (N_11081,N_10630,N_10068);
or U11082 (N_11082,N_10292,N_10842);
nor U11083 (N_11083,N_10525,N_10628);
xor U11084 (N_11084,N_10261,N_10643);
or U11085 (N_11085,N_10972,N_10360);
nor U11086 (N_11086,N_10601,N_10191);
and U11087 (N_11087,N_10616,N_10910);
nor U11088 (N_11088,N_10271,N_10996);
nor U11089 (N_11089,N_10463,N_10829);
or U11090 (N_11090,N_10872,N_10313);
and U11091 (N_11091,N_10283,N_10527);
nand U11092 (N_11092,N_10803,N_10162);
nand U11093 (N_11093,N_10344,N_10907);
nand U11094 (N_11094,N_10582,N_10322);
nor U11095 (N_11095,N_10297,N_10401);
xor U11096 (N_11096,N_10129,N_10726);
nor U11097 (N_11097,N_10955,N_10913);
nor U11098 (N_11098,N_10874,N_10427);
or U11099 (N_11099,N_10690,N_10417);
nor U11100 (N_11100,N_10037,N_10839);
or U11101 (N_11101,N_10153,N_10649);
nor U11102 (N_11102,N_10379,N_10267);
nand U11103 (N_11103,N_10665,N_10531);
nand U11104 (N_11104,N_10731,N_10759);
or U11105 (N_11105,N_10909,N_10123);
and U11106 (N_11106,N_10863,N_10652);
and U11107 (N_11107,N_10013,N_10378);
or U11108 (N_11108,N_10888,N_10494);
nand U11109 (N_11109,N_10609,N_10999);
xor U11110 (N_11110,N_10537,N_10291);
or U11111 (N_11111,N_10034,N_10774);
or U11112 (N_11112,N_10983,N_10285);
nand U11113 (N_11113,N_10078,N_10859);
nand U11114 (N_11114,N_10651,N_10785);
and U11115 (N_11115,N_10747,N_10758);
and U11116 (N_11116,N_10688,N_10981);
nor U11117 (N_11117,N_10978,N_10356);
nand U11118 (N_11118,N_10806,N_10051);
xor U11119 (N_11119,N_10583,N_10122);
and U11120 (N_11120,N_10368,N_10138);
nor U11121 (N_11121,N_10273,N_10456);
xnor U11122 (N_11122,N_10925,N_10047);
or U11123 (N_11123,N_10089,N_10049);
or U11124 (N_11124,N_10033,N_10305);
xor U11125 (N_11125,N_10059,N_10928);
or U11126 (N_11126,N_10765,N_10656);
nor U11127 (N_11127,N_10937,N_10526);
nor U11128 (N_11128,N_10359,N_10735);
xor U11129 (N_11129,N_10433,N_10258);
or U11130 (N_11130,N_10622,N_10195);
xor U11131 (N_11131,N_10779,N_10498);
xor U11132 (N_11132,N_10658,N_10997);
nand U11133 (N_11133,N_10569,N_10756);
xor U11134 (N_11134,N_10431,N_10255);
or U11135 (N_11135,N_10495,N_10067);
nor U11136 (N_11136,N_10439,N_10788);
nand U11137 (N_11137,N_10411,N_10099);
nor U11138 (N_11138,N_10448,N_10634);
xnor U11139 (N_11139,N_10310,N_10931);
or U11140 (N_11140,N_10396,N_10336);
xor U11141 (N_11141,N_10398,N_10740);
nand U11142 (N_11142,N_10082,N_10745);
or U11143 (N_11143,N_10746,N_10592);
and U11144 (N_11144,N_10199,N_10659);
xnor U11145 (N_11145,N_10024,N_10597);
and U11146 (N_11146,N_10449,N_10470);
or U11147 (N_11147,N_10174,N_10511);
xnor U11148 (N_11148,N_10063,N_10580);
or U11149 (N_11149,N_10799,N_10602);
xnor U11150 (N_11150,N_10642,N_10466);
xor U11151 (N_11151,N_10306,N_10702);
xor U11152 (N_11152,N_10464,N_10270);
nor U11153 (N_11153,N_10975,N_10281);
xnor U11154 (N_11154,N_10905,N_10355);
and U11155 (N_11155,N_10572,N_10852);
nor U11156 (N_11156,N_10514,N_10370);
nand U11157 (N_11157,N_10492,N_10314);
or U11158 (N_11158,N_10465,N_10738);
or U11159 (N_11159,N_10932,N_10019);
and U11160 (N_11160,N_10670,N_10753);
or U11161 (N_11161,N_10927,N_10460);
nor U11162 (N_11162,N_10175,N_10898);
nand U11163 (N_11163,N_10341,N_10085);
nand U11164 (N_11164,N_10394,N_10600);
xor U11165 (N_11165,N_10831,N_10181);
nand U11166 (N_11166,N_10298,N_10613);
and U11167 (N_11167,N_10402,N_10007);
or U11168 (N_11168,N_10407,N_10482);
xnor U11169 (N_11169,N_10239,N_10069);
or U11170 (N_11170,N_10563,N_10393);
xor U11171 (N_11171,N_10707,N_10538);
or U11172 (N_11172,N_10854,N_10923);
or U11173 (N_11173,N_10290,N_10025);
nand U11174 (N_11174,N_10948,N_10751);
or U11175 (N_11175,N_10868,N_10994);
or U11176 (N_11176,N_10269,N_10554);
or U11177 (N_11177,N_10775,N_10809);
or U11178 (N_11178,N_10166,N_10125);
and U11179 (N_11179,N_10415,N_10160);
xnor U11180 (N_11180,N_10777,N_10211);
or U11181 (N_11181,N_10251,N_10071);
xor U11182 (N_11182,N_10512,N_10246);
xnor U11183 (N_11183,N_10677,N_10787);
or U11184 (N_11184,N_10705,N_10621);
nand U11185 (N_11185,N_10995,N_10004);
xor U11186 (N_11186,N_10681,N_10508);
xnor U11187 (N_11187,N_10331,N_10184);
or U11188 (N_11188,N_10856,N_10094);
or U11189 (N_11189,N_10757,N_10743);
and U11190 (N_11190,N_10327,N_10061);
xnor U11191 (N_11191,N_10354,N_10611);
nand U11192 (N_11192,N_10136,N_10535);
or U11193 (N_11193,N_10533,N_10031);
and U11194 (N_11194,N_10197,N_10486);
xor U11195 (N_11195,N_10915,N_10084);
and U11196 (N_11196,N_10828,N_10077);
nor U11197 (N_11197,N_10882,N_10458);
and U11198 (N_11198,N_10302,N_10443);
nand U11199 (N_11199,N_10097,N_10374);
nor U11200 (N_11200,N_10647,N_10752);
nand U11201 (N_11201,N_10424,N_10631);
or U11202 (N_11202,N_10834,N_10447);
and U11203 (N_11203,N_10311,N_10823);
and U11204 (N_11204,N_10991,N_10971);
nor U11205 (N_11205,N_10265,N_10661);
nor U11206 (N_11206,N_10770,N_10887);
nor U11207 (N_11207,N_10423,N_10115);
nor U11208 (N_11208,N_10667,N_10549);
nor U11209 (N_11209,N_10605,N_10568);
nand U11210 (N_11210,N_10507,N_10412);
and U11211 (N_11211,N_10657,N_10586);
nand U11212 (N_11212,N_10692,N_10012);
nand U11213 (N_11213,N_10452,N_10858);
xnor U11214 (N_11214,N_10760,N_10233);
or U11215 (N_11215,N_10718,N_10674);
nand U11216 (N_11216,N_10504,N_10536);
or U11217 (N_11217,N_10426,N_10221);
nand U11218 (N_11218,N_10748,N_10729);
xnor U11219 (N_11219,N_10154,N_10190);
nand U11220 (N_11220,N_10708,N_10838);
and U11221 (N_11221,N_10933,N_10489);
nor U11222 (N_11222,N_10903,N_10654);
xor U11223 (N_11223,N_10080,N_10772);
nand U11224 (N_11224,N_10544,N_10695);
and U11225 (N_11225,N_10791,N_10827);
nand U11226 (N_11226,N_10950,N_10349);
or U11227 (N_11227,N_10074,N_10704);
nor U11228 (N_11228,N_10876,N_10880);
and U11229 (N_11229,N_10889,N_10698);
and U11230 (N_11230,N_10282,N_10176);
nor U11231 (N_11231,N_10053,N_10057);
xnor U11232 (N_11232,N_10976,N_10979);
nand U11233 (N_11233,N_10241,N_10144);
and U11234 (N_11234,N_10713,N_10202);
and U11235 (N_11235,N_10435,N_10867);
nor U11236 (N_11236,N_10339,N_10384);
xnor U11237 (N_11237,N_10902,N_10625);
and U11238 (N_11238,N_10103,N_10227);
and U11239 (N_11239,N_10660,N_10802);
xor U11240 (N_11240,N_10576,N_10546);
and U11241 (N_11241,N_10883,N_10096);
xnor U11242 (N_11242,N_10266,N_10646);
xnor U11243 (N_11243,N_10410,N_10141);
nand U11244 (N_11244,N_10633,N_10721);
nand U11245 (N_11245,N_10262,N_10471);
or U11246 (N_11246,N_10052,N_10516);
xor U11247 (N_11247,N_10687,N_10977);
nand U11248 (N_11248,N_10217,N_10167);
xnor U11249 (N_11249,N_10814,N_10041);
nand U11250 (N_11250,N_10895,N_10408);
and U11251 (N_11251,N_10234,N_10079);
nand U11252 (N_11252,N_10173,N_10672);
nand U11253 (N_11253,N_10943,N_10365);
or U11254 (N_11254,N_10381,N_10505);
nor U11255 (N_11255,N_10627,N_10142);
nand U11256 (N_11256,N_10371,N_10185);
and U11257 (N_11257,N_10151,N_10086);
nand U11258 (N_11258,N_10253,N_10553);
and U11259 (N_11259,N_10107,N_10866);
or U11260 (N_11260,N_10496,N_10973);
or U11261 (N_11261,N_10250,N_10524);
and U11262 (N_11262,N_10724,N_10316);
and U11263 (N_11263,N_10145,N_10334);
nor U11264 (N_11264,N_10120,N_10720);
and U11265 (N_11265,N_10780,N_10881);
xor U11266 (N_11266,N_10992,N_10924);
or U11267 (N_11267,N_10404,N_10300);
xor U11268 (N_11268,N_10848,N_10219);
and U11269 (N_11269,N_10497,N_10329);
xnor U11270 (N_11270,N_10350,N_10886);
nor U11271 (N_11271,N_10792,N_10087);
xnor U11272 (N_11272,N_10457,N_10446);
or U11273 (N_11273,N_10294,N_10044);
nor U11274 (N_11274,N_10000,N_10143);
or U11275 (N_11275,N_10590,N_10884);
nand U11276 (N_11276,N_10348,N_10567);
or U11277 (N_11277,N_10459,N_10472);
nor U11278 (N_11278,N_10104,N_10147);
nor U11279 (N_11279,N_10767,N_10490);
nor U11280 (N_11280,N_10132,N_10532);
or U11281 (N_11281,N_10798,N_10683);
and U11282 (N_11282,N_10952,N_10970);
and U11283 (N_11283,N_10897,N_10837);
and U11284 (N_11284,N_10338,N_10990);
and U11285 (N_11285,N_10229,N_10844);
or U11286 (N_11286,N_10284,N_10440);
nor U11287 (N_11287,N_10418,N_10958);
nand U11288 (N_11288,N_10409,N_10252);
nand U11289 (N_11289,N_10986,N_10437);
and U11290 (N_11290,N_10560,N_10055);
nor U11291 (N_11291,N_10890,N_10686);
or U11292 (N_11292,N_10635,N_10669);
xor U11293 (N_11293,N_10542,N_10824);
and U11294 (N_11294,N_10029,N_10161);
xor U11295 (N_11295,N_10121,N_10030);
and U11296 (N_11296,N_10304,N_10650);
nand U11297 (N_11297,N_10694,N_10373);
xnor U11298 (N_11298,N_10878,N_10392);
xor U11299 (N_11299,N_10441,N_10817);
and U11300 (N_11300,N_10818,N_10425);
xnor U11301 (N_11301,N_10422,N_10766);
xor U11302 (N_11302,N_10790,N_10170);
nor U11303 (N_11303,N_10820,N_10709);
or U11304 (N_11304,N_10864,N_10213);
and U11305 (N_11305,N_10277,N_10163);
or U11306 (N_11306,N_10557,N_10414);
or U11307 (N_11307,N_10101,N_10124);
nand U11308 (N_11308,N_10581,N_10565);
or U11309 (N_11309,N_10632,N_10664);
or U11310 (N_11310,N_10244,N_10912);
and U11311 (N_11311,N_10454,N_10615);
or U11312 (N_11312,N_10959,N_10861);
nand U11313 (N_11313,N_10610,N_10938);
nand U11314 (N_11314,N_10014,N_10478);
nor U11315 (N_11315,N_10026,N_10501);
nor U11316 (N_11316,N_10678,N_10795);
nand U11317 (N_11317,N_10091,N_10130);
xor U11318 (N_11318,N_10502,N_10040);
or U11319 (N_11319,N_10619,N_10009);
xor U11320 (N_11320,N_10968,N_10624);
nand U11321 (N_11321,N_10474,N_10797);
and U11322 (N_11322,N_10862,N_10969);
and U11323 (N_11323,N_10286,N_10075);
xor U11324 (N_11324,N_10951,N_10367);
and U11325 (N_11325,N_10476,N_10242);
xnor U11326 (N_11326,N_10873,N_10137);
xnor U11327 (N_11327,N_10555,N_10725);
nor U11328 (N_11328,N_10194,N_10781);
and U11329 (N_11329,N_10825,N_10988);
nor U11330 (N_11330,N_10894,N_10315);
and U11331 (N_11331,N_10395,N_10830);
nor U11332 (N_11332,N_10140,N_10763);
nand U11333 (N_11333,N_10764,N_10732);
or U11334 (N_11334,N_10021,N_10114);
and U11335 (N_11335,N_10946,N_10146);
nor U11336 (N_11336,N_10351,N_10256);
xor U11337 (N_11337,N_10750,N_10608);
xnor U11338 (N_11338,N_10222,N_10607);
and U11339 (N_11339,N_10940,N_10626);
and U11340 (N_11340,N_10280,N_10278);
and U11341 (N_11341,N_10680,N_10183);
nor U11342 (N_11342,N_10187,N_10011);
and U11343 (N_11343,N_10406,N_10919);
or U11344 (N_11344,N_10324,N_10345);
or U11345 (N_11345,N_10488,N_10467);
or U11346 (N_11346,N_10200,N_10003);
nor U11347 (N_11347,N_10358,N_10118);
nand U11348 (N_11348,N_10438,N_10293);
and U11349 (N_11349,N_10755,N_10761);
nand U11350 (N_11350,N_10742,N_10728);
nor U11351 (N_11351,N_10899,N_10254);
xnor U11352 (N_11352,N_10865,N_10171);
and U11353 (N_11353,N_10450,N_10963);
nand U11354 (N_11354,N_10218,N_10127);
xnor U11355 (N_11355,N_10620,N_10685);
nor U11356 (N_11356,N_10673,N_10429);
xnor U11357 (N_11357,N_10551,N_10547);
or U11358 (N_11358,N_10110,N_10822);
and U11359 (N_11359,N_10871,N_10962);
nor U11360 (N_11360,N_10585,N_10796);
nand U11361 (N_11361,N_10741,N_10691);
and U11362 (N_11362,N_10230,N_10299);
nor U11363 (N_11363,N_10513,N_10432);
and U11364 (N_11364,N_10896,N_10556);
and U11365 (N_11365,N_10575,N_10196);
xnor U11366 (N_11366,N_10921,N_10090);
nor U11367 (N_11367,N_10045,N_10027);
nor U11368 (N_11368,N_10020,N_10993);
nor U11369 (N_11369,N_10066,N_10966);
nand U11370 (N_11370,N_10939,N_10832);
or U11371 (N_11371,N_10220,N_10566);
and U11372 (N_11372,N_10203,N_10891);
nand U11373 (N_11373,N_10212,N_10070);
and U11374 (N_11374,N_10249,N_10870);
and U11375 (N_11375,N_10272,N_10420);
xnor U11376 (N_11376,N_10419,N_10596);
or U11377 (N_11377,N_10072,N_10481);
and U11378 (N_11378,N_10475,N_10444);
and U11379 (N_11379,N_10093,N_10376);
and U11380 (N_11380,N_10469,N_10599);
nand U11381 (N_11381,N_10390,N_10679);
nor U11382 (N_11382,N_10893,N_10500);
and U11383 (N_11383,N_10287,N_10054);
nor U11384 (N_11384,N_10804,N_10539);
or U11385 (N_11385,N_10982,N_10754);
xnor U11386 (N_11386,N_10028,N_10156);
or U11387 (N_11387,N_10710,N_10917);
nor U11388 (N_11388,N_10663,N_10321);
nand U11389 (N_11389,N_10042,N_10914);
and U11390 (N_11390,N_10158,N_10023);
nand U11391 (N_11391,N_10612,N_10387);
nand U11392 (N_11392,N_10984,N_10317);
xnor U11393 (N_11393,N_10043,N_10662);
nand U11394 (N_11394,N_10320,N_10519);
and U11395 (N_11395,N_10152,N_10606);
xor U11396 (N_11396,N_10303,N_10342);
and U11397 (N_11397,N_10813,N_10189);
and U11398 (N_11398,N_10257,N_10517);
or U11399 (N_11399,N_10480,N_10060);
or U11400 (N_11400,N_10468,N_10216);
or U11401 (N_11401,N_10849,N_10518);
nor U11402 (N_11402,N_10295,N_10434);
nand U11403 (N_11403,N_10623,N_10214);
nor U11404 (N_11404,N_10929,N_10364);
or U11405 (N_11405,N_10477,N_10237);
and U11406 (N_11406,N_10784,N_10840);
nor U11407 (N_11407,N_10352,N_10243);
nor U11408 (N_11408,N_10209,N_10719);
nand U11409 (N_11409,N_10240,N_10892);
nand U11410 (N_11410,N_10001,N_10105);
and U11411 (N_11411,N_10400,N_10050);
or U11412 (N_11412,N_10436,N_10591);
and U11413 (N_11413,N_10100,N_10377);
and U11414 (N_11414,N_10198,N_10815);
and U11415 (N_11415,N_10510,N_10319);
nor U11416 (N_11416,N_10111,N_10380);
xnor U11417 (N_11417,N_10180,N_10205);
and U11418 (N_11418,N_10288,N_10076);
and U11419 (N_11419,N_10330,N_10421);
nand U11420 (N_11420,N_10847,N_10192);
or U11421 (N_11421,N_10528,N_10617);
and U11422 (N_11422,N_10065,N_10812);
nand U11423 (N_11423,N_10493,N_10413);
xor U11424 (N_11424,N_10574,N_10794);
nor U11425 (N_11425,N_10260,N_10264);
or U11426 (N_11426,N_10133,N_10911);
nor U11427 (N_11427,N_10786,N_10570);
and U11428 (N_11428,N_10587,N_10487);
or U11429 (N_11429,N_10835,N_10523);
nand U11430 (N_11430,N_10325,N_10268);
and U11431 (N_11431,N_10399,N_10357);
xnor U11432 (N_11432,N_10540,N_10552);
xnor U11433 (N_11433,N_10961,N_10901);
xnor U11434 (N_11434,N_10312,N_10139);
nand U11435 (N_11435,N_10577,N_10855);
nor U11436 (N_11436,N_10155,N_10945);
and U11437 (N_11437,N_10935,N_10821);
nor U11438 (N_11438,N_10109,N_10461);
or U11439 (N_11439,N_10793,N_10956);
xnor U11440 (N_11440,N_10588,N_10875);
nand U11441 (N_11441,N_10039,N_10231);
and U11442 (N_11442,N_10479,N_10614);
xnor U11443 (N_11443,N_10201,N_10128);
nand U11444 (N_11444,N_10263,N_10727);
nor U11445 (N_11445,N_10782,N_10860);
and U11446 (N_11446,N_10098,N_10908);
and U11447 (N_11447,N_10885,N_10430);
nor U11448 (N_11448,N_10916,N_10279);
nand U11449 (N_11449,N_10451,N_10372);
nor U11450 (N_11450,N_10712,N_10953);
nand U11451 (N_11451,N_10595,N_10545);
xor U11452 (N_11452,N_10930,N_10035);
and U11453 (N_11453,N_10593,N_10668);
or U11454 (N_11454,N_10206,N_10807);
nor U11455 (N_11455,N_10603,N_10589);
nand U11456 (N_11456,N_10816,N_10850);
and U11457 (N_11457,N_10833,N_10405);
or U11458 (N_11458,N_10644,N_10346);
or U11459 (N_11459,N_10289,N_10274);
or U11460 (N_11460,N_10362,N_10337);
xor U11461 (N_11461,N_10232,N_10204);
nor U11462 (N_11462,N_10648,N_10900);
xnor U11463 (N_11463,N_10168,N_10736);
nand U11464 (N_11464,N_10106,N_10598);
or U11465 (N_11465,N_10131,N_10998);
xor U11466 (N_11466,N_10416,N_10717);
nor U11467 (N_11467,N_10095,N_10165);
and U11468 (N_11468,N_10318,N_10002);
nor U11469 (N_11469,N_10186,N_10046);
nand U11470 (N_11470,N_10879,N_10744);
or U11471 (N_11471,N_10126,N_10706);
or U11472 (N_11472,N_10769,N_10157);
and U11473 (N_11473,N_10326,N_10010);
nor U11474 (N_11474,N_10640,N_10666);
nand U11475 (N_11475,N_10309,N_10904);
xnor U11476 (N_11476,N_10015,N_10215);
and U11477 (N_11477,N_10715,N_10164);
nor U11478 (N_11478,N_10543,N_10558);
and U11479 (N_11479,N_10323,N_10918);
nand U11480 (N_11480,N_10789,N_10210);
nor U11481 (N_11481,N_10150,N_10036);
nand U11482 (N_11482,N_10869,N_10453);
or U11483 (N_11483,N_10985,N_10102);
nand U11484 (N_11484,N_10366,N_10934);
and U11485 (N_11485,N_10957,N_10017);
nand U11486 (N_11486,N_10506,N_10188);
xor U11487 (N_11487,N_10851,N_10936);
nand U11488 (N_11488,N_10800,N_10473);
nor U11489 (N_11489,N_10730,N_10722);
and U11490 (N_11490,N_10703,N_10737);
and U11491 (N_11491,N_10520,N_10259);
nand U11492 (N_11492,N_10521,N_10048);
nand U11493 (N_11493,N_10503,N_10989);
xnor U11494 (N_11494,N_10092,N_10618);
and U11495 (N_11495,N_10149,N_10006);
nor U11496 (N_11496,N_10245,N_10148);
and U11497 (N_11497,N_10335,N_10056);
xnor U11498 (N_11498,N_10857,N_10182);
and U11499 (N_11499,N_10579,N_10491);
xor U11500 (N_11500,N_10484,N_10749);
nor U11501 (N_11501,N_10724,N_10725);
nor U11502 (N_11502,N_10037,N_10173);
or U11503 (N_11503,N_10126,N_10792);
and U11504 (N_11504,N_10678,N_10348);
or U11505 (N_11505,N_10055,N_10298);
nand U11506 (N_11506,N_10024,N_10444);
and U11507 (N_11507,N_10700,N_10420);
nand U11508 (N_11508,N_10780,N_10524);
and U11509 (N_11509,N_10662,N_10658);
and U11510 (N_11510,N_10561,N_10126);
and U11511 (N_11511,N_10137,N_10513);
nor U11512 (N_11512,N_10206,N_10776);
xnor U11513 (N_11513,N_10123,N_10526);
xor U11514 (N_11514,N_10783,N_10482);
and U11515 (N_11515,N_10128,N_10782);
nor U11516 (N_11516,N_10217,N_10231);
and U11517 (N_11517,N_10784,N_10410);
nor U11518 (N_11518,N_10548,N_10261);
xnor U11519 (N_11519,N_10040,N_10295);
nor U11520 (N_11520,N_10135,N_10808);
and U11521 (N_11521,N_10435,N_10136);
nand U11522 (N_11522,N_10009,N_10804);
and U11523 (N_11523,N_10107,N_10173);
xnor U11524 (N_11524,N_10917,N_10355);
xor U11525 (N_11525,N_10244,N_10171);
nand U11526 (N_11526,N_10592,N_10458);
or U11527 (N_11527,N_10735,N_10392);
nand U11528 (N_11528,N_10454,N_10114);
and U11529 (N_11529,N_10183,N_10321);
or U11530 (N_11530,N_10513,N_10064);
and U11531 (N_11531,N_10106,N_10935);
nand U11532 (N_11532,N_10432,N_10948);
or U11533 (N_11533,N_10675,N_10869);
and U11534 (N_11534,N_10471,N_10442);
and U11535 (N_11535,N_10841,N_10862);
nor U11536 (N_11536,N_10261,N_10336);
nor U11537 (N_11537,N_10796,N_10222);
xor U11538 (N_11538,N_10121,N_10696);
xnor U11539 (N_11539,N_10027,N_10904);
and U11540 (N_11540,N_10995,N_10095);
and U11541 (N_11541,N_10535,N_10811);
and U11542 (N_11542,N_10009,N_10127);
nand U11543 (N_11543,N_10004,N_10360);
and U11544 (N_11544,N_10506,N_10207);
xor U11545 (N_11545,N_10003,N_10767);
nor U11546 (N_11546,N_10957,N_10747);
or U11547 (N_11547,N_10933,N_10530);
and U11548 (N_11548,N_10289,N_10313);
and U11549 (N_11549,N_10890,N_10728);
and U11550 (N_11550,N_10429,N_10692);
and U11551 (N_11551,N_10873,N_10562);
xor U11552 (N_11552,N_10253,N_10318);
xor U11553 (N_11553,N_10405,N_10259);
and U11554 (N_11554,N_10104,N_10656);
or U11555 (N_11555,N_10072,N_10203);
nor U11556 (N_11556,N_10354,N_10669);
nand U11557 (N_11557,N_10777,N_10674);
nand U11558 (N_11558,N_10562,N_10302);
nor U11559 (N_11559,N_10653,N_10538);
nand U11560 (N_11560,N_10196,N_10182);
nand U11561 (N_11561,N_10036,N_10760);
and U11562 (N_11562,N_10445,N_10755);
nor U11563 (N_11563,N_10962,N_10052);
and U11564 (N_11564,N_10931,N_10471);
and U11565 (N_11565,N_10146,N_10058);
xor U11566 (N_11566,N_10672,N_10473);
nand U11567 (N_11567,N_10930,N_10212);
nand U11568 (N_11568,N_10406,N_10257);
xnor U11569 (N_11569,N_10896,N_10669);
or U11570 (N_11570,N_10706,N_10837);
or U11571 (N_11571,N_10088,N_10010);
and U11572 (N_11572,N_10683,N_10742);
or U11573 (N_11573,N_10981,N_10067);
nand U11574 (N_11574,N_10833,N_10083);
and U11575 (N_11575,N_10888,N_10394);
nand U11576 (N_11576,N_10099,N_10345);
or U11577 (N_11577,N_10566,N_10823);
nor U11578 (N_11578,N_10375,N_10645);
nor U11579 (N_11579,N_10708,N_10367);
or U11580 (N_11580,N_10886,N_10060);
and U11581 (N_11581,N_10307,N_10712);
nor U11582 (N_11582,N_10830,N_10773);
and U11583 (N_11583,N_10615,N_10480);
or U11584 (N_11584,N_10387,N_10774);
nor U11585 (N_11585,N_10253,N_10483);
and U11586 (N_11586,N_10025,N_10591);
and U11587 (N_11587,N_10984,N_10290);
xor U11588 (N_11588,N_10897,N_10942);
and U11589 (N_11589,N_10673,N_10557);
and U11590 (N_11590,N_10281,N_10395);
or U11591 (N_11591,N_10558,N_10841);
and U11592 (N_11592,N_10740,N_10930);
and U11593 (N_11593,N_10091,N_10541);
or U11594 (N_11594,N_10883,N_10038);
xnor U11595 (N_11595,N_10340,N_10542);
xor U11596 (N_11596,N_10060,N_10558);
xnor U11597 (N_11597,N_10740,N_10753);
xnor U11598 (N_11598,N_10815,N_10100);
xnor U11599 (N_11599,N_10118,N_10002);
xnor U11600 (N_11600,N_10461,N_10943);
nand U11601 (N_11601,N_10243,N_10437);
and U11602 (N_11602,N_10247,N_10448);
nand U11603 (N_11603,N_10951,N_10065);
or U11604 (N_11604,N_10755,N_10473);
nor U11605 (N_11605,N_10829,N_10750);
xor U11606 (N_11606,N_10792,N_10733);
and U11607 (N_11607,N_10339,N_10166);
xor U11608 (N_11608,N_10343,N_10255);
nor U11609 (N_11609,N_10707,N_10698);
nor U11610 (N_11610,N_10306,N_10725);
or U11611 (N_11611,N_10884,N_10710);
or U11612 (N_11612,N_10173,N_10955);
xnor U11613 (N_11613,N_10073,N_10107);
nor U11614 (N_11614,N_10720,N_10894);
nand U11615 (N_11615,N_10344,N_10661);
and U11616 (N_11616,N_10655,N_10111);
nand U11617 (N_11617,N_10509,N_10255);
nor U11618 (N_11618,N_10559,N_10584);
nand U11619 (N_11619,N_10879,N_10905);
nand U11620 (N_11620,N_10728,N_10678);
xnor U11621 (N_11621,N_10022,N_10431);
xnor U11622 (N_11622,N_10865,N_10505);
nor U11623 (N_11623,N_10773,N_10496);
xnor U11624 (N_11624,N_10737,N_10589);
xor U11625 (N_11625,N_10381,N_10251);
xnor U11626 (N_11626,N_10065,N_10080);
nand U11627 (N_11627,N_10749,N_10550);
and U11628 (N_11628,N_10226,N_10980);
nor U11629 (N_11629,N_10831,N_10744);
nand U11630 (N_11630,N_10566,N_10799);
or U11631 (N_11631,N_10710,N_10509);
nand U11632 (N_11632,N_10305,N_10198);
and U11633 (N_11633,N_10402,N_10523);
nand U11634 (N_11634,N_10084,N_10151);
nand U11635 (N_11635,N_10559,N_10907);
or U11636 (N_11636,N_10795,N_10812);
and U11637 (N_11637,N_10252,N_10177);
nand U11638 (N_11638,N_10225,N_10556);
xor U11639 (N_11639,N_10487,N_10006);
or U11640 (N_11640,N_10235,N_10138);
and U11641 (N_11641,N_10591,N_10855);
and U11642 (N_11642,N_10908,N_10065);
and U11643 (N_11643,N_10456,N_10237);
or U11644 (N_11644,N_10148,N_10118);
or U11645 (N_11645,N_10220,N_10427);
nand U11646 (N_11646,N_10701,N_10503);
xnor U11647 (N_11647,N_10108,N_10137);
or U11648 (N_11648,N_10704,N_10070);
nand U11649 (N_11649,N_10896,N_10737);
or U11650 (N_11650,N_10787,N_10589);
xnor U11651 (N_11651,N_10195,N_10802);
xor U11652 (N_11652,N_10082,N_10526);
xor U11653 (N_11653,N_10163,N_10276);
nand U11654 (N_11654,N_10448,N_10957);
and U11655 (N_11655,N_10205,N_10653);
nand U11656 (N_11656,N_10970,N_10372);
nand U11657 (N_11657,N_10699,N_10324);
and U11658 (N_11658,N_10899,N_10627);
nor U11659 (N_11659,N_10308,N_10478);
and U11660 (N_11660,N_10853,N_10378);
and U11661 (N_11661,N_10613,N_10167);
nand U11662 (N_11662,N_10579,N_10128);
nand U11663 (N_11663,N_10592,N_10132);
xor U11664 (N_11664,N_10657,N_10526);
nor U11665 (N_11665,N_10739,N_10654);
nor U11666 (N_11666,N_10346,N_10300);
nor U11667 (N_11667,N_10068,N_10929);
and U11668 (N_11668,N_10181,N_10548);
nand U11669 (N_11669,N_10827,N_10480);
nand U11670 (N_11670,N_10993,N_10092);
nor U11671 (N_11671,N_10079,N_10614);
xnor U11672 (N_11672,N_10857,N_10059);
nand U11673 (N_11673,N_10854,N_10029);
nand U11674 (N_11674,N_10371,N_10639);
or U11675 (N_11675,N_10857,N_10855);
or U11676 (N_11676,N_10527,N_10680);
or U11677 (N_11677,N_10464,N_10173);
xnor U11678 (N_11678,N_10792,N_10894);
xor U11679 (N_11679,N_10242,N_10614);
or U11680 (N_11680,N_10046,N_10769);
and U11681 (N_11681,N_10725,N_10304);
nor U11682 (N_11682,N_10481,N_10053);
or U11683 (N_11683,N_10945,N_10938);
and U11684 (N_11684,N_10611,N_10911);
and U11685 (N_11685,N_10363,N_10802);
xor U11686 (N_11686,N_10962,N_10881);
nand U11687 (N_11687,N_10424,N_10157);
nand U11688 (N_11688,N_10768,N_10578);
nor U11689 (N_11689,N_10863,N_10777);
xnor U11690 (N_11690,N_10966,N_10674);
nand U11691 (N_11691,N_10643,N_10169);
xnor U11692 (N_11692,N_10735,N_10950);
and U11693 (N_11693,N_10071,N_10907);
or U11694 (N_11694,N_10197,N_10404);
nor U11695 (N_11695,N_10818,N_10815);
nor U11696 (N_11696,N_10762,N_10071);
and U11697 (N_11697,N_10692,N_10878);
or U11698 (N_11698,N_10285,N_10243);
nor U11699 (N_11699,N_10548,N_10801);
nand U11700 (N_11700,N_10081,N_10951);
and U11701 (N_11701,N_10080,N_10928);
xnor U11702 (N_11702,N_10458,N_10589);
nand U11703 (N_11703,N_10055,N_10850);
xnor U11704 (N_11704,N_10951,N_10217);
and U11705 (N_11705,N_10677,N_10374);
nor U11706 (N_11706,N_10630,N_10685);
nor U11707 (N_11707,N_10352,N_10189);
and U11708 (N_11708,N_10518,N_10031);
or U11709 (N_11709,N_10581,N_10538);
nor U11710 (N_11710,N_10630,N_10869);
nor U11711 (N_11711,N_10733,N_10897);
xor U11712 (N_11712,N_10550,N_10539);
and U11713 (N_11713,N_10117,N_10364);
xnor U11714 (N_11714,N_10141,N_10500);
or U11715 (N_11715,N_10908,N_10838);
xor U11716 (N_11716,N_10837,N_10031);
xor U11717 (N_11717,N_10494,N_10601);
or U11718 (N_11718,N_10854,N_10311);
nand U11719 (N_11719,N_10950,N_10518);
or U11720 (N_11720,N_10155,N_10030);
and U11721 (N_11721,N_10080,N_10505);
nand U11722 (N_11722,N_10930,N_10647);
and U11723 (N_11723,N_10053,N_10438);
nor U11724 (N_11724,N_10433,N_10415);
nor U11725 (N_11725,N_10534,N_10170);
nor U11726 (N_11726,N_10602,N_10471);
or U11727 (N_11727,N_10641,N_10067);
nand U11728 (N_11728,N_10474,N_10901);
nand U11729 (N_11729,N_10462,N_10854);
nand U11730 (N_11730,N_10617,N_10276);
xor U11731 (N_11731,N_10474,N_10069);
nor U11732 (N_11732,N_10152,N_10690);
and U11733 (N_11733,N_10366,N_10847);
and U11734 (N_11734,N_10270,N_10304);
and U11735 (N_11735,N_10481,N_10287);
xnor U11736 (N_11736,N_10622,N_10138);
xor U11737 (N_11737,N_10835,N_10498);
xnor U11738 (N_11738,N_10031,N_10439);
nor U11739 (N_11739,N_10232,N_10838);
nor U11740 (N_11740,N_10012,N_10713);
nor U11741 (N_11741,N_10513,N_10604);
nand U11742 (N_11742,N_10138,N_10666);
xnor U11743 (N_11743,N_10462,N_10779);
nand U11744 (N_11744,N_10093,N_10768);
nor U11745 (N_11745,N_10452,N_10998);
nand U11746 (N_11746,N_10350,N_10896);
xor U11747 (N_11747,N_10578,N_10163);
nor U11748 (N_11748,N_10422,N_10669);
or U11749 (N_11749,N_10615,N_10911);
nand U11750 (N_11750,N_10412,N_10068);
nand U11751 (N_11751,N_10912,N_10513);
nor U11752 (N_11752,N_10216,N_10802);
xor U11753 (N_11753,N_10378,N_10863);
xor U11754 (N_11754,N_10457,N_10134);
or U11755 (N_11755,N_10479,N_10360);
nor U11756 (N_11756,N_10832,N_10710);
nand U11757 (N_11757,N_10063,N_10254);
nand U11758 (N_11758,N_10129,N_10923);
or U11759 (N_11759,N_10888,N_10382);
xnor U11760 (N_11760,N_10981,N_10629);
and U11761 (N_11761,N_10531,N_10332);
or U11762 (N_11762,N_10461,N_10610);
nor U11763 (N_11763,N_10481,N_10767);
and U11764 (N_11764,N_10335,N_10478);
nand U11765 (N_11765,N_10902,N_10426);
xor U11766 (N_11766,N_10754,N_10228);
nor U11767 (N_11767,N_10602,N_10525);
nor U11768 (N_11768,N_10920,N_10498);
or U11769 (N_11769,N_10067,N_10915);
or U11770 (N_11770,N_10827,N_10520);
or U11771 (N_11771,N_10469,N_10578);
nand U11772 (N_11772,N_10935,N_10144);
nand U11773 (N_11773,N_10891,N_10281);
xor U11774 (N_11774,N_10640,N_10102);
nor U11775 (N_11775,N_10799,N_10110);
or U11776 (N_11776,N_10777,N_10818);
nor U11777 (N_11777,N_10856,N_10911);
and U11778 (N_11778,N_10028,N_10408);
or U11779 (N_11779,N_10600,N_10264);
or U11780 (N_11780,N_10485,N_10747);
xnor U11781 (N_11781,N_10517,N_10404);
and U11782 (N_11782,N_10531,N_10997);
or U11783 (N_11783,N_10331,N_10495);
xnor U11784 (N_11784,N_10370,N_10343);
or U11785 (N_11785,N_10934,N_10962);
nor U11786 (N_11786,N_10375,N_10576);
nand U11787 (N_11787,N_10688,N_10729);
nor U11788 (N_11788,N_10722,N_10389);
nand U11789 (N_11789,N_10907,N_10763);
xnor U11790 (N_11790,N_10934,N_10555);
or U11791 (N_11791,N_10422,N_10900);
and U11792 (N_11792,N_10420,N_10617);
and U11793 (N_11793,N_10593,N_10561);
nor U11794 (N_11794,N_10523,N_10160);
and U11795 (N_11795,N_10985,N_10310);
xor U11796 (N_11796,N_10440,N_10409);
or U11797 (N_11797,N_10949,N_10998);
xor U11798 (N_11798,N_10726,N_10435);
and U11799 (N_11799,N_10732,N_10311);
xnor U11800 (N_11800,N_10730,N_10774);
and U11801 (N_11801,N_10895,N_10331);
nor U11802 (N_11802,N_10179,N_10162);
or U11803 (N_11803,N_10446,N_10897);
nand U11804 (N_11804,N_10976,N_10680);
nor U11805 (N_11805,N_10385,N_10747);
xnor U11806 (N_11806,N_10811,N_10291);
or U11807 (N_11807,N_10324,N_10913);
xor U11808 (N_11808,N_10067,N_10553);
nand U11809 (N_11809,N_10588,N_10263);
nor U11810 (N_11810,N_10007,N_10635);
nand U11811 (N_11811,N_10678,N_10134);
xor U11812 (N_11812,N_10153,N_10588);
nand U11813 (N_11813,N_10482,N_10828);
and U11814 (N_11814,N_10279,N_10346);
nand U11815 (N_11815,N_10540,N_10736);
xnor U11816 (N_11816,N_10416,N_10755);
xor U11817 (N_11817,N_10022,N_10754);
or U11818 (N_11818,N_10664,N_10363);
nand U11819 (N_11819,N_10406,N_10422);
nand U11820 (N_11820,N_10421,N_10667);
nor U11821 (N_11821,N_10530,N_10260);
nand U11822 (N_11822,N_10614,N_10483);
nand U11823 (N_11823,N_10704,N_10217);
nand U11824 (N_11824,N_10045,N_10627);
or U11825 (N_11825,N_10294,N_10891);
nor U11826 (N_11826,N_10349,N_10605);
or U11827 (N_11827,N_10984,N_10715);
nor U11828 (N_11828,N_10341,N_10082);
nor U11829 (N_11829,N_10455,N_10973);
nand U11830 (N_11830,N_10491,N_10019);
xnor U11831 (N_11831,N_10169,N_10912);
or U11832 (N_11832,N_10688,N_10427);
and U11833 (N_11833,N_10644,N_10208);
or U11834 (N_11834,N_10460,N_10939);
nand U11835 (N_11835,N_10936,N_10733);
and U11836 (N_11836,N_10436,N_10296);
nand U11837 (N_11837,N_10106,N_10168);
nand U11838 (N_11838,N_10191,N_10600);
nand U11839 (N_11839,N_10558,N_10981);
or U11840 (N_11840,N_10166,N_10608);
or U11841 (N_11841,N_10377,N_10418);
xor U11842 (N_11842,N_10963,N_10693);
nand U11843 (N_11843,N_10376,N_10231);
and U11844 (N_11844,N_10349,N_10967);
and U11845 (N_11845,N_10392,N_10775);
and U11846 (N_11846,N_10228,N_10801);
or U11847 (N_11847,N_10978,N_10103);
xnor U11848 (N_11848,N_10489,N_10068);
nor U11849 (N_11849,N_10769,N_10212);
xor U11850 (N_11850,N_10935,N_10462);
or U11851 (N_11851,N_10285,N_10231);
nand U11852 (N_11852,N_10867,N_10066);
and U11853 (N_11853,N_10783,N_10330);
xor U11854 (N_11854,N_10144,N_10763);
and U11855 (N_11855,N_10117,N_10593);
or U11856 (N_11856,N_10072,N_10932);
nor U11857 (N_11857,N_10700,N_10830);
nor U11858 (N_11858,N_10892,N_10081);
nand U11859 (N_11859,N_10233,N_10501);
nand U11860 (N_11860,N_10335,N_10524);
or U11861 (N_11861,N_10579,N_10063);
xnor U11862 (N_11862,N_10362,N_10132);
nor U11863 (N_11863,N_10895,N_10492);
xnor U11864 (N_11864,N_10733,N_10928);
nand U11865 (N_11865,N_10543,N_10101);
and U11866 (N_11866,N_10315,N_10947);
nand U11867 (N_11867,N_10583,N_10598);
nor U11868 (N_11868,N_10192,N_10368);
nor U11869 (N_11869,N_10706,N_10854);
and U11870 (N_11870,N_10185,N_10058);
and U11871 (N_11871,N_10302,N_10752);
and U11872 (N_11872,N_10065,N_10623);
xnor U11873 (N_11873,N_10304,N_10471);
nand U11874 (N_11874,N_10786,N_10723);
nand U11875 (N_11875,N_10179,N_10686);
and U11876 (N_11876,N_10060,N_10786);
nand U11877 (N_11877,N_10619,N_10161);
or U11878 (N_11878,N_10014,N_10514);
xor U11879 (N_11879,N_10380,N_10578);
nor U11880 (N_11880,N_10496,N_10781);
nand U11881 (N_11881,N_10799,N_10199);
and U11882 (N_11882,N_10280,N_10540);
xnor U11883 (N_11883,N_10255,N_10404);
xor U11884 (N_11884,N_10706,N_10352);
xnor U11885 (N_11885,N_10956,N_10475);
and U11886 (N_11886,N_10224,N_10531);
nand U11887 (N_11887,N_10460,N_10201);
and U11888 (N_11888,N_10481,N_10292);
nand U11889 (N_11889,N_10977,N_10628);
and U11890 (N_11890,N_10671,N_10593);
nor U11891 (N_11891,N_10067,N_10788);
or U11892 (N_11892,N_10763,N_10745);
or U11893 (N_11893,N_10471,N_10466);
and U11894 (N_11894,N_10260,N_10674);
nor U11895 (N_11895,N_10773,N_10871);
xnor U11896 (N_11896,N_10410,N_10964);
xnor U11897 (N_11897,N_10588,N_10373);
or U11898 (N_11898,N_10256,N_10721);
xnor U11899 (N_11899,N_10373,N_10102);
or U11900 (N_11900,N_10249,N_10574);
nor U11901 (N_11901,N_10933,N_10095);
nand U11902 (N_11902,N_10702,N_10609);
xor U11903 (N_11903,N_10800,N_10036);
nor U11904 (N_11904,N_10645,N_10209);
or U11905 (N_11905,N_10220,N_10669);
and U11906 (N_11906,N_10724,N_10500);
nor U11907 (N_11907,N_10424,N_10183);
or U11908 (N_11908,N_10501,N_10925);
or U11909 (N_11909,N_10679,N_10060);
and U11910 (N_11910,N_10693,N_10589);
or U11911 (N_11911,N_10455,N_10865);
or U11912 (N_11912,N_10223,N_10080);
and U11913 (N_11913,N_10933,N_10652);
nor U11914 (N_11914,N_10204,N_10117);
or U11915 (N_11915,N_10789,N_10622);
xor U11916 (N_11916,N_10296,N_10447);
xnor U11917 (N_11917,N_10142,N_10330);
or U11918 (N_11918,N_10655,N_10081);
or U11919 (N_11919,N_10837,N_10170);
or U11920 (N_11920,N_10866,N_10704);
xor U11921 (N_11921,N_10809,N_10759);
nor U11922 (N_11922,N_10988,N_10104);
nand U11923 (N_11923,N_10038,N_10419);
nand U11924 (N_11924,N_10913,N_10742);
xor U11925 (N_11925,N_10544,N_10405);
xor U11926 (N_11926,N_10130,N_10529);
or U11927 (N_11927,N_10643,N_10273);
xor U11928 (N_11928,N_10671,N_10403);
nand U11929 (N_11929,N_10863,N_10576);
xor U11930 (N_11930,N_10124,N_10110);
xor U11931 (N_11931,N_10791,N_10941);
and U11932 (N_11932,N_10913,N_10756);
or U11933 (N_11933,N_10811,N_10544);
and U11934 (N_11934,N_10828,N_10407);
xor U11935 (N_11935,N_10768,N_10113);
nand U11936 (N_11936,N_10504,N_10425);
and U11937 (N_11937,N_10810,N_10130);
and U11938 (N_11938,N_10852,N_10724);
or U11939 (N_11939,N_10441,N_10179);
and U11940 (N_11940,N_10418,N_10822);
nand U11941 (N_11941,N_10307,N_10412);
or U11942 (N_11942,N_10194,N_10181);
and U11943 (N_11943,N_10682,N_10075);
xnor U11944 (N_11944,N_10610,N_10781);
nor U11945 (N_11945,N_10349,N_10773);
or U11946 (N_11946,N_10349,N_10166);
nand U11947 (N_11947,N_10974,N_10607);
xnor U11948 (N_11948,N_10602,N_10978);
and U11949 (N_11949,N_10439,N_10052);
nor U11950 (N_11950,N_10133,N_10278);
and U11951 (N_11951,N_10725,N_10873);
nand U11952 (N_11952,N_10137,N_10237);
and U11953 (N_11953,N_10217,N_10576);
and U11954 (N_11954,N_10341,N_10709);
xnor U11955 (N_11955,N_10097,N_10023);
nor U11956 (N_11956,N_10917,N_10519);
nor U11957 (N_11957,N_10594,N_10115);
nor U11958 (N_11958,N_10167,N_10875);
and U11959 (N_11959,N_10064,N_10230);
or U11960 (N_11960,N_10865,N_10321);
and U11961 (N_11961,N_10677,N_10082);
nor U11962 (N_11962,N_10836,N_10077);
xor U11963 (N_11963,N_10095,N_10888);
xor U11964 (N_11964,N_10872,N_10096);
nor U11965 (N_11965,N_10271,N_10004);
xnor U11966 (N_11966,N_10575,N_10414);
nor U11967 (N_11967,N_10791,N_10414);
or U11968 (N_11968,N_10675,N_10087);
or U11969 (N_11969,N_10128,N_10826);
nor U11970 (N_11970,N_10055,N_10631);
nor U11971 (N_11971,N_10413,N_10216);
nor U11972 (N_11972,N_10389,N_10100);
xnor U11973 (N_11973,N_10278,N_10455);
nor U11974 (N_11974,N_10016,N_10313);
nand U11975 (N_11975,N_10777,N_10140);
nor U11976 (N_11976,N_10998,N_10892);
and U11977 (N_11977,N_10851,N_10771);
nor U11978 (N_11978,N_10381,N_10368);
and U11979 (N_11979,N_10207,N_10499);
nor U11980 (N_11980,N_10487,N_10136);
or U11981 (N_11981,N_10577,N_10046);
or U11982 (N_11982,N_10497,N_10133);
nor U11983 (N_11983,N_10746,N_10779);
or U11984 (N_11984,N_10009,N_10711);
nand U11985 (N_11985,N_10836,N_10745);
nand U11986 (N_11986,N_10674,N_10121);
or U11987 (N_11987,N_10992,N_10894);
and U11988 (N_11988,N_10911,N_10210);
xnor U11989 (N_11989,N_10555,N_10178);
nor U11990 (N_11990,N_10951,N_10482);
or U11991 (N_11991,N_10217,N_10799);
nor U11992 (N_11992,N_10856,N_10609);
or U11993 (N_11993,N_10884,N_10000);
nand U11994 (N_11994,N_10858,N_10674);
nand U11995 (N_11995,N_10877,N_10058);
nand U11996 (N_11996,N_10332,N_10982);
nor U11997 (N_11997,N_10051,N_10496);
and U11998 (N_11998,N_10558,N_10948);
or U11999 (N_11999,N_10263,N_10697);
nor U12000 (N_12000,N_11384,N_11478);
xnor U12001 (N_12001,N_11794,N_11744);
and U12002 (N_12002,N_11515,N_11319);
xnor U12003 (N_12003,N_11006,N_11029);
xor U12004 (N_12004,N_11623,N_11456);
xor U12005 (N_12005,N_11322,N_11308);
xnor U12006 (N_12006,N_11187,N_11805);
xor U12007 (N_12007,N_11171,N_11775);
or U12008 (N_12008,N_11757,N_11525);
xnor U12009 (N_12009,N_11050,N_11530);
nor U12010 (N_12010,N_11682,N_11060);
and U12011 (N_12011,N_11130,N_11237);
and U12012 (N_12012,N_11025,N_11020);
nand U12013 (N_12013,N_11164,N_11353);
or U12014 (N_12014,N_11637,N_11523);
and U12015 (N_12015,N_11486,N_11166);
or U12016 (N_12016,N_11061,N_11449);
xor U12017 (N_12017,N_11192,N_11728);
xnor U12018 (N_12018,N_11548,N_11428);
or U12019 (N_12019,N_11616,N_11337);
nor U12020 (N_12020,N_11552,N_11712);
xor U12021 (N_12021,N_11748,N_11786);
or U12022 (N_12022,N_11475,N_11640);
nor U12023 (N_12023,N_11247,N_11904);
xor U12024 (N_12024,N_11188,N_11070);
nor U12025 (N_12025,N_11159,N_11819);
or U12026 (N_12026,N_11887,N_11612);
or U12027 (N_12027,N_11069,N_11348);
or U12028 (N_12028,N_11088,N_11709);
or U12029 (N_12029,N_11971,N_11807);
xor U12030 (N_12030,N_11176,N_11831);
nor U12031 (N_12031,N_11420,N_11660);
or U12032 (N_12032,N_11442,N_11719);
nand U12033 (N_12033,N_11964,N_11080);
xnor U12034 (N_12034,N_11511,N_11751);
nor U12035 (N_12035,N_11778,N_11367);
and U12036 (N_12036,N_11139,N_11376);
nor U12037 (N_12037,N_11415,N_11095);
or U12038 (N_12038,N_11865,N_11032);
nor U12039 (N_12039,N_11386,N_11163);
nor U12040 (N_12040,N_11126,N_11555);
and U12041 (N_12041,N_11395,N_11848);
and U12042 (N_12042,N_11871,N_11365);
nor U12043 (N_12043,N_11368,N_11856);
xor U12044 (N_12044,N_11675,N_11059);
nand U12045 (N_12045,N_11306,N_11950);
and U12046 (N_12046,N_11972,N_11470);
nor U12047 (N_12047,N_11736,N_11764);
nor U12048 (N_12048,N_11068,N_11575);
nor U12049 (N_12049,N_11944,N_11214);
xnor U12050 (N_12050,N_11746,N_11557);
and U12051 (N_12051,N_11499,N_11699);
xnor U12052 (N_12052,N_11947,N_11364);
nor U12053 (N_12053,N_11978,N_11646);
and U12054 (N_12054,N_11577,N_11324);
or U12055 (N_12055,N_11143,N_11042);
nor U12056 (N_12056,N_11418,N_11158);
nand U12057 (N_12057,N_11927,N_11627);
xnor U12058 (N_12058,N_11878,N_11148);
and U12059 (N_12059,N_11402,N_11284);
xor U12060 (N_12060,N_11033,N_11326);
or U12061 (N_12061,N_11867,N_11618);
xor U12062 (N_12062,N_11081,N_11624);
nor U12063 (N_12063,N_11544,N_11250);
nand U12064 (N_12064,N_11372,N_11474);
nor U12065 (N_12065,N_11593,N_11174);
nor U12066 (N_12066,N_11168,N_11708);
nand U12067 (N_12067,N_11318,N_11452);
or U12068 (N_12068,N_11361,N_11213);
nand U12069 (N_12069,N_11467,N_11241);
xnor U12070 (N_12070,N_11272,N_11731);
nand U12071 (N_12071,N_11431,N_11203);
nand U12072 (N_12072,N_11404,N_11524);
xor U12073 (N_12073,N_11201,N_11795);
xor U12074 (N_12074,N_11890,N_11275);
or U12075 (N_12075,N_11399,N_11255);
nor U12076 (N_12076,N_11980,N_11836);
nor U12077 (N_12077,N_11363,N_11790);
and U12078 (N_12078,N_11263,N_11849);
nand U12079 (N_12079,N_11044,N_11129);
nand U12080 (N_12080,N_11521,N_11082);
or U12081 (N_12081,N_11816,N_11468);
nand U12082 (N_12082,N_11864,N_11335);
and U12083 (N_12083,N_11641,N_11939);
and U12084 (N_12084,N_11462,N_11313);
nor U12085 (N_12085,N_11099,N_11868);
or U12086 (N_12086,N_11052,N_11953);
and U12087 (N_12087,N_11409,N_11833);
nand U12088 (N_12088,N_11289,N_11608);
or U12089 (N_12089,N_11986,N_11750);
nor U12090 (N_12090,N_11687,N_11110);
xor U12091 (N_12091,N_11488,N_11962);
or U12092 (N_12092,N_11128,N_11948);
or U12093 (N_12093,N_11569,N_11253);
nand U12094 (N_12094,N_11051,N_11926);
xnor U12095 (N_12095,N_11038,N_11869);
and U12096 (N_12096,N_11131,N_11889);
nand U12097 (N_12097,N_11850,N_11259);
xor U12098 (N_12098,N_11056,N_11842);
xor U12099 (N_12099,N_11261,N_11861);
xnor U12100 (N_12100,N_11560,N_11279);
nand U12101 (N_12101,N_11196,N_11875);
or U12102 (N_12102,N_11483,N_11940);
nor U12103 (N_12103,N_11340,N_11600);
or U12104 (N_12104,N_11329,N_11508);
xnor U12105 (N_12105,N_11305,N_11469);
and U12106 (N_12106,N_11223,N_11678);
or U12107 (N_12107,N_11346,N_11460);
or U12108 (N_12108,N_11244,N_11934);
nor U12109 (N_12109,N_11249,N_11763);
xnor U12110 (N_12110,N_11929,N_11700);
nand U12111 (N_12111,N_11437,N_11681);
nand U12112 (N_12112,N_11233,N_11632);
nor U12113 (N_12113,N_11723,N_11743);
xor U12114 (N_12114,N_11388,N_11382);
xnor U12115 (N_12115,N_11767,N_11136);
nand U12116 (N_12116,N_11598,N_11717);
nand U12117 (N_12117,N_11662,N_11771);
or U12118 (N_12118,N_11278,N_11380);
or U12119 (N_12119,N_11208,N_11121);
and U12120 (N_12120,N_11776,N_11107);
and U12121 (N_12121,N_11015,N_11998);
nor U12122 (N_12122,N_11605,N_11315);
nand U12123 (N_12123,N_11299,N_11977);
xor U12124 (N_12124,N_11023,N_11286);
or U12125 (N_12125,N_11602,N_11410);
xnor U12126 (N_12126,N_11374,N_11839);
nand U12127 (N_12127,N_11103,N_11979);
nand U12128 (N_12128,N_11574,N_11144);
or U12129 (N_12129,N_11898,N_11425);
xor U12130 (N_12130,N_11584,N_11447);
nand U12131 (N_12131,N_11390,N_11693);
or U12132 (N_12132,N_11484,N_11886);
nand U12133 (N_12133,N_11993,N_11269);
nor U12134 (N_12134,N_11942,N_11943);
nor U12135 (N_12135,N_11297,N_11028);
nor U12136 (N_12136,N_11761,N_11609);
or U12137 (N_12137,N_11827,N_11561);
and U12138 (N_12138,N_11595,N_11918);
xor U12139 (N_12139,N_11938,N_11156);
nor U12140 (N_12140,N_11446,N_11601);
nor U12141 (N_12141,N_11243,N_11277);
nor U12142 (N_12142,N_11046,N_11747);
nand U12143 (N_12143,N_11245,N_11925);
or U12144 (N_12144,N_11722,N_11303);
or U12145 (N_12145,N_11455,N_11800);
xnor U12146 (N_12146,N_11445,N_11405);
and U12147 (N_12147,N_11782,N_11298);
or U12148 (N_12148,N_11408,N_11969);
xor U12149 (N_12149,N_11599,N_11064);
nand U12150 (N_12150,N_11016,N_11300);
xnor U12151 (N_12151,N_11293,N_11003);
xor U12152 (N_12152,N_11539,N_11434);
or U12153 (N_12153,N_11184,N_11222);
xor U12154 (N_12154,N_11282,N_11251);
xor U12155 (N_12155,N_11650,N_11888);
and U12156 (N_12156,N_11783,N_11177);
xor U12157 (N_12157,N_11529,N_11606);
nor U12158 (N_12158,N_11098,N_11360);
xnor U12159 (N_12159,N_11497,N_11076);
or U12160 (N_12160,N_11866,N_11369);
nor U12161 (N_12161,N_11073,N_11851);
nand U12162 (N_12162,N_11494,N_11914);
or U12163 (N_12163,N_11565,N_11965);
and U12164 (N_12164,N_11151,N_11847);
xnor U12165 (N_12165,N_11840,N_11145);
and U12166 (N_12166,N_11031,N_11493);
and U12167 (N_12167,N_11085,N_11652);
nand U12168 (N_12168,N_11506,N_11354);
nand U12169 (N_12169,N_11997,N_11371);
nand U12170 (N_12170,N_11160,N_11667);
xnor U12171 (N_12171,N_11570,N_11949);
or U12172 (N_12172,N_11491,N_11695);
and U12173 (N_12173,N_11824,N_11172);
and U12174 (N_12174,N_11457,N_11412);
or U12175 (N_12175,N_11629,N_11119);
and U12176 (N_12176,N_11818,N_11647);
nand U12177 (N_12177,N_11215,N_11919);
or U12178 (N_12178,N_11067,N_11973);
nor U12179 (N_12179,N_11772,N_11901);
nand U12180 (N_12180,N_11239,N_11635);
xor U12181 (N_12181,N_11473,N_11175);
nor U12182 (N_12182,N_11820,N_11932);
or U12183 (N_12183,N_11443,N_11806);
xnor U12184 (N_12184,N_11075,N_11127);
xor U12185 (N_12185,N_11909,N_11009);
or U12186 (N_12186,N_11150,N_11673);
xnor U12187 (N_12187,N_11799,N_11663);
xnor U12188 (N_12188,N_11122,N_11435);
xnor U12189 (N_12189,N_11454,N_11910);
xor U12190 (N_12190,N_11536,N_11458);
xnor U12191 (N_12191,N_11894,N_11347);
nand U12192 (N_12192,N_11302,N_11310);
or U12193 (N_12193,N_11375,N_11974);
nand U12194 (N_12194,N_11661,N_11716);
nand U12195 (N_12195,N_11876,N_11373);
xor U12196 (N_12196,N_11622,N_11210);
nand U12197 (N_12197,N_11516,N_11242);
or U12198 (N_12198,N_11787,N_11017);
and U12199 (N_12199,N_11492,N_11113);
xnor U12200 (N_12200,N_11729,N_11796);
xor U12201 (N_12201,N_11216,N_11720);
nor U12202 (N_12202,N_11568,N_11562);
xor U12203 (N_12203,N_11835,N_11656);
and U12204 (N_12204,N_11742,N_11180);
and U12205 (N_12205,N_11558,N_11264);
xnor U12206 (N_12206,N_11047,N_11007);
or U12207 (N_12207,N_11262,N_11958);
xor U12208 (N_12208,N_11270,N_11877);
or U12209 (N_12209,N_11636,N_11520);
nor U12210 (N_12210,N_11753,N_11906);
nand U12211 (N_12211,N_11960,N_11022);
or U12212 (N_12212,N_11970,N_11741);
nand U12213 (N_12213,N_11923,N_11413);
and U12214 (N_12214,N_11967,N_11692);
or U12215 (N_12215,N_11838,N_11749);
or U12216 (N_12216,N_11086,N_11765);
xor U12217 (N_12217,N_11035,N_11117);
and U12218 (N_12218,N_11549,N_11430);
nor U12219 (N_12219,N_11698,N_11792);
nand U12220 (N_12220,N_11785,N_11981);
nand U12221 (N_12221,N_11448,N_11394);
and U12222 (N_12222,N_11968,N_11352);
and U12223 (N_12223,N_11533,N_11634);
and U12224 (N_12224,N_11345,N_11218);
xnor U12225 (N_12225,N_11651,N_11436);
and U12226 (N_12226,N_11014,N_11167);
and U12227 (N_12227,N_11162,N_11359);
and U12228 (N_12228,N_11951,N_11846);
xnor U12229 (N_12229,N_11908,N_11758);
nand U12230 (N_12230,N_11519,N_11774);
nor U12231 (N_12231,N_11671,N_11205);
or U12232 (N_12232,N_11730,N_11476);
and U12233 (N_12233,N_11542,N_11190);
nand U12234 (N_12234,N_11803,N_11226);
nand U12235 (N_12235,N_11200,N_11316);
xor U12236 (N_12236,N_11391,N_11759);
or U12237 (N_12237,N_11071,N_11400);
and U12238 (N_12238,N_11439,N_11578);
or U12239 (N_12239,N_11267,N_11477);
nor U12240 (N_12240,N_11004,N_11451);
xor U12241 (N_12241,N_11461,N_11355);
nor U12242 (N_12242,N_11726,N_11490);
xnor U12243 (N_12243,N_11897,N_11781);
nor U12244 (N_12244,N_11387,N_11857);
or U12245 (N_12245,N_11639,N_11132);
or U12246 (N_12246,N_11224,N_11703);
nand U12247 (N_12247,N_11021,N_11685);
nand U12248 (N_12248,N_11586,N_11591);
and U12249 (N_12249,N_11826,N_11766);
xor U12250 (N_12250,N_11920,N_11106);
and U12251 (N_12251,N_11679,N_11809);
nor U12252 (N_12252,N_11621,N_11713);
and U12253 (N_12253,N_11238,N_11854);
xnor U12254 (N_12254,N_11714,N_11696);
nor U12255 (N_12255,N_11266,N_11913);
and U12256 (N_12256,N_11414,N_11545);
nand U12257 (N_12257,N_11024,N_11845);
nand U12258 (N_12258,N_11810,N_11221);
nor U12259 (N_12259,N_11027,N_11874);
xnor U12260 (N_12260,N_11690,N_11582);
nand U12261 (N_12261,N_11770,N_11522);
nor U12262 (N_12262,N_11327,N_11105);
or U12263 (N_12263,N_11668,N_11401);
or U12264 (N_12264,N_11994,N_11509);
xor U12265 (N_12265,N_11202,N_11538);
or U12266 (N_12266,N_11514,N_11546);
xnor U12267 (N_12267,N_11916,N_11220);
or U12268 (N_12268,N_11320,N_11392);
and U12269 (N_12269,N_11396,N_11333);
and U12270 (N_12270,N_11377,N_11737);
nor U12271 (N_12271,N_11350,N_11768);
xor U12272 (N_12272,N_11655,N_11195);
xnor U12273 (N_12273,N_11183,N_11053);
and U12274 (N_12274,N_11732,N_11231);
and U12275 (N_12275,N_11645,N_11048);
xor U12276 (N_12276,N_11141,N_11610);
xnor U12277 (N_12277,N_11983,N_11881);
nand U12278 (N_12278,N_11248,N_11344);
xor U12279 (N_12279,N_11513,N_11198);
or U12280 (N_12280,N_11534,N_11686);
and U12281 (N_12281,N_11094,N_11579);
or U12282 (N_12282,N_11411,N_11169);
or U12283 (N_12283,N_11225,N_11922);
nand U12284 (N_12284,N_11419,N_11961);
xnor U12285 (N_12285,N_11417,N_11466);
and U12286 (N_12286,N_11273,N_11501);
and U12287 (N_12287,N_11294,N_11532);
xor U12288 (N_12288,N_11587,N_11931);
nor U12289 (N_12289,N_11657,N_11459);
and U12290 (N_12290,N_11531,N_11311);
xor U12291 (N_12291,N_11915,N_11946);
and U12292 (N_12292,N_11055,N_11444);
xnor U12293 (N_12293,N_11423,N_11788);
xor U12294 (N_12294,N_11090,N_11398);
xor U12295 (N_12295,N_11096,N_11342);
nand U12296 (N_12296,N_11312,N_11065);
xnor U12297 (N_12297,N_11832,N_11339);
and U12298 (N_12298,N_11093,N_11626);
xnor U12299 (N_12299,N_11011,N_11590);
or U12300 (N_12300,N_11290,N_11072);
nand U12301 (N_12301,N_11860,N_11450);
nand U12302 (N_12302,N_11999,N_11734);
or U12303 (N_12303,N_11821,N_11844);
or U12304 (N_12304,N_11049,N_11706);
nor U12305 (N_12305,N_11937,N_11037);
and U12306 (N_12306,N_11254,N_11236);
nor U12307 (N_12307,N_11291,N_11882);
and U12308 (N_12308,N_11019,N_11873);
and U12309 (N_12309,N_11589,N_11870);
xnor U12310 (N_12310,N_11186,N_11995);
nand U12311 (N_12311,N_11625,N_11982);
nand U12312 (N_12312,N_11791,N_11379);
nor U12313 (N_12313,N_11825,N_11204);
xor U12314 (N_12314,N_11041,N_11550);
nor U12315 (N_12315,N_11537,N_11100);
nand U12316 (N_12316,N_11683,N_11553);
nand U12317 (N_12317,N_11274,N_11672);
and U12318 (N_12318,N_11872,N_11331);
nor U12319 (N_12319,N_11966,N_11615);
xnor U12320 (N_12320,N_11991,N_11941);
nand U12321 (N_12321,N_11863,N_11830);
and U12322 (N_12322,N_11109,N_11822);
or U12323 (N_12323,N_11510,N_11936);
nand U12324 (N_12324,N_11573,N_11314);
or U12325 (N_12325,N_11370,N_11433);
nor U12326 (N_12326,N_11138,N_11271);
nor U12327 (N_12327,N_11594,N_11912);
and U12328 (N_12328,N_11114,N_11724);
and U12329 (N_12329,N_11665,N_11118);
or U12330 (N_12330,N_11045,N_11489);
nand U12331 (N_12331,N_11855,N_11030);
xnor U12332 (N_12332,N_11815,N_11309);
xor U12333 (N_12333,N_11843,N_11620);
nand U12334 (N_12334,N_11691,N_11793);
xnor U12335 (N_12335,N_11209,N_11924);
or U12336 (N_12336,N_11780,N_11258);
xor U12337 (N_12337,N_11407,N_11659);
xnor U12338 (N_12338,N_11811,N_11762);
nor U12339 (N_12339,N_11240,N_11108);
nand U12340 (N_12340,N_11232,N_11643);
xnor U12341 (N_12341,N_11984,N_11323);
nor U12342 (N_12342,N_11554,N_11194);
or U12343 (N_12343,N_11252,N_11089);
xor U12344 (N_12344,N_11633,N_11985);
nand U12345 (N_12345,N_11517,N_11893);
and U12346 (N_12346,N_11954,N_11104);
or U12347 (N_12347,N_11234,N_11694);
nand U12348 (N_12348,N_11596,N_11173);
or U12349 (N_12349,N_11518,N_11644);
xnor U12350 (N_12350,N_11178,N_11638);
xor U12351 (N_12351,N_11140,N_11432);
or U12352 (N_12352,N_11721,N_11823);
or U12353 (N_12353,N_11120,N_11260);
or U12354 (N_12354,N_11101,N_11197);
nor U12355 (N_12355,N_11504,N_11841);
nand U12356 (N_12356,N_11181,N_11976);
or U12357 (N_12357,N_11341,N_11066);
nand U12358 (N_12358,N_11862,N_11317);
nor U12359 (N_12359,N_11642,N_11078);
nand U12360 (N_12360,N_11684,N_11834);
xor U12361 (N_12361,N_11325,N_11349);
or U12362 (N_12362,N_11357,N_11817);
xor U12363 (N_12363,N_11670,N_11858);
nor U12364 (N_12364,N_11779,N_11097);
nor U12365 (N_12365,N_11149,N_11769);
or U12366 (N_12366,N_11566,N_11191);
or U12367 (N_12367,N_11057,N_11812);
and U12368 (N_12368,N_11091,N_11828);
nor U12369 (N_12369,N_11988,N_11124);
xnor U12370 (N_12370,N_11406,N_11281);
or U12371 (N_12371,N_11301,N_11631);
nand U12372 (N_12372,N_11334,N_11733);
or U12373 (N_12373,N_11421,N_11512);
nand U12374 (N_12374,N_11987,N_11885);
nor U12375 (N_12375,N_11572,N_11356);
nor U12376 (N_12376,N_11351,N_11649);
xor U12377 (N_12377,N_11911,N_11480);
xnor U12378 (N_12378,N_11182,N_11959);
and U12379 (N_12379,N_11125,N_11735);
xnor U12380 (N_12380,N_11040,N_11664);
and U12381 (N_12381,N_11592,N_11654);
nand U12382 (N_12382,N_11453,N_11393);
nor U12383 (N_12383,N_11503,N_11283);
and U12384 (N_12384,N_11705,N_11362);
xor U12385 (N_12385,N_11482,N_11597);
and U12386 (N_12386,N_11837,N_11427);
xor U12387 (N_12387,N_11185,N_11471);
or U12388 (N_12388,N_11465,N_11666);
or U12389 (N_12389,N_11674,N_11111);
nand U12390 (N_12390,N_11199,N_11507);
nand U12391 (N_12391,N_11378,N_11495);
nand U12392 (N_12392,N_11102,N_11063);
or U12393 (N_12393,N_11852,N_11963);
and U12394 (N_12394,N_11535,N_11797);
nor U12395 (N_12395,N_11385,N_11039);
xnor U12396 (N_12396,N_11296,N_11715);
nand U12397 (N_12397,N_11358,N_11676);
xor U12398 (N_12398,N_11527,N_11256);
nand U12399 (N_12399,N_11727,N_11784);
or U12400 (N_12400,N_11739,N_11292);
nand U12401 (N_12401,N_11990,N_11902);
or U12402 (N_12402,N_11268,N_11952);
nor U12403 (N_12403,N_11212,N_11740);
and U12404 (N_12404,N_11808,N_11134);
nand U12405 (N_12405,N_11933,N_11155);
or U12406 (N_12406,N_11630,N_11229);
xnor U12407 (N_12407,N_11583,N_11043);
nand U12408 (N_12408,N_11907,N_11669);
or U12409 (N_12409,N_11752,N_11115);
nor U12410 (N_12410,N_11528,N_11896);
nor U12411 (N_12411,N_11010,N_11680);
xor U12412 (N_12412,N_11227,N_11760);
nor U12413 (N_12413,N_11087,N_11219);
or U12414 (N_12414,N_11658,N_11502);
and U12415 (N_12415,N_11276,N_11677);
nor U12416 (N_12416,N_11718,N_11648);
xnor U12417 (N_12417,N_11883,N_11905);
nand U12418 (N_12418,N_11193,N_11814);
nor U12419 (N_12419,N_11170,N_11604);
nor U12420 (N_12420,N_11957,N_11416);
xnor U12421 (N_12421,N_11332,N_11580);
nor U12422 (N_12422,N_11899,N_11738);
nor U12423 (N_12423,N_11154,N_11802);
or U12424 (N_12424,N_11804,N_11133);
and U12425 (N_12425,N_11389,N_11496);
or U12426 (N_12426,N_11903,N_11829);
xor U12427 (N_12427,N_11207,N_11152);
or U12428 (N_12428,N_11567,N_11628);
and U12429 (N_12429,N_11813,N_11479);
and U12430 (N_12430,N_11230,N_11321);
or U12431 (N_12431,N_11077,N_11383);
nand U12432 (N_12432,N_11745,N_11343);
and U12433 (N_12433,N_11304,N_11054);
and U12434 (N_12434,N_11137,N_11702);
xor U12435 (N_12435,N_11556,N_11008);
or U12436 (N_12436,N_11955,N_11366);
xnor U12437 (N_12437,N_11996,N_11074);
nand U12438 (N_12438,N_11704,N_11551);
or U12439 (N_12439,N_11288,N_11725);
and U12440 (N_12440,N_11500,N_11058);
nor U12441 (N_12441,N_11485,N_11498);
and U12442 (N_12442,N_11062,N_11754);
or U12443 (N_12443,N_11756,N_11928);
xor U12444 (N_12444,N_11426,N_11859);
and U12445 (N_12445,N_11755,N_11189);
nor U12446 (N_12446,N_11710,N_11607);
or U12447 (N_12447,N_11992,N_11801);
nor U12448 (N_12448,N_11547,N_11989);
nand U12449 (N_12449,N_11034,N_11935);
nand U12450 (N_12450,N_11559,N_11526);
nor U12451 (N_12451,N_11285,N_11880);
xnor U12452 (N_12452,N_11930,N_11257);
or U12453 (N_12453,N_11879,N_11328);
or U12454 (N_12454,N_11472,N_11921);
nor U12455 (N_12455,N_11381,N_11481);
or U12456 (N_12456,N_11228,N_11707);
or U12457 (N_12457,N_11287,N_11330);
nor U12458 (N_12458,N_11689,N_11161);
nand U12459 (N_12459,N_11614,N_11112);
or U12460 (N_12460,N_11956,N_11917);
xor U12461 (N_12461,N_11798,N_11135);
nor U12462 (N_12462,N_11585,N_11146);
and U12463 (N_12463,N_11853,N_11588);
and U12464 (N_12464,N_11895,N_11711);
and U12465 (N_12465,N_11116,N_11777);
and U12466 (N_12466,N_11945,N_11611);
xor U12467 (N_12467,N_11211,N_11789);
and U12468 (N_12468,N_11026,N_11697);
nor U12469 (N_12469,N_11541,N_11688);
nor U12470 (N_12470,N_11084,N_11295);
nor U12471 (N_12471,N_11000,N_11179);
nor U12472 (N_12472,N_11036,N_11892);
xnor U12473 (N_12473,N_11013,N_11092);
nor U12474 (N_12474,N_11336,N_11338);
or U12475 (N_12475,N_11123,N_11773);
nor U12476 (N_12476,N_11884,N_11619);
or U12477 (N_12477,N_11002,N_11564);
xor U12478 (N_12478,N_11206,N_11012);
nor U12479 (N_12479,N_11018,N_11975);
or U12480 (N_12480,N_11280,N_11563);
nand U12481 (N_12481,N_11307,N_11083);
nand U12482 (N_12482,N_11005,N_11246);
xnor U12483 (N_12483,N_11571,N_11438);
xor U12484 (N_12484,N_11653,N_11543);
nor U12485 (N_12485,N_11464,N_11617);
nor U12486 (N_12486,N_11165,N_11147);
nand U12487 (N_12487,N_11900,N_11463);
xor U12488 (N_12488,N_11603,N_11441);
xnor U12489 (N_12489,N_11422,N_11891);
nand U12490 (N_12490,N_11265,N_11429);
nand U12491 (N_12491,N_11157,N_11505);
nand U12492 (N_12492,N_11576,N_11403);
nand U12493 (N_12493,N_11581,N_11701);
xor U12494 (N_12494,N_11487,N_11540);
nor U12495 (N_12495,N_11235,N_11079);
nand U12496 (N_12496,N_11440,N_11424);
nor U12497 (N_12497,N_11217,N_11153);
and U12498 (N_12498,N_11613,N_11001);
nand U12499 (N_12499,N_11397,N_11142);
xnor U12500 (N_12500,N_11369,N_11719);
nor U12501 (N_12501,N_11484,N_11547);
and U12502 (N_12502,N_11814,N_11848);
nor U12503 (N_12503,N_11431,N_11384);
xnor U12504 (N_12504,N_11584,N_11153);
xor U12505 (N_12505,N_11083,N_11971);
xnor U12506 (N_12506,N_11115,N_11432);
nor U12507 (N_12507,N_11920,N_11581);
and U12508 (N_12508,N_11529,N_11458);
xor U12509 (N_12509,N_11491,N_11176);
nor U12510 (N_12510,N_11751,N_11868);
nor U12511 (N_12511,N_11084,N_11165);
or U12512 (N_12512,N_11040,N_11284);
nor U12513 (N_12513,N_11935,N_11845);
nor U12514 (N_12514,N_11600,N_11707);
and U12515 (N_12515,N_11269,N_11110);
xor U12516 (N_12516,N_11985,N_11416);
nand U12517 (N_12517,N_11384,N_11079);
or U12518 (N_12518,N_11731,N_11208);
xor U12519 (N_12519,N_11451,N_11491);
and U12520 (N_12520,N_11145,N_11499);
nor U12521 (N_12521,N_11078,N_11652);
nor U12522 (N_12522,N_11350,N_11860);
nand U12523 (N_12523,N_11080,N_11336);
or U12524 (N_12524,N_11750,N_11829);
or U12525 (N_12525,N_11587,N_11046);
xor U12526 (N_12526,N_11429,N_11010);
nand U12527 (N_12527,N_11753,N_11048);
xor U12528 (N_12528,N_11772,N_11250);
nand U12529 (N_12529,N_11095,N_11017);
nor U12530 (N_12530,N_11135,N_11741);
xor U12531 (N_12531,N_11135,N_11054);
or U12532 (N_12532,N_11441,N_11275);
nor U12533 (N_12533,N_11486,N_11009);
xnor U12534 (N_12534,N_11672,N_11114);
or U12535 (N_12535,N_11858,N_11980);
nand U12536 (N_12536,N_11444,N_11643);
and U12537 (N_12537,N_11202,N_11910);
nor U12538 (N_12538,N_11311,N_11582);
or U12539 (N_12539,N_11026,N_11236);
nor U12540 (N_12540,N_11499,N_11824);
xor U12541 (N_12541,N_11014,N_11163);
and U12542 (N_12542,N_11321,N_11297);
and U12543 (N_12543,N_11734,N_11625);
xor U12544 (N_12544,N_11046,N_11428);
nor U12545 (N_12545,N_11884,N_11273);
or U12546 (N_12546,N_11129,N_11254);
and U12547 (N_12547,N_11706,N_11538);
xnor U12548 (N_12548,N_11887,N_11134);
nand U12549 (N_12549,N_11568,N_11563);
or U12550 (N_12550,N_11102,N_11971);
nor U12551 (N_12551,N_11483,N_11126);
and U12552 (N_12552,N_11362,N_11145);
nor U12553 (N_12553,N_11421,N_11091);
nand U12554 (N_12554,N_11727,N_11524);
and U12555 (N_12555,N_11276,N_11054);
or U12556 (N_12556,N_11577,N_11905);
nor U12557 (N_12557,N_11602,N_11708);
and U12558 (N_12558,N_11318,N_11137);
and U12559 (N_12559,N_11353,N_11497);
nand U12560 (N_12560,N_11810,N_11535);
nor U12561 (N_12561,N_11797,N_11558);
and U12562 (N_12562,N_11305,N_11285);
xnor U12563 (N_12563,N_11231,N_11841);
nand U12564 (N_12564,N_11398,N_11063);
xor U12565 (N_12565,N_11411,N_11601);
or U12566 (N_12566,N_11569,N_11818);
or U12567 (N_12567,N_11453,N_11710);
nand U12568 (N_12568,N_11326,N_11428);
nor U12569 (N_12569,N_11701,N_11490);
xor U12570 (N_12570,N_11703,N_11781);
xor U12571 (N_12571,N_11208,N_11960);
or U12572 (N_12572,N_11035,N_11008);
and U12573 (N_12573,N_11002,N_11870);
and U12574 (N_12574,N_11620,N_11953);
nor U12575 (N_12575,N_11785,N_11761);
nand U12576 (N_12576,N_11100,N_11683);
or U12577 (N_12577,N_11673,N_11033);
nand U12578 (N_12578,N_11115,N_11435);
xor U12579 (N_12579,N_11874,N_11503);
xnor U12580 (N_12580,N_11625,N_11353);
nand U12581 (N_12581,N_11264,N_11670);
xnor U12582 (N_12582,N_11976,N_11486);
and U12583 (N_12583,N_11064,N_11564);
xor U12584 (N_12584,N_11551,N_11624);
nor U12585 (N_12585,N_11356,N_11438);
xor U12586 (N_12586,N_11299,N_11554);
xnor U12587 (N_12587,N_11808,N_11009);
and U12588 (N_12588,N_11003,N_11004);
and U12589 (N_12589,N_11172,N_11154);
xnor U12590 (N_12590,N_11791,N_11765);
xor U12591 (N_12591,N_11569,N_11010);
nor U12592 (N_12592,N_11009,N_11709);
xnor U12593 (N_12593,N_11826,N_11502);
or U12594 (N_12594,N_11325,N_11084);
and U12595 (N_12595,N_11691,N_11564);
or U12596 (N_12596,N_11923,N_11447);
nor U12597 (N_12597,N_11589,N_11178);
and U12598 (N_12598,N_11127,N_11100);
nand U12599 (N_12599,N_11397,N_11484);
and U12600 (N_12600,N_11586,N_11837);
or U12601 (N_12601,N_11601,N_11804);
nor U12602 (N_12602,N_11680,N_11026);
and U12603 (N_12603,N_11810,N_11923);
or U12604 (N_12604,N_11856,N_11656);
nand U12605 (N_12605,N_11700,N_11246);
and U12606 (N_12606,N_11809,N_11068);
nor U12607 (N_12607,N_11832,N_11763);
xnor U12608 (N_12608,N_11078,N_11127);
nand U12609 (N_12609,N_11276,N_11094);
and U12610 (N_12610,N_11268,N_11493);
nor U12611 (N_12611,N_11031,N_11169);
and U12612 (N_12612,N_11729,N_11122);
nand U12613 (N_12613,N_11676,N_11722);
and U12614 (N_12614,N_11048,N_11195);
nand U12615 (N_12615,N_11270,N_11012);
xnor U12616 (N_12616,N_11734,N_11214);
or U12617 (N_12617,N_11707,N_11630);
and U12618 (N_12618,N_11038,N_11414);
and U12619 (N_12619,N_11091,N_11831);
and U12620 (N_12620,N_11338,N_11348);
nand U12621 (N_12621,N_11020,N_11223);
or U12622 (N_12622,N_11871,N_11046);
xnor U12623 (N_12623,N_11532,N_11190);
nand U12624 (N_12624,N_11837,N_11450);
or U12625 (N_12625,N_11020,N_11957);
xor U12626 (N_12626,N_11765,N_11685);
and U12627 (N_12627,N_11327,N_11810);
xnor U12628 (N_12628,N_11573,N_11198);
and U12629 (N_12629,N_11218,N_11315);
or U12630 (N_12630,N_11098,N_11426);
and U12631 (N_12631,N_11046,N_11192);
xnor U12632 (N_12632,N_11807,N_11116);
nor U12633 (N_12633,N_11325,N_11358);
nand U12634 (N_12634,N_11149,N_11789);
and U12635 (N_12635,N_11537,N_11829);
or U12636 (N_12636,N_11314,N_11007);
nand U12637 (N_12637,N_11214,N_11486);
xor U12638 (N_12638,N_11825,N_11259);
and U12639 (N_12639,N_11243,N_11298);
xnor U12640 (N_12640,N_11387,N_11176);
nand U12641 (N_12641,N_11269,N_11547);
nand U12642 (N_12642,N_11196,N_11453);
nand U12643 (N_12643,N_11799,N_11573);
and U12644 (N_12644,N_11554,N_11894);
nand U12645 (N_12645,N_11684,N_11529);
xor U12646 (N_12646,N_11102,N_11744);
nor U12647 (N_12647,N_11630,N_11967);
nand U12648 (N_12648,N_11732,N_11373);
nand U12649 (N_12649,N_11984,N_11557);
and U12650 (N_12650,N_11072,N_11990);
and U12651 (N_12651,N_11146,N_11685);
xnor U12652 (N_12652,N_11760,N_11158);
nand U12653 (N_12653,N_11499,N_11421);
or U12654 (N_12654,N_11243,N_11683);
and U12655 (N_12655,N_11463,N_11268);
and U12656 (N_12656,N_11267,N_11595);
or U12657 (N_12657,N_11202,N_11577);
xor U12658 (N_12658,N_11987,N_11312);
nor U12659 (N_12659,N_11958,N_11649);
and U12660 (N_12660,N_11902,N_11361);
and U12661 (N_12661,N_11888,N_11484);
and U12662 (N_12662,N_11790,N_11677);
nor U12663 (N_12663,N_11234,N_11751);
nor U12664 (N_12664,N_11584,N_11645);
and U12665 (N_12665,N_11192,N_11196);
nor U12666 (N_12666,N_11924,N_11918);
nor U12667 (N_12667,N_11299,N_11441);
or U12668 (N_12668,N_11179,N_11282);
xor U12669 (N_12669,N_11308,N_11996);
or U12670 (N_12670,N_11037,N_11192);
nor U12671 (N_12671,N_11264,N_11041);
nand U12672 (N_12672,N_11115,N_11364);
nor U12673 (N_12673,N_11576,N_11948);
or U12674 (N_12674,N_11734,N_11033);
nor U12675 (N_12675,N_11387,N_11328);
nand U12676 (N_12676,N_11831,N_11768);
nor U12677 (N_12677,N_11730,N_11432);
nand U12678 (N_12678,N_11187,N_11451);
nand U12679 (N_12679,N_11098,N_11053);
and U12680 (N_12680,N_11376,N_11566);
xnor U12681 (N_12681,N_11434,N_11852);
xor U12682 (N_12682,N_11898,N_11607);
and U12683 (N_12683,N_11662,N_11354);
xnor U12684 (N_12684,N_11001,N_11541);
xor U12685 (N_12685,N_11459,N_11802);
nand U12686 (N_12686,N_11346,N_11782);
xnor U12687 (N_12687,N_11987,N_11092);
and U12688 (N_12688,N_11857,N_11580);
nor U12689 (N_12689,N_11016,N_11565);
nor U12690 (N_12690,N_11414,N_11219);
and U12691 (N_12691,N_11619,N_11468);
and U12692 (N_12692,N_11009,N_11033);
nand U12693 (N_12693,N_11537,N_11826);
nand U12694 (N_12694,N_11828,N_11363);
or U12695 (N_12695,N_11375,N_11390);
nor U12696 (N_12696,N_11616,N_11088);
xnor U12697 (N_12697,N_11423,N_11741);
or U12698 (N_12698,N_11258,N_11579);
or U12699 (N_12699,N_11755,N_11708);
xor U12700 (N_12700,N_11242,N_11190);
xnor U12701 (N_12701,N_11487,N_11987);
and U12702 (N_12702,N_11957,N_11692);
nor U12703 (N_12703,N_11918,N_11711);
or U12704 (N_12704,N_11996,N_11832);
or U12705 (N_12705,N_11173,N_11540);
nand U12706 (N_12706,N_11280,N_11648);
xnor U12707 (N_12707,N_11741,N_11672);
xnor U12708 (N_12708,N_11786,N_11505);
and U12709 (N_12709,N_11702,N_11781);
and U12710 (N_12710,N_11518,N_11546);
and U12711 (N_12711,N_11533,N_11235);
xnor U12712 (N_12712,N_11120,N_11272);
nor U12713 (N_12713,N_11541,N_11602);
and U12714 (N_12714,N_11005,N_11195);
nand U12715 (N_12715,N_11922,N_11549);
xor U12716 (N_12716,N_11769,N_11274);
nand U12717 (N_12717,N_11337,N_11344);
xnor U12718 (N_12718,N_11562,N_11505);
xnor U12719 (N_12719,N_11938,N_11222);
or U12720 (N_12720,N_11562,N_11188);
xor U12721 (N_12721,N_11146,N_11035);
xnor U12722 (N_12722,N_11835,N_11869);
or U12723 (N_12723,N_11136,N_11093);
nor U12724 (N_12724,N_11818,N_11337);
or U12725 (N_12725,N_11975,N_11778);
nand U12726 (N_12726,N_11342,N_11418);
or U12727 (N_12727,N_11613,N_11493);
and U12728 (N_12728,N_11884,N_11633);
or U12729 (N_12729,N_11948,N_11686);
nand U12730 (N_12730,N_11245,N_11311);
xnor U12731 (N_12731,N_11686,N_11101);
xor U12732 (N_12732,N_11573,N_11733);
nor U12733 (N_12733,N_11641,N_11969);
xor U12734 (N_12734,N_11560,N_11146);
or U12735 (N_12735,N_11018,N_11687);
and U12736 (N_12736,N_11555,N_11179);
nand U12737 (N_12737,N_11216,N_11999);
or U12738 (N_12738,N_11628,N_11892);
and U12739 (N_12739,N_11768,N_11458);
xor U12740 (N_12740,N_11883,N_11289);
or U12741 (N_12741,N_11232,N_11300);
nor U12742 (N_12742,N_11293,N_11666);
and U12743 (N_12743,N_11619,N_11516);
xnor U12744 (N_12744,N_11875,N_11212);
nand U12745 (N_12745,N_11867,N_11403);
and U12746 (N_12746,N_11401,N_11351);
and U12747 (N_12747,N_11672,N_11828);
or U12748 (N_12748,N_11050,N_11783);
or U12749 (N_12749,N_11957,N_11778);
xor U12750 (N_12750,N_11436,N_11790);
nand U12751 (N_12751,N_11765,N_11435);
and U12752 (N_12752,N_11721,N_11480);
and U12753 (N_12753,N_11741,N_11218);
xor U12754 (N_12754,N_11183,N_11176);
or U12755 (N_12755,N_11809,N_11677);
and U12756 (N_12756,N_11097,N_11788);
or U12757 (N_12757,N_11475,N_11972);
and U12758 (N_12758,N_11652,N_11509);
or U12759 (N_12759,N_11804,N_11281);
and U12760 (N_12760,N_11227,N_11775);
nor U12761 (N_12761,N_11561,N_11559);
xor U12762 (N_12762,N_11835,N_11697);
nand U12763 (N_12763,N_11028,N_11515);
and U12764 (N_12764,N_11289,N_11714);
and U12765 (N_12765,N_11573,N_11753);
nand U12766 (N_12766,N_11549,N_11402);
xnor U12767 (N_12767,N_11863,N_11301);
xnor U12768 (N_12768,N_11606,N_11549);
nor U12769 (N_12769,N_11067,N_11736);
nor U12770 (N_12770,N_11964,N_11176);
nand U12771 (N_12771,N_11568,N_11616);
nand U12772 (N_12772,N_11217,N_11463);
and U12773 (N_12773,N_11734,N_11144);
nand U12774 (N_12774,N_11827,N_11463);
xor U12775 (N_12775,N_11568,N_11467);
xor U12776 (N_12776,N_11667,N_11798);
and U12777 (N_12777,N_11817,N_11985);
nand U12778 (N_12778,N_11858,N_11081);
and U12779 (N_12779,N_11663,N_11056);
and U12780 (N_12780,N_11701,N_11279);
xnor U12781 (N_12781,N_11596,N_11815);
nand U12782 (N_12782,N_11442,N_11853);
and U12783 (N_12783,N_11904,N_11638);
xnor U12784 (N_12784,N_11593,N_11099);
and U12785 (N_12785,N_11112,N_11708);
and U12786 (N_12786,N_11963,N_11516);
nor U12787 (N_12787,N_11792,N_11620);
nand U12788 (N_12788,N_11730,N_11667);
nor U12789 (N_12789,N_11257,N_11626);
nand U12790 (N_12790,N_11963,N_11858);
nand U12791 (N_12791,N_11002,N_11592);
or U12792 (N_12792,N_11559,N_11723);
nor U12793 (N_12793,N_11401,N_11638);
or U12794 (N_12794,N_11816,N_11298);
nand U12795 (N_12795,N_11300,N_11602);
or U12796 (N_12796,N_11696,N_11087);
or U12797 (N_12797,N_11474,N_11419);
and U12798 (N_12798,N_11880,N_11980);
and U12799 (N_12799,N_11487,N_11360);
xnor U12800 (N_12800,N_11830,N_11056);
and U12801 (N_12801,N_11121,N_11043);
nor U12802 (N_12802,N_11114,N_11891);
and U12803 (N_12803,N_11176,N_11238);
xor U12804 (N_12804,N_11553,N_11783);
or U12805 (N_12805,N_11190,N_11054);
xor U12806 (N_12806,N_11846,N_11379);
nand U12807 (N_12807,N_11305,N_11237);
nand U12808 (N_12808,N_11467,N_11523);
nor U12809 (N_12809,N_11944,N_11244);
and U12810 (N_12810,N_11185,N_11338);
nand U12811 (N_12811,N_11906,N_11765);
nand U12812 (N_12812,N_11487,N_11576);
and U12813 (N_12813,N_11555,N_11757);
xor U12814 (N_12814,N_11593,N_11006);
xnor U12815 (N_12815,N_11334,N_11247);
nor U12816 (N_12816,N_11486,N_11492);
nand U12817 (N_12817,N_11079,N_11741);
nand U12818 (N_12818,N_11692,N_11293);
nor U12819 (N_12819,N_11391,N_11771);
xnor U12820 (N_12820,N_11780,N_11962);
or U12821 (N_12821,N_11549,N_11357);
nand U12822 (N_12822,N_11737,N_11342);
xor U12823 (N_12823,N_11730,N_11217);
or U12824 (N_12824,N_11192,N_11776);
or U12825 (N_12825,N_11031,N_11819);
xor U12826 (N_12826,N_11651,N_11795);
nand U12827 (N_12827,N_11518,N_11098);
nand U12828 (N_12828,N_11185,N_11870);
xor U12829 (N_12829,N_11072,N_11005);
or U12830 (N_12830,N_11664,N_11951);
nand U12831 (N_12831,N_11910,N_11490);
nor U12832 (N_12832,N_11938,N_11374);
xor U12833 (N_12833,N_11621,N_11040);
xnor U12834 (N_12834,N_11834,N_11330);
nand U12835 (N_12835,N_11564,N_11858);
nand U12836 (N_12836,N_11204,N_11192);
nand U12837 (N_12837,N_11854,N_11362);
nor U12838 (N_12838,N_11426,N_11428);
nor U12839 (N_12839,N_11502,N_11617);
xor U12840 (N_12840,N_11328,N_11985);
nor U12841 (N_12841,N_11178,N_11030);
xor U12842 (N_12842,N_11134,N_11546);
nor U12843 (N_12843,N_11865,N_11026);
xnor U12844 (N_12844,N_11291,N_11180);
xor U12845 (N_12845,N_11405,N_11050);
or U12846 (N_12846,N_11252,N_11170);
or U12847 (N_12847,N_11417,N_11858);
nand U12848 (N_12848,N_11792,N_11209);
or U12849 (N_12849,N_11375,N_11831);
nand U12850 (N_12850,N_11314,N_11189);
nor U12851 (N_12851,N_11349,N_11079);
nand U12852 (N_12852,N_11738,N_11902);
xor U12853 (N_12853,N_11960,N_11523);
xnor U12854 (N_12854,N_11353,N_11785);
or U12855 (N_12855,N_11057,N_11690);
nand U12856 (N_12856,N_11284,N_11421);
and U12857 (N_12857,N_11760,N_11266);
xnor U12858 (N_12858,N_11866,N_11344);
nand U12859 (N_12859,N_11720,N_11117);
nand U12860 (N_12860,N_11849,N_11404);
xor U12861 (N_12861,N_11637,N_11339);
xor U12862 (N_12862,N_11272,N_11759);
and U12863 (N_12863,N_11664,N_11282);
nor U12864 (N_12864,N_11075,N_11659);
or U12865 (N_12865,N_11697,N_11264);
xor U12866 (N_12866,N_11023,N_11353);
xnor U12867 (N_12867,N_11027,N_11096);
nor U12868 (N_12868,N_11526,N_11692);
or U12869 (N_12869,N_11580,N_11915);
nor U12870 (N_12870,N_11417,N_11743);
nor U12871 (N_12871,N_11669,N_11622);
and U12872 (N_12872,N_11064,N_11052);
and U12873 (N_12873,N_11308,N_11720);
or U12874 (N_12874,N_11313,N_11402);
nor U12875 (N_12875,N_11252,N_11966);
xnor U12876 (N_12876,N_11402,N_11026);
xor U12877 (N_12877,N_11146,N_11918);
nor U12878 (N_12878,N_11526,N_11650);
and U12879 (N_12879,N_11138,N_11977);
xnor U12880 (N_12880,N_11939,N_11476);
or U12881 (N_12881,N_11546,N_11816);
and U12882 (N_12882,N_11080,N_11059);
and U12883 (N_12883,N_11660,N_11681);
xor U12884 (N_12884,N_11942,N_11129);
xnor U12885 (N_12885,N_11481,N_11658);
or U12886 (N_12886,N_11593,N_11612);
nor U12887 (N_12887,N_11714,N_11806);
nor U12888 (N_12888,N_11261,N_11666);
or U12889 (N_12889,N_11435,N_11239);
or U12890 (N_12890,N_11007,N_11758);
nand U12891 (N_12891,N_11960,N_11240);
nand U12892 (N_12892,N_11789,N_11658);
or U12893 (N_12893,N_11663,N_11521);
or U12894 (N_12894,N_11372,N_11128);
nor U12895 (N_12895,N_11587,N_11281);
nand U12896 (N_12896,N_11744,N_11508);
and U12897 (N_12897,N_11327,N_11470);
nor U12898 (N_12898,N_11231,N_11421);
and U12899 (N_12899,N_11314,N_11141);
xnor U12900 (N_12900,N_11321,N_11066);
nand U12901 (N_12901,N_11562,N_11391);
nand U12902 (N_12902,N_11488,N_11923);
nand U12903 (N_12903,N_11671,N_11448);
and U12904 (N_12904,N_11600,N_11913);
nand U12905 (N_12905,N_11648,N_11966);
nand U12906 (N_12906,N_11851,N_11797);
nand U12907 (N_12907,N_11924,N_11361);
and U12908 (N_12908,N_11329,N_11138);
xor U12909 (N_12909,N_11537,N_11902);
nand U12910 (N_12910,N_11046,N_11787);
xnor U12911 (N_12911,N_11999,N_11989);
and U12912 (N_12912,N_11300,N_11849);
xor U12913 (N_12913,N_11199,N_11586);
and U12914 (N_12914,N_11105,N_11319);
xnor U12915 (N_12915,N_11763,N_11461);
or U12916 (N_12916,N_11629,N_11965);
nand U12917 (N_12917,N_11181,N_11448);
xor U12918 (N_12918,N_11092,N_11654);
nor U12919 (N_12919,N_11889,N_11218);
nand U12920 (N_12920,N_11516,N_11597);
xnor U12921 (N_12921,N_11570,N_11295);
xor U12922 (N_12922,N_11318,N_11266);
xnor U12923 (N_12923,N_11621,N_11787);
xor U12924 (N_12924,N_11229,N_11050);
and U12925 (N_12925,N_11594,N_11907);
and U12926 (N_12926,N_11181,N_11633);
nor U12927 (N_12927,N_11973,N_11741);
nand U12928 (N_12928,N_11171,N_11509);
nand U12929 (N_12929,N_11122,N_11537);
nand U12930 (N_12930,N_11608,N_11314);
xor U12931 (N_12931,N_11001,N_11479);
xor U12932 (N_12932,N_11520,N_11181);
and U12933 (N_12933,N_11700,N_11096);
xor U12934 (N_12934,N_11440,N_11330);
or U12935 (N_12935,N_11620,N_11856);
xor U12936 (N_12936,N_11576,N_11115);
and U12937 (N_12937,N_11532,N_11420);
nand U12938 (N_12938,N_11715,N_11751);
nand U12939 (N_12939,N_11149,N_11817);
nand U12940 (N_12940,N_11913,N_11987);
or U12941 (N_12941,N_11931,N_11484);
nand U12942 (N_12942,N_11948,N_11115);
xnor U12943 (N_12943,N_11390,N_11699);
nor U12944 (N_12944,N_11946,N_11591);
nor U12945 (N_12945,N_11890,N_11912);
nand U12946 (N_12946,N_11729,N_11391);
nand U12947 (N_12947,N_11950,N_11966);
nand U12948 (N_12948,N_11339,N_11596);
or U12949 (N_12949,N_11296,N_11838);
or U12950 (N_12950,N_11784,N_11963);
and U12951 (N_12951,N_11204,N_11293);
nor U12952 (N_12952,N_11754,N_11825);
xnor U12953 (N_12953,N_11135,N_11669);
or U12954 (N_12954,N_11517,N_11217);
nand U12955 (N_12955,N_11513,N_11721);
or U12956 (N_12956,N_11072,N_11319);
nand U12957 (N_12957,N_11364,N_11705);
nor U12958 (N_12958,N_11275,N_11104);
or U12959 (N_12959,N_11884,N_11545);
and U12960 (N_12960,N_11257,N_11410);
xor U12961 (N_12961,N_11192,N_11180);
xor U12962 (N_12962,N_11881,N_11022);
or U12963 (N_12963,N_11290,N_11446);
nand U12964 (N_12964,N_11719,N_11621);
xnor U12965 (N_12965,N_11826,N_11732);
nor U12966 (N_12966,N_11056,N_11540);
and U12967 (N_12967,N_11484,N_11920);
nand U12968 (N_12968,N_11948,N_11193);
nand U12969 (N_12969,N_11363,N_11163);
and U12970 (N_12970,N_11997,N_11486);
nand U12971 (N_12971,N_11173,N_11912);
nand U12972 (N_12972,N_11972,N_11415);
nor U12973 (N_12973,N_11611,N_11789);
xnor U12974 (N_12974,N_11624,N_11127);
xnor U12975 (N_12975,N_11638,N_11430);
xnor U12976 (N_12976,N_11277,N_11381);
nand U12977 (N_12977,N_11801,N_11820);
and U12978 (N_12978,N_11873,N_11224);
nand U12979 (N_12979,N_11327,N_11020);
nor U12980 (N_12980,N_11113,N_11165);
nand U12981 (N_12981,N_11580,N_11602);
or U12982 (N_12982,N_11792,N_11893);
xnor U12983 (N_12983,N_11750,N_11446);
nor U12984 (N_12984,N_11240,N_11672);
nand U12985 (N_12985,N_11012,N_11055);
nand U12986 (N_12986,N_11567,N_11550);
xor U12987 (N_12987,N_11622,N_11218);
nor U12988 (N_12988,N_11034,N_11912);
nand U12989 (N_12989,N_11187,N_11286);
xor U12990 (N_12990,N_11457,N_11308);
or U12991 (N_12991,N_11450,N_11220);
or U12992 (N_12992,N_11579,N_11343);
or U12993 (N_12993,N_11110,N_11897);
nor U12994 (N_12994,N_11199,N_11580);
xnor U12995 (N_12995,N_11845,N_11988);
or U12996 (N_12996,N_11746,N_11251);
or U12997 (N_12997,N_11076,N_11104);
nor U12998 (N_12998,N_11457,N_11194);
xor U12999 (N_12999,N_11886,N_11417);
or U13000 (N_13000,N_12229,N_12350);
or U13001 (N_13001,N_12462,N_12062);
nor U13002 (N_13002,N_12367,N_12885);
or U13003 (N_13003,N_12443,N_12594);
xnor U13004 (N_13004,N_12656,N_12976);
nand U13005 (N_13005,N_12328,N_12822);
and U13006 (N_13006,N_12803,N_12863);
xnor U13007 (N_13007,N_12572,N_12403);
nor U13008 (N_13008,N_12301,N_12813);
nand U13009 (N_13009,N_12986,N_12456);
xnor U13010 (N_13010,N_12472,N_12398);
xnor U13011 (N_13011,N_12578,N_12374);
nor U13012 (N_13012,N_12510,N_12162);
nor U13013 (N_13013,N_12774,N_12867);
or U13014 (N_13014,N_12120,N_12587);
nor U13015 (N_13015,N_12382,N_12104);
and U13016 (N_13016,N_12529,N_12676);
nand U13017 (N_13017,N_12596,N_12818);
nand U13018 (N_13018,N_12408,N_12371);
nor U13019 (N_13019,N_12233,N_12297);
xor U13020 (N_13020,N_12571,N_12075);
and U13021 (N_13021,N_12722,N_12618);
and U13022 (N_13022,N_12261,N_12670);
and U13023 (N_13023,N_12092,N_12216);
or U13024 (N_13024,N_12061,N_12714);
nor U13025 (N_13025,N_12474,N_12019);
or U13026 (N_13026,N_12138,N_12673);
or U13027 (N_13027,N_12772,N_12256);
nand U13028 (N_13028,N_12479,N_12645);
xnor U13029 (N_13029,N_12097,N_12943);
and U13030 (N_13030,N_12900,N_12751);
or U13031 (N_13031,N_12991,N_12484);
or U13032 (N_13032,N_12210,N_12005);
nand U13033 (N_13033,N_12801,N_12276);
nor U13034 (N_13034,N_12202,N_12548);
and U13035 (N_13035,N_12190,N_12044);
xnor U13036 (N_13036,N_12154,N_12112);
nand U13037 (N_13037,N_12440,N_12808);
and U13038 (N_13038,N_12681,N_12070);
and U13039 (N_13039,N_12300,N_12105);
nor U13040 (N_13040,N_12150,N_12320);
nand U13041 (N_13041,N_12675,N_12013);
xnor U13042 (N_13042,N_12362,N_12195);
nor U13043 (N_13043,N_12607,N_12208);
nor U13044 (N_13044,N_12537,N_12568);
and U13045 (N_13045,N_12346,N_12585);
nor U13046 (N_13046,N_12661,N_12080);
nor U13047 (N_13047,N_12996,N_12187);
and U13048 (N_13048,N_12394,N_12789);
nand U13049 (N_13049,N_12875,N_12004);
nand U13050 (N_13050,N_12999,N_12836);
nand U13051 (N_13051,N_12145,N_12575);
nand U13052 (N_13052,N_12762,N_12515);
or U13053 (N_13053,N_12207,N_12816);
xor U13054 (N_13054,N_12299,N_12153);
nor U13055 (N_13055,N_12020,N_12255);
or U13056 (N_13056,N_12824,N_12418);
or U13057 (N_13057,N_12071,N_12878);
or U13058 (N_13058,N_12805,N_12702);
nand U13059 (N_13059,N_12550,N_12122);
and U13060 (N_13060,N_12014,N_12054);
xnor U13061 (N_13061,N_12000,N_12630);
nor U13062 (N_13062,N_12228,N_12570);
nor U13063 (N_13063,N_12525,N_12118);
xnor U13064 (N_13064,N_12345,N_12002);
or U13065 (N_13065,N_12205,N_12627);
nand U13066 (N_13066,N_12965,N_12954);
or U13067 (N_13067,N_12703,N_12903);
nor U13068 (N_13068,N_12876,N_12874);
nand U13069 (N_13069,N_12017,N_12414);
xnor U13070 (N_13070,N_12533,N_12919);
xnor U13071 (N_13071,N_12284,N_12921);
xnor U13072 (N_13072,N_12471,N_12436);
nand U13073 (N_13073,N_12639,N_12599);
xnor U13074 (N_13074,N_12098,N_12700);
xnor U13075 (N_13075,N_12896,N_12707);
xnor U13076 (N_13076,N_12450,N_12696);
nor U13077 (N_13077,N_12370,N_12623);
and U13078 (N_13078,N_12087,N_12952);
nor U13079 (N_13079,N_12901,N_12073);
nor U13080 (N_13080,N_12756,N_12137);
xor U13081 (N_13081,N_12736,N_12956);
and U13082 (N_13082,N_12657,N_12308);
nor U13083 (N_13083,N_12333,N_12492);
nor U13084 (N_13084,N_12704,N_12468);
or U13085 (N_13085,N_12183,N_12877);
xnor U13086 (N_13086,N_12754,N_12306);
xor U13087 (N_13087,N_12163,N_12518);
or U13088 (N_13088,N_12846,N_12995);
nor U13089 (N_13089,N_12144,N_12953);
or U13090 (N_13090,N_12724,N_12304);
or U13091 (N_13091,N_12902,N_12633);
or U13092 (N_13092,N_12043,N_12650);
and U13093 (N_13093,N_12771,N_12680);
and U13094 (N_13094,N_12264,N_12740);
nand U13095 (N_13095,N_12540,N_12409);
and U13096 (N_13096,N_12384,N_12318);
xnor U13097 (N_13097,N_12981,N_12984);
nand U13098 (N_13098,N_12348,N_12536);
nand U13099 (N_13099,N_12465,N_12620);
nand U13100 (N_13100,N_12884,N_12880);
or U13101 (N_13101,N_12313,N_12742);
xor U13102 (N_13102,N_12032,N_12835);
nand U13103 (N_13103,N_12966,N_12252);
and U13104 (N_13104,N_12402,N_12692);
xor U13105 (N_13105,N_12767,N_12850);
or U13106 (N_13106,N_12106,N_12904);
and U13107 (N_13107,N_12937,N_12231);
xor U13108 (N_13108,N_12438,N_12602);
and U13109 (N_13109,N_12505,N_12040);
nand U13110 (N_13110,N_12315,N_12164);
and U13111 (N_13111,N_12033,N_12725);
nor U13112 (N_13112,N_12082,N_12636);
or U13113 (N_13113,N_12491,N_12101);
or U13114 (N_13114,N_12432,N_12539);
nand U13115 (N_13115,N_12612,N_12891);
and U13116 (N_13116,N_12227,N_12616);
xnor U13117 (N_13117,N_12797,N_12871);
and U13118 (N_13118,N_12084,N_12589);
and U13119 (N_13119,N_12385,N_12041);
and U13120 (N_13120,N_12157,N_12528);
or U13121 (N_13121,N_12938,N_12775);
nand U13122 (N_13122,N_12509,N_12982);
nand U13123 (N_13123,N_12974,N_12972);
nand U13124 (N_13124,N_12064,N_12343);
xor U13125 (N_13125,N_12893,N_12679);
or U13126 (N_13126,N_12219,N_12830);
and U13127 (N_13127,N_12729,N_12460);
nand U13128 (N_13128,N_12928,N_12522);
nand U13129 (N_13129,N_12372,N_12457);
nor U13130 (N_13130,N_12785,N_12842);
and U13131 (N_13131,N_12720,N_12425);
nand U13132 (N_13132,N_12360,N_12147);
or U13133 (N_13133,N_12269,N_12251);
nand U13134 (N_13134,N_12286,N_12314);
nand U13135 (N_13135,N_12834,N_12215);
or U13136 (N_13136,N_12429,N_12807);
nand U13137 (N_13137,N_12547,N_12095);
nor U13138 (N_13138,N_12086,N_12180);
nor U13139 (N_13139,N_12669,N_12794);
nor U13140 (N_13140,N_12427,N_12331);
xor U13141 (N_13141,N_12796,N_12191);
and U13142 (N_13142,N_12694,N_12790);
and U13143 (N_13143,N_12685,N_12591);
or U13144 (N_13144,N_12151,N_12827);
nor U13145 (N_13145,N_12977,N_12378);
and U13146 (N_13146,N_12201,N_12747);
nand U13147 (N_13147,N_12173,N_12667);
or U13148 (N_13148,N_12065,N_12873);
nor U13149 (N_13149,N_12373,N_12036);
nand U13150 (N_13150,N_12366,N_12665);
or U13151 (N_13151,N_12341,N_12584);
nor U13152 (N_13152,N_12496,N_12718);
and U13153 (N_13153,N_12689,N_12609);
or U13154 (N_13154,N_12279,N_12200);
nand U13155 (N_13155,N_12400,N_12214);
xor U13156 (N_13156,N_12464,N_12752);
xor U13157 (N_13157,N_12165,N_12294);
and U13158 (N_13158,N_12504,N_12149);
xor U13159 (N_13159,N_12375,N_12812);
xnor U13160 (N_13160,N_12424,N_12778);
or U13161 (N_13161,N_12833,N_12254);
and U13162 (N_13162,N_12038,N_12635);
xor U13163 (N_13163,N_12381,N_12380);
and U13164 (N_13164,N_12125,N_12579);
or U13165 (N_13165,N_12107,N_12532);
xnor U13166 (N_13166,N_12887,N_12483);
nor U13167 (N_13167,N_12798,N_12148);
nand U13168 (N_13168,N_12335,N_12705);
xor U13169 (N_13169,N_12793,N_12644);
xor U13170 (N_13170,N_12079,N_12845);
xnor U13171 (N_13171,N_12419,N_12853);
nand U13172 (N_13172,N_12407,N_12161);
or U13173 (N_13173,N_12349,N_12783);
xor U13174 (N_13174,N_12899,N_12625);
xor U13175 (N_13175,N_12950,N_12958);
or U13176 (N_13176,N_12037,N_12170);
or U13177 (N_13177,N_12434,N_12970);
nor U13178 (N_13178,N_12222,N_12121);
nand U13179 (N_13179,N_12908,N_12776);
and U13180 (N_13180,N_12668,N_12734);
nand U13181 (N_13181,N_12291,N_12114);
or U13182 (N_13182,N_12906,N_12624);
nand U13183 (N_13183,N_12626,N_12099);
nand U13184 (N_13184,N_12964,N_12021);
nand U13185 (N_13185,N_12699,N_12749);
nand U13186 (N_13186,N_12124,N_12993);
or U13187 (N_13187,N_12733,N_12588);
nand U13188 (N_13188,N_12259,N_12779);
xnor U13189 (N_13189,N_12199,N_12486);
nand U13190 (N_13190,N_12482,N_12865);
or U13191 (N_13191,N_12898,N_12327);
nand U13192 (N_13192,N_12185,N_12915);
xor U13193 (N_13193,N_12662,N_12193);
nor U13194 (N_13194,N_12177,N_12340);
xnor U13195 (N_13195,N_12130,N_12544);
nor U13196 (N_13196,N_12946,N_12879);
xor U13197 (N_13197,N_12174,N_12473);
or U13198 (N_13198,N_12136,N_12049);
nor U13199 (N_13199,N_12171,N_12452);
or U13200 (N_13200,N_12693,N_12849);
or U13201 (N_13201,N_12586,N_12866);
nor U13202 (N_13202,N_12811,N_12060);
xor U13203 (N_13203,N_12111,N_12059);
and U13204 (N_13204,N_12344,N_12182);
nand U13205 (N_13205,N_12412,N_12444);
nand U13206 (N_13206,N_12316,N_12085);
nand U13207 (N_13207,N_12988,N_12234);
xnor U13208 (N_13208,N_12067,N_12319);
nand U13209 (N_13209,N_12446,N_12016);
nand U13210 (N_13210,N_12433,N_12860);
xor U13211 (N_13211,N_12422,N_12451);
or U13212 (N_13212,N_12249,N_12029);
nand U13213 (N_13213,N_12709,N_12129);
and U13214 (N_13214,N_12851,N_12166);
and U13215 (N_13215,N_12477,N_12562);
nor U13216 (N_13216,N_12244,N_12167);
or U13217 (N_13217,N_12189,N_12078);
nand U13218 (N_13218,N_12501,N_12194);
nor U13219 (N_13219,N_12514,N_12405);
nor U13220 (N_13220,N_12302,N_12310);
and U13221 (N_13221,N_12777,N_12421);
nand U13222 (N_13222,N_12628,N_12695);
xnor U13223 (N_13223,N_12574,N_12337);
xnor U13224 (N_13224,N_12746,N_12218);
xor U13225 (N_13225,N_12453,N_12632);
nand U13226 (N_13226,N_12782,N_12738);
or U13227 (N_13227,N_12159,N_12534);
nand U13228 (N_13228,N_12927,N_12848);
nand U13229 (N_13229,N_12417,N_12888);
xor U13230 (N_13230,N_12963,N_12292);
nand U13231 (N_13231,N_12930,N_12076);
xnor U13232 (N_13232,N_12828,N_12862);
and U13233 (N_13233,N_12712,N_12911);
or U13234 (N_13234,N_12238,N_12933);
nand U13235 (N_13235,N_12006,N_12897);
nand U13236 (N_13236,N_12806,N_12196);
nand U13237 (N_13237,N_12882,N_12719);
xor U13238 (N_13238,N_12223,N_12241);
nor U13239 (N_13239,N_12230,N_12128);
and U13240 (N_13240,N_12047,N_12455);
and U13241 (N_13241,N_12942,N_12117);
and U13242 (N_13242,N_12271,N_12442);
xnor U13243 (N_13243,N_12131,N_12389);
and U13244 (N_13244,N_12913,N_12413);
and U13245 (N_13245,N_12357,N_12437);
nand U13246 (N_13246,N_12723,N_12192);
or U13247 (N_13247,N_12593,N_12945);
or U13248 (N_13248,N_12905,N_12659);
or U13249 (N_13249,N_12998,N_12478);
and U13250 (N_13250,N_12449,N_12387);
nand U13251 (N_13251,N_12133,N_12975);
and U13252 (N_13252,N_12369,N_12935);
xnor U13253 (N_13253,N_12081,N_12728);
nor U13254 (N_13254,N_12758,N_12135);
and U13255 (N_13255,N_12245,N_12353);
and U13256 (N_13256,N_12861,N_12463);
nand U13257 (N_13257,N_12494,N_12072);
or U13258 (N_13258,N_12990,N_12495);
nor U13259 (N_13259,N_12557,N_12603);
and U13260 (N_13260,N_12856,N_12441);
or U13261 (N_13261,N_12717,N_12521);
nand U13262 (N_13262,N_12654,N_12088);
nand U13263 (N_13263,N_12426,N_12221);
nor U13264 (N_13264,N_12430,N_12595);
xor U13265 (N_13265,N_12889,N_12293);
or U13266 (N_13266,N_12027,N_12140);
nand U13267 (N_13267,N_12641,N_12209);
and U13268 (N_13268,N_12045,N_12459);
nor U13269 (N_13269,N_12831,N_12466);
nand U13270 (N_13270,N_12947,N_12487);
and U13271 (N_13271,N_12103,N_12590);
nor U13272 (N_13272,N_12172,N_12894);
nor U13273 (N_13273,N_12461,N_12892);
nand U13274 (N_13274,N_12090,N_12610);
and U13275 (N_13275,N_12858,N_12715);
nand U13276 (N_13276,N_12920,N_12325);
xor U13277 (N_13277,N_12934,N_12428);
nand U13278 (N_13278,N_12277,N_12458);
xnor U13279 (N_13279,N_12566,N_12141);
xor U13280 (N_13280,N_12158,N_12697);
nand U13281 (N_13281,N_12666,N_12820);
nand U13282 (N_13282,N_12010,N_12500);
or U13283 (N_13283,N_12576,N_12924);
and U13284 (N_13284,N_12439,N_12220);
nor U13285 (N_13285,N_12470,N_12770);
nand U13286 (N_13286,N_12268,N_12094);
nand U13287 (N_13287,N_12926,N_12755);
xnor U13288 (N_13288,N_12569,N_12211);
xnor U13289 (N_13289,N_12787,N_12476);
nor U13290 (N_13290,N_12731,N_12007);
or U13291 (N_13291,N_12139,N_12317);
xor U13292 (N_13292,N_12792,N_12802);
nor U13293 (N_13293,N_12295,N_12146);
nand U13294 (N_13294,N_12653,N_12334);
xor U13295 (N_13295,N_12288,N_12647);
or U13296 (N_13296,N_12757,N_12561);
nand U13297 (N_13297,N_12730,N_12169);
xor U13298 (N_13298,N_12281,N_12795);
or U13299 (N_13299,N_12753,N_12025);
and U13300 (N_13300,N_12677,N_12614);
or U13301 (N_13301,N_12634,N_12022);
and U13302 (N_13302,N_12324,N_12030);
nand U13303 (N_13303,N_12556,N_12186);
and U13304 (N_13304,N_12311,N_12872);
or U13305 (N_13305,N_12018,N_12265);
and U13306 (N_13306,N_12939,N_12212);
nor U13307 (N_13307,N_12026,N_12663);
xnor U13308 (N_13308,N_12052,N_12621);
and U13309 (N_13309,N_12608,N_12322);
and U13310 (N_13310,N_12870,N_12411);
nor U13311 (N_13311,N_12638,N_12431);
nand U13312 (N_13312,N_12989,N_12985);
nor U13313 (N_13313,N_12386,N_12881);
or U13314 (N_13314,N_12664,N_12352);
and U13315 (N_13315,N_12829,N_12339);
or U13316 (N_13316,N_12282,N_12960);
nor U13317 (N_13317,N_12857,N_12267);
nor U13318 (N_13318,N_12309,N_12713);
xnor U13319 (N_13319,N_12936,N_12840);
xnor U13320 (N_13320,N_12296,N_12356);
xor U13321 (N_13321,N_12330,N_12711);
or U13322 (N_13322,N_12489,N_12617);
xor U13323 (N_13323,N_12968,N_12069);
nor U13324 (N_13324,N_12012,N_12395);
and U13325 (N_13325,N_12406,N_12217);
or U13326 (N_13326,N_12825,N_12706);
or U13327 (N_13327,N_12009,N_12321);
nor U13328 (N_13328,N_12601,N_12275);
nor U13329 (N_13329,N_12181,N_12855);
and U13330 (N_13330,N_12629,N_12535);
nor U13331 (N_13331,N_12542,N_12074);
or U13332 (N_13332,N_12961,N_12499);
xor U13333 (N_13333,N_12583,N_12929);
or U13334 (N_13334,N_12615,N_12143);
xor U13335 (N_13335,N_12179,N_12710);
and U13336 (N_13336,N_12741,N_12132);
nand U13337 (N_13337,N_12978,N_12110);
nand U13338 (N_13338,N_12839,N_12910);
nand U13339 (N_13339,N_12962,N_12931);
nor U13340 (N_13340,N_12916,N_12864);
xor U13341 (N_13341,N_12001,N_12526);
or U13342 (N_13342,N_12726,N_12015);
or U13343 (N_13343,N_12655,N_12788);
and U13344 (N_13344,N_12843,N_12404);
nand U13345 (N_13345,N_12979,N_12034);
xor U13346 (N_13346,N_12011,N_12160);
xnor U13347 (N_13347,N_12410,N_12298);
or U13348 (N_13348,N_12435,N_12769);
or U13349 (N_13349,N_12914,N_12469);
xor U13350 (N_13350,N_12347,N_12511);
xnor U13351 (N_13351,N_12113,N_12361);
and U13352 (N_13352,N_12203,N_12134);
nor U13353 (N_13353,N_12396,N_12716);
nand U13354 (N_13354,N_12498,N_12246);
or U13355 (N_13355,N_12605,N_12804);
nor U13356 (N_13356,N_12683,N_12280);
and U13357 (N_13357,N_12581,N_12109);
or U13358 (N_13358,N_12832,N_12543);
and U13359 (N_13359,N_12213,N_12648);
nand U13360 (N_13360,N_12643,N_12250);
or U13361 (N_13361,N_12949,N_12688);
nor U13362 (N_13362,N_12721,N_12024);
and U13363 (N_13363,N_12155,N_12563);
xor U13364 (N_13364,N_12156,N_12102);
xnor U13365 (N_13365,N_12368,N_12243);
nor U13366 (N_13366,N_12508,N_12997);
nor U13367 (N_13367,N_12600,N_12278);
or U13368 (N_13368,N_12423,N_12671);
and U13369 (N_13369,N_12582,N_12690);
or U13370 (N_13370,N_12055,N_12948);
or U13371 (N_13371,N_12342,N_12819);
xnor U13372 (N_13372,N_12119,N_12239);
nand U13373 (N_13373,N_12674,N_12549);
nor U13374 (N_13374,N_12445,N_12480);
and U13375 (N_13375,N_12257,N_12743);
xor U13376 (N_13376,N_12454,N_12285);
nor U13377 (N_13377,N_12258,N_12305);
nor U13378 (N_13378,N_12115,N_12565);
xor U13379 (N_13379,N_12523,N_12980);
or U13380 (N_13380,N_12517,N_12791);
xor U13381 (N_13381,N_12520,N_12142);
nand U13382 (N_13382,N_12089,N_12003);
xor U13383 (N_13383,N_12058,N_12558);
and U13384 (N_13384,N_12039,N_12739);
nand U13385 (N_13385,N_12503,N_12555);
nor U13386 (N_13386,N_12527,N_12682);
xnor U13387 (N_13387,N_12691,N_12519);
nand U13388 (N_13388,N_12814,N_12765);
and U13389 (N_13389,N_12242,N_12289);
nor U13390 (N_13390,N_12925,N_12050);
xor U13391 (N_13391,N_12392,N_12750);
nor U13392 (N_13392,N_12168,N_12053);
or U13393 (N_13393,N_12598,N_12351);
or U13394 (N_13394,N_12323,N_12091);
and U13395 (N_13395,N_12266,N_12823);
and U13396 (N_13396,N_12274,N_12485);
and U13397 (N_13397,N_12573,N_12108);
and U13398 (N_13398,N_12096,N_12773);
xnor U13399 (N_13399,N_12761,N_12658);
xnor U13400 (N_13400,N_12048,N_12290);
nor U13401 (N_13401,N_12708,N_12068);
nor U13402 (N_13402,N_12987,N_12909);
and U13403 (N_13403,N_12760,N_12329);
and U13404 (N_13404,N_12401,N_12809);
and U13405 (N_13405,N_12057,N_12868);
nand U13406 (N_13406,N_12184,N_12838);
xnor U13407 (N_13407,N_12388,N_12225);
xor U13408 (N_13408,N_12545,N_12604);
and U13409 (N_13409,N_12237,N_12737);
or U13410 (N_13410,N_12530,N_12507);
nor U13411 (N_13411,N_12852,N_12907);
and U13412 (N_13412,N_12152,N_12992);
or U13413 (N_13413,N_12379,N_12895);
and U13414 (N_13414,N_12126,N_12232);
and U13415 (N_13415,N_12969,N_12475);
and U13416 (N_13416,N_12262,N_12732);
nand U13417 (N_13417,N_12748,N_12859);
xnor U13418 (N_13418,N_12397,N_12886);
or U13419 (N_13419,N_12056,N_12248);
xor U13420 (N_13420,N_12008,N_12235);
and U13421 (N_13421,N_12226,N_12844);
nor U13422 (N_13422,N_12567,N_12178);
nand U13423 (N_13423,N_12890,N_12516);
xor U13424 (N_13424,N_12497,N_12488);
or U13425 (N_13425,N_12869,N_12272);
or U13426 (N_13426,N_12263,N_12815);
and U13427 (N_13427,N_12780,N_12955);
xor U13428 (N_13428,N_12744,N_12512);
and U13429 (N_13429,N_12355,N_12642);
or U13430 (N_13430,N_12100,N_12240);
or U13431 (N_13431,N_12944,N_12932);
and U13432 (N_13432,N_12083,N_12764);
nor U13433 (N_13433,N_12391,N_12821);
nand U13434 (N_13434,N_12312,N_12784);
or U13435 (N_13435,N_12918,N_12541);
or U13436 (N_13436,N_12260,N_12678);
and U13437 (N_13437,N_12698,N_12253);
or U13438 (N_13438,N_12390,N_12383);
nor U13439 (N_13439,N_12652,N_12983);
or U13440 (N_13440,N_12538,N_12766);
and U13441 (N_13441,N_12051,N_12560);
and U13442 (N_13442,N_12273,N_12553);
nor U13443 (N_13443,N_12416,N_12420);
and U13444 (N_13444,N_12236,N_12377);
and U13445 (N_13445,N_12359,N_12922);
and U13446 (N_13446,N_12524,N_12967);
nand U13447 (N_13447,N_12204,N_12447);
xnor U13448 (N_13448,N_12364,N_12399);
nand U13449 (N_13449,N_12660,N_12684);
nand U13450 (N_13450,N_12551,N_12847);
xor U13451 (N_13451,N_12768,N_12837);
nand U13452 (N_13452,N_12606,N_12613);
xnor U13453 (N_13453,N_12363,N_12365);
nand U13454 (N_13454,N_12631,N_12611);
nor U13455 (N_13455,N_12940,N_12735);
nor U13456 (N_13456,N_12559,N_12123);
and U13457 (N_13457,N_12448,N_12687);
nor U13458 (N_13458,N_12197,N_12854);
or U13459 (N_13459,N_12959,N_12646);
and U13460 (N_13460,N_12307,N_12176);
nor U13461 (N_13461,N_12619,N_12912);
and U13462 (N_13462,N_12354,N_12127);
nor U13463 (N_13463,N_12467,N_12188);
xor U13464 (N_13464,N_12941,N_12332);
xor U13465 (N_13465,N_12031,N_12810);
nor U13466 (N_13466,N_12637,N_12336);
and U13467 (N_13467,N_12554,N_12923);
nand U13468 (N_13468,N_12577,N_12303);
and U13469 (N_13469,N_12649,N_12531);
and U13470 (N_13470,N_12622,N_12066);
nor U13471 (N_13471,N_12973,N_12490);
and U13472 (N_13472,N_12415,N_12994);
nand U13473 (N_13473,N_12358,N_12917);
nand U13474 (N_13474,N_12786,N_12493);
and U13475 (N_13475,N_12841,N_12781);
xor U13476 (N_13476,N_12763,N_12376);
nor U13477 (N_13477,N_12028,N_12338);
and U13478 (N_13478,N_12826,N_12745);
and U13479 (N_13479,N_12502,N_12580);
nand U13480 (N_13480,N_12883,N_12564);
xor U13481 (N_13481,N_12077,N_12971);
nor U13482 (N_13482,N_12393,N_12175);
nor U13483 (N_13483,N_12546,N_12951);
xor U13484 (N_13484,N_12287,N_12759);
nor U13485 (N_13485,N_12701,N_12206);
and U13486 (N_13486,N_12063,N_12817);
nor U13487 (N_13487,N_12597,N_12042);
nor U13488 (N_13488,N_12023,N_12116);
nor U13489 (N_13489,N_12270,N_12727);
and U13490 (N_13490,N_12481,N_12640);
xor U13491 (N_13491,N_12592,N_12093);
xor U13492 (N_13492,N_12035,N_12326);
and U13493 (N_13493,N_12513,N_12799);
xnor U13494 (N_13494,N_12552,N_12800);
xor U13495 (N_13495,N_12283,N_12046);
or U13496 (N_13496,N_12957,N_12506);
nor U13497 (N_13497,N_12672,N_12651);
nor U13498 (N_13498,N_12686,N_12247);
nand U13499 (N_13499,N_12198,N_12224);
nor U13500 (N_13500,N_12394,N_12382);
nor U13501 (N_13501,N_12797,N_12306);
nor U13502 (N_13502,N_12299,N_12719);
or U13503 (N_13503,N_12755,N_12365);
or U13504 (N_13504,N_12372,N_12177);
nor U13505 (N_13505,N_12761,N_12150);
xor U13506 (N_13506,N_12753,N_12314);
nor U13507 (N_13507,N_12748,N_12201);
nor U13508 (N_13508,N_12336,N_12698);
xnor U13509 (N_13509,N_12618,N_12711);
xor U13510 (N_13510,N_12106,N_12768);
xnor U13511 (N_13511,N_12643,N_12665);
or U13512 (N_13512,N_12147,N_12947);
nand U13513 (N_13513,N_12385,N_12415);
xnor U13514 (N_13514,N_12304,N_12161);
or U13515 (N_13515,N_12323,N_12453);
or U13516 (N_13516,N_12483,N_12334);
and U13517 (N_13517,N_12241,N_12529);
xnor U13518 (N_13518,N_12208,N_12860);
xor U13519 (N_13519,N_12079,N_12099);
nand U13520 (N_13520,N_12752,N_12071);
nand U13521 (N_13521,N_12245,N_12588);
xor U13522 (N_13522,N_12141,N_12204);
and U13523 (N_13523,N_12761,N_12931);
and U13524 (N_13524,N_12843,N_12409);
or U13525 (N_13525,N_12923,N_12752);
and U13526 (N_13526,N_12486,N_12352);
xnor U13527 (N_13527,N_12393,N_12821);
or U13528 (N_13528,N_12708,N_12194);
or U13529 (N_13529,N_12395,N_12298);
xnor U13530 (N_13530,N_12779,N_12571);
and U13531 (N_13531,N_12664,N_12896);
and U13532 (N_13532,N_12986,N_12271);
nand U13533 (N_13533,N_12733,N_12554);
and U13534 (N_13534,N_12511,N_12127);
xnor U13535 (N_13535,N_12172,N_12601);
or U13536 (N_13536,N_12292,N_12781);
or U13537 (N_13537,N_12378,N_12980);
xor U13538 (N_13538,N_12235,N_12674);
nand U13539 (N_13539,N_12730,N_12408);
xor U13540 (N_13540,N_12205,N_12802);
nand U13541 (N_13541,N_12099,N_12402);
nor U13542 (N_13542,N_12955,N_12333);
or U13543 (N_13543,N_12197,N_12583);
and U13544 (N_13544,N_12494,N_12982);
xor U13545 (N_13545,N_12135,N_12731);
or U13546 (N_13546,N_12249,N_12790);
xor U13547 (N_13547,N_12748,N_12091);
nand U13548 (N_13548,N_12427,N_12894);
nor U13549 (N_13549,N_12355,N_12083);
nand U13550 (N_13550,N_12656,N_12220);
and U13551 (N_13551,N_12935,N_12487);
and U13552 (N_13552,N_12752,N_12380);
xnor U13553 (N_13553,N_12204,N_12700);
and U13554 (N_13554,N_12044,N_12049);
or U13555 (N_13555,N_12416,N_12774);
nor U13556 (N_13556,N_12075,N_12552);
nor U13557 (N_13557,N_12147,N_12862);
nand U13558 (N_13558,N_12343,N_12090);
nand U13559 (N_13559,N_12112,N_12741);
or U13560 (N_13560,N_12391,N_12141);
nor U13561 (N_13561,N_12469,N_12676);
nand U13562 (N_13562,N_12579,N_12869);
xnor U13563 (N_13563,N_12418,N_12120);
xnor U13564 (N_13564,N_12384,N_12370);
and U13565 (N_13565,N_12721,N_12729);
and U13566 (N_13566,N_12535,N_12961);
xnor U13567 (N_13567,N_12986,N_12988);
and U13568 (N_13568,N_12159,N_12415);
nor U13569 (N_13569,N_12921,N_12947);
nand U13570 (N_13570,N_12107,N_12030);
or U13571 (N_13571,N_12710,N_12012);
xnor U13572 (N_13572,N_12332,N_12280);
nand U13573 (N_13573,N_12859,N_12596);
or U13574 (N_13574,N_12711,N_12417);
or U13575 (N_13575,N_12692,N_12345);
or U13576 (N_13576,N_12864,N_12551);
or U13577 (N_13577,N_12241,N_12340);
and U13578 (N_13578,N_12777,N_12687);
or U13579 (N_13579,N_12553,N_12645);
nor U13580 (N_13580,N_12928,N_12728);
and U13581 (N_13581,N_12996,N_12957);
or U13582 (N_13582,N_12037,N_12513);
nor U13583 (N_13583,N_12172,N_12761);
or U13584 (N_13584,N_12918,N_12304);
and U13585 (N_13585,N_12703,N_12126);
xor U13586 (N_13586,N_12472,N_12590);
and U13587 (N_13587,N_12924,N_12403);
and U13588 (N_13588,N_12600,N_12810);
nand U13589 (N_13589,N_12731,N_12720);
or U13590 (N_13590,N_12489,N_12156);
xor U13591 (N_13591,N_12018,N_12840);
and U13592 (N_13592,N_12613,N_12142);
or U13593 (N_13593,N_12441,N_12168);
nand U13594 (N_13594,N_12527,N_12058);
or U13595 (N_13595,N_12551,N_12715);
nand U13596 (N_13596,N_12024,N_12846);
nor U13597 (N_13597,N_12428,N_12523);
or U13598 (N_13598,N_12640,N_12435);
xnor U13599 (N_13599,N_12124,N_12754);
nand U13600 (N_13600,N_12114,N_12502);
nor U13601 (N_13601,N_12426,N_12682);
and U13602 (N_13602,N_12721,N_12020);
or U13603 (N_13603,N_12525,N_12693);
xor U13604 (N_13604,N_12185,N_12289);
nand U13605 (N_13605,N_12723,N_12646);
or U13606 (N_13606,N_12380,N_12811);
or U13607 (N_13607,N_12992,N_12853);
xor U13608 (N_13608,N_12259,N_12227);
xnor U13609 (N_13609,N_12032,N_12067);
and U13610 (N_13610,N_12198,N_12168);
or U13611 (N_13611,N_12199,N_12237);
xnor U13612 (N_13612,N_12930,N_12588);
nand U13613 (N_13613,N_12830,N_12805);
nand U13614 (N_13614,N_12727,N_12476);
or U13615 (N_13615,N_12762,N_12755);
and U13616 (N_13616,N_12026,N_12217);
nand U13617 (N_13617,N_12636,N_12625);
nor U13618 (N_13618,N_12825,N_12153);
or U13619 (N_13619,N_12510,N_12908);
and U13620 (N_13620,N_12092,N_12218);
or U13621 (N_13621,N_12772,N_12602);
nand U13622 (N_13622,N_12839,N_12395);
and U13623 (N_13623,N_12798,N_12653);
nor U13624 (N_13624,N_12589,N_12273);
nor U13625 (N_13625,N_12382,N_12118);
or U13626 (N_13626,N_12351,N_12241);
or U13627 (N_13627,N_12301,N_12017);
nor U13628 (N_13628,N_12281,N_12932);
and U13629 (N_13629,N_12676,N_12749);
xnor U13630 (N_13630,N_12802,N_12920);
xnor U13631 (N_13631,N_12545,N_12421);
and U13632 (N_13632,N_12189,N_12507);
nand U13633 (N_13633,N_12617,N_12470);
or U13634 (N_13634,N_12191,N_12487);
or U13635 (N_13635,N_12604,N_12948);
nand U13636 (N_13636,N_12665,N_12543);
or U13637 (N_13637,N_12455,N_12865);
xor U13638 (N_13638,N_12874,N_12664);
nor U13639 (N_13639,N_12321,N_12738);
or U13640 (N_13640,N_12417,N_12270);
nand U13641 (N_13641,N_12689,N_12361);
or U13642 (N_13642,N_12266,N_12564);
xor U13643 (N_13643,N_12720,N_12224);
nand U13644 (N_13644,N_12587,N_12689);
xor U13645 (N_13645,N_12058,N_12719);
xnor U13646 (N_13646,N_12722,N_12309);
and U13647 (N_13647,N_12069,N_12687);
xor U13648 (N_13648,N_12853,N_12896);
or U13649 (N_13649,N_12042,N_12522);
and U13650 (N_13650,N_12646,N_12236);
and U13651 (N_13651,N_12439,N_12958);
xnor U13652 (N_13652,N_12236,N_12221);
nand U13653 (N_13653,N_12743,N_12945);
and U13654 (N_13654,N_12801,N_12381);
xnor U13655 (N_13655,N_12694,N_12979);
xor U13656 (N_13656,N_12602,N_12192);
nand U13657 (N_13657,N_12483,N_12226);
nand U13658 (N_13658,N_12485,N_12748);
nand U13659 (N_13659,N_12516,N_12884);
and U13660 (N_13660,N_12180,N_12380);
nand U13661 (N_13661,N_12680,N_12141);
xor U13662 (N_13662,N_12684,N_12011);
xnor U13663 (N_13663,N_12838,N_12572);
nand U13664 (N_13664,N_12511,N_12392);
or U13665 (N_13665,N_12411,N_12496);
nor U13666 (N_13666,N_12459,N_12086);
or U13667 (N_13667,N_12307,N_12853);
nor U13668 (N_13668,N_12318,N_12624);
nand U13669 (N_13669,N_12654,N_12364);
nor U13670 (N_13670,N_12166,N_12425);
nor U13671 (N_13671,N_12259,N_12297);
nor U13672 (N_13672,N_12115,N_12666);
nand U13673 (N_13673,N_12207,N_12784);
and U13674 (N_13674,N_12536,N_12710);
xor U13675 (N_13675,N_12441,N_12955);
and U13676 (N_13676,N_12709,N_12438);
and U13677 (N_13677,N_12264,N_12776);
or U13678 (N_13678,N_12826,N_12322);
xnor U13679 (N_13679,N_12364,N_12558);
nand U13680 (N_13680,N_12178,N_12239);
or U13681 (N_13681,N_12785,N_12571);
and U13682 (N_13682,N_12837,N_12699);
nor U13683 (N_13683,N_12370,N_12452);
or U13684 (N_13684,N_12276,N_12587);
nor U13685 (N_13685,N_12290,N_12688);
or U13686 (N_13686,N_12738,N_12680);
nand U13687 (N_13687,N_12813,N_12418);
nor U13688 (N_13688,N_12948,N_12354);
or U13689 (N_13689,N_12066,N_12872);
xnor U13690 (N_13690,N_12564,N_12118);
xnor U13691 (N_13691,N_12103,N_12682);
nand U13692 (N_13692,N_12197,N_12816);
nor U13693 (N_13693,N_12541,N_12367);
nor U13694 (N_13694,N_12215,N_12524);
or U13695 (N_13695,N_12179,N_12566);
xnor U13696 (N_13696,N_12897,N_12306);
nand U13697 (N_13697,N_12119,N_12949);
xor U13698 (N_13698,N_12319,N_12162);
nand U13699 (N_13699,N_12722,N_12864);
xnor U13700 (N_13700,N_12927,N_12581);
xor U13701 (N_13701,N_12761,N_12874);
nor U13702 (N_13702,N_12520,N_12800);
xor U13703 (N_13703,N_12161,N_12072);
and U13704 (N_13704,N_12665,N_12574);
nand U13705 (N_13705,N_12178,N_12216);
nand U13706 (N_13706,N_12812,N_12282);
nand U13707 (N_13707,N_12638,N_12458);
nand U13708 (N_13708,N_12949,N_12856);
or U13709 (N_13709,N_12267,N_12330);
or U13710 (N_13710,N_12626,N_12369);
xor U13711 (N_13711,N_12440,N_12754);
nor U13712 (N_13712,N_12398,N_12609);
nor U13713 (N_13713,N_12459,N_12327);
or U13714 (N_13714,N_12342,N_12517);
nand U13715 (N_13715,N_12950,N_12207);
nor U13716 (N_13716,N_12122,N_12560);
and U13717 (N_13717,N_12116,N_12884);
nand U13718 (N_13718,N_12743,N_12564);
or U13719 (N_13719,N_12828,N_12432);
or U13720 (N_13720,N_12272,N_12435);
or U13721 (N_13721,N_12618,N_12841);
or U13722 (N_13722,N_12490,N_12478);
xor U13723 (N_13723,N_12507,N_12893);
nor U13724 (N_13724,N_12601,N_12938);
nor U13725 (N_13725,N_12544,N_12565);
nor U13726 (N_13726,N_12365,N_12720);
nand U13727 (N_13727,N_12776,N_12795);
and U13728 (N_13728,N_12548,N_12405);
xor U13729 (N_13729,N_12014,N_12506);
and U13730 (N_13730,N_12834,N_12134);
or U13731 (N_13731,N_12804,N_12451);
nand U13732 (N_13732,N_12676,N_12896);
nor U13733 (N_13733,N_12974,N_12291);
nor U13734 (N_13734,N_12318,N_12424);
or U13735 (N_13735,N_12454,N_12868);
nand U13736 (N_13736,N_12509,N_12228);
nor U13737 (N_13737,N_12419,N_12607);
nand U13738 (N_13738,N_12603,N_12310);
and U13739 (N_13739,N_12630,N_12391);
and U13740 (N_13740,N_12303,N_12833);
nand U13741 (N_13741,N_12611,N_12901);
nand U13742 (N_13742,N_12658,N_12535);
xor U13743 (N_13743,N_12180,N_12561);
nor U13744 (N_13744,N_12169,N_12096);
and U13745 (N_13745,N_12234,N_12695);
and U13746 (N_13746,N_12688,N_12991);
or U13747 (N_13747,N_12742,N_12632);
nor U13748 (N_13748,N_12093,N_12860);
nor U13749 (N_13749,N_12829,N_12479);
nor U13750 (N_13750,N_12483,N_12098);
xnor U13751 (N_13751,N_12827,N_12953);
nand U13752 (N_13752,N_12110,N_12235);
nor U13753 (N_13753,N_12485,N_12553);
and U13754 (N_13754,N_12049,N_12366);
and U13755 (N_13755,N_12273,N_12261);
xnor U13756 (N_13756,N_12300,N_12305);
xor U13757 (N_13757,N_12957,N_12207);
and U13758 (N_13758,N_12958,N_12831);
nand U13759 (N_13759,N_12185,N_12656);
xor U13760 (N_13760,N_12712,N_12575);
or U13761 (N_13761,N_12821,N_12524);
and U13762 (N_13762,N_12370,N_12216);
and U13763 (N_13763,N_12882,N_12611);
nand U13764 (N_13764,N_12734,N_12757);
and U13765 (N_13765,N_12428,N_12353);
and U13766 (N_13766,N_12426,N_12274);
xnor U13767 (N_13767,N_12467,N_12222);
nor U13768 (N_13768,N_12308,N_12576);
xor U13769 (N_13769,N_12517,N_12782);
nor U13770 (N_13770,N_12432,N_12082);
nor U13771 (N_13771,N_12165,N_12888);
or U13772 (N_13772,N_12756,N_12440);
or U13773 (N_13773,N_12021,N_12925);
or U13774 (N_13774,N_12275,N_12529);
and U13775 (N_13775,N_12803,N_12407);
and U13776 (N_13776,N_12353,N_12930);
nand U13777 (N_13777,N_12648,N_12461);
nor U13778 (N_13778,N_12539,N_12490);
or U13779 (N_13779,N_12482,N_12064);
and U13780 (N_13780,N_12100,N_12454);
nand U13781 (N_13781,N_12180,N_12774);
nand U13782 (N_13782,N_12258,N_12261);
xnor U13783 (N_13783,N_12477,N_12154);
or U13784 (N_13784,N_12488,N_12893);
nand U13785 (N_13785,N_12617,N_12590);
or U13786 (N_13786,N_12863,N_12258);
xor U13787 (N_13787,N_12456,N_12009);
xnor U13788 (N_13788,N_12770,N_12958);
and U13789 (N_13789,N_12396,N_12057);
or U13790 (N_13790,N_12701,N_12043);
nand U13791 (N_13791,N_12466,N_12302);
nor U13792 (N_13792,N_12245,N_12475);
nor U13793 (N_13793,N_12939,N_12655);
and U13794 (N_13794,N_12523,N_12135);
and U13795 (N_13795,N_12374,N_12598);
xnor U13796 (N_13796,N_12529,N_12479);
nand U13797 (N_13797,N_12742,N_12723);
nor U13798 (N_13798,N_12218,N_12801);
nor U13799 (N_13799,N_12481,N_12088);
nand U13800 (N_13800,N_12788,N_12519);
nor U13801 (N_13801,N_12223,N_12274);
xor U13802 (N_13802,N_12380,N_12903);
nand U13803 (N_13803,N_12982,N_12422);
and U13804 (N_13804,N_12882,N_12018);
nor U13805 (N_13805,N_12797,N_12763);
xor U13806 (N_13806,N_12675,N_12476);
and U13807 (N_13807,N_12771,N_12751);
or U13808 (N_13808,N_12741,N_12576);
or U13809 (N_13809,N_12583,N_12644);
or U13810 (N_13810,N_12408,N_12805);
or U13811 (N_13811,N_12742,N_12012);
nor U13812 (N_13812,N_12384,N_12472);
and U13813 (N_13813,N_12917,N_12216);
or U13814 (N_13814,N_12338,N_12399);
or U13815 (N_13815,N_12979,N_12250);
nand U13816 (N_13816,N_12258,N_12850);
nand U13817 (N_13817,N_12724,N_12704);
xor U13818 (N_13818,N_12631,N_12646);
nor U13819 (N_13819,N_12790,N_12091);
xnor U13820 (N_13820,N_12910,N_12608);
or U13821 (N_13821,N_12334,N_12142);
and U13822 (N_13822,N_12069,N_12672);
xnor U13823 (N_13823,N_12589,N_12378);
and U13824 (N_13824,N_12351,N_12994);
xnor U13825 (N_13825,N_12189,N_12269);
or U13826 (N_13826,N_12614,N_12555);
nor U13827 (N_13827,N_12847,N_12092);
nand U13828 (N_13828,N_12919,N_12468);
nand U13829 (N_13829,N_12268,N_12406);
and U13830 (N_13830,N_12260,N_12006);
and U13831 (N_13831,N_12934,N_12391);
xnor U13832 (N_13832,N_12512,N_12590);
xor U13833 (N_13833,N_12043,N_12536);
xor U13834 (N_13834,N_12109,N_12494);
or U13835 (N_13835,N_12145,N_12613);
nor U13836 (N_13836,N_12995,N_12747);
xnor U13837 (N_13837,N_12566,N_12889);
or U13838 (N_13838,N_12221,N_12165);
or U13839 (N_13839,N_12153,N_12879);
and U13840 (N_13840,N_12951,N_12767);
xnor U13841 (N_13841,N_12502,N_12206);
or U13842 (N_13842,N_12949,N_12995);
nand U13843 (N_13843,N_12455,N_12333);
xnor U13844 (N_13844,N_12044,N_12393);
nor U13845 (N_13845,N_12793,N_12762);
nor U13846 (N_13846,N_12909,N_12865);
or U13847 (N_13847,N_12917,N_12353);
xnor U13848 (N_13848,N_12199,N_12071);
nand U13849 (N_13849,N_12255,N_12436);
or U13850 (N_13850,N_12480,N_12778);
xnor U13851 (N_13851,N_12339,N_12375);
nor U13852 (N_13852,N_12606,N_12852);
nor U13853 (N_13853,N_12878,N_12780);
or U13854 (N_13854,N_12096,N_12194);
and U13855 (N_13855,N_12663,N_12267);
nor U13856 (N_13856,N_12625,N_12601);
xor U13857 (N_13857,N_12741,N_12187);
and U13858 (N_13858,N_12891,N_12115);
nand U13859 (N_13859,N_12542,N_12610);
nand U13860 (N_13860,N_12207,N_12885);
xnor U13861 (N_13861,N_12848,N_12824);
nor U13862 (N_13862,N_12184,N_12587);
and U13863 (N_13863,N_12057,N_12977);
nand U13864 (N_13864,N_12287,N_12085);
and U13865 (N_13865,N_12456,N_12252);
nor U13866 (N_13866,N_12791,N_12477);
nand U13867 (N_13867,N_12398,N_12905);
nor U13868 (N_13868,N_12256,N_12509);
and U13869 (N_13869,N_12006,N_12593);
xnor U13870 (N_13870,N_12612,N_12471);
nor U13871 (N_13871,N_12567,N_12090);
xor U13872 (N_13872,N_12803,N_12876);
or U13873 (N_13873,N_12919,N_12817);
xor U13874 (N_13874,N_12212,N_12583);
or U13875 (N_13875,N_12990,N_12356);
nor U13876 (N_13876,N_12848,N_12620);
xnor U13877 (N_13877,N_12459,N_12467);
xor U13878 (N_13878,N_12928,N_12231);
xor U13879 (N_13879,N_12823,N_12817);
nand U13880 (N_13880,N_12918,N_12232);
nor U13881 (N_13881,N_12502,N_12191);
nand U13882 (N_13882,N_12588,N_12446);
nor U13883 (N_13883,N_12728,N_12799);
nand U13884 (N_13884,N_12301,N_12111);
nand U13885 (N_13885,N_12975,N_12035);
or U13886 (N_13886,N_12172,N_12704);
and U13887 (N_13887,N_12526,N_12819);
or U13888 (N_13888,N_12542,N_12411);
nor U13889 (N_13889,N_12064,N_12523);
or U13890 (N_13890,N_12940,N_12545);
nand U13891 (N_13891,N_12985,N_12721);
xor U13892 (N_13892,N_12574,N_12517);
nor U13893 (N_13893,N_12421,N_12177);
nand U13894 (N_13894,N_12219,N_12109);
and U13895 (N_13895,N_12048,N_12175);
nand U13896 (N_13896,N_12281,N_12535);
xnor U13897 (N_13897,N_12642,N_12370);
or U13898 (N_13898,N_12564,N_12085);
or U13899 (N_13899,N_12647,N_12216);
nand U13900 (N_13900,N_12526,N_12684);
nor U13901 (N_13901,N_12017,N_12688);
xnor U13902 (N_13902,N_12406,N_12711);
xnor U13903 (N_13903,N_12939,N_12314);
and U13904 (N_13904,N_12384,N_12030);
nor U13905 (N_13905,N_12770,N_12136);
nor U13906 (N_13906,N_12196,N_12790);
or U13907 (N_13907,N_12929,N_12899);
nor U13908 (N_13908,N_12220,N_12922);
xor U13909 (N_13909,N_12773,N_12675);
xor U13910 (N_13910,N_12508,N_12183);
xnor U13911 (N_13911,N_12369,N_12165);
xor U13912 (N_13912,N_12369,N_12681);
nand U13913 (N_13913,N_12473,N_12544);
nor U13914 (N_13914,N_12674,N_12428);
nor U13915 (N_13915,N_12217,N_12192);
nand U13916 (N_13916,N_12994,N_12756);
xnor U13917 (N_13917,N_12023,N_12914);
and U13918 (N_13918,N_12955,N_12254);
nand U13919 (N_13919,N_12703,N_12077);
and U13920 (N_13920,N_12441,N_12230);
nand U13921 (N_13921,N_12195,N_12414);
nand U13922 (N_13922,N_12728,N_12977);
nor U13923 (N_13923,N_12582,N_12187);
or U13924 (N_13924,N_12795,N_12831);
nand U13925 (N_13925,N_12511,N_12956);
xnor U13926 (N_13926,N_12151,N_12089);
or U13927 (N_13927,N_12649,N_12427);
or U13928 (N_13928,N_12460,N_12787);
xor U13929 (N_13929,N_12883,N_12845);
nor U13930 (N_13930,N_12906,N_12570);
and U13931 (N_13931,N_12746,N_12664);
and U13932 (N_13932,N_12698,N_12450);
xor U13933 (N_13933,N_12267,N_12755);
nor U13934 (N_13934,N_12346,N_12163);
and U13935 (N_13935,N_12515,N_12541);
xor U13936 (N_13936,N_12221,N_12189);
or U13937 (N_13937,N_12492,N_12709);
nor U13938 (N_13938,N_12271,N_12584);
nand U13939 (N_13939,N_12145,N_12826);
nand U13940 (N_13940,N_12259,N_12109);
and U13941 (N_13941,N_12225,N_12686);
nand U13942 (N_13942,N_12537,N_12010);
and U13943 (N_13943,N_12704,N_12046);
and U13944 (N_13944,N_12179,N_12275);
nor U13945 (N_13945,N_12911,N_12901);
nand U13946 (N_13946,N_12198,N_12097);
nand U13947 (N_13947,N_12338,N_12598);
or U13948 (N_13948,N_12663,N_12953);
nand U13949 (N_13949,N_12673,N_12457);
and U13950 (N_13950,N_12559,N_12119);
nand U13951 (N_13951,N_12002,N_12386);
xnor U13952 (N_13952,N_12735,N_12088);
nand U13953 (N_13953,N_12789,N_12366);
or U13954 (N_13954,N_12940,N_12289);
and U13955 (N_13955,N_12811,N_12694);
nand U13956 (N_13956,N_12469,N_12023);
nor U13957 (N_13957,N_12765,N_12198);
and U13958 (N_13958,N_12639,N_12422);
and U13959 (N_13959,N_12013,N_12578);
nand U13960 (N_13960,N_12115,N_12182);
nor U13961 (N_13961,N_12932,N_12939);
nor U13962 (N_13962,N_12189,N_12428);
nand U13963 (N_13963,N_12255,N_12626);
nor U13964 (N_13964,N_12529,N_12911);
nand U13965 (N_13965,N_12467,N_12461);
xnor U13966 (N_13966,N_12113,N_12554);
xor U13967 (N_13967,N_12086,N_12640);
or U13968 (N_13968,N_12016,N_12191);
xor U13969 (N_13969,N_12936,N_12588);
nor U13970 (N_13970,N_12248,N_12836);
nor U13971 (N_13971,N_12154,N_12341);
or U13972 (N_13972,N_12128,N_12751);
nor U13973 (N_13973,N_12273,N_12950);
xor U13974 (N_13974,N_12878,N_12352);
xnor U13975 (N_13975,N_12376,N_12711);
or U13976 (N_13976,N_12299,N_12896);
nand U13977 (N_13977,N_12552,N_12804);
or U13978 (N_13978,N_12091,N_12742);
nand U13979 (N_13979,N_12100,N_12395);
or U13980 (N_13980,N_12551,N_12064);
xor U13981 (N_13981,N_12016,N_12139);
nand U13982 (N_13982,N_12394,N_12562);
or U13983 (N_13983,N_12487,N_12675);
nand U13984 (N_13984,N_12262,N_12645);
or U13985 (N_13985,N_12505,N_12594);
and U13986 (N_13986,N_12299,N_12932);
nand U13987 (N_13987,N_12900,N_12366);
xnor U13988 (N_13988,N_12205,N_12776);
or U13989 (N_13989,N_12544,N_12102);
nor U13990 (N_13990,N_12754,N_12338);
and U13991 (N_13991,N_12251,N_12704);
nor U13992 (N_13992,N_12691,N_12810);
or U13993 (N_13993,N_12261,N_12598);
nor U13994 (N_13994,N_12284,N_12755);
nor U13995 (N_13995,N_12439,N_12519);
nor U13996 (N_13996,N_12032,N_12073);
xnor U13997 (N_13997,N_12490,N_12187);
nor U13998 (N_13998,N_12017,N_12200);
xor U13999 (N_13999,N_12076,N_12005);
or U14000 (N_14000,N_13181,N_13326);
or U14001 (N_14001,N_13586,N_13761);
xor U14002 (N_14002,N_13697,N_13995);
nor U14003 (N_14003,N_13526,N_13513);
and U14004 (N_14004,N_13100,N_13113);
nand U14005 (N_14005,N_13422,N_13267);
xnor U14006 (N_14006,N_13082,N_13673);
xor U14007 (N_14007,N_13200,N_13774);
and U14008 (N_14008,N_13150,N_13911);
xnor U14009 (N_14009,N_13579,N_13373);
nor U14010 (N_14010,N_13202,N_13437);
nor U14011 (N_14011,N_13295,N_13313);
nand U14012 (N_14012,N_13936,N_13155);
xor U14013 (N_14013,N_13432,N_13890);
nor U14014 (N_14014,N_13368,N_13271);
nand U14015 (N_14015,N_13087,N_13490);
or U14016 (N_14016,N_13751,N_13947);
xor U14017 (N_14017,N_13042,N_13979);
xnor U14018 (N_14018,N_13694,N_13862);
nand U14019 (N_14019,N_13552,N_13131);
nand U14020 (N_14020,N_13211,N_13341);
nor U14021 (N_14021,N_13493,N_13417);
or U14022 (N_14022,N_13978,N_13532);
and U14023 (N_14023,N_13980,N_13838);
or U14024 (N_14024,N_13455,N_13550);
xnor U14025 (N_14025,N_13201,N_13576);
and U14026 (N_14026,N_13057,N_13010);
or U14027 (N_14027,N_13677,N_13463);
nand U14028 (N_14028,N_13725,N_13356);
xor U14029 (N_14029,N_13991,N_13452);
or U14030 (N_14030,N_13842,N_13050);
xor U14031 (N_14031,N_13606,N_13310);
nand U14032 (N_14032,N_13036,N_13334);
nand U14033 (N_14033,N_13291,N_13610);
or U14034 (N_14034,N_13811,N_13982);
and U14035 (N_14035,N_13145,N_13702);
nor U14036 (N_14036,N_13955,N_13758);
nand U14037 (N_14037,N_13912,N_13617);
nor U14038 (N_14038,N_13435,N_13235);
or U14039 (N_14039,N_13301,N_13512);
xnor U14040 (N_14040,N_13296,N_13534);
or U14041 (N_14041,N_13255,N_13439);
nand U14042 (N_14042,N_13132,N_13571);
and U14043 (N_14043,N_13340,N_13221);
or U14044 (N_14044,N_13247,N_13360);
nor U14045 (N_14045,N_13799,N_13025);
nand U14046 (N_14046,N_13674,N_13961);
nand U14047 (N_14047,N_13063,N_13404);
xnor U14048 (N_14048,N_13733,N_13342);
nor U14049 (N_14049,N_13119,N_13768);
xor U14050 (N_14050,N_13027,N_13167);
nor U14051 (N_14051,N_13693,N_13314);
nand U14052 (N_14052,N_13399,N_13861);
xor U14053 (N_14053,N_13248,N_13661);
xor U14054 (N_14054,N_13092,N_13485);
and U14055 (N_14055,N_13782,N_13074);
and U14056 (N_14056,N_13017,N_13644);
nand U14057 (N_14057,N_13350,N_13400);
xor U14058 (N_14058,N_13277,N_13604);
xnor U14059 (N_14059,N_13195,N_13937);
and U14060 (N_14060,N_13450,N_13877);
nand U14061 (N_14061,N_13946,N_13690);
nor U14062 (N_14062,N_13773,N_13070);
nor U14063 (N_14063,N_13517,N_13016);
nand U14064 (N_14064,N_13728,N_13664);
or U14065 (N_14065,N_13871,N_13727);
nor U14066 (N_14066,N_13065,N_13323);
and U14067 (N_14067,N_13335,N_13832);
nand U14068 (N_14068,N_13405,N_13919);
nand U14069 (N_14069,N_13032,N_13581);
nand U14070 (N_14070,N_13207,N_13444);
nand U14071 (N_14071,N_13574,N_13709);
nor U14072 (N_14072,N_13086,N_13851);
or U14073 (N_14073,N_13352,N_13764);
nor U14074 (N_14074,N_13898,N_13654);
or U14075 (N_14075,N_13069,N_13907);
and U14076 (N_14076,N_13110,N_13044);
or U14077 (N_14077,N_13480,N_13481);
xnor U14078 (N_14078,N_13218,N_13021);
and U14079 (N_14079,N_13177,N_13308);
xnor U14080 (N_14080,N_13064,N_13459);
and U14081 (N_14081,N_13000,N_13943);
or U14082 (N_14082,N_13007,N_13881);
nand U14083 (N_14083,N_13749,N_13988);
nor U14084 (N_14084,N_13284,N_13484);
nand U14085 (N_14085,N_13942,N_13495);
or U14086 (N_14086,N_13037,N_13864);
and U14087 (N_14087,N_13114,N_13243);
xnor U14088 (N_14088,N_13795,N_13105);
and U14089 (N_14089,N_13977,N_13168);
or U14090 (N_14090,N_13927,N_13873);
nand U14091 (N_14091,N_13544,N_13591);
nand U14092 (N_14092,N_13797,N_13822);
nor U14093 (N_14093,N_13511,N_13306);
xor U14094 (N_14094,N_13077,N_13788);
or U14095 (N_14095,N_13231,N_13887);
and U14096 (N_14096,N_13396,N_13724);
or U14097 (N_14097,N_13297,N_13361);
and U14098 (N_14098,N_13962,N_13164);
nand U14099 (N_14099,N_13228,N_13078);
nor U14100 (N_14100,N_13425,N_13895);
and U14101 (N_14101,N_13847,N_13353);
nand U14102 (N_14102,N_13573,N_13712);
and U14103 (N_14103,N_13940,N_13142);
or U14104 (N_14104,N_13753,N_13095);
or U14105 (N_14105,N_13566,N_13117);
and U14106 (N_14106,N_13288,N_13473);
xor U14107 (N_14107,N_13115,N_13424);
or U14108 (N_14108,N_13222,N_13789);
nand U14109 (N_14109,N_13096,N_13685);
or U14110 (N_14110,N_13865,N_13680);
and U14111 (N_14111,N_13794,N_13650);
or U14112 (N_14112,N_13054,N_13190);
xnor U14113 (N_14113,N_13060,N_13626);
and U14114 (N_14114,N_13780,N_13302);
and U14115 (N_14115,N_13798,N_13196);
or U14116 (N_14116,N_13382,N_13398);
xnor U14117 (N_14117,N_13224,N_13347);
xor U14118 (N_14118,N_13333,N_13939);
nor U14119 (N_14119,N_13236,N_13623);
nand U14120 (N_14120,N_13922,N_13790);
nor U14121 (N_14121,N_13850,N_13910);
nand U14122 (N_14122,N_13009,N_13125);
or U14123 (N_14123,N_13406,N_13648);
and U14124 (N_14124,N_13309,N_13545);
or U14125 (N_14125,N_13281,N_13730);
xor U14126 (N_14126,N_13003,N_13250);
and U14127 (N_14127,N_13537,N_13427);
or U14128 (N_14128,N_13602,N_13233);
nor U14129 (N_14129,N_13215,N_13769);
xor U14130 (N_14130,N_13853,N_13682);
and U14131 (N_14131,N_13796,N_13641);
or U14132 (N_14132,N_13583,N_13921);
xor U14133 (N_14133,N_13428,N_13263);
xor U14134 (N_14134,N_13020,N_13594);
or U14135 (N_14135,N_13713,N_13558);
nor U14136 (N_14136,N_13061,N_13950);
nand U14137 (N_14137,N_13152,N_13525);
and U14138 (N_14138,N_13553,N_13038);
and U14139 (N_14139,N_13635,N_13521);
nand U14140 (N_14140,N_13578,N_13963);
nor U14141 (N_14141,N_13676,N_13934);
nand U14142 (N_14142,N_13646,N_13671);
or U14143 (N_14143,N_13029,N_13944);
nor U14144 (N_14144,N_13374,N_13959);
xor U14145 (N_14145,N_13567,N_13073);
or U14146 (N_14146,N_13966,N_13516);
nand U14147 (N_14147,N_13539,N_13123);
nor U14148 (N_14148,N_13157,N_13869);
and U14149 (N_14149,N_13212,N_13144);
xor U14150 (N_14150,N_13148,N_13475);
or U14151 (N_14151,N_13540,N_13529);
and U14152 (N_14152,N_13464,N_13863);
or U14153 (N_14153,N_13121,N_13371);
or U14154 (N_14154,N_13343,N_13412);
and U14155 (N_14155,N_13531,N_13756);
or U14156 (N_14156,N_13740,N_13739);
or U14157 (N_14157,N_13787,N_13651);
nand U14158 (N_14158,N_13194,N_13182);
and U14159 (N_14159,N_13376,N_13729);
or U14160 (N_14160,N_13820,N_13320);
xnor U14161 (N_14161,N_13443,N_13018);
nand U14162 (N_14162,N_13462,N_13603);
and U14163 (N_14163,N_13741,N_13191);
and U14164 (N_14164,N_13708,N_13745);
nor U14165 (N_14165,N_13908,N_13059);
nand U14166 (N_14166,N_13486,N_13246);
xor U14167 (N_14167,N_13278,N_13561);
and U14168 (N_14168,N_13325,N_13099);
xnor U14169 (N_14169,N_13408,N_13718);
nor U14170 (N_14170,N_13330,N_13755);
xnor U14171 (N_14171,N_13109,N_13754);
nor U14172 (N_14172,N_13965,N_13023);
and U14173 (N_14173,N_13008,N_13319);
or U14174 (N_14174,N_13924,N_13434);
or U14175 (N_14175,N_13011,N_13839);
xnor U14176 (N_14176,N_13595,N_13687);
and U14177 (N_14177,N_13828,N_13533);
and U14178 (N_14178,N_13589,N_13714);
xor U14179 (N_14179,N_13090,N_13914);
and U14180 (N_14180,N_13732,N_13500);
nor U14181 (N_14181,N_13389,N_13262);
nand U14182 (N_14182,N_13226,N_13506);
nand U14183 (N_14183,N_13630,N_13487);
xor U14184 (N_14184,N_13520,N_13840);
nand U14185 (N_14185,N_13106,N_13994);
xor U14186 (N_14186,N_13476,N_13094);
and U14187 (N_14187,N_13655,N_13104);
or U14188 (N_14188,N_13835,N_13688);
nand U14189 (N_14189,N_13193,N_13625);
and U14190 (N_14190,N_13458,N_13638);
and U14191 (N_14191,N_13891,N_13438);
and U14192 (N_14192,N_13888,N_13624);
or U14193 (N_14193,N_13577,N_13375);
nand U14194 (N_14194,N_13139,N_13809);
nand U14195 (N_14195,N_13261,N_13770);
xor U14196 (N_14196,N_13156,N_13945);
and U14197 (N_14197,N_13679,N_13442);
nor U14198 (N_14198,N_13479,N_13598);
nor U14199 (N_14199,N_13418,N_13609);
xnor U14200 (N_14200,N_13205,N_13771);
xor U14201 (N_14201,N_13785,N_13383);
xor U14202 (N_14202,N_13904,N_13543);
nand U14203 (N_14203,N_13477,N_13746);
nand U14204 (N_14204,N_13546,N_13868);
xnor U14205 (N_14205,N_13670,N_13711);
nor U14206 (N_14206,N_13784,N_13209);
and U14207 (N_14207,N_13781,N_13006);
nor U14208 (N_14208,N_13762,N_13524);
or U14209 (N_14209,N_13700,N_13245);
and U14210 (N_14210,N_13127,N_13830);
nor U14211 (N_14211,N_13146,N_13413);
and U14212 (N_14212,N_13564,N_13457);
nor U14213 (N_14213,N_13289,N_13518);
xor U14214 (N_14214,N_13403,N_13509);
xor U14215 (N_14215,N_13112,N_13456);
nor U14216 (N_14216,N_13362,N_13560);
xnor U14217 (N_14217,N_13071,N_13143);
nand U14218 (N_14218,N_13667,N_13683);
or U14219 (N_14219,N_13556,N_13256);
and U14220 (N_14220,N_13752,N_13372);
xor U14221 (N_14221,N_13897,N_13660);
or U14222 (N_14222,N_13478,N_13266);
and U14223 (N_14223,N_13615,N_13258);
xor U14224 (N_14224,N_13831,N_13040);
nor U14225 (N_14225,N_13004,N_13097);
or U14226 (N_14226,N_13715,N_13311);
or U14227 (N_14227,N_13453,N_13147);
nand U14228 (N_14228,N_13197,N_13590);
and U14229 (N_14229,N_13187,N_13707);
and U14230 (N_14230,N_13721,N_13068);
and U14231 (N_14231,N_13259,N_13367);
and U14232 (N_14232,N_13045,N_13203);
xnor U14233 (N_14233,N_13244,N_13241);
or U14234 (N_14234,N_13351,N_13293);
and U14235 (N_14235,N_13274,N_13158);
xor U14236 (N_14236,N_13766,N_13703);
nand U14237 (N_14237,N_13938,N_13019);
or U14238 (N_14238,N_13080,N_13468);
nor U14239 (N_14239,N_13920,N_13970);
nor U14240 (N_14240,N_13916,N_13565);
xnor U14241 (N_14241,N_13185,N_13821);
nand U14242 (N_14242,N_13159,N_13307);
or U14243 (N_14243,N_13491,N_13093);
or U14244 (N_14244,N_13569,N_13841);
nand U14245 (N_14245,N_13161,N_13804);
nand U14246 (N_14246,N_13254,N_13969);
nor U14247 (N_14247,N_13759,N_13137);
and U14248 (N_14248,N_13562,N_13572);
nor U14249 (N_14249,N_13391,N_13836);
and U14250 (N_14250,N_13812,N_13964);
or U14251 (N_14251,N_13691,N_13731);
and U14252 (N_14252,N_13772,N_13716);
nand U14253 (N_14253,N_13409,N_13318);
or U14254 (N_14254,N_13393,N_13555);
nand U14255 (N_14255,N_13359,N_13767);
nand U14256 (N_14256,N_13033,N_13878);
xor U14257 (N_14257,N_13217,N_13906);
or U14258 (N_14258,N_13672,N_13696);
or U14259 (N_14259,N_13166,N_13722);
nor U14260 (N_14260,N_13172,N_13275);
nand U14261 (N_14261,N_13055,N_13686);
or U14262 (N_14262,N_13570,N_13743);
or U14263 (N_14263,N_13299,N_13014);
nor U14264 (N_14264,N_13681,N_13260);
nand U14265 (N_14265,N_13067,N_13501);
nand U14266 (N_14266,N_13760,N_13706);
xnor U14267 (N_14267,N_13058,N_13303);
and U14268 (N_14268,N_13684,N_13678);
xor U14269 (N_14269,N_13859,N_13381);
or U14270 (N_14270,N_13536,N_13300);
xor U14271 (N_14271,N_13173,N_13649);
nand U14272 (N_14272,N_13883,N_13926);
nor U14273 (N_14273,N_13996,N_13206);
nor U14274 (N_14274,N_13363,N_13129);
nand U14275 (N_14275,N_13441,N_13637);
nor U14276 (N_14276,N_13857,N_13502);
xnor U14277 (N_14277,N_13659,N_13229);
nand U14278 (N_14278,N_13792,N_13802);
or U14279 (N_14279,N_13631,N_13584);
and U14280 (N_14280,N_13507,N_13251);
nand U14281 (N_14281,N_13102,N_13328);
and U14282 (N_14282,N_13286,N_13332);
and U14283 (N_14283,N_13541,N_13429);
nand U14284 (N_14284,N_13163,N_13647);
xor U14285 (N_14285,N_13879,N_13188);
or U14286 (N_14286,N_13433,N_13198);
or U14287 (N_14287,N_13726,N_13582);
nand U14288 (N_14288,N_13813,N_13607);
nor U14289 (N_14289,N_13913,N_13636);
nor U14290 (N_14290,N_13046,N_13527);
xor U14291 (N_14291,N_13614,N_13817);
nand U14292 (N_14292,N_13701,N_13975);
nor U14293 (N_14293,N_13514,N_13952);
and U14294 (N_14294,N_13178,N_13953);
nor U14295 (N_14295,N_13416,N_13049);
nand U14296 (N_14296,N_13750,N_13385);
nor U14297 (N_14297,N_13689,N_13549);
nand U14298 (N_14298,N_13355,N_13776);
xnor U14299 (N_14299,N_13596,N_13987);
or U14300 (N_14300,N_13431,N_13508);
or U14301 (N_14301,N_13948,N_13339);
or U14302 (N_14302,N_13053,N_13162);
nand U14303 (N_14303,N_13345,N_13130);
nor U14304 (N_14304,N_13580,N_13327);
xor U14305 (N_14305,N_13470,N_13949);
or U14306 (N_14306,N_13354,N_13223);
and U14307 (N_14307,N_13902,N_13783);
or U14308 (N_14308,N_13960,N_13778);
xnor U14309 (N_14309,N_13107,N_13472);
or U14310 (N_14310,N_13808,N_13829);
nor U14311 (N_14311,N_13272,N_13918);
nor U14312 (N_14312,N_13632,N_13084);
nor U14313 (N_14313,N_13814,N_13738);
or U14314 (N_14314,N_13930,N_13925);
xor U14315 (N_14315,N_13825,N_13022);
and U14316 (N_14316,N_13621,N_13257);
nand U14317 (N_14317,N_13242,N_13232);
and U14318 (N_14318,N_13662,N_13585);
xnor U14319 (N_14319,N_13668,N_13387);
and U14320 (N_14320,N_13079,N_13081);
nand U14321 (N_14321,N_13496,N_13454);
or U14322 (N_14322,N_13805,N_13349);
and U14323 (N_14323,N_13298,N_13154);
or U14324 (N_14324,N_13174,N_13051);
and U14325 (N_14325,N_13357,N_13826);
or U14326 (N_14326,N_13968,N_13557);
nor U14327 (N_14327,N_13645,N_13083);
or U14328 (N_14328,N_13886,N_13030);
xor U14329 (N_14329,N_13214,N_13620);
nor U14330 (N_14330,N_13034,N_13896);
nor U14331 (N_14331,N_13108,N_13024);
nand U14332 (N_14332,N_13467,N_13929);
xor U14333 (N_14333,N_13504,N_13465);
nand U14334 (N_14334,N_13220,N_13043);
and U14335 (N_14335,N_13860,N_13613);
and U14336 (N_14336,N_13931,N_13954);
nand U14337 (N_14337,N_13336,N_13331);
and U14338 (N_14338,N_13515,N_13884);
xor U14339 (N_14339,N_13551,N_13199);
or U14340 (N_14340,N_13779,N_13559);
nor U14341 (N_14341,N_13253,N_13149);
nor U14342 (N_14342,N_13482,N_13449);
nand U14343 (N_14343,N_13627,N_13249);
nor U14344 (N_14344,N_13324,N_13337);
xor U14345 (N_14345,N_13366,N_13415);
and U14346 (N_14346,N_13528,N_13270);
nand U14347 (N_14347,N_13338,N_13775);
xnor U14348 (N_14348,N_13628,N_13608);
nand U14349 (N_14349,N_13547,N_13999);
nand U14350 (N_14350,N_13204,N_13171);
nand U14351 (N_14351,N_13698,N_13039);
or U14352 (N_14352,N_13901,N_13136);
xnor U14353 (N_14353,N_13041,N_13675);
xor U14354 (N_14354,N_13234,N_13225);
nor U14355 (N_14355,N_13189,N_13282);
xnor U14356 (N_14356,N_13138,N_13269);
nor U14357 (N_14357,N_13981,N_13322);
xor U14358 (N_14358,N_13986,N_13855);
xor U14359 (N_14359,N_13348,N_13592);
nor U14360 (N_14360,N_13984,N_13088);
or U14361 (N_14361,N_13469,N_13587);
nand U14362 (N_14362,N_13846,N_13395);
nor U14363 (N_14363,N_13013,N_13239);
nor U14364 (N_14364,N_13134,N_13522);
nand U14365 (N_14365,N_13252,N_13892);
or U14366 (N_14366,N_13317,N_13219);
xnor U14367 (N_14367,N_13880,N_13186);
xor U14368 (N_14368,N_13292,N_13806);
or U14369 (N_14369,N_13990,N_13498);
and U14370 (N_14370,N_13656,N_13710);
xor U14371 (N_14371,N_13238,N_13923);
xnor U14372 (N_14372,N_13141,N_13066);
nor U14373 (N_14373,N_13748,N_13101);
xor U14374 (N_14374,N_13447,N_13548);
xor U14375 (N_14375,N_13510,N_13365);
or U14376 (N_14376,N_13705,N_13414);
or U14377 (N_14377,N_13992,N_13663);
xor U14378 (N_14378,N_13622,N_13227);
nand U14379 (N_14379,N_13494,N_13128);
or U14380 (N_14380,N_13793,N_13801);
nand U14381 (N_14381,N_13133,N_13419);
nor U14382 (N_14382,N_13720,N_13026);
nor U14383 (N_14383,N_13184,N_13619);
xnor U14384 (N_14384,N_13983,N_13126);
nand U14385 (N_14385,N_13140,N_13974);
nand U14386 (N_14386,N_13344,N_13237);
xnor U14387 (N_14387,N_13072,N_13423);
or U14388 (N_14388,N_13734,N_13653);
or U14389 (N_14389,N_13287,N_13001);
and U14390 (N_14390,N_13380,N_13563);
nand U14391 (N_14391,N_13390,N_13736);
nand U14392 (N_14392,N_13815,N_13047);
and U14393 (N_14393,N_13165,N_13633);
nor U14394 (N_14394,N_13876,N_13179);
or U14395 (N_14395,N_13791,N_13666);
nand U14396 (N_14396,N_13276,N_13503);
and U14397 (N_14397,N_13120,N_13213);
nor U14398 (N_14398,N_13377,N_13461);
xor U14399 (N_14399,N_13305,N_13160);
nand U14400 (N_14400,N_13210,N_13176);
nand U14401 (N_14401,N_13695,N_13180);
nand U14402 (N_14402,N_13699,N_13285);
xor U14403 (N_14403,N_13757,N_13854);
nand U14404 (N_14404,N_13958,N_13056);
nor U14405 (N_14405,N_13849,N_13364);
xnor U14406 (N_14406,N_13279,N_13170);
or U14407 (N_14407,N_13091,N_13446);
xnor U14408 (N_14408,N_13917,N_13379);
nor U14409 (N_14409,N_13998,N_13872);
xnor U14410 (N_14410,N_13971,N_13411);
or U14411 (N_14411,N_13858,N_13903);
and U14412 (N_14412,N_13489,N_13474);
and U14413 (N_14413,N_13230,N_13466);
nor U14414 (N_14414,N_13807,N_13002);
xor U14415 (N_14415,N_13597,N_13240);
xor U14416 (N_14416,N_13599,N_13265);
and U14417 (N_14417,N_13273,N_13600);
nand U14418 (N_14418,N_13283,N_13397);
xnor U14419 (N_14419,N_13175,N_13492);
and U14420 (N_14420,N_13483,N_13005);
xor U14421 (N_14421,N_13436,N_13048);
and U14422 (N_14422,N_13642,N_13401);
nand U14423 (N_14423,N_13652,N_13658);
xor U14424 (N_14424,N_13856,N_13629);
nand U14425 (N_14425,N_13593,N_13744);
and U14426 (N_14426,N_13723,N_13098);
nor U14427 (N_14427,N_13889,N_13928);
xor U14428 (N_14428,N_13505,N_13394);
and U14429 (N_14429,N_13208,N_13900);
nor U14430 (N_14430,N_13800,N_13392);
and U14431 (N_14431,N_13665,N_13407);
or U14432 (N_14432,N_13870,N_13116);
nand U14433 (N_14433,N_13618,N_13616);
nor U14434 (N_14434,N_13899,N_13384);
nand U14435 (N_14435,N_13315,N_13894);
and U14436 (N_14436,N_13031,N_13704);
xnor U14437 (N_14437,N_13530,N_13803);
or U14438 (N_14438,N_13135,N_13216);
nor U14439 (N_14439,N_13692,N_13818);
xnor U14440 (N_14440,N_13369,N_13845);
nand U14441 (N_14441,N_13378,N_13440);
xor U14442 (N_14442,N_13993,N_13909);
nand U14443 (N_14443,N_13089,N_13833);
or U14444 (N_14444,N_13951,N_13568);
nand U14445 (N_14445,N_13497,N_13410);
nor U14446 (N_14446,N_13012,N_13386);
or U14447 (N_14447,N_13941,N_13915);
and U14448 (N_14448,N_13151,N_13777);
or U14449 (N_14449,N_13471,N_13304);
or U14450 (N_14450,N_13169,N_13765);
nand U14451 (N_14451,N_13823,N_13448);
or U14452 (N_14452,N_13810,N_13657);
or U14453 (N_14453,N_13280,N_13290);
nand U14454 (N_14454,N_13819,N_13601);
nand U14455 (N_14455,N_13640,N_13848);
and U14456 (N_14456,N_13735,N_13153);
and U14457 (N_14457,N_13866,N_13316);
or U14458 (N_14458,N_13329,N_13827);
or U14459 (N_14459,N_13643,N_13192);
or U14460 (N_14460,N_13426,N_13972);
nor U14461 (N_14461,N_13956,N_13062);
or U14462 (N_14462,N_13997,N_13111);
nand U14463 (N_14463,N_13076,N_13358);
and U14464 (N_14464,N_13575,N_13015);
and U14465 (N_14465,N_13388,N_13882);
nor U14466 (N_14466,N_13763,N_13183);
xor U14467 (N_14467,N_13852,N_13035);
and U14468 (N_14468,N_13028,N_13634);
xor U14469 (N_14469,N_13294,N_13430);
nand U14470 (N_14470,N_13445,N_13538);
xor U14471 (N_14471,N_13421,N_13118);
xnor U14472 (N_14472,N_13837,N_13554);
or U14473 (N_14473,N_13321,N_13719);
nor U14474 (N_14474,N_13523,N_13122);
xor U14475 (N_14475,N_13885,N_13935);
nand U14476 (N_14476,N_13893,N_13933);
and U14477 (N_14477,N_13264,N_13967);
and U14478 (N_14478,N_13612,N_13075);
xor U14479 (N_14479,N_13957,N_13268);
xor U14480 (N_14480,N_13843,N_13085);
nand U14481 (N_14481,N_13844,N_13905);
nand U14482 (N_14482,N_13312,N_13605);
and U14483 (N_14483,N_13499,N_13976);
and U14484 (N_14484,N_13989,N_13985);
and U14485 (N_14485,N_13420,N_13973);
nor U14486 (N_14486,N_13535,N_13816);
and U14487 (N_14487,N_13542,N_13932);
and U14488 (N_14488,N_13588,N_13747);
and U14489 (N_14489,N_13737,N_13451);
nand U14490 (N_14490,N_13717,N_13874);
and U14491 (N_14491,N_13867,N_13346);
nand U14492 (N_14492,N_13124,N_13460);
xor U14493 (N_14493,N_13639,N_13824);
nand U14494 (N_14494,N_13370,N_13103);
and U14495 (N_14495,N_13519,N_13786);
xor U14496 (N_14496,N_13669,N_13834);
nor U14497 (N_14497,N_13488,N_13402);
xnor U14498 (N_14498,N_13052,N_13875);
nand U14499 (N_14499,N_13742,N_13611);
nor U14500 (N_14500,N_13738,N_13157);
and U14501 (N_14501,N_13893,N_13730);
nand U14502 (N_14502,N_13379,N_13667);
xor U14503 (N_14503,N_13752,N_13700);
or U14504 (N_14504,N_13254,N_13121);
or U14505 (N_14505,N_13339,N_13763);
xnor U14506 (N_14506,N_13418,N_13779);
or U14507 (N_14507,N_13652,N_13969);
and U14508 (N_14508,N_13706,N_13798);
and U14509 (N_14509,N_13775,N_13726);
nor U14510 (N_14510,N_13832,N_13595);
nor U14511 (N_14511,N_13241,N_13630);
and U14512 (N_14512,N_13883,N_13932);
nor U14513 (N_14513,N_13778,N_13354);
xor U14514 (N_14514,N_13679,N_13993);
nor U14515 (N_14515,N_13404,N_13595);
or U14516 (N_14516,N_13171,N_13243);
xor U14517 (N_14517,N_13228,N_13793);
xor U14518 (N_14518,N_13407,N_13477);
nor U14519 (N_14519,N_13795,N_13948);
or U14520 (N_14520,N_13289,N_13169);
or U14521 (N_14521,N_13308,N_13130);
or U14522 (N_14522,N_13311,N_13666);
or U14523 (N_14523,N_13979,N_13230);
and U14524 (N_14524,N_13173,N_13822);
nand U14525 (N_14525,N_13364,N_13857);
xor U14526 (N_14526,N_13515,N_13502);
nand U14527 (N_14527,N_13792,N_13510);
and U14528 (N_14528,N_13832,N_13010);
nor U14529 (N_14529,N_13158,N_13875);
xnor U14530 (N_14530,N_13177,N_13075);
and U14531 (N_14531,N_13114,N_13782);
nand U14532 (N_14532,N_13112,N_13549);
xnor U14533 (N_14533,N_13966,N_13852);
nor U14534 (N_14534,N_13187,N_13922);
nand U14535 (N_14535,N_13124,N_13476);
nand U14536 (N_14536,N_13830,N_13762);
nor U14537 (N_14537,N_13566,N_13798);
nor U14538 (N_14538,N_13255,N_13657);
nor U14539 (N_14539,N_13307,N_13267);
nand U14540 (N_14540,N_13095,N_13998);
nor U14541 (N_14541,N_13464,N_13317);
nand U14542 (N_14542,N_13247,N_13618);
nand U14543 (N_14543,N_13412,N_13623);
nor U14544 (N_14544,N_13695,N_13766);
or U14545 (N_14545,N_13195,N_13272);
or U14546 (N_14546,N_13108,N_13187);
nand U14547 (N_14547,N_13577,N_13676);
nand U14548 (N_14548,N_13196,N_13708);
and U14549 (N_14549,N_13751,N_13937);
nand U14550 (N_14550,N_13534,N_13636);
nor U14551 (N_14551,N_13560,N_13949);
and U14552 (N_14552,N_13346,N_13507);
xor U14553 (N_14553,N_13811,N_13444);
and U14554 (N_14554,N_13659,N_13936);
or U14555 (N_14555,N_13124,N_13569);
nor U14556 (N_14556,N_13615,N_13330);
nor U14557 (N_14557,N_13717,N_13418);
xnor U14558 (N_14558,N_13961,N_13660);
nand U14559 (N_14559,N_13018,N_13456);
or U14560 (N_14560,N_13052,N_13119);
and U14561 (N_14561,N_13871,N_13951);
xnor U14562 (N_14562,N_13571,N_13075);
nor U14563 (N_14563,N_13659,N_13089);
nand U14564 (N_14564,N_13948,N_13029);
nor U14565 (N_14565,N_13983,N_13139);
or U14566 (N_14566,N_13661,N_13551);
or U14567 (N_14567,N_13060,N_13024);
xor U14568 (N_14568,N_13445,N_13616);
and U14569 (N_14569,N_13928,N_13275);
nand U14570 (N_14570,N_13860,N_13229);
xnor U14571 (N_14571,N_13508,N_13595);
or U14572 (N_14572,N_13934,N_13261);
and U14573 (N_14573,N_13588,N_13420);
and U14574 (N_14574,N_13292,N_13608);
xnor U14575 (N_14575,N_13018,N_13447);
nand U14576 (N_14576,N_13858,N_13249);
or U14577 (N_14577,N_13997,N_13503);
nand U14578 (N_14578,N_13494,N_13569);
nor U14579 (N_14579,N_13952,N_13425);
nand U14580 (N_14580,N_13520,N_13625);
and U14581 (N_14581,N_13833,N_13129);
or U14582 (N_14582,N_13611,N_13236);
nor U14583 (N_14583,N_13130,N_13586);
and U14584 (N_14584,N_13722,N_13420);
nand U14585 (N_14585,N_13775,N_13875);
and U14586 (N_14586,N_13235,N_13064);
or U14587 (N_14587,N_13120,N_13745);
nor U14588 (N_14588,N_13677,N_13901);
xor U14589 (N_14589,N_13544,N_13235);
nor U14590 (N_14590,N_13807,N_13855);
and U14591 (N_14591,N_13933,N_13969);
xor U14592 (N_14592,N_13455,N_13742);
nor U14593 (N_14593,N_13260,N_13073);
and U14594 (N_14594,N_13261,N_13190);
or U14595 (N_14595,N_13678,N_13399);
or U14596 (N_14596,N_13551,N_13512);
xnor U14597 (N_14597,N_13840,N_13801);
nand U14598 (N_14598,N_13912,N_13883);
and U14599 (N_14599,N_13081,N_13808);
xnor U14600 (N_14600,N_13808,N_13405);
nand U14601 (N_14601,N_13441,N_13245);
xor U14602 (N_14602,N_13754,N_13287);
or U14603 (N_14603,N_13864,N_13807);
or U14604 (N_14604,N_13166,N_13665);
and U14605 (N_14605,N_13137,N_13929);
or U14606 (N_14606,N_13545,N_13373);
nor U14607 (N_14607,N_13064,N_13682);
nor U14608 (N_14608,N_13432,N_13748);
and U14609 (N_14609,N_13990,N_13775);
or U14610 (N_14610,N_13971,N_13181);
nand U14611 (N_14611,N_13646,N_13475);
and U14612 (N_14612,N_13065,N_13249);
and U14613 (N_14613,N_13322,N_13174);
nor U14614 (N_14614,N_13564,N_13293);
nor U14615 (N_14615,N_13369,N_13789);
and U14616 (N_14616,N_13159,N_13096);
and U14617 (N_14617,N_13100,N_13419);
and U14618 (N_14618,N_13987,N_13395);
nand U14619 (N_14619,N_13907,N_13600);
and U14620 (N_14620,N_13035,N_13937);
nor U14621 (N_14621,N_13556,N_13299);
or U14622 (N_14622,N_13794,N_13006);
or U14623 (N_14623,N_13697,N_13112);
nor U14624 (N_14624,N_13939,N_13303);
xor U14625 (N_14625,N_13845,N_13716);
and U14626 (N_14626,N_13041,N_13955);
xnor U14627 (N_14627,N_13090,N_13577);
or U14628 (N_14628,N_13272,N_13948);
and U14629 (N_14629,N_13059,N_13312);
or U14630 (N_14630,N_13695,N_13248);
nor U14631 (N_14631,N_13533,N_13219);
nor U14632 (N_14632,N_13584,N_13937);
or U14633 (N_14633,N_13348,N_13095);
xnor U14634 (N_14634,N_13709,N_13805);
or U14635 (N_14635,N_13588,N_13863);
nand U14636 (N_14636,N_13710,N_13836);
nand U14637 (N_14637,N_13485,N_13150);
or U14638 (N_14638,N_13757,N_13074);
xnor U14639 (N_14639,N_13541,N_13462);
xor U14640 (N_14640,N_13384,N_13818);
nand U14641 (N_14641,N_13399,N_13340);
xnor U14642 (N_14642,N_13340,N_13285);
or U14643 (N_14643,N_13032,N_13163);
nor U14644 (N_14644,N_13663,N_13138);
and U14645 (N_14645,N_13135,N_13632);
xnor U14646 (N_14646,N_13554,N_13566);
nor U14647 (N_14647,N_13362,N_13973);
and U14648 (N_14648,N_13035,N_13383);
or U14649 (N_14649,N_13100,N_13117);
or U14650 (N_14650,N_13201,N_13415);
and U14651 (N_14651,N_13203,N_13735);
xor U14652 (N_14652,N_13777,N_13336);
xor U14653 (N_14653,N_13788,N_13515);
nand U14654 (N_14654,N_13428,N_13373);
xor U14655 (N_14655,N_13259,N_13864);
nor U14656 (N_14656,N_13753,N_13463);
nor U14657 (N_14657,N_13255,N_13709);
or U14658 (N_14658,N_13353,N_13228);
and U14659 (N_14659,N_13001,N_13359);
nand U14660 (N_14660,N_13001,N_13343);
xnor U14661 (N_14661,N_13185,N_13442);
nand U14662 (N_14662,N_13107,N_13866);
nor U14663 (N_14663,N_13818,N_13197);
xor U14664 (N_14664,N_13062,N_13020);
and U14665 (N_14665,N_13462,N_13961);
and U14666 (N_14666,N_13169,N_13582);
and U14667 (N_14667,N_13773,N_13754);
or U14668 (N_14668,N_13192,N_13986);
or U14669 (N_14669,N_13384,N_13064);
nand U14670 (N_14670,N_13908,N_13558);
xor U14671 (N_14671,N_13759,N_13555);
or U14672 (N_14672,N_13663,N_13345);
xnor U14673 (N_14673,N_13159,N_13756);
or U14674 (N_14674,N_13646,N_13531);
xnor U14675 (N_14675,N_13408,N_13514);
xnor U14676 (N_14676,N_13438,N_13628);
and U14677 (N_14677,N_13323,N_13762);
nand U14678 (N_14678,N_13349,N_13991);
xnor U14679 (N_14679,N_13129,N_13338);
xnor U14680 (N_14680,N_13420,N_13402);
or U14681 (N_14681,N_13187,N_13142);
xnor U14682 (N_14682,N_13560,N_13257);
nand U14683 (N_14683,N_13134,N_13159);
xor U14684 (N_14684,N_13971,N_13802);
or U14685 (N_14685,N_13348,N_13860);
nand U14686 (N_14686,N_13907,N_13864);
xnor U14687 (N_14687,N_13737,N_13576);
nor U14688 (N_14688,N_13694,N_13478);
nor U14689 (N_14689,N_13577,N_13823);
xor U14690 (N_14690,N_13240,N_13110);
and U14691 (N_14691,N_13557,N_13993);
nand U14692 (N_14692,N_13878,N_13830);
or U14693 (N_14693,N_13384,N_13532);
xor U14694 (N_14694,N_13579,N_13721);
or U14695 (N_14695,N_13805,N_13706);
nor U14696 (N_14696,N_13016,N_13905);
and U14697 (N_14697,N_13864,N_13144);
xnor U14698 (N_14698,N_13649,N_13304);
or U14699 (N_14699,N_13487,N_13846);
nor U14700 (N_14700,N_13480,N_13018);
nand U14701 (N_14701,N_13300,N_13225);
nand U14702 (N_14702,N_13580,N_13690);
nand U14703 (N_14703,N_13094,N_13722);
and U14704 (N_14704,N_13847,N_13600);
xnor U14705 (N_14705,N_13069,N_13766);
and U14706 (N_14706,N_13548,N_13805);
nand U14707 (N_14707,N_13520,N_13475);
xnor U14708 (N_14708,N_13328,N_13630);
xor U14709 (N_14709,N_13665,N_13479);
nor U14710 (N_14710,N_13081,N_13911);
nor U14711 (N_14711,N_13308,N_13748);
nor U14712 (N_14712,N_13592,N_13471);
nand U14713 (N_14713,N_13478,N_13964);
nand U14714 (N_14714,N_13845,N_13491);
nor U14715 (N_14715,N_13387,N_13923);
xnor U14716 (N_14716,N_13660,N_13696);
nand U14717 (N_14717,N_13851,N_13470);
or U14718 (N_14718,N_13426,N_13468);
xor U14719 (N_14719,N_13977,N_13670);
xnor U14720 (N_14720,N_13995,N_13557);
nand U14721 (N_14721,N_13064,N_13754);
and U14722 (N_14722,N_13950,N_13913);
nor U14723 (N_14723,N_13400,N_13601);
nor U14724 (N_14724,N_13283,N_13932);
xor U14725 (N_14725,N_13798,N_13215);
or U14726 (N_14726,N_13433,N_13400);
or U14727 (N_14727,N_13384,N_13387);
or U14728 (N_14728,N_13203,N_13931);
or U14729 (N_14729,N_13126,N_13698);
nand U14730 (N_14730,N_13907,N_13201);
nor U14731 (N_14731,N_13490,N_13393);
xnor U14732 (N_14732,N_13114,N_13545);
xor U14733 (N_14733,N_13190,N_13738);
nand U14734 (N_14734,N_13262,N_13763);
and U14735 (N_14735,N_13110,N_13131);
nand U14736 (N_14736,N_13726,N_13601);
nand U14737 (N_14737,N_13946,N_13587);
nand U14738 (N_14738,N_13155,N_13709);
nand U14739 (N_14739,N_13004,N_13329);
xnor U14740 (N_14740,N_13683,N_13465);
nor U14741 (N_14741,N_13381,N_13773);
and U14742 (N_14742,N_13421,N_13347);
xor U14743 (N_14743,N_13161,N_13296);
nand U14744 (N_14744,N_13645,N_13735);
xnor U14745 (N_14745,N_13967,N_13905);
nand U14746 (N_14746,N_13196,N_13366);
and U14747 (N_14747,N_13300,N_13273);
and U14748 (N_14748,N_13276,N_13329);
xnor U14749 (N_14749,N_13335,N_13750);
xor U14750 (N_14750,N_13664,N_13984);
or U14751 (N_14751,N_13736,N_13080);
xnor U14752 (N_14752,N_13935,N_13350);
nor U14753 (N_14753,N_13419,N_13770);
or U14754 (N_14754,N_13204,N_13322);
and U14755 (N_14755,N_13834,N_13284);
xor U14756 (N_14756,N_13442,N_13362);
nor U14757 (N_14757,N_13757,N_13669);
xor U14758 (N_14758,N_13117,N_13253);
xor U14759 (N_14759,N_13148,N_13407);
nand U14760 (N_14760,N_13757,N_13688);
or U14761 (N_14761,N_13049,N_13370);
nand U14762 (N_14762,N_13557,N_13871);
and U14763 (N_14763,N_13820,N_13239);
or U14764 (N_14764,N_13828,N_13880);
or U14765 (N_14765,N_13855,N_13705);
or U14766 (N_14766,N_13848,N_13432);
nand U14767 (N_14767,N_13030,N_13765);
and U14768 (N_14768,N_13819,N_13611);
or U14769 (N_14769,N_13095,N_13023);
nand U14770 (N_14770,N_13162,N_13219);
and U14771 (N_14771,N_13783,N_13191);
or U14772 (N_14772,N_13668,N_13462);
nand U14773 (N_14773,N_13597,N_13677);
xor U14774 (N_14774,N_13238,N_13760);
or U14775 (N_14775,N_13959,N_13528);
nand U14776 (N_14776,N_13397,N_13355);
xor U14777 (N_14777,N_13043,N_13319);
xnor U14778 (N_14778,N_13278,N_13318);
nand U14779 (N_14779,N_13851,N_13051);
nand U14780 (N_14780,N_13092,N_13491);
xor U14781 (N_14781,N_13131,N_13876);
and U14782 (N_14782,N_13602,N_13745);
and U14783 (N_14783,N_13665,N_13442);
or U14784 (N_14784,N_13016,N_13393);
xor U14785 (N_14785,N_13961,N_13354);
and U14786 (N_14786,N_13019,N_13951);
or U14787 (N_14787,N_13765,N_13535);
or U14788 (N_14788,N_13276,N_13959);
nand U14789 (N_14789,N_13345,N_13629);
or U14790 (N_14790,N_13967,N_13552);
xnor U14791 (N_14791,N_13870,N_13089);
and U14792 (N_14792,N_13530,N_13034);
or U14793 (N_14793,N_13796,N_13183);
xnor U14794 (N_14794,N_13648,N_13962);
or U14795 (N_14795,N_13035,N_13961);
xnor U14796 (N_14796,N_13038,N_13304);
or U14797 (N_14797,N_13617,N_13274);
or U14798 (N_14798,N_13958,N_13095);
nand U14799 (N_14799,N_13689,N_13408);
nor U14800 (N_14800,N_13177,N_13808);
nand U14801 (N_14801,N_13034,N_13023);
xnor U14802 (N_14802,N_13367,N_13913);
nand U14803 (N_14803,N_13469,N_13318);
or U14804 (N_14804,N_13301,N_13493);
xnor U14805 (N_14805,N_13198,N_13340);
xnor U14806 (N_14806,N_13725,N_13261);
nor U14807 (N_14807,N_13190,N_13503);
nor U14808 (N_14808,N_13565,N_13933);
and U14809 (N_14809,N_13964,N_13489);
nor U14810 (N_14810,N_13221,N_13456);
or U14811 (N_14811,N_13774,N_13720);
or U14812 (N_14812,N_13678,N_13396);
nand U14813 (N_14813,N_13943,N_13969);
or U14814 (N_14814,N_13467,N_13541);
nand U14815 (N_14815,N_13327,N_13471);
or U14816 (N_14816,N_13939,N_13992);
or U14817 (N_14817,N_13183,N_13784);
and U14818 (N_14818,N_13351,N_13950);
or U14819 (N_14819,N_13976,N_13285);
or U14820 (N_14820,N_13170,N_13039);
and U14821 (N_14821,N_13417,N_13622);
and U14822 (N_14822,N_13302,N_13035);
nand U14823 (N_14823,N_13047,N_13701);
and U14824 (N_14824,N_13241,N_13309);
and U14825 (N_14825,N_13233,N_13178);
xor U14826 (N_14826,N_13994,N_13753);
nand U14827 (N_14827,N_13834,N_13253);
nor U14828 (N_14828,N_13922,N_13515);
xor U14829 (N_14829,N_13180,N_13064);
xor U14830 (N_14830,N_13933,N_13916);
or U14831 (N_14831,N_13592,N_13664);
or U14832 (N_14832,N_13829,N_13501);
nor U14833 (N_14833,N_13175,N_13292);
nor U14834 (N_14834,N_13071,N_13208);
and U14835 (N_14835,N_13721,N_13346);
nor U14836 (N_14836,N_13910,N_13455);
nand U14837 (N_14837,N_13701,N_13072);
or U14838 (N_14838,N_13633,N_13534);
nand U14839 (N_14839,N_13912,N_13274);
nor U14840 (N_14840,N_13366,N_13567);
and U14841 (N_14841,N_13107,N_13321);
or U14842 (N_14842,N_13102,N_13927);
and U14843 (N_14843,N_13746,N_13632);
and U14844 (N_14844,N_13990,N_13236);
nand U14845 (N_14845,N_13902,N_13834);
and U14846 (N_14846,N_13284,N_13845);
nand U14847 (N_14847,N_13211,N_13832);
xor U14848 (N_14848,N_13840,N_13031);
xnor U14849 (N_14849,N_13100,N_13414);
or U14850 (N_14850,N_13531,N_13492);
and U14851 (N_14851,N_13887,N_13960);
or U14852 (N_14852,N_13635,N_13725);
nor U14853 (N_14853,N_13765,N_13400);
nor U14854 (N_14854,N_13958,N_13225);
or U14855 (N_14855,N_13990,N_13689);
nand U14856 (N_14856,N_13935,N_13889);
and U14857 (N_14857,N_13358,N_13459);
nand U14858 (N_14858,N_13374,N_13837);
nor U14859 (N_14859,N_13849,N_13228);
xnor U14860 (N_14860,N_13529,N_13669);
nor U14861 (N_14861,N_13428,N_13223);
xor U14862 (N_14862,N_13704,N_13525);
and U14863 (N_14863,N_13244,N_13396);
and U14864 (N_14864,N_13936,N_13902);
nand U14865 (N_14865,N_13140,N_13049);
nand U14866 (N_14866,N_13675,N_13519);
nor U14867 (N_14867,N_13602,N_13414);
and U14868 (N_14868,N_13638,N_13597);
nor U14869 (N_14869,N_13421,N_13158);
or U14870 (N_14870,N_13830,N_13239);
nand U14871 (N_14871,N_13320,N_13716);
and U14872 (N_14872,N_13446,N_13317);
nand U14873 (N_14873,N_13688,N_13179);
nor U14874 (N_14874,N_13651,N_13246);
nor U14875 (N_14875,N_13338,N_13701);
nand U14876 (N_14876,N_13235,N_13372);
or U14877 (N_14877,N_13097,N_13145);
or U14878 (N_14878,N_13913,N_13563);
xnor U14879 (N_14879,N_13317,N_13306);
or U14880 (N_14880,N_13752,N_13661);
nor U14881 (N_14881,N_13363,N_13025);
nand U14882 (N_14882,N_13982,N_13856);
xor U14883 (N_14883,N_13080,N_13542);
xnor U14884 (N_14884,N_13045,N_13834);
and U14885 (N_14885,N_13723,N_13417);
or U14886 (N_14886,N_13547,N_13047);
or U14887 (N_14887,N_13255,N_13115);
xnor U14888 (N_14888,N_13166,N_13658);
xor U14889 (N_14889,N_13929,N_13363);
nor U14890 (N_14890,N_13379,N_13009);
or U14891 (N_14891,N_13226,N_13532);
nor U14892 (N_14892,N_13317,N_13576);
nor U14893 (N_14893,N_13775,N_13724);
and U14894 (N_14894,N_13060,N_13253);
nor U14895 (N_14895,N_13627,N_13512);
nor U14896 (N_14896,N_13849,N_13285);
nor U14897 (N_14897,N_13533,N_13091);
nand U14898 (N_14898,N_13853,N_13715);
or U14899 (N_14899,N_13370,N_13783);
nor U14900 (N_14900,N_13318,N_13128);
nor U14901 (N_14901,N_13047,N_13779);
xor U14902 (N_14902,N_13163,N_13172);
xnor U14903 (N_14903,N_13301,N_13237);
xnor U14904 (N_14904,N_13338,N_13158);
nand U14905 (N_14905,N_13022,N_13154);
or U14906 (N_14906,N_13504,N_13687);
nand U14907 (N_14907,N_13826,N_13922);
or U14908 (N_14908,N_13681,N_13711);
and U14909 (N_14909,N_13212,N_13662);
nor U14910 (N_14910,N_13577,N_13368);
nor U14911 (N_14911,N_13654,N_13674);
nor U14912 (N_14912,N_13399,N_13368);
nor U14913 (N_14913,N_13161,N_13217);
or U14914 (N_14914,N_13232,N_13645);
or U14915 (N_14915,N_13526,N_13146);
xor U14916 (N_14916,N_13701,N_13418);
or U14917 (N_14917,N_13635,N_13152);
nand U14918 (N_14918,N_13359,N_13392);
nor U14919 (N_14919,N_13047,N_13534);
nor U14920 (N_14920,N_13848,N_13761);
or U14921 (N_14921,N_13113,N_13977);
nand U14922 (N_14922,N_13849,N_13772);
and U14923 (N_14923,N_13789,N_13739);
and U14924 (N_14924,N_13119,N_13954);
xnor U14925 (N_14925,N_13817,N_13363);
or U14926 (N_14926,N_13049,N_13134);
and U14927 (N_14927,N_13966,N_13041);
nand U14928 (N_14928,N_13087,N_13246);
nor U14929 (N_14929,N_13956,N_13666);
and U14930 (N_14930,N_13149,N_13130);
and U14931 (N_14931,N_13831,N_13949);
and U14932 (N_14932,N_13370,N_13366);
nand U14933 (N_14933,N_13035,N_13357);
and U14934 (N_14934,N_13054,N_13022);
xor U14935 (N_14935,N_13382,N_13236);
nand U14936 (N_14936,N_13733,N_13427);
xnor U14937 (N_14937,N_13417,N_13448);
xnor U14938 (N_14938,N_13419,N_13068);
xor U14939 (N_14939,N_13548,N_13892);
nand U14940 (N_14940,N_13778,N_13746);
nand U14941 (N_14941,N_13853,N_13501);
or U14942 (N_14942,N_13316,N_13513);
nor U14943 (N_14943,N_13187,N_13923);
and U14944 (N_14944,N_13702,N_13947);
or U14945 (N_14945,N_13277,N_13820);
nand U14946 (N_14946,N_13886,N_13548);
nor U14947 (N_14947,N_13628,N_13604);
and U14948 (N_14948,N_13473,N_13465);
xor U14949 (N_14949,N_13699,N_13595);
and U14950 (N_14950,N_13884,N_13987);
nor U14951 (N_14951,N_13948,N_13587);
nor U14952 (N_14952,N_13096,N_13351);
nand U14953 (N_14953,N_13526,N_13359);
nand U14954 (N_14954,N_13737,N_13715);
and U14955 (N_14955,N_13630,N_13702);
and U14956 (N_14956,N_13159,N_13082);
nand U14957 (N_14957,N_13504,N_13403);
nor U14958 (N_14958,N_13784,N_13474);
and U14959 (N_14959,N_13279,N_13398);
or U14960 (N_14960,N_13742,N_13814);
xnor U14961 (N_14961,N_13432,N_13891);
or U14962 (N_14962,N_13357,N_13618);
or U14963 (N_14963,N_13018,N_13584);
xnor U14964 (N_14964,N_13908,N_13360);
nand U14965 (N_14965,N_13509,N_13796);
or U14966 (N_14966,N_13391,N_13585);
or U14967 (N_14967,N_13018,N_13911);
nand U14968 (N_14968,N_13830,N_13428);
and U14969 (N_14969,N_13975,N_13410);
or U14970 (N_14970,N_13232,N_13729);
and U14971 (N_14971,N_13365,N_13950);
nor U14972 (N_14972,N_13756,N_13938);
or U14973 (N_14973,N_13782,N_13346);
and U14974 (N_14974,N_13766,N_13001);
or U14975 (N_14975,N_13986,N_13199);
and U14976 (N_14976,N_13341,N_13671);
or U14977 (N_14977,N_13745,N_13037);
and U14978 (N_14978,N_13037,N_13972);
xnor U14979 (N_14979,N_13126,N_13531);
and U14980 (N_14980,N_13668,N_13881);
and U14981 (N_14981,N_13873,N_13911);
and U14982 (N_14982,N_13386,N_13310);
nand U14983 (N_14983,N_13255,N_13916);
xor U14984 (N_14984,N_13592,N_13564);
and U14985 (N_14985,N_13934,N_13750);
nand U14986 (N_14986,N_13156,N_13634);
and U14987 (N_14987,N_13080,N_13719);
xnor U14988 (N_14988,N_13212,N_13646);
xor U14989 (N_14989,N_13086,N_13483);
nor U14990 (N_14990,N_13224,N_13832);
or U14991 (N_14991,N_13706,N_13735);
or U14992 (N_14992,N_13153,N_13238);
and U14993 (N_14993,N_13445,N_13618);
nand U14994 (N_14994,N_13166,N_13466);
nand U14995 (N_14995,N_13136,N_13541);
xnor U14996 (N_14996,N_13847,N_13790);
and U14997 (N_14997,N_13137,N_13499);
and U14998 (N_14998,N_13753,N_13770);
and U14999 (N_14999,N_13263,N_13064);
xnor UO_0 (O_0,N_14225,N_14547);
and UO_1 (O_1,N_14360,N_14365);
nor UO_2 (O_2,N_14172,N_14155);
nor UO_3 (O_3,N_14859,N_14196);
and UO_4 (O_4,N_14983,N_14495);
nand UO_5 (O_5,N_14799,N_14074);
nor UO_6 (O_6,N_14683,N_14181);
nor UO_7 (O_7,N_14791,N_14845);
and UO_8 (O_8,N_14284,N_14209);
or UO_9 (O_9,N_14819,N_14414);
xnor UO_10 (O_10,N_14733,N_14251);
and UO_11 (O_11,N_14352,N_14182);
and UO_12 (O_12,N_14956,N_14383);
nand UO_13 (O_13,N_14496,N_14295);
or UO_14 (O_14,N_14067,N_14356);
and UO_15 (O_15,N_14232,N_14484);
nor UO_16 (O_16,N_14347,N_14389);
and UO_17 (O_17,N_14185,N_14823);
and UO_18 (O_18,N_14513,N_14612);
and UO_19 (O_19,N_14237,N_14587);
or UO_20 (O_20,N_14221,N_14787);
xor UO_21 (O_21,N_14243,N_14623);
nand UO_22 (O_22,N_14061,N_14380);
or UO_23 (O_23,N_14491,N_14811);
xnor UO_24 (O_24,N_14813,N_14624);
nand UO_25 (O_25,N_14009,N_14081);
or UO_26 (O_26,N_14563,N_14311);
nor UO_27 (O_27,N_14667,N_14040);
nand UO_28 (O_28,N_14660,N_14218);
nand UO_29 (O_29,N_14766,N_14674);
or UO_30 (O_30,N_14903,N_14871);
nand UO_31 (O_31,N_14960,N_14493);
xor UO_32 (O_32,N_14384,N_14482);
nand UO_33 (O_33,N_14275,N_14179);
nand UO_34 (O_34,N_14515,N_14934);
and UO_35 (O_35,N_14720,N_14304);
or UO_36 (O_36,N_14643,N_14933);
and UO_37 (O_37,N_14989,N_14600);
nand UO_38 (O_38,N_14200,N_14068);
and UO_39 (O_39,N_14235,N_14456);
nor UO_40 (O_40,N_14052,N_14533);
nand UO_41 (O_41,N_14313,N_14682);
nand UO_42 (O_42,N_14827,N_14062);
xor UO_43 (O_43,N_14096,N_14373);
and UO_44 (O_44,N_14930,N_14854);
or UO_45 (O_45,N_14162,N_14400);
nand UO_46 (O_46,N_14214,N_14160);
and UO_47 (O_47,N_14509,N_14542);
xor UO_48 (O_48,N_14034,N_14281);
nor UO_49 (O_49,N_14511,N_14986);
or UO_50 (O_50,N_14696,N_14878);
nand UO_51 (O_51,N_14844,N_14135);
or UO_52 (O_52,N_14023,N_14118);
nor UO_53 (O_53,N_14578,N_14599);
xnor UO_54 (O_54,N_14064,N_14216);
xnor UO_55 (O_55,N_14171,N_14724);
and UO_56 (O_56,N_14539,N_14601);
and UO_57 (O_57,N_14357,N_14111);
nand UO_58 (O_58,N_14280,N_14525);
or UO_59 (O_59,N_14288,N_14589);
nor UO_60 (O_60,N_14749,N_14969);
nor UO_61 (O_61,N_14371,N_14714);
nand UO_62 (O_62,N_14671,N_14409);
nor UO_63 (O_63,N_14688,N_14302);
nand UO_64 (O_64,N_14398,N_14085);
nand UO_65 (O_65,N_14133,N_14173);
nand UO_66 (O_66,N_14194,N_14189);
xor UO_67 (O_67,N_14026,N_14211);
xor UO_68 (O_68,N_14432,N_14917);
nand UO_69 (O_69,N_14337,N_14928);
nand UO_70 (O_70,N_14348,N_14834);
xnor UO_71 (O_71,N_14943,N_14018);
nand UO_72 (O_72,N_14261,N_14838);
nor UO_73 (O_73,N_14388,N_14748);
nor UO_74 (O_74,N_14494,N_14988);
nand UO_75 (O_75,N_14810,N_14359);
xnor UO_76 (O_76,N_14982,N_14307);
nand UO_77 (O_77,N_14056,N_14148);
xor UO_78 (O_78,N_14907,N_14492);
nand UO_79 (O_79,N_14490,N_14806);
or UO_80 (O_80,N_14726,N_14761);
or UO_81 (O_81,N_14752,N_14922);
nand UO_82 (O_82,N_14408,N_14792);
and UO_83 (O_83,N_14676,N_14168);
nor UO_84 (O_84,N_14508,N_14099);
xnor UO_85 (O_85,N_14422,N_14774);
nand UO_86 (O_86,N_14809,N_14438);
and UO_87 (O_87,N_14603,N_14962);
and UO_88 (O_88,N_14729,N_14620);
or UO_89 (O_89,N_14426,N_14912);
nand UO_90 (O_90,N_14004,N_14655);
nor UO_91 (O_91,N_14979,N_14025);
nor UO_92 (O_92,N_14807,N_14385);
nor UO_93 (O_93,N_14535,N_14124);
nand UO_94 (O_94,N_14376,N_14022);
nand UO_95 (O_95,N_14001,N_14862);
nor UO_96 (O_96,N_14691,N_14929);
xor UO_97 (O_97,N_14268,N_14763);
nor UO_98 (O_98,N_14139,N_14233);
nor UO_99 (O_99,N_14522,N_14372);
nor UO_100 (O_100,N_14657,N_14727);
xnor UO_101 (O_101,N_14543,N_14773);
and UO_102 (O_102,N_14919,N_14648);
or UO_103 (O_103,N_14101,N_14636);
nand UO_104 (O_104,N_14379,N_14978);
xor UO_105 (O_105,N_14423,N_14204);
xor UO_106 (O_106,N_14941,N_14707);
or UO_107 (O_107,N_14421,N_14606);
xnor UO_108 (O_108,N_14569,N_14320);
nand UO_109 (O_109,N_14427,N_14220);
and UO_110 (O_110,N_14402,N_14367);
or UO_111 (O_111,N_14802,N_14132);
and UO_112 (O_112,N_14458,N_14293);
or UO_113 (O_113,N_14800,N_14972);
xor UO_114 (O_114,N_14425,N_14825);
and UO_115 (O_115,N_14574,N_14528);
xor UO_116 (O_116,N_14954,N_14159);
xor UO_117 (O_117,N_14805,N_14127);
and UO_118 (O_118,N_14417,N_14582);
nor UO_119 (O_119,N_14897,N_14297);
xor UO_120 (O_120,N_14430,N_14997);
and UO_121 (O_121,N_14650,N_14397);
and UO_122 (O_122,N_14286,N_14548);
xor UO_123 (O_123,N_14245,N_14571);
nand UO_124 (O_124,N_14579,N_14663);
or UO_125 (O_125,N_14649,N_14622);
nand UO_126 (O_126,N_14681,N_14700);
and UO_127 (O_127,N_14830,N_14479);
or UO_128 (O_128,N_14735,N_14814);
nor UO_129 (O_129,N_14291,N_14345);
and UO_130 (O_130,N_14044,N_14103);
nand UO_131 (O_131,N_14049,N_14770);
nor UO_132 (O_132,N_14699,N_14977);
or UO_133 (O_133,N_14002,N_14043);
or UO_134 (O_134,N_14836,N_14324);
and UO_135 (O_135,N_14222,N_14795);
nand UO_136 (O_136,N_14784,N_14684);
nor UO_137 (O_137,N_14303,N_14391);
nand UO_138 (O_138,N_14153,N_14079);
and UO_139 (O_139,N_14029,N_14147);
and UO_140 (O_140,N_14829,N_14666);
and UO_141 (O_141,N_14927,N_14771);
and UO_142 (O_142,N_14070,N_14236);
and UO_143 (O_143,N_14312,N_14607);
nand UO_144 (O_144,N_14234,N_14856);
or UO_145 (O_145,N_14860,N_14888);
or UO_146 (O_146,N_14412,N_14690);
or UO_147 (O_147,N_14781,N_14219);
and UO_148 (O_148,N_14947,N_14405);
nand UO_149 (O_149,N_14102,N_14531);
xor UO_150 (O_150,N_14580,N_14306);
and UO_151 (O_151,N_14595,N_14499);
or UO_152 (O_152,N_14540,N_14920);
nor UO_153 (O_153,N_14488,N_14551);
nor UO_154 (O_154,N_14410,N_14713);
nor UO_155 (O_155,N_14377,N_14190);
nor UO_156 (O_156,N_14392,N_14014);
nand UO_157 (O_157,N_14276,N_14449);
and UO_158 (O_158,N_14180,N_14154);
or UO_159 (O_159,N_14705,N_14646);
nand UO_160 (O_160,N_14487,N_14723);
xnor UO_161 (O_161,N_14901,N_14529);
nand UO_162 (O_162,N_14635,N_14776);
nand UO_163 (O_163,N_14461,N_14407);
nand UO_164 (O_164,N_14145,N_14550);
and UO_165 (O_165,N_14831,N_14489);
nand UO_166 (O_166,N_14537,N_14501);
and UO_167 (O_167,N_14904,N_14704);
or UO_168 (O_168,N_14203,N_14249);
nor UO_169 (O_169,N_14339,N_14327);
nor UO_170 (O_170,N_14703,N_14980);
or UO_171 (O_171,N_14273,N_14137);
nand UO_172 (O_172,N_14712,N_14740);
or UO_173 (O_173,N_14474,N_14966);
nor UO_174 (O_174,N_14082,N_14305);
nand UO_175 (O_175,N_14861,N_14891);
xor UO_176 (O_176,N_14653,N_14785);
or UO_177 (O_177,N_14875,N_14072);
nand UO_178 (O_178,N_14030,N_14151);
xnor UO_179 (O_179,N_14007,N_14626);
or UO_180 (O_180,N_14931,N_14374);
xor UO_181 (O_181,N_14323,N_14149);
and UO_182 (O_182,N_14129,N_14368);
or UO_183 (O_183,N_14677,N_14447);
or UO_184 (O_184,N_14801,N_14957);
nand UO_185 (O_185,N_14885,N_14546);
nand UO_186 (O_186,N_14812,N_14575);
nor UO_187 (O_187,N_14640,N_14621);
nand UO_188 (O_188,N_14538,N_14981);
nor UO_189 (O_189,N_14566,N_14473);
nor UO_190 (O_190,N_14448,N_14033);
or UO_191 (O_191,N_14270,N_14775);
xnor UO_192 (O_192,N_14892,N_14326);
nor UO_193 (O_193,N_14021,N_14946);
nand UO_194 (O_194,N_14319,N_14170);
xnor UO_195 (O_195,N_14843,N_14224);
and UO_196 (O_196,N_14950,N_14316);
xor UO_197 (O_197,N_14475,N_14262);
nand UO_198 (O_198,N_14876,N_14338);
or UO_199 (O_199,N_14116,N_14877);
nand UO_200 (O_200,N_14695,N_14485);
nand UO_201 (O_201,N_14730,N_14586);
nand UO_202 (O_202,N_14758,N_14738);
nand UO_203 (O_203,N_14340,N_14736);
nor UO_204 (O_204,N_14864,N_14751);
and UO_205 (O_205,N_14017,N_14290);
nor UO_206 (O_206,N_14750,N_14363);
nand UO_207 (O_207,N_14793,N_14047);
nand UO_208 (O_208,N_14241,N_14144);
xor UO_209 (O_209,N_14138,N_14207);
and UO_210 (O_210,N_14974,N_14136);
or UO_211 (O_211,N_14767,N_14822);
nand UO_212 (O_212,N_14764,N_14000);
and UO_213 (O_213,N_14431,N_14527);
or UO_214 (O_214,N_14470,N_14742);
xor UO_215 (O_215,N_14433,N_14143);
xnor UO_216 (O_216,N_14651,N_14900);
xnor UO_217 (O_217,N_14344,N_14559);
xnor UO_218 (O_218,N_14045,N_14743);
nor UO_219 (O_219,N_14369,N_14746);
xnor UO_220 (O_220,N_14741,N_14006);
nand UO_221 (O_221,N_14213,N_14121);
and UO_222 (O_222,N_14734,N_14274);
nand UO_223 (O_223,N_14076,N_14205);
nand UO_224 (O_224,N_14027,N_14759);
or UO_225 (O_225,N_14505,N_14038);
and UO_226 (O_226,N_14668,N_14396);
and UO_227 (O_227,N_14887,N_14465);
nand UO_228 (O_228,N_14685,N_14973);
or UO_229 (O_229,N_14665,N_14012);
or UO_230 (O_230,N_14353,N_14625);
xnor UO_231 (O_231,N_14769,N_14544);
xor UO_232 (O_232,N_14087,N_14105);
nor UO_233 (O_233,N_14906,N_14015);
nor UO_234 (O_234,N_14454,N_14697);
xor UO_235 (O_235,N_14619,N_14710);
or UO_236 (O_236,N_14277,N_14238);
xor UO_237 (O_237,N_14177,N_14639);
nand UO_238 (O_238,N_14024,N_14406);
and UO_239 (O_239,N_14112,N_14504);
or UO_240 (O_240,N_14679,N_14754);
or UO_241 (O_241,N_14558,N_14174);
xnor UO_242 (O_242,N_14782,N_14628);
xnor UO_243 (O_243,N_14967,N_14924);
nor UO_244 (O_244,N_14593,N_14768);
and UO_245 (O_245,N_14991,N_14197);
nand UO_246 (O_246,N_14602,N_14965);
or UO_247 (O_247,N_14336,N_14552);
xor UO_248 (O_248,N_14739,N_14790);
nand UO_249 (O_249,N_14199,N_14868);
or UO_250 (O_250,N_14202,N_14898);
nor UO_251 (O_251,N_14325,N_14945);
nor UO_252 (O_252,N_14872,N_14106);
or UO_253 (O_253,N_14926,N_14851);
xor UO_254 (O_254,N_14053,N_14016);
and UO_255 (O_255,N_14899,N_14075);
nand UO_256 (O_256,N_14287,N_14242);
nand UO_257 (O_257,N_14618,N_14258);
or UO_258 (O_258,N_14446,N_14497);
or UO_259 (O_259,N_14554,N_14778);
nand UO_260 (O_260,N_14637,N_14048);
nand UO_261 (O_261,N_14510,N_14902);
or UO_262 (O_262,N_14436,N_14869);
nand UO_263 (O_263,N_14706,N_14250);
or UO_264 (O_264,N_14330,N_14178);
nor UO_265 (O_265,N_14013,N_14095);
and UO_266 (O_266,N_14131,N_14835);
nor UO_267 (O_267,N_14915,N_14317);
xor UO_268 (O_268,N_14894,N_14630);
nor UO_269 (O_269,N_14298,N_14999);
and UO_270 (O_270,N_14477,N_14963);
or UO_271 (O_271,N_14632,N_14937);
xor UO_272 (O_272,N_14032,N_14094);
and UO_273 (O_273,N_14597,N_14942);
and UO_274 (O_274,N_14987,N_14254);
nand UO_275 (O_275,N_14523,N_14731);
xor UO_276 (O_276,N_14158,N_14737);
xnor UO_277 (O_277,N_14150,N_14516);
nand UO_278 (O_278,N_14351,N_14584);
and UO_279 (O_279,N_14610,N_14721);
nor UO_280 (O_280,N_14354,N_14362);
xnor UO_281 (O_281,N_14483,N_14654);
xnor UO_282 (O_282,N_14279,N_14985);
and UO_283 (O_283,N_14512,N_14698);
or UO_284 (O_284,N_14517,N_14944);
or UO_285 (O_285,N_14975,N_14964);
nand UO_286 (O_286,N_14005,N_14702);
nand UO_287 (O_287,N_14780,N_14169);
or UO_288 (O_288,N_14718,N_14108);
nor UO_289 (O_289,N_14824,N_14914);
or UO_290 (O_290,N_14210,N_14100);
nor UO_291 (O_291,N_14318,N_14846);
and UO_292 (O_292,N_14530,N_14532);
nor UO_293 (O_293,N_14450,N_14455);
nand UO_294 (O_294,N_14553,N_14193);
nor UO_295 (O_295,N_14853,N_14577);
xnor UO_296 (O_296,N_14227,N_14109);
or UO_297 (O_297,N_14083,N_14267);
xnor UO_298 (O_298,N_14228,N_14804);
xor UO_299 (O_299,N_14673,N_14609);
and UO_300 (O_300,N_14886,N_14728);
or UO_301 (O_301,N_14858,N_14452);
nor UO_302 (O_302,N_14428,N_14939);
xnor UO_303 (O_303,N_14059,N_14998);
or UO_304 (O_304,N_14188,N_14300);
nor UO_305 (O_305,N_14166,N_14925);
and UO_306 (O_306,N_14037,N_14818);
nor UO_307 (O_307,N_14289,N_14870);
nand UO_308 (O_308,N_14255,N_14263);
or UO_309 (O_309,N_14073,N_14366);
or UO_310 (O_310,N_14215,N_14745);
xnor UO_311 (O_311,N_14570,N_14451);
and UO_312 (O_312,N_14549,N_14918);
and UO_313 (O_313,N_14019,N_14386);
or UO_314 (O_314,N_14594,N_14265);
or UO_315 (O_315,N_14541,N_14747);
nor UO_316 (O_316,N_14208,N_14175);
nor UO_317 (O_317,N_14156,N_14343);
and UO_318 (O_318,N_14206,N_14309);
or UO_319 (O_319,N_14585,N_14744);
xor UO_320 (O_320,N_14832,N_14874);
or UO_321 (O_321,N_14011,N_14756);
or UO_322 (O_322,N_14916,N_14641);
nand UO_323 (O_323,N_14990,N_14050);
nor UO_324 (O_324,N_14692,N_14908);
nand UO_325 (O_325,N_14664,N_14534);
and UO_326 (O_326,N_14370,N_14439);
and UO_327 (O_327,N_14857,N_14656);
and UO_328 (O_328,N_14058,N_14350);
and UO_329 (O_329,N_14355,N_14520);
nor UO_330 (O_330,N_14468,N_14266);
nor UO_331 (O_331,N_14481,N_14244);
or UO_332 (O_332,N_14036,N_14847);
xnor UO_333 (O_333,N_14349,N_14562);
or UO_334 (O_334,N_14722,N_14993);
nor UO_335 (O_335,N_14051,N_14271);
xnor UO_336 (O_336,N_14608,N_14789);
and UO_337 (O_337,N_14157,N_14441);
or UO_338 (O_338,N_14278,N_14066);
nand UO_339 (O_339,N_14949,N_14069);
nand UO_340 (O_340,N_14041,N_14198);
xnor UO_341 (O_341,N_14335,N_14502);
nor UO_342 (O_342,N_14462,N_14457);
nor UO_343 (O_343,N_14896,N_14557);
nor UO_344 (O_344,N_14765,N_14467);
and UO_345 (O_345,N_14680,N_14252);
nand UO_346 (O_346,N_14732,N_14088);
nand UO_347 (O_347,N_14123,N_14596);
xor UO_348 (O_348,N_14678,N_14940);
or UO_349 (O_349,N_14498,N_14097);
nand UO_350 (O_350,N_14644,N_14820);
nor UO_351 (O_351,N_14849,N_14672);
or UO_352 (O_352,N_14686,N_14378);
nor UO_353 (O_353,N_14796,N_14140);
nand UO_354 (O_354,N_14500,N_14333);
xor UO_355 (O_355,N_14779,N_14223);
nand UO_356 (O_356,N_14192,N_14694);
nor UO_357 (O_357,N_14880,N_14115);
nand UO_358 (O_358,N_14693,N_14296);
nand UO_359 (O_359,N_14797,N_14953);
or UO_360 (O_360,N_14701,N_14994);
nor UO_361 (O_361,N_14039,N_14658);
nor UO_362 (O_362,N_14633,N_14840);
nor UO_363 (O_363,N_14092,N_14020);
nor UO_364 (O_364,N_14952,N_14913);
nand UO_365 (O_365,N_14078,N_14478);
or UO_366 (O_366,N_14852,N_14788);
xnor UO_367 (O_367,N_14110,N_14976);
nand UO_368 (O_368,N_14615,N_14889);
xnor UO_369 (O_369,N_14401,N_14867);
and UO_370 (O_370,N_14322,N_14364);
or UO_371 (O_371,N_14716,N_14709);
xnor UO_372 (O_372,N_14717,N_14055);
or UO_373 (O_373,N_14938,N_14031);
and UO_374 (O_374,N_14555,N_14472);
nand UO_375 (O_375,N_14444,N_14089);
nand UO_376 (O_376,N_14605,N_14134);
xnor UO_377 (O_377,N_14315,N_14893);
nor UO_378 (O_378,N_14661,N_14598);
nor UO_379 (O_379,N_14329,N_14996);
nor UO_380 (O_380,N_14560,N_14411);
nor UO_381 (O_381,N_14866,N_14260);
or UO_382 (O_382,N_14629,N_14890);
xor UO_383 (O_383,N_14884,N_14239);
nand UO_384 (O_384,N_14689,N_14480);
nor UO_385 (O_385,N_14808,N_14572);
and UO_386 (O_386,N_14403,N_14662);
nor UO_387 (O_387,N_14046,N_14346);
xnor UO_388 (O_388,N_14453,N_14460);
or UO_389 (O_389,N_14757,N_14521);
nor UO_390 (O_390,N_14164,N_14264);
and UO_391 (O_391,N_14212,N_14091);
nor UO_392 (O_392,N_14098,N_14259);
or UO_393 (O_393,N_14923,N_14471);
nand UO_394 (O_394,N_14591,N_14503);
nor UO_395 (O_395,N_14573,N_14301);
nand UO_396 (O_396,N_14299,N_14815);
xor UO_397 (O_397,N_14670,N_14613);
or UO_398 (O_398,N_14008,N_14163);
nor UO_399 (O_399,N_14564,N_14435);
xor UO_400 (O_400,N_14627,N_14093);
or UO_401 (O_401,N_14486,N_14381);
nand UO_402 (O_402,N_14762,N_14948);
and UO_403 (O_403,N_14616,N_14445);
nor UO_404 (O_404,N_14711,N_14959);
or UO_405 (O_405,N_14394,N_14565);
nor UO_406 (O_406,N_14833,N_14556);
nor UO_407 (O_407,N_14951,N_14060);
or UO_408 (O_408,N_14090,N_14590);
nor UO_409 (O_409,N_14253,N_14321);
or UO_410 (O_410,N_14839,N_14375);
and UO_411 (O_411,N_14561,N_14631);
or UO_412 (O_412,N_14187,N_14936);
nand UO_413 (O_413,N_14248,N_14798);
or UO_414 (O_414,N_14247,N_14420);
or UO_415 (O_415,N_14971,N_14294);
xnor UO_416 (O_416,N_14536,N_14652);
and UO_417 (O_417,N_14416,N_14424);
nand UO_418 (O_418,N_14328,N_14310);
or UO_419 (O_419,N_14126,N_14958);
nor UO_420 (O_420,N_14581,N_14035);
and UO_421 (O_421,N_14466,N_14463);
xor UO_422 (O_422,N_14399,N_14783);
and UO_423 (O_423,N_14935,N_14413);
nand UO_424 (O_424,N_14229,N_14777);
nor UO_425 (O_425,N_14063,N_14634);
xnor UO_426 (O_426,N_14583,N_14176);
or UO_427 (O_427,N_14507,N_14873);
nor UO_428 (O_428,N_14057,N_14186);
nor UO_429 (O_429,N_14146,N_14476);
nand UO_430 (O_430,N_14195,N_14642);
or UO_431 (O_431,N_14459,N_14120);
and UO_432 (O_432,N_14183,N_14167);
nor UO_433 (O_433,N_14909,N_14961);
nand UO_434 (O_434,N_14675,N_14010);
nor UO_435 (O_435,N_14119,N_14955);
xor UO_436 (O_436,N_14130,N_14545);
nand UO_437 (O_437,N_14841,N_14257);
and UO_438 (O_438,N_14382,N_14117);
or UO_439 (O_439,N_14231,N_14440);
or UO_440 (O_440,N_14201,N_14821);
and UO_441 (O_441,N_14269,N_14080);
and UO_442 (O_442,N_14341,N_14995);
and UO_443 (O_443,N_14418,N_14842);
and UO_444 (O_444,N_14895,N_14794);
nand UO_445 (O_445,N_14256,N_14992);
nand UO_446 (O_446,N_14604,N_14434);
xor UO_447 (O_447,N_14065,N_14443);
nor UO_448 (O_448,N_14230,N_14715);
and UO_449 (O_449,N_14828,N_14647);
xnor UO_450 (O_450,N_14645,N_14863);
and UO_451 (O_451,N_14358,N_14576);
or UO_452 (O_452,N_14283,N_14524);
or UO_453 (O_453,N_14442,N_14638);
nor UO_454 (O_454,N_14113,N_14469);
and UO_455 (O_455,N_14003,N_14141);
nand UO_456 (O_456,N_14865,N_14708);
xnor UO_457 (O_457,N_14077,N_14054);
nor UO_458 (O_458,N_14419,N_14519);
nand UO_459 (O_459,N_14882,N_14042);
or UO_460 (O_460,N_14240,N_14415);
and UO_461 (O_461,N_14968,N_14282);
and UO_462 (O_462,N_14165,N_14334);
nand UO_463 (O_463,N_14816,N_14850);
nand UO_464 (O_464,N_14308,N_14879);
xor UO_465 (O_465,N_14837,N_14332);
nand UO_466 (O_466,N_14826,N_14387);
nor UO_467 (O_467,N_14314,N_14687);
xnor UO_468 (O_468,N_14342,N_14437);
nand UO_469 (O_469,N_14755,N_14393);
xnor UO_470 (O_470,N_14331,N_14125);
and UO_471 (O_471,N_14905,N_14292);
nand UO_472 (O_472,N_14725,N_14429);
xnor UO_473 (O_473,N_14285,N_14669);
xnor UO_474 (O_474,N_14786,N_14772);
and UO_475 (O_475,N_14760,N_14404);
nor UO_476 (O_476,N_14753,N_14526);
xor UO_477 (O_477,N_14514,N_14659);
xnor UO_478 (O_478,N_14361,N_14617);
xnor UO_479 (O_479,N_14817,N_14128);
xor UO_480 (O_480,N_14084,N_14246);
and UO_481 (O_481,N_14142,N_14226);
nand UO_482 (O_482,N_14611,N_14567);
xnor UO_483 (O_483,N_14921,N_14719);
xor UO_484 (O_484,N_14883,N_14568);
nor UO_485 (O_485,N_14086,N_14161);
or UO_486 (O_486,N_14217,N_14984);
nand UO_487 (O_487,N_14184,N_14588);
and UO_488 (O_488,N_14114,N_14518);
nor UO_489 (O_489,N_14028,N_14122);
and UO_490 (O_490,N_14614,N_14395);
or UO_491 (O_491,N_14803,N_14910);
nor UO_492 (O_492,N_14152,N_14506);
nand UO_493 (O_493,N_14104,N_14107);
nand UO_494 (O_494,N_14071,N_14272);
xor UO_495 (O_495,N_14390,N_14970);
nand UO_496 (O_496,N_14848,N_14191);
nor UO_497 (O_497,N_14881,N_14464);
and UO_498 (O_498,N_14855,N_14932);
and UO_499 (O_499,N_14592,N_14911);
nand UO_500 (O_500,N_14376,N_14641);
nor UO_501 (O_501,N_14618,N_14944);
nor UO_502 (O_502,N_14446,N_14221);
xor UO_503 (O_503,N_14580,N_14970);
or UO_504 (O_504,N_14643,N_14826);
nor UO_505 (O_505,N_14311,N_14045);
xor UO_506 (O_506,N_14853,N_14261);
and UO_507 (O_507,N_14645,N_14968);
xor UO_508 (O_508,N_14459,N_14142);
xor UO_509 (O_509,N_14924,N_14237);
xnor UO_510 (O_510,N_14771,N_14127);
nand UO_511 (O_511,N_14051,N_14187);
nand UO_512 (O_512,N_14565,N_14925);
nor UO_513 (O_513,N_14516,N_14521);
or UO_514 (O_514,N_14855,N_14730);
or UO_515 (O_515,N_14520,N_14952);
nor UO_516 (O_516,N_14052,N_14836);
xnor UO_517 (O_517,N_14379,N_14446);
nor UO_518 (O_518,N_14817,N_14402);
or UO_519 (O_519,N_14400,N_14671);
or UO_520 (O_520,N_14151,N_14131);
or UO_521 (O_521,N_14498,N_14136);
xor UO_522 (O_522,N_14720,N_14896);
and UO_523 (O_523,N_14887,N_14012);
nand UO_524 (O_524,N_14400,N_14252);
nor UO_525 (O_525,N_14545,N_14472);
or UO_526 (O_526,N_14599,N_14179);
or UO_527 (O_527,N_14029,N_14520);
xor UO_528 (O_528,N_14845,N_14912);
nand UO_529 (O_529,N_14498,N_14272);
xor UO_530 (O_530,N_14179,N_14567);
nand UO_531 (O_531,N_14685,N_14573);
nand UO_532 (O_532,N_14752,N_14935);
nand UO_533 (O_533,N_14213,N_14939);
xor UO_534 (O_534,N_14596,N_14762);
or UO_535 (O_535,N_14901,N_14196);
nor UO_536 (O_536,N_14159,N_14026);
and UO_537 (O_537,N_14487,N_14240);
and UO_538 (O_538,N_14447,N_14682);
nand UO_539 (O_539,N_14334,N_14272);
nand UO_540 (O_540,N_14377,N_14521);
xor UO_541 (O_541,N_14125,N_14615);
nand UO_542 (O_542,N_14632,N_14538);
nand UO_543 (O_543,N_14984,N_14465);
nor UO_544 (O_544,N_14795,N_14214);
nor UO_545 (O_545,N_14491,N_14091);
nand UO_546 (O_546,N_14451,N_14393);
xnor UO_547 (O_547,N_14907,N_14737);
nor UO_548 (O_548,N_14263,N_14615);
nand UO_549 (O_549,N_14403,N_14172);
xor UO_550 (O_550,N_14564,N_14699);
and UO_551 (O_551,N_14219,N_14268);
nor UO_552 (O_552,N_14555,N_14185);
or UO_553 (O_553,N_14705,N_14452);
and UO_554 (O_554,N_14918,N_14072);
nand UO_555 (O_555,N_14811,N_14965);
nor UO_556 (O_556,N_14476,N_14819);
xor UO_557 (O_557,N_14335,N_14284);
or UO_558 (O_558,N_14226,N_14483);
nand UO_559 (O_559,N_14530,N_14077);
nand UO_560 (O_560,N_14097,N_14995);
nand UO_561 (O_561,N_14325,N_14420);
or UO_562 (O_562,N_14590,N_14695);
xor UO_563 (O_563,N_14340,N_14012);
or UO_564 (O_564,N_14048,N_14359);
nor UO_565 (O_565,N_14703,N_14074);
and UO_566 (O_566,N_14135,N_14254);
nand UO_567 (O_567,N_14091,N_14431);
nand UO_568 (O_568,N_14710,N_14378);
or UO_569 (O_569,N_14231,N_14611);
nand UO_570 (O_570,N_14705,N_14225);
nor UO_571 (O_571,N_14729,N_14621);
and UO_572 (O_572,N_14034,N_14248);
xnor UO_573 (O_573,N_14072,N_14854);
or UO_574 (O_574,N_14719,N_14873);
or UO_575 (O_575,N_14052,N_14694);
and UO_576 (O_576,N_14991,N_14988);
xor UO_577 (O_577,N_14344,N_14916);
and UO_578 (O_578,N_14291,N_14635);
and UO_579 (O_579,N_14717,N_14555);
xnor UO_580 (O_580,N_14725,N_14559);
and UO_581 (O_581,N_14813,N_14761);
xnor UO_582 (O_582,N_14163,N_14269);
and UO_583 (O_583,N_14711,N_14568);
nor UO_584 (O_584,N_14326,N_14105);
or UO_585 (O_585,N_14982,N_14596);
nor UO_586 (O_586,N_14118,N_14180);
or UO_587 (O_587,N_14242,N_14223);
or UO_588 (O_588,N_14489,N_14763);
xnor UO_589 (O_589,N_14670,N_14432);
nand UO_590 (O_590,N_14045,N_14481);
nand UO_591 (O_591,N_14760,N_14464);
nand UO_592 (O_592,N_14287,N_14384);
nand UO_593 (O_593,N_14972,N_14913);
or UO_594 (O_594,N_14809,N_14313);
xor UO_595 (O_595,N_14237,N_14483);
nand UO_596 (O_596,N_14851,N_14728);
and UO_597 (O_597,N_14033,N_14870);
xnor UO_598 (O_598,N_14664,N_14862);
xnor UO_599 (O_599,N_14948,N_14621);
or UO_600 (O_600,N_14151,N_14398);
nand UO_601 (O_601,N_14880,N_14702);
and UO_602 (O_602,N_14710,N_14239);
and UO_603 (O_603,N_14360,N_14242);
xor UO_604 (O_604,N_14599,N_14748);
nor UO_605 (O_605,N_14826,N_14949);
nor UO_606 (O_606,N_14582,N_14391);
nand UO_607 (O_607,N_14348,N_14283);
and UO_608 (O_608,N_14952,N_14644);
nand UO_609 (O_609,N_14476,N_14247);
nor UO_610 (O_610,N_14399,N_14987);
and UO_611 (O_611,N_14113,N_14082);
and UO_612 (O_612,N_14430,N_14154);
and UO_613 (O_613,N_14278,N_14204);
xnor UO_614 (O_614,N_14926,N_14182);
nor UO_615 (O_615,N_14200,N_14831);
and UO_616 (O_616,N_14402,N_14606);
nand UO_617 (O_617,N_14053,N_14145);
xor UO_618 (O_618,N_14053,N_14165);
and UO_619 (O_619,N_14815,N_14074);
or UO_620 (O_620,N_14940,N_14306);
nand UO_621 (O_621,N_14626,N_14599);
xnor UO_622 (O_622,N_14668,N_14448);
nor UO_623 (O_623,N_14997,N_14089);
or UO_624 (O_624,N_14514,N_14605);
or UO_625 (O_625,N_14010,N_14189);
nor UO_626 (O_626,N_14405,N_14395);
and UO_627 (O_627,N_14383,N_14367);
or UO_628 (O_628,N_14100,N_14954);
or UO_629 (O_629,N_14401,N_14283);
and UO_630 (O_630,N_14682,N_14925);
or UO_631 (O_631,N_14215,N_14516);
xnor UO_632 (O_632,N_14624,N_14281);
or UO_633 (O_633,N_14155,N_14539);
or UO_634 (O_634,N_14807,N_14490);
and UO_635 (O_635,N_14489,N_14513);
xnor UO_636 (O_636,N_14714,N_14320);
or UO_637 (O_637,N_14880,N_14261);
nor UO_638 (O_638,N_14491,N_14197);
nor UO_639 (O_639,N_14589,N_14299);
and UO_640 (O_640,N_14831,N_14080);
nor UO_641 (O_641,N_14944,N_14726);
nor UO_642 (O_642,N_14506,N_14793);
nor UO_643 (O_643,N_14209,N_14522);
xor UO_644 (O_644,N_14315,N_14801);
xor UO_645 (O_645,N_14215,N_14213);
nand UO_646 (O_646,N_14095,N_14766);
and UO_647 (O_647,N_14344,N_14673);
xnor UO_648 (O_648,N_14743,N_14212);
nand UO_649 (O_649,N_14670,N_14833);
xor UO_650 (O_650,N_14737,N_14531);
nor UO_651 (O_651,N_14773,N_14344);
nand UO_652 (O_652,N_14940,N_14774);
xnor UO_653 (O_653,N_14026,N_14906);
nand UO_654 (O_654,N_14602,N_14589);
and UO_655 (O_655,N_14949,N_14166);
nand UO_656 (O_656,N_14187,N_14850);
and UO_657 (O_657,N_14517,N_14753);
xor UO_658 (O_658,N_14981,N_14110);
nor UO_659 (O_659,N_14331,N_14857);
nand UO_660 (O_660,N_14802,N_14694);
nand UO_661 (O_661,N_14386,N_14045);
nor UO_662 (O_662,N_14897,N_14278);
xor UO_663 (O_663,N_14628,N_14075);
nand UO_664 (O_664,N_14892,N_14113);
xor UO_665 (O_665,N_14984,N_14127);
nand UO_666 (O_666,N_14280,N_14176);
or UO_667 (O_667,N_14912,N_14178);
nand UO_668 (O_668,N_14998,N_14895);
xor UO_669 (O_669,N_14799,N_14108);
nand UO_670 (O_670,N_14786,N_14631);
or UO_671 (O_671,N_14263,N_14246);
or UO_672 (O_672,N_14301,N_14729);
nand UO_673 (O_673,N_14719,N_14436);
xnor UO_674 (O_674,N_14918,N_14463);
and UO_675 (O_675,N_14158,N_14744);
nor UO_676 (O_676,N_14314,N_14125);
nor UO_677 (O_677,N_14417,N_14128);
or UO_678 (O_678,N_14883,N_14305);
or UO_679 (O_679,N_14866,N_14537);
xor UO_680 (O_680,N_14938,N_14214);
xnor UO_681 (O_681,N_14356,N_14744);
nand UO_682 (O_682,N_14762,N_14379);
nor UO_683 (O_683,N_14492,N_14717);
or UO_684 (O_684,N_14876,N_14994);
and UO_685 (O_685,N_14699,N_14543);
xnor UO_686 (O_686,N_14865,N_14864);
or UO_687 (O_687,N_14910,N_14044);
and UO_688 (O_688,N_14869,N_14382);
nor UO_689 (O_689,N_14797,N_14781);
or UO_690 (O_690,N_14904,N_14677);
or UO_691 (O_691,N_14355,N_14081);
and UO_692 (O_692,N_14456,N_14759);
nand UO_693 (O_693,N_14367,N_14597);
nand UO_694 (O_694,N_14566,N_14844);
and UO_695 (O_695,N_14503,N_14489);
xor UO_696 (O_696,N_14945,N_14625);
and UO_697 (O_697,N_14331,N_14804);
xor UO_698 (O_698,N_14958,N_14835);
and UO_699 (O_699,N_14545,N_14674);
and UO_700 (O_700,N_14072,N_14943);
and UO_701 (O_701,N_14623,N_14038);
and UO_702 (O_702,N_14744,N_14619);
and UO_703 (O_703,N_14088,N_14059);
xnor UO_704 (O_704,N_14997,N_14571);
nor UO_705 (O_705,N_14306,N_14894);
and UO_706 (O_706,N_14766,N_14940);
xor UO_707 (O_707,N_14853,N_14341);
xor UO_708 (O_708,N_14305,N_14214);
or UO_709 (O_709,N_14300,N_14315);
and UO_710 (O_710,N_14648,N_14178);
or UO_711 (O_711,N_14282,N_14448);
xnor UO_712 (O_712,N_14570,N_14617);
nand UO_713 (O_713,N_14144,N_14199);
xor UO_714 (O_714,N_14156,N_14755);
xor UO_715 (O_715,N_14041,N_14858);
nand UO_716 (O_716,N_14432,N_14550);
or UO_717 (O_717,N_14555,N_14388);
nor UO_718 (O_718,N_14231,N_14401);
or UO_719 (O_719,N_14609,N_14028);
nand UO_720 (O_720,N_14369,N_14034);
or UO_721 (O_721,N_14745,N_14504);
nor UO_722 (O_722,N_14744,N_14013);
nor UO_723 (O_723,N_14189,N_14923);
or UO_724 (O_724,N_14995,N_14532);
xnor UO_725 (O_725,N_14957,N_14746);
xnor UO_726 (O_726,N_14321,N_14429);
nor UO_727 (O_727,N_14221,N_14977);
or UO_728 (O_728,N_14661,N_14784);
or UO_729 (O_729,N_14220,N_14962);
or UO_730 (O_730,N_14066,N_14926);
and UO_731 (O_731,N_14169,N_14171);
nand UO_732 (O_732,N_14247,N_14248);
xor UO_733 (O_733,N_14353,N_14626);
xnor UO_734 (O_734,N_14635,N_14654);
xor UO_735 (O_735,N_14547,N_14590);
nor UO_736 (O_736,N_14945,N_14373);
nand UO_737 (O_737,N_14552,N_14479);
or UO_738 (O_738,N_14860,N_14791);
nor UO_739 (O_739,N_14022,N_14840);
nor UO_740 (O_740,N_14577,N_14139);
nor UO_741 (O_741,N_14717,N_14512);
nor UO_742 (O_742,N_14376,N_14604);
or UO_743 (O_743,N_14640,N_14801);
nand UO_744 (O_744,N_14879,N_14473);
xnor UO_745 (O_745,N_14725,N_14827);
or UO_746 (O_746,N_14121,N_14781);
or UO_747 (O_747,N_14834,N_14401);
or UO_748 (O_748,N_14607,N_14644);
and UO_749 (O_749,N_14488,N_14821);
nand UO_750 (O_750,N_14181,N_14429);
xnor UO_751 (O_751,N_14034,N_14867);
nand UO_752 (O_752,N_14489,N_14648);
or UO_753 (O_753,N_14489,N_14983);
or UO_754 (O_754,N_14079,N_14381);
nand UO_755 (O_755,N_14637,N_14231);
nand UO_756 (O_756,N_14548,N_14230);
or UO_757 (O_757,N_14686,N_14148);
and UO_758 (O_758,N_14175,N_14297);
or UO_759 (O_759,N_14179,N_14683);
and UO_760 (O_760,N_14109,N_14321);
and UO_761 (O_761,N_14025,N_14518);
nor UO_762 (O_762,N_14754,N_14806);
xor UO_763 (O_763,N_14002,N_14326);
and UO_764 (O_764,N_14041,N_14993);
nand UO_765 (O_765,N_14617,N_14907);
or UO_766 (O_766,N_14587,N_14461);
and UO_767 (O_767,N_14245,N_14483);
or UO_768 (O_768,N_14582,N_14765);
nand UO_769 (O_769,N_14406,N_14365);
or UO_770 (O_770,N_14631,N_14215);
and UO_771 (O_771,N_14181,N_14368);
or UO_772 (O_772,N_14770,N_14246);
xnor UO_773 (O_773,N_14108,N_14227);
nand UO_774 (O_774,N_14811,N_14412);
nand UO_775 (O_775,N_14484,N_14292);
nand UO_776 (O_776,N_14151,N_14132);
nor UO_777 (O_777,N_14520,N_14643);
and UO_778 (O_778,N_14005,N_14210);
nor UO_779 (O_779,N_14161,N_14699);
nor UO_780 (O_780,N_14875,N_14438);
nor UO_781 (O_781,N_14366,N_14361);
and UO_782 (O_782,N_14641,N_14549);
and UO_783 (O_783,N_14540,N_14806);
xnor UO_784 (O_784,N_14180,N_14625);
or UO_785 (O_785,N_14486,N_14603);
nor UO_786 (O_786,N_14856,N_14015);
nor UO_787 (O_787,N_14482,N_14165);
nand UO_788 (O_788,N_14374,N_14314);
or UO_789 (O_789,N_14078,N_14379);
xnor UO_790 (O_790,N_14069,N_14427);
nor UO_791 (O_791,N_14165,N_14509);
xnor UO_792 (O_792,N_14224,N_14854);
xor UO_793 (O_793,N_14349,N_14861);
nor UO_794 (O_794,N_14425,N_14057);
nand UO_795 (O_795,N_14836,N_14096);
xnor UO_796 (O_796,N_14817,N_14745);
nand UO_797 (O_797,N_14729,N_14483);
and UO_798 (O_798,N_14079,N_14190);
xor UO_799 (O_799,N_14410,N_14525);
nand UO_800 (O_800,N_14249,N_14487);
nor UO_801 (O_801,N_14105,N_14346);
nand UO_802 (O_802,N_14011,N_14034);
or UO_803 (O_803,N_14571,N_14635);
nand UO_804 (O_804,N_14981,N_14994);
nor UO_805 (O_805,N_14727,N_14875);
nand UO_806 (O_806,N_14863,N_14256);
nand UO_807 (O_807,N_14315,N_14923);
and UO_808 (O_808,N_14675,N_14463);
or UO_809 (O_809,N_14435,N_14761);
and UO_810 (O_810,N_14882,N_14561);
nand UO_811 (O_811,N_14462,N_14052);
xor UO_812 (O_812,N_14463,N_14779);
or UO_813 (O_813,N_14138,N_14274);
or UO_814 (O_814,N_14669,N_14457);
or UO_815 (O_815,N_14788,N_14456);
nor UO_816 (O_816,N_14316,N_14713);
xor UO_817 (O_817,N_14412,N_14261);
or UO_818 (O_818,N_14837,N_14971);
xor UO_819 (O_819,N_14305,N_14532);
or UO_820 (O_820,N_14228,N_14807);
nand UO_821 (O_821,N_14893,N_14493);
nor UO_822 (O_822,N_14255,N_14380);
nand UO_823 (O_823,N_14274,N_14607);
nor UO_824 (O_824,N_14432,N_14316);
nand UO_825 (O_825,N_14790,N_14008);
or UO_826 (O_826,N_14812,N_14274);
nor UO_827 (O_827,N_14531,N_14054);
xnor UO_828 (O_828,N_14401,N_14247);
and UO_829 (O_829,N_14143,N_14632);
and UO_830 (O_830,N_14069,N_14780);
and UO_831 (O_831,N_14699,N_14656);
or UO_832 (O_832,N_14849,N_14548);
nor UO_833 (O_833,N_14833,N_14735);
and UO_834 (O_834,N_14157,N_14181);
nor UO_835 (O_835,N_14047,N_14918);
or UO_836 (O_836,N_14724,N_14577);
nand UO_837 (O_837,N_14597,N_14221);
xnor UO_838 (O_838,N_14016,N_14352);
nand UO_839 (O_839,N_14550,N_14116);
nor UO_840 (O_840,N_14305,N_14284);
and UO_841 (O_841,N_14084,N_14937);
or UO_842 (O_842,N_14486,N_14392);
and UO_843 (O_843,N_14240,N_14715);
nor UO_844 (O_844,N_14027,N_14352);
and UO_845 (O_845,N_14007,N_14410);
xor UO_846 (O_846,N_14559,N_14530);
nor UO_847 (O_847,N_14824,N_14434);
or UO_848 (O_848,N_14942,N_14612);
nor UO_849 (O_849,N_14896,N_14109);
nor UO_850 (O_850,N_14658,N_14160);
nand UO_851 (O_851,N_14308,N_14223);
xnor UO_852 (O_852,N_14064,N_14537);
nand UO_853 (O_853,N_14778,N_14027);
and UO_854 (O_854,N_14002,N_14049);
and UO_855 (O_855,N_14725,N_14912);
and UO_856 (O_856,N_14457,N_14673);
xor UO_857 (O_857,N_14715,N_14965);
nand UO_858 (O_858,N_14846,N_14225);
or UO_859 (O_859,N_14790,N_14578);
or UO_860 (O_860,N_14381,N_14839);
xnor UO_861 (O_861,N_14632,N_14012);
or UO_862 (O_862,N_14013,N_14297);
nand UO_863 (O_863,N_14895,N_14182);
or UO_864 (O_864,N_14575,N_14169);
nand UO_865 (O_865,N_14904,N_14427);
xnor UO_866 (O_866,N_14018,N_14531);
or UO_867 (O_867,N_14273,N_14576);
nor UO_868 (O_868,N_14306,N_14001);
xnor UO_869 (O_869,N_14968,N_14414);
or UO_870 (O_870,N_14125,N_14887);
nor UO_871 (O_871,N_14938,N_14542);
nand UO_872 (O_872,N_14343,N_14008);
nand UO_873 (O_873,N_14991,N_14806);
nand UO_874 (O_874,N_14806,N_14642);
and UO_875 (O_875,N_14977,N_14997);
and UO_876 (O_876,N_14287,N_14551);
nor UO_877 (O_877,N_14047,N_14694);
nand UO_878 (O_878,N_14399,N_14344);
nand UO_879 (O_879,N_14697,N_14589);
or UO_880 (O_880,N_14829,N_14021);
and UO_881 (O_881,N_14683,N_14562);
nand UO_882 (O_882,N_14626,N_14369);
nor UO_883 (O_883,N_14812,N_14636);
nand UO_884 (O_884,N_14665,N_14852);
xor UO_885 (O_885,N_14915,N_14137);
nor UO_886 (O_886,N_14334,N_14734);
nor UO_887 (O_887,N_14358,N_14244);
and UO_888 (O_888,N_14641,N_14353);
or UO_889 (O_889,N_14359,N_14081);
and UO_890 (O_890,N_14351,N_14620);
nor UO_891 (O_891,N_14477,N_14390);
nand UO_892 (O_892,N_14636,N_14736);
xor UO_893 (O_893,N_14694,N_14722);
nor UO_894 (O_894,N_14300,N_14589);
xnor UO_895 (O_895,N_14904,N_14133);
and UO_896 (O_896,N_14468,N_14920);
nor UO_897 (O_897,N_14389,N_14011);
nand UO_898 (O_898,N_14986,N_14153);
xnor UO_899 (O_899,N_14327,N_14050);
nand UO_900 (O_900,N_14048,N_14666);
and UO_901 (O_901,N_14493,N_14564);
nand UO_902 (O_902,N_14806,N_14465);
and UO_903 (O_903,N_14514,N_14267);
and UO_904 (O_904,N_14776,N_14795);
or UO_905 (O_905,N_14958,N_14280);
and UO_906 (O_906,N_14115,N_14594);
or UO_907 (O_907,N_14967,N_14788);
nor UO_908 (O_908,N_14563,N_14744);
and UO_909 (O_909,N_14708,N_14264);
or UO_910 (O_910,N_14627,N_14279);
and UO_911 (O_911,N_14697,N_14075);
nor UO_912 (O_912,N_14259,N_14573);
nand UO_913 (O_913,N_14856,N_14919);
and UO_914 (O_914,N_14623,N_14639);
nand UO_915 (O_915,N_14544,N_14823);
xor UO_916 (O_916,N_14269,N_14464);
or UO_917 (O_917,N_14620,N_14974);
or UO_918 (O_918,N_14545,N_14032);
xor UO_919 (O_919,N_14834,N_14721);
nand UO_920 (O_920,N_14534,N_14362);
xor UO_921 (O_921,N_14445,N_14099);
and UO_922 (O_922,N_14564,N_14048);
and UO_923 (O_923,N_14265,N_14882);
xnor UO_924 (O_924,N_14929,N_14748);
xor UO_925 (O_925,N_14328,N_14493);
or UO_926 (O_926,N_14214,N_14285);
xor UO_927 (O_927,N_14743,N_14419);
xnor UO_928 (O_928,N_14809,N_14324);
nor UO_929 (O_929,N_14778,N_14000);
nand UO_930 (O_930,N_14489,N_14974);
and UO_931 (O_931,N_14939,N_14122);
xor UO_932 (O_932,N_14415,N_14483);
xor UO_933 (O_933,N_14419,N_14407);
and UO_934 (O_934,N_14507,N_14062);
nor UO_935 (O_935,N_14027,N_14126);
and UO_936 (O_936,N_14422,N_14359);
and UO_937 (O_937,N_14859,N_14323);
nor UO_938 (O_938,N_14865,N_14196);
nand UO_939 (O_939,N_14464,N_14214);
xnor UO_940 (O_940,N_14705,N_14322);
or UO_941 (O_941,N_14017,N_14967);
and UO_942 (O_942,N_14769,N_14547);
xnor UO_943 (O_943,N_14421,N_14816);
nand UO_944 (O_944,N_14569,N_14542);
and UO_945 (O_945,N_14605,N_14748);
or UO_946 (O_946,N_14738,N_14547);
nor UO_947 (O_947,N_14276,N_14093);
nand UO_948 (O_948,N_14388,N_14269);
or UO_949 (O_949,N_14504,N_14608);
nand UO_950 (O_950,N_14854,N_14828);
or UO_951 (O_951,N_14571,N_14901);
and UO_952 (O_952,N_14856,N_14054);
nor UO_953 (O_953,N_14974,N_14724);
nor UO_954 (O_954,N_14870,N_14490);
nor UO_955 (O_955,N_14541,N_14363);
and UO_956 (O_956,N_14219,N_14130);
and UO_957 (O_957,N_14299,N_14537);
nand UO_958 (O_958,N_14468,N_14672);
nor UO_959 (O_959,N_14958,N_14557);
nor UO_960 (O_960,N_14943,N_14887);
and UO_961 (O_961,N_14510,N_14929);
xnor UO_962 (O_962,N_14050,N_14415);
or UO_963 (O_963,N_14108,N_14943);
nor UO_964 (O_964,N_14293,N_14520);
nor UO_965 (O_965,N_14032,N_14675);
or UO_966 (O_966,N_14117,N_14230);
nand UO_967 (O_967,N_14966,N_14719);
or UO_968 (O_968,N_14578,N_14844);
nand UO_969 (O_969,N_14803,N_14993);
and UO_970 (O_970,N_14242,N_14979);
nor UO_971 (O_971,N_14391,N_14136);
nand UO_972 (O_972,N_14792,N_14000);
nor UO_973 (O_973,N_14138,N_14660);
or UO_974 (O_974,N_14693,N_14116);
and UO_975 (O_975,N_14741,N_14863);
nand UO_976 (O_976,N_14456,N_14588);
nor UO_977 (O_977,N_14485,N_14109);
xor UO_978 (O_978,N_14261,N_14770);
or UO_979 (O_979,N_14863,N_14173);
xnor UO_980 (O_980,N_14254,N_14553);
and UO_981 (O_981,N_14787,N_14780);
xor UO_982 (O_982,N_14368,N_14269);
and UO_983 (O_983,N_14923,N_14470);
nor UO_984 (O_984,N_14994,N_14519);
or UO_985 (O_985,N_14596,N_14427);
xor UO_986 (O_986,N_14582,N_14197);
xnor UO_987 (O_987,N_14226,N_14819);
and UO_988 (O_988,N_14879,N_14686);
nand UO_989 (O_989,N_14109,N_14252);
and UO_990 (O_990,N_14370,N_14685);
or UO_991 (O_991,N_14679,N_14402);
nor UO_992 (O_992,N_14703,N_14244);
and UO_993 (O_993,N_14469,N_14451);
and UO_994 (O_994,N_14362,N_14751);
or UO_995 (O_995,N_14322,N_14969);
nand UO_996 (O_996,N_14791,N_14470);
xor UO_997 (O_997,N_14945,N_14229);
nand UO_998 (O_998,N_14115,N_14791);
and UO_999 (O_999,N_14478,N_14440);
nand UO_1000 (O_1000,N_14817,N_14502);
xnor UO_1001 (O_1001,N_14704,N_14014);
nand UO_1002 (O_1002,N_14385,N_14524);
or UO_1003 (O_1003,N_14330,N_14575);
nand UO_1004 (O_1004,N_14086,N_14028);
or UO_1005 (O_1005,N_14425,N_14744);
xor UO_1006 (O_1006,N_14543,N_14301);
nor UO_1007 (O_1007,N_14978,N_14862);
nor UO_1008 (O_1008,N_14673,N_14265);
and UO_1009 (O_1009,N_14108,N_14860);
nand UO_1010 (O_1010,N_14997,N_14348);
and UO_1011 (O_1011,N_14346,N_14861);
nand UO_1012 (O_1012,N_14203,N_14801);
xor UO_1013 (O_1013,N_14437,N_14578);
nor UO_1014 (O_1014,N_14044,N_14094);
and UO_1015 (O_1015,N_14698,N_14458);
xor UO_1016 (O_1016,N_14102,N_14619);
nor UO_1017 (O_1017,N_14550,N_14918);
or UO_1018 (O_1018,N_14174,N_14976);
nor UO_1019 (O_1019,N_14598,N_14089);
nor UO_1020 (O_1020,N_14374,N_14768);
nor UO_1021 (O_1021,N_14376,N_14152);
xnor UO_1022 (O_1022,N_14447,N_14303);
or UO_1023 (O_1023,N_14313,N_14353);
and UO_1024 (O_1024,N_14209,N_14396);
or UO_1025 (O_1025,N_14261,N_14082);
nand UO_1026 (O_1026,N_14143,N_14567);
nor UO_1027 (O_1027,N_14973,N_14346);
nor UO_1028 (O_1028,N_14080,N_14587);
nor UO_1029 (O_1029,N_14532,N_14803);
nor UO_1030 (O_1030,N_14529,N_14488);
and UO_1031 (O_1031,N_14932,N_14759);
nor UO_1032 (O_1032,N_14472,N_14320);
nand UO_1033 (O_1033,N_14382,N_14276);
and UO_1034 (O_1034,N_14148,N_14303);
nand UO_1035 (O_1035,N_14618,N_14088);
xnor UO_1036 (O_1036,N_14505,N_14887);
xor UO_1037 (O_1037,N_14741,N_14723);
and UO_1038 (O_1038,N_14612,N_14688);
and UO_1039 (O_1039,N_14281,N_14914);
nor UO_1040 (O_1040,N_14873,N_14238);
or UO_1041 (O_1041,N_14635,N_14752);
nand UO_1042 (O_1042,N_14894,N_14889);
and UO_1043 (O_1043,N_14829,N_14071);
and UO_1044 (O_1044,N_14840,N_14898);
nor UO_1045 (O_1045,N_14298,N_14416);
nor UO_1046 (O_1046,N_14561,N_14253);
or UO_1047 (O_1047,N_14126,N_14035);
xnor UO_1048 (O_1048,N_14093,N_14077);
nor UO_1049 (O_1049,N_14325,N_14433);
and UO_1050 (O_1050,N_14110,N_14073);
and UO_1051 (O_1051,N_14248,N_14638);
nor UO_1052 (O_1052,N_14143,N_14247);
xnor UO_1053 (O_1053,N_14851,N_14580);
or UO_1054 (O_1054,N_14373,N_14155);
xnor UO_1055 (O_1055,N_14590,N_14027);
nor UO_1056 (O_1056,N_14879,N_14734);
nand UO_1057 (O_1057,N_14738,N_14500);
xor UO_1058 (O_1058,N_14882,N_14842);
and UO_1059 (O_1059,N_14587,N_14927);
nand UO_1060 (O_1060,N_14041,N_14482);
or UO_1061 (O_1061,N_14862,N_14520);
nor UO_1062 (O_1062,N_14199,N_14975);
xor UO_1063 (O_1063,N_14125,N_14780);
nand UO_1064 (O_1064,N_14651,N_14490);
or UO_1065 (O_1065,N_14805,N_14750);
or UO_1066 (O_1066,N_14903,N_14254);
or UO_1067 (O_1067,N_14646,N_14119);
nand UO_1068 (O_1068,N_14903,N_14572);
or UO_1069 (O_1069,N_14184,N_14806);
nand UO_1070 (O_1070,N_14310,N_14365);
or UO_1071 (O_1071,N_14587,N_14217);
xor UO_1072 (O_1072,N_14951,N_14992);
nor UO_1073 (O_1073,N_14239,N_14120);
or UO_1074 (O_1074,N_14440,N_14249);
xnor UO_1075 (O_1075,N_14616,N_14086);
nor UO_1076 (O_1076,N_14306,N_14254);
and UO_1077 (O_1077,N_14735,N_14785);
xor UO_1078 (O_1078,N_14300,N_14659);
xor UO_1079 (O_1079,N_14950,N_14499);
nand UO_1080 (O_1080,N_14457,N_14426);
and UO_1081 (O_1081,N_14052,N_14174);
or UO_1082 (O_1082,N_14798,N_14593);
nor UO_1083 (O_1083,N_14698,N_14831);
nand UO_1084 (O_1084,N_14290,N_14332);
nor UO_1085 (O_1085,N_14381,N_14571);
nand UO_1086 (O_1086,N_14971,N_14192);
nor UO_1087 (O_1087,N_14226,N_14728);
nand UO_1088 (O_1088,N_14286,N_14161);
xnor UO_1089 (O_1089,N_14049,N_14229);
xor UO_1090 (O_1090,N_14303,N_14605);
or UO_1091 (O_1091,N_14812,N_14236);
nor UO_1092 (O_1092,N_14047,N_14190);
nor UO_1093 (O_1093,N_14860,N_14926);
or UO_1094 (O_1094,N_14677,N_14509);
nand UO_1095 (O_1095,N_14918,N_14478);
xor UO_1096 (O_1096,N_14682,N_14886);
xor UO_1097 (O_1097,N_14350,N_14459);
nand UO_1098 (O_1098,N_14576,N_14144);
and UO_1099 (O_1099,N_14630,N_14521);
nand UO_1100 (O_1100,N_14285,N_14036);
xor UO_1101 (O_1101,N_14600,N_14877);
xor UO_1102 (O_1102,N_14607,N_14906);
xor UO_1103 (O_1103,N_14816,N_14574);
xor UO_1104 (O_1104,N_14041,N_14809);
xor UO_1105 (O_1105,N_14779,N_14437);
and UO_1106 (O_1106,N_14111,N_14042);
xnor UO_1107 (O_1107,N_14191,N_14086);
nand UO_1108 (O_1108,N_14834,N_14803);
or UO_1109 (O_1109,N_14619,N_14513);
and UO_1110 (O_1110,N_14956,N_14009);
nor UO_1111 (O_1111,N_14226,N_14767);
nor UO_1112 (O_1112,N_14872,N_14855);
xnor UO_1113 (O_1113,N_14338,N_14744);
nor UO_1114 (O_1114,N_14903,N_14267);
nor UO_1115 (O_1115,N_14335,N_14297);
or UO_1116 (O_1116,N_14999,N_14245);
nor UO_1117 (O_1117,N_14856,N_14346);
and UO_1118 (O_1118,N_14181,N_14738);
or UO_1119 (O_1119,N_14556,N_14324);
xnor UO_1120 (O_1120,N_14922,N_14311);
and UO_1121 (O_1121,N_14252,N_14255);
xor UO_1122 (O_1122,N_14569,N_14864);
xor UO_1123 (O_1123,N_14301,N_14981);
or UO_1124 (O_1124,N_14772,N_14210);
or UO_1125 (O_1125,N_14458,N_14175);
or UO_1126 (O_1126,N_14003,N_14780);
nor UO_1127 (O_1127,N_14395,N_14358);
and UO_1128 (O_1128,N_14854,N_14412);
nor UO_1129 (O_1129,N_14564,N_14459);
or UO_1130 (O_1130,N_14580,N_14249);
xor UO_1131 (O_1131,N_14032,N_14909);
and UO_1132 (O_1132,N_14169,N_14853);
and UO_1133 (O_1133,N_14683,N_14809);
xnor UO_1134 (O_1134,N_14686,N_14511);
or UO_1135 (O_1135,N_14542,N_14272);
nor UO_1136 (O_1136,N_14869,N_14513);
or UO_1137 (O_1137,N_14644,N_14673);
nor UO_1138 (O_1138,N_14654,N_14262);
nor UO_1139 (O_1139,N_14643,N_14214);
or UO_1140 (O_1140,N_14196,N_14132);
nor UO_1141 (O_1141,N_14203,N_14572);
xnor UO_1142 (O_1142,N_14335,N_14498);
or UO_1143 (O_1143,N_14777,N_14948);
xor UO_1144 (O_1144,N_14504,N_14310);
or UO_1145 (O_1145,N_14877,N_14053);
nor UO_1146 (O_1146,N_14337,N_14908);
nand UO_1147 (O_1147,N_14960,N_14579);
and UO_1148 (O_1148,N_14312,N_14150);
nor UO_1149 (O_1149,N_14762,N_14628);
or UO_1150 (O_1150,N_14704,N_14112);
nand UO_1151 (O_1151,N_14195,N_14440);
xor UO_1152 (O_1152,N_14266,N_14079);
nor UO_1153 (O_1153,N_14535,N_14396);
or UO_1154 (O_1154,N_14132,N_14536);
nor UO_1155 (O_1155,N_14654,N_14516);
xor UO_1156 (O_1156,N_14053,N_14624);
and UO_1157 (O_1157,N_14501,N_14342);
nor UO_1158 (O_1158,N_14104,N_14384);
and UO_1159 (O_1159,N_14077,N_14003);
nand UO_1160 (O_1160,N_14728,N_14844);
nand UO_1161 (O_1161,N_14441,N_14848);
and UO_1162 (O_1162,N_14689,N_14100);
nand UO_1163 (O_1163,N_14700,N_14347);
nor UO_1164 (O_1164,N_14270,N_14933);
and UO_1165 (O_1165,N_14147,N_14512);
and UO_1166 (O_1166,N_14386,N_14197);
nand UO_1167 (O_1167,N_14979,N_14228);
and UO_1168 (O_1168,N_14710,N_14853);
nor UO_1169 (O_1169,N_14883,N_14248);
or UO_1170 (O_1170,N_14830,N_14191);
and UO_1171 (O_1171,N_14471,N_14951);
nand UO_1172 (O_1172,N_14190,N_14049);
nor UO_1173 (O_1173,N_14334,N_14001);
nor UO_1174 (O_1174,N_14821,N_14121);
xnor UO_1175 (O_1175,N_14586,N_14646);
nor UO_1176 (O_1176,N_14926,N_14811);
and UO_1177 (O_1177,N_14033,N_14533);
nor UO_1178 (O_1178,N_14084,N_14916);
nor UO_1179 (O_1179,N_14699,N_14403);
and UO_1180 (O_1180,N_14496,N_14894);
or UO_1181 (O_1181,N_14009,N_14499);
nor UO_1182 (O_1182,N_14407,N_14124);
and UO_1183 (O_1183,N_14873,N_14534);
nand UO_1184 (O_1184,N_14273,N_14514);
nand UO_1185 (O_1185,N_14967,N_14592);
or UO_1186 (O_1186,N_14868,N_14234);
nor UO_1187 (O_1187,N_14528,N_14360);
nor UO_1188 (O_1188,N_14771,N_14332);
or UO_1189 (O_1189,N_14367,N_14692);
xnor UO_1190 (O_1190,N_14075,N_14078);
or UO_1191 (O_1191,N_14875,N_14674);
nor UO_1192 (O_1192,N_14834,N_14120);
or UO_1193 (O_1193,N_14291,N_14840);
xor UO_1194 (O_1194,N_14463,N_14843);
and UO_1195 (O_1195,N_14101,N_14095);
and UO_1196 (O_1196,N_14746,N_14126);
xnor UO_1197 (O_1197,N_14643,N_14409);
and UO_1198 (O_1198,N_14868,N_14248);
xnor UO_1199 (O_1199,N_14741,N_14243);
xor UO_1200 (O_1200,N_14742,N_14799);
xnor UO_1201 (O_1201,N_14749,N_14852);
and UO_1202 (O_1202,N_14892,N_14447);
and UO_1203 (O_1203,N_14115,N_14655);
nor UO_1204 (O_1204,N_14074,N_14304);
and UO_1205 (O_1205,N_14987,N_14077);
nand UO_1206 (O_1206,N_14560,N_14536);
nor UO_1207 (O_1207,N_14124,N_14000);
xor UO_1208 (O_1208,N_14133,N_14948);
xor UO_1209 (O_1209,N_14295,N_14805);
and UO_1210 (O_1210,N_14241,N_14377);
or UO_1211 (O_1211,N_14251,N_14759);
or UO_1212 (O_1212,N_14320,N_14615);
xnor UO_1213 (O_1213,N_14849,N_14439);
nor UO_1214 (O_1214,N_14100,N_14712);
xnor UO_1215 (O_1215,N_14409,N_14364);
or UO_1216 (O_1216,N_14126,N_14024);
nor UO_1217 (O_1217,N_14161,N_14946);
or UO_1218 (O_1218,N_14137,N_14070);
and UO_1219 (O_1219,N_14193,N_14492);
xnor UO_1220 (O_1220,N_14231,N_14240);
nor UO_1221 (O_1221,N_14760,N_14929);
or UO_1222 (O_1222,N_14508,N_14802);
or UO_1223 (O_1223,N_14185,N_14076);
nand UO_1224 (O_1224,N_14510,N_14110);
nand UO_1225 (O_1225,N_14768,N_14080);
or UO_1226 (O_1226,N_14939,N_14181);
nor UO_1227 (O_1227,N_14326,N_14550);
or UO_1228 (O_1228,N_14442,N_14906);
and UO_1229 (O_1229,N_14289,N_14729);
and UO_1230 (O_1230,N_14859,N_14804);
and UO_1231 (O_1231,N_14648,N_14082);
and UO_1232 (O_1232,N_14877,N_14552);
nor UO_1233 (O_1233,N_14125,N_14078);
and UO_1234 (O_1234,N_14664,N_14176);
nand UO_1235 (O_1235,N_14495,N_14918);
and UO_1236 (O_1236,N_14714,N_14733);
and UO_1237 (O_1237,N_14336,N_14708);
nand UO_1238 (O_1238,N_14256,N_14019);
or UO_1239 (O_1239,N_14963,N_14087);
or UO_1240 (O_1240,N_14515,N_14297);
and UO_1241 (O_1241,N_14122,N_14236);
and UO_1242 (O_1242,N_14935,N_14391);
and UO_1243 (O_1243,N_14207,N_14622);
nand UO_1244 (O_1244,N_14780,N_14577);
nand UO_1245 (O_1245,N_14958,N_14041);
and UO_1246 (O_1246,N_14977,N_14743);
and UO_1247 (O_1247,N_14685,N_14247);
nand UO_1248 (O_1248,N_14060,N_14869);
and UO_1249 (O_1249,N_14756,N_14360);
and UO_1250 (O_1250,N_14452,N_14897);
nor UO_1251 (O_1251,N_14253,N_14697);
nor UO_1252 (O_1252,N_14470,N_14822);
nor UO_1253 (O_1253,N_14078,N_14815);
nor UO_1254 (O_1254,N_14496,N_14999);
or UO_1255 (O_1255,N_14882,N_14832);
or UO_1256 (O_1256,N_14859,N_14739);
xor UO_1257 (O_1257,N_14285,N_14736);
nand UO_1258 (O_1258,N_14914,N_14530);
nand UO_1259 (O_1259,N_14008,N_14974);
nor UO_1260 (O_1260,N_14884,N_14921);
nor UO_1261 (O_1261,N_14491,N_14274);
nand UO_1262 (O_1262,N_14284,N_14836);
or UO_1263 (O_1263,N_14206,N_14968);
and UO_1264 (O_1264,N_14869,N_14006);
and UO_1265 (O_1265,N_14524,N_14748);
nor UO_1266 (O_1266,N_14690,N_14503);
nor UO_1267 (O_1267,N_14057,N_14518);
nand UO_1268 (O_1268,N_14266,N_14308);
nand UO_1269 (O_1269,N_14909,N_14506);
xnor UO_1270 (O_1270,N_14070,N_14605);
nand UO_1271 (O_1271,N_14306,N_14133);
xor UO_1272 (O_1272,N_14460,N_14833);
nor UO_1273 (O_1273,N_14941,N_14802);
and UO_1274 (O_1274,N_14837,N_14208);
xor UO_1275 (O_1275,N_14471,N_14377);
or UO_1276 (O_1276,N_14162,N_14775);
and UO_1277 (O_1277,N_14459,N_14964);
or UO_1278 (O_1278,N_14540,N_14719);
xor UO_1279 (O_1279,N_14000,N_14371);
xnor UO_1280 (O_1280,N_14199,N_14755);
and UO_1281 (O_1281,N_14909,N_14829);
nand UO_1282 (O_1282,N_14195,N_14847);
and UO_1283 (O_1283,N_14605,N_14551);
nor UO_1284 (O_1284,N_14882,N_14205);
nor UO_1285 (O_1285,N_14499,N_14187);
nand UO_1286 (O_1286,N_14191,N_14953);
and UO_1287 (O_1287,N_14629,N_14359);
nand UO_1288 (O_1288,N_14164,N_14380);
nor UO_1289 (O_1289,N_14586,N_14259);
nand UO_1290 (O_1290,N_14640,N_14957);
or UO_1291 (O_1291,N_14646,N_14078);
nor UO_1292 (O_1292,N_14879,N_14058);
and UO_1293 (O_1293,N_14959,N_14891);
nand UO_1294 (O_1294,N_14890,N_14223);
and UO_1295 (O_1295,N_14226,N_14604);
or UO_1296 (O_1296,N_14441,N_14223);
xnor UO_1297 (O_1297,N_14189,N_14292);
nor UO_1298 (O_1298,N_14416,N_14212);
nand UO_1299 (O_1299,N_14388,N_14065);
or UO_1300 (O_1300,N_14596,N_14750);
or UO_1301 (O_1301,N_14926,N_14994);
and UO_1302 (O_1302,N_14979,N_14918);
nor UO_1303 (O_1303,N_14563,N_14297);
or UO_1304 (O_1304,N_14941,N_14437);
and UO_1305 (O_1305,N_14897,N_14085);
nor UO_1306 (O_1306,N_14091,N_14755);
or UO_1307 (O_1307,N_14418,N_14308);
or UO_1308 (O_1308,N_14177,N_14228);
xnor UO_1309 (O_1309,N_14144,N_14706);
or UO_1310 (O_1310,N_14653,N_14535);
nand UO_1311 (O_1311,N_14735,N_14698);
and UO_1312 (O_1312,N_14542,N_14695);
xor UO_1313 (O_1313,N_14074,N_14684);
nor UO_1314 (O_1314,N_14710,N_14479);
nor UO_1315 (O_1315,N_14399,N_14362);
and UO_1316 (O_1316,N_14838,N_14670);
nand UO_1317 (O_1317,N_14883,N_14965);
nand UO_1318 (O_1318,N_14824,N_14400);
or UO_1319 (O_1319,N_14513,N_14158);
xor UO_1320 (O_1320,N_14763,N_14777);
or UO_1321 (O_1321,N_14324,N_14167);
nand UO_1322 (O_1322,N_14531,N_14425);
nor UO_1323 (O_1323,N_14415,N_14313);
nor UO_1324 (O_1324,N_14436,N_14954);
or UO_1325 (O_1325,N_14410,N_14438);
and UO_1326 (O_1326,N_14830,N_14331);
or UO_1327 (O_1327,N_14836,N_14490);
nor UO_1328 (O_1328,N_14089,N_14709);
or UO_1329 (O_1329,N_14269,N_14562);
or UO_1330 (O_1330,N_14975,N_14092);
and UO_1331 (O_1331,N_14358,N_14000);
or UO_1332 (O_1332,N_14078,N_14017);
nand UO_1333 (O_1333,N_14433,N_14832);
or UO_1334 (O_1334,N_14636,N_14848);
nand UO_1335 (O_1335,N_14823,N_14755);
nor UO_1336 (O_1336,N_14427,N_14365);
nor UO_1337 (O_1337,N_14005,N_14959);
nor UO_1338 (O_1338,N_14562,N_14807);
and UO_1339 (O_1339,N_14940,N_14037);
and UO_1340 (O_1340,N_14599,N_14245);
nor UO_1341 (O_1341,N_14601,N_14645);
and UO_1342 (O_1342,N_14166,N_14767);
xor UO_1343 (O_1343,N_14601,N_14995);
or UO_1344 (O_1344,N_14293,N_14765);
nand UO_1345 (O_1345,N_14803,N_14858);
xor UO_1346 (O_1346,N_14142,N_14739);
nand UO_1347 (O_1347,N_14187,N_14589);
or UO_1348 (O_1348,N_14735,N_14732);
or UO_1349 (O_1349,N_14782,N_14332);
or UO_1350 (O_1350,N_14820,N_14915);
or UO_1351 (O_1351,N_14752,N_14918);
and UO_1352 (O_1352,N_14046,N_14208);
or UO_1353 (O_1353,N_14536,N_14830);
xor UO_1354 (O_1354,N_14738,N_14877);
and UO_1355 (O_1355,N_14971,N_14533);
and UO_1356 (O_1356,N_14151,N_14702);
nand UO_1357 (O_1357,N_14955,N_14253);
and UO_1358 (O_1358,N_14353,N_14727);
or UO_1359 (O_1359,N_14945,N_14703);
or UO_1360 (O_1360,N_14273,N_14946);
xor UO_1361 (O_1361,N_14822,N_14537);
and UO_1362 (O_1362,N_14414,N_14259);
and UO_1363 (O_1363,N_14148,N_14972);
nor UO_1364 (O_1364,N_14870,N_14831);
xnor UO_1365 (O_1365,N_14315,N_14131);
and UO_1366 (O_1366,N_14969,N_14845);
xor UO_1367 (O_1367,N_14241,N_14454);
and UO_1368 (O_1368,N_14806,N_14429);
or UO_1369 (O_1369,N_14832,N_14065);
and UO_1370 (O_1370,N_14690,N_14435);
nand UO_1371 (O_1371,N_14328,N_14921);
nor UO_1372 (O_1372,N_14380,N_14212);
nand UO_1373 (O_1373,N_14431,N_14102);
xnor UO_1374 (O_1374,N_14344,N_14895);
nor UO_1375 (O_1375,N_14243,N_14115);
nor UO_1376 (O_1376,N_14350,N_14619);
or UO_1377 (O_1377,N_14665,N_14418);
xor UO_1378 (O_1378,N_14737,N_14860);
nand UO_1379 (O_1379,N_14430,N_14325);
nand UO_1380 (O_1380,N_14837,N_14438);
nor UO_1381 (O_1381,N_14452,N_14644);
nand UO_1382 (O_1382,N_14463,N_14089);
nor UO_1383 (O_1383,N_14694,N_14821);
nor UO_1384 (O_1384,N_14471,N_14480);
or UO_1385 (O_1385,N_14461,N_14223);
xor UO_1386 (O_1386,N_14793,N_14574);
or UO_1387 (O_1387,N_14520,N_14427);
or UO_1388 (O_1388,N_14063,N_14740);
xor UO_1389 (O_1389,N_14957,N_14510);
nand UO_1390 (O_1390,N_14744,N_14947);
nor UO_1391 (O_1391,N_14496,N_14218);
or UO_1392 (O_1392,N_14315,N_14610);
xor UO_1393 (O_1393,N_14523,N_14029);
nor UO_1394 (O_1394,N_14467,N_14222);
nand UO_1395 (O_1395,N_14169,N_14641);
xnor UO_1396 (O_1396,N_14534,N_14532);
and UO_1397 (O_1397,N_14036,N_14931);
and UO_1398 (O_1398,N_14399,N_14227);
xor UO_1399 (O_1399,N_14606,N_14158);
nor UO_1400 (O_1400,N_14477,N_14427);
nor UO_1401 (O_1401,N_14995,N_14474);
or UO_1402 (O_1402,N_14712,N_14809);
nor UO_1403 (O_1403,N_14336,N_14389);
nor UO_1404 (O_1404,N_14836,N_14568);
nand UO_1405 (O_1405,N_14060,N_14153);
nor UO_1406 (O_1406,N_14738,N_14399);
and UO_1407 (O_1407,N_14427,N_14225);
nor UO_1408 (O_1408,N_14284,N_14355);
nand UO_1409 (O_1409,N_14361,N_14689);
and UO_1410 (O_1410,N_14439,N_14326);
nand UO_1411 (O_1411,N_14782,N_14703);
nor UO_1412 (O_1412,N_14338,N_14856);
and UO_1413 (O_1413,N_14205,N_14706);
or UO_1414 (O_1414,N_14545,N_14348);
nor UO_1415 (O_1415,N_14990,N_14337);
nand UO_1416 (O_1416,N_14513,N_14453);
xor UO_1417 (O_1417,N_14307,N_14162);
and UO_1418 (O_1418,N_14482,N_14696);
and UO_1419 (O_1419,N_14690,N_14871);
nor UO_1420 (O_1420,N_14633,N_14475);
nor UO_1421 (O_1421,N_14664,N_14365);
nand UO_1422 (O_1422,N_14522,N_14682);
and UO_1423 (O_1423,N_14114,N_14446);
xor UO_1424 (O_1424,N_14986,N_14426);
or UO_1425 (O_1425,N_14488,N_14732);
and UO_1426 (O_1426,N_14758,N_14633);
nand UO_1427 (O_1427,N_14371,N_14500);
or UO_1428 (O_1428,N_14116,N_14742);
xor UO_1429 (O_1429,N_14056,N_14747);
nor UO_1430 (O_1430,N_14463,N_14526);
xor UO_1431 (O_1431,N_14549,N_14526);
nor UO_1432 (O_1432,N_14210,N_14773);
or UO_1433 (O_1433,N_14352,N_14643);
nor UO_1434 (O_1434,N_14356,N_14891);
xnor UO_1435 (O_1435,N_14009,N_14351);
or UO_1436 (O_1436,N_14819,N_14495);
xnor UO_1437 (O_1437,N_14363,N_14378);
or UO_1438 (O_1438,N_14933,N_14392);
xnor UO_1439 (O_1439,N_14396,N_14533);
nand UO_1440 (O_1440,N_14691,N_14636);
xor UO_1441 (O_1441,N_14349,N_14088);
nor UO_1442 (O_1442,N_14503,N_14060);
and UO_1443 (O_1443,N_14075,N_14040);
xor UO_1444 (O_1444,N_14513,N_14424);
xor UO_1445 (O_1445,N_14502,N_14212);
and UO_1446 (O_1446,N_14035,N_14610);
nor UO_1447 (O_1447,N_14982,N_14910);
nor UO_1448 (O_1448,N_14688,N_14420);
and UO_1449 (O_1449,N_14619,N_14273);
nor UO_1450 (O_1450,N_14046,N_14173);
xnor UO_1451 (O_1451,N_14010,N_14248);
and UO_1452 (O_1452,N_14295,N_14106);
nand UO_1453 (O_1453,N_14543,N_14115);
and UO_1454 (O_1454,N_14172,N_14382);
nor UO_1455 (O_1455,N_14276,N_14721);
and UO_1456 (O_1456,N_14746,N_14153);
and UO_1457 (O_1457,N_14024,N_14912);
or UO_1458 (O_1458,N_14376,N_14733);
and UO_1459 (O_1459,N_14922,N_14592);
nor UO_1460 (O_1460,N_14194,N_14942);
nand UO_1461 (O_1461,N_14804,N_14446);
nor UO_1462 (O_1462,N_14106,N_14828);
and UO_1463 (O_1463,N_14559,N_14874);
xor UO_1464 (O_1464,N_14433,N_14155);
xor UO_1465 (O_1465,N_14436,N_14483);
xnor UO_1466 (O_1466,N_14717,N_14676);
xnor UO_1467 (O_1467,N_14260,N_14057);
xor UO_1468 (O_1468,N_14014,N_14235);
or UO_1469 (O_1469,N_14438,N_14477);
nand UO_1470 (O_1470,N_14533,N_14211);
and UO_1471 (O_1471,N_14602,N_14663);
and UO_1472 (O_1472,N_14141,N_14580);
nor UO_1473 (O_1473,N_14326,N_14490);
or UO_1474 (O_1474,N_14406,N_14301);
nand UO_1475 (O_1475,N_14091,N_14095);
nor UO_1476 (O_1476,N_14573,N_14500);
nor UO_1477 (O_1477,N_14553,N_14701);
or UO_1478 (O_1478,N_14417,N_14681);
and UO_1479 (O_1479,N_14496,N_14335);
nand UO_1480 (O_1480,N_14735,N_14437);
nand UO_1481 (O_1481,N_14340,N_14326);
nor UO_1482 (O_1482,N_14645,N_14265);
nand UO_1483 (O_1483,N_14976,N_14812);
nor UO_1484 (O_1484,N_14806,N_14672);
nand UO_1485 (O_1485,N_14649,N_14345);
nand UO_1486 (O_1486,N_14266,N_14544);
or UO_1487 (O_1487,N_14042,N_14588);
or UO_1488 (O_1488,N_14965,N_14088);
xor UO_1489 (O_1489,N_14171,N_14794);
and UO_1490 (O_1490,N_14166,N_14354);
nor UO_1491 (O_1491,N_14666,N_14365);
nand UO_1492 (O_1492,N_14011,N_14923);
xnor UO_1493 (O_1493,N_14414,N_14379);
or UO_1494 (O_1494,N_14303,N_14282);
nor UO_1495 (O_1495,N_14763,N_14494);
or UO_1496 (O_1496,N_14669,N_14863);
nor UO_1497 (O_1497,N_14259,N_14520);
nand UO_1498 (O_1498,N_14575,N_14771);
nand UO_1499 (O_1499,N_14629,N_14030);
and UO_1500 (O_1500,N_14312,N_14250);
or UO_1501 (O_1501,N_14965,N_14723);
or UO_1502 (O_1502,N_14730,N_14790);
or UO_1503 (O_1503,N_14290,N_14026);
and UO_1504 (O_1504,N_14664,N_14368);
nor UO_1505 (O_1505,N_14202,N_14983);
nand UO_1506 (O_1506,N_14366,N_14935);
or UO_1507 (O_1507,N_14777,N_14652);
xor UO_1508 (O_1508,N_14875,N_14576);
or UO_1509 (O_1509,N_14695,N_14004);
xor UO_1510 (O_1510,N_14129,N_14252);
nand UO_1511 (O_1511,N_14429,N_14326);
nand UO_1512 (O_1512,N_14493,N_14977);
or UO_1513 (O_1513,N_14841,N_14554);
and UO_1514 (O_1514,N_14097,N_14136);
nand UO_1515 (O_1515,N_14376,N_14204);
and UO_1516 (O_1516,N_14201,N_14940);
and UO_1517 (O_1517,N_14654,N_14449);
xnor UO_1518 (O_1518,N_14527,N_14320);
and UO_1519 (O_1519,N_14924,N_14039);
and UO_1520 (O_1520,N_14967,N_14007);
xnor UO_1521 (O_1521,N_14143,N_14361);
nor UO_1522 (O_1522,N_14541,N_14636);
and UO_1523 (O_1523,N_14020,N_14504);
xnor UO_1524 (O_1524,N_14898,N_14755);
or UO_1525 (O_1525,N_14354,N_14720);
and UO_1526 (O_1526,N_14611,N_14627);
or UO_1527 (O_1527,N_14711,N_14031);
nand UO_1528 (O_1528,N_14471,N_14341);
nand UO_1529 (O_1529,N_14689,N_14795);
or UO_1530 (O_1530,N_14749,N_14229);
nand UO_1531 (O_1531,N_14370,N_14560);
and UO_1532 (O_1532,N_14461,N_14728);
and UO_1533 (O_1533,N_14183,N_14247);
nand UO_1534 (O_1534,N_14191,N_14995);
xor UO_1535 (O_1535,N_14032,N_14683);
nor UO_1536 (O_1536,N_14168,N_14793);
xor UO_1537 (O_1537,N_14902,N_14253);
and UO_1538 (O_1538,N_14428,N_14555);
and UO_1539 (O_1539,N_14817,N_14912);
xnor UO_1540 (O_1540,N_14984,N_14336);
xor UO_1541 (O_1541,N_14523,N_14236);
nand UO_1542 (O_1542,N_14118,N_14588);
and UO_1543 (O_1543,N_14695,N_14096);
or UO_1544 (O_1544,N_14214,N_14232);
nor UO_1545 (O_1545,N_14759,N_14173);
xor UO_1546 (O_1546,N_14840,N_14661);
or UO_1547 (O_1547,N_14923,N_14901);
or UO_1548 (O_1548,N_14126,N_14106);
nand UO_1549 (O_1549,N_14254,N_14539);
xor UO_1550 (O_1550,N_14134,N_14871);
and UO_1551 (O_1551,N_14124,N_14251);
xnor UO_1552 (O_1552,N_14823,N_14851);
nor UO_1553 (O_1553,N_14377,N_14253);
or UO_1554 (O_1554,N_14496,N_14098);
nor UO_1555 (O_1555,N_14562,N_14449);
or UO_1556 (O_1556,N_14829,N_14827);
and UO_1557 (O_1557,N_14094,N_14336);
xnor UO_1558 (O_1558,N_14125,N_14468);
nand UO_1559 (O_1559,N_14812,N_14467);
xnor UO_1560 (O_1560,N_14437,N_14457);
and UO_1561 (O_1561,N_14976,N_14911);
xnor UO_1562 (O_1562,N_14881,N_14645);
or UO_1563 (O_1563,N_14657,N_14955);
xor UO_1564 (O_1564,N_14196,N_14648);
and UO_1565 (O_1565,N_14800,N_14957);
nor UO_1566 (O_1566,N_14903,N_14753);
xnor UO_1567 (O_1567,N_14897,N_14550);
or UO_1568 (O_1568,N_14753,N_14547);
xor UO_1569 (O_1569,N_14891,N_14762);
nor UO_1570 (O_1570,N_14751,N_14616);
and UO_1571 (O_1571,N_14302,N_14222);
nand UO_1572 (O_1572,N_14205,N_14572);
nand UO_1573 (O_1573,N_14807,N_14944);
nor UO_1574 (O_1574,N_14897,N_14365);
nand UO_1575 (O_1575,N_14736,N_14136);
or UO_1576 (O_1576,N_14615,N_14403);
nand UO_1577 (O_1577,N_14135,N_14539);
nand UO_1578 (O_1578,N_14881,N_14622);
nand UO_1579 (O_1579,N_14670,N_14443);
or UO_1580 (O_1580,N_14049,N_14047);
and UO_1581 (O_1581,N_14443,N_14472);
xnor UO_1582 (O_1582,N_14151,N_14854);
nor UO_1583 (O_1583,N_14696,N_14318);
nor UO_1584 (O_1584,N_14569,N_14868);
nor UO_1585 (O_1585,N_14083,N_14440);
or UO_1586 (O_1586,N_14231,N_14579);
xor UO_1587 (O_1587,N_14926,N_14765);
or UO_1588 (O_1588,N_14919,N_14619);
or UO_1589 (O_1589,N_14204,N_14553);
xnor UO_1590 (O_1590,N_14371,N_14648);
xor UO_1591 (O_1591,N_14010,N_14184);
xnor UO_1592 (O_1592,N_14188,N_14692);
and UO_1593 (O_1593,N_14023,N_14473);
xor UO_1594 (O_1594,N_14812,N_14998);
nor UO_1595 (O_1595,N_14090,N_14252);
and UO_1596 (O_1596,N_14288,N_14169);
nand UO_1597 (O_1597,N_14193,N_14322);
or UO_1598 (O_1598,N_14636,N_14404);
or UO_1599 (O_1599,N_14392,N_14067);
nor UO_1600 (O_1600,N_14169,N_14689);
or UO_1601 (O_1601,N_14468,N_14958);
or UO_1602 (O_1602,N_14792,N_14279);
xor UO_1603 (O_1603,N_14566,N_14989);
and UO_1604 (O_1604,N_14787,N_14047);
or UO_1605 (O_1605,N_14357,N_14889);
and UO_1606 (O_1606,N_14157,N_14701);
nor UO_1607 (O_1607,N_14820,N_14554);
or UO_1608 (O_1608,N_14713,N_14014);
or UO_1609 (O_1609,N_14561,N_14502);
xnor UO_1610 (O_1610,N_14334,N_14621);
nand UO_1611 (O_1611,N_14837,N_14747);
xor UO_1612 (O_1612,N_14142,N_14883);
xnor UO_1613 (O_1613,N_14044,N_14527);
nand UO_1614 (O_1614,N_14485,N_14627);
and UO_1615 (O_1615,N_14527,N_14522);
or UO_1616 (O_1616,N_14446,N_14094);
nand UO_1617 (O_1617,N_14752,N_14506);
and UO_1618 (O_1618,N_14846,N_14192);
nand UO_1619 (O_1619,N_14097,N_14896);
and UO_1620 (O_1620,N_14087,N_14310);
or UO_1621 (O_1621,N_14703,N_14756);
xor UO_1622 (O_1622,N_14516,N_14853);
nor UO_1623 (O_1623,N_14857,N_14140);
and UO_1624 (O_1624,N_14853,N_14157);
or UO_1625 (O_1625,N_14645,N_14784);
or UO_1626 (O_1626,N_14199,N_14346);
or UO_1627 (O_1627,N_14303,N_14091);
or UO_1628 (O_1628,N_14428,N_14524);
xor UO_1629 (O_1629,N_14266,N_14661);
xnor UO_1630 (O_1630,N_14308,N_14491);
and UO_1631 (O_1631,N_14306,N_14439);
and UO_1632 (O_1632,N_14963,N_14490);
and UO_1633 (O_1633,N_14330,N_14959);
nand UO_1634 (O_1634,N_14076,N_14016);
nand UO_1635 (O_1635,N_14854,N_14395);
nor UO_1636 (O_1636,N_14173,N_14223);
nand UO_1637 (O_1637,N_14158,N_14895);
or UO_1638 (O_1638,N_14770,N_14232);
or UO_1639 (O_1639,N_14875,N_14814);
nor UO_1640 (O_1640,N_14490,N_14772);
xor UO_1641 (O_1641,N_14685,N_14377);
nor UO_1642 (O_1642,N_14112,N_14595);
xor UO_1643 (O_1643,N_14567,N_14545);
nor UO_1644 (O_1644,N_14084,N_14061);
and UO_1645 (O_1645,N_14176,N_14626);
nand UO_1646 (O_1646,N_14703,N_14792);
or UO_1647 (O_1647,N_14713,N_14329);
nor UO_1648 (O_1648,N_14226,N_14577);
xnor UO_1649 (O_1649,N_14452,N_14913);
or UO_1650 (O_1650,N_14454,N_14695);
nand UO_1651 (O_1651,N_14457,N_14045);
nor UO_1652 (O_1652,N_14876,N_14632);
nor UO_1653 (O_1653,N_14714,N_14309);
nand UO_1654 (O_1654,N_14800,N_14155);
nor UO_1655 (O_1655,N_14295,N_14273);
or UO_1656 (O_1656,N_14796,N_14823);
xnor UO_1657 (O_1657,N_14074,N_14422);
and UO_1658 (O_1658,N_14169,N_14757);
or UO_1659 (O_1659,N_14665,N_14389);
xor UO_1660 (O_1660,N_14672,N_14324);
or UO_1661 (O_1661,N_14186,N_14915);
or UO_1662 (O_1662,N_14065,N_14722);
or UO_1663 (O_1663,N_14599,N_14136);
or UO_1664 (O_1664,N_14629,N_14449);
xnor UO_1665 (O_1665,N_14906,N_14304);
and UO_1666 (O_1666,N_14791,N_14866);
nand UO_1667 (O_1667,N_14673,N_14061);
nor UO_1668 (O_1668,N_14827,N_14943);
xor UO_1669 (O_1669,N_14959,N_14810);
nor UO_1670 (O_1670,N_14044,N_14464);
nor UO_1671 (O_1671,N_14791,N_14024);
nand UO_1672 (O_1672,N_14020,N_14605);
and UO_1673 (O_1673,N_14086,N_14024);
nand UO_1674 (O_1674,N_14203,N_14467);
or UO_1675 (O_1675,N_14222,N_14710);
xnor UO_1676 (O_1676,N_14994,N_14877);
or UO_1677 (O_1677,N_14224,N_14765);
nor UO_1678 (O_1678,N_14211,N_14591);
nand UO_1679 (O_1679,N_14843,N_14389);
nor UO_1680 (O_1680,N_14091,N_14001);
nor UO_1681 (O_1681,N_14756,N_14753);
and UO_1682 (O_1682,N_14816,N_14397);
nand UO_1683 (O_1683,N_14240,N_14787);
or UO_1684 (O_1684,N_14969,N_14153);
or UO_1685 (O_1685,N_14506,N_14969);
xnor UO_1686 (O_1686,N_14435,N_14668);
and UO_1687 (O_1687,N_14803,N_14457);
or UO_1688 (O_1688,N_14125,N_14383);
or UO_1689 (O_1689,N_14740,N_14246);
or UO_1690 (O_1690,N_14135,N_14551);
nor UO_1691 (O_1691,N_14888,N_14273);
nor UO_1692 (O_1692,N_14545,N_14632);
xnor UO_1693 (O_1693,N_14290,N_14647);
or UO_1694 (O_1694,N_14950,N_14509);
xnor UO_1695 (O_1695,N_14490,N_14979);
or UO_1696 (O_1696,N_14378,N_14471);
or UO_1697 (O_1697,N_14434,N_14953);
xnor UO_1698 (O_1698,N_14711,N_14299);
nor UO_1699 (O_1699,N_14150,N_14701);
xnor UO_1700 (O_1700,N_14357,N_14920);
or UO_1701 (O_1701,N_14322,N_14528);
nand UO_1702 (O_1702,N_14065,N_14417);
or UO_1703 (O_1703,N_14297,N_14716);
or UO_1704 (O_1704,N_14452,N_14031);
xor UO_1705 (O_1705,N_14093,N_14750);
or UO_1706 (O_1706,N_14977,N_14741);
and UO_1707 (O_1707,N_14643,N_14416);
nor UO_1708 (O_1708,N_14023,N_14216);
nand UO_1709 (O_1709,N_14206,N_14106);
nor UO_1710 (O_1710,N_14772,N_14860);
nor UO_1711 (O_1711,N_14966,N_14257);
nand UO_1712 (O_1712,N_14340,N_14411);
and UO_1713 (O_1713,N_14259,N_14690);
or UO_1714 (O_1714,N_14342,N_14566);
xnor UO_1715 (O_1715,N_14997,N_14383);
and UO_1716 (O_1716,N_14910,N_14293);
and UO_1717 (O_1717,N_14167,N_14127);
nand UO_1718 (O_1718,N_14920,N_14669);
and UO_1719 (O_1719,N_14500,N_14227);
nor UO_1720 (O_1720,N_14184,N_14429);
and UO_1721 (O_1721,N_14506,N_14154);
xor UO_1722 (O_1722,N_14623,N_14081);
or UO_1723 (O_1723,N_14156,N_14128);
and UO_1724 (O_1724,N_14774,N_14299);
or UO_1725 (O_1725,N_14481,N_14476);
or UO_1726 (O_1726,N_14662,N_14073);
and UO_1727 (O_1727,N_14577,N_14904);
nand UO_1728 (O_1728,N_14852,N_14114);
nor UO_1729 (O_1729,N_14864,N_14279);
xnor UO_1730 (O_1730,N_14798,N_14857);
nor UO_1731 (O_1731,N_14948,N_14891);
nor UO_1732 (O_1732,N_14246,N_14647);
or UO_1733 (O_1733,N_14078,N_14728);
xor UO_1734 (O_1734,N_14667,N_14373);
and UO_1735 (O_1735,N_14183,N_14921);
xor UO_1736 (O_1736,N_14834,N_14792);
or UO_1737 (O_1737,N_14504,N_14161);
and UO_1738 (O_1738,N_14398,N_14587);
and UO_1739 (O_1739,N_14709,N_14610);
and UO_1740 (O_1740,N_14723,N_14132);
nand UO_1741 (O_1741,N_14590,N_14058);
nor UO_1742 (O_1742,N_14438,N_14761);
or UO_1743 (O_1743,N_14526,N_14927);
nand UO_1744 (O_1744,N_14646,N_14336);
nand UO_1745 (O_1745,N_14562,N_14118);
xnor UO_1746 (O_1746,N_14363,N_14563);
or UO_1747 (O_1747,N_14774,N_14267);
xnor UO_1748 (O_1748,N_14431,N_14124);
or UO_1749 (O_1749,N_14301,N_14182);
nand UO_1750 (O_1750,N_14536,N_14884);
or UO_1751 (O_1751,N_14550,N_14879);
nand UO_1752 (O_1752,N_14874,N_14472);
nor UO_1753 (O_1753,N_14872,N_14656);
and UO_1754 (O_1754,N_14037,N_14055);
nand UO_1755 (O_1755,N_14659,N_14052);
and UO_1756 (O_1756,N_14640,N_14090);
nand UO_1757 (O_1757,N_14248,N_14694);
nand UO_1758 (O_1758,N_14728,N_14746);
and UO_1759 (O_1759,N_14568,N_14061);
or UO_1760 (O_1760,N_14812,N_14534);
and UO_1761 (O_1761,N_14527,N_14907);
xor UO_1762 (O_1762,N_14397,N_14954);
nor UO_1763 (O_1763,N_14932,N_14886);
or UO_1764 (O_1764,N_14287,N_14854);
nor UO_1765 (O_1765,N_14107,N_14106);
or UO_1766 (O_1766,N_14143,N_14851);
or UO_1767 (O_1767,N_14867,N_14189);
xnor UO_1768 (O_1768,N_14620,N_14851);
or UO_1769 (O_1769,N_14647,N_14254);
nand UO_1770 (O_1770,N_14857,N_14205);
and UO_1771 (O_1771,N_14754,N_14192);
nand UO_1772 (O_1772,N_14217,N_14799);
nor UO_1773 (O_1773,N_14923,N_14982);
nor UO_1774 (O_1774,N_14870,N_14481);
or UO_1775 (O_1775,N_14188,N_14683);
nor UO_1776 (O_1776,N_14198,N_14689);
xor UO_1777 (O_1777,N_14662,N_14226);
or UO_1778 (O_1778,N_14603,N_14510);
and UO_1779 (O_1779,N_14856,N_14102);
nor UO_1780 (O_1780,N_14971,N_14820);
xnor UO_1781 (O_1781,N_14310,N_14565);
and UO_1782 (O_1782,N_14184,N_14620);
nand UO_1783 (O_1783,N_14650,N_14074);
and UO_1784 (O_1784,N_14081,N_14502);
nand UO_1785 (O_1785,N_14067,N_14937);
nand UO_1786 (O_1786,N_14681,N_14423);
or UO_1787 (O_1787,N_14418,N_14958);
or UO_1788 (O_1788,N_14599,N_14130);
or UO_1789 (O_1789,N_14890,N_14099);
and UO_1790 (O_1790,N_14058,N_14628);
nor UO_1791 (O_1791,N_14741,N_14659);
and UO_1792 (O_1792,N_14800,N_14187);
and UO_1793 (O_1793,N_14128,N_14761);
xnor UO_1794 (O_1794,N_14225,N_14345);
and UO_1795 (O_1795,N_14512,N_14859);
nor UO_1796 (O_1796,N_14113,N_14171);
and UO_1797 (O_1797,N_14049,N_14796);
xor UO_1798 (O_1798,N_14380,N_14101);
nor UO_1799 (O_1799,N_14992,N_14200);
and UO_1800 (O_1800,N_14897,N_14606);
or UO_1801 (O_1801,N_14338,N_14079);
nand UO_1802 (O_1802,N_14125,N_14346);
and UO_1803 (O_1803,N_14515,N_14238);
or UO_1804 (O_1804,N_14652,N_14013);
nor UO_1805 (O_1805,N_14791,N_14603);
and UO_1806 (O_1806,N_14677,N_14921);
nor UO_1807 (O_1807,N_14624,N_14404);
xnor UO_1808 (O_1808,N_14560,N_14334);
and UO_1809 (O_1809,N_14701,N_14614);
nand UO_1810 (O_1810,N_14930,N_14850);
or UO_1811 (O_1811,N_14085,N_14124);
and UO_1812 (O_1812,N_14515,N_14601);
or UO_1813 (O_1813,N_14114,N_14445);
nor UO_1814 (O_1814,N_14909,N_14548);
nand UO_1815 (O_1815,N_14305,N_14208);
and UO_1816 (O_1816,N_14833,N_14101);
and UO_1817 (O_1817,N_14641,N_14181);
xor UO_1818 (O_1818,N_14307,N_14548);
nand UO_1819 (O_1819,N_14573,N_14043);
or UO_1820 (O_1820,N_14502,N_14067);
and UO_1821 (O_1821,N_14675,N_14775);
nor UO_1822 (O_1822,N_14563,N_14642);
nand UO_1823 (O_1823,N_14701,N_14589);
xor UO_1824 (O_1824,N_14468,N_14217);
and UO_1825 (O_1825,N_14616,N_14677);
or UO_1826 (O_1826,N_14850,N_14098);
and UO_1827 (O_1827,N_14816,N_14551);
or UO_1828 (O_1828,N_14057,N_14770);
nand UO_1829 (O_1829,N_14421,N_14511);
nor UO_1830 (O_1830,N_14256,N_14100);
or UO_1831 (O_1831,N_14519,N_14041);
nor UO_1832 (O_1832,N_14853,N_14694);
and UO_1833 (O_1833,N_14923,N_14909);
or UO_1834 (O_1834,N_14794,N_14320);
nand UO_1835 (O_1835,N_14696,N_14881);
or UO_1836 (O_1836,N_14745,N_14917);
nor UO_1837 (O_1837,N_14073,N_14603);
or UO_1838 (O_1838,N_14300,N_14005);
and UO_1839 (O_1839,N_14534,N_14150);
nor UO_1840 (O_1840,N_14032,N_14554);
nor UO_1841 (O_1841,N_14961,N_14911);
xnor UO_1842 (O_1842,N_14102,N_14605);
nor UO_1843 (O_1843,N_14690,N_14310);
or UO_1844 (O_1844,N_14063,N_14028);
and UO_1845 (O_1845,N_14905,N_14846);
or UO_1846 (O_1846,N_14911,N_14008);
nand UO_1847 (O_1847,N_14608,N_14560);
nand UO_1848 (O_1848,N_14567,N_14857);
or UO_1849 (O_1849,N_14746,N_14143);
or UO_1850 (O_1850,N_14515,N_14799);
nand UO_1851 (O_1851,N_14815,N_14458);
nand UO_1852 (O_1852,N_14917,N_14813);
nand UO_1853 (O_1853,N_14919,N_14686);
nand UO_1854 (O_1854,N_14734,N_14666);
xnor UO_1855 (O_1855,N_14732,N_14231);
nand UO_1856 (O_1856,N_14260,N_14405);
and UO_1857 (O_1857,N_14723,N_14180);
nor UO_1858 (O_1858,N_14987,N_14495);
nor UO_1859 (O_1859,N_14284,N_14245);
xor UO_1860 (O_1860,N_14914,N_14294);
or UO_1861 (O_1861,N_14346,N_14229);
nor UO_1862 (O_1862,N_14603,N_14511);
nor UO_1863 (O_1863,N_14503,N_14939);
and UO_1864 (O_1864,N_14525,N_14702);
or UO_1865 (O_1865,N_14646,N_14313);
or UO_1866 (O_1866,N_14464,N_14399);
or UO_1867 (O_1867,N_14080,N_14231);
xor UO_1868 (O_1868,N_14307,N_14251);
nand UO_1869 (O_1869,N_14290,N_14359);
nor UO_1870 (O_1870,N_14526,N_14795);
and UO_1871 (O_1871,N_14498,N_14263);
and UO_1872 (O_1872,N_14319,N_14632);
and UO_1873 (O_1873,N_14858,N_14302);
or UO_1874 (O_1874,N_14977,N_14589);
nand UO_1875 (O_1875,N_14288,N_14502);
nand UO_1876 (O_1876,N_14712,N_14872);
or UO_1877 (O_1877,N_14880,N_14882);
and UO_1878 (O_1878,N_14784,N_14773);
xor UO_1879 (O_1879,N_14926,N_14673);
nor UO_1880 (O_1880,N_14072,N_14907);
nor UO_1881 (O_1881,N_14790,N_14070);
nor UO_1882 (O_1882,N_14520,N_14904);
and UO_1883 (O_1883,N_14996,N_14908);
nor UO_1884 (O_1884,N_14763,N_14609);
or UO_1885 (O_1885,N_14353,N_14185);
and UO_1886 (O_1886,N_14592,N_14187);
nor UO_1887 (O_1887,N_14018,N_14575);
or UO_1888 (O_1888,N_14272,N_14157);
nor UO_1889 (O_1889,N_14163,N_14138);
nand UO_1890 (O_1890,N_14146,N_14191);
and UO_1891 (O_1891,N_14880,N_14612);
and UO_1892 (O_1892,N_14362,N_14929);
xor UO_1893 (O_1893,N_14395,N_14108);
and UO_1894 (O_1894,N_14231,N_14516);
xor UO_1895 (O_1895,N_14922,N_14630);
xnor UO_1896 (O_1896,N_14139,N_14316);
and UO_1897 (O_1897,N_14776,N_14152);
or UO_1898 (O_1898,N_14641,N_14576);
nor UO_1899 (O_1899,N_14846,N_14924);
nor UO_1900 (O_1900,N_14392,N_14141);
nor UO_1901 (O_1901,N_14142,N_14134);
nand UO_1902 (O_1902,N_14450,N_14033);
nand UO_1903 (O_1903,N_14689,N_14997);
or UO_1904 (O_1904,N_14000,N_14091);
and UO_1905 (O_1905,N_14466,N_14302);
nand UO_1906 (O_1906,N_14177,N_14881);
nor UO_1907 (O_1907,N_14893,N_14202);
nand UO_1908 (O_1908,N_14546,N_14483);
xor UO_1909 (O_1909,N_14809,N_14323);
xor UO_1910 (O_1910,N_14563,N_14683);
or UO_1911 (O_1911,N_14676,N_14303);
xor UO_1912 (O_1912,N_14003,N_14011);
nand UO_1913 (O_1913,N_14121,N_14260);
or UO_1914 (O_1914,N_14245,N_14084);
nand UO_1915 (O_1915,N_14183,N_14174);
and UO_1916 (O_1916,N_14256,N_14635);
or UO_1917 (O_1917,N_14773,N_14186);
xor UO_1918 (O_1918,N_14331,N_14121);
xnor UO_1919 (O_1919,N_14369,N_14055);
and UO_1920 (O_1920,N_14982,N_14688);
nand UO_1921 (O_1921,N_14787,N_14092);
nor UO_1922 (O_1922,N_14066,N_14932);
nor UO_1923 (O_1923,N_14314,N_14024);
or UO_1924 (O_1924,N_14516,N_14446);
and UO_1925 (O_1925,N_14446,N_14974);
nand UO_1926 (O_1926,N_14211,N_14661);
and UO_1927 (O_1927,N_14319,N_14927);
nand UO_1928 (O_1928,N_14338,N_14086);
xor UO_1929 (O_1929,N_14621,N_14684);
and UO_1930 (O_1930,N_14920,N_14495);
nand UO_1931 (O_1931,N_14128,N_14217);
nor UO_1932 (O_1932,N_14792,N_14149);
nor UO_1933 (O_1933,N_14471,N_14995);
xnor UO_1934 (O_1934,N_14282,N_14417);
xor UO_1935 (O_1935,N_14211,N_14711);
and UO_1936 (O_1936,N_14136,N_14818);
xnor UO_1937 (O_1937,N_14023,N_14326);
xnor UO_1938 (O_1938,N_14091,N_14368);
nor UO_1939 (O_1939,N_14936,N_14840);
xnor UO_1940 (O_1940,N_14770,N_14211);
and UO_1941 (O_1941,N_14690,N_14555);
nor UO_1942 (O_1942,N_14199,N_14825);
and UO_1943 (O_1943,N_14139,N_14518);
nand UO_1944 (O_1944,N_14373,N_14981);
and UO_1945 (O_1945,N_14610,N_14805);
xor UO_1946 (O_1946,N_14066,N_14175);
or UO_1947 (O_1947,N_14385,N_14443);
or UO_1948 (O_1948,N_14647,N_14432);
nor UO_1949 (O_1949,N_14531,N_14049);
or UO_1950 (O_1950,N_14815,N_14209);
or UO_1951 (O_1951,N_14252,N_14835);
nand UO_1952 (O_1952,N_14477,N_14734);
nor UO_1953 (O_1953,N_14480,N_14388);
xnor UO_1954 (O_1954,N_14548,N_14808);
xnor UO_1955 (O_1955,N_14215,N_14670);
nand UO_1956 (O_1956,N_14256,N_14533);
xor UO_1957 (O_1957,N_14718,N_14092);
nor UO_1958 (O_1958,N_14173,N_14514);
or UO_1959 (O_1959,N_14298,N_14887);
xnor UO_1960 (O_1960,N_14999,N_14904);
and UO_1961 (O_1961,N_14252,N_14381);
or UO_1962 (O_1962,N_14080,N_14075);
and UO_1963 (O_1963,N_14163,N_14029);
xor UO_1964 (O_1964,N_14247,N_14438);
and UO_1965 (O_1965,N_14646,N_14583);
nor UO_1966 (O_1966,N_14924,N_14391);
nand UO_1967 (O_1967,N_14511,N_14058);
or UO_1968 (O_1968,N_14418,N_14473);
nand UO_1969 (O_1969,N_14047,N_14399);
xnor UO_1970 (O_1970,N_14052,N_14869);
or UO_1971 (O_1971,N_14375,N_14003);
or UO_1972 (O_1972,N_14111,N_14299);
nor UO_1973 (O_1973,N_14232,N_14190);
or UO_1974 (O_1974,N_14569,N_14888);
or UO_1975 (O_1975,N_14593,N_14788);
or UO_1976 (O_1976,N_14555,N_14586);
nor UO_1977 (O_1977,N_14051,N_14992);
or UO_1978 (O_1978,N_14783,N_14439);
nand UO_1979 (O_1979,N_14172,N_14776);
and UO_1980 (O_1980,N_14450,N_14911);
xnor UO_1981 (O_1981,N_14328,N_14582);
xor UO_1982 (O_1982,N_14519,N_14679);
xor UO_1983 (O_1983,N_14706,N_14785);
nor UO_1984 (O_1984,N_14776,N_14604);
nor UO_1985 (O_1985,N_14432,N_14801);
and UO_1986 (O_1986,N_14607,N_14005);
or UO_1987 (O_1987,N_14673,N_14642);
xor UO_1988 (O_1988,N_14024,N_14725);
xor UO_1989 (O_1989,N_14830,N_14077);
or UO_1990 (O_1990,N_14802,N_14619);
and UO_1991 (O_1991,N_14227,N_14094);
nand UO_1992 (O_1992,N_14494,N_14987);
xnor UO_1993 (O_1993,N_14057,N_14553);
xor UO_1994 (O_1994,N_14214,N_14384);
nand UO_1995 (O_1995,N_14537,N_14769);
xnor UO_1996 (O_1996,N_14137,N_14684);
or UO_1997 (O_1997,N_14894,N_14010);
nor UO_1998 (O_1998,N_14996,N_14625);
nor UO_1999 (O_1999,N_14165,N_14593);
endmodule