module basic_1000_10000_1500_10_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_294,In_358);
nand U1 (N_1,In_759,In_981);
or U2 (N_2,In_910,In_502);
and U3 (N_3,In_987,In_181);
nor U4 (N_4,In_685,In_8);
or U5 (N_5,In_606,In_832);
nor U6 (N_6,In_947,In_104);
or U7 (N_7,In_737,In_422);
nand U8 (N_8,In_211,In_419);
nor U9 (N_9,In_913,In_403);
nor U10 (N_10,In_518,In_545);
nand U11 (N_11,In_595,In_377);
nor U12 (N_12,In_508,In_875);
or U13 (N_13,In_806,In_564);
nor U14 (N_14,In_282,In_465);
or U15 (N_15,In_519,In_989);
nand U16 (N_16,In_958,In_82);
nor U17 (N_17,In_186,In_299);
nand U18 (N_18,In_676,In_451);
nor U19 (N_19,In_479,In_201);
or U20 (N_20,In_919,In_674);
and U21 (N_21,In_311,In_399);
nand U22 (N_22,In_648,In_322);
nor U23 (N_23,In_598,In_743);
nand U24 (N_24,In_251,In_51);
nand U25 (N_25,In_705,In_29);
nor U26 (N_26,In_90,In_318);
nand U27 (N_27,In_15,In_787);
nand U28 (N_28,In_939,In_242);
nand U29 (N_29,In_94,In_857);
nand U30 (N_30,In_547,In_383);
and U31 (N_31,In_49,In_456);
and U32 (N_32,In_470,In_380);
nor U33 (N_33,In_930,In_960);
or U34 (N_34,In_991,In_656);
nand U35 (N_35,In_878,In_900);
or U36 (N_36,In_530,In_315);
and U37 (N_37,In_385,In_701);
nor U38 (N_38,In_852,In_611);
or U39 (N_39,In_692,In_753);
nand U40 (N_40,In_397,In_973);
or U41 (N_41,In_307,In_480);
nand U42 (N_42,In_733,In_744);
and U43 (N_43,In_174,In_16);
nand U44 (N_44,In_749,In_509);
nor U45 (N_45,In_190,In_241);
nand U46 (N_46,In_56,In_75);
and U47 (N_47,In_940,In_199);
or U48 (N_48,In_526,In_452);
or U49 (N_49,In_630,In_130);
nand U50 (N_50,In_466,In_129);
nand U51 (N_51,In_459,In_253);
nor U52 (N_52,In_928,In_936);
nand U53 (N_53,In_952,In_226);
or U54 (N_54,In_810,In_881);
nand U55 (N_55,In_325,In_690);
or U56 (N_56,In_162,In_2);
and U57 (N_57,In_487,In_212);
nand U58 (N_58,In_37,In_788);
and U59 (N_59,In_99,In_70);
nand U60 (N_60,In_636,In_43);
xor U61 (N_61,In_142,In_567);
and U62 (N_62,In_227,In_781);
and U63 (N_63,In_147,In_388);
nand U64 (N_64,In_483,In_861);
nand U65 (N_65,In_120,In_264);
nor U66 (N_66,In_645,In_571);
nand U67 (N_67,In_516,In_12);
nor U68 (N_68,In_402,In_409);
nand U69 (N_69,In_180,In_341);
nor U70 (N_70,In_557,In_491);
or U71 (N_71,In_204,In_895);
and U72 (N_72,In_735,In_851);
and U73 (N_73,In_945,In_712);
nor U74 (N_74,In_905,In_833);
nand U75 (N_75,In_664,In_379);
or U76 (N_76,In_644,In_245);
or U77 (N_77,In_198,In_720);
nor U78 (N_78,In_624,In_304);
and U79 (N_79,In_501,In_706);
nand U80 (N_80,In_969,In_757);
nor U81 (N_81,In_755,In_448);
nor U82 (N_82,In_924,In_638);
and U83 (N_83,In_356,In_351);
nor U84 (N_84,In_196,In_133);
and U85 (N_85,In_923,In_751);
nor U86 (N_86,In_903,In_175);
and U87 (N_87,In_782,In_734);
xnor U88 (N_88,In_95,In_141);
or U89 (N_89,In_192,In_262);
or U90 (N_90,In_992,In_440);
or U91 (N_91,In_343,In_985);
or U92 (N_92,In_561,In_689);
nand U93 (N_93,In_821,In_955);
or U94 (N_94,In_223,In_899);
or U95 (N_95,In_844,In_31);
nor U96 (N_96,In_885,In_641);
nor U97 (N_97,In_71,In_261);
or U98 (N_98,In_728,In_69);
nand U99 (N_99,In_36,In_877);
xor U100 (N_100,In_461,In_627);
or U101 (N_101,In_436,In_804);
nand U102 (N_102,In_775,In_584);
nor U103 (N_103,In_121,In_702);
and U104 (N_104,In_184,In_21);
and U105 (N_105,In_244,In_313);
and U106 (N_106,In_283,In_27);
nor U107 (N_107,In_658,In_125);
and U108 (N_108,In_297,In_615);
or U109 (N_109,In_32,In_964);
nand U110 (N_110,In_937,In_58);
nand U111 (N_111,In_462,In_953);
nand U112 (N_112,In_965,In_391);
nand U113 (N_113,In_783,In_314);
nor U114 (N_114,In_990,In_866);
or U115 (N_115,In_63,In_770);
and U116 (N_116,In_13,In_4);
nor U117 (N_117,In_879,In_655);
and U118 (N_118,In_273,In_962);
or U119 (N_119,In_441,In_902);
or U120 (N_120,In_772,In_836);
nor U121 (N_121,In_335,In_96);
or U122 (N_122,In_842,In_333);
nand U123 (N_123,In_476,In_277);
and U124 (N_124,In_276,In_219);
nand U125 (N_125,In_73,In_118);
and U126 (N_126,In_258,In_997);
and U127 (N_127,In_976,In_552);
nand U128 (N_128,In_709,In_270);
nand U129 (N_129,In_376,In_26);
and U130 (N_130,In_532,In_579);
and U131 (N_131,In_725,In_815);
or U132 (N_132,In_24,In_616);
nand U133 (N_133,In_748,In_809);
or U134 (N_134,In_959,In_123);
nand U135 (N_135,In_726,In_346);
nand U136 (N_136,In_865,In_368);
nand U137 (N_137,In_353,In_256);
nor U138 (N_138,In_767,In_247);
and U139 (N_139,In_637,In_617);
xor U140 (N_140,In_386,In_670);
nor U141 (N_141,In_537,In_574);
and U142 (N_142,In_298,In_352);
nor U143 (N_143,In_891,In_978);
nand U144 (N_144,In_289,In_536);
nand U145 (N_145,In_850,In_10);
or U146 (N_146,In_257,In_633);
or U147 (N_147,In_541,In_477);
nor U148 (N_148,In_546,In_185);
or U149 (N_149,In_429,In_215);
nor U150 (N_150,In_485,In_275);
and U151 (N_151,In_66,In_796);
and U152 (N_152,In_236,In_824);
nor U153 (N_153,In_115,In_102);
nor U154 (N_154,In_326,In_986);
and U155 (N_155,In_158,In_825);
nor U156 (N_156,In_568,In_999);
nand U157 (N_157,In_507,In_797);
xor U158 (N_158,In_588,In_620);
and U159 (N_159,In_166,In_840);
and U160 (N_160,In_621,In_442);
and U161 (N_161,In_418,In_450);
or U162 (N_162,In_40,In_375);
nand U163 (N_163,In_387,In_478);
nand U164 (N_164,In_623,In_635);
nor U165 (N_165,In_979,In_332);
and U166 (N_166,In_540,In_424);
nand U167 (N_167,In_908,In_854);
nand U168 (N_168,In_453,In_416);
nand U169 (N_169,In_18,In_570);
nand U170 (N_170,In_41,In_179);
nand U171 (N_171,In_372,In_826);
nand U172 (N_172,In_800,In_604);
and U173 (N_173,In_355,In_946);
nand U174 (N_174,In_330,In_417);
and U175 (N_175,In_931,In_699);
or U176 (N_176,In_197,In_493);
nand U177 (N_177,In_243,In_874);
nor U178 (N_178,In_533,In_163);
and U179 (N_179,In_608,In_592);
and U180 (N_180,In_160,In_415);
nand U181 (N_181,In_367,In_126);
and U182 (N_182,In_287,In_880);
nand U183 (N_183,In_148,In_867);
and U184 (N_184,In_57,In_35);
nand U185 (N_185,In_444,In_228);
nor U186 (N_186,In_848,In_543);
nor U187 (N_187,In_182,In_950);
nor U188 (N_188,In_700,In_378);
nor U189 (N_189,In_432,In_187);
nor U190 (N_190,In_619,In_773);
nor U191 (N_191,In_205,In_194);
nor U192 (N_192,In_935,In_534);
and U193 (N_193,In_156,In_200);
and U194 (N_194,In_968,In_14);
xor U195 (N_195,In_739,In_252);
or U196 (N_196,In_464,In_413);
or U197 (N_197,In_414,In_293);
nor U198 (N_198,In_914,In_774);
nand U199 (N_199,In_88,In_538);
nand U200 (N_200,In_183,In_89);
nor U201 (N_201,In_319,In_25);
nand U202 (N_202,In_601,In_662);
or U203 (N_203,In_607,In_993);
nand U204 (N_204,In_439,In_827);
nand U205 (N_205,In_746,In_549);
nor U206 (N_206,In_423,In_151);
nor U207 (N_207,In_625,In_67);
and U208 (N_208,In_678,In_437);
nor U209 (N_209,In_631,In_60);
nand U210 (N_210,In_281,In_535);
nand U211 (N_211,In_85,In_272);
nor U212 (N_212,In_994,In_814);
nor U213 (N_213,In_578,In_680);
nor U214 (N_214,In_525,In_512);
and U215 (N_215,In_941,In_687);
nand U216 (N_216,In_593,In_114);
or U217 (N_217,In_134,In_505);
xor U218 (N_218,In_371,In_855);
or U219 (N_219,In_722,In_742);
nand U220 (N_220,In_932,In_240);
nor U221 (N_221,In_468,In_915);
and U222 (N_222,In_168,In_718);
xnor U223 (N_223,In_539,In_511);
or U224 (N_224,In_711,In_818);
nand U225 (N_225,In_847,In_78);
nand U226 (N_226,In_929,In_345);
nand U227 (N_227,In_404,In_154);
nor U228 (N_228,In_5,In_410);
or U229 (N_229,In_87,In_308);
and U230 (N_230,In_805,In_317);
nand U231 (N_231,In_92,In_406);
nor U232 (N_232,In_754,In_150);
nand U233 (N_233,In_271,In_207);
nand U234 (N_234,In_135,In_472);
nor U235 (N_235,In_425,In_292);
nand U236 (N_236,In_612,In_50);
or U237 (N_237,In_823,In_471);
and U238 (N_238,In_221,In_911);
nor U239 (N_239,In_618,In_366);
and U240 (N_240,In_431,In_360);
nand U241 (N_241,In_747,In_122);
nor U242 (N_242,In_305,In_514);
or U243 (N_243,In_917,In_176);
and U244 (N_244,In_9,In_693);
and U245 (N_245,In_892,In_822);
or U246 (N_246,In_614,In_336);
or U247 (N_247,In_338,In_652);
or U248 (N_248,In_408,In_752);
and U249 (N_249,In_750,In_907);
or U250 (N_250,In_136,In_972);
nand U251 (N_251,In_11,In_523);
nand U252 (N_252,In_124,In_771);
nor U253 (N_253,In_398,In_698);
and U254 (N_254,In_691,In_428);
and U255 (N_255,In_789,In_819);
or U256 (N_256,In_177,In_369);
nand U257 (N_257,In_337,In_597);
nand U258 (N_258,In_284,In_629);
and U259 (N_259,In_155,In_862);
nor U260 (N_260,In_927,In_603);
or U261 (N_261,In_52,In_808);
nand U262 (N_262,In_544,In_449);
or U263 (N_263,In_237,In_684);
or U264 (N_264,In_33,In_503);
nor U265 (N_265,In_551,In_229);
nor U266 (N_266,In_859,In_626);
nand U267 (N_267,In_721,In_686);
and U268 (N_268,In_663,In_967);
nand U269 (N_269,In_602,In_48);
or U270 (N_270,In_671,In_364);
nor U271 (N_271,In_517,In_107);
and U272 (N_272,In_764,In_839);
nand U273 (N_273,In_171,In_249);
nand U274 (N_274,In_756,In_646);
or U275 (N_275,In_768,In_421);
nand U276 (N_276,In_695,In_886);
and U277 (N_277,In_843,In_816);
or U278 (N_278,In_576,In_113);
or U279 (N_279,In_494,In_586);
or U280 (N_280,In_72,In_301);
nor U281 (N_281,In_195,In_666);
and U282 (N_282,In_217,In_394);
nor U283 (N_283,In_795,In_361);
or U284 (N_284,In_741,In_661);
nand U285 (N_285,In_675,In_765);
nor U286 (N_286,In_393,In_220);
nor U287 (N_287,In_17,In_39);
or U288 (N_288,In_395,In_389);
or U289 (N_289,In_558,In_382);
nand U290 (N_290,In_527,In_834);
or U291 (N_291,In_285,In_715);
nor U292 (N_292,In_396,In_786);
or U293 (N_293,In_613,In_893);
and U294 (N_294,In_901,In_871);
and U295 (N_295,In_454,In_224);
nor U296 (N_296,In_486,In_44);
nand U297 (N_297,In_573,In_563);
nor U298 (N_298,In_169,In_776);
nor U299 (N_299,In_250,In_1);
xor U300 (N_300,In_951,In_498);
nand U301 (N_301,In_23,In_344);
and U302 (N_302,In_912,In_373);
or U303 (N_303,In_149,In_707);
nand U304 (N_304,In_599,In_777);
nand U305 (N_305,In_600,In_898);
and U306 (N_306,In_622,In_554);
nor U307 (N_307,In_873,In_112);
or U308 (N_308,In_132,In_34);
and U309 (N_309,In_77,In_736);
nand U310 (N_310,In_350,In_970);
nor U311 (N_311,In_357,In_696);
and U312 (N_312,In_339,In_374);
and U313 (N_313,In_323,In_996);
and U314 (N_314,In_269,In_469);
or U315 (N_315,In_84,In_384);
or U316 (N_316,In_665,In_434);
and U317 (N_317,In_327,In_80);
or U318 (N_318,In_673,In_938);
nor U319 (N_319,In_222,In_164);
nand U320 (N_320,In_111,In_274);
nand U321 (N_321,In_841,In_575);
nand U322 (N_322,In_798,In_802);
nor U323 (N_323,In_697,In_758);
nand U324 (N_324,In_870,In_933);
and U325 (N_325,In_916,In_831);
nand U326 (N_326,In_86,In_650);
nand U327 (N_327,In_320,In_731);
or U328 (N_328,In_191,In_81);
and U329 (N_329,In_101,In_206);
nor U330 (N_330,In_324,In_580);
nand U331 (N_331,In_888,In_583);
nand U332 (N_332,In_813,In_137);
xnor U333 (N_333,In_254,In_458);
nor U334 (N_334,In_628,In_553);
or U335 (N_335,In_980,In_55);
and U336 (N_336,In_433,In_145);
and U337 (N_337,In_766,In_172);
and U338 (N_338,In_455,In_110);
nor U339 (N_339,In_500,In_589);
or U340 (N_340,In_203,In_988);
nor U341 (N_341,In_312,In_956);
nor U342 (N_342,In_286,In_811);
nand U343 (N_343,In_407,In_869);
nand U344 (N_344,In_660,In_559);
and U345 (N_345,In_504,In_828);
and U346 (N_346,In_42,In_232);
or U347 (N_347,In_348,In_897);
nor U348 (N_348,In_143,In_643);
nor U349 (N_349,In_146,In_548);
and U350 (N_350,In_189,In_647);
nand U351 (N_351,In_529,In_128);
or U352 (N_352,In_587,In_7);
nand U353 (N_353,In_265,In_19);
and U354 (N_354,In_291,In_381);
and U355 (N_355,In_830,In_708);
nand U356 (N_356,In_642,In_460);
or U357 (N_357,In_426,In_723);
nand U358 (N_358,In_926,In_596);
and U359 (N_359,In_846,In_316);
and U360 (N_360,In_727,In_430);
nand U361 (N_361,In_288,In_259);
or U362 (N_362,In_780,In_340);
nor U363 (N_363,In_679,In_463);
and U364 (N_364,In_79,In_651);
or U365 (N_365,In_496,In_310);
or U366 (N_366,In_520,In_853);
nor U367 (N_367,In_858,In_173);
nand U368 (N_368,In_820,In_225);
nor U369 (N_369,In_904,In_882);
or U370 (N_370,In_446,In_303);
or U371 (N_371,In_942,In_681);
and U372 (N_372,In_710,In_729);
nand U373 (N_373,In_524,In_672);
nand U374 (N_374,In_740,In_778);
nor U375 (N_375,In_975,In_263);
nor U376 (N_376,In_457,In_762);
nand U377 (N_377,In_522,In_210);
or U378 (N_378,In_260,In_248);
nand U379 (N_379,In_634,In_334);
nor U380 (N_380,In_694,In_105);
or U381 (N_381,In_246,In_390);
nor U382 (N_382,In_983,In_639);
nand U383 (N_383,In_515,In_209);
or U384 (N_384,In_216,In_640);
nand U385 (N_385,In_47,In_682);
nand U386 (N_386,In_920,In_817);
nor U387 (N_387,In_349,In_610);
nor U388 (N_388,In_295,In_239);
or U389 (N_389,In_108,In_876);
or U390 (N_390,In_714,In_560);
or U391 (N_391,In_447,In_302);
nand U392 (N_392,In_278,In_61);
or U393 (N_393,In_6,In_632);
nand U394 (N_394,In_745,In_268);
nor U395 (N_395,In_963,In_144);
nand U396 (N_396,In_957,In_769);
nand U397 (N_397,In_889,In_91);
xnor U398 (N_398,In_473,In_412);
nor U399 (N_399,In_45,In_83);
nor U400 (N_400,In_863,In_482);
and U401 (N_401,In_513,In_909);
nand U402 (N_402,In_562,In_234);
nor U403 (N_403,In_296,In_760);
and U404 (N_404,In_669,In_542);
nand U405 (N_405,In_812,In_329);
or U406 (N_406,In_838,In_793);
nand U407 (N_407,In_677,In_331);
and U408 (N_408,In_214,In_427);
nand U409 (N_409,In_309,In_279);
or U410 (N_410,In_170,In_556);
and U411 (N_411,In_127,In_400);
nor U412 (N_412,In_683,In_974);
or U413 (N_413,In_884,In_738);
nand U414 (N_414,In_943,In_188);
or U415 (N_415,In_954,In_392);
xnor U416 (N_416,In_474,In_138);
nand U417 (N_417,In_719,In_300);
nand U418 (N_418,In_792,In_845);
and U419 (N_419,In_347,In_467);
and U420 (N_420,In_202,In_497);
nand U421 (N_421,In_521,In_761);
xor U422 (N_422,In_116,In_688);
nand U423 (N_423,In_157,In_490);
nor U424 (N_424,In_492,In_717);
xnor U425 (N_425,In_76,In_54);
nand U426 (N_426,In_306,In_555);
nor U427 (N_427,In_435,In_948);
nor U428 (N_428,In_38,In_481);
and U429 (N_429,In_65,In_582);
and U430 (N_430,In_609,In_837);
nor U431 (N_431,In_791,In_165);
nor U432 (N_432,In_966,In_894);
and U433 (N_433,In_605,In_208);
nor U434 (N_434,In_117,In_103);
nor U435 (N_435,In_732,In_657);
nor U436 (N_436,In_531,In_100);
nand U437 (N_437,In_238,In_131);
nand U438 (N_438,In_654,In_420);
nor U439 (N_439,In_506,In_475);
nor U440 (N_440,In_109,In_401);
nand U441 (N_441,In_230,In_3);
or U442 (N_442,In_550,In_161);
nand U443 (N_443,In_585,In_918);
nand U444 (N_444,In_984,In_140);
or U445 (N_445,In_30,In_566);
and U446 (N_446,In_98,In_233);
nor U447 (N_447,In_74,In_971);
nand U448 (N_448,In_577,In_794);
nor U449 (N_449,In_887,In_569);
and U450 (N_450,In_20,In_290);
nor U451 (N_451,In_46,In_28);
or U452 (N_452,In_835,In_411);
nor U453 (N_453,In_925,In_235);
or U454 (N_454,In_59,In_724);
nand U455 (N_455,In_213,In_849);
nor U456 (N_456,In_438,In_572);
nand U457 (N_457,In_949,In_119);
nand U458 (N_458,In_445,In_668);
nor U459 (N_459,In_495,In_864);
and U460 (N_460,In_590,In_488);
nand U461 (N_461,In_591,In_594);
or U462 (N_462,In_218,In_362);
nand U463 (N_463,In_510,In_896);
nand U464 (N_464,In_53,In_565);
or U465 (N_465,In_365,In_93);
nand U466 (N_466,In_649,In_659);
nor U467 (N_467,In_255,In_667);
and U468 (N_468,In_883,In_801);
or U469 (N_469,In_763,In_159);
and U470 (N_470,In_328,In_499);
and U471 (N_471,In_342,In_653);
nand U472 (N_472,In_152,In_489);
and U473 (N_473,In_784,In_22);
nor U474 (N_474,In_906,In_730);
or U475 (N_475,In_484,In_443);
xnor U476 (N_476,In_704,In_267);
nor U477 (N_477,In_995,In_703);
or U478 (N_478,In_934,In_982);
nor U479 (N_479,In_779,In_860);
nand U480 (N_480,In_890,In_799);
or U481 (N_481,In_178,In_167);
and U482 (N_482,In_829,In_280);
nand U483 (N_483,In_528,In_807);
or U484 (N_484,In_321,In_64);
nand U485 (N_485,In_977,In_359);
or U486 (N_486,In_153,In_856);
or U487 (N_487,In_872,In_922);
or U488 (N_488,In_231,In_193);
and U489 (N_489,In_106,In_713);
and U490 (N_490,In_266,In_785);
nor U491 (N_491,In_68,In_921);
nand U492 (N_492,In_581,In_998);
or U493 (N_493,In_363,In_0);
nand U494 (N_494,In_405,In_868);
and U495 (N_495,In_97,In_354);
and U496 (N_496,In_803,In_139);
or U497 (N_497,In_62,In_790);
and U498 (N_498,In_961,In_944);
nand U499 (N_499,In_370,In_716);
and U500 (N_500,In_238,In_552);
nand U501 (N_501,In_757,In_827);
xnor U502 (N_502,In_84,In_40);
and U503 (N_503,In_207,In_286);
nand U504 (N_504,In_587,In_627);
and U505 (N_505,In_848,In_497);
or U506 (N_506,In_561,In_988);
and U507 (N_507,In_108,In_240);
or U508 (N_508,In_621,In_391);
nor U509 (N_509,In_566,In_155);
nand U510 (N_510,In_215,In_512);
and U511 (N_511,In_377,In_895);
or U512 (N_512,In_753,In_298);
and U513 (N_513,In_934,In_936);
xor U514 (N_514,In_533,In_802);
nor U515 (N_515,In_221,In_138);
or U516 (N_516,In_357,In_225);
and U517 (N_517,In_956,In_811);
and U518 (N_518,In_31,In_882);
nor U519 (N_519,In_883,In_721);
nand U520 (N_520,In_283,In_460);
or U521 (N_521,In_718,In_963);
and U522 (N_522,In_976,In_558);
or U523 (N_523,In_574,In_653);
and U524 (N_524,In_115,In_308);
and U525 (N_525,In_147,In_459);
and U526 (N_526,In_606,In_884);
and U527 (N_527,In_836,In_357);
and U528 (N_528,In_473,In_890);
or U529 (N_529,In_510,In_743);
or U530 (N_530,In_188,In_95);
xor U531 (N_531,In_112,In_398);
nand U532 (N_532,In_876,In_489);
nand U533 (N_533,In_188,In_246);
nand U534 (N_534,In_595,In_861);
and U535 (N_535,In_334,In_651);
nor U536 (N_536,In_545,In_396);
xnor U537 (N_537,In_88,In_509);
or U538 (N_538,In_30,In_2);
nand U539 (N_539,In_443,In_659);
and U540 (N_540,In_269,In_878);
or U541 (N_541,In_542,In_768);
and U542 (N_542,In_856,In_891);
and U543 (N_543,In_132,In_857);
or U544 (N_544,In_205,In_163);
nor U545 (N_545,In_252,In_566);
or U546 (N_546,In_256,In_504);
nand U547 (N_547,In_510,In_46);
or U548 (N_548,In_817,In_33);
nor U549 (N_549,In_636,In_822);
and U550 (N_550,In_29,In_155);
nor U551 (N_551,In_191,In_639);
nor U552 (N_552,In_42,In_76);
nand U553 (N_553,In_35,In_328);
or U554 (N_554,In_649,In_796);
nor U555 (N_555,In_922,In_841);
nor U556 (N_556,In_875,In_392);
or U557 (N_557,In_679,In_653);
nor U558 (N_558,In_197,In_308);
and U559 (N_559,In_745,In_968);
or U560 (N_560,In_313,In_438);
and U561 (N_561,In_43,In_214);
nor U562 (N_562,In_80,In_246);
or U563 (N_563,In_269,In_539);
or U564 (N_564,In_627,In_611);
nand U565 (N_565,In_673,In_65);
nand U566 (N_566,In_907,In_973);
or U567 (N_567,In_419,In_152);
nor U568 (N_568,In_381,In_423);
and U569 (N_569,In_242,In_758);
and U570 (N_570,In_711,In_146);
and U571 (N_571,In_935,In_142);
nand U572 (N_572,In_427,In_80);
and U573 (N_573,In_668,In_997);
and U574 (N_574,In_743,In_235);
nand U575 (N_575,In_495,In_366);
and U576 (N_576,In_778,In_346);
or U577 (N_577,In_231,In_256);
and U578 (N_578,In_441,In_973);
and U579 (N_579,In_545,In_511);
and U580 (N_580,In_8,In_84);
nor U581 (N_581,In_912,In_819);
nand U582 (N_582,In_829,In_401);
nor U583 (N_583,In_69,In_217);
nand U584 (N_584,In_849,In_972);
and U585 (N_585,In_149,In_701);
nand U586 (N_586,In_87,In_965);
nand U587 (N_587,In_379,In_328);
nor U588 (N_588,In_82,In_593);
and U589 (N_589,In_804,In_468);
nand U590 (N_590,In_247,In_306);
and U591 (N_591,In_910,In_320);
or U592 (N_592,In_176,In_593);
and U593 (N_593,In_398,In_690);
and U594 (N_594,In_441,In_127);
or U595 (N_595,In_770,In_995);
or U596 (N_596,In_993,In_709);
and U597 (N_597,In_161,In_485);
or U598 (N_598,In_465,In_757);
and U599 (N_599,In_821,In_395);
and U600 (N_600,In_330,In_695);
nand U601 (N_601,In_182,In_400);
or U602 (N_602,In_583,In_669);
and U603 (N_603,In_99,In_349);
nor U604 (N_604,In_167,In_40);
and U605 (N_605,In_291,In_166);
nand U606 (N_606,In_234,In_907);
and U607 (N_607,In_182,In_281);
or U608 (N_608,In_6,In_984);
nor U609 (N_609,In_499,In_799);
nand U610 (N_610,In_137,In_734);
nor U611 (N_611,In_746,In_619);
or U612 (N_612,In_683,In_830);
and U613 (N_613,In_498,In_233);
nor U614 (N_614,In_775,In_685);
nand U615 (N_615,In_247,In_42);
and U616 (N_616,In_437,In_674);
nor U617 (N_617,In_33,In_521);
nand U618 (N_618,In_934,In_626);
nor U619 (N_619,In_838,In_8);
nor U620 (N_620,In_212,In_747);
nand U621 (N_621,In_16,In_748);
nand U622 (N_622,In_835,In_451);
and U623 (N_623,In_237,In_462);
nor U624 (N_624,In_573,In_549);
and U625 (N_625,In_907,In_0);
and U626 (N_626,In_567,In_300);
nand U627 (N_627,In_226,In_957);
or U628 (N_628,In_661,In_21);
or U629 (N_629,In_136,In_975);
and U630 (N_630,In_896,In_681);
nand U631 (N_631,In_668,In_890);
nand U632 (N_632,In_790,In_492);
and U633 (N_633,In_149,In_697);
and U634 (N_634,In_611,In_983);
or U635 (N_635,In_820,In_120);
and U636 (N_636,In_740,In_990);
or U637 (N_637,In_693,In_174);
nor U638 (N_638,In_929,In_281);
nand U639 (N_639,In_298,In_635);
and U640 (N_640,In_47,In_879);
nor U641 (N_641,In_644,In_590);
nor U642 (N_642,In_378,In_43);
nor U643 (N_643,In_614,In_240);
or U644 (N_644,In_867,In_405);
or U645 (N_645,In_958,In_599);
nand U646 (N_646,In_963,In_322);
nor U647 (N_647,In_660,In_344);
nand U648 (N_648,In_86,In_921);
nor U649 (N_649,In_96,In_543);
nor U650 (N_650,In_174,In_116);
or U651 (N_651,In_516,In_681);
and U652 (N_652,In_165,In_754);
and U653 (N_653,In_303,In_405);
and U654 (N_654,In_252,In_428);
nand U655 (N_655,In_667,In_555);
and U656 (N_656,In_51,In_370);
nor U657 (N_657,In_829,In_490);
nor U658 (N_658,In_406,In_829);
nor U659 (N_659,In_239,In_893);
and U660 (N_660,In_401,In_0);
nand U661 (N_661,In_683,In_487);
and U662 (N_662,In_51,In_40);
or U663 (N_663,In_444,In_727);
xnor U664 (N_664,In_824,In_676);
nor U665 (N_665,In_771,In_556);
or U666 (N_666,In_444,In_821);
or U667 (N_667,In_930,In_277);
and U668 (N_668,In_746,In_255);
or U669 (N_669,In_932,In_569);
nand U670 (N_670,In_638,In_942);
nor U671 (N_671,In_666,In_98);
and U672 (N_672,In_887,In_158);
and U673 (N_673,In_83,In_49);
nor U674 (N_674,In_330,In_944);
or U675 (N_675,In_292,In_911);
nand U676 (N_676,In_721,In_109);
nand U677 (N_677,In_314,In_538);
and U678 (N_678,In_30,In_315);
and U679 (N_679,In_551,In_973);
nand U680 (N_680,In_272,In_311);
or U681 (N_681,In_738,In_53);
nand U682 (N_682,In_61,In_566);
or U683 (N_683,In_297,In_283);
or U684 (N_684,In_328,In_16);
and U685 (N_685,In_351,In_831);
xor U686 (N_686,In_810,In_320);
or U687 (N_687,In_222,In_849);
nand U688 (N_688,In_85,In_351);
and U689 (N_689,In_159,In_352);
nor U690 (N_690,In_323,In_805);
nand U691 (N_691,In_504,In_976);
nor U692 (N_692,In_328,In_588);
nor U693 (N_693,In_463,In_234);
nand U694 (N_694,In_682,In_142);
or U695 (N_695,In_913,In_225);
or U696 (N_696,In_450,In_142);
and U697 (N_697,In_413,In_534);
nand U698 (N_698,In_870,In_970);
nor U699 (N_699,In_124,In_303);
nand U700 (N_700,In_493,In_232);
nand U701 (N_701,In_233,In_410);
or U702 (N_702,In_512,In_117);
nor U703 (N_703,In_993,In_84);
or U704 (N_704,In_346,In_897);
or U705 (N_705,In_520,In_624);
and U706 (N_706,In_788,In_412);
or U707 (N_707,In_255,In_72);
nand U708 (N_708,In_961,In_222);
and U709 (N_709,In_886,In_870);
and U710 (N_710,In_654,In_485);
and U711 (N_711,In_141,In_226);
or U712 (N_712,In_966,In_712);
and U713 (N_713,In_415,In_950);
or U714 (N_714,In_314,In_792);
or U715 (N_715,In_493,In_135);
and U716 (N_716,In_449,In_662);
nand U717 (N_717,In_129,In_295);
or U718 (N_718,In_951,In_122);
nand U719 (N_719,In_704,In_785);
and U720 (N_720,In_612,In_650);
and U721 (N_721,In_222,In_591);
or U722 (N_722,In_567,In_283);
nor U723 (N_723,In_734,In_818);
and U724 (N_724,In_854,In_749);
or U725 (N_725,In_674,In_567);
nand U726 (N_726,In_816,In_572);
and U727 (N_727,In_112,In_417);
xnor U728 (N_728,In_995,In_266);
and U729 (N_729,In_486,In_529);
nand U730 (N_730,In_652,In_493);
and U731 (N_731,In_695,In_20);
or U732 (N_732,In_126,In_886);
and U733 (N_733,In_395,In_918);
nand U734 (N_734,In_592,In_927);
nor U735 (N_735,In_597,In_436);
nor U736 (N_736,In_710,In_892);
and U737 (N_737,In_511,In_33);
and U738 (N_738,In_370,In_831);
nor U739 (N_739,In_920,In_932);
and U740 (N_740,In_442,In_33);
and U741 (N_741,In_899,In_158);
and U742 (N_742,In_705,In_394);
nor U743 (N_743,In_282,In_373);
and U744 (N_744,In_723,In_542);
xnor U745 (N_745,In_525,In_13);
and U746 (N_746,In_722,In_58);
nor U747 (N_747,In_724,In_540);
nor U748 (N_748,In_744,In_508);
nor U749 (N_749,In_611,In_887);
nand U750 (N_750,In_557,In_559);
nor U751 (N_751,In_454,In_783);
and U752 (N_752,In_183,In_464);
and U753 (N_753,In_489,In_838);
or U754 (N_754,In_819,In_604);
and U755 (N_755,In_994,In_295);
nand U756 (N_756,In_999,In_574);
and U757 (N_757,In_979,In_595);
and U758 (N_758,In_958,In_949);
nor U759 (N_759,In_681,In_383);
or U760 (N_760,In_526,In_759);
and U761 (N_761,In_404,In_662);
nand U762 (N_762,In_366,In_253);
or U763 (N_763,In_64,In_95);
or U764 (N_764,In_595,In_285);
and U765 (N_765,In_958,In_876);
or U766 (N_766,In_17,In_648);
and U767 (N_767,In_663,In_953);
or U768 (N_768,In_27,In_42);
nand U769 (N_769,In_689,In_156);
nand U770 (N_770,In_446,In_798);
nor U771 (N_771,In_129,In_126);
or U772 (N_772,In_193,In_880);
nor U773 (N_773,In_170,In_965);
nand U774 (N_774,In_877,In_842);
or U775 (N_775,In_152,In_771);
and U776 (N_776,In_203,In_165);
and U777 (N_777,In_259,In_849);
or U778 (N_778,In_939,In_108);
or U779 (N_779,In_352,In_679);
and U780 (N_780,In_753,In_563);
nand U781 (N_781,In_874,In_344);
or U782 (N_782,In_443,In_26);
and U783 (N_783,In_68,In_394);
and U784 (N_784,In_350,In_299);
nand U785 (N_785,In_716,In_118);
nor U786 (N_786,In_344,In_183);
or U787 (N_787,In_971,In_497);
nor U788 (N_788,In_7,In_8);
or U789 (N_789,In_718,In_951);
nor U790 (N_790,In_452,In_975);
and U791 (N_791,In_618,In_289);
nor U792 (N_792,In_701,In_486);
or U793 (N_793,In_976,In_435);
nand U794 (N_794,In_979,In_87);
nand U795 (N_795,In_228,In_879);
nand U796 (N_796,In_496,In_831);
and U797 (N_797,In_213,In_574);
and U798 (N_798,In_117,In_768);
nand U799 (N_799,In_828,In_930);
nand U800 (N_800,In_535,In_385);
nor U801 (N_801,In_984,In_72);
and U802 (N_802,In_127,In_885);
and U803 (N_803,In_438,In_186);
nor U804 (N_804,In_695,In_315);
nand U805 (N_805,In_536,In_993);
nor U806 (N_806,In_521,In_544);
and U807 (N_807,In_36,In_369);
and U808 (N_808,In_450,In_343);
or U809 (N_809,In_91,In_180);
nor U810 (N_810,In_412,In_842);
or U811 (N_811,In_602,In_307);
and U812 (N_812,In_425,In_478);
nor U813 (N_813,In_81,In_959);
nand U814 (N_814,In_43,In_116);
nor U815 (N_815,In_649,In_197);
or U816 (N_816,In_720,In_284);
or U817 (N_817,In_2,In_122);
nand U818 (N_818,In_42,In_704);
or U819 (N_819,In_794,In_645);
nor U820 (N_820,In_352,In_387);
or U821 (N_821,In_924,In_157);
nand U822 (N_822,In_178,In_777);
nand U823 (N_823,In_308,In_868);
or U824 (N_824,In_391,In_160);
and U825 (N_825,In_311,In_389);
and U826 (N_826,In_438,In_945);
nor U827 (N_827,In_714,In_361);
or U828 (N_828,In_671,In_383);
and U829 (N_829,In_70,In_897);
or U830 (N_830,In_156,In_813);
or U831 (N_831,In_784,In_144);
nand U832 (N_832,In_849,In_536);
or U833 (N_833,In_595,In_310);
nand U834 (N_834,In_390,In_258);
and U835 (N_835,In_400,In_749);
and U836 (N_836,In_111,In_217);
nor U837 (N_837,In_176,In_453);
nand U838 (N_838,In_816,In_28);
and U839 (N_839,In_250,In_962);
and U840 (N_840,In_689,In_339);
or U841 (N_841,In_44,In_941);
nand U842 (N_842,In_883,In_984);
nor U843 (N_843,In_630,In_876);
nand U844 (N_844,In_275,In_142);
and U845 (N_845,In_540,In_745);
nand U846 (N_846,In_225,In_158);
nand U847 (N_847,In_455,In_225);
nand U848 (N_848,In_546,In_688);
nor U849 (N_849,In_748,In_623);
nand U850 (N_850,In_138,In_959);
or U851 (N_851,In_565,In_635);
or U852 (N_852,In_212,In_451);
nor U853 (N_853,In_549,In_68);
nor U854 (N_854,In_16,In_973);
nand U855 (N_855,In_287,In_707);
nand U856 (N_856,In_703,In_384);
nor U857 (N_857,In_4,In_202);
nand U858 (N_858,In_761,In_235);
nor U859 (N_859,In_20,In_326);
nor U860 (N_860,In_120,In_898);
nand U861 (N_861,In_287,In_824);
and U862 (N_862,In_423,In_590);
nand U863 (N_863,In_515,In_762);
and U864 (N_864,In_764,In_451);
and U865 (N_865,In_364,In_77);
nand U866 (N_866,In_936,In_316);
nand U867 (N_867,In_15,In_896);
and U868 (N_868,In_126,In_697);
nor U869 (N_869,In_220,In_975);
or U870 (N_870,In_3,In_120);
nor U871 (N_871,In_139,In_64);
or U872 (N_872,In_485,In_302);
and U873 (N_873,In_620,In_744);
nor U874 (N_874,In_594,In_686);
and U875 (N_875,In_499,In_864);
and U876 (N_876,In_951,In_918);
nor U877 (N_877,In_572,In_220);
nand U878 (N_878,In_490,In_945);
or U879 (N_879,In_534,In_752);
nand U880 (N_880,In_433,In_498);
nand U881 (N_881,In_954,In_226);
and U882 (N_882,In_330,In_674);
nor U883 (N_883,In_545,In_342);
nor U884 (N_884,In_9,In_69);
xnor U885 (N_885,In_416,In_677);
or U886 (N_886,In_629,In_449);
nor U887 (N_887,In_534,In_669);
xnor U888 (N_888,In_198,In_90);
nand U889 (N_889,In_702,In_332);
nand U890 (N_890,In_874,In_312);
nor U891 (N_891,In_187,In_689);
and U892 (N_892,In_209,In_112);
and U893 (N_893,In_766,In_459);
and U894 (N_894,In_931,In_649);
and U895 (N_895,In_330,In_561);
or U896 (N_896,In_16,In_153);
and U897 (N_897,In_68,In_103);
and U898 (N_898,In_499,In_972);
and U899 (N_899,In_622,In_514);
or U900 (N_900,In_540,In_458);
nor U901 (N_901,In_426,In_792);
or U902 (N_902,In_678,In_701);
nand U903 (N_903,In_911,In_669);
and U904 (N_904,In_478,In_409);
and U905 (N_905,In_695,In_156);
nor U906 (N_906,In_754,In_604);
or U907 (N_907,In_728,In_974);
or U908 (N_908,In_375,In_42);
nand U909 (N_909,In_95,In_849);
nor U910 (N_910,In_199,In_67);
nand U911 (N_911,In_466,In_679);
or U912 (N_912,In_292,In_584);
nand U913 (N_913,In_777,In_704);
or U914 (N_914,In_317,In_603);
or U915 (N_915,In_286,In_414);
or U916 (N_916,In_323,In_164);
or U917 (N_917,In_736,In_490);
and U918 (N_918,In_630,In_5);
nand U919 (N_919,In_477,In_408);
nand U920 (N_920,In_496,In_842);
and U921 (N_921,In_178,In_502);
nor U922 (N_922,In_696,In_532);
nand U923 (N_923,In_72,In_826);
and U924 (N_924,In_941,In_765);
and U925 (N_925,In_225,In_312);
and U926 (N_926,In_38,In_239);
and U927 (N_927,In_679,In_944);
and U928 (N_928,In_110,In_287);
nor U929 (N_929,In_635,In_152);
nor U930 (N_930,In_928,In_893);
nand U931 (N_931,In_419,In_109);
or U932 (N_932,In_361,In_868);
and U933 (N_933,In_857,In_505);
and U934 (N_934,In_316,In_431);
or U935 (N_935,In_807,In_433);
nand U936 (N_936,In_782,In_118);
nor U937 (N_937,In_594,In_576);
nand U938 (N_938,In_435,In_259);
nor U939 (N_939,In_551,In_952);
nor U940 (N_940,In_268,In_264);
or U941 (N_941,In_770,In_293);
nor U942 (N_942,In_73,In_666);
nand U943 (N_943,In_757,In_631);
nand U944 (N_944,In_6,In_611);
nand U945 (N_945,In_483,In_870);
nor U946 (N_946,In_695,In_96);
nor U947 (N_947,In_440,In_590);
nand U948 (N_948,In_607,In_837);
or U949 (N_949,In_695,In_579);
nand U950 (N_950,In_116,In_307);
nor U951 (N_951,In_64,In_533);
nor U952 (N_952,In_527,In_426);
and U953 (N_953,In_283,In_423);
nand U954 (N_954,In_416,In_39);
nor U955 (N_955,In_600,In_740);
and U956 (N_956,In_789,In_527);
or U957 (N_957,In_958,In_154);
or U958 (N_958,In_380,In_94);
nand U959 (N_959,In_126,In_272);
nand U960 (N_960,In_819,In_286);
or U961 (N_961,In_826,In_708);
or U962 (N_962,In_10,In_193);
and U963 (N_963,In_415,In_423);
and U964 (N_964,In_648,In_948);
nand U965 (N_965,In_808,In_385);
and U966 (N_966,In_906,In_792);
nand U967 (N_967,In_979,In_422);
nor U968 (N_968,In_728,In_779);
nand U969 (N_969,In_132,In_883);
and U970 (N_970,In_294,In_493);
nand U971 (N_971,In_586,In_73);
nand U972 (N_972,In_131,In_305);
nand U973 (N_973,In_731,In_582);
and U974 (N_974,In_752,In_765);
or U975 (N_975,In_843,In_889);
nand U976 (N_976,In_380,In_647);
nand U977 (N_977,In_945,In_18);
and U978 (N_978,In_61,In_316);
and U979 (N_979,In_73,In_193);
and U980 (N_980,In_366,In_553);
nand U981 (N_981,In_103,In_282);
nor U982 (N_982,In_752,In_656);
and U983 (N_983,In_501,In_707);
and U984 (N_984,In_946,In_412);
nor U985 (N_985,In_146,In_886);
nor U986 (N_986,In_419,In_649);
and U987 (N_987,In_697,In_452);
and U988 (N_988,In_599,In_279);
and U989 (N_989,In_350,In_481);
nor U990 (N_990,In_284,In_403);
nand U991 (N_991,In_727,In_924);
or U992 (N_992,In_297,In_722);
nand U993 (N_993,In_812,In_617);
nor U994 (N_994,In_232,In_527);
and U995 (N_995,In_646,In_350);
nand U996 (N_996,In_139,In_299);
and U997 (N_997,In_835,In_386);
nor U998 (N_998,In_0,In_652);
and U999 (N_999,In_603,In_386);
nand U1000 (N_1000,N_389,N_256);
or U1001 (N_1001,N_843,N_957);
or U1002 (N_1002,N_665,N_833);
or U1003 (N_1003,N_262,N_537);
nand U1004 (N_1004,N_752,N_917);
nand U1005 (N_1005,N_453,N_188);
nor U1006 (N_1006,N_786,N_557);
and U1007 (N_1007,N_423,N_189);
and U1008 (N_1008,N_754,N_133);
nand U1009 (N_1009,N_2,N_689);
or U1010 (N_1010,N_125,N_456);
nor U1011 (N_1011,N_599,N_912);
nor U1012 (N_1012,N_675,N_584);
xor U1013 (N_1013,N_885,N_919);
or U1014 (N_1014,N_753,N_911);
and U1015 (N_1015,N_305,N_749);
nand U1016 (N_1016,N_949,N_964);
or U1017 (N_1017,N_445,N_197);
or U1018 (N_1018,N_535,N_914);
nand U1019 (N_1019,N_386,N_206);
and U1020 (N_1020,N_935,N_761);
or U1021 (N_1021,N_996,N_924);
and U1022 (N_1022,N_551,N_569);
nor U1023 (N_1023,N_104,N_37);
or U1024 (N_1024,N_866,N_764);
nand U1025 (N_1025,N_598,N_940);
and U1026 (N_1026,N_883,N_208);
and U1027 (N_1027,N_713,N_524);
or U1028 (N_1028,N_719,N_162);
or U1029 (N_1029,N_775,N_172);
nand U1030 (N_1030,N_857,N_154);
nand U1031 (N_1031,N_650,N_659);
and U1032 (N_1032,N_789,N_132);
nor U1033 (N_1033,N_717,N_48);
and U1034 (N_1034,N_120,N_332);
or U1035 (N_1035,N_449,N_576);
and U1036 (N_1036,N_552,N_800);
nand U1037 (N_1037,N_871,N_634);
or U1038 (N_1038,N_331,N_491);
nand U1039 (N_1039,N_304,N_908);
nand U1040 (N_1040,N_874,N_784);
or U1041 (N_1041,N_954,N_341);
or U1042 (N_1042,N_235,N_321);
nand U1043 (N_1043,N_745,N_258);
nand U1044 (N_1044,N_54,N_284);
nor U1045 (N_1045,N_270,N_968);
and U1046 (N_1046,N_110,N_203);
and U1047 (N_1047,N_296,N_907);
and U1048 (N_1048,N_399,N_47);
or U1049 (N_1049,N_149,N_865);
nand U1050 (N_1050,N_329,N_268);
nand U1051 (N_1051,N_625,N_404);
nand U1052 (N_1052,N_999,N_716);
or U1053 (N_1053,N_187,N_226);
nor U1054 (N_1054,N_704,N_131);
or U1055 (N_1055,N_565,N_152);
nor U1056 (N_1056,N_623,N_632);
or U1057 (N_1057,N_813,N_680);
and U1058 (N_1058,N_0,N_35);
nand U1059 (N_1059,N_830,N_867);
nor U1060 (N_1060,N_477,N_394);
and U1061 (N_1061,N_53,N_556);
and U1062 (N_1062,N_220,N_910);
or U1063 (N_1063,N_45,N_333);
or U1064 (N_1064,N_246,N_604);
or U1065 (N_1065,N_820,N_315);
nor U1066 (N_1066,N_359,N_266);
nor U1067 (N_1067,N_514,N_84);
nor U1068 (N_1068,N_750,N_488);
and U1069 (N_1069,N_506,N_610);
nand U1070 (N_1070,N_111,N_701);
nand U1071 (N_1071,N_578,N_723);
nor U1072 (N_1072,N_442,N_878);
nor U1073 (N_1073,N_517,N_854);
and U1074 (N_1074,N_970,N_976);
and U1075 (N_1075,N_771,N_592);
or U1076 (N_1076,N_762,N_290);
nor U1077 (N_1077,N_714,N_734);
or U1078 (N_1078,N_763,N_906);
and U1079 (N_1079,N_356,N_620);
nand U1080 (N_1080,N_799,N_895);
nand U1081 (N_1081,N_402,N_654);
or U1082 (N_1082,N_903,N_112);
nor U1083 (N_1083,N_21,N_894);
nand U1084 (N_1084,N_580,N_192);
and U1085 (N_1085,N_371,N_840);
nor U1086 (N_1086,N_748,N_265);
or U1087 (N_1087,N_463,N_715);
and U1088 (N_1088,N_500,N_85);
nor U1089 (N_1089,N_845,N_222);
or U1090 (N_1090,N_978,N_64);
nand U1091 (N_1091,N_168,N_902);
nand U1092 (N_1092,N_278,N_231);
or U1093 (N_1093,N_340,N_959);
nand U1094 (N_1094,N_336,N_482);
nor U1095 (N_1095,N_109,N_554);
nor U1096 (N_1096,N_57,N_502);
or U1097 (N_1097,N_496,N_484);
nor U1098 (N_1098,N_90,N_615);
nand U1099 (N_1099,N_160,N_76);
nor U1100 (N_1100,N_746,N_436);
or U1101 (N_1101,N_52,N_633);
and U1102 (N_1102,N_264,N_915);
nand U1103 (N_1103,N_619,N_309);
nor U1104 (N_1104,N_405,N_718);
or U1105 (N_1105,N_791,N_9);
and U1106 (N_1106,N_898,N_916);
nand U1107 (N_1107,N_648,N_147);
or U1108 (N_1108,N_124,N_43);
nor U1109 (N_1109,N_119,N_848);
nand U1110 (N_1110,N_828,N_319);
or U1111 (N_1111,N_663,N_859);
nand U1112 (N_1112,N_26,N_728);
and U1113 (N_1113,N_96,N_966);
nand U1114 (N_1114,N_587,N_881);
and U1115 (N_1115,N_175,N_13);
nand U1116 (N_1116,N_641,N_825);
and U1117 (N_1117,N_115,N_400);
nor U1118 (N_1118,N_536,N_148);
nor U1119 (N_1119,N_367,N_1);
or U1120 (N_1120,N_370,N_299);
and U1121 (N_1121,N_581,N_59);
and U1122 (N_1122,N_541,N_932);
nor U1123 (N_1123,N_695,N_727);
or U1124 (N_1124,N_724,N_548);
nand U1125 (N_1125,N_920,N_640);
nor U1126 (N_1126,N_409,N_937);
and U1127 (N_1127,N_489,N_794);
or U1128 (N_1128,N_328,N_655);
and U1129 (N_1129,N_563,N_68);
or U1130 (N_1130,N_652,N_292);
nand U1131 (N_1131,N_571,N_236);
nor U1132 (N_1132,N_944,N_74);
nor U1133 (N_1133,N_91,N_67);
nand U1134 (N_1134,N_71,N_317);
nor U1135 (N_1135,N_239,N_138);
or U1136 (N_1136,N_550,N_721);
and U1137 (N_1137,N_585,N_46);
nor U1138 (N_1138,N_905,N_269);
nand U1139 (N_1139,N_480,N_614);
and U1140 (N_1140,N_165,N_674);
and U1141 (N_1141,N_681,N_447);
or U1142 (N_1142,N_969,N_824);
nor U1143 (N_1143,N_60,N_17);
or U1144 (N_1144,N_956,N_822);
nor U1145 (N_1145,N_72,N_286);
nand U1146 (N_1146,N_766,N_291);
nor U1147 (N_1147,N_989,N_980);
nor U1148 (N_1148,N_238,N_692);
nand U1149 (N_1149,N_401,N_280);
or U1150 (N_1150,N_186,N_39);
nor U1151 (N_1151,N_275,N_428);
and U1152 (N_1152,N_967,N_863);
nand U1153 (N_1153,N_676,N_839);
nor U1154 (N_1154,N_30,N_851);
nor U1155 (N_1155,N_841,N_391);
nor U1156 (N_1156,N_973,N_872);
or U1157 (N_1157,N_758,N_708);
or U1158 (N_1158,N_519,N_145);
and U1159 (N_1159,N_855,N_809);
and U1160 (N_1160,N_568,N_136);
or U1161 (N_1161,N_815,N_322);
or U1162 (N_1162,N_808,N_483);
nand U1163 (N_1163,N_942,N_215);
nand U1164 (N_1164,N_744,N_923);
nand U1165 (N_1165,N_785,N_756);
nor U1166 (N_1166,N_80,N_586);
nand U1167 (N_1167,N_913,N_591);
nand U1168 (N_1168,N_693,N_507);
and U1169 (N_1169,N_156,N_129);
and U1170 (N_1170,N_459,N_948);
or U1171 (N_1171,N_107,N_850);
and U1172 (N_1172,N_971,N_547);
or U1173 (N_1173,N_510,N_559);
nor U1174 (N_1174,N_433,N_657);
or U1175 (N_1175,N_142,N_575);
and U1176 (N_1176,N_922,N_879);
or U1177 (N_1177,N_558,N_995);
or U1178 (N_1178,N_630,N_732);
nand U1179 (N_1179,N_376,N_972);
nor U1180 (N_1180,N_34,N_475);
or U1181 (N_1181,N_670,N_274);
xor U1182 (N_1182,N_958,N_116);
and U1183 (N_1183,N_56,N_667);
nand U1184 (N_1184,N_14,N_691);
nand U1185 (N_1185,N_382,N_737);
nor U1186 (N_1186,N_306,N_298);
nor U1187 (N_1187,N_358,N_330);
and U1188 (N_1188,N_62,N_457);
nand U1189 (N_1189,N_993,N_271);
or U1190 (N_1190,N_934,N_49);
or U1191 (N_1191,N_658,N_918);
nor U1192 (N_1192,N_823,N_590);
and U1193 (N_1193,N_960,N_117);
nand U1194 (N_1194,N_22,N_896);
or U1195 (N_1195,N_395,N_255);
nor U1196 (N_1196,N_3,N_144);
or U1197 (N_1197,N_832,N_501);
nor U1198 (N_1198,N_860,N_503);
and U1199 (N_1199,N_807,N_101);
and U1200 (N_1200,N_438,N_928);
and U1201 (N_1201,N_97,N_643);
or U1202 (N_1202,N_415,N_28);
or U1203 (N_1203,N_444,N_962);
nand U1204 (N_1204,N_351,N_406);
nor U1205 (N_1205,N_601,N_703);
or U1206 (N_1206,N_312,N_529);
nor U1207 (N_1207,N_801,N_323);
or U1208 (N_1208,N_849,N_221);
or U1209 (N_1209,N_555,N_837);
or U1210 (N_1210,N_466,N_32);
nand U1211 (N_1211,N_261,N_364);
nor U1212 (N_1212,N_666,N_486);
nand U1213 (N_1213,N_873,N_983);
nand U1214 (N_1214,N_864,N_781);
nand U1215 (N_1215,N_185,N_245);
nor U1216 (N_1216,N_248,N_396);
and U1217 (N_1217,N_530,N_326);
nor U1218 (N_1218,N_41,N_526);
or U1219 (N_1219,N_617,N_412);
and U1220 (N_1220,N_253,N_900);
nor U1221 (N_1221,N_403,N_320);
nor U1222 (N_1222,N_847,N_65);
and U1223 (N_1223,N_465,N_314);
nand U1224 (N_1224,N_660,N_69);
and U1225 (N_1225,N_527,N_285);
or U1226 (N_1226,N_40,N_181);
and U1227 (N_1227,N_884,N_776);
nand U1228 (N_1228,N_953,N_595);
or U1229 (N_1229,N_137,N_738);
nor U1230 (N_1230,N_730,N_515);
nand U1231 (N_1231,N_342,N_739);
nor U1232 (N_1232,N_720,N_982);
and U1233 (N_1233,N_542,N_656);
xnor U1234 (N_1234,N_612,N_20);
nand U1235 (N_1235,N_696,N_780);
and U1236 (N_1236,N_408,N_725);
nor U1237 (N_1237,N_325,N_366);
and U1238 (N_1238,N_435,N_504);
and U1239 (N_1239,N_38,N_250);
nor U1240 (N_1240,N_493,N_741);
nand U1241 (N_1241,N_505,N_15);
nor U1242 (N_1242,N_86,N_796);
nand U1243 (N_1243,N_627,N_687);
nor U1244 (N_1244,N_207,N_930);
nor U1245 (N_1245,N_887,N_194);
or U1246 (N_1246,N_88,N_698);
and U1247 (N_1247,N_407,N_988);
nor U1248 (N_1248,N_19,N_51);
or U1249 (N_1249,N_77,N_779);
or U1250 (N_1250,N_307,N_310);
and U1251 (N_1251,N_205,N_577);
nor U1252 (N_1252,N_182,N_212);
or U1253 (N_1253,N_434,N_974);
nor U1254 (N_1254,N_827,N_143);
nand U1255 (N_1255,N_603,N_499);
nand U1256 (N_1256,N_157,N_417);
nand U1257 (N_1257,N_567,N_856);
and U1258 (N_1258,N_368,N_705);
nand U1259 (N_1259,N_965,N_316);
nor U1260 (N_1260,N_668,N_994);
or U1261 (N_1261,N_963,N_852);
or U1262 (N_1262,N_726,N_36);
nor U1263 (N_1263,N_826,N_777);
and U1264 (N_1264,N_227,N_685);
nor U1265 (N_1265,N_198,N_237);
and U1266 (N_1266,N_904,N_452);
and U1267 (N_1267,N_230,N_936);
xor U1268 (N_1268,N_209,N_446);
nand U1269 (N_1269,N_429,N_199);
nand U1270 (N_1270,N_219,N_254);
xor U1271 (N_1271,N_75,N_78);
nand U1272 (N_1272,N_594,N_6);
or U1273 (N_1273,N_50,N_882);
nor U1274 (N_1274,N_909,N_398);
nor U1275 (N_1275,N_579,N_276);
nand U1276 (N_1276,N_113,N_294);
and U1277 (N_1277,N_606,N_374);
nand U1278 (N_1278,N_740,N_939);
and U1279 (N_1279,N_862,N_931);
nand U1280 (N_1280,N_516,N_961);
or U1281 (N_1281,N_573,N_164);
nor U1282 (N_1282,N_335,N_392);
or U1283 (N_1283,N_324,N_121);
nor U1284 (N_1284,N_73,N_211);
or U1285 (N_1285,N_25,N_393);
or U1286 (N_1286,N_544,N_492);
nand U1287 (N_1287,N_66,N_722);
nor U1288 (N_1288,N_252,N_362);
or U1289 (N_1289,N_348,N_427);
nor U1290 (N_1290,N_812,N_202);
or U1291 (N_1291,N_352,N_947);
nor U1292 (N_1292,N_540,N_490);
nand U1293 (N_1293,N_811,N_369);
or U1294 (N_1294,N_814,N_984);
or U1295 (N_1295,N_682,N_639);
or U1296 (N_1296,N_522,N_471);
and U1297 (N_1297,N_876,N_651);
and U1298 (N_1298,N_108,N_952);
and U1299 (N_1299,N_669,N_411);
and U1300 (N_1300,N_891,N_7);
nor U1301 (N_1301,N_139,N_539);
nor U1302 (N_1302,N_177,N_842);
nand U1303 (N_1303,N_699,N_24);
or U1304 (N_1304,N_562,N_345);
or U1305 (N_1305,N_63,N_282);
or U1306 (N_1306,N_773,N_134);
nand U1307 (N_1307,N_380,N_975);
nand U1308 (N_1308,N_831,N_778);
and U1309 (N_1309,N_170,N_118);
or U1310 (N_1310,N_729,N_945);
or U1311 (N_1311,N_191,N_479);
xnor U1312 (N_1312,N_998,N_834);
or U1313 (N_1313,N_163,N_93);
or U1314 (N_1314,N_613,N_512);
nand U1315 (N_1315,N_61,N_94);
or U1316 (N_1316,N_990,N_217);
nand U1317 (N_1317,N_570,N_293);
nor U1318 (N_1318,N_943,N_249);
and U1319 (N_1319,N_712,N_360);
nand U1320 (N_1320,N_283,N_12);
nand U1321 (N_1321,N_844,N_528);
or U1322 (N_1322,N_287,N_98);
nand U1323 (N_1323,N_99,N_783);
or U1324 (N_1324,N_508,N_127);
or U1325 (N_1325,N_337,N_810);
nand U1326 (N_1326,N_432,N_653);
nor U1327 (N_1327,N_802,N_161);
nand U1328 (N_1328,N_169,N_683);
nor U1329 (N_1329,N_277,N_677);
or U1330 (N_1330,N_173,N_247);
nand U1331 (N_1331,N_636,N_372);
and U1332 (N_1332,N_806,N_251);
and U1333 (N_1333,N_213,N_889);
nand U1334 (N_1334,N_572,N_214);
and U1335 (N_1335,N_263,N_986);
nor U1336 (N_1336,N_731,N_390);
nor U1337 (N_1337,N_183,N_821);
xnor U1338 (N_1338,N_135,N_769);
and U1339 (N_1339,N_228,N_350);
xor U1340 (N_1340,N_311,N_422);
nand U1341 (N_1341,N_941,N_673);
nand U1342 (N_1342,N_629,N_803);
nor U1343 (N_1343,N_538,N_804);
or U1344 (N_1344,N_901,N_128);
nand U1345 (N_1345,N_419,N_858);
and U1346 (N_1346,N_481,N_87);
or U1347 (N_1347,N_795,N_384);
and U1348 (N_1348,N_257,N_702);
and U1349 (N_1349,N_709,N_977);
and U1350 (N_1350,N_174,N_8);
or U1351 (N_1351,N_838,N_511);
nand U1352 (N_1352,N_520,N_819);
or U1353 (N_1353,N_464,N_431);
or U1354 (N_1354,N_338,N_546);
nor U1355 (N_1355,N_289,N_200);
or U1356 (N_1356,N_880,N_609);
or U1357 (N_1357,N_440,N_295);
nor U1358 (N_1358,N_458,N_760);
or U1359 (N_1359,N_755,N_597);
and U1360 (N_1360,N_103,N_997);
or U1361 (N_1361,N_588,N_624);
or U1362 (N_1362,N_818,N_743);
nand U1363 (N_1363,N_166,N_151);
nor U1364 (N_1364,N_987,N_532);
nand U1365 (N_1365,N_388,N_105);
nor U1366 (N_1366,N_545,N_664);
and U1367 (N_1367,N_241,N_229);
or U1368 (N_1368,N_621,N_950);
or U1369 (N_1369,N_846,N_711);
nor U1370 (N_1370,N_886,N_180);
nand U1371 (N_1371,N_622,N_593);
nor U1372 (N_1372,N_130,N_44);
xnor U1373 (N_1373,N_343,N_89);
or U1374 (N_1374,N_373,N_765);
nor U1375 (N_1375,N_608,N_159);
and U1376 (N_1376,N_561,N_979);
or U1377 (N_1377,N_985,N_448);
or U1378 (N_1378,N_353,N_981);
and U1379 (N_1379,N_533,N_835);
or U1380 (N_1380,N_589,N_757);
xor U1381 (N_1381,N_742,N_992);
nand U1382 (N_1382,N_600,N_684);
nand U1383 (N_1383,N_216,N_55);
nand U1384 (N_1384,N_176,N_123);
and U1385 (N_1385,N_272,N_141);
nor U1386 (N_1386,N_955,N_790);
and U1387 (N_1387,N_421,N_751);
and U1388 (N_1388,N_793,N_611);
and U1389 (N_1389,N_888,N_23);
nand U1390 (N_1390,N_497,N_383);
nor U1391 (N_1391,N_234,N_179);
nand U1392 (N_1392,N_626,N_853);
and U1393 (N_1393,N_596,N_153);
nor U1394 (N_1394,N_733,N_774);
nor U1395 (N_1395,N_4,N_167);
or U1396 (N_1396,N_193,N_210);
and U1397 (N_1397,N_574,N_279);
nor U1398 (N_1398,N_281,N_690);
nor U1399 (N_1399,N_470,N_455);
and U1400 (N_1400,N_355,N_897);
and U1401 (N_1401,N_642,N_645);
and U1402 (N_1402,N_646,N_425);
or U1403 (N_1403,N_543,N_787);
and U1404 (N_1404,N_672,N_195);
and U1405 (N_1405,N_225,N_339);
or U1406 (N_1406,N_921,N_441);
xnor U1407 (N_1407,N_549,N_671);
or U1408 (N_1408,N_81,N_318);
nand U1409 (N_1409,N_302,N_300);
or U1410 (N_1410,N_560,N_223);
or U1411 (N_1411,N_416,N_870);
or U1412 (N_1412,N_31,N_381);
and U1413 (N_1413,N_836,N_868);
nor U1414 (N_1414,N_100,N_92);
nand U1415 (N_1415,N_468,N_303);
nor U1416 (N_1416,N_893,N_782);
nand U1417 (N_1417,N_375,N_631);
and U1418 (N_1418,N_410,N_933);
and U1419 (N_1419,N_476,N_313);
nor U1420 (N_1420,N_451,N_938);
and U1421 (N_1421,N_439,N_553);
or U1422 (N_1422,N_385,N_523);
or U1423 (N_1423,N_114,N_308);
or U1424 (N_1424,N_140,N_797);
nand U1425 (N_1425,N_566,N_861);
nor U1426 (N_1426,N_525,N_498);
or U1427 (N_1427,N_736,N_478);
nor U1428 (N_1428,N_184,N_473);
and U1429 (N_1429,N_196,N_649);
and U1430 (N_1430,N_259,N_424);
or U1431 (N_1431,N_70,N_346);
nand U1432 (N_1432,N_564,N_472);
or U1433 (N_1433,N_991,N_426);
or U1434 (N_1434,N_155,N_487);
or U1435 (N_1435,N_816,N_150);
or U1436 (N_1436,N_420,N_260);
and U1437 (N_1437,N_469,N_710);
or U1438 (N_1438,N_951,N_204);
nor U1439 (N_1439,N_42,N_102);
nor U1440 (N_1440,N_686,N_628);
and U1441 (N_1441,N_534,N_605);
and U1442 (N_1442,N_759,N_697);
or U1443 (N_1443,N_10,N_106);
nand U1444 (N_1444,N_768,N_877);
and U1445 (N_1445,N_243,N_27);
nor U1446 (N_1446,N_363,N_201);
or U1447 (N_1447,N_454,N_767);
or U1448 (N_1448,N_521,N_644);
nor U1449 (N_1449,N_365,N_178);
nand U1450 (N_1450,N_875,N_288);
and U1451 (N_1451,N_772,N_461);
nand U1452 (N_1452,N_706,N_735);
nor U1453 (N_1453,N_146,N_661);
or U1454 (N_1454,N_616,N_349);
and U1455 (N_1455,N_509,N_926);
or U1456 (N_1456,N_233,N_95);
nand U1457 (N_1457,N_679,N_485);
nand U1458 (N_1458,N_11,N_805);
or U1459 (N_1459,N_377,N_82);
nor U1460 (N_1460,N_18,N_397);
or U1461 (N_1461,N_232,N_437);
nor U1462 (N_1462,N_869,N_462);
nor U1463 (N_1463,N_244,N_334);
nand U1464 (N_1464,N_582,N_297);
nand U1465 (N_1465,N_792,N_327);
or U1466 (N_1466,N_218,N_79);
or U1467 (N_1467,N_700,N_929);
or U1468 (N_1468,N_899,N_224);
nor U1469 (N_1469,N_443,N_946);
and U1470 (N_1470,N_190,N_16);
nand U1471 (N_1471,N_301,N_583);
nor U1472 (N_1472,N_387,N_267);
or U1473 (N_1473,N_892,N_347);
and U1474 (N_1474,N_242,N_927);
or U1475 (N_1475,N_770,N_33);
nand U1476 (N_1476,N_158,N_122);
and U1477 (N_1477,N_647,N_662);
nor U1478 (N_1478,N_29,N_925);
nand U1479 (N_1479,N_344,N_788);
nand U1480 (N_1480,N_635,N_378);
nand U1481 (N_1481,N_430,N_798);
or U1482 (N_1482,N_450,N_361);
nor U1483 (N_1483,N_357,N_678);
or U1484 (N_1484,N_494,N_618);
nor U1485 (N_1485,N_418,N_694);
or U1486 (N_1486,N_240,N_467);
nand U1487 (N_1487,N_688,N_890);
or U1488 (N_1488,N_707,N_460);
and U1489 (N_1489,N_531,N_171);
nand U1490 (N_1490,N_354,N_747);
and U1491 (N_1491,N_829,N_602);
nand U1492 (N_1492,N_474,N_379);
nor U1493 (N_1493,N_817,N_126);
nand U1494 (N_1494,N_518,N_637);
and U1495 (N_1495,N_414,N_413);
and U1496 (N_1496,N_273,N_607);
and U1497 (N_1497,N_495,N_83);
and U1498 (N_1498,N_638,N_58);
or U1499 (N_1499,N_513,N_5);
nor U1500 (N_1500,N_720,N_594);
and U1501 (N_1501,N_645,N_319);
or U1502 (N_1502,N_429,N_856);
and U1503 (N_1503,N_735,N_896);
or U1504 (N_1504,N_482,N_77);
and U1505 (N_1505,N_662,N_239);
nor U1506 (N_1506,N_727,N_380);
or U1507 (N_1507,N_35,N_438);
nand U1508 (N_1508,N_889,N_674);
and U1509 (N_1509,N_774,N_111);
nor U1510 (N_1510,N_175,N_209);
or U1511 (N_1511,N_890,N_581);
and U1512 (N_1512,N_717,N_204);
nor U1513 (N_1513,N_735,N_28);
nand U1514 (N_1514,N_960,N_799);
and U1515 (N_1515,N_996,N_690);
nor U1516 (N_1516,N_93,N_90);
nor U1517 (N_1517,N_919,N_816);
nor U1518 (N_1518,N_808,N_931);
nor U1519 (N_1519,N_627,N_967);
or U1520 (N_1520,N_569,N_689);
nor U1521 (N_1521,N_204,N_872);
and U1522 (N_1522,N_328,N_207);
or U1523 (N_1523,N_520,N_621);
or U1524 (N_1524,N_979,N_98);
nor U1525 (N_1525,N_772,N_392);
nand U1526 (N_1526,N_488,N_811);
and U1527 (N_1527,N_631,N_11);
nor U1528 (N_1528,N_964,N_157);
nor U1529 (N_1529,N_445,N_900);
nand U1530 (N_1530,N_254,N_724);
nand U1531 (N_1531,N_261,N_186);
and U1532 (N_1532,N_685,N_408);
or U1533 (N_1533,N_697,N_251);
or U1534 (N_1534,N_390,N_424);
nand U1535 (N_1535,N_713,N_272);
nor U1536 (N_1536,N_12,N_454);
and U1537 (N_1537,N_651,N_531);
or U1538 (N_1538,N_413,N_647);
and U1539 (N_1539,N_66,N_454);
and U1540 (N_1540,N_313,N_252);
nand U1541 (N_1541,N_478,N_514);
and U1542 (N_1542,N_92,N_728);
and U1543 (N_1543,N_776,N_451);
or U1544 (N_1544,N_993,N_885);
xor U1545 (N_1545,N_935,N_141);
and U1546 (N_1546,N_467,N_971);
nor U1547 (N_1547,N_617,N_975);
and U1548 (N_1548,N_167,N_599);
or U1549 (N_1549,N_692,N_739);
and U1550 (N_1550,N_349,N_312);
and U1551 (N_1551,N_923,N_30);
nand U1552 (N_1552,N_729,N_239);
or U1553 (N_1553,N_465,N_164);
nor U1554 (N_1554,N_315,N_832);
nand U1555 (N_1555,N_778,N_880);
and U1556 (N_1556,N_367,N_441);
nor U1557 (N_1557,N_455,N_807);
or U1558 (N_1558,N_360,N_114);
nand U1559 (N_1559,N_960,N_267);
nor U1560 (N_1560,N_564,N_307);
or U1561 (N_1561,N_369,N_639);
or U1562 (N_1562,N_212,N_694);
nand U1563 (N_1563,N_672,N_682);
nor U1564 (N_1564,N_876,N_569);
nor U1565 (N_1565,N_980,N_528);
nand U1566 (N_1566,N_718,N_327);
and U1567 (N_1567,N_536,N_102);
nor U1568 (N_1568,N_692,N_481);
or U1569 (N_1569,N_574,N_327);
nor U1570 (N_1570,N_593,N_677);
and U1571 (N_1571,N_501,N_290);
or U1572 (N_1572,N_836,N_550);
and U1573 (N_1573,N_625,N_917);
nand U1574 (N_1574,N_961,N_144);
nand U1575 (N_1575,N_850,N_458);
nand U1576 (N_1576,N_745,N_675);
and U1577 (N_1577,N_850,N_46);
nor U1578 (N_1578,N_904,N_694);
nor U1579 (N_1579,N_845,N_894);
nor U1580 (N_1580,N_968,N_7);
and U1581 (N_1581,N_271,N_143);
and U1582 (N_1582,N_72,N_474);
nand U1583 (N_1583,N_538,N_509);
or U1584 (N_1584,N_162,N_58);
nor U1585 (N_1585,N_594,N_77);
or U1586 (N_1586,N_60,N_312);
nand U1587 (N_1587,N_726,N_898);
or U1588 (N_1588,N_183,N_541);
nand U1589 (N_1589,N_584,N_688);
or U1590 (N_1590,N_582,N_708);
nor U1591 (N_1591,N_605,N_443);
or U1592 (N_1592,N_522,N_369);
nand U1593 (N_1593,N_542,N_111);
or U1594 (N_1594,N_537,N_749);
nand U1595 (N_1595,N_440,N_77);
and U1596 (N_1596,N_550,N_534);
nor U1597 (N_1597,N_811,N_332);
nand U1598 (N_1598,N_204,N_353);
nand U1599 (N_1599,N_43,N_945);
and U1600 (N_1600,N_210,N_337);
nor U1601 (N_1601,N_399,N_518);
nand U1602 (N_1602,N_818,N_136);
nor U1603 (N_1603,N_580,N_254);
and U1604 (N_1604,N_178,N_44);
nand U1605 (N_1605,N_855,N_443);
or U1606 (N_1606,N_257,N_119);
nor U1607 (N_1607,N_569,N_152);
and U1608 (N_1608,N_898,N_408);
or U1609 (N_1609,N_242,N_667);
nor U1610 (N_1610,N_710,N_718);
nor U1611 (N_1611,N_929,N_12);
nor U1612 (N_1612,N_355,N_128);
nor U1613 (N_1613,N_366,N_246);
and U1614 (N_1614,N_845,N_196);
nand U1615 (N_1615,N_320,N_331);
nand U1616 (N_1616,N_608,N_951);
nor U1617 (N_1617,N_865,N_229);
or U1618 (N_1618,N_70,N_554);
or U1619 (N_1619,N_449,N_361);
or U1620 (N_1620,N_999,N_659);
and U1621 (N_1621,N_385,N_681);
nor U1622 (N_1622,N_962,N_344);
nor U1623 (N_1623,N_296,N_46);
nor U1624 (N_1624,N_401,N_172);
or U1625 (N_1625,N_29,N_674);
and U1626 (N_1626,N_166,N_608);
nand U1627 (N_1627,N_588,N_244);
nand U1628 (N_1628,N_715,N_656);
or U1629 (N_1629,N_446,N_35);
nor U1630 (N_1630,N_544,N_957);
and U1631 (N_1631,N_4,N_120);
or U1632 (N_1632,N_367,N_703);
nor U1633 (N_1633,N_310,N_35);
or U1634 (N_1634,N_231,N_450);
nand U1635 (N_1635,N_485,N_602);
nand U1636 (N_1636,N_511,N_563);
and U1637 (N_1637,N_229,N_658);
or U1638 (N_1638,N_805,N_661);
nand U1639 (N_1639,N_37,N_175);
nand U1640 (N_1640,N_152,N_834);
nor U1641 (N_1641,N_797,N_6);
nor U1642 (N_1642,N_106,N_335);
and U1643 (N_1643,N_588,N_572);
nor U1644 (N_1644,N_601,N_636);
nor U1645 (N_1645,N_99,N_237);
nor U1646 (N_1646,N_865,N_364);
nor U1647 (N_1647,N_808,N_49);
or U1648 (N_1648,N_531,N_1);
and U1649 (N_1649,N_409,N_318);
or U1650 (N_1650,N_893,N_367);
or U1651 (N_1651,N_164,N_307);
and U1652 (N_1652,N_435,N_138);
or U1653 (N_1653,N_17,N_22);
nor U1654 (N_1654,N_549,N_861);
or U1655 (N_1655,N_806,N_463);
and U1656 (N_1656,N_296,N_399);
and U1657 (N_1657,N_261,N_32);
nor U1658 (N_1658,N_391,N_426);
and U1659 (N_1659,N_973,N_435);
and U1660 (N_1660,N_813,N_936);
and U1661 (N_1661,N_315,N_779);
nor U1662 (N_1662,N_992,N_317);
nand U1663 (N_1663,N_816,N_232);
and U1664 (N_1664,N_306,N_936);
nor U1665 (N_1665,N_2,N_798);
nand U1666 (N_1666,N_728,N_777);
nand U1667 (N_1667,N_654,N_702);
nor U1668 (N_1668,N_626,N_117);
and U1669 (N_1669,N_357,N_346);
or U1670 (N_1670,N_496,N_651);
or U1671 (N_1671,N_235,N_564);
or U1672 (N_1672,N_735,N_562);
nor U1673 (N_1673,N_841,N_355);
or U1674 (N_1674,N_379,N_1);
or U1675 (N_1675,N_841,N_184);
and U1676 (N_1676,N_871,N_509);
or U1677 (N_1677,N_777,N_136);
or U1678 (N_1678,N_722,N_427);
and U1679 (N_1679,N_914,N_269);
nand U1680 (N_1680,N_265,N_357);
nor U1681 (N_1681,N_416,N_348);
and U1682 (N_1682,N_858,N_575);
nand U1683 (N_1683,N_386,N_400);
nor U1684 (N_1684,N_439,N_700);
or U1685 (N_1685,N_137,N_262);
nor U1686 (N_1686,N_309,N_646);
nor U1687 (N_1687,N_957,N_2);
nand U1688 (N_1688,N_381,N_342);
and U1689 (N_1689,N_767,N_127);
nand U1690 (N_1690,N_58,N_412);
nand U1691 (N_1691,N_163,N_210);
nor U1692 (N_1692,N_947,N_732);
nand U1693 (N_1693,N_583,N_964);
and U1694 (N_1694,N_127,N_248);
nor U1695 (N_1695,N_331,N_508);
and U1696 (N_1696,N_754,N_466);
nand U1697 (N_1697,N_988,N_147);
or U1698 (N_1698,N_392,N_618);
or U1699 (N_1699,N_995,N_533);
nand U1700 (N_1700,N_978,N_826);
nand U1701 (N_1701,N_117,N_374);
nand U1702 (N_1702,N_663,N_930);
nor U1703 (N_1703,N_665,N_681);
nand U1704 (N_1704,N_289,N_130);
or U1705 (N_1705,N_838,N_904);
or U1706 (N_1706,N_198,N_317);
xor U1707 (N_1707,N_427,N_433);
nand U1708 (N_1708,N_948,N_573);
or U1709 (N_1709,N_36,N_292);
and U1710 (N_1710,N_856,N_889);
or U1711 (N_1711,N_866,N_161);
nand U1712 (N_1712,N_39,N_800);
or U1713 (N_1713,N_532,N_92);
nor U1714 (N_1714,N_210,N_199);
nand U1715 (N_1715,N_396,N_350);
nand U1716 (N_1716,N_767,N_191);
or U1717 (N_1717,N_602,N_608);
nand U1718 (N_1718,N_90,N_162);
and U1719 (N_1719,N_574,N_504);
nor U1720 (N_1720,N_228,N_430);
nand U1721 (N_1721,N_845,N_901);
and U1722 (N_1722,N_76,N_373);
or U1723 (N_1723,N_573,N_637);
and U1724 (N_1724,N_313,N_702);
nand U1725 (N_1725,N_569,N_355);
or U1726 (N_1726,N_403,N_609);
nor U1727 (N_1727,N_259,N_552);
and U1728 (N_1728,N_446,N_93);
nor U1729 (N_1729,N_118,N_565);
and U1730 (N_1730,N_776,N_374);
and U1731 (N_1731,N_27,N_383);
or U1732 (N_1732,N_387,N_850);
nand U1733 (N_1733,N_452,N_35);
and U1734 (N_1734,N_150,N_88);
nor U1735 (N_1735,N_297,N_576);
nor U1736 (N_1736,N_960,N_82);
nor U1737 (N_1737,N_964,N_675);
nand U1738 (N_1738,N_734,N_343);
nor U1739 (N_1739,N_715,N_534);
nand U1740 (N_1740,N_926,N_280);
or U1741 (N_1741,N_784,N_448);
or U1742 (N_1742,N_104,N_925);
and U1743 (N_1743,N_799,N_212);
or U1744 (N_1744,N_561,N_254);
and U1745 (N_1745,N_350,N_553);
nand U1746 (N_1746,N_387,N_655);
nor U1747 (N_1747,N_539,N_155);
nor U1748 (N_1748,N_861,N_793);
or U1749 (N_1749,N_719,N_31);
nand U1750 (N_1750,N_943,N_938);
or U1751 (N_1751,N_250,N_652);
nand U1752 (N_1752,N_273,N_73);
and U1753 (N_1753,N_677,N_947);
nand U1754 (N_1754,N_402,N_641);
nand U1755 (N_1755,N_589,N_746);
nor U1756 (N_1756,N_4,N_490);
nor U1757 (N_1757,N_902,N_721);
nand U1758 (N_1758,N_486,N_790);
nand U1759 (N_1759,N_726,N_541);
or U1760 (N_1760,N_832,N_335);
nor U1761 (N_1761,N_864,N_682);
or U1762 (N_1762,N_318,N_481);
and U1763 (N_1763,N_463,N_372);
and U1764 (N_1764,N_607,N_124);
nand U1765 (N_1765,N_861,N_611);
nor U1766 (N_1766,N_319,N_698);
and U1767 (N_1767,N_716,N_396);
nor U1768 (N_1768,N_367,N_87);
nand U1769 (N_1769,N_445,N_816);
or U1770 (N_1770,N_258,N_974);
nand U1771 (N_1771,N_329,N_706);
and U1772 (N_1772,N_657,N_549);
or U1773 (N_1773,N_72,N_643);
nor U1774 (N_1774,N_309,N_540);
or U1775 (N_1775,N_719,N_391);
or U1776 (N_1776,N_656,N_706);
or U1777 (N_1777,N_209,N_793);
nor U1778 (N_1778,N_13,N_603);
xnor U1779 (N_1779,N_229,N_987);
nand U1780 (N_1780,N_620,N_57);
nor U1781 (N_1781,N_898,N_845);
nand U1782 (N_1782,N_5,N_941);
nor U1783 (N_1783,N_882,N_987);
nand U1784 (N_1784,N_133,N_940);
nand U1785 (N_1785,N_467,N_844);
nor U1786 (N_1786,N_782,N_302);
nor U1787 (N_1787,N_412,N_367);
nand U1788 (N_1788,N_208,N_461);
or U1789 (N_1789,N_720,N_411);
nand U1790 (N_1790,N_922,N_4);
and U1791 (N_1791,N_706,N_958);
and U1792 (N_1792,N_212,N_845);
and U1793 (N_1793,N_197,N_487);
or U1794 (N_1794,N_572,N_596);
nand U1795 (N_1795,N_71,N_700);
nand U1796 (N_1796,N_417,N_924);
and U1797 (N_1797,N_676,N_833);
or U1798 (N_1798,N_882,N_401);
and U1799 (N_1799,N_786,N_645);
or U1800 (N_1800,N_656,N_417);
xnor U1801 (N_1801,N_571,N_688);
nor U1802 (N_1802,N_985,N_643);
nand U1803 (N_1803,N_614,N_523);
nor U1804 (N_1804,N_654,N_607);
and U1805 (N_1805,N_642,N_201);
nand U1806 (N_1806,N_206,N_455);
or U1807 (N_1807,N_648,N_961);
nor U1808 (N_1808,N_17,N_910);
or U1809 (N_1809,N_484,N_720);
and U1810 (N_1810,N_213,N_986);
nand U1811 (N_1811,N_591,N_508);
nand U1812 (N_1812,N_536,N_476);
nand U1813 (N_1813,N_928,N_341);
nand U1814 (N_1814,N_808,N_308);
xor U1815 (N_1815,N_374,N_835);
and U1816 (N_1816,N_106,N_156);
nor U1817 (N_1817,N_620,N_289);
or U1818 (N_1818,N_785,N_248);
or U1819 (N_1819,N_703,N_417);
or U1820 (N_1820,N_53,N_943);
nor U1821 (N_1821,N_871,N_70);
nand U1822 (N_1822,N_250,N_682);
nor U1823 (N_1823,N_832,N_528);
nor U1824 (N_1824,N_420,N_6);
and U1825 (N_1825,N_883,N_105);
and U1826 (N_1826,N_188,N_1);
or U1827 (N_1827,N_890,N_423);
and U1828 (N_1828,N_309,N_771);
or U1829 (N_1829,N_727,N_493);
nand U1830 (N_1830,N_699,N_910);
nor U1831 (N_1831,N_866,N_181);
nor U1832 (N_1832,N_524,N_304);
or U1833 (N_1833,N_585,N_742);
nand U1834 (N_1834,N_922,N_576);
or U1835 (N_1835,N_54,N_249);
or U1836 (N_1836,N_876,N_495);
nor U1837 (N_1837,N_417,N_736);
nand U1838 (N_1838,N_475,N_11);
nand U1839 (N_1839,N_197,N_754);
or U1840 (N_1840,N_627,N_981);
nor U1841 (N_1841,N_820,N_163);
nor U1842 (N_1842,N_706,N_966);
and U1843 (N_1843,N_531,N_461);
and U1844 (N_1844,N_733,N_353);
nand U1845 (N_1845,N_20,N_362);
or U1846 (N_1846,N_712,N_624);
nand U1847 (N_1847,N_753,N_886);
or U1848 (N_1848,N_615,N_951);
or U1849 (N_1849,N_824,N_433);
or U1850 (N_1850,N_243,N_600);
nand U1851 (N_1851,N_158,N_690);
or U1852 (N_1852,N_54,N_77);
or U1853 (N_1853,N_275,N_525);
nand U1854 (N_1854,N_500,N_716);
and U1855 (N_1855,N_557,N_859);
and U1856 (N_1856,N_882,N_782);
and U1857 (N_1857,N_238,N_368);
and U1858 (N_1858,N_13,N_750);
and U1859 (N_1859,N_364,N_9);
and U1860 (N_1860,N_824,N_197);
nor U1861 (N_1861,N_7,N_367);
nor U1862 (N_1862,N_89,N_36);
and U1863 (N_1863,N_928,N_962);
or U1864 (N_1864,N_637,N_66);
nand U1865 (N_1865,N_651,N_934);
nor U1866 (N_1866,N_838,N_83);
nand U1867 (N_1867,N_58,N_750);
nor U1868 (N_1868,N_953,N_279);
and U1869 (N_1869,N_911,N_808);
nor U1870 (N_1870,N_277,N_638);
nand U1871 (N_1871,N_650,N_699);
and U1872 (N_1872,N_478,N_855);
or U1873 (N_1873,N_813,N_986);
and U1874 (N_1874,N_415,N_998);
and U1875 (N_1875,N_827,N_648);
and U1876 (N_1876,N_842,N_565);
and U1877 (N_1877,N_313,N_670);
nor U1878 (N_1878,N_500,N_866);
nand U1879 (N_1879,N_620,N_12);
and U1880 (N_1880,N_64,N_13);
nand U1881 (N_1881,N_397,N_202);
nand U1882 (N_1882,N_647,N_959);
or U1883 (N_1883,N_888,N_815);
nand U1884 (N_1884,N_82,N_328);
and U1885 (N_1885,N_847,N_923);
or U1886 (N_1886,N_313,N_992);
nand U1887 (N_1887,N_317,N_325);
nand U1888 (N_1888,N_350,N_688);
nand U1889 (N_1889,N_499,N_814);
nor U1890 (N_1890,N_348,N_454);
nor U1891 (N_1891,N_872,N_941);
nand U1892 (N_1892,N_487,N_43);
nor U1893 (N_1893,N_305,N_785);
or U1894 (N_1894,N_761,N_896);
nor U1895 (N_1895,N_980,N_24);
nand U1896 (N_1896,N_500,N_153);
and U1897 (N_1897,N_999,N_30);
and U1898 (N_1898,N_618,N_243);
or U1899 (N_1899,N_193,N_842);
or U1900 (N_1900,N_170,N_520);
and U1901 (N_1901,N_981,N_932);
or U1902 (N_1902,N_393,N_77);
nor U1903 (N_1903,N_679,N_8);
nand U1904 (N_1904,N_627,N_332);
nor U1905 (N_1905,N_245,N_449);
and U1906 (N_1906,N_652,N_788);
or U1907 (N_1907,N_213,N_706);
nor U1908 (N_1908,N_916,N_201);
nor U1909 (N_1909,N_59,N_564);
and U1910 (N_1910,N_904,N_216);
nor U1911 (N_1911,N_271,N_532);
nand U1912 (N_1912,N_640,N_91);
or U1913 (N_1913,N_837,N_680);
nor U1914 (N_1914,N_930,N_876);
or U1915 (N_1915,N_799,N_301);
nand U1916 (N_1916,N_311,N_834);
nor U1917 (N_1917,N_814,N_516);
nor U1918 (N_1918,N_901,N_969);
xnor U1919 (N_1919,N_355,N_164);
or U1920 (N_1920,N_645,N_340);
nor U1921 (N_1921,N_841,N_545);
or U1922 (N_1922,N_402,N_79);
or U1923 (N_1923,N_481,N_371);
nor U1924 (N_1924,N_548,N_331);
or U1925 (N_1925,N_358,N_412);
or U1926 (N_1926,N_728,N_280);
and U1927 (N_1927,N_899,N_572);
and U1928 (N_1928,N_881,N_405);
or U1929 (N_1929,N_316,N_544);
nand U1930 (N_1930,N_769,N_866);
and U1931 (N_1931,N_537,N_551);
or U1932 (N_1932,N_286,N_508);
or U1933 (N_1933,N_55,N_664);
nand U1934 (N_1934,N_299,N_359);
or U1935 (N_1935,N_890,N_75);
or U1936 (N_1936,N_589,N_741);
nor U1937 (N_1937,N_752,N_532);
nor U1938 (N_1938,N_935,N_332);
and U1939 (N_1939,N_777,N_869);
or U1940 (N_1940,N_891,N_666);
nand U1941 (N_1941,N_828,N_515);
nor U1942 (N_1942,N_811,N_930);
nand U1943 (N_1943,N_171,N_144);
nand U1944 (N_1944,N_399,N_860);
or U1945 (N_1945,N_334,N_396);
nor U1946 (N_1946,N_492,N_242);
or U1947 (N_1947,N_89,N_420);
nand U1948 (N_1948,N_660,N_729);
nor U1949 (N_1949,N_582,N_626);
nor U1950 (N_1950,N_811,N_274);
and U1951 (N_1951,N_65,N_233);
nor U1952 (N_1952,N_876,N_126);
nor U1953 (N_1953,N_309,N_660);
or U1954 (N_1954,N_7,N_4);
or U1955 (N_1955,N_692,N_986);
or U1956 (N_1956,N_421,N_475);
nand U1957 (N_1957,N_170,N_543);
and U1958 (N_1958,N_234,N_638);
nand U1959 (N_1959,N_959,N_301);
nand U1960 (N_1960,N_40,N_776);
nand U1961 (N_1961,N_425,N_691);
nand U1962 (N_1962,N_882,N_800);
and U1963 (N_1963,N_222,N_162);
nand U1964 (N_1964,N_188,N_392);
or U1965 (N_1965,N_609,N_109);
and U1966 (N_1966,N_142,N_772);
nand U1967 (N_1967,N_865,N_394);
nor U1968 (N_1968,N_478,N_725);
nor U1969 (N_1969,N_841,N_401);
xor U1970 (N_1970,N_661,N_458);
nor U1971 (N_1971,N_463,N_764);
and U1972 (N_1972,N_157,N_301);
and U1973 (N_1973,N_115,N_93);
xor U1974 (N_1974,N_18,N_41);
nor U1975 (N_1975,N_150,N_513);
nand U1976 (N_1976,N_303,N_391);
nor U1977 (N_1977,N_233,N_483);
nand U1978 (N_1978,N_855,N_556);
nand U1979 (N_1979,N_386,N_946);
nor U1980 (N_1980,N_234,N_351);
nor U1981 (N_1981,N_864,N_742);
nand U1982 (N_1982,N_745,N_895);
nand U1983 (N_1983,N_925,N_737);
nand U1984 (N_1984,N_323,N_425);
nor U1985 (N_1985,N_613,N_886);
nor U1986 (N_1986,N_581,N_732);
nor U1987 (N_1987,N_589,N_165);
or U1988 (N_1988,N_857,N_372);
nand U1989 (N_1989,N_123,N_588);
nor U1990 (N_1990,N_516,N_485);
or U1991 (N_1991,N_22,N_780);
and U1992 (N_1992,N_799,N_179);
or U1993 (N_1993,N_644,N_900);
and U1994 (N_1994,N_789,N_130);
or U1995 (N_1995,N_364,N_117);
nor U1996 (N_1996,N_394,N_429);
and U1997 (N_1997,N_718,N_431);
nand U1998 (N_1998,N_753,N_592);
and U1999 (N_1999,N_551,N_585);
and U2000 (N_2000,N_1212,N_1300);
nor U2001 (N_2001,N_1642,N_1098);
nor U2002 (N_2002,N_1352,N_1563);
xor U2003 (N_2003,N_1675,N_1518);
and U2004 (N_2004,N_1745,N_1885);
or U2005 (N_2005,N_1981,N_1325);
and U2006 (N_2006,N_1035,N_1827);
nor U2007 (N_2007,N_1186,N_1086);
or U2008 (N_2008,N_1151,N_1206);
and U2009 (N_2009,N_1811,N_1595);
nand U2010 (N_2010,N_1892,N_1621);
nor U2011 (N_2011,N_1271,N_1336);
and U2012 (N_2012,N_1247,N_1366);
and U2013 (N_2013,N_1862,N_1765);
nor U2014 (N_2014,N_1315,N_1729);
nor U2015 (N_2015,N_1492,N_1200);
or U2016 (N_2016,N_1115,N_1180);
or U2017 (N_2017,N_1719,N_1252);
and U2018 (N_2018,N_1871,N_1565);
or U2019 (N_2019,N_1910,N_1726);
and U2020 (N_2020,N_1161,N_1288);
or U2021 (N_2021,N_1639,N_1465);
nand U2022 (N_2022,N_1464,N_1144);
nor U2023 (N_2023,N_1607,N_1654);
and U2024 (N_2024,N_1808,N_1660);
and U2025 (N_2025,N_1686,N_1333);
nand U2026 (N_2026,N_1994,N_1506);
and U2027 (N_2027,N_1880,N_1969);
or U2028 (N_2028,N_1743,N_1911);
or U2029 (N_2029,N_1323,N_1680);
or U2030 (N_2030,N_1917,N_1961);
nand U2031 (N_2031,N_1401,N_1459);
or U2032 (N_2032,N_1079,N_1174);
nand U2033 (N_2033,N_1580,N_1353);
or U2034 (N_2034,N_1795,N_1407);
nor U2035 (N_2035,N_1444,N_1205);
or U2036 (N_2036,N_1915,N_1165);
nand U2037 (N_2037,N_1410,N_1504);
nor U2038 (N_2038,N_1062,N_1409);
nand U2039 (N_2039,N_1239,N_1731);
or U2040 (N_2040,N_1559,N_1583);
nor U2041 (N_2041,N_1154,N_1546);
and U2042 (N_2042,N_1462,N_1370);
and U2043 (N_2043,N_1319,N_1725);
and U2044 (N_2044,N_1002,N_1950);
and U2045 (N_2045,N_1782,N_1983);
nand U2046 (N_2046,N_1221,N_1520);
and U2047 (N_2047,N_1657,N_1088);
or U2048 (N_2048,N_1176,N_1490);
or U2049 (N_2049,N_1228,N_1476);
or U2050 (N_2050,N_1667,N_1960);
and U2051 (N_2051,N_1209,N_1996);
and U2052 (N_2052,N_1946,N_1799);
nor U2053 (N_2053,N_1641,N_1394);
or U2054 (N_2054,N_1722,N_1131);
nand U2055 (N_2055,N_1412,N_1800);
and U2056 (N_2056,N_1438,N_1978);
and U2057 (N_2057,N_1674,N_1349);
nand U2058 (N_2058,N_1185,N_1399);
and U2059 (N_2059,N_1501,N_1877);
or U2060 (N_2060,N_1099,N_1012);
and U2061 (N_2061,N_1344,N_1486);
and U2062 (N_2062,N_1691,N_1619);
nor U2063 (N_2063,N_1682,N_1967);
nand U2064 (N_2064,N_1096,N_1890);
or U2065 (N_2065,N_1295,N_1290);
or U2066 (N_2066,N_1466,N_1661);
or U2067 (N_2067,N_1244,N_1780);
or U2068 (N_2068,N_1702,N_1510);
nand U2069 (N_2069,N_1508,N_1326);
and U2070 (N_2070,N_1669,N_1838);
nor U2071 (N_2071,N_1630,N_1939);
and U2072 (N_2072,N_1664,N_1928);
or U2073 (N_2073,N_1106,N_1867);
nand U2074 (N_2074,N_1920,N_1427);
nor U2075 (N_2075,N_1907,N_1446);
or U2076 (N_2076,N_1544,N_1817);
or U2077 (N_2077,N_1431,N_1945);
or U2078 (N_2078,N_1478,N_1178);
or U2079 (N_2079,N_1070,N_1162);
or U2080 (N_2080,N_1710,N_1814);
nand U2081 (N_2081,N_1944,N_1269);
and U2082 (N_2082,N_1530,N_1602);
nor U2083 (N_2083,N_1119,N_1777);
or U2084 (N_2084,N_1449,N_1701);
nand U2085 (N_2085,N_1140,N_1219);
nand U2086 (N_2086,N_1111,N_1004);
nor U2087 (N_2087,N_1285,N_1570);
nor U2088 (N_2088,N_1084,N_1526);
or U2089 (N_2089,N_1949,N_1953);
nor U2090 (N_2090,N_1739,N_1328);
and U2091 (N_2091,N_1037,N_1029);
nand U2092 (N_2092,N_1965,N_1679);
nor U2093 (N_2093,N_1255,N_1554);
nor U2094 (N_2094,N_1977,N_1477);
nand U2095 (N_2095,N_1282,N_1748);
nand U2096 (N_2096,N_1324,N_1321);
nor U2097 (N_2097,N_1975,N_1600);
nor U2098 (N_2098,N_1638,N_1397);
or U2099 (N_2099,N_1395,N_1887);
nand U2100 (N_2100,N_1312,N_1117);
nor U2101 (N_2101,N_1505,N_1644);
or U2102 (N_2102,N_1258,N_1534);
or U2103 (N_2103,N_1145,N_1104);
nand U2104 (N_2104,N_1519,N_1207);
or U2105 (N_2105,N_1440,N_1441);
and U2106 (N_2106,N_1329,N_1061);
nor U2107 (N_2107,N_1481,N_1773);
and U2108 (N_2108,N_1385,N_1776);
and U2109 (N_2109,N_1980,N_1606);
and U2110 (N_2110,N_1687,N_1331);
and U2111 (N_2111,N_1539,N_1372);
or U2112 (N_2112,N_1021,N_1418);
nor U2113 (N_2113,N_1381,N_1046);
nor U2114 (N_2114,N_1371,N_1601);
nand U2115 (N_2115,N_1134,N_1812);
nor U2116 (N_2116,N_1191,N_1286);
nor U2117 (N_2117,N_1284,N_1845);
nor U2118 (N_2118,N_1217,N_1986);
nor U2119 (N_2119,N_1335,N_1868);
or U2120 (N_2120,N_1482,N_1059);
nor U2121 (N_2121,N_1298,N_1820);
nor U2122 (N_2122,N_1789,N_1495);
and U2123 (N_2123,N_1704,N_1802);
nor U2124 (N_2124,N_1358,N_1724);
nor U2125 (N_2125,N_1576,N_1112);
and U2126 (N_2126,N_1738,N_1493);
nor U2127 (N_2127,N_1413,N_1668);
nand U2128 (N_2128,N_1141,N_1224);
and U2129 (N_2129,N_1901,N_1652);
nand U2130 (N_2130,N_1875,N_1826);
or U2131 (N_2131,N_1226,N_1631);
nor U2132 (N_2132,N_1833,N_1008);
and U2133 (N_2133,N_1376,N_1433);
nand U2134 (N_2134,N_1806,N_1883);
nor U2135 (N_2135,N_1753,N_1163);
nand U2136 (N_2136,N_1850,N_1732);
and U2137 (N_2137,N_1955,N_1929);
nand U2138 (N_2138,N_1645,N_1699);
or U2139 (N_2139,N_1153,N_1435);
nand U2140 (N_2140,N_1750,N_1952);
nor U2141 (N_2141,N_1582,N_1190);
or U2142 (N_2142,N_1545,N_1010);
nand U2143 (N_2143,N_1605,N_1623);
or U2144 (N_2144,N_1968,N_1696);
nor U2145 (N_2145,N_1487,N_1166);
or U2146 (N_2146,N_1542,N_1707);
nand U2147 (N_2147,N_1865,N_1304);
nand U2148 (N_2148,N_1825,N_1374);
and U2149 (N_2149,N_1881,N_1836);
nor U2150 (N_2150,N_1128,N_1683);
and U2151 (N_2151,N_1237,N_1741);
or U2152 (N_2152,N_1053,N_1499);
and U2153 (N_2153,N_1429,N_1659);
nor U2154 (N_2154,N_1591,N_1618);
or U2155 (N_2155,N_1175,N_1201);
and U2156 (N_2156,N_1422,N_1756);
nor U2157 (N_2157,N_1309,N_1234);
or U2158 (N_2158,N_1168,N_1172);
nand U2159 (N_2159,N_1337,N_1124);
and U2160 (N_2160,N_1218,N_1019);
nand U2161 (N_2161,N_1467,N_1818);
and U2162 (N_2162,N_1633,N_1067);
and U2163 (N_2163,N_1041,N_1824);
nand U2164 (N_2164,N_1058,N_1251);
or U2165 (N_2165,N_1898,N_1405);
and U2166 (N_2166,N_1541,N_1527);
nor U2167 (N_2167,N_1024,N_1020);
and U2168 (N_2168,N_1786,N_1677);
nand U2169 (N_2169,N_1573,N_1844);
or U2170 (N_2170,N_1509,N_1231);
nor U2171 (N_2171,N_1609,N_1211);
or U2172 (N_2172,N_1297,N_1489);
nor U2173 (N_2173,N_1671,N_1853);
nor U2174 (N_2174,N_1246,N_1320);
and U2175 (N_2175,N_1210,N_1164);
or U2176 (N_2176,N_1060,N_1423);
nand U2177 (N_2177,N_1143,N_1022);
nand U2178 (N_2178,N_1751,N_1543);
and U2179 (N_2179,N_1148,N_1045);
or U2180 (N_2180,N_1610,N_1962);
and U2181 (N_2181,N_1943,N_1406);
nand U2182 (N_2182,N_1289,N_1972);
or U2183 (N_2183,N_1785,N_1215);
xnor U2184 (N_2184,N_1569,N_1832);
and U2185 (N_2185,N_1771,N_1620);
and U2186 (N_2186,N_1819,N_1941);
nor U2187 (N_2187,N_1936,N_1643);
and U2188 (N_2188,N_1866,N_1872);
nor U2189 (N_2189,N_1524,N_1085);
nor U2190 (N_2190,N_1564,N_1856);
and U2191 (N_2191,N_1142,N_1223);
and U2192 (N_2192,N_1229,N_1556);
or U2193 (N_2193,N_1450,N_1895);
or U2194 (N_2194,N_1759,N_1150);
nand U2195 (N_2195,N_1050,N_1193);
or U2196 (N_2196,N_1127,N_1281);
nor U2197 (N_2197,N_1547,N_1456);
nor U2198 (N_2198,N_1919,N_1241);
or U2199 (N_2199,N_1711,N_1733);
or U2200 (N_2200,N_1049,N_1500);
nand U2201 (N_2201,N_1039,N_1473);
and U2202 (N_2202,N_1959,N_1888);
or U2203 (N_2203,N_1721,N_1964);
nand U2204 (N_2204,N_1834,N_1781);
nor U2205 (N_2205,N_1970,N_1801);
xnor U2206 (N_2206,N_1133,N_1485);
nor U2207 (N_2207,N_1453,N_1730);
and U2208 (N_2208,N_1663,N_1637);
nand U2209 (N_2209,N_1689,N_1275);
and U2210 (N_2210,N_1742,N_1636);
or U2211 (N_2211,N_1574,N_1757);
nor U2212 (N_2212,N_1828,N_1359);
or U2213 (N_2213,N_1717,N_1187);
and U2214 (N_2214,N_1114,N_1973);
nor U2215 (N_2215,N_1109,N_1558);
or U2216 (N_2216,N_1925,N_1640);
and U2217 (N_2217,N_1684,N_1391);
nor U2218 (N_2218,N_1420,N_1314);
nor U2219 (N_2219,N_1400,N_1015);
nor U2220 (N_2220,N_1313,N_1425);
nor U2221 (N_2221,N_1647,N_1308);
or U2222 (N_2222,N_1517,N_1030);
and U2223 (N_2223,N_1723,N_1798);
nand U2224 (N_2224,N_1382,N_1108);
nor U2225 (N_2225,N_1238,N_1204);
and U2226 (N_2226,N_1402,N_1598);
nor U2227 (N_2227,N_1149,N_1129);
and U2228 (N_2228,N_1577,N_1656);
and U2229 (N_2229,N_1028,N_1531);
nor U2230 (N_2230,N_1854,N_1227);
or U2231 (N_2231,N_1005,N_1192);
nand U2232 (N_2232,N_1779,N_1997);
nor U2233 (N_2233,N_1334,N_1013);
and U2234 (N_2234,N_1136,N_1208);
nor U2235 (N_2235,N_1551,N_1179);
nor U2236 (N_2236,N_1159,N_1305);
nand U2237 (N_2237,N_1171,N_1373);
or U2238 (N_2238,N_1572,N_1327);
or U2239 (N_2239,N_1987,N_1522);
and U2240 (N_2240,N_1727,N_1097);
and U2241 (N_2241,N_1317,N_1548);
and U2242 (N_2242,N_1183,N_1470);
and U2243 (N_2243,N_1199,N_1810);
nand U2244 (N_2244,N_1038,N_1762);
or U2245 (N_2245,N_1296,N_1507);
and U2246 (N_2246,N_1276,N_1170);
or U2247 (N_2247,N_1502,N_1649);
nor U2248 (N_2248,N_1581,N_1345);
and U2249 (N_2249,N_1474,N_1864);
or U2250 (N_2250,N_1389,N_1624);
nor U2251 (N_2251,N_1746,N_1403);
nor U2252 (N_2252,N_1794,N_1072);
and U2253 (N_2253,N_1078,N_1396);
nor U2254 (N_2254,N_1714,N_1700);
or U2255 (N_2255,N_1240,N_1471);
and U2256 (N_2256,N_1051,N_1788);
or U2257 (N_2257,N_1843,N_1626);
or U2258 (N_2258,N_1475,N_1803);
nor U2259 (N_2259,N_1956,N_1587);
nand U2260 (N_2260,N_1672,N_1347);
or U2261 (N_2261,N_1705,N_1066);
or U2262 (N_2262,N_1658,N_1796);
nand U2263 (N_2263,N_1135,N_1194);
nand U2264 (N_2264,N_1787,N_1216);
nor U2265 (N_2265,N_1918,N_1057);
or U2266 (N_2266,N_1695,N_1082);
and U2267 (N_2267,N_1628,N_1468);
and U2268 (N_2268,N_1622,N_1937);
and U2269 (N_2269,N_1951,N_1536);
nor U2270 (N_2270,N_1392,N_1043);
nand U2271 (N_2271,N_1612,N_1365);
or U2272 (N_2272,N_1860,N_1560);
nand U2273 (N_2273,N_1356,N_1934);
nor U2274 (N_2274,N_1708,N_1483);
or U2275 (N_2275,N_1455,N_1555);
and U2276 (N_2276,N_1461,N_1829);
or U2277 (N_2277,N_1198,N_1398);
nand U2278 (N_2278,N_1350,N_1966);
or U2279 (N_2279,N_1380,N_1805);
nor U2280 (N_2280,N_1414,N_1254);
or U2281 (N_2281,N_1823,N_1177);
and U2282 (N_2282,N_1584,N_1566);
xnor U2283 (N_2283,N_1528,N_1138);
or U2284 (N_2284,N_1930,N_1614);
and U2285 (N_2285,N_1635,N_1342);
or U2286 (N_2286,N_1755,N_1681);
nand U2287 (N_2287,N_1203,N_1256);
nor U2288 (N_2288,N_1747,N_1767);
or U2289 (N_2289,N_1993,N_1763);
and U2290 (N_2290,N_1393,N_1589);
or U2291 (N_2291,N_1585,N_1855);
and U2292 (N_2292,N_1263,N_1575);
or U2293 (N_2293,N_1387,N_1749);
or U2294 (N_2294,N_1744,N_1849);
nand U2295 (N_2295,N_1089,N_1454);
nand U2296 (N_2296,N_1311,N_1879);
and U2297 (N_2297,N_1503,N_1047);
nor U2298 (N_2298,N_1242,N_1369);
nand U2299 (N_2299,N_1213,N_1457);
nor U2300 (N_2300,N_1235,N_1257);
and U2301 (N_2301,N_1125,N_1302);
or U2302 (N_2302,N_1291,N_1430);
and U2303 (N_2303,N_1835,N_1693);
nand U2304 (N_2304,N_1513,N_1137);
nand U2305 (N_2305,N_1330,N_1735);
nand U2306 (N_2306,N_1995,N_1837);
or U2307 (N_2307,N_1891,N_1615);
and U2308 (N_2308,N_1469,N_1913);
nand U2309 (N_2309,N_1388,N_1783);
or U2310 (N_2310,N_1354,N_1886);
nand U2311 (N_2311,N_1442,N_1230);
and U2312 (N_2312,N_1417,N_1073);
and U2313 (N_2313,N_1740,N_1222);
nand U2314 (N_2314,N_1197,N_1123);
nor U2315 (N_2315,N_1157,N_1809);
nor U2316 (N_2316,N_1511,N_1090);
nor U2317 (N_2317,N_1797,N_1361);
nand U2318 (N_2318,N_1270,N_1122);
and U2319 (N_2319,N_1232,N_1404);
nand U2320 (N_2320,N_1593,N_1355);
or U2321 (N_2321,N_1195,N_1971);
and U2322 (N_2322,N_1611,N_1260);
or U2323 (N_2323,N_1550,N_1032);
nor U2324 (N_2324,N_1902,N_1225);
nand U2325 (N_2325,N_1307,N_1292);
and U2326 (N_2326,N_1998,N_1958);
nor U2327 (N_2327,N_1274,N_1516);
or U2328 (N_2328,N_1367,N_1065);
nor U2329 (N_2329,N_1279,N_1259);
nand U2330 (N_2330,N_1521,N_1093);
nand U2331 (N_2331,N_1384,N_1126);
nand U2332 (N_2332,N_1497,N_1364);
nor U2333 (N_2333,N_1293,N_1588);
and U2334 (N_2334,N_1734,N_1863);
or U2335 (N_2335,N_1596,N_1512);
nor U2336 (N_2336,N_1648,N_1332);
and U2337 (N_2337,N_1006,N_1909);
and U2338 (N_2338,N_1031,N_1666);
nand U2339 (N_2339,N_1018,N_1793);
nor U2340 (N_2340,N_1113,N_1306);
or U2341 (N_2341,N_1139,N_1214);
nor U2342 (N_2342,N_1592,N_1650);
nor U2343 (N_2343,N_1419,N_1884);
nor U2344 (N_2344,N_1390,N_1338);
nor U2345 (N_2345,N_1979,N_1923);
nor U2346 (N_2346,N_1807,N_1264);
nor U2347 (N_2347,N_1718,N_1760);
nand U2348 (N_2348,N_1940,N_1561);
nor U2349 (N_2349,N_1452,N_1976);
nor U2350 (N_2350,N_1432,N_1525);
or U2351 (N_2351,N_1017,N_1822);
nor U2352 (N_2352,N_1688,N_1957);
or U2353 (N_2353,N_1245,N_1272);
or U2354 (N_2354,N_1676,N_1932);
nand U2355 (N_2355,N_1054,N_1784);
nor U2356 (N_2356,N_1152,N_1105);
nand U2357 (N_2357,N_1590,N_1906);
or U2358 (N_2358,N_1772,N_1250);
nand U2359 (N_2359,N_1988,N_1287);
nor U2360 (N_2360,N_1662,N_1651);
nand U2361 (N_2361,N_1273,N_1278);
nand U2362 (N_2362,N_1001,N_1922);
and U2363 (N_2363,N_1102,N_1715);
nor U2364 (N_2364,N_1146,N_1301);
nor U2365 (N_2365,N_1056,N_1599);
or U2366 (N_2366,N_1839,N_1277);
or U2367 (N_2367,N_1603,N_1014);
nand U2368 (N_2368,N_1678,N_1552);
or U2369 (N_2369,N_1617,N_1848);
nand U2370 (N_2370,N_1874,N_1873);
or U2371 (N_2371,N_1351,N_1488);
nor U2372 (N_2372,N_1713,N_1737);
nor U2373 (N_2373,N_1169,N_1770);
nand U2374 (N_2374,N_1173,N_1608);
or U2375 (N_2375,N_1882,N_1383);
nand U2376 (N_2376,N_1445,N_1578);
or U2377 (N_2377,N_1692,N_1665);
nand U2378 (N_2378,N_1484,N_1386);
nor U2379 (N_2379,N_1160,N_1120);
nor U2380 (N_2380,N_1766,N_1447);
nor U2381 (N_2381,N_1158,N_1876);
nand U2382 (N_2382,N_1894,N_1984);
nor U2383 (N_2383,N_1156,N_1627);
and U2384 (N_2384,N_1632,N_1299);
nor U2385 (N_2385,N_1071,N_1904);
nor U2386 (N_2386,N_1931,N_1092);
nor U2387 (N_2387,N_1537,N_1316);
nor U2388 (N_2388,N_1343,N_1992);
nand U2389 (N_2389,N_1948,N_1424);
nand U2390 (N_2390,N_1804,N_1553);
nand U2391 (N_2391,N_1963,N_1322);
nand U2392 (N_2392,N_1974,N_1908);
or U2393 (N_2393,N_1861,N_1899);
or U2394 (N_2394,N_1016,N_1790);
nand U2395 (N_2395,N_1460,N_1549);
or U2396 (N_2396,N_1858,N_1847);
and U2397 (N_2397,N_1100,N_1670);
and U2398 (N_2398,N_1025,N_1942);
nand U2399 (N_2399,N_1080,N_1815);
or U2400 (N_2400,N_1878,N_1924);
nand U2401 (N_2401,N_1491,N_1905);
nor U2402 (N_2402,N_1896,N_1761);
or U2403 (N_2403,N_1991,N_1816);
nand U2404 (N_2404,N_1118,N_1167);
nand U2405 (N_2405,N_1036,N_1181);
nand U2406 (N_2406,N_1052,N_1912);
nand U2407 (N_2407,N_1716,N_1754);
and U2408 (N_2408,N_1044,N_1033);
nor U2409 (N_2409,N_1375,N_1339);
and U2410 (N_2410,N_1261,N_1515);
or U2411 (N_2411,N_1533,N_1698);
or U2412 (N_2412,N_1220,N_1437);
nor U2413 (N_2413,N_1266,N_1523);
or U2414 (N_2414,N_1758,N_1443);
and U2415 (N_2415,N_1498,N_1893);
and U2416 (N_2416,N_1532,N_1709);
and U2417 (N_2417,N_1377,N_1378);
nand U2418 (N_2418,N_1416,N_1557);
nor U2419 (N_2419,N_1625,N_1357);
nand U2420 (N_2420,N_1346,N_1116);
and U2421 (N_2421,N_1653,N_1752);
or U2422 (N_2422,N_1706,N_1236);
and U2423 (N_2423,N_1567,N_1363);
xnor U2424 (N_2424,N_1095,N_1496);
and U2425 (N_2425,N_1294,N_1009);
nand U2426 (N_2426,N_1027,N_1703);
or U2427 (N_2427,N_1935,N_1472);
xnor U2428 (N_2428,N_1985,N_1673);
or U2429 (N_2429,N_1267,N_1571);
nand U2430 (N_2430,N_1933,N_1914);
and U2431 (N_2431,N_1411,N_1026);
or U2432 (N_2432,N_1697,N_1846);
nor U2433 (N_2433,N_1458,N_1068);
or U2434 (N_2434,N_1479,N_1921);
nand U2435 (N_2435,N_1248,N_1712);
and U2436 (N_2436,N_1830,N_1064);
or U2437 (N_2437,N_1529,N_1132);
and U2438 (N_2438,N_1870,N_1101);
nor U2439 (N_2439,N_1243,N_1434);
and U2440 (N_2440,N_1728,N_1857);
and U2441 (N_2441,N_1428,N_1094);
or U2442 (N_2442,N_1426,N_1616);
nand U2443 (N_2443,N_1063,N_1121);
nand U2444 (N_2444,N_1463,N_1077);
or U2445 (N_2445,N_1629,N_1990);
nor U2446 (N_2446,N_1023,N_1448);
or U2447 (N_2447,N_1075,N_1764);
or U2448 (N_2448,N_1360,N_1318);
or U2449 (N_2449,N_1869,N_1233);
nand U2450 (N_2450,N_1451,N_1034);
nand U2451 (N_2451,N_1646,N_1694);
and U2452 (N_2452,N_1999,N_1415);
and U2453 (N_2453,N_1091,N_1249);
nand U2454 (N_2454,N_1083,N_1989);
nor U2455 (N_2455,N_1947,N_1690);
or U2456 (N_2456,N_1436,N_1188);
or U2457 (N_2457,N_1011,N_1147);
or U2458 (N_2458,N_1774,N_1368);
and U2459 (N_2459,N_1842,N_1791);
nor U2460 (N_2460,N_1494,N_1655);
nand U2461 (N_2461,N_1927,N_1926);
nand U2462 (N_2462,N_1362,N_1087);
nor U2463 (N_2463,N_1604,N_1720);
nor U2464 (N_2464,N_1903,N_1076);
nand U2465 (N_2465,N_1778,N_1634);
nor U2466 (N_2466,N_1155,N_1048);
or U2467 (N_2467,N_1184,N_1340);
and U2468 (N_2468,N_1982,N_1007);
nor U2469 (N_2469,N_1586,N_1081);
or U2470 (N_2470,N_1074,N_1841);
and U2471 (N_2471,N_1736,N_1568);
or U2472 (N_2472,N_1685,N_1813);
and U2473 (N_2473,N_1262,N_1594);
or U2474 (N_2474,N_1310,N_1859);
and U2475 (N_2475,N_1253,N_1268);
nand U2476 (N_2476,N_1852,N_1938);
or U2477 (N_2477,N_1202,N_1768);
and U2478 (N_2478,N_1535,N_1514);
and U2479 (N_2479,N_1954,N_1069);
nor U2480 (N_2480,N_1775,N_1110);
and U2481 (N_2481,N_1055,N_1831);
nand U2482 (N_2482,N_1130,N_1821);
nand U2483 (N_2483,N_1897,N_1562);
nor U2484 (N_2484,N_1040,N_1042);
or U2485 (N_2485,N_1900,N_1916);
nor U2486 (N_2486,N_1597,N_1439);
nand U2487 (N_2487,N_1189,N_1283);
nor U2488 (N_2488,N_1421,N_1379);
or U2489 (N_2489,N_1341,N_1613);
and U2490 (N_2490,N_1280,N_1792);
or U2491 (N_2491,N_1107,N_1348);
or U2492 (N_2492,N_1265,N_1538);
and U2493 (N_2493,N_1540,N_1889);
nand U2494 (N_2494,N_1103,N_1182);
or U2495 (N_2495,N_1840,N_1196);
nor U2496 (N_2496,N_1408,N_1000);
and U2497 (N_2497,N_1769,N_1579);
and U2498 (N_2498,N_1480,N_1851);
nor U2499 (N_2499,N_1003,N_1303);
and U2500 (N_2500,N_1454,N_1951);
or U2501 (N_2501,N_1331,N_1789);
and U2502 (N_2502,N_1214,N_1949);
or U2503 (N_2503,N_1931,N_1107);
or U2504 (N_2504,N_1765,N_1289);
nand U2505 (N_2505,N_1676,N_1315);
or U2506 (N_2506,N_1125,N_1317);
and U2507 (N_2507,N_1523,N_1157);
nand U2508 (N_2508,N_1057,N_1002);
and U2509 (N_2509,N_1083,N_1723);
and U2510 (N_2510,N_1144,N_1958);
and U2511 (N_2511,N_1437,N_1164);
or U2512 (N_2512,N_1697,N_1605);
or U2513 (N_2513,N_1733,N_1597);
or U2514 (N_2514,N_1273,N_1566);
and U2515 (N_2515,N_1942,N_1961);
nand U2516 (N_2516,N_1784,N_1662);
nor U2517 (N_2517,N_1039,N_1751);
and U2518 (N_2518,N_1996,N_1853);
nor U2519 (N_2519,N_1807,N_1559);
nand U2520 (N_2520,N_1725,N_1833);
and U2521 (N_2521,N_1997,N_1105);
and U2522 (N_2522,N_1722,N_1351);
nor U2523 (N_2523,N_1427,N_1357);
nand U2524 (N_2524,N_1174,N_1002);
and U2525 (N_2525,N_1806,N_1175);
and U2526 (N_2526,N_1573,N_1859);
nand U2527 (N_2527,N_1970,N_1836);
and U2528 (N_2528,N_1500,N_1493);
nand U2529 (N_2529,N_1007,N_1200);
and U2530 (N_2530,N_1127,N_1571);
and U2531 (N_2531,N_1953,N_1140);
nand U2532 (N_2532,N_1049,N_1565);
nand U2533 (N_2533,N_1582,N_1102);
and U2534 (N_2534,N_1684,N_1926);
nor U2535 (N_2535,N_1254,N_1205);
nor U2536 (N_2536,N_1941,N_1360);
or U2537 (N_2537,N_1811,N_1433);
or U2538 (N_2538,N_1518,N_1230);
nand U2539 (N_2539,N_1472,N_1090);
or U2540 (N_2540,N_1955,N_1010);
nor U2541 (N_2541,N_1192,N_1449);
and U2542 (N_2542,N_1239,N_1401);
nand U2543 (N_2543,N_1573,N_1222);
or U2544 (N_2544,N_1100,N_1902);
or U2545 (N_2545,N_1303,N_1700);
or U2546 (N_2546,N_1295,N_1151);
or U2547 (N_2547,N_1567,N_1351);
and U2548 (N_2548,N_1684,N_1970);
nor U2549 (N_2549,N_1499,N_1959);
or U2550 (N_2550,N_1851,N_1225);
and U2551 (N_2551,N_1541,N_1866);
or U2552 (N_2552,N_1904,N_1892);
nor U2553 (N_2553,N_1187,N_1353);
or U2554 (N_2554,N_1475,N_1480);
and U2555 (N_2555,N_1799,N_1954);
nand U2556 (N_2556,N_1188,N_1279);
or U2557 (N_2557,N_1039,N_1712);
or U2558 (N_2558,N_1432,N_1270);
nor U2559 (N_2559,N_1747,N_1425);
or U2560 (N_2560,N_1632,N_1845);
and U2561 (N_2561,N_1860,N_1225);
nand U2562 (N_2562,N_1960,N_1599);
nand U2563 (N_2563,N_1933,N_1343);
nand U2564 (N_2564,N_1210,N_1851);
nor U2565 (N_2565,N_1052,N_1920);
and U2566 (N_2566,N_1399,N_1986);
nand U2567 (N_2567,N_1098,N_1583);
nor U2568 (N_2568,N_1352,N_1443);
and U2569 (N_2569,N_1377,N_1741);
or U2570 (N_2570,N_1206,N_1186);
or U2571 (N_2571,N_1982,N_1871);
nand U2572 (N_2572,N_1334,N_1060);
or U2573 (N_2573,N_1515,N_1616);
or U2574 (N_2574,N_1048,N_1353);
or U2575 (N_2575,N_1624,N_1429);
and U2576 (N_2576,N_1872,N_1247);
nor U2577 (N_2577,N_1523,N_1120);
nor U2578 (N_2578,N_1766,N_1520);
or U2579 (N_2579,N_1207,N_1186);
and U2580 (N_2580,N_1638,N_1838);
or U2581 (N_2581,N_1611,N_1381);
and U2582 (N_2582,N_1851,N_1565);
and U2583 (N_2583,N_1707,N_1748);
nand U2584 (N_2584,N_1358,N_1792);
nor U2585 (N_2585,N_1103,N_1466);
xor U2586 (N_2586,N_1104,N_1456);
and U2587 (N_2587,N_1011,N_1332);
nand U2588 (N_2588,N_1863,N_1393);
nor U2589 (N_2589,N_1134,N_1161);
or U2590 (N_2590,N_1617,N_1371);
or U2591 (N_2591,N_1093,N_1918);
nand U2592 (N_2592,N_1913,N_1455);
and U2593 (N_2593,N_1831,N_1616);
nand U2594 (N_2594,N_1340,N_1485);
and U2595 (N_2595,N_1047,N_1838);
nand U2596 (N_2596,N_1918,N_1271);
nand U2597 (N_2597,N_1936,N_1818);
nand U2598 (N_2598,N_1954,N_1152);
nand U2599 (N_2599,N_1908,N_1832);
nor U2600 (N_2600,N_1523,N_1745);
nor U2601 (N_2601,N_1822,N_1308);
and U2602 (N_2602,N_1223,N_1946);
and U2603 (N_2603,N_1545,N_1648);
nor U2604 (N_2604,N_1298,N_1853);
and U2605 (N_2605,N_1081,N_1519);
or U2606 (N_2606,N_1596,N_1786);
nor U2607 (N_2607,N_1563,N_1675);
nor U2608 (N_2608,N_1640,N_1556);
nor U2609 (N_2609,N_1909,N_1188);
nand U2610 (N_2610,N_1662,N_1513);
nand U2611 (N_2611,N_1249,N_1481);
nand U2612 (N_2612,N_1921,N_1395);
and U2613 (N_2613,N_1820,N_1774);
nand U2614 (N_2614,N_1034,N_1525);
nor U2615 (N_2615,N_1234,N_1022);
nand U2616 (N_2616,N_1074,N_1717);
or U2617 (N_2617,N_1798,N_1138);
and U2618 (N_2618,N_1254,N_1630);
and U2619 (N_2619,N_1478,N_1169);
nand U2620 (N_2620,N_1384,N_1832);
or U2621 (N_2621,N_1872,N_1898);
nand U2622 (N_2622,N_1590,N_1946);
nand U2623 (N_2623,N_1957,N_1034);
or U2624 (N_2624,N_1307,N_1062);
nor U2625 (N_2625,N_1829,N_1863);
and U2626 (N_2626,N_1696,N_1278);
and U2627 (N_2627,N_1707,N_1774);
nand U2628 (N_2628,N_1202,N_1681);
nand U2629 (N_2629,N_1484,N_1138);
nor U2630 (N_2630,N_1403,N_1076);
nand U2631 (N_2631,N_1784,N_1473);
or U2632 (N_2632,N_1426,N_1055);
and U2633 (N_2633,N_1950,N_1308);
and U2634 (N_2634,N_1197,N_1069);
or U2635 (N_2635,N_1906,N_1920);
nand U2636 (N_2636,N_1229,N_1522);
and U2637 (N_2637,N_1616,N_1765);
or U2638 (N_2638,N_1282,N_1380);
nand U2639 (N_2639,N_1564,N_1039);
nor U2640 (N_2640,N_1270,N_1326);
and U2641 (N_2641,N_1523,N_1919);
nand U2642 (N_2642,N_1647,N_1699);
nand U2643 (N_2643,N_1873,N_1363);
nor U2644 (N_2644,N_1894,N_1545);
nand U2645 (N_2645,N_1947,N_1595);
nor U2646 (N_2646,N_1147,N_1861);
nand U2647 (N_2647,N_1381,N_1943);
or U2648 (N_2648,N_1008,N_1212);
or U2649 (N_2649,N_1222,N_1293);
or U2650 (N_2650,N_1480,N_1387);
nor U2651 (N_2651,N_1590,N_1984);
or U2652 (N_2652,N_1712,N_1678);
nor U2653 (N_2653,N_1490,N_1479);
nor U2654 (N_2654,N_1214,N_1327);
nand U2655 (N_2655,N_1048,N_1415);
or U2656 (N_2656,N_1168,N_1010);
nand U2657 (N_2657,N_1504,N_1999);
and U2658 (N_2658,N_1761,N_1972);
nand U2659 (N_2659,N_1982,N_1584);
nor U2660 (N_2660,N_1262,N_1303);
or U2661 (N_2661,N_1956,N_1021);
or U2662 (N_2662,N_1582,N_1827);
or U2663 (N_2663,N_1696,N_1793);
or U2664 (N_2664,N_1295,N_1256);
nand U2665 (N_2665,N_1358,N_1802);
nor U2666 (N_2666,N_1871,N_1922);
nand U2667 (N_2667,N_1609,N_1914);
nor U2668 (N_2668,N_1110,N_1818);
nand U2669 (N_2669,N_1941,N_1844);
and U2670 (N_2670,N_1749,N_1707);
nor U2671 (N_2671,N_1180,N_1632);
and U2672 (N_2672,N_1302,N_1733);
and U2673 (N_2673,N_1629,N_1155);
and U2674 (N_2674,N_1549,N_1389);
nand U2675 (N_2675,N_1736,N_1041);
or U2676 (N_2676,N_1975,N_1034);
nor U2677 (N_2677,N_1310,N_1889);
nand U2678 (N_2678,N_1768,N_1327);
nand U2679 (N_2679,N_1753,N_1685);
nand U2680 (N_2680,N_1320,N_1704);
and U2681 (N_2681,N_1634,N_1739);
or U2682 (N_2682,N_1715,N_1165);
or U2683 (N_2683,N_1148,N_1186);
nor U2684 (N_2684,N_1934,N_1997);
and U2685 (N_2685,N_1229,N_1652);
or U2686 (N_2686,N_1933,N_1038);
or U2687 (N_2687,N_1046,N_1635);
nor U2688 (N_2688,N_1677,N_1293);
or U2689 (N_2689,N_1798,N_1477);
and U2690 (N_2690,N_1974,N_1811);
or U2691 (N_2691,N_1307,N_1193);
and U2692 (N_2692,N_1753,N_1514);
and U2693 (N_2693,N_1886,N_1674);
and U2694 (N_2694,N_1143,N_1581);
and U2695 (N_2695,N_1093,N_1302);
nor U2696 (N_2696,N_1078,N_1937);
and U2697 (N_2697,N_1698,N_1408);
nand U2698 (N_2698,N_1208,N_1128);
nand U2699 (N_2699,N_1864,N_1578);
nand U2700 (N_2700,N_1719,N_1724);
nand U2701 (N_2701,N_1806,N_1520);
or U2702 (N_2702,N_1109,N_1912);
and U2703 (N_2703,N_1915,N_1029);
or U2704 (N_2704,N_1830,N_1354);
nor U2705 (N_2705,N_1026,N_1792);
nor U2706 (N_2706,N_1078,N_1651);
nor U2707 (N_2707,N_1001,N_1453);
or U2708 (N_2708,N_1022,N_1432);
or U2709 (N_2709,N_1773,N_1918);
and U2710 (N_2710,N_1385,N_1943);
nor U2711 (N_2711,N_1666,N_1343);
nand U2712 (N_2712,N_1887,N_1127);
and U2713 (N_2713,N_1575,N_1626);
nor U2714 (N_2714,N_1299,N_1896);
nor U2715 (N_2715,N_1179,N_1870);
or U2716 (N_2716,N_1786,N_1784);
or U2717 (N_2717,N_1605,N_1309);
or U2718 (N_2718,N_1463,N_1167);
nor U2719 (N_2719,N_1984,N_1810);
or U2720 (N_2720,N_1897,N_1778);
or U2721 (N_2721,N_1105,N_1812);
or U2722 (N_2722,N_1609,N_1372);
nand U2723 (N_2723,N_1309,N_1659);
and U2724 (N_2724,N_1752,N_1987);
and U2725 (N_2725,N_1687,N_1424);
nor U2726 (N_2726,N_1223,N_1782);
or U2727 (N_2727,N_1711,N_1856);
or U2728 (N_2728,N_1693,N_1538);
or U2729 (N_2729,N_1932,N_1547);
nor U2730 (N_2730,N_1068,N_1588);
nand U2731 (N_2731,N_1503,N_1758);
or U2732 (N_2732,N_1117,N_1056);
or U2733 (N_2733,N_1774,N_1952);
nor U2734 (N_2734,N_1043,N_1506);
and U2735 (N_2735,N_1036,N_1109);
nand U2736 (N_2736,N_1081,N_1324);
nor U2737 (N_2737,N_1185,N_1443);
and U2738 (N_2738,N_1539,N_1012);
and U2739 (N_2739,N_1336,N_1833);
nand U2740 (N_2740,N_1292,N_1610);
and U2741 (N_2741,N_1906,N_1160);
or U2742 (N_2742,N_1216,N_1376);
or U2743 (N_2743,N_1123,N_1507);
nor U2744 (N_2744,N_1418,N_1063);
or U2745 (N_2745,N_1186,N_1407);
or U2746 (N_2746,N_1424,N_1816);
nor U2747 (N_2747,N_1494,N_1460);
and U2748 (N_2748,N_1278,N_1978);
nor U2749 (N_2749,N_1042,N_1737);
and U2750 (N_2750,N_1834,N_1646);
nor U2751 (N_2751,N_1901,N_1283);
nor U2752 (N_2752,N_1555,N_1939);
nor U2753 (N_2753,N_1131,N_1830);
and U2754 (N_2754,N_1397,N_1921);
or U2755 (N_2755,N_1701,N_1609);
and U2756 (N_2756,N_1005,N_1270);
nor U2757 (N_2757,N_1680,N_1787);
nor U2758 (N_2758,N_1737,N_1850);
nand U2759 (N_2759,N_1775,N_1025);
and U2760 (N_2760,N_1882,N_1518);
or U2761 (N_2761,N_1446,N_1431);
or U2762 (N_2762,N_1816,N_1090);
and U2763 (N_2763,N_1621,N_1384);
nand U2764 (N_2764,N_1724,N_1356);
and U2765 (N_2765,N_1387,N_1741);
or U2766 (N_2766,N_1049,N_1765);
nor U2767 (N_2767,N_1416,N_1434);
or U2768 (N_2768,N_1918,N_1835);
nor U2769 (N_2769,N_1560,N_1762);
nand U2770 (N_2770,N_1556,N_1548);
nor U2771 (N_2771,N_1558,N_1598);
and U2772 (N_2772,N_1053,N_1455);
nand U2773 (N_2773,N_1343,N_1746);
or U2774 (N_2774,N_1875,N_1155);
or U2775 (N_2775,N_1126,N_1514);
nand U2776 (N_2776,N_1748,N_1286);
nand U2777 (N_2777,N_1496,N_1837);
or U2778 (N_2778,N_1904,N_1918);
nor U2779 (N_2779,N_1175,N_1325);
or U2780 (N_2780,N_1260,N_1027);
nand U2781 (N_2781,N_1365,N_1692);
or U2782 (N_2782,N_1329,N_1334);
or U2783 (N_2783,N_1648,N_1830);
nand U2784 (N_2784,N_1763,N_1468);
nor U2785 (N_2785,N_1687,N_1722);
nand U2786 (N_2786,N_1142,N_1464);
and U2787 (N_2787,N_1772,N_1932);
or U2788 (N_2788,N_1101,N_1802);
nand U2789 (N_2789,N_1034,N_1838);
nand U2790 (N_2790,N_1326,N_1317);
nand U2791 (N_2791,N_1203,N_1744);
or U2792 (N_2792,N_1543,N_1169);
nand U2793 (N_2793,N_1179,N_1571);
and U2794 (N_2794,N_1351,N_1876);
nor U2795 (N_2795,N_1210,N_1413);
and U2796 (N_2796,N_1806,N_1903);
nor U2797 (N_2797,N_1539,N_1908);
or U2798 (N_2798,N_1614,N_1309);
and U2799 (N_2799,N_1671,N_1712);
nand U2800 (N_2800,N_1854,N_1861);
or U2801 (N_2801,N_1273,N_1978);
nor U2802 (N_2802,N_1199,N_1377);
nor U2803 (N_2803,N_1655,N_1462);
nor U2804 (N_2804,N_1613,N_1926);
and U2805 (N_2805,N_1565,N_1235);
nand U2806 (N_2806,N_1948,N_1011);
or U2807 (N_2807,N_1215,N_1223);
nand U2808 (N_2808,N_1252,N_1968);
or U2809 (N_2809,N_1061,N_1603);
or U2810 (N_2810,N_1323,N_1775);
nor U2811 (N_2811,N_1032,N_1059);
nand U2812 (N_2812,N_1278,N_1581);
nand U2813 (N_2813,N_1482,N_1416);
and U2814 (N_2814,N_1353,N_1027);
or U2815 (N_2815,N_1901,N_1927);
nor U2816 (N_2816,N_1172,N_1604);
nor U2817 (N_2817,N_1754,N_1810);
nor U2818 (N_2818,N_1361,N_1635);
nor U2819 (N_2819,N_1717,N_1532);
nand U2820 (N_2820,N_1092,N_1783);
xnor U2821 (N_2821,N_1034,N_1217);
nor U2822 (N_2822,N_1312,N_1996);
or U2823 (N_2823,N_1650,N_1551);
nand U2824 (N_2824,N_1635,N_1501);
and U2825 (N_2825,N_1339,N_1081);
nand U2826 (N_2826,N_1947,N_1530);
nand U2827 (N_2827,N_1489,N_1623);
and U2828 (N_2828,N_1631,N_1606);
nor U2829 (N_2829,N_1668,N_1016);
nand U2830 (N_2830,N_1804,N_1312);
or U2831 (N_2831,N_1876,N_1666);
or U2832 (N_2832,N_1092,N_1286);
and U2833 (N_2833,N_1492,N_1608);
nand U2834 (N_2834,N_1329,N_1732);
and U2835 (N_2835,N_1545,N_1513);
and U2836 (N_2836,N_1847,N_1623);
or U2837 (N_2837,N_1213,N_1240);
nand U2838 (N_2838,N_1091,N_1436);
or U2839 (N_2839,N_1384,N_1159);
nand U2840 (N_2840,N_1586,N_1627);
nor U2841 (N_2841,N_1720,N_1494);
nand U2842 (N_2842,N_1330,N_1571);
nand U2843 (N_2843,N_1980,N_1818);
nand U2844 (N_2844,N_1485,N_1516);
nor U2845 (N_2845,N_1335,N_1004);
nand U2846 (N_2846,N_1496,N_1939);
or U2847 (N_2847,N_1771,N_1702);
or U2848 (N_2848,N_1805,N_1338);
and U2849 (N_2849,N_1734,N_1046);
nand U2850 (N_2850,N_1435,N_1596);
nor U2851 (N_2851,N_1994,N_1315);
nor U2852 (N_2852,N_1969,N_1588);
and U2853 (N_2853,N_1606,N_1783);
or U2854 (N_2854,N_1122,N_1913);
or U2855 (N_2855,N_1861,N_1980);
nand U2856 (N_2856,N_1883,N_1076);
nor U2857 (N_2857,N_1674,N_1606);
nand U2858 (N_2858,N_1539,N_1066);
nand U2859 (N_2859,N_1576,N_1374);
nand U2860 (N_2860,N_1293,N_1282);
or U2861 (N_2861,N_1679,N_1657);
or U2862 (N_2862,N_1174,N_1687);
or U2863 (N_2863,N_1706,N_1626);
nor U2864 (N_2864,N_1519,N_1913);
or U2865 (N_2865,N_1518,N_1453);
or U2866 (N_2866,N_1669,N_1935);
nor U2867 (N_2867,N_1422,N_1373);
nor U2868 (N_2868,N_1686,N_1017);
and U2869 (N_2869,N_1454,N_1433);
nand U2870 (N_2870,N_1213,N_1906);
nor U2871 (N_2871,N_1555,N_1986);
nor U2872 (N_2872,N_1916,N_1040);
nor U2873 (N_2873,N_1957,N_1369);
nand U2874 (N_2874,N_1557,N_1452);
nand U2875 (N_2875,N_1793,N_1908);
nor U2876 (N_2876,N_1781,N_1937);
nor U2877 (N_2877,N_1451,N_1576);
nor U2878 (N_2878,N_1032,N_1514);
nor U2879 (N_2879,N_1429,N_1045);
nand U2880 (N_2880,N_1146,N_1304);
nand U2881 (N_2881,N_1283,N_1508);
nor U2882 (N_2882,N_1056,N_1143);
and U2883 (N_2883,N_1234,N_1991);
nor U2884 (N_2884,N_1857,N_1318);
nor U2885 (N_2885,N_1766,N_1185);
nor U2886 (N_2886,N_1374,N_1080);
and U2887 (N_2887,N_1897,N_1719);
or U2888 (N_2888,N_1221,N_1262);
or U2889 (N_2889,N_1765,N_1897);
and U2890 (N_2890,N_1834,N_1824);
and U2891 (N_2891,N_1214,N_1809);
nor U2892 (N_2892,N_1756,N_1701);
nor U2893 (N_2893,N_1270,N_1670);
nand U2894 (N_2894,N_1743,N_1918);
or U2895 (N_2895,N_1339,N_1646);
nor U2896 (N_2896,N_1881,N_1773);
nor U2897 (N_2897,N_1168,N_1455);
or U2898 (N_2898,N_1812,N_1920);
and U2899 (N_2899,N_1385,N_1415);
or U2900 (N_2900,N_1685,N_1370);
and U2901 (N_2901,N_1947,N_1836);
or U2902 (N_2902,N_1844,N_1967);
nand U2903 (N_2903,N_1872,N_1382);
and U2904 (N_2904,N_1784,N_1581);
or U2905 (N_2905,N_1055,N_1150);
or U2906 (N_2906,N_1808,N_1613);
nand U2907 (N_2907,N_1878,N_1124);
and U2908 (N_2908,N_1574,N_1191);
or U2909 (N_2909,N_1879,N_1208);
or U2910 (N_2910,N_1868,N_1684);
nand U2911 (N_2911,N_1638,N_1364);
or U2912 (N_2912,N_1656,N_1549);
nor U2913 (N_2913,N_1788,N_1588);
nand U2914 (N_2914,N_1681,N_1612);
or U2915 (N_2915,N_1887,N_1014);
and U2916 (N_2916,N_1392,N_1113);
nand U2917 (N_2917,N_1121,N_1324);
nand U2918 (N_2918,N_1196,N_1397);
or U2919 (N_2919,N_1127,N_1031);
nand U2920 (N_2920,N_1276,N_1708);
nand U2921 (N_2921,N_1292,N_1852);
and U2922 (N_2922,N_1299,N_1708);
nor U2923 (N_2923,N_1988,N_1198);
and U2924 (N_2924,N_1221,N_1795);
nand U2925 (N_2925,N_1574,N_1275);
and U2926 (N_2926,N_1439,N_1728);
or U2927 (N_2927,N_1437,N_1256);
nand U2928 (N_2928,N_1179,N_1374);
or U2929 (N_2929,N_1006,N_1573);
nand U2930 (N_2930,N_1326,N_1969);
nor U2931 (N_2931,N_1437,N_1459);
nand U2932 (N_2932,N_1943,N_1874);
and U2933 (N_2933,N_1313,N_1386);
nor U2934 (N_2934,N_1552,N_1670);
and U2935 (N_2935,N_1607,N_1359);
or U2936 (N_2936,N_1826,N_1398);
nor U2937 (N_2937,N_1014,N_1613);
nor U2938 (N_2938,N_1128,N_1217);
or U2939 (N_2939,N_1551,N_1665);
nand U2940 (N_2940,N_1838,N_1024);
nand U2941 (N_2941,N_1610,N_1794);
nand U2942 (N_2942,N_1627,N_1723);
or U2943 (N_2943,N_1706,N_1016);
and U2944 (N_2944,N_1386,N_1747);
nor U2945 (N_2945,N_1375,N_1594);
nand U2946 (N_2946,N_1623,N_1431);
and U2947 (N_2947,N_1383,N_1827);
or U2948 (N_2948,N_1813,N_1856);
nand U2949 (N_2949,N_1100,N_1611);
and U2950 (N_2950,N_1510,N_1445);
and U2951 (N_2951,N_1247,N_1582);
or U2952 (N_2952,N_1065,N_1526);
nor U2953 (N_2953,N_1689,N_1957);
nand U2954 (N_2954,N_1260,N_1182);
nor U2955 (N_2955,N_1735,N_1341);
nand U2956 (N_2956,N_1976,N_1831);
nand U2957 (N_2957,N_1786,N_1054);
and U2958 (N_2958,N_1658,N_1249);
nor U2959 (N_2959,N_1754,N_1657);
and U2960 (N_2960,N_1923,N_1870);
and U2961 (N_2961,N_1300,N_1887);
nor U2962 (N_2962,N_1202,N_1973);
and U2963 (N_2963,N_1182,N_1414);
nor U2964 (N_2964,N_1678,N_1254);
or U2965 (N_2965,N_1065,N_1312);
and U2966 (N_2966,N_1111,N_1631);
nor U2967 (N_2967,N_1374,N_1681);
and U2968 (N_2968,N_1167,N_1423);
nor U2969 (N_2969,N_1144,N_1962);
nor U2970 (N_2970,N_1632,N_1469);
nand U2971 (N_2971,N_1528,N_1860);
and U2972 (N_2972,N_1847,N_1582);
nor U2973 (N_2973,N_1801,N_1391);
or U2974 (N_2974,N_1658,N_1758);
and U2975 (N_2975,N_1721,N_1460);
nand U2976 (N_2976,N_1762,N_1108);
or U2977 (N_2977,N_1415,N_1395);
nor U2978 (N_2978,N_1650,N_1802);
and U2979 (N_2979,N_1026,N_1865);
and U2980 (N_2980,N_1394,N_1827);
and U2981 (N_2981,N_1784,N_1933);
nor U2982 (N_2982,N_1356,N_1576);
nand U2983 (N_2983,N_1172,N_1665);
nand U2984 (N_2984,N_1995,N_1610);
and U2985 (N_2985,N_1467,N_1120);
nand U2986 (N_2986,N_1985,N_1512);
nor U2987 (N_2987,N_1152,N_1886);
and U2988 (N_2988,N_1652,N_1098);
nand U2989 (N_2989,N_1512,N_1152);
or U2990 (N_2990,N_1973,N_1170);
nand U2991 (N_2991,N_1974,N_1952);
or U2992 (N_2992,N_1931,N_1304);
and U2993 (N_2993,N_1812,N_1119);
nor U2994 (N_2994,N_1352,N_1313);
nand U2995 (N_2995,N_1191,N_1342);
nor U2996 (N_2996,N_1228,N_1991);
or U2997 (N_2997,N_1365,N_1177);
or U2998 (N_2998,N_1194,N_1915);
or U2999 (N_2999,N_1147,N_1763);
and U3000 (N_3000,N_2563,N_2644);
nand U3001 (N_3001,N_2979,N_2266);
nand U3002 (N_3002,N_2945,N_2334);
nor U3003 (N_3003,N_2865,N_2360);
or U3004 (N_3004,N_2798,N_2253);
nand U3005 (N_3005,N_2633,N_2053);
nor U3006 (N_3006,N_2961,N_2713);
and U3007 (N_3007,N_2920,N_2349);
and U3008 (N_3008,N_2246,N_2948);
and U3009 (N_3009,N_2696,N_2174);
and U3010 (N_3010,N_2373,N_2482);
nand U3011 (N_3011,N_2306,N_2512);
and U3012 (N_3012,N_2113,N_2216);
nand U3013 (N_3013,N_2523,N_2890);
or U3014 (N_3014,N_2518,N_2107);
nand U3015 (N_3015,N_2045,N_2269);
or U3016 (N_3016,N_2338,N_2263);
or U3017 (N_3017,N_2019,N_2176);
and U3018 (N_3018,N_2683,N_2316);
nor U3019 (N_3019,N_2913,N_2640);
and U3020 (N_3020,N_2483,N_2270);
or U3021 (N_3021,N_2943,N_2885);
or U3022 (N_3022,N_2503,N_2564);
nor U3023 (N_3023,N_2905,N_2576);
or U3024 (N_3024,N_2043,N_2211);
nand U3025 (N_3025,N_2379,N_2268);
or U3026 (N_3026,N_2023,N_2934);
nand U3027 (N_3027,N_2522,N_2343);
nor U3028 (N_3028,N_2685,N_2687);
nand U3029 (N_3029,N_2720,N_2042);
nand U3030 (N_3030,N_2093,N_2299);
nand U3031 (N_3031,N_2565,N_2327);
nor U3032 (N_3032,N_2096,N_2897);
nand U3033 (N_3033,N_2089,N_2131);
nor U3034 (N_3034,N_2645,N_2745);
or U3035 (N_3035,N_2006,N_2758);
nor U3036 (N_3036,N_2276,N_2147);
nor U3037 (N_3037,N_2915,N_2997);
nor U3038 (N_3038,N_2498,N_2212);
xnor U3039 (N_3039,N_2062,N_2097);
and U3040 (N_3040,N_2539,N_2844);
or U3041 (N_3041,N_2668,N_2724);
nand U3042 (N_3042,N_2110,N_2830);
nand U3043 (N_3043,N_2025,N_2846);
nand U3044 (N_3044,N_2970,N_2262);
nand U3045 (N_3045,N_2387,N_2479);
nand U3046 (N_3046,N_2529,N_2031);
and U3047 (N_3047,N_2455,N_2284);
nor U3048 (N_3048,N_2092,N_2257);
nand U3049 (N_3049,N_2021,N_2707);
or U3050 (N_3050,N_2350,N_2662);
or U3051 (N_3051,N_2091,N_2038);
and U3052 (N_3052,N_2171,N_2458);
and U3053 (N_3053,N_2793,N_2209);
and U3054 (N_3054,N_2572,N_2240);
nand U3055 (N_3055,N_2542,N_2590);
nand U3056 (N_3056,N_2095,N_2207);
and U3057 (N_3057,N_2944,N_2837);
and U3058 (N_3058,N_2872,N_2192);
nor U3059 (N_3059,N_2533,N_2695);
nor U3060 (N_3060,N_2251,N_2605);
and U3061 (N_3061,N_2610,N_2852);
or U3062 (N_3062,N_2868,N_2962);
nand U3063 (N_3063,N_2239,N_2421);
nor U3064 (N_3064,N_2549,N_2494);
or U3065 (N_3065,N_2362,N_2442);
and U3066 (N_3066,N_2711,N_2916);
and U3067 (N_3067,N_2666,N_2775);
and U3068 (N_3068,N_2465,N_2734);
or U3069 (N_3069,N_2799,N_2586);
nand U3070 (N_3070,N_2957,N_2649);
or U3071 (N_3071,N_2608,N_2675);
or U3072 (N_3072,N_2402,N_2480);
or U3073 (N_3073,N_2450,N_2892);
and U3074 (N_3074,N_2870,N_2908);
or U3075 (N_3075,N_2757,N_2861);
nor U3076 (N_3076,N_2098,N_2430);
nor U3077 (N_3077,N_2848,N_2158);
nand U3078 (N_3078,N_2302,N_2909);
nand U3079 (N_3079,N_2814,N_2635);
nand U3080 (N_3080,N_2462,N_2433);
and U3081 (N_3081,N_2500,N_2604);
and U3082 (N_3082,N_2028,N_2778);
and U3083 (N_3083,N_2153,N_2435);
nand U3084 (N_3084,N_2423,N_2030);
and U3085 (N_3085,N_2887,N_2833);
and U3086 (N_3086,N_2544,N_2759);
and U3087 (N_3087,N_2272,N_2161);
or U3088 (N_3088,N_2393,N_2700);
and U3089 (N_3089,N_2222,N_2034);
or U3090 (N_3090,N_2723,N_2762);
and U3091 (N_3091,N_2447,N_2806);
and U3092 (N_3092,N_2278,N_2352);
or U3093 (N_3093,N_2571,N_2875);
and U3094 (N_3094,N_2509,N_2477);
nor U3095 (N_3095,N_2203,N_2835);
nand U3096 (N_3096,N_2124,N_2754);
nand U3097 (N_3097,N_2871,N_2591);
or U3098 (N_3098,N_2528,N_2087);
or U3099 (N_3099,N_2172,N_2715);
and U3100 (N_3100,N_2893,N_2233);
nor U3101 (N_3101,N_2652,N_2204);
nor U3102 (N_3102,N_2526,N_2205);
and U3103 (N_3103,N_2156,N_2056);
xnor U3104 (N_3104,N_2150,N_2308);
or U3105 (N_3105,N_2128,N_2790);
nand U3106 (N_3106,N_2525,N_2785);
nor U3107 (N_3107,N_2543,N_2339);
nor U3108 (N_3108,N_2358,N_2927);
nand U3109 (N_3109,N_2322,N_2145);
nand U3110 (N_3110,N_2923,N_2742);
nand U3111 (N_3111,N_2795,N_2390);
and U3112 (N_3112,N_2653,N_2149);
nand U3113 (N_3113,N_2747,N_2285);
or U3114 (N_3114,N_2628,N_2142);
nor U3115 (N_3115,N_2002,N_2622);
or U3116 (N_3116,N_2228,N_2324);
and U3117 (N_3117,N_2751,N_2551);
or U3118 (N_3118,N_2679,N_2459);
nand U3119 (N_3119,N_2347,N_2736);
or U3120 (N_3120,N_2419,N_2527);
nor U3121 (N_3121,N_2474,N_2468);
nor U3122 (N_3122,N_2326,N_2954);
nand U3123 (N_3123,N_2295,N_2234);
nor U3124 (N_3124,N_2236,N_2705);
or U3125 (N_3125,N_2779,N_2190);
nand U3126 (N_3126,N_2189,N_2827);
or U3127 (N_3127,N_2426,N_2112);
nor U3128 (N_3128,N_2618,N_2063);
or U3129 (N_3129,N_2464,N_2496);
nand U3130 (N_3130,N_2606,N_2184);
or U3131 (N_3131,N_2703,N_2904);
nand U3132 (N_3132,N_2788,N_2587);
and U3133 (N_3133,N_2981,N_2655);
nor U3134 (N_3134,N_2810,N_2507);
or U3135 (N_3135,N_2422,N_2267);
or U3136 (N_3136,N_2414,N_2749);
or U3137 (N_3137,N_2227,N_2825);
or U3138 (N_3138,N_2561,N_2689);
nor U3139 (N_3139,N_2621,N_2613);
and U3140 (N_3140,N_2157,N_2667);
xnor U3141 (N_3141,N_2119,N_2508);
nor U3142 (N_3142,N_2714,N_2077);
nor U3143 (N_3143,N_2005,N_2701);
or U3144 (N_3144,N_2654,N_2947);
and U3145 (N_3145,N_2946,N_2824);
nor U3146 (N_3146,N_2213,N_2279);
nor U3147 (N_3147,N_2210,N_2804);
or U3148 (N_3148,N_2646,N_2869);
nand U3149 (N_3149,N_2173,N_2664);
nor U3150 (N_3150,N_2336,N_2318);
or U3151 (N_3151,N_2122,N_2364);
or U3152 (N_3152,N_2678,N_2601);
nand U3153 (N_3153,N_2004,N_2127);
or U3154 (N_3154,N_2039,N_2307);
nand U3155 (N_3155,N_2291,N_2412);
and U3156 (N_3156,N_2983,N_2388);
nand U3157 (N_3157,N_2047,N_2310);
nor U3158 (N_3158,N_2321,N_2155);
or U3159 (N_3159,N_2879,N_2367);
nor U3160 (N_3160,N_2922,N_2951);
and U3161 (N_3161,N_2688,N_2669);
nand U3162 (N_3162,N_2167,N_2037);
nor U3163 (N_3163,N_2116,N_2136);
or U3164 (N_3164,N_2193,N_2956);
and U3165 (N_3165,N_2516,N_2286);
and U3166 (N_3166,N_2218,N_2578);
nand U3167 (N_3167,N_2391,N_2287);
nor U3168 (N_3168,N_2152,N_2146);
nor U3169 (N_3169,N_2105,N_2012);
nor U3170 (N_3170,N_2860,N_2049);
nor U3171 (N_3171,N_2708,N_2650);
or U3172 (N_3172,N_2162,N_2449);
nor U3173 (N_3173,N_2581,N_2074);
nand U3174 (N_3174,N_2356,N_2394);
and U3175 (N_3175,N_2986,N_2050);
and U3176 (N_3176,N_2569,N_2014);
or U3177 (N_3177,N_2114,N_2169);
nand U3178 (N_3178,N_2020,N_2641);
nand U3179 (N_3179,N_2282,N_2382);
nand U3180 (N_3180,N_2540,N_2057);
and U3181 (N_3181,N_2598,N_2242);
or U3182 (N_3182,N_2249,N_2086);
and U3183 (N_3183,N_2671,N_2428);
or U3184 (N_3184,N_2882,N_2873);
or U3185 (N_3185,N_2822,N_2900);
nor U3186 (N_3186,N_2651,N_2936);
and U3187 (N_3187,N_2899,N_2809);
or U3188 (N_3188,N_2254,N_2225);
or U3189 (N_3189,N_2770,N_2118);
or U3190 (N_3190,N_2980,N_2933);
or U3191 (N_3191,N_2370,N_2315);
nor U3192 (N_3192,N_2492,N_2984);
or U3193 (N_3193,N_2369,N_2968);
nor U3194 (N_3194,N_2932,N_2530);
or U3195 (N_3195,N_2427,N_2235);
and U3196 (N_3196,N_2553,N_2763);
or U3197 (N_3197,N_2520,N_2015);
or U3198 (N_3198,N_2312,N_2230);
nor U3199 (N_3199,N_2555,N_2550);
nor U3200 (N_3200,N_2842,N_2612);
and U3201 (N_3201,N_2955,N_2958);
nor U3202 (N_3202,N_2300,N_2366);
nand U3203 (N_3203,N_2281,N_2994);
nor U3204 (N_3204,N_2656,N_2490);
nand U3205 (N_3205,N_2966,N_2752);
nand U3206 (N_3206,N_2297,N_2616);
nand U3207 (N_3207,N_2055,N_2374);
and U3208 (N_3208,N_2776,N_2241);
and U3209 (N_3209,N_2686,N_2126);
or U3210 (N_3210,N_2941,N_2461);
nand U3211 (N_3211,N_2260,N_2560);
or U3212 (N_3212,N_2454,N_2117);
nand U3213 (N_3213,N_2643,N_2780);
or U3214 (N_3214,N_2129,N_2987);
or U3215 (N_3215,N_2499,N_2008);
nor U3216 (N_3216,N_2907,N_2401);
nand U3217 (N_3217,N_2912,N_2585);
nand U3218 (N_3218,N_2371,N_2682);
or U3219 (N_3219,N_2817,N_2659);
or U3220 (N_3220,N_2631,N_2451);
and U3221 (N_3221,N_2769,N_2397);
and U3222 (N_3222,N_2022,N_2491);
nor U3223 (N_3223,N_2052,N_2416);
nor U3224 (N_3224,N_2130,N_2342);
nor U3225 (N_3225,N_2275,N_2384);
nand U3226 (N_3226,N_2629,N_2800);
and U3227 (N_3227,N_2739,N_2085);
nand U3228 (N_3228,N_2385,N_2383);
nand U3229 (N_3229,N_2977,N_2502);
or U3230 (N_3230,N_2903,N_2314);
nand U3231 (N_3231,N_2985,N_2960);
nand U3232 (N_3232,N_2568,N_2485);
nor U3233 (N_3233,N_2398,N_2144);
nand U3234 (N_3234,N_2989,N_2504);
nand U3235 (N_3235,N_2721,N_2058);
nand U3236 (N_3236,N_2988,N_2760);
or U3237 (N_3237,N_2570,N_2969);
nor U3238 (N_3238,N_2514,N_2791);
or U3239 (N_3239,N_2104,N_2737);
nand U3240 (N_3240,N_2313,N_2471);
or U3241 (N_3241,N_2993,N_2886);
or U3242 (N_3242,N_2141,N_2330);
nor U3243 (N_3243,N_2917,N_2614);
or U3244 (N_3244,N_2926,N_2726);
or U3245 (N_3245,N_2940,N_2493);
nand U3246 (N_3246,N_2148,N_2789);
or U3247 (N_3247,N_2888,N_2972);
nor U3248 (N_3248,N_2250,N_2575);
nor U3249 (N_3249,N_2594,N_2431);
and U3250 (N_3250,N_2611,N_2009);
nor U3251 (N_3251,N_2853,N_2625);
and U3252 (N_3252,N_2513,N_2756);
nor U3253 (N_3253,N_2335,N_2901);
and U3254 (N_3254,N_2252,N_2200);
nor U3255 (N_3255,N_2208,N_2929);
and U3256 (N_3256,N_2381,N_2185);
nand U3257 (N_3257,N_2935,N_2556);
or U3258 (N_3258,N_2186,N_2636);
and U3259 (N_3259,N_2329,N_2774);
or U3260 (N_3260,N_2247,N_2510);
nand U3261 (N_3261,N_2548,N_2079);
nand U3262 (N_3262,N_2854,N_2180);
and U3263 (N_3263,N_2755,N_2773);
or U3264 (N_3264,N_2473,N_2071);
nand U3265 (N_3265,N_2841,N_2928);
nand U3266 (N_3266,N_2624,N_2223);
and U3267 (N_3267,N_2102,N_2054);
nand U3268 (N_3268,N_2803,N_2201);
nand U3269 (N_3269,N_2365,N_2395);
nor U3270 (N_3270,N_2991,N_2566);
or U3271 (N_3271,N_2638,N_2998);
nor U3272 (N_3272,N_2567,N_2277);
or U3273 (N_3273,N_2206,N_2577);
nor U3274 (N_3274,N_2229,N_2851);
nor U3275 (N_3275,N_2432,N_2953);
nor U3276 (N_3276,N_2466,N_2469);
and U3277 (N_3277,N_2661,N_2690);
and U3278 (N_3278,N_2607,N_2066);
nand U3279 (N_3279,N_2821,N_2750);
nor U3280 (N_3280,N_2434,N_2084);
or U3281 (N_3281,N_2812,N_2697);
nand U3282 (N_3282,N_2163,N_2003);
or U3283 (N_3283,N_2475,N_2716);
and U3284 (N_3284,N_2808,N_2978);
and U3285 (N_3285,N_2215,N_2866);
nand U3286 (N_3286,N_2534,N_2709);
nand U3287 (N_3287,N_2733,N_2238);
and U3288 (N_3288,N_2036,N_2197);
nand U3289 (N_3289,N_2580,N_2761);
nor U3290 (N_3290,N_2202,N_2506);
nand U3291 (N_3291,N_2456,N_2748);
nand U3292 (N_3292,N_2328,N_2317);
nand U3293 (N_3293,N_2782,N_2883);
nor U3294 (N_3294,N_2546,N_2862);
nor U3295 (N_3295,N_2444,N_2361);
nor U3296 (N_3296,N_2858,N_2351);
nor U3297 (N_3297,N_2065,N_2845);
and U3298 (N_3298,N_2179,N_2354);
and U3299 (N_3299,N_2452,N_2293);
nor U3300 (N_3300,N_2348,N_2305);
nor U3301 (N_3301,N_2952,N_2368);
nor U3302 (N_3302,N_2040,N_2029);
nor U3303 (N_3303,N_2813,N_2424);
nor U3304 (N_3304,N_2674,N_2771);
nand U3305 (N_3305,N_2850,N_2392);
xnor U3306 (N_3306,N_2160,N_2436);
nand U3307 (N_3307,N_2467,N_2891);
and U3308 (N_3308,N_2959,N_2219);
nand U3309 (N_3309,N_2729,N_2072);
or U3310 (N_3310,N_2843,N_2289);
nor U3311 (N_3311,N_2874,N_2309);
nand U3312 (N_3312,N_2881,N_2670);
nor U3313 (N_3313,N_2743,N_2080);
or U3314 (N_3314,N_2797,N_2992);
or U3315 (N_3315,N_2898,N_2660);
nand U3316 (N_3316,N_2232,N_2376);
or U3317 (N_3317,N_2884,N_2088);
nor U3318 (N_3318,N_2864,N_2949);
nand U3319 (N_3319,N_2805,N_2115);
and U3320 (N_3320,N_2559,N_2722);
or U3321 (N_3321,N_2792,N_2880);
or U3322 (N_3322,N_2519,N_2658);
nor U3323 (N_3323,N_2133,N_2304);
nand U3324 (N_3324,N_2111,N_2290);
and U3325 (N_3325,N_2786,N_2386);
nand U3326 (N_3326,N_2914,N_2818);
or U3327 (N_3327,N_2815,N_2832);
nand U3328 (N_3328,N_2070,N_2017);
nor U3329 (N_3329,N_2829,N_2396);
nand U3330 (N_3330,N_2221,N_2271);
or U3331 (N_3331,N_2495,N_2630);
nor U3332 (N_3332,N_2692,N_2406);
or U3333 (N_3333,N_2712,N_2857);
nor U3334 (N_3334,N_2069,N_2060);
nor U3335 (N_3335,N_2637,N_2138);
and U3336 (N_3336,N_2151,N_2446);
and U3337 (N_3337,N_2178,N_2541);
nor U3338 (N_3338,N_2767,N_2831);
and U3339 (N_3339,N_2024,N_2083);
or U3340 (N_3340,N_2735,N_2521);
and U3341 (N_3341,N_2081,N_2856);
and U3342 (N_3342,N_2108,N_2663);
nor U3343 (N_3343,N_2413,N_2840);
or U3344 (N_3344,N_2226,N_2634);
nand U3345 (N_3345,N_2801,N_2274);
and U3346 (N_3346,N_2768,N_2702);
nand U3347 (N_3347,N_2681,N_2439);
nand U3348 (N_3348,N_2965,N_2602);
and U3349 (N_3349,N_2296,N_2501);
and U3350 (N_3350,N_2220,N_2007);
or U3351 (N_3351,N_2794,N_2517);
nand U3352 (N_3352,N_2265,N_2823);
or U3353 (N_3353,N_2481,N_2930);
or U3354 (N_3354,N_2429,N_2470);
nor U3355 (N_3355,N_2375,N_2411);
nor U3356 (N_3356,N_2632,N_2547);
and U3357 (N_3357,N_2438,N_2320);
and U3358 (N_3358,N_2018,N_2440);
nor U3359 (N_3359,N_2256,N_2583);
or U3360 (N_3360,N_2048,N_2694);
nand U3361 (N_3361,N_2013,N_2137);
or U3362 (N_3362,N_2340,N_2288);
and U3363 (N_3363,N_2710,N_2311);
or U3364 (N_3364,N_2698,N_2033);
nand U3365 (N_3365,N_2990,N_2816);
or U3366 (N_3366,N_2046,N_2363);
nand U3367 (N_3367,N_2766,N_2294);
and U3368 (N_3368,N_2380,N_2486);
or U3369 (N_3369,N_2532,N_2140);
or U3370 (N_3370,N_2731,N_2531);
nor U3371 (N_3371,N_2918,N_2472);
and U3372 (N_3372,N_2123,N_2337);
nand U3373 (N_3373,N_2906,N_2323);
or U3374 (N_3374,N_2772,N_2182);
nand U3375 (N_3375,N_2876,N_2214);
nand U3376 (N_3376,N_2836,N_2159);
nor U3377 (N_3377,N_2399,N_2963);
nand U3378 (N_3378,N_2718,N_2325);
or U3379 (N_3379,N_2691,N_2082);
and U3380 (N_3380,N_2765,N_2967);
and U3381 (N_3381,N_2258,N_2198);
nor U3382 (N_3382,N_2895,N_2199);
or U3383 (N_3383,N_2011,N_2417);
xnor U3384 (N_3384,N_2620,N_2244);
or U3385 (N_3385,N_2684,N_2976);
or U3386 (N_3386,N_2680,N_2725);
or U3387 (N_3387,N_2623,N_2041);
nor U3388 (N_3388,N_2068,N_2855);
and U3389 (N_3389,N_2188,N_2657);
nand U3390 (N_3390,N_2027,N_2164);
nand U3391 (N_3391,N_2699,N_2595);
or U3392 (N_3392,N_2125,N_2557);
nand U3393 (N_3393,N_2292,N_2971);
and U3394 (N_3394,N_2059,N_2617);
and U3395 (N_3395,N_2950,N_2728);
and U3396 (N_3396,N_2044,N_2443);
or U3397 (N_3397,N_2593,N_2919);
nor U3398 (N_3398,N_2974,N_2599);
or U3399 (N_3399,N_2582,N_2746);
or U3400 (N_3400,N_2341,N_2706);
nand U3401 (N_3401,N_2574,N_2896);
and U3402 (N_3402,N_2727,N_2497);
or U3403 (N_3403,N_2704,N_2937);
or U3404 (N_3404,N_2964,N_2925);
and U3405 (N_3405,N_2181,N_2921);
or U3406 (N_3406,N_2407,N_2639);
nand U3407 (N_3407,N_2484,N_2404);
nand U3408 (N_3408,N_2784,N_2120);
or U3409 (N_3409,N_2717,N_2828);
nor U3410 (N_3410,N_2359,N_2811);
or U3411 (N_3411,N_2243,N_2740);
nand U3412 (N_3412,N_2448,N_2524);
nand U3413 (N_3413,N_2353,N_2408);
nor U3414 (N_3414,N_2648,N_2942);
and U3415 (N_3415,N_2168,N_2738);
and U3416 (N_3416,N_2303,N_2996);
nand U3417 (N_3417,N_2558,N_2777);
nor U3418 (N_3418,N_2463,N_2418);
and U3419 (N_3419,N_2536,N_2597);
nand U3420 (N_3420,N_2103,N_2035);
or U3421 (N_3421,N_2819,N_2121);
nand U3422 (N_3422,N_2061,N_2999);
or U3423 (N_3423,N_2245,N_2511);
and U3424 (N_3424,N_2894,N_2378);
xnor U3425 (N_3425,N_2478,N_2787);
and U3426 (N_3426,N_2647,N_2377);
and U3427 (N_3427,N_2554,N_2672);
or U3428 (N_3428,N_2345,N_2280);
or U3429 (N_3429,N_2802,N_2902);
and U3430 (N_3430,N_2863,N_2589);
nand U3431 (N_3431,N_2409,N_2333);
or U3432 (N_3432,N_2489,N_2154);
nand U3433 (N_3433,N_2596,N_2165);
and U3434 (N_3434,N_2457,N_2826);
and U3435 (N_3435,N_2515,N_2372);
or U3436 (N_3436,N_2357,N_2217);
nor U3437 (N_3437,N_2859,N_2783);
nor U3438 (N_3438,N_2346,N_2973);
nand U3439 (N_3439,N_2183,N_2051);
nor U3440 (N_3440,N_2505,N_2139);
or U3441 (N_3441,N_2237,N_2231);
or U3442 (N_3442,N_2441,N_2255);
and U3443 (N_3443,N_2642,N_2588);
nand U3444 (N_3444,N_2283,N_2403);
and U3445 (N_3445,N_2938,N_2834);
nor U3446 (N_3446,N_2400,N_2191);
and U3447 (N_3447,N_2562,N_2807);
and U3448 (N_3448,N_2796,N_2545);
nor U3449 (N_3449,N_2273,N_2355);
nand U3450 (N_3450,N_2298,N_2248);
nand U3451 (N_3451,N_2878,N_2719);
nor U3452 (N_3452,N_2109,N_2910);
nor U3453 (N_3453,N_2820,N_2078);
nand U3454 (N_3454,N_2982,N_2741);
or U3455 (N_3455,N_2838,N_2101);
nor U3456 (N_3456,N_2626,N_2665);
nand U3457 (N_3457,N_2301,N_2445);
nand U3458 (N_3458,N_2732,N_2143);
or U3459 (N_3459,N_2744,N_2753);
nor U3460 (N_3460,N_2537,N_2389);
nor U3461 (N_3461,N_2259,N_2877);
or U3462 (N_3462,N_2405,N_2781);
and U3463 (N_3463,N_2420,N_2332);
nor U3464 (N_3464,N_2839,N_2619);
nor U3465 (N_3465,N_2135,N_2924);
nor U3466 (N_3466,N_2195,N_2194);
nand U3467 (N_3467,N_2488,N_2975);
or U3468 (N_3468,N_2187,N_2166);
or U3469 (N_3469,N_2693,N_2073);
nand U3470 (N_3470,N_2175,N_2931);
and U3471 (N_3471,N_2331,N_2592);
or U3472 (N_3472,N_2170,N_2132);
nor U3473 (N_3473,N_2026,N_2579);
and U3474 (N_3474,N_2261,N_2196);
nor U3475 (N_3475,N_2425,N_2867);
nor U3476 (N_3476,N_2911,N_2476);
nor U3477 (N_3477,N_2615,N_2076);
or U3478 (N_3478,N_2487,N_2677);
or U3479 (N_3479,N_2538,N_2415);
and U3480 (N_3480,N_2224,N_2090);
nand U3481 (N_3481,N_2460,N_2000);
nand U3482 (N_3482,N_2410,N_2344);
or U3483 (N_3483,N_2064,N_2603);
nand U3484 (N_3484,N_2453,N_2075);
nand U3485 (N_3485,N_2177,N_2995);
nor U3486 (N_3486,N_2535,N_2627);
nand U3487 (N_3487,N_2889,N_2010);
nand U3488 (N_3488,N_2100,N_2032);
and U3489 (N_3489,N_2067,N_2094);
and U3490 (N_3490,N_2584,N_2016);
nand U3491 (N_3491,N_2673,N_2849);
nand U3492 (N_3492,N_2573,N_2134);
and U3493 (N_3493,N_2847,N_2437);
nand U3494 (N_3494,N_2939,N_2001);
or U3495 (N_3495,N_2106,N_2099);
and U3496 (N_3496,N_2552,N_2264);
nand U3497 (N_3497,N_2609,N_2676);
nor U3498 (N_3498,N_2600,N_2319);
and U3499 (N_3499,N_2764,N_2730);
nand U3500 (N_3500,N_2535,N_2224);
or U3501 (N_3501,N_2609,N_2145);
nor U3502 (N_3502,N_2595,N_2826);
and U3503 (N_3503,N_2191,N_2671);
or U3504 (N_3504,N_2624,N_2694);
nor U3505 (N_3505,N_2518,N_2509);
or U3506 (N_3506,N_2670,N_2100);
nor U3507 (N_3507,N_2968,N_2102);
or U3508 (N_3508,N_2029,N_2893);
nand U3509 (N_3509,N_2343,N_2896);
nand U3510 (N_3510,N_2037,N_2168);
nor U3511 (N_3511,N_2385,N_2619);
and U3512 (N_3512,N_2055,N_2362);
nand U3513 (N_3513,N_2346,N_2790);
and U3514 (N_3514,N_2576,N_2873);
or U3515 (N_3515,N_2365,N_2559);
nor U3516 (N_3516,N_2142,N_2215);
or U3517 (N_3517,N_2236,N_2533);
and U3518 (N_3518,N_2772,N_2284);
nor U3519 (N_3519,N_2924,N_2489);
nor U3520 (N_3520,N_2880,N_2509);
nor U3521 (N_3521,N_2566,N_2800);
nand U3522 (N_3522,N_2351,N_2433);
and U3523 (N_3523,N_2306,N_2621);
or U3524 (N_3524,N_2283,N_2974);
nand U3525 (N_3525,N_2023,N_2003);
and U3526 (N_3526,N_2327,N_2461);
nor U3527 (N_3527,N_2605,N_2811);
and U3528 (N_3528,N_2910,N_2387);
and U3529 (N_3529,N_2560,N_2377);
nor U3530 (N_3530,N_2921,N_2133);
nand U3531 (N_3531,N_2340,N_2649);
nand U3532 (N_3532,N_2770,N_2558);
nand U3533 (N_3533,N_2148,N_2264);
or U3534 (N_3534,N_2069,N_2829);
and U3535 (N_3535,N_2333,N_2189);
nor U3536 (N_3536,N_2619,N_2866);
and U3537 (N_3537,N_2005,N_2810);
nor U3538 (N_3538,N_2580,N_2276);
nor U3539 (N_3539,N_2110,N_2315);
nor U3540 (N_3540,N_2720,N_2398);
or U3541 (N_3541,N_2363,N_2594);
or U3542 (N_3542,N_2732,N_2454);
nor U3543 (N_3543,N_2175,N_2582);
nor U3544 (N_3544,N_2375,N_2271);
or U3545 (N_3545,N_2955,N_2920);
nand U3546 (N_3546,N_2499,N_2095);
nor U3547 (N_3547,N_2630,N_2018);
nand U3548 (N_3548,N_2858,N_2503);
or U3549 (N_3549,N_2463,N_2081);
and U3550 (N_3550,N_2462,N_2668);
and U3551 (N_3551,N_2536,N_2450);
nand U3552 (N_3552,N_2019,N_2084);
nand U3553 (N_3553,N_2325,N_2461);
or U3554 (N_3554,N_2578,N_2425);
and U3555 (N_3555,N_2347,N_2031);
nor U3556 (N_3556,N_2399,N_2820);
or U3557 (N_3557,N_2017,N_2720);
nand U3558 (N_3558,N_2598,N_2903);
or U3559 (N_3559,N_2315,N_2213);
nor U3560 (N_3560,N_2915,N_2333);
or U3561 (N_3561,N_2505,N_2238);
or U3562 (N_3562,N_2008,N_2301);
nand U3563 (N_3563,N_2862,N_2058);
or U3564 (N_3564,N_2101,N_2753);
or U3565 (N_3565,N_2047,N_2392);
and U3566 (N_3566,N_2039,N_2273);
nand U3567 (N_3567,N_2688,N_2853);
nor U3568 (N_3568,N_2126,N_2897);
or U3569 (N_3569,N_2216,N_2001);
nor U3570 (N_3570,N_2476,N_2101);
xnor U3571 (N_3571,N_2061,N_2616);
or U3572 (N_3572,N_2183,N_2064);
and U3573 (N_3573,N_2909,N_2748);
or U3574 (N_3574,N_2895,N_2702);
and U3575 (N_3575,N_2742,N_2709);
nand U3576 (N_3576,N_2080,N_2591);
nand U3577 (N_3577,N_2238,N_2443);
or U3578 (N_3578,N_2215,N_2809);
nand U3579 (N_3579,N_2498,N_2660);
nor U3580 (N_3580,N_2161,N_2580);
nand U3581 (N_3581,N_2404,N_2897);
nor U3582 (N_3582,N_2215,N_2041);
or U3583 (N_3583,N_2588,N_2118);
and U3584 (N_3584,N_2384,N_2200);
and U3585 (N_3585,N_2689,N_2150);
nand U3586 (N_3586,N_2147,N_2021);
and U3587 (N_3587,N_2690,N_2480);
nor U3588 (N_3588,N_2573,N_2252);
or U3589 (N_3589,N_2875,N_2835);
and U3590 (N_3590,N_2797,N_2204);
nand U3591 (N_3591,N_2680,N_2796);
nor U3592 (N_3592,N_2094,N_2980);
nand U3593 (N_3593,N_2217,N_2899);
nand U3594 (N_3594,N_2079,N_2334);
or U3595 (N_3595,N_2393,N_2812);
and U3596 (N_3596,N_2405,N_2114);
nor U3597 (N_3597,N_2230,N_2155);
nand U3598 (N_3598,N_2294,N_2205);
or U3599 (N_3599,N_2134,N_2831);
nor U3600 (N_3600,N_2284,N_2138);
and U3601 (N_3601,N_2413,N_2995);
nand U3602 (N_3602,N_2533,N_2089);
and U3603 (N_3603,N_2703,N_2753);
nand U3604 (N_3604,N_2981,N_2535);
nor U3605 (N_3605,N_2219,N_2583);
or U3606 (N_3606,N_2600,N_2141);
or U3607 (N_3607,N_2369,N_2785);
nand U3608 (N_3608,N_2266,N_2537);
and U3609 (N_3609,N_2968,N_2757);
nand U3610 (N_3610,N_2329,N_2775);
or U3611 (N_3611,N_2948,N_2814);
nand U3612 (N_3612,N_2958,N_2213);
nand U3613 (N_3613,N_2150,N_2041);
nand U3614 (N_3614,N_2853,N_2822);
or U3615 (N_3615,N_2667,N_2670);
and U3616 (N_3616,N_2512,N_2231);
or U3617 (N_3617,N_2702,N_2422);
nor U3618 (N_3618,N_2462,N_2239);
nand U3619 (N_3619,N_2331,N_2926);
nor U3620 (N_3620,N_2354,N_2898);
and U3621 (N_3621,N_2990,N_2919);
nor U3622 (N_3622,N_2913,N_2129);
or U3623 (N_3623,N_2351,N_2225);
and U3624 (N_3624,N_2283,N_2316);
nor U3625 (N_3625,N_2086,N_2568);
nand U3626 (N_3626,N_2112,N_2061);
nor U3627 (N_3627,N_2899,N_2712);
or U3628 (N_3628,N_2429,N_2867);
and U3629 (N_3629,N_2608,N_2519);
and U3630 (N_3630,N_2570,N_2109);
or U3631 (N_3631,N_2084,N_2459);
xor U3632 (N_3632,N_2722,N_2493);
nor U3633 (N_3633,N_2309,N_2317);
or U3634 (N_3634,N_2563,N_2109);
or U3635 (N_3635,N_2638,N_2957);
and U3636 (N_3636,N_2891,N_2544);
nor U3637 (N_3637,N_2485,N_2633);
and U3638 (N_3638,N_2645,N_2963);
or U3639 (N_3639,N_2180,N_2706);
or U3640 (N_3640,N_2582,N_2758);
and U3641 (N_3641,N_2668,N_2310);
and U3642 (N_3642,N_2477,N_2859);
nor U3643 (N_3643,N_2651,N_2136);
nand U3644 (N_3644,N_2261,N_2105);
nor U3645 (N_3645,N_2422,N_2175);
nand U3646 (N_3646,N_2200,N_2367);
nor U3647 (N_3647,N_2809,N_2415);
or U3648 (N_3648,N_2266,N_2543);
and U3649 (N_3649,N_2649,N_2388);
xnor U3650 (N_3650,N_2414,N_2512);
nor U3651 (N_3651,N_2375,N_2040);
nor U3652 (N_3652,N_2590,N_2742);
nor U3653 (N_3653,N_2024,N_2899);
nor U3654 (N_3654,N_2007,N_2605);
and U3655 (N_3655,N_2083,N_2453);
and U3656 (N_3656,N_2451,N_2619);
and U3657 (N_3657,N_2007,N_2296);
and U3658 (N_3658,N_2093,N_2350);
or U3659 (N_3659,N_2222,N_2775);
nand U3660 (N_3660,N_2694,N_2268);
nor U3661 (N_3661,N_2420,N_2359);
nand U3662 (N_3662,N_2938,N_2059);
nand U3663 (N_3663,N_2602,N_2296);
nor U3664 (N_3664,N_2825,N_2466);
nand U3665 (N_3665,N_2538,N_2064);
or U3666 (N_3666,N_2283,N_2246);
nor U3667 (N_3667,N_2542,N_2749);
nand U3668 (N_3668,N_2452,N_2017);
nand U3669 (N_3669,N_2467,N_2091);
nor U3670 (N_3670,N_2558,N_2097);
nor U3671 (N_3671,N_2412,N_2601);
and U3672 (N_3672,N_2442,N_2115);
and U3673 (N_3673,N_2205,N_2004);
nand U3674 (N_3674,N_2034,N_2411);
or U3675 (N_3675,N_2523,N_2491);
nor U3676 (N_3676,N_2898,N_2454);
and U3677 (N_3677,N_2306,N_2981);
and U3678 (N_3678,N_2208,N_2020);
nor U3679 (N_3679,N_2407,N_2929);
nor U3680 (N_3680,N_2910,N_2798);
nor U3681 (N_3681,N_2812,N_2461);
nor U3682 (N_3682,N_2914,N_2499);
nand U3683 (N_3683,N_2985,N_2282);
or U3684 (N_3684,N_2030,N_2314);
and U3685 (N_3685,N_2641,N_2601);
nor U3686 (N_3686,N_2913,N_2806);
nand U3687 (N_3687,N_2915,N_2316);
or U3688 (N_3688,N_2976,N_2920);
or U3689 (N_3689,N_2096,N_2068);
nand U3690 (N_3690,N_2545,N_2403);
and U3691 (N_3691,N_2495,N_2755);
nor U3692 (N_3692,N_2482,N_2182);
and U3693 (N_3693,N_2542,N_2473);
or U3694 (N_3694,N_2296,N_2200);
nand U3695 (N_3695,N_2798,N_2448);
nand U3696 (N_3696,N_2027,N_2110);
nand U3697 (N_3697,N_2336,N_2152);
nand U3698 (N_3698,N_2382,N_2850);
nand U3699 (N_3699,N_2130,N_2542);
nor U3700 (N_3700,N_2965,N_2610);
nand U3701 (N_3701,N_2221,N_2716);
nor U3702 (N_3702,N_2327,N_2788);
or U3703 (N_3703,N_2594,N_2129);
or U3704 (N_3704,N_2279,N_2319);
nor U3705 (N_3705,N_2285,N_2473);
or U3706 (N_3706,N_2707,N_2868);
nor U3707 (N_3707,N_2641,N_2893);
and U3708 (N_3708,N_2783,N_2991);
nor U3709 (N_3709,N_2039,N_2777);
or U3710 (N_3710,N_2209,N_2812);
or U3711 (N_3711,N_2014,N_2161);
or U3712 (N_3712,N_2650,N_2677);
or U3713 (N_3713,N_2124,N_2686);
nor U3714 (N_3714,N_2486,N_2534);
or U3715 (N_3715,N_2909,N_2841);
xnor U3716 (N_3716,N_2839,N_2648);
and U3717 (N_3717,N_2852,N_2047);
and U3718 (N_3718,N_2207,N_2432);
and U3719 (N_3719,N_2708,N_2566);
nor U3720 (N_3720,N_2314,N_2039);
nand U3721 (N_3721,N_2909,N_2967);
nor U3722 (N_3722,N_2184,N_2506);
nand U3723 (N_3723,N_2078,N_2900);
and U3724 (N_3724,N_2003,N_2220);
nor U3725 (N_3725,N_2224,N_2789);
nor U3726 (N_3726,N_2600,N_2515);
nor U3727 (N_3727,N_2778,N_2736);
and U3728 (N_3728,N_2320,N_2493);
nand U3729 (N_3729,N_2755,N_2129);
or U3730 (N_3730,N_2448,N_2881);
nor U3731 (N_3731,N_2155,N_2627);
or U3732 (N_3732,N_2836,N_2739);
nor U3733 (N_3733,N_2845,N_2037);
nand U3734 (N_3734,N_2702,N_2799);
or U3735 (N_3735,N_2045,N_2786);
nor U3736 (N_3736,N_2689,N_2297);
nor U3737 (N_3737,N_2694,N_2188);
or U3738 (N_3738,N_2008,N_2105);
and U3739 (N_3739,N_2222,N_2995);
nand U3740 (N_3740,N_2075,N_2554);
nor U3741 (N_3741,N_2874,N_2769);
nand U3742 (N_3742,N_2344,N_2697);
nand U3743 (N_3743,N_2430,N_2122);
or U3744 (N_3744,N_2791,N_2419);
nor U3745 (N_3745,N_2058,N_2826);
and U3746 (N_3746,N_2520,N_2121);
nand U3747 (N_3747,N_2191,N_2957);
nor U3748 (N_3748,N_2496,N_2105);
nor U3749 (N_3749,N_2311,N_2233);
and U3750 (N_3750,N_2087,N_2332);
nand U3751 (N_3751,N_2869,N_2828);
nand U3752 (N_3752,N_2776,N_2247);
nor U3753 (N_3753,N_2486,N_2213);
nor U3754 (N_3754,N_2647,N_2284);
nand U3755 (N_3755,N_2236,N_2093);
and U3756 (N_3756,N_2217,N_2684);
and U3757 (N_3757,N_2845,N_2251);
and U3758 (N_3758,N_2194,N_2607);
nand U3759 (N_3759,N_2342,N_2419);
nor U3760 (N_3760,N_2870,N_2880);
or U3761 (N_3761,N_2922,N_2744);
nand U3762 (N_3762,N_2234,N_2592);
nor U3763 (N_3763,N_2520,N_2715);
or U3764 (N_3764,N_2380,N_2291);
or U3765 (N_3765,N_2565,N_2912);
nor U3766 (N_3766,N_2619,N_2555);
and U3767 (N_3767,N_2857,N_2682);
and U3768 (N_3768,N_2233,N_2354);
and U3769 (N_3769,N_2989,N_2342);
or U3770 (N_3770,N_2427,N_2238);
nand U3771 (N_3771,N_2429,N_2347);
or U3772 (N_3772,N_2262,N_2406);
and U3773 (N_3773,N_2010,N_2311);
and U3774 (N_3774,N_2203,N_2576);
nand U3775 (N_3775,N_2588,N_2499);
and U3776 (N_3776,N_2822,N_2763);
or U3777 (N_3777,N_2402,N_2564);
or U3778 (N_3778,N_2855,N_2990);
or U3779 (N_3779,N_2712,N_2086);
nand U3780 (N_3780,N_2435,N_2396);
nor U3781 (N_3781,N_2409,N_2628);
and U3782 (N_3782,N_2290,N_2506);
nand U3783 (N_3783,N_2838,N_2085);
or U3784 (N_3784,N_2193,N_2004);
nor U3785 (N_3785,N_2929,N_2031);
nor U3786 (N_3786,N_2629,N_2009);
and U3787 (N_3787,N_2978,N_2958);
or U3788 (N_3788,N_2303,N_2334);
nand U3789 (N_3789,N_2186,N_2008);
nor U3790 (N_3790,N_2252,N_2067);
and U3791 (N_3791,N_2096,N_2257);
or U3792 (N_3792,N_2611,N_2952);
nor U3793 (N_3793,N_2133,N_2033);
nor U3794 (N_3794,N_2074,N_2918);
and U3795 (N_3795,N_2690,N_2775);
or U3796 (N_3796,N_2295,N_2198);
nor U3797 (N_3797,N_2151,N_2126);
or U3798 (N_3798,N_2971,N_2509);
xnor U3799 (N_3799,N_2463,N_2572);
or U3800 (N_3800,N_2494,N_2586);
or U3801 (N_3801,N_2739,N_2632);
nor U3802 (N_3802,N_2336,N_2896);
or U3803 (N_3803,N_2761,N_2462);
nand U3804 (N_3804,N_2928,N_2027);
or U3805 (N_3805,N_2603,N_2363);
nand U3806 (N_3806,N_2077,N_2195);
nand U3807 (N_3807,N_2143,N_2020);
nand U3808 (N_3808,N_2564,N_2236);
or U3809 (N_3809,N_2552,N_2886);
or U3810 (N_3810,N_2168,N_2543);
nor U3811 (N_3811,N_2108,N_2466);
and U3812 (N_3812,N_2436,N_2446);
nand U3813 (N_3813,N_2969,N_2794);
or U3814 (N_3814,N_2737,N_2448);
or U3815 (N_3815,N_2810,N_2768);
and U3816 (N_3816,N_2280,N_2499);
or U3817 (N_3817,N_2860,N_2217);
or U3818 (N_3818,N_2780,N_2184);
and U3819 (N_3819,N_2204,N_2234);
nand U3820 (N_3820,N_2730,N_2440);
nand U3821 (N_3821,N_2409,N_2494);
or U3822 (N_3822,N_2055,N_2095);
and U3823 (N_3823,N_2590,N_2534);
xor U3824 (N_3824,N_2700,N_2915);
or U3825 (N_3825,N_2294,N_2549);
or U3826 (N_3826,N_2572,N_2393);
nand U3827 (N_3827,N_2515,N_2013);
nor U3828 (N_3828,N_2436,N_2832);
or U3829 (N_3829,N_2034,N_2731);
nand U3830 (N_3830,N_2204,N_2724);
or U3831 (N_3831,N_2301,N_2681);
and U3832 (N_3832,N_2804,N_2672);
nor U3833 (N_3833,N_2749,N_2086);
nand U3834 (N_3834,N_2490,N_2013);
and U3835 (N_3835,N_2045,N_2977);
or U3836 (N_3836,N_2710,N_2016);
or U3837 (N_3837,N_2899,N_2041);
and U3838 (N_3838,N_2970,N_2643);
or U3839 (N_3839,N_2434,N_2936);
nand U3840 (N_3840,N_2604,N_2171);
and U3841 (N_3841,N_2968,N_2786);
and U3842 (N_3842,N_2539,N_2258);
or U3843 (N_3843,N_2002,N_2164);
or U3844 (N_3844,N_2296,N_2054);
nand U3845 (N_3845,N_2030,N_2021);
nand U3846 (N_3846,N_2805,N_2681);
nand U3847 (N_3847,N_2244,N_2378);
nor U3848 (N_3848,N_2526,N_2822);
nor U3849 (N_3849,N_2072,N_2756);
nor U3850 (N_3850,N_2236,N_2864);
and U3851 (N_3851,N_2107,N_2655);
nor U3852 (N_3852,N_2591,N_2975);
nor U3853 (N_3853,N_2610,N_2951);
nor U3854 (N_3854,N_2085,N_2805);
nor U3855 (N_3855,N_2027,N_2216);
or U3856 (N_3856,N_2216,N_2500);
and U3857 (N_3857,N_2215,N_2515);
nor U3858 (N_3858,N_2759,N_2804);
nand U3859 (N_3859,N_2592,N_2808);
nor U3860 (N_3860,N_2967,N_2177);
and U3861 (N_3861,N_2588,N_2771);
nor U3862 (N_3862,N_2273,N_2304);
or U3863 (N_3863,N_2124,N_2759);
nand U3864 (N_3864,N_2629,N_2417);
or U3865 (N_3865,N_2469,N_2135);
or U3866 (N_3866,N_2660,N_2897);
or U3867 (N_3867,N_2653,N_2660);
nor U3868 (N_3868,N_2153,N_2023);
and U3869 (N_3869,N_2109,N_2922);
nor U3870 (N_3870,N_2657,N_2413);
and U3871 (N_3871,N_2152,N_2363);
nor U3872 (N_3872,N_2946,N_2792);
nor U3873 (N_3873,N_2884,N_2639);
nor U3874 (N_3874,N_2873,N_2974);
nor U3875 (N_3875,N_2568,N_2896);
or U3876 (N_3876,N_2267,N_2530);
or U3877 (N_3877,N_2513,N_2090);
nor U3878 (N_3878,N_2180,N_2196);
or U3879 (N_3879,N_2857,N_2830);
and U3880 (N_3880,N_2104,N_2330);
nor U3881 (N_3881,N_2015,N_2583);
and U3882 (N_3882,N_2661,N_2898);
nor U3883 (N_3883,N_2953,N_2797);
and U3884 (N_3884,N_2041,N_2036);
and U3885 (N_3885,N_2788,N_2485);
or U3886 (N_3886,N_2085,N_2220);
nand U3887 (N_3887,N_2661,N_2745);
nor U3888 (N_3888,N_2341,N_2088);
or U3889 (N_3889,N_2120,N_2466);
and U3890 (N_3890,N_2819,N_2959);
and U3891 (N_3891,N_2521,N_2284);
and U3892 (N_3892,N_2821,N_2855);
nand U3893 (N_3893,N_2854,N_2120);
and U3894 (N_3894,N_2649,N_2721);
nand U3895 (N_3895,N_2036,N_2004);
and U3896 (N_3896,N_2206,N_2189);
nor U3897 (N_3897,N_2770,N_2975);
and U3898 (N_3898,N_2110,N_2142);
and U3899 (N_3899,N_2664,N_2114);
nor U3900 (N_3900,N_2422,N_2898);
nand U3901 (N_3901,N_2280,N_2166);
nor U3902 (N_3902,N_2730,N_2777);
or U3903 (N_3903,N_2377,N_2549);
or U3904 (N_3904,N_2246,N_2724);
or U3905 (N_3905,N_2239,N_2242);
nor U3906 (N_3906,N_2414,N_2443);
nor U3907 (N_3907,N_2827,N_2536);
nor U3908 (N_3908,N_2827,N_2413);
and U3909 (N_3909,N_2685,N_2923);
and U3910 (N_3910,N_2426,N_2754);
and U3911 (N_3911,N_2919,N_2208);
nand U3912 (N_3912,N_2292,N_2470);
or U3913 (N_3913,N_2287,N_2070);
nor U3914 (N_3914,N_2526,N_2435);
nand U3915 (N_3915,N_2736,N_2132);
nand U3916 (N_3916,N_2238,N_2831);
nor U3917 (N_3917,N_2155,N_2723);
and U3918 (N_3918,N_2979,N_2366);
nor U3919 (N_3919,N_2205,N_2859);
or U3920 (N_3920,N_2408,N_2469);
nor U3921 (N_3921,N_2162,N_2810);
nand U3922 (N_3922,N_2019,N_2751);
or U3923 (N_3923,N_2432,N_2296);
and U3924 (N_3924,N_2051,N_2200);
or U3925 (N_3925,N_2304,N_2270);
and U3926 (N_3926,N_2626,N_2988);
or U3927 (N_3927,N_2653,N_2368);
nor U3928 (N_3928,N_2839,N_2313);
nand U3929 (N_3929,N_2620,N_2248);
and U3930 (N_3930,N_2769,N_2786);
nor U3931 (N_3931,N_2022,N_2822);
and U3932 (N_3932,N_2023,N_2901);
xor U3933 (N_3933,N_2495,N_2954);
and U3934 (N_3934,N_2179,N_2233);
nor U3935 (N_3935,N_2756,N_2041);
or U3936 (N_3936,N_2695,N_2335);
nor U3937 (N_3937,N_2219,N_2530);
or U3938 (N_3938,N_2882,N_2157);
or U3939 (N_3939,N_2187,N_2231);
or U3940 (N_3940,N_2515,N_2562);
or U3941 (N_3941,N_2096,N_2457);
nand U3942 (N_3942,N_2750,N_2988);
nand U3943 (N_3943,N_2050,N_2715);
nand U3944 (N_3944,N_2724,N_2281);
nor U3945 (N_3945,N_2769,N_2100);
nand U3946 (N_3946,N_2234,N_2855);
nor U3947 (N_3947,N_2437,N_2172);
nor U3948 (N_3948,N_2315,N_2361);
nor U3949 (N_3949,N_2594,N_2002);
or U3950 (N_3950,N_2207,N_2076);
nand U3951 (N_3951,N_2150,N_2847);
or U3952 (N_3952,N_2204,N_2285);
nor U3953 (N_3953,N_2666,N_2989);
nor U3954 (N_3954,N_2231,N_2038);
nor U3955 (N_3955,N_2819,N_2507);
nor U3956 (N_3956,N_2152,N_2171);
and U3957 (N_3957,N_2746,N_2190);
and U3958 (N_3958,N_2307,N_2806);
or U3959 (N_3959,N_2777,N_2144);
and U3960 (N_3960,N_2902,N_2302);
nand U3961 (N_3961,N_2881,N_2160);
nor U3962 (N_3962,N_2910,N_2191);
and U3963 (N_3963,N_2837,N_2402);
nand U3964 (N_3964,N_2472,N_2542);
or U3965 (N_3965,N_2438,N_2887);
and U3966 (N_3966,N_2085,N_2440);
or U3967 (N_3967,N_2961,N_2788);
or U3968 (N_3968,N_2948,N_2236);
and U3969 (N_3969,N_2083,N_2914);
nor U3970 (N_3970,N_2382,N_2216);
nand U3971 (N_3971,N_2850,N_2512);
nor U3972 (N_3972,N_2186,N_2072);
nand U3973 (N_3973,N_2900,N_2211);
and U3974 (N_3974,N_2839,N_2986);
or U3975 (N_3975,N_2432,N_2033);
nand U3976 (N_3976,N_2908,N_2880);
nand U3977 (N_3977,N_2528,N_2369);
and U3978 (N_3978,N_2326,N_2379);
nor U3979 (N_3979,N_2452,N_2750);
nand U3980 (N_3980,N_2668,N_2023);
nor U3981 (N_3981,N_2632,N_2088);
nand U3982 (N_3982,N_2191,N_2643);
or U3983 (N_3983,N_2458,N_2742);
nand U3984 (N_3984,N_2844,N_2598);
and U3985 (N_3985,N_2688,N_2761);
nor U3986 (N_3986,N_2634,N_2668);
or U3987 (N_3987,N_2301,N_2320);
nor U3988 (N_3988,N_2236,N_2000);
or U3989 (N_3989,N_2029,N_2057);
nand U3990 (N_3990,N_2048,N_2584);
and U3991 (N_3991,N_2234,N_2307);
nand U3992 (N_3992,N_2638,N_2594);
and U3993 (N_3993,N_2051,N_2889);
or U3994 (N_3994,N_2840,N_2858);
nand U3995 (N_3995,N_2967,N_2921);
or U3996 (N_3996,N_2638,N_2507);
nand U3997 (N_3997,N_2875,N_2500);
nor U3998 (N_3998,N_2251,N_2770);
xnor U3999 (N_3999,N_2512,N_2904);
or U4000 (N_4000,N_3479,N_3069);
or U4001 (N_4001,N_3303,N_3317);
nor U4002 (N_4002,N_3223,N_3851);
or U4003 (N_4003,N_3427,N_3762);
and U4004 (N_4004,N_3122,N_3170);
nor U4005 (N_4005,N_3281,N_3319);
nor U4006 (N_4006,N_3769,N_3434);
nor U4007 (N_4007,N_3128,N_3617);
nor U4008 (N_4008,N_3049,N_3875);
or U4009 (N_4009,N_3857,N_3698);
nor U4010 (N_4010,N_3094,N_3076);
and U4011 (N_4011,N_3750,N_3089);
and U4012 (N_4012,N_3370,N_3057);
nor U4013 (N_4013,N_3347,N_3705);
nand U4014 (N_4014,N_3313,N_3763);
or U4015 (N_4015,N_3299,N_3568);
nor U4016 (N_4016,N_3213,N_3001);
and U4017 (N_4017,N_3247,N_3258);
nand U4018 (N_4018,N_3235,N_3039);
nor U4019 (N_4019,N_3598,N_3367);
nor U4020 (N_4020,N_3563,N_3808);
and U4021 (N_4021,N_3083,N_3713);
and U4022 (N_4022,N_3834,N_3318);
nand U4023 (N_4023,N_3623,N_3830);
nor U4024 (N_4024,N_3664,N_3594);
and U4025 (N_4025,N_3788,N_3900);
nand U4026 (N_4026,N_3804,N_3382);
nor U4027 (N_4027,N_3245,N_3234);
or U4028 (N_4028,N_3754,N_3154);
or U4029 (N_4029,N_3835,N_3937);
nor U4030 (N_4030,N_3656,N_3183);
or U4031 (N_4031,N_3114,N_3841);
or U4032 (N_4032,N_3936,N_3351);
or U4033 (N_4033,N_3519,N_3322);
and U4034 (N_4034,N_3181,N_3504);
nand U4035 (N_4035,N_3155,N_3574);
or U4036 (N_4036,N_3681,N_3759);
nor U4037 (N_4037,N_3944,N_3931);
and U4038 (N_4038,N_3659,N_3696);
and U4039 (N_4039,N_3473,N_3206);
or U4040 (N_4040,N_3606,N_3184);
and U4041 (N_4041,N_3468,N_3325);
and U4042 (N_4042,N_3220,N_3477);
or U4043 (N_4043,N_3671,N_3978);
and U4044 (N_4044,N_3774,N_3676);
or U4045 (N_4045,N_3356,N_3328);
nor U4046 (N_4046,N_3558,N_3193);
nand U4047 (N_4047,N_3239,N_3605);
nand U4048 (N_4048,N_3077,N_3670);
and U4049 (N_4049,N_3003,N_3876);
or U4050 (N_4050,N_3555,N_3257);
and U4051 (N_4051,N_3324,N_3962);
nand U4052 (N_4052,N_3216,N_3161);
nor U4053 (N_4053,N_3253,N_3663);
nor U4054 (N_4054,N_3631,N_3567);
nor U4055 (N_4055,N_3217,N_3095);
nand U4056 (N_4056,N_3715,N_3772);
nand U4057 (N_4057,N_3514,N_3585);
nor U4058 (N_4058,N_3126,N_3593);
and U4059 (N_4059,N_3811,N_3453);
nand U4060 (N_4060,N_3815,N_3259);
or U4061 (N_4061,N_3334,N_3645);
nor U4062 (N_4062,N_3959,N_3188);
xor U4063 (N_4063,N_3037,N_3162);
nand U4064 (N_4064,N_3901,N_3544);
nand U4065 (N_4065,N_3203,N_3792);
and U4066 (N_4066,N_3789,N_3982);
and U4067 (N_4067,N_3165,N_3355);
or U4068 (N_4068,N_3046,N_3443);
or U4069 (N_4069,N_3595,N_3907);
or U4070 (N_4070,N_3930,N_3706);
nor U4071 (N_4071,N_3127,N_3465);
and U4072 (N_4072,N_3752,N_3524);
nor U4073 (N_4073,N_3892,N_3158);
and U4074 (N_4074,N_3784,N_3411);
or U4075 (N_4075,N_3724,N_3485);
nand U4076 (N_4076,N_3899,N_3994);
nor U4077 (N_4077,N_3886,N_3391);
and U4078 (N_4078,N_3932,N_3949);
nand U4079 (N_4079,N_3358,N_3496);
nor U4080 (N_4080,N_3837,N_3960);
nor U4081 (N_4081,N_3734,N_3480);
or U4082 (N_4082,N_3372,N_3662);
nor U4083 (N_4083,N_3934,N_3539);
nor U4084 (N_4084,N_3674,N_3588);
or U4085 (N_4085,N_3753,N_3080);
nand U4086 (N_4086,N_3580,N_3343);
nand U4087 (N_4087,N_3445,N_3433);
nor U4088 (N_4088,N_3349,N_3371);
and U4089 (N_4089,N_3646,N_3228);
and U4090 (N_4090,N_3614,N_3885);
nand U4091 (N_4091,N_3836,N_3726);
nand U4092 (N_4092,N_3723,N_3529);
and U4093 (N_4093,N_3787,N_3208);
and U4094 (N_4094,N_3133,N_3141);
nand U4095 (N_4095,N_3736,N_3346);
or U4096 (N_4096,N_3252,N_3817);
or U4097 (N_4097,N_3357,N_3483);
or U4098 (N_4098,N_3063,N_3913);
and U4099 (N_4099,N_3010,N_3416);
nand U4100 (N_4100,N_3112,N_3549);
nand U4101 (N_4101,N_3068,N_3441);
nand U4102 (N_4102,N_3502,N_3704);
and U4103 (N_4103,N_3897,N_3320);
and U4104 (N_4104,N_3831,N_3694);
and U4105 (N_4105,N_3178,N_3569);
nand U4106 (N_4106,N_3498,N_3148);
or U4107 (N_4107,N_3012,N_3398);
nand U4108 (N_4108,N_3725,N_3729);
and U4109 (N_4109,N_3047,N_3022);
and U4110 (N_4110,N_3442,N_3489);
nand U4111 (N_4111,N_3961,N_3909);
and U4112 (N_4112,N_3336,N_3028);
nand U4113 (N_4113,N_3300,N_3438);
nor U4114 (N_4114,N_3570,N_3056);
nand U4115 (N_4115,N_3030,N_3703);
nand U4116 (N_4116,N_3560,N_3180);
nor U4117 (N_4117,N_3616,N_3390);
nor U4118 (N_4118,N_3020,N_3854);
xor U4119 (N_4119,N_3065,N_3394);
nand U4120 (N_4120,N_3110,N_3535);
and U4121 (N_4121,N_3136,N_3501);
or U4122 (N_4122,N_3942,N_3840);
nand U4123 (N_4123,N_3634,N_3064);
and U4124 (N_4124,N_3261,N_3666);
nand U4125 (N_4125,N_3297,N_3655);
and U4126 (N_4126,N_3929,N_3693);
or U4127 (N_4127,N_3013,N_3098);
and U4128 (N_4128,N_3891,N_3805);
or U4129 (N_4129,N_3985,N_3244);
nor U4130 (N_4130,N_3768,N_3491);
nor U4131 (N_4131,N_3541,N_3345);
and U4132 (N_4132,N_3439,N_3517);
and U4133 (N_4133,N_3744,N_3669);
or U4134 (N_4134,N_3081,N_3939);
nand U4135 (N_4135,N_3249,N_3199);
and U4136 (N_4136,N_3632,N_3981);
nand U4137 (N_4137,N_3418,N_3458);
or U4138 (N_4138,N_3209,N_3414);
or U4139 (N_4139,N_3302,N_3627);
or U4140 (N_4140,N_3924,N_3509);
nand U4141 (N_4141,N_3791,N_3194);
or U4142 (N_4142,N_3896,N_3066);
nand U4143 (N_4143,N_3388,N_3229);
or U4144 (N_4144,N_3435,N_3866);
nand U4145 (N_4145,N_3849,N_3816);
and U4146 (N_4146,N_3182,N_3115);
and U4147 (N_4147,N_3254,N_3389);
nor U4148 (N_4148,N_3576,N_3147);
and U4149 (N_4149,N_3340,N_3137);
nand U4150 (N_4150,N_3255,N_3121);
and U4151 (N_4151,N_3971,N_3902);
and U4152 (N_4152,N_3448,N_3212);
nand U4153 (N_4153,N_3423,N_3649);
nand U4154 (N_4154,N_3888,N_3643);
and U4155 (N_4155,N_3469,N_3904);
and U4156 (N_4156,N_3305,N_3470);
or U4157 (N_4157,N_3903,N_3583);
and U4158 (N_4158,N_3451,N_3884);
nor U4159 (N_4159,N_3270,N_3820);
and U4160 (N_4160,N_3260,N_3461);
nor U4161 (N_4161,N_3809,N_3174);
nand U4162 (N_4162,N_3604,N_3758);
nand U4163 (N_4163,N_3230,N_3384);
or U4164 (N_4164,N_3187,N_3874);
nand U4165 (N_4165,N_3072,N_3051);
or U4166 (N_4166,N_3279,N_3550);
nand U4167 (N_4167,N_3185,N_3238);
nand U4168 (N_4168,N_3581,N_3843);
and U4169 (N_4169,N_3626,N_3457);
nand U4170 (N_4170,N_3419,N_3381);
or U4171 (N_4171,N_3586,N_3471);
nand U4172 (N_4172,N_3612,N_3553);
nor U4173 (N_4173,N_3027,N_3284);
nand U4174 (N_4174,N_3452,N_3906);
nor U4175 (N_4175,N_3677,N_3198);
nand U4176 (N_4176,N_3038,N_3100);
nor U4177 (N_4177,N_3017,N_3742);
nor U4178 (N_4178,N_3085,N_3740);
nand U4179 (N_4179,N_3506,N_3315);
or U4180 (N_4180,N_3149,N_3362);
nand U4181 (N_4181,N_3084,N_3999);
nor U4182 (N_4182,N_3379,N_3146);
and U4183 (N_4183,N_3945,N_3251);
and U4184 (N_4184,N_3309,N_3887);
and U4185 (N_4185,N_3968,N_3807);
and U4186 (N_4186,N_3425,N_3856);
nand U4187 (N_4187,N_3339,N_3404);
nor U4188 (N_4188,N_3877,N_3781);
nor U4189 (N_4189,N_3500,N_3380);
or U4190 (N_4190,N_3482,N_3168);
nand U4191 (N_4191,N_3396,N_3954);
nor U4192 (N_4192,N_3237,N_3973);
or U4193 (N_4193,N_3002,N_3823);
or U4194 (N_4194,N_3975,N_3033);
nor U4195 (N_4195,N_3926,N_3437);
and U4196 (N_4196,N_3720,N_3761);
nor U4197 (N_4197,N_3641,N_3354);
or U4198 (N_4198,N_3430,N_3974);
and U4199 (N_4199,N_3846,N_3803);
nor U4200 (N_4200,N_3977,N_3364);
nor U4201 (N_4201,N_3035,N_3546);
xnor U4202 (N_4202,N_3119,N_3782);
nor U4203 (N_4203,N_3352,N_3175);
nor U4204 (N_4204,N_3618,N_3475);
nand U4205 (N_4205,N_3658,N_3692);
and U4206 (N_4206,N_3839,N_3608);
nand U4207 (N_4207,N_3403,N_3218);
nand U4208 (N_4208,N_3310,N_3344);
or U4209 (N_4209,N_3493,N_3861);
nor U4210 (N_4210,N_3847,N_3104);
nor U4211 (N_4211,N_3579,N_3474);
or U4212 (N_4212,N_3741,N_3086);
nor U4213 (N_4213,N_3824,N_3408);
and U4214 (N_4214,N_3620,N_3288);
or U4215 (N_4215,N_3368,N_3597);
or U4216 (N_4216,N_3997,N_3467);
or U4217 (N_4217,N_3554,N_3650);
xor U4218 (N_4218,N_3547,N_3917);
and U4219 (N_4219,N_3103,N_3409);
and U4220 (N_4220,N_3231,N_3045);
or U4221 (N_4221,N_3093,N_3116);
nor U4222 (N_4222,N_3842,N_3979);
nand U4223 (N_4223,N_3786,N_3635);
nor U4224 (N_4224,N_3599,N_3191);
nand U4225 (N_4225,N_3397,N_3138);
and U4226 (N_4226,N_3683,N_3195);
or U4227 (N_4227,N_3088,N_3428);
or U4228 (N_4228,N_3812,N_3505);
nand U4229 (N_4229,N_3348,N_3025);
nor U4230 (N_4230,N_3476,N_3628);
nand U4231 (N_4231,N_3523,N_3629);
nor U4232 (N_4232,N_3559,N_3156);
and U4233 (N_4233,N_3923,N_3177);
nand U4234 (N_4234,N_3879,N_3828);
or U4235 (N_4235,N_3431,N_3413);
or U4236 (N_4236,N_3893,N_3602);
nand U4237 (N_4237,N_3233,N_3853);
nand U4238 (N_4238,N_3201,N_3625);
nand U4239 (N_4239,N_3009,N_3240);
and U4240 (N_4240,N_3665,N_3611);
nor U4241 (N_4241,N_3950,N_3619);
nand U4242 (N_4242,N_3023,N_3459);
nor U4243 (N_4243,N_3813,N_3144);
or U4244 (N_4244,N_3283,N_3363);
and U4245 (N_4245,N_3711,N_3622);
and U4246 (N_4246,N_3532,N_3196);
nor U4247 (N_4247,N_3731,N_3296);
nand U4248 (N_4248,N_3415,N_3660);
or U4249 (N_4249,N_3798,N_3079);
or U4250 (N_4250,N_3911,N_3644);
nor U4251 (N_4251,N_3984,N_3207);
and U4252 (N_4252,N_3746,N_3243);
nor U4253 (N_4253,N_3624,N_3957);
and U4254 (N_4254,N_3822,N_3783);
nand U4255 (N_4255,N_3487,N_3832);
and U4256 (N_4256,N_3990,N_3205);
nor U4257 (N_4257,N_3702,N_3337);
or U4258 (N_4258,N_3735,N_3176);
nor U4259 (N_4259,N_3685,N_3745);
or U4260 (N_4260,N_3511,N_3508);
nor U4261 (N_4261,N_3918,N_3755);
nor U4262 (N_4262,N_3969,N_3298);
nor U4263 (N_4263,N_3044,N_3332);
and U4264 (N_4264,N_3169,N_3621);
and U4265 (N_4265,N_3091,N_3938);
or U4266 (N_4266,N_3738,N_3527);
nor U4267 (N_4267,N_3872,N_3436);
and U4268 (N_4268,N_3536,N_3914);
or U4269 (N_4269,N_3573,N_3881);
and U4270 (N_4270,N_3862,N_3818);
nand U4271 (N_4271,N_3190,N_3780);
nor U4272 (N_4272,N_3041,N_3680);
and U4273 (N_4273,N_3765,N_3531);
nand U4274 (N_4274,N_3087,N_3327);
or U4275 (N_4275,N_3272,N_3466);
nand U4276 (N_4276,N_3684,N_3402);
nor U4277 (N_4277,N_3572,N_3308);
or U4278 (N_4278,N_3312,N_3712);
nor U4279 (N_4279,N_3829,N_3360);
or U4280 (N_4280,N_3157,N_3654);
or U4281 (N_4281,N_3053,N_3970);
nor U4282 (N_4282,N_3189,N_3717);
or U4283 (N_4283,N_3778,N_3412);
nand U4284 (N_4284,N_3171,N_3225);
nor U4285 (N_4285,N_3099,N_3518);
nor U4286 (N_4286,N_3109,N_3290);
nor U4287 (N_4287,N_3743,N_3365);
or U4288 (N_4288,N_3905,N_3700);
or U4289 (N_4289,N_3967,N_3565);
or U4290 (N_4290,N_3395,N_3492);
nor U4291 (N_4291,N_3062,N_3444);
nand U4292 (N_4292,N_3152,N_3958);
nand U4293 (N_4293,N_3578,N_3739);
nand U4294 (N_4294,N_3951,N_3264);
and U4295 (N_4295,N_3941,N_3040);
nor U4296 (N_4296,N_3050,N_3749);
nor U4297 (N_4297,N_3728,N_3678);
or U4298 (N_4298,N_3271,N_3338);
nor U4299 (N_4299,N_3108,N_3266);
nor U4300 (N_4300,N_3202,N_3246);
and U4301 (N_4301,N_3280,N_3293);
nand U4302 (N_4302,N_3639,N_3779);
nor U4303 (N_4303,N_3564,N_3894);
nor U4304 (N_4304,N_3016,N_3718);
nand U4305 (N_4305,N_3852,N_3073);
xnor U4306 (N_4306,N_3150,N_3640);
and U4307 (N_4307,N_3802,N_3916);
and U4308 (N_4308,N_3186,N_3214);
and U4309 (N_4309,N_3799,N_3463);
and U4310 (N_4310,N_3167,N_3987);
nor U4311 (N_4311,N_3859,N_3661);
or U4312 (N_4312,N_3764,N_3067);
nor U4313 (N_4313,N_3691,N_3486);
and U4314 (N_4314,N_3701,N_3797);
nand U4315 (N_4315,N_3933,N_3256);
and U4316 (N_4316,N_3793,N_3719);
nor U4317 (N_4317,N_3908,N_3070);
or U4318 (N_4318,N_3131,N_3869);
nor U4319 (N_4319,N_3197,N_3771);
nor U4320 (N_4320,N_3946,N_3697);
nand U4321 (N_4321,N_3111,N_3392);
nand U4322 (N_4322,N_3587,N_3401);
and U4323 (N_4323,N_3575,N_3795);
and U4324 (N_4324,N_3610,N_3350);
nand U4325 (N_4325,N_3675,N_3601);
nor U4326 (N_4326,N_3335,N_3915);
or U4327 (N_4327,N_3928,N_3850);
nor U4328 (N_4328,N_3510,N_3285);
nor U4329 (N_4329,N_3316,N_3417);
and U4330 (N_4330,N_3732,N_3890);
nor U4331 (N_4331,N_3801,N_3034);
nor U4332 (N_4332,N_3454,N_3673);
and U4333 (N_4333,N_3562,N_3727);
nor U4334 (N_4334,N_3385,N_3838);
or U4335 (N_4335,N_3151,N_3052);
and U4336 (N_4336,N_3160,N_3375);
and U4337 (N_4337,N_3642,N_3455);
nor U4338 (N_4338,N_3232,N_3106);
nand U4339 (N_4339,N_3102,N_3988);
and U4340 (N_4340,N_3609,N_3263);
or U4341 (N_4341,N_3542,N_3690);
nand U4342 (N_4342,N_3140,N_3855);
or U4343 (N_4343,N_3353,N_3200);
and U4344 (N_4344,N_3007,N_3653);
and U4345 (N_4345,N_3015,N_3989);
nand U4346 (N_4346,N_3026,N_3329);
and U4347 (N_4347,N_3860,N_3163);
nand U4348 (N_4348,N_3992,N_3497);
nand U4349 (N_4349,N_3029,N_3777);
nor U4350 (N_4350,N_3577,N_3449);
nor U4351 (N_4351,N_3082,N_3943);
nor U4352 (N_4352,N_3326,N_3366);
nand U4353 (N_4353,N_3236,N_3827);
nand U4354 (N_4354,N_3596,N_3426);
and U4355 (N_4355,N_3014,N_3129);
nand U4356 (N_4356,N_3276,N_3868);
nor U4357 (N_4357,N_3770,N_3668);
xnor U4358 (N_4358,N_3361,N_3964);
or U4359 (N_4359,N_3166,N_3767);
or U4360 (N_4360,N_3748,N_3460);
or U4361 (N_4361,N_3224,N_3966);
nand U4362 (N_4362,N_3630,N_3273);
or U4363 (N_4363,N_3953,N_3311);
or U4364 (N_4364,N_3922,N_3582);
nand U4365 (N_4365,N_3494,N_3773);
nand U4366 (N_4366,N_3387,N_3421);
nand U4367 (N_4367,N_3775,N_3410);
nand U4368 (N_4368,N_3867,N_3386);
nand U4369 (N_4369,N_3672,N_3757);
and U4370 (N_4370,N_3242,N_3130);
nor U4371 (N_4371,N_3589,N_3277);
nor U4372 (N_4372,N_3870,N_3295);
nand U4373 (N_4373,N_3980,N_3330);
nand U4374 (N_4374,N_3709,N_3376);
nor U4375 (N_4375,N_3955,N_3543);
nor U4376 (N_4376,N_3525,N_3520);
nand U4377 (N_4377,N_3993,N_3399);
nor U4378 (N_4378,N_3464,N_3819);
or U4379 (N_4379,N_3566,N_3533);
and U4380 (N_4380,N_3018,N_3889);
or U4381 (N_4381,N_3507,N_3592);
nor U4382 (N_4382,N_3374,N_3733);
or U4383 (N_4383,N_3863,N_3873);
nor U4384 (N_4384,N_3250,N_3024);
nand U4385 (N_4385,N_3008,N_3210);
nor U4386 (N_4386,N_3307,N_3516);
nand U4387 (N_4387,N_3737,N_3006);
nand U4388 (N_4388,N_3341,N_3055);
nand U4389 (N_4389,N_3286,N_3895);
and U4390 (N_4390,N_3996,N_3695);
nand U4391 (N_4391,N_3882,N_3552);
and U4392 (N_4392,N_3306,N_3513);
and U4393 (N_4393,N_3107,N_3825);
or U4394 (N_4394,N_3688,N_3120);
nor U4395 (N_4395,N_3528,N_3032);
or U4396 (N_4396,N_3912,N_3682);
and U4397 (N_4397,N_3521,N_3383);
or U4398 (N_4398,N_3667,N_3534);
and U4399 (N_4399,N_3456,N_3059);
or U4400 (N_4400,N_3657,N_3021);
nor U4401 (N_4401,N_3490,N_3848);
nand U4402 (N_4402,N_3301,N_3090);
or U4403 (N_4403,N_3865,N_3429);
and U4404 (N_4404,N_3274,N_3548);
nor U4405 (N_4405,N_3800,N_3910);
nand U4406 (N_4406,N_3806,N_3603);
and U4407 (N_4407,N_3495,N_3031);
nor U4408 (N_4408,N_3481,N_3686);
nand U4409 (N_4409,N_3078,N_3556);
or U4410 (N_4410,N_3648,N_3651);
and U4411 (N_4411,N_3192,N_3406);
nand U4412 (N_4412,N_3113,N_3400);
nand U4413 (N_4413,N_3998,N_3794);
nor U4414 (N_4414,N_3074,N_3935);
or U4415 (N_4415,N_3143,N_3551);
or U4416 (N_4416,N_3420,N_3215);
and U4417 (N_4417,N_3226,N_3515);
or U4418 (N_4418,N_3153,N_3241);
nor U4419 (N_4419,N_3048,N_3730);
and U4420 (N_4420,N_3584,N_3275);
nand U4421 (N_4421,N_3135,N_3976);
or U4422 (N_4422,N_3118,N_3139);
or U4423 (N_4423,N_3826,N_3092);
nand U4424 (N_4424,N_3446,N_3219);
and U4425 (N_4425,N_3995,N_3845);
and U4426 (N_4426,N_3919,N_3561);
nor U4427 (N_4427,N_3972,N_3132);
and U4428 (N_4428,N_3125,N_3637);
or U4429 (N_4429,N_3814,N_3488);
and U4430 (N_4430,N_3097,N_3880);
nor U4431 (N_4431,N_3019,N_3359);
and U4432 (N_4432,N_3145,N_3462);
nor U4433 (N_4433,N_3921,N_3883);
nor U4434 (N_4434,N_3687,N_3607);
nand U4435 (N_4435,N_3304,N_3499);
nor U4436 (N_4436,N_3289,N_3940);
or U4437 (N_4437,N_3878,N_3833);
nand U4438 (N_4438,N_3096,N_3638);
or U4439 (N_4439,N_3407,N_3075);
or U4440 (N_4440,N_3537,N_3751);
and U4441 (N_4441,N_3714,N_3790);
nand U4442 (N_4442,N_3042,N_3378);
nand U4443 (N_4443,N_3269,N_3716);
or U4444 (N_4444,N_3858,N_3333);
nor U4445 (N_4445,N_3265,N_3927);
nand U4446 (N_4446,N_3054,N_3267);
and U4447 (N_4447,N_3221,N_3538);
and U4448 (N_4448,N_3294,N_3952);
and U4449 (N_4449,N_3991,N_3821);
nand U4450 (N_4450,N_3179,N_3004);
xor U4451 (N_4451,N_3011,N_3472);
nor U4452 (N_4452,N_3963,N_3613);
nor U4453 (N_4453,N_3422,N_3314);
nand U4454 (N_4454,N_3965,N_3785);
and U4455 (N_4455,N_3211,N_3331);
nor U4456 (N_4456,N_3282,N_3699);
nand U4457 (N_4457,N_3321,N_3503);
nor U4458 (N_4458,N_3287,N_3036);
nand U4459 (N_4459,N_3871,N_3707);
and U4460 (N_4460,N_3373,N_3636);
or U4461 (N_4461,N_3000,N_3440);
nor U4462 (N_4462,N_3920,N_3557);
and U4463 (N_4463,N_3134,N_3142);
or U4464 (N_4464,N_3061,N_3545);
or U4465 (N_4465,N_3721,N_3173);
nor U4466 (N_4466,N_3647,N_3123);
nor U4467 (N_4467,N_3591,N_3722);
nand U4468 (N_4468,N_3484,N_3747);
or U4469 (N_4469,N_3776,N_3268);
or U4470 (N_4470,N_3124,N_3058);
and U4471 (N_4471,N_3710,N_3071);
or U4472 (N_4472,N_3323,N_3986);
or U4473 (N_4473,N_3530,N_3060);
nand U4474 (N_4474,N_3948,N_3956);
or U4475 (N_4475,N_3405,N_3864);
or U4476 (N_4476,N_3278,N_3222);
nor U4477 (N_4477,N_3043,N_3633);
or U4478 (N_4478,N_3925,N_3172);
nand U4479 (N_4479,N_3615,N_3652);
or U4480 (N_4480,N_3571,N_3424);
nor U4481 (N_4481,N_3369,N_3600);
and U4482 (N_4482,N_3227,N_3159);
and U4483 (N_4483,N_3760,N_3291);
nand U4484 (N_4484,N_3101,N_3689);
nand U4485 (N_4485,N_3947,N_3248);
nand U4486 (N_4486,N_3117,N_3796);
nor U4487 (N_4487,N_3292,N_3204);
or U4488 (N_4488,N_3447,N_3105);
nor U4489 (N_4489,N_3679,N_3512);
and U4490 (N_4490,N_3590,N_3005);
nor U4491 (N_4491,N_3450,N_3377);
or U4492 (N_4492,N_3844,N_3262);
nand U4493 (N_4493,N_3393,N_3766);
and U4494 (N_4494,N_3708,N_3540);
nand U4495 (N_4495,N_3898,N_3342);
nor U4496 (N_4496,N_3526,N_3478);
nor U4497 (N_4497,N_3810,N_3164);
and U4498 (N_4498,N_3522,N_3756);
or U4499 (N_4499,N_3983,N_3432);
nand U4500 (N_4500,N_3729,N_3739);
and U4501 (N_4501,N_3417,N_3797);
nor U4502 (N_4502,N_3588,N_3458);
and U4503 (N_4503,N_3263,N_3532);
and U4504 (N_4504,N_3127,N_3441);
nand U4505 (N_4505,N_3532,N_3186);
and U4506 (N_4506,N_3865,N_3489);
or U4507 (N_4507,N_3959,N_3767);
nor U4508 (N_4508,N_3382,N_3826);
or U4509 (N_4509,N_3881,N_3814);
nand U4510 (N_4510,N_3813,N_3228);
nand U4511 (N_4511,N_3424,N_3696);
nor U4512 (N_4512,N_3488,N_3449);
xor U4513 (N_4513,N_3402,N_3823);
or U4514 (N_4514,N_3250,N_3287);
and U4515 (N_4515,N_3437,N_3190);
nor U4516 (N_4516,N_3104,N_3572);
or U4517 (N_4517,N_3769,N_3734);
or U4518 (N_4518,N_3713,N_3506);
or U4519 (N_4519,N_3431,N_3191);
or U4520 (N_4520,N_3222,N_3973);
or U4521 (N_4521,N_3060,N_3933);
or U4522 (N_4522,N_3978,N_3879);
and U4523 (N_4523,N_3036,N_3871);
nor U4524 (N_4524,N_3544,N_3004);
xor U4525 (N_4525,N_3652,N_3167);
nor U4526 (N_4526,N_3437,N_3013);
nand U4527 (N_4527,N_3082,N_3100);
nand U4528 (N_4528,N_3041,N_3982);
and U4529 (N_4529,N_3010,N_3969);
nand U4530 (N_4530,N_3845,N_3152);
nor U4531 (N_4531,N_3788,N_3312);
nand U4532 (N_4532,N_3634,N_3676);
and U4533 (N_4533,N_3164,N_3502);
nand U4534 (N_4534,N_3604,N_3575);
or U4535 (N_4535,N_3274,N_3022);
nand U4536 (N_4536,N_3220,N_3608);
and U4537 (N_4537,N_3424,N_3067);
or U4538 (N_4538,N_3399,N_3459);
nor U4539 (N_4539,N_3635,N_3103);
nor U4540 (N_4540,N_3289,N_3017);
nor U4541 (N_4541,N_3638,N_3994);
or U4542 (N_4542,N_3831,N_3504);
nor U4543 (N_4543,N_3066,N_3580);
nand U4544 (N_4544,N_3419,N_3119);
nand U4545 (N_4545,N_3653,N_3528);
and U4546 (N_4546,N_3082,N_3382);
or U4547 (N_4547,N_3900,N_3086);
and U4548 (N_4548,N_3922,N_3045);
or U4549 (N_4549,N_3496,N_3964);
and U4550 (N_4550,N_3689,N_3516);
nand U4551 (N_4551,N_3780,N_3493);
and U4552 (N_4552,N_3247,N_3823);
or U4553 (N_4553,N_3438,N_3558);
nand U4554 (N_4554,N_3680,N_3157);
nand U4555 (N_4555,N_3206,N_3502);
and U4556 (N_4556,N_3441,N_3782);
and U4557 (N_4557,N_3682,N_3259);
nor U4558 (N_4558,N_3669,N_3260);
nor U4559 (N_4559,N_3881,N_3119);
or U4560 (N_4560,N_3919,N_3249);
nand U4561 (N_4561,N_3091,N_3537);
or U4562 (N_4562,N_3263,N_3505);
nand U4563 (N_4563,N_3179,N_3079);
or U4564 (N_4564,N_3435,N_3888);
or U4565 (N_4565,N_3953,N_3407);
or U4566 (N_4566,N_3170,N_3278);
nor U4567 (N_4567,N_3161,N_3693);
nor U4568 (N_4568,N_3383,N_3328);
nand U4569 (N_4569,N_3221,N_3451);
or U4570 (N_4570,N_3037,N_3801);
and U4571 (N_4571,N_3333,N_3577);
nand U4572 (N_4572,N_3503,N_3097);
and U4573 (N_4573,N_3201,N_3135);
nor U4574 (N_4574,N_3415,N_3569);
nand U4575 (N_4575,N_3084,N_3285);
nand U4576 (N_4576,N_3021,N_3755);
nor U4577 (N_4577,N_3880,N_3231);
and U4578 (N_4578,N_3517,N_3266);
nand U4579 (N_4579,N_3232,N_3365);
or U4580 (N_4580,N_3768,N_3761);
or U4581 (N_4581,N_3255,N_3754);
and U4582 (N_4582,N_3688,N_3667);
xnor U4583 (N_4583,N_3069,N_3115);
nand U4584 (N_4584,N_3772,N_3158);
or U4585 (N_4585,N_3711,N_3837);
nand U4586 (N_4586,N_3331,N_3882);
or U4587 (N_4587,N_3216,N_3132);
nor U4588 (N_4588,N_3857,N_3783);
or U4589 (N_4589,N_3938,N_3373);
nand U4590 (N_4590,N_3808,N_3421);
xnor U4591 (N_4591,N_3164,N_3186);
or U4592 (N_4592,N_3561,N_3548);
or U4593 (N_4593,N_3498,N_3881);
and U4594 (N_4594,N_3691,N_3656);
or U4595 (N_4595,N_3929,N_3718);
nor U4596 (N_4596,N_3369,N_3760);
nand U4597 (N_4597,N_3766,N_3493);
and U4598 (N_4598,N_3876,N_3675);
or U4599 (N_4599,N_3559,N_3235);
and U4600 (N_4600,N_3379,N_3198);
xor U4601 (N_4601,N_3337,N_3199);
nor U4602 (N_4602,N_3403,N_3168);
or U4603 (N_4603,N_3650,N_3698);
nand U4604 (N_4604,N_3488,N_3028);
nand U4605 (N_4605,N_3125,N_3803);
and U4606 (N_4606,N_3282,N_3499);
nand U4607 (N_4607,N_3019,N_3805);
nor U4608 (N_4608,N_3005,N_3069);
and U4609 (N_4609,N_3228,N_3103);
or U4610 (N_4610,N_3607,N_3968);
and U4611 (N_4611,N_3267,N_3701);
or U4612 (N_4612,N_3286,N_3389);
and U4613 (N_4613,N_3515,N_3057);
nor U4614 (N_4614,N_3576,N_3817);
and U4615 (N_4615,N_3026,N_3553);
or U4616 (N_4616,N_3667,N_3205);
nor U4617 (N_4617,N_3083,N_3220);
and U4618 (N_4618,N_3587,N_3450);
nand U4619 (N_4619,N_3462,N_3596);
nand U4620 (N_4620,N_3653,N_3011);
or U4621 (N_4621,N_3925,N_3931);
or U4622 (N_4622,N_3651,N_3833);
or U4623 (N_4623,N_3212,N_3372);
and U4624 (N_4624,N_3278,N_3335);
and U4625 (N_4625,N_3274,N_3012);
or U4626 (N_4626,N_3039,N_3719);
and U4627 (N_4627,N_3278,N_3495);
nor U4628 (N_4628,N_3720,N_3861);
nor U4629 (N_4629,N_3891,N_3401);
and U4630 (N_4630,N_3638,N_3348);
or U4631 (N_4631,N_3066,N_3803);
or U4632 (N_4632,N_3172,N_3732);
xor U4633 (N_4633,N_3033,N_3427);
nand U4634 (N_4634,N_3539,N_3162);
nor U4635 (N_4635,N_3278,N_3839);
nor U4636 (N_4636,N_3295,N_3807);
and U4637 (N_4637,N_3697,N_3113);
or U4638 (N_4638,N_3647,N_3498);
or U4639 (N_4639,N_3839,N_3075);
or U4640 (N_4640,N_3382,N_3945);
nand U4641 (N_4641,N_3164,N_3045);
nor U4642 (N_4642,N_3379,N_3114);
nor U4643 (N_4643,N_3252,N_3692);
nand U4644 (N_4644,N_3305,N_3533);
and U4645 (N_4645,N_3233,N_3542);
nor U4646 (N_4646,N_3929,N_3924);
or U4647 (N_4647,N_3510,N_3484);
and U4648 (N_4648,N_3591,N_3322);
and U4649 (N_4649,N_3282,N_3675);
nor U4650 (N_4650,N_3229,N_3246);
nor U4651 (N_4651,N_3661,N_3326);
nand U4652 (N_4652,N_3428,N_3398);
nor U4653 (N_4653,N_3884,N_3571);
nand U4654 (N_4654,N_3820,N_3960);
or U4655 (N_4655,N_3265,N_3194);
or U4656 (N_4656,N_3219,N_3827);
or U4657 (N_4657,N_3188,N_3293);
nor U4658 (N_4658,N_3483,N_3621);
and U4659 (N_4659,N_3926,N_3297);
nor U4660 (N_4660,N_3589,N_3342);
nand U4661 (N_4661,N_3995,N_3323);
and U4662 (N_4662,N_3504,N_3080);
nor U4663 (N_4663,N_3586,N_3955);
and U4664 (N_4664,N_3606,N_3093);
nand U4665 (N_4665,N_3722,N_3342);
and U4666 (N_4666,N_3185,N_3886);
and U4667 (N_4667,N_3438,N_3835);
or U4668 (N_4668,N_3815,N_3237);
or U4669 (N_4669,N_3410,N_3643);
nand U4670 (N_4670,N_3633,N_3585);
and U4671 (N_4671,N_3848,N_3319);
and U4672 (N_4672,N_3698,N_3803);
and U4673 (N_4673,N_3521,N_3569);
nand U4674 (N_4674,N_3564,N_3031);
nand U4675 (N_4675,N_3133,N_3361);
and U4676 (N_4676,N_3963,N_3606);
or U4677 (N_4677,N_3025,N_3938);
nand U4678 (N_4678,N_3921,N_3276);
nand U4679 (N_4679,N_3216,N_3583);
nand U4680 (N_4680,N_3777,N_3898);
nor U4681 (N_4681,N_3377,N_3511);
nor U4682 (N_4682,N_3054,N_3645);
and U4683 (N_4683,N_3129,N_3130);
xnor U4684 (N_4684,N_3225,N_3360);
nand U4685 (N_4685,N_3642,N_3292);
and U4686 (N_4686,N_3267,N_3941);
nand U4687 (N_4687,N_3654,N_3592);
or U4688 (N_4688,N_3140,N_3239);
nor U4689 (N_4689,N_3890,N_3645);
nor U4690 (N_4690,N_3626,N_3833);
and U4691 (N_4691,N_3203,N_3544);
or U4692 (N_4692,N_3550,N_3777);
nand U4693 (N_4693,N_3562,N_3306);
and U4694 (N_4694,N_3197,N_3723);
and U4695 (N_4695,N_3451,N_3689);
nand U4696 (N_4696,N_3840,N_3789);
and U4697 (N_4697,N_3021,N_3350);
nor U4698 (N_4698,N_3138,N_3443);
or U4699 (N_4699,N_3276,N_3097);
or U4700 (N_4700,N_3953,N_3864);
nand U4701 (N_4701,N_3220,N_3612);
and U4702 (N_4702,N_3028,N_3403);
nand U4703 (N_4703,N_3822,N_3937);
nand U4704 (N_4704,N_3862,N_3640);
nand U4705 (N_4705,N_3538,N_3623);
nor U4706 (N_4706,N_3739,N_3095);
nand U4707 (N_4707,N_3271,N_3019);
or U4708 (N_4708,N_3837,N_3212);
and U4709 (N_4709,N_3731,N_3598);
nor U4710 (N_4710,N_3868,N_3989);
nor U4711 (N_4711,N_3605,N_3891);
and U4712 (N_4712,N_3929,N_3118);
and U4713 (N_4713,N_3695,N_3722);
and U4714 (N_4714,N_3228,N_3183);
nor U4715 (N_4715,N_3146,N_3983);
nand U4716 (N_4716,N_3277,N_3415);
and U4717 (N_4717,N_3225,N_3123);
and U4718 (N_4718,N_3044,N_3394);
nor U4719 (N_4719,N_3419,N_3952);
nor U4720 (N_4720,N_3756,N_3420);
and U4721 (N_4721,N_3248,N_3873);
and U4722 (N_4722,N_3557,N_3380);
or U4723 (N_4723,N_3938,N_3155);
and U4724 (N_4724,N_3126,N_3432);
nor U4725 (N_4725,N_3587,N_3419);
and U4726 (N_4726,N_3490,N_3680);
and U4727 (N_4727,N_3368,N_3413);
nor U4728 (N_4728,N_3643,N_3365);
or U4729 (N_4729,N_3944,N_3825);
nand U4730 (N_4730,N_3345,N_3680);
and U4731 (N_4731,N_3667,N_3374);
and U4732 (N_4732,N_3192,N_3946);
and U4733 (N_4733,N_3048,N_3940);
or U4734 (N_4734,N_3110,N_3534);
and U4735 (N_4735,N_3704,N_3449);
nor U4736 (N_4736,N_3714,N_3282);
or U4737 (N_4737,N_3629,N_3498);
nor U4738 (N_4738,N_3568,N_3762);
nor U4739 (N_4739,N_3659,N_3926);
or U4740 (N_4740,N_3456,N_3967);
nand U4741 (N_4741,N_3862,N_3249);
and U4742 (N_4742,N_3729,N_3169);
nand U4743 (N_4743,N_3374,N_3255);
nor U4744 (N_4744,N_3116,N_3728);
nand U4745 (N_4745,N_3256,N_3686);
and U4746 (N_4746,N_3112,N_3068);
nor U4747 (N_4747,N_3371,N_3960);
or U4748 (N_4748,N_3302,N_3253);
and U4749 (N_4749,N_3007,N_3065);
or U4750 (N_4750,N_3820,N_3564);
nand U4751 (N_4751,N_3488,N_3738);
nand U4752 (N_4752,N_3486,N_3045);
or U4753 (N_4753,N_3744,N_3504);
nand U4754 (N_4754,N_3111,N_3233);
and U4755 (N_4755,N_3462,N_3473);
and U4756 (N_4756,N_3701,N_3865);
or U4757 (N_4757,N_3911,N_3569);
nand U4758 (N_4758,N_3338,N_3004);
and U4759 (N_4759,N_3895,N_3605);
and U4760 (N_4760,N_3167,N_3835);
nand U4761 (N_4761,N_3291,N_3926);
or U4762 (N_4762,N_3899,N_3457);
nand U4763 (N_4763,N_3685,N_3963);
and U4764 (N_4764,N_3389,N_3369);
nand U4765 (N_4765,N_3221,N_3704);
nand U4766 (N_4766,N_3702,N_3959);
or U4767 (N_4767,N_3506,N_3967);
or U4768 (N_4768,N_3815,N_3369);
nor U4769 (N_4769,N_3303,N_3431);
or U4770 (N_4770,N_3440,N_3768);
and U4771 (N_4771,N_3022,N_3508);
and U4772 (N_4772,N_3141,N_3577);
and U4773 (N_4773,N_3196,N_3065);
nand U4774 (N_4774,N_3173,N_3386);
or U4775 (N_4775,N_3135,N_3615);
nand U4776 (N_4776,N_3041,N_3587);
nand U4777 (N_4777,N_3011,N_3971);
or U4778 (N_4778,N_3633,N_3852);
nor U4779 (N_4779,N_3327,N_3105);
nor U4780 (N_4780,N_3015,N_3780);
and U4781 (N_4781,N_3576,N_3245);
nand U4782 (N_4782,N_3839,N_3399);
nand U4783 (N_4783,N_3132,N_3924);
and U4784 (N_4784,N_3874,N_3843);
nand U4785 (N_4785,N_3115,N_3477);
or U4786 (N_4786,N_3813,N_3651);
nor U4787 (N_4787,N_3998,N_3191);
nand U4788 (N_4788,N_3153,N_3985);
nand U4789 (N_4789,N_3011,N_3066);
and U4790 (N_4790,N_3108,N_3092);
or U4791 (N_4791,N_3377,N_3421);
or U4792 (N_4792,N_3385,N_3851);
and U4793 (N_4793,N_3241,N_3148);
and U4794 (N_4794,N_3924,N_3562);
xor U4795 (N_4795,N_3290,N_3881);
nand U4796 (N_4796,N_3614,N_3851);
nand U4797 (N_4797,N_3132,N_3011);
or U4798 (N_4798,N_3935,N_3653);
nand U4799 (N_4799,N_3217,N_3156);
nand U4800 (N_4800,N_3754,N_3550);
and U4801 (N_4801,N_3064,N_3971);
nor U4802 (N_4802,N_3137,N_3711);
nor U4803 (N_4803,N_3578,N_3636);
nor U4804 (N_4804,N_3183,N_3919);
nor U4805 (N_4805,N_3669,N_3568);
or U4806 (N_4806,N_3624,N_3356);
nor U4807 (N_4807,N_3445,N_3199);
nand U4808 (N_4808,N_3166,N_3535);
nand U4809 (N_4809,N_3481,N_3417);
nand U4810 (N_4810,N_3038,N_3612);
and U4811 (N_4811,N_3585,N_3979);
nor U4812 (N_4812,N_3722,N_3176);
and U4813 (N_4813,N_3337,N_3419);
or U4814 (N_4814,N_3017,N_3540);
and U4815 (N_4815,N_3915,N_3688);
and U4816 (N_4816,N_3928,N_3147);
nor U4817 (N_4817,N_3262,N_3258);
or U4818 (N_4818,N_3270,N_3383);
nand U4819 (N_4819,N_3016,N_3832);
nand U4820 (N_4820,N_3202,N_3494);
or U4821 (N_4821,N_3536,N_3671);
nor U4822 (N_4822,N_3532,N_3158);
or U4823 (N_4823,N_3147,N_3986);
or U4824 (N_4824,N_3081,N_3472);
nor U4825 (N_4825,N_3048,N_3568);
and U4826 (N_4826,N_3883,N_3215);
nand U4827 (N_4827,N_3699,N_3451);
or U4828 (N_4828,N_3086,N_3051);
nor U4829 (N_4829,N_3951,N_3481);
nand U4830 (N_4830,N_3463,N_3083);
nand U4831 (N_4831,N_3738,N_3433);
and U4832 (N_4832,N_3984,N_3452);
nand U4833 (N_4833,N_3970,N_3674);
nor U4834 (N_4834,N_3658,N_3731);
or U4835 (N_4835,N_3879,N_3213);
nand U4836 (N_4836,N_3905,N_3617);
or U4837 (N_4837,N_3592,N_3704);
or U4838 (N_4838,N_3524,N_3582);
nand U4839 (N_4839,N_3352,N_3745);
nor U4840 (N_4840,N_3622,N_3814);
or U4841 (N_4841,N_3799,N_3390);
and U4842 (N_4842,N_3400,N_3635);
nand U4843 (N_4843,N_3510,N_3453);
or U4844 (N_4844,N_3106,N_3370);
or U4845 (N_4845,N_3891,N_3698);
and U4846 (N_4846,N_3586,N_3957);
or U4847 (N_4847,N_3505,N_3198);
nand U4848 (N_4848,N_3935,N_3081);
nand U4849 (N_4849,N_3811,N_3101);
nand U4850 (N_4850,N_3669,N_3178);
nand U4851 (N_4851,N_3044,N_3347);
and U4852 (N_4852,N_3988,N_3692);
and U4853 (N_4853,N_3591,N_3605);
nand U4854 (N_4854,N_3478,N_3132);
and U4855 (N_4855,N_3998,N_3335);
and U4856 (N_4856,N_3771,N_3765);
nor U4857 (N_4857,N_3848,N_3112);
and U4858 (N_4858,N_3102,N_3190);
and U4859 (N_4859,N_3817,N_3277);
nand U4860 (N_4860,N_3403,N_3956);
xor U4861 (N_4861,N_3049,N_3086);
and U4862 (N_4862,N_3525,N_3933);
nor U4863 (N_4863,N_3652,N_3749);
or U4864 (N_4864,N_3256,N_3862);
or U4865 (N_4865,N_3799,N_3215);
and U4866 (N_4866,N_3889,N_3555);
nand U4867 (N_4867,N_3976,N_3233);
and U4868 (N_4868,N_3829,N_3986);
and U4869 (N_4869,N_3871,N_3513);
nor U4870 (N_4870,N_3323,N_3773);
nand U4871 (N_4871,N_3030,N_3904);
nor U4872 (N_4872,N_3929,N_3291);
and U4873 (N_4873,N_3975,N_3769);
and U4874 (N_4874,N_3445,N_3274);
or U4875 (N_4875,N_3471,N_3223);
nand U4876 (N_4876,N_3042,N_3235);
nor U4877 (N_4877,N_3339,N_3388);
and U4878 (N_4878,N_3630,N_3675);
or U4879 (N_4879,N_3244,N_3834);
nand U4880 (N_4880,N_3690,N_3108);
nor U4881 (N_4881,N_3583,N_3379);
or U4882 (N_4882,N_3674,N_3719);
or U4883 (N_4883,N_3526,N_3179);
nand U4884 (N_4884,N_3350,N_3418);
and U4885 (N_4885,N_3261,N_3365);
nand U4886 (N_4886,N_3217,N_3803);
and U4887 (N_4887,N_3955,N_3002);
nand U4888 (N_4888,N_3350,N_3172);
nand U4889 (N_4889,N_3843,N_3290);
and U4890 (N_4890,N_3927,N_3612);
and U4891 (N_4891,N_3273,N_3070);
or U4892 (N_4892,N_3226,N_3002);
nor U4893 (N_4893,N_3267,N_3432);
and U4894 (N_4894,N_3330,N_3536);
nor U4895 (N_4895,N_3881,N_3295);
nor U4896 (N_4896,N_3176,N_3524);
nand U4897 (N_4897,N_3802,N_3829);
nor U4898 (N_4898,N_3512,N_3839);
or U4899 (N_4899,N_3620,N_3038);
nor U4900 (N_4900,N_3105,N_3302);
and U4901 (N_4901,N_3210,N_3433);
and U4902 (N_4902,N_3403,N_3823);
or U4903 (N_4903,N_3564,N_3228);
or U4904 (N_4904,N_3650,N_3131);
or U4905 (N_4905,N_3919,N_3870);
or U4906 (N_4906,N_3827,N_3925);
and U4907 (N_4907,N_3480,N_3617);
or U4908 (N_4908,N_3226,N_3263);
or U4909 (N_4909,N_3875,N_3711);
nand U4910 (N_4910,N_3717,N_3679);
and U4911 (N_4911,N_3249,N_3874);
and U4912 (N_4912,N_3354,N_3842);
xor U4913 (N_4913,N_3437,N_3925);
and U4914 (N_4914,N_3593,N_3260);
nand U4915 (N_4915,N_3067,N_3546);
or U4916 (N_4916,N_3057,N_3651);
nor U4917 (N_4917,N_3889,N_3216);
nand U4918 (N_4918,N_3619,N_3587);
nand U4919 (N_4919,N_3120,N_3256);
or U4920 (N_4920,N_3416,N_3013);
nand U4921 (N_4921,N_3296,N_3697);
and U4922 (N_4922,N_3353,N_3402);
nand U4923 (N_4923,N_3097,N_3838);
nand U4924 (N_4924,N_3342,N_3852);
nand U4925 (N_4925,N_3216,N_3104);
nor U4926 (N_4926,N_3822,N_3895);
or U4927 (N_4927,N_3570,N_3106);
nand U4928 (N_4928,N_3607,N_3569);
or U4929 (N_4929,N_3227,N_3285);
and U4930 (N_4930,N_3859,N_3464);
and U4931 (N_4931,N_3103,N_3759);
nand U4932 (N_4932,N_3724,N_3248);
or U4933 (N_4933,N_3793,N_3589);
and U4934 (N_4934,N_3023,N_3183);
or U4935 (N_4935,N_3934,N_3951);
and U4936 (N_4936,N_3034,N_3833);
and U4937 (N_4937,N_3593,N_3606);
nor U4938 (N_4938,N_3409,N_3697);
and U4939 (N_4939,N_3006,N_3785);
or U4940 (N_4940,N_3323,N_3255);
nand U4941 (N_4941,N_3065,N_3515);
and U4942 (N_4942,N_3288,N_3417);
nand U4943 (N_4943,N_3174,N_3880);
or U4944 (N_4944,N_3897,N_3333);
nor U4945 (N_4945,N_3661,N_3261);
nand U4946 (N_4946,N_3209,N_3831);
nand U4947 (N_4947,N_3264,N_3048);
nand U4948 (N_4948,N_3599,N_3633);
and U4949 (N_4949,N_3469,N_3269);
or U4950 (N_4950,N_3773,N_3163);
nor U4951 (N_4951,N_3712,N_3504);
or U4952 (N_4952,N_3128,N_3301);
or U4953 (N_4953,N_3750,N_3230);
nor U4954 (N_4954,N_3109,N_3207);
nand U4955 (N_4955,N_3649,N_3138);
xor U4956 (N_4956,N_3250,N_3145);
nor U4957 (N_4957,N_3436,N_3723);
nor U4958 (N_4958,N_3328,N_3734);
and U4959 (N_4959,N_3716,N_3215);
and U4960 (N_4960,N_3594,N_3331);
nand U4961 (N_4961,N_3745,N_3693);
nand U4962 (N_4962,N_3742,N_3025);
nor U4963 (N_4963,N_3175,N_3357);
or U4964 (N_4964,N_3735,N_3198);
nand U4965 (N_4965,N_3108,N_3774);
or U4966 (N_4966,N_3661,N_3071);
and U4967 (N_4967,N_3416,N_3339);
or U4968 (N_4968,N_3542,N_3332);
nand U4969 (N_4969,N_3105,N_3889);
nand U4970 (N_4970,N_3925,N_3501);
nand U4971 (N_4971,N_3574,N_3984);
nor U4972 (N_4972,N_3073,N_3343);
xnor U4973 (N_4973,N_3356,N_3668);
and U4974 (N_4974,N_3541,N_3846);
or U4975 (N_4975,N_3755,N_3055);
and U4976 (N_4976,N_3415,N_3902);
nand U4977 (N_4977,N_3680,N_3249);
nand U4978 (N_4978,N_3689,N_3843);
or U4979 (N_4979,N_3191,N_3750);
nor U4980 (N_4980,N_3773,N_3457);
or U4981 (N_4981,N_3433,N_3143);
and U4982 (N_4982,N_3091,N_3817);
or U4983 (N_4983,N_3454,N_3076);
nand U4984 (N_4984,N_3111,N_3206);
nor U4985 (N_4985,N_3208,N_3672);
or U4986 (N_4986,N_3817,N_3660);
nand U4987 (N_4987,N_3451,N_3750);
nor U4988 (N_4988,N_3782,N_3869);
and U4989 (N_4989,N_3889,N_3558);
or U4990 (N_4990,N_3657,N_3388);
nor U4991 (N_4991,N_3234,N_3577);
or U4992 (N_4992,N_3926,N_3841);
xnor U4993 (N_4993,N_3850,N_3574);
nor U4994 (N_4994,N_3138,N_3510);
or U4995 (N_4995,N_3616,N_3851);
and U4996 (N_4996,N_3122,N_3815);
or U4997 (N_4997,N_3832,N_3273);
nor U4998 (N_4998,N_3563,N_3371);
nor U4999 (N_4999,N_3810,N_3611);
nor U5000 (N_5000,N_4867,N_4531);
nor U5001 (N_5001,N_4170,N_4772);
or U5002 (N_5002,N_4947,N_4380);
or U5003 (N_5003,N_4568,N_4451);
or U5004 (N_5004,N_4882,N_4542);
or U5005 (N_5005,N_4786,N_4626);
nor U5006 (N_5006,N_4888,N_4712);
xor U5007 (N_5007,N_4713,N_4738);
nor U5008 (N_5008,N_4570,N_4832);
or U5009 (N_5009,N_4364,N_4447);
nand U5010 (N_5010,N_4472,N_4311);
or U5011 (N_5011,N_4111,N_4749);
nand U5012 (N_5012,N_4850,N_4413);
nor U5013 (N_5013,N_4303,N_4351);
or U5014 (N_5014,N_4317,N_4774);
or U5015 (N_5015,N_4457,N_4366);
nand U5016 (N_5016,N_4191,N_4758);
and U5017 (N_5017,N_4824,N_4766);
nand U5018 (N_5018,N_4225,N_4160);
nand U5019 (N_5019,N_4704,N_4708);
nand U5020 (N_5020,N_4982,N_4794);
and U5021 (N_5021,N_4228,N_4623);
nand U5022 (N_5022,N_4473,N_4927);
and U5023 (N_5023,N_4916,N_4432);
nor U5024 (N_5024,N_4625,N_4847);
or U5025 (N_5025,N_4983,N_4929);
and U5026 (N_5026,N_4498,N_4501);
and U5027 (N_5027,N_4067,N_4230);
nor U5028 (N_5028,N_4492,N_4723);
or U5029 (N_5029,N_4653,N_4593);
and U5030 (N_5030,N_4068,N_4171);
and U5031 (N_5031,N_4254,N_4592);
nand U5032 (N_5032,N_4322,N_4372);
and U5033 (N_5033,N_4149,N_4316);
and U5034 (N_5034,N_4085,N_4384);
and U5035 (N_5035,N_4392,N_4352);
and U5036 (N_5036,N_4659,N_4865);
nor U5037 (N_5037,N_4703,N_4962);
and U5038 (N_5038,N_4206,N_4591);
and U5039 (N_5039,N_4894,N_4797);
or U5040 (N_5040,N_4602,N_4657);
or U5041 (N_5041,N_4101,N_4032);
nor U5042 (N_5042,N_4527,N_4891);
nor U5043 (N_5043,N_4331,N_4016);
or U5044 (N_5044,N_4561,N_4686);
and U5045 (N_5045,N_4275,N_4378);
or U5046 (N_5046,N_4907,N_4603);
and U5047 (N_5047,N_4862,N_4386);
nand U5048 (N_5048,N_4123,N_4197);
or U5049 (N_5049,N_4036,N_4724);
nor U5050 (N_5050,N_4409,N_4544);
or U5051 (N_5051,N_4244,N_4585);
and U5052 (N_5052,N_4655,N_4512);
and U5053 (N_5053,N_4672,N_4822);
nor U5054 (N_5054,N_4779,N_4283);
xor U5055 (N_5055,N_4614,N_4465);
and U5056 (N_5056,N_4966,N_4554);
and U5057 (N_5057,N_4575,N_4428);
and U5058 (N_5058,N_4956,N_4854);
and U5059 (N_5059,N_4363,N_4619);
nor U5060 (N_5060,N_4484,N_4391);
and U5061 (N_5061,N_4096,N_4470);
or U5062 (N_5062,N_4532,N_4058);
and U5063 (N_5063,N_4759,N_4462);
nand U5064 (N_5064,N_4569,N_4833);
nor U5065 (N_5065,N_4654,N_4350);
nor U5066 (N_5066,N_4937,N_4715);
nand U5067 (N_5067,N_4019,N_4787);
nor U5068 (N_5068,N_4541,N_4651);
or U5069 (N_5069,N_4770,N_4629);
nand U5070 (N_5070,N_4471,N_4106);
and U5071 (N_5071,N_4248,N_4995);
or U5072 (N_5072,N_4271,N_4388);
or U5073 (N_5073,N_4130,N_4688);
nor U5074 (N_5074,N_4204,N_4714);
nor U5075 (N_5075,N_4518,N_4120);
and U5076 (N_5076,N_4645,N_4941);
nor U5077 (N_5077,N_4503,N_4908);
nand U5078 (N_5078,N_4341,N_4073);
or U5079 (N_5079,N_4985,N_4436);
nand U5080 (N_5080,N_4219,N_4513);
and U5081 (N_5081,N_4773,N_4439);
and U5082 (N_5082,N_4805,N_4356);
or U5083 (N_5083,N_4475,N_4474);
nand U5084 (N_5084,N_4009,N_4520);
and U5085 (N_5085,N_4940,N_4666);
or U5086 (N_5086,N_4030,N_4948);
nor U5087 (N_5087,N_4987,N_4615);
and U5088 (N_5088,N_4493,N_4636);
nor U5089 (N_5089,N_4329,N_4419);
or U5090 (N_5090,N_4334,N_4266);
nand U5091 (N_5091,N_4379,N_4646);
nor U5092 (N_5092,N_4014,N_4294);
nor U5093 (N_5093,N_4040,N_4321);
nor U5094 (N_5094,N_4309,N_4567);
nor U5095 (N_5095,N_4718,N_4878);
or U5096 (N_5096,N_4705,N_4820);
nand U5097 (N_5097,N_4722,N_4214);
nand U5098 (N_5098,N_4288,N_4885);
nand U5099 (N_5099,N_4263,N_4818);
nand U5100 (N_5100,N_4670,N_4935);
and U5101 (N_5101,N_4902,N_4959);
and U5102 (N_5102,N_4611,N_4583);
nor U5103 (N_5103,N_4369,N_4678);
and U5104 (N_5104,N_4216,N_4018);
nor U5105 (N_5105,N_4652,N_4119);
or U5106 (N_5106,N_4280,N_4381);
and U5107 (N_5107,N_4113,N_4740);
and U5108 (N_5108,N_4576,N_4840);
or U5109 (N_5109,N_4958,N_4564);
nand U5110 (N_5110,N_4084,N_4869);
nor U5111 (N_5111,N_4523,N_4530);
nor U5112 (N_5112,N_4154,N_4207);
or U5113 (N_5113,N_4621,N_4024);
nand U5114 (N_5114,N_4889,N_4559);
nor U5115 (N_5115,N_4269,N_4855);
nor U5116 (N_5116,N_4826,N_4563);
and U5117 (N_5117,N_4199,N_4033);
or U5118 (N_5118,N_4081,N_4557);
and U5119 (N_5119,N_4047,N_4755);
nor U5120 (N_5120,N_4168,N_4600);
nor U5121 (N_5121,N_4080,N_4013);
nand U5122 (N_5122,N_4857,N_4744);
nand U5123 (N_5123,N_4326,N_4796);
and U5124 (N_5124,N_4782,N_4397);
nand U5125 (N_5125,N_4696,N_4692);
nor U5126 (N_5126,N_4343,N_4990);
or U5127 (N_5127,N_4886,N_4267);
or U5128 (N_5128,N_4203,N_4618);
nand U5129 (N_5129,N_4522,N_4701);
nor U5130 (N_5130,N_4565,N_4582);
nand U5131 (N_5131,N_4211,N_4890);
nor U5132 (N_5132,N_4868,N_4620);
nor U5133 (N_5133,N_4529,N_4789);
nand U5134 (N_5134,N_4859,N_4421);
and U5135 (N_5135,N_4028,N_4955);
or U5136 (N_5136,N_4074,N_4763);
nand U5137 (N_5137,N_4534,N_4144);
nand U5138 (N_5138,N_4920,N_4368);
and U5139 (N_5139,N_4848,N_4035);
or U5140 (N_5140,N_4778,N_4416);
or U5141 (N_5141,N_4577,N_4543);
or U5142 (N_5142,N_4217,N_4183);
nor U5143 (N_5143,N_4540,N_4764);
and U5144 (N_5144,N_4390,N_4803);
nor U5145 (N_5145,N_4812,N_4861);
or U5146 (N_5146,N_4190,N_4637);
nor U5147 (N_5147,N_4994,N_4122);
nor U5148 (N_5148,N_4748,N_4076);
or U5149 (N_5149,N_4946,N_4328);
and U5150 (N_5150,N_4105,N_4877);
and U5151 (N_5151,N_4739,N_4727);
nand U5152 (N_5152,N_4992,N_4781);
nand U5153 (N_5153,N_4834,N_4580);
nand U5154 (N_5154,N_4806,N_4353);
nand U5155 (N_5155,N_4466,N_4059);
nand U5156 (N_5156,N_4936,N_4173);
nor U5157 (N_5157,N_4300,N_4307);
and U5158 (N_5158,N_4976,N_4574);
or U5159 (N_5159,N_4463,N_4771);
or U5160 (N_5160,N_4135,N_4256);
or U5161 (N_5161,N_4731,N_4142);
or U5162 (N_5162,N_4247,N_4338);
nor U5163 (N_5163,N_4658,N_4417);
nand U5164 (N_5164,N_4240,N_4427);
or U5165 (N_5165,N_4661,N_4488);
or U5166 (N_5166,N_4586,N_4752);
or U5167 (N_5167,N_4044,N_4856);
and U5168 (N_5168,N_4049,N_4091);
and U5169 (N_5169,N_4737,N_4305);
nand U5170 (N_5170,N_4196,N_4566);
nor U5171 (N_5171,N_4093,N_4761);
xor U5172 (N_5172,N_4286,N_4747);
and U5173 (N_5173,N_4944,N_4038);
nor U5174 (N_5174,N_4065,N_4006);
and U5175 (N_5175,N_4952,N_4604);
and U5176 (N_5176,N_4784,N_4118);
nand U5177 (N_5177,N_4114,N_4487);
nor U5178 (N_5178,N_4278,N_4768);
or U5179 (N_5179,N_4141,N_4802);
and U5180 (N_5180,N_4631,N_4632);
nor U5181 (N_5181,N_4819,N_4993);
nand U5182 (N_5182,N_4634,N_4053);
nor U5183 (N_5183,N_4552,N_4968);
nand U5184 (N_5184,N_4418,N_4178);
or U5185 (N_5185,N_4296,N_4975);
nor U5186 (N_5186,N_4839,N_4989);
nand U5187 (N_5187,N_4255,N_4627);
and U5188 (N_5188,N_4274,N_4965);
nand U5189 (N_5189,N_4444,N_4229);
and U5190 (N_5190,N_4679,N_4546);
or U5191 (N_5191,N_4550,N_4200);
nor U5192 (N_5192,N_4308,N_4485);
nand U5193 (N_5193,N_4525,N_4361);
nor U5194 (N_5194,N_4681,N_4751);
and U5195 (N_5195,N_4157,N_4996);
nand U5196 (N_5196,N_4125,N_4660);
or U5197 (N_5197,N_4056,N_4639);
nor U5198 (N_5198,N_4584,N_4598);
and U5199 (N_5199,N_4235,N_4745);
or U5200 (N_5200,N_4194,N_4717);
nor U5201 (N_5201,N_4015,N_4825);
nor U5202 (N_5202,N_4026,N_4360);
or U5203 (N_5203,N_4063,N_4395);
or U5204 (N_5204,N_4510,N_4450);
xor U5205 (N_5205,N_4601,N_4310);
nand U5206 (N_5206,N_4469,N_4769);
nand U5207 (N_5207,N_4181,N_4480);
nand U5208 (N_5208,N_4725,N_4268);
or U5209 (N_5209,N_4579,N_4385);
and U5210 (N_5210,N_4589,N_4187);
nor U5211 (N_5211,N_4249,N_4934);
and U5212 (N_5212,N_4339,N_4257);
or U5213 (N_5213,N_4849,N_4939);
or U5214 (N_5214,N_4342,N_4798);
or U5215 (N_5215,N_4060,N_4816);
nor U5216 (N_5216,N_4282,N_4972);
or U5217 (N_5217,N_4988,N_4648);
xnor U5218 (N_5218,N_4829,N_4949);
or U5219 (N_5219,N_4613,N_4259);
and U5220 (N_5220,N_4359,N_4333);
nor U5221 (N_5221,N_4514,N_4124);
nor U5222 (N_5222,N_4845,N_4545);
and U5223 (N_5223,N_4046,N_4134);
and U5224 (N_5224,N_4760,N_4468);
nor U5225 (N_5225,N_4588,N_4998);
nand U5226 (N_5226,N_4336,N_4838);
or U5227 (N_5227,N_4842,N_4633);
or U5228 (N_5228,N_4729,N_4597);
xnor U5229 (N_5229,N_4005,N_4176);
or U5230 (N_5230,N_4964,N_4365);
nor U5231 (N_5231,N_4398,N_4276);
and U5232 (N_5232,N_4511,N_4880);
nor U5233 (N_5233,N_4431,N_4594);
nor U5234 (N_5234,N_4180,N_4152);
nor U5235 (N_5235,N_4377,N_4314);
or U5236 (N_5236,N_4719,N_4813);
nor U5237 (N_5237,N_4950,N_4279);
nand U5238 (N_5238,N_4693,N_4136);
nand U5239 (N_5239,N_4479,N_4756);
and U5240 (N_5240,N_4224,N_4898);
xor U5241 (N_5241,N_4753,N_4151);
and U5242 (N_5242,N_4978,N_4330);
and U5243 (N_5243,N_4245,N_4892);
and U5244 (N_5244,N_4293,N_4780);
or U5245 (N_5245,N_4158,N_4066);
or U5246 (N_5246,N_4689,N_4201);
and U5247 (N_5247,N_4414,N_4879);
and U5248 (N_5248,N_4486,N_4500);
xor U5249 (N_5249,N_4698,N_4246);
and U5250 (N_5250,N_4707,N_4401);
or U5251 (N_5251,N_4437,N_4442);
and U5252 (N_5252,N_4860,N_4804);
or U5253 (N_5253,N_4393,N_4345);
and U5254 (N_5254,N_4117,N_4456);
or U5255 (N_5255,N_4808,N_4823);
and U5256 (N_5256,N_4926,N_4460);
nor U5257 (N_5257,N_4057,N_4277);
or U5258 (N_5258,N_4481,N_4710);
nor U5259 (N_5259,N_4167,N_4507);
or U5260 (N_5260,N_4521,N_4362);
or U5261 (N_5261,N_4641,N_4807);
nand U5262 (N_5262,N_4370,N_4578);
nor U5263 (N_5263,N_4502,N_4967);
or U5264 (N_5264,N_4355,N_4742);
nor U5265 (N_5265,N_4139,N_4922);
nor U5266 (N_5266,N_4494,N_4260);
nor U5267 (N_5267,N_4107,N_4656);
and U5268 (N_5268,N_4031,N_4793);
and U5269 (N_5269,N_4086,N_4238);
nor U5270 (N_5270,N_4979,N_4312);
nand U5271 (N_5271,N_4095,N_4367);
nand U5272 (N_5272,N_4943,N_4508);
or U5273 (N_5273,N_4638,N_4673);
nand U5274 (N_5274,N_4017,N_4635);
nand U5275 (N_5275,N_4020,N_4008);
nor U5276 (N_5276,N_4156,N_4932);
and U5277 (N_5277,N_4938,N_4299);
nand U5278 (N_5278,N_4509,N_4337);
nand U5279 (N_5279,N_4458,N_4213);
nor U5280 (N_5280,N_4684,N_4163);
nand U5281 (N_5281,N_4287,N_4347);
or U5282 (N_5282,N_4298,N_4411);
and U5283 (N_5283,N_4121,N_4928);
and U5284 (N_5284,N_4438,N_4148);
and U5285 (N_5285,N_4827,N_4243);
nand U5286 (N_5286,N_4528,N_4045);
nor U5287 (N_5287,N_4250,N_4129);
nor U5288 (N_5288,N_4691,N_4547);
nand U5289 (N_5289,N_4864,N_4587);
or U5290 (N_5290,N_4153,N_4261);
and U5291 (N_5291,N_4695,N_4373);
nor U5292 (N_5292,N_4108,N_4709);
or U5293 (N_5293,N_4841,N_4970);
or U5294 (N_5294,N_4918,N_4210);
nor U5295 (N_5295,N_4184,N_4387);
nand U5296 (N_5296,N_4663,N_4027);
and U5297 (N_5297,N_4415,N_4034);
nor U5298 (N_5298,N_4164,N_4133);
and U5299 (N_5299,N_4161,N_4986);
xnor U5300 (N_5300,N_4951,N_4801);
nand U5301 (N_5301,N_4991,N_4116);
nor U5302 (N_5302,N_4733,N_4304);
nand U5303 (N_5303,N_4115,N_4029);
nand U5304 (N_5304,N_4349,N_4223);
nand U5305 (N_5305,N_4205,N_4765);
nor U5306 (N_5306,N_4412,N_4306);
nand U5307 (N_5307,N_4917,N_4750);
or U5308 (N_5308,N_4910,N_4874);
nor U5309 (N_5309,N_4082,N_4143);
nand U5310 (N_5310,N_4075,N_4089);
nand U5311 (N_5311,N_4179,N_4165);
or U5312 (N_5312,N_4923,N_4186);
nor U5313 (N_5313,N_4220,N_4021);
nand U5314 (N_5314,N_4140,N_4003);
nor U5315 (N_5315,N_4555,N_4612);
nor U5316 (N_5316,N_4464,N_4110);
nand U5317 (N_5317,N_4558,N_4270);
or U5318 (N_5318,N_4650,N_4872);
nand U5319 (N_5319,N_4517,N_4630);
or U5320 (N_5320,N_4981,N_4072);
and U5321 (N_5321,N_4676,N_4757);
nand U5322 (N_5322,N_4446,N_4429);
nand U5323 (N_5323,N_4599,N_4358);
nor U5324 (N_5324,N_4548,N_4721);
nand U5325 (N_5325,N_4810,N_4374);
and U5326 (N_5326,N_4145,N_4174);
xor U5327 (N_5327,N_4628,N_4252);
nor U5328 (N_5328,N_4571,N_4665);
and U5329 (N_5329,N_4997,N_4251);
or U5330 (N_5330,N_4402,N_4933);
or U5331 (N_5331,N_4039,N_4595);
nor U5332 (N_5332,N_4895,N_4871);
nand U5333 (N_5333,N_4182,N_4999);
and U5334 (N_5334,N_4383,N_4682);
and U5335 (N_5335,N_4426,N_4461);
or U5336 (N_5336,N_4011,N_4835);
nor U5337 (N_5337,N_4327,N_4062);
or U5338 (N_5338,N_4969,N_4945);
nand U5339 (N_5339,N_4192,N_4443);
nand U5340 (N_5340,N_4324,N_4931);
or U5341 (N_5341,N_4258,N_4903);
nand U5342 (N_5342,N_4408,N_4285);
and U5343 (N_5343,N_4138,N_4609);
nand U5344 (N_5344,N_4410,N_4785);
nor U5345 (N_5345,N_4896,N_4974);
nand U5346 (N_5346,N_4128,N_4858);
nor U5347 (N_5347,N_4234,N_4497);
nor U5348 (N_5348,N_4734,N_4325);
nand U5349 (N_5349,N_4087,N_4232);
nor U5350 (N_5350,N_4150,N_4539);
and U5351 (N_5351,N_4846,N_4911);
or U5352 (N_5352,N_4876,N_4218);
and U5353 (N_5353,N_4098,N_4054);
nor U5354 (N_5354,N_4828,N_4643);
and U5355 (N_5355,N_4605,N_4132);
nand U5356 (N_5356,N_4332,N_4055);
nor U5357 (N_5357,N_4624,N_4357);
xnor U5358 (N_5358,N_4921,N_4403);
or U5359 (N_5359,N_4198,N_4253);
and U5360 (N_5360,N_4622,N_4866);
and U5361 (N_5361,N_4209,N_4071);
or U5362 (N_5362,N_4792,N_4422);
and U5363 (N_5363,N_4112,N_4445);
xor U5364 (N_5364,N_4440,N_4496);
nand U5365 (N_5365,N_4159,N_4478);
and U5366 (N_5366,N_4177,N_4851);
nand U5367 (N_5367,N_4610,N_4083);
or U5368 (N_5368,N_4700,N_4004);
nand U5369 (N_5369,N_4690,N_4195);
or U5370 (N_5370,N_4504,N_4126);
nand U5371 (N_5371,N_4536,N_4454);
nand U5372 (N_5372,N_4791,N_4884);
and U5373 (N_5373,N_4452,N_4843);
or U5374 (N_5374,N_4323,N_4137);
or U5375 (N_5375,N_4900,N_4899);
or U5376 (N_5376,N_4919,N_4448);
and U5377 (N_5377,N_4435,N_4424);
nand U5378 (N_5378,N_4732,N_4242);
and U5379 (N_5379,N_4697,N_4175);
and U5380 (N_5380,N_4208,N_4906);
nor U5381 (N_5381,N_4549,N_4425);
and U5382 (N_5382,N_4313,N_4767);
nor U5383 (N_5383,N_4320,N_4348);
or U5384 (N_5384,N_4957,N_4776);
and U5385 (N_5385,N_4389,N_4809);
or U5386 (N_5386,N_4953,N_4775);
nor U5387 (N_5387,N_4685,N_4099);
or U5388 (N_5388,N_4346,N_4668);
nand U5389 (N_5389,N_4077,N_4538);
nand U5390 (N_5390,N_4103,N_4726);
nand U5391 (N_5391,N_4743,N_4489);
or U5392 (N_5392,N_4335,N_4706);
nor U5393 (N_5393,N_4669,N_4795);
nor U5394 (N_5394,N_4495,N_4264);
and U5395 (N_5395,N_4783,N_4459);
or U5396 (N_5396,N_4984,N_4505);
and U5397 (N_5397,N_4477,N_4491);
or U5398 (N_5398,N_4844,N_4001);
or U5399 (N_5399,N_4394,N_4893);
nand U5400 (N_5400,N_4533,N_4420);
nor U5401 (N_5401,N_4711,N_4371);
and U5402 (N_5402,N_4499,N_4185);
or U5403 (N_5403,N_4674,N_4687);
or U5404 (N_5404,N_4730,N_4301);
nand U5405 (N_5405,N_4735,N_4925);
and U5406 (N_5406,N_4799,N_4694);
nor U5407 (N_5407,N_4455,N_4042);
or U5408 (N_5408,N_4960,N_4537);
nand U5409 (N_5409,N_4079,N_4404);
nand U5410 (N_5410,N_4052,N_4051);
xor U5411 (N_5411,N_4399,N_4212);
or U5412 (N_5412,N_4483,N_4172);
and U5413 (N_5413,N_4596,N_4434);
nand U5414 (N_5414,N_4284,N_4642);
and U5415 (N_5415,N_4777,N_4954);
nor U5416 (N_5416,N_4002,N_4736);
nor U5417 (N_5417,N_4406,N_4010);
nand U5418 (N_5418,N_4562,N_4400);
nand U5419 (N_5419,N_4295,N_4640);
nand U5420 (N_5420,N_4607,N_4649);
or U5421 (N_5421,N_4980,N_4762);
nand U5422 (N_5422,N_4515,N_4560);
and U5423 (N_5423,N_4396,N_4215);
nor U5424 (N_5424,N_4519,N_4169);
nor U5425 (N_5425,N_4606,N_4617);
and U5426 (N_5426,N_4716,N_4023);
and U5427 (N_5427,N_4930,N_4581);
nor U5428 (N_5428,N_4022,N_4815);
nor U5429 (N_5429,N_4667,N_4788);
nor U5430 (N_5430,N_4837,N_4664);
nor U5431 (N_5431,N_4375,N_4746);
or U5432 (N_5432,N_4092,N_4423);
nor U5433 (N_5433,N_4647,N_4887);
or U5434 (N_5434,N_4319,N_4811);
and U5435 (N_5435,N_4873,N_4094);
nand U5436 (N_5436,N_4915,N_4644);
and U5437 (N_5437,N_4821,N_4482);
and U5438 (N_5438,N_4226,N_4699);
and U5439 (N_5439,N_4449,N_4061);
nor U5440 (N_5440,N_4476,N_4572);
nand U5441 (N_5441,N_4430,N_4441);
nand U5442 (N_5442,N_4516,N_4490);
nor U5443 (N_5443,N_4162,N_4007);
or U5444 (N_5444,N_4382,N_4037);
nor U5445 (N_5445,N_4467,N_4340);
nand U5446 (N_5446,N_4616,N_4102);
nor U5447 (N_5447,N_4909,N_4506);
and U5448 (N_5448,N_4924,N_4147);
nand U5449 (N_5449,N_4297,N_4453);
nor U5450 (N_5450,N_4025,N_4202);
nand U5451 (N_5451,N_4273,N_4109);
or U5452 (N_5452,N_4146,N_4971);
nor U5453 (N_5453,N_4231,N_4675);
nand U5454 (N_5454,N_4556,N_4942);
or U5455 (N_5455,N_4189,N_4043);
and U5456 (N_5456,N_4237,N_4830);
nand U5457 (N_5457,N_4790,N_4870);
or U5458 (N_5458,N_4265,N_4608);
and U5459 (N_5459,N_4754,N_4535);
nand U5460 (N_5460,N_4680,N_4800);
or U5461 (N_5461,N_4262,N_4904);
nor U5462 (N_5462,N_4590,N_4127);
nor U5463 (N_5463,N_4881,N_4836);
nand U5464 (N_5464,N_4901,N_4064);
and U5465 (N_5465,N_4166,N_4302);
nor U5466 (N_5466,N_4239,N_4221);
or U5467 (N_5467,N_4573,N_4193);
and U5468 (N_5468,N_4272,N_4405);
and U5469 (N_5469,N_4526,N_4551);
or U5470 (N_5470,N_4078,N_4897);
nand U5471 (N_5471,N_4315,N_4292);
or U5472 (N_5472,N_4875,N_4728);
nand U5473 (N_5473,N_4671,N_4233);
xnor U5474 (N_5474,N_4973,N_4069);
nand U5475 (N_5475,N_4050,N_4961);
nand U5476 (N_5476,N_4289,N_4720);
and U5477 (N_5477,N_4188,N_4236);
nand U5478 (N_5478,N_4088,N_4912);
nor U5479 (N_5479,N_4963,N_4407);
nor U5480 (N_5480,N_4155,N_4041);
or U5481 (N_5481,N_4814,N_4097);
or U5482 (N_5482,N_4831,N_4090);
xnor U5483 (N_5483,N_4702,N_4318);
or U5484 (N_5484,N_4070,N_4376);
nand U5485 (N_5485,N_4131,N_4524);
or U5486 (N_5486,N_4913,N_4853);
nand U5487 (N_5487,N_4852,N_4291);
or U5488 (N_5488,N_4817,N_4905);
nand U5489 (N_5489,N_4012,N_4553);
nand U5490 (N_5490,N_4863,N_4433);
or U5491 (N_5491,N_4662,N_4290);
nand U5492 (N_5492,N_4344,N_4241);
or U5493 (N_5493,N_4977,N_4914);
or U5494 (N_5494,N_4000,N_4048);
nand U5495 (N_5495,N_4677,N_4100);
or U5496 (N_5496,N_4281,N_4683);
nand U5497 (N_5497,N_4222,N_4104);
and U5498 (N_5498,N_4883,N_4227);
nor U5499 (N_5499,N_4354,N_4741);
nor U5500 (N_5500,N_4539,N_4094);
or U5501 (N_5501,N_4674,N_4789);
xor U5502 (N_5502,N_4526,N_4569);
nor U5503 (N_5503,N_4829,N_4881);
and U5504 (N_5504,N_4841,N_4590);
nor U5505 (N_5505,N_4948,N_4739);
nand U5506 (N_5506,N_4270,N_4737);
and U5507 (N_5507,N_4996,N_4249);
nor U5508 (N_5508,N_4924,N_4710);
and U5509 (N_5509,N_4171,N_4358);
nand U5510 (N_5510,N_4648,N_4156);
or U5511 (N_5511,N_4941,N_4679);
nand U5512 (N_5512,N_4930,N_4100);
and U5513 (N_5513,N_4686,N_4676);
nor U5514 (N_5514,N_4785,N_4108);
and U5515 (N_5515,N_4242,N_4117);
and U5516 (N_5516,N_4701,N_4642);
nor U5517 (N_5517,N_4400,N_4836);
nor U5518 (N_5518,N_4659,N_4320);
and U5519 (N_5519,N_4846,N_4088);
or U5520 (N_5520,N_4515,N_4450);
nand U5521 (N_5521,N_4573,N_4752);
nor U5522 (N_5522,N_4046,N_4451);
nand U5523 (N_5523,N_4053,N_4346);
nand U5524 (N_5524,N_4359,N_4861);
nor U5525 (N_5525,N_4819,N_4424);
or U5526 (N_5526,N_4509,N_4114);
and U5527 (N_5527,N_4537,N_4590);
or U5528 (N_5528,N_4292,N_4919);
or U5529 (N_5529,N_4486,N_4340);
nor U5530 (N_5530,N_4685,N_4868);
nand U5531 (N_5531,N_4362,N_4852);
nor U5532 (N_5532,N_4300,N_4921);
or U5533 (N_5533,N_4947,N_4668);
and U5534 (N_5534,N_4287,N_4703);
nand U5535 (N_5535,N_4480,N_4241);
or U5536 (N_5536,N_4078,N_4703);
nand U5537 (N_5537,N_4026,N_4482);
nor U5538 (N_5538,N_4710,N_4174);
nand U5539 (N_5539,N_4727,N_4188);
and U5540 (N_5540,N_4114,N_4759);
and U5541 (N_5541,N_4162,N_4960);
nand U5542 (N_5542,N_4351,N_4574);
and U5543 (N_5543,N_4777,N_4319);
nor U5544 (N_5544,N_4843,N_4375);
nor U5545 (N_5545,N_4855,N_4904);
or U5546 (N_5546,N_4640,N_4534);
and U5547 (N_5547,N_4425,N_4933);
nor U5548 (N_5548,N_4468,N_4210);
nand U5549 (N_5549,N_4036,N_4317);
or U5550 (N_5550,N_4650,N_4975);
and U5551 (N_5551,N_4674,N_4520);
or U5552 (N_5552,N_4768,N_4388);
nor U5553 (N_5553,N_4912,N_4227);
and U5554 (N_5554,N_4370,N_4143);
nor U5555 (N_5555,N_4253,N_4606);
xor U5556 (N_5556,N_4462,N_4355);
nor U5557 (N_5557,N_4349,N_4895);
or U5558 (N_5558,N_4955,N_4115);
nor U5559 (N_5559,N_4969,N_4998);
nand U5560 (N_5560,N_4820,N_4452);
and U5561 (N_5561,N_4318,N_4709);
nor U5562 (N_5562,N_4866,N_4810);
nor U5563 (N_5563,N_4219,N_4265);
or U5564 (N_5564,N_4489,N_4351);
and U5565 (N_5565,N_4762,N_4247);
nor U5566 (N_5566,N_4861,N_4902);
nor U5567 (N_5567,N_4687,N_4575);
nor U5568 (N_5568,N_4122,N_4151);
nand U5569 (N_5569,N_4336,N_4579);
nor U5570 (N_5570,N_4446,N_4377);
nand U5571 (N_5571,N_4559,N_4516);
and U5572 (N_5572,N_4925,N_4608);
or U5573 (N_5573,N_4739,N_4664);
or U5574 (N_5574,N_4929,N_4683);
nor U5575 (N_5575,N_4708,N_4835);
nand U5576 (N_5576,N_4120,N_4766);
nor U5577 (N_5577,N_4262,N_4959);
nand U5578 (N_5578,N_4584,N_4486);
or U5579 (N_5579,N_4625,N_4011);
or U5580 (N_5580,N_4582,N_4978);
nor U5581 (N_5581,N_4813,N_4232);
nand U5582 (N_5582,N_4066,N_4946);
nand U5583 (N_5583,N_4543,N_4695);
nand U5584 (N_5584,N_4692,N_4288);
and U5585 (N_5585,N_4663,N_4273);
or U5586 (N_5586,N_4286,N_4762);
nand U5587 (N_5587,N_4926,N_4775);
or U5588 (N_5588,N_4086,N_4068);
and U5589 (N_5589,N_4238,N_4211);
and U5590 (N_5590,N_4366,N_4250);
nor U5591 (N_5591,N_4493,N_4242);
nor U5592 (N_5592,N_4643,N_4649);
nand U5593 (N_5593,N_4087,N_4242);
and U5594 (N_5594,N_4753,N_4894);
or U5595 (N_5595,N_4344,N_4356);
xnor U5596 (N_5596,N_4628,N_4643);
nor U5597 (N_5597,N_4513,N_4545);
or U5598 (N_5598,N_4207,N_4986);
nor U5599 (N_5599,N_4264,N_4193);
or U5600 (N_5600,N_4897,N_4604);
or U5601 (N_5601,N_4473,N_4207);
or U5602 (N_5602,N_4282,N_4695);
nor U5603 (N_5603,N_4445,N_4942);
and U5604 (N_5604,N_4662,N_4383);
or U5605 (N_5605,N_4000,N_4280);
and U5606 (N_5606,N_4144,N_4433);
nand U5607 (N_5607,N_4192,N_4794);
and U5608 (N_5608,N_4709,N_4889);
or U5609 (N_5609,N_4372,N_4846);
nand U5610 (N_5610,N_4025,N_4831);
and U5611 (N_5611,N_4609,N_4192);
nor U5612 (N_5612,N_4483,N_4489);
nor U5613 (N_5613,N_4349,N_4464);
nand U5614 (N_5614,N_4130,N_4170);
nand U5615 (N_5615,N_4628,N_4310);
and U5616 (N_5616,N_4319,N_4932);
or U5617 (N_5617,N_4828,N_4263);
or U5618 (N_5618,N_4406,N_4252);
nand U5619 (N_5619,N_4905,N_4678);
or U5620 (N_5620,N_4163,N_4177);
or U5621 (N_5621,N_4026,N_4866);
or U5622 (N_5622,N_4005,N_4863);
and U5623 (N_5623,N_4116,N_4740);
or U5624 (N_5624,N_4634,N_4042);
xor U5625 (N_5625,N_4999,N_4228);
xnor U5626 (N_5626,N_4272,N_4834);
nor U5627 (N_5627,N_4403,N_4021);
and U5628 (N_5628,N_4371,N_4712);
and U5629 (N_5629,N_4439,N_4081);
nand U5630 (N_5630,N_4057,N_4539);
or U5631 (N_5631,N_4352,N_4731);
or U5632 (N_5632,N_4766,N_4670);
nor U5633 (N_5633,N_4017,N_4015);
and U5634 (N_5634,N_4777,N_4879);
xnor U5635 (N_5635,N_4967,N_4862);
nand U5636 (N_5636,N_4352,N_4451);
and U5637 (N_5637,N_4991,N_4449);
and U5638 (N_5638,N_4437,N_4133);
nand U5639 (N_5639,N_4215,N_4472);
nand U5640 (N_5640,N_4468,N_4562);
nand U5641 (N_5641,N_4615,N_4111);
and U5642 (N_5642,N_4237,N_4288);
or U5643 (N_5643,N_4315,N_4714);
nand U5644 (N_5644,N_4739,N_4372);
or U5645 (N_5645,N_4451,N_4038);
or U5646 (N_5646,N_4243,N_4824);
nand U5647 (N_5647,N_4319,N_4361);
nor U5648 (N_5648,N_4828,N_4612);
or U5649 (N_5649,N_4493,N_4519);
and U5650 (N_5650,N_4403,N_4378);
nand U5651 (N_5651,N_4913,N_4968);
or U5652 (N_5652,N_4074,N_4079);
or U5653 (N_5653,N_4426,N_4181);
or U5654 (N_5654,N_4678,N_4063);
or U5655 (N_5655,N_4521,N_4636);
nor U5656 (N_5656,N_4083,N_4189);
and U5657 (N_5657,N_4335,N_4283);
and U5658 (N_5658,N_4899,N_4856);
nor U5659 (N_5659,N_4730,N_4735);
nand U5660 (N_5660,N_4890,N_4342);
and U5661 (N_5661,N_4943,N_4986);
nand U5662 (N_5662,N_4471,N_4085);
nor U5663 (N_5663,N_4726,N_4003);
nand U5664 (N_5664,N_4214,N_4314);
or U5665 (N_5665,N_4708,N_4383);
nand U5666 (N_5666,N_4105,N_4233);
or U5667 (N_5667,N_4532,N_4809);
nand U5668 (N_5668,N_4836,N_4607);
nand U5669 (N_5669,N_4814,N_4892);
or U5670 (N_5670,N_4116,N_4182);
nand U5671 (N_5671,N_4189,N_4839);
and U5672 (N_5672,N_4705,N_4371);
nand U5673 (N_5673,N_4568,N_4690);
nor U5674 (N_5674,N_4213,N_4314);
or U5675 (N_5675,N_4053,N_4844);
or U5676 (N_5676,N_4340,N_4212);
and U5677 (N_5677,N_4806,N_4840);
and U5678 (N_5678,N_4438,N_4325);
nor U5679 (N_5679,N_4479,N_4548);
nand U5680 (N_5680,N_4659,N_4612);
or U5681 (N_5681,N_4688,N_4180);
nand U5682 (N_5682,N_4879,N_4063);
nand U5683 (N_5683,N_4876,N_4867);
nand U5684 (N_5684,N_4827,N_4386);
nand U5685 (N_5685,N_4755,N_4954);
xnor U5686 (N_5686,N_4937,N_4483);
or U5687 (N_5687,N_4205,N_4039);
or U5688 (N_5688,N_4148,N_4788);
nand U5689 (N_5689,N_4039,N_4867);
or U5690 (N_5690,N_4030,N_4651);
nand U5691 (N_5691,N_4701,N_4066);
or U5692 (N_5692,N_4166,N_4212);
xnor U5693 (N_5693,N_4113,N_4549);
or U5694 (N_5694,N_4401,N_4594);
nor U5695 (N_5695,N_4727,N_4166);
and U5696 (N_5696,N_4088,N_4600);
and U5697 (N_5697,N_4255,N_4292);
or U5698 (N_5698,N_4694,N_4778);
nor U5699 (N_5699,N_4658,N_4486);
xnor U5700 (N_5700,N_4458,N_4384);
nand U5701 (N_5701,N_4780,N_4618);
nand U5702 (N_5702,N_4968,N_4311);
or U5703 (N_5703,N_4089,N_4463);
nor U5704 (N_5704,N_4593,N_4569);
or U5705 (N_5705,N_4537,N_4972);
nor U5706 (N_5706,N_4626,N_4870);
and U5707 (N_5707,N_4480,N_4507);
or U5708 (N_5708,N_4267,N_4535);
nand U5709 (N_5709,N_4380,N_4767);
and U5710 (N_5710,N_4286,N_4317);
nand U5711 (N_5711,N_4163,N_4060);
or U5712 (N_5712,N_4750,N_4032);
and U5713 (N_5713,N_4406,N_4922);
or U5714 (N_5714,N_4188,N_4260);
or U5715 (N_5715,N_4497,N_4125);
or U5716 (N_5716,N_4904,N_4479);
or U5717 (N_5717,N_4936,N_4820);
and U5718 (N_5718,N_4841,N_4737);
nor U5719 (N_5719,N_4164,N_4277);
or U5720 (N_5720,N_4504,N_4263);
nor U5721 (N_5721,N_4527,N_4751);
and U5722 (N_5722,N_4709,N_4433);
and U5723 (N_5723,N_4899,N_4969);
nand U5724 (N_5724,N_4201,N_4090);
nor U5725 (N_5725,N_4585,N_4292);
nor U5726 (N_5726,N_4442,N_4476);
xor U5727 (N_5727,N_4634,N_4344);
and U5728 (N_5728,N_4096,N_4081);
and U5729 (N_5729,N_4442,N_4841);
nand U5730 (N_5730,N_4680,N_4196);
or U5731 (N_5731,N_4703,N_4602);
nor U5732 (N_5732,N_4170,N_4269);
or U5733 (N_5733,N_4817,N_4708);
nor U5734 (N_5734,N_4495,N_4932);
nor U5735 (N_5735,N_4222,N_4274);
nand U5736 (N_5736,N_4579,N_4057);
and U5737 (N_5737,N_4976,N_4784);
and U5738 (N_5738,N_4443,N_4622);
or U5739 (N_5739,N_4120,N_4928);
and U5740 (N_5740,N_4195,N_4696);
and U5741 (N_5741,N_4888,N_4388);
xnor U5742 (N_5742,N_4082,N_4787);
nand U5743 (N_5743,N_4689,N_4054);
nor U5744 (N_5744,N_4714,N_4372);
or U5745 (N_5745,N_4370,N_4585);
or U5746 (N_5746,N_4487,N_4579);
nor U5747 (N_5747,N_4855,N_4092);
nor U5748 (N_5748,N_4316,N_4934);
nand U5749 (N_5749,N_4609,N_4890);
or U5750 (N_5750,N_4380,N_4427);
nor U5751 (N_5751,N_4280,N_4639);
or U5752 (N_5752,N_4771,N_4077);
nor U5753 (N_5753,N_4850,N_4059);
nor U5754 (N_5754,N_4634,N_4289);
nor U5755 (N_5755,N_4359,N_4407);
or U5756 (N_5756,N_4263,N_4611);
nand U5757 (N_5757,N_4379,N_4363);
nand U5758 (N_5758,N_4221,N_4016);
or U5759 (N_5759,N_4345,N_4303);
and U5760 (N_5760,N_4743,N_4224);
nand U5761 (N_5761,N_4036,N_4026);
nand U5762 (N_5762,N_4757,N_4863);
or U5763 (N_5763,N_4023,N_4912);
or U5764 (N_5764,N_4988,N_4592);
and U5765 (N_5765,N_4448,N_4934);
and U5766 (N_5766,N_4950,N_4846);
nor U5767 (N_5767,N_4772,N_4026);
or U5768 (N_5768,N_4783,N_4137);
nand U5769 (N_5769,N_4232,N_4750);
nor U5770 (N_5770,N_4847,N_4204);
or U5771 (N_5771,N_4969,N_4263);
and U5772 (N_5772,N_4848,N_4147);
and U5773 (N_5773,N_4958,N_4043);
nor U5774 (N_5774,N_4323,N_4099);
nand U5775 (N_5775,N_4521,N_4150);
nor U5776 (N_5776,N_4829,N_4672);
nor U5777 (N_5777,N_4814,N_4083);
nor U5778 (N_5778,N_4095,N_4057);
and U5779 (N_5779,N_4811,N_4905);
or U5780 (N_5780,N_4497,N_4891);
and U5781 (N_5781,N_4811,N_4637);
nand U5782 (N_5782,N_4521,N_4583);
and U5783 (N_5783,N_4356,N_4842);
or U5784 (N_5784,N_4561,N_4565);
nand U5785 (N_5785,N_4104,N_4191);
nand U5786 (N_5786,N_4612,N_4494);
or U5787 (N_5787,N_4874,N_4913);
and U5788 (N_5788,N_4943,N_4989);
nor U5789 (N_5789,N_4877,N_4064);
nor U5790 (N_5790,N_4143,N_4356);
xor U5791 (N_5791,N_4685,N_4087);
nand U5792 (N_5792,N_4576,N_4735);
nand U5793 (N_5793,N_4411,N_4901);
nand U5794 (N_5794,N_4077,N_4027);
nand U5795 (N_5795,N_4992,N_4083);
or U5796 (N_5796,N_4266,N_4883);
nor U5797 (N_5797,N_4191,N_4277);
nor U5798 (N_5798,N_4815,N_4869);
and U5799 (N_5799,N_4621,N_4363);
nor U5800 (N_5800,N_4338,N_4517);
and U5801 (N_5801,N_4666,N_4170);
and U5802 (N_5802,N_4387,N_4130);
and U5803 (N_5803,N_4696,N_4927);
and U5804 (N_5804,N_4734,N_4281);
nor U5805 (N_5805,N_4672,N_4292);
nor U5806 (N_5806,N_4057,N_4445);
nand U5807 (N_5807,N_4913,N_4441);
and U5808 (N_5808,N_4605,N_4405);
nor U5809 (N_5809,N_4644,N_4396);
and U5810 (N_5810,N_4685,N_4857);
and U5811 (N_5811,N_4415,N_4646);
and U5812 (N_5812,N_4389,N_4721);
and U5813 (N_5813,N_4589,N_4105);
or U5814 (N_5814,N_4694,N_4257);
nand U5815 (N_5815,N_4639,N_4344);
nor U5816 (N_5816,N_4978,N_4153);
nor U5817 (N_5817,N_4889,N_4000);
and U5818 (N_5818,N_4818,N_4227);
and U5819 (N_5819,N_4385,N_4218);
or U5820 (N_5820,N_4830,N_4465);
nand U5821 (N_5821,N_4561,N_4323);
nor U5822 (N_5822,N_4941,N_4358);
nor U5823 (N_5823,N_4556,N_4040);
or U5824 (N_5824,N_4229,N_4941);
nor U5825 (N_5825,N_4905,N_4916);
and U5826 (N_5826,N_4957,N_4544);
nand U5827 (N_5827,N_4252,N_4912);
or U5828 (N_5828,N_4500,N_4903);
and U5829 (N_5829,N_4908,N_4235);
and U5830 (N_5830,N_4601,N_4848);
or U5831 (N_5831,N_4692,N_4824);
and U5832 (N_5832,N_4787,N_4673);
nor U5833 (N_5833,N_4920,N_4507);
or U5834 (N_5834,N_4399,N_4843);
and U5835 (N_5835,N_4937,N_4312);
nand U5836 (N_5836,N_4957,N_4842);
nor U5837 (N_5837,N_4385,N_4495);
and U5838 (N_5838,N_4087,N_4009);
nor U5839 (N_5839,N_4832,N_4120);
nand U5840 (N_5840,N_4976,N_4067);
nor U5841 (N_5841,N_4651,N_4164);
or U5842 (N_5842,N_4636,N_4718);
nor U5843 (N_5843,N_4009,N_4855);
nor U5844 (N_5844,N_4693,N_4970);
nand U5845 (N_5845,N_4401,N_4899);
nand U5846 (N_5846,N_4623,N_4143);
and U5847 (N_5847,N_4634,N_4537);
nor U5848 (N_5848,N_4596,N_4494);
nor U5849 (N_5849,N_4942,N_4968);
and U5850 (N_5850,N_4088,N_4296);
nand U5851 (N_5851,N_4205,N_4154);
nor U5852 (N_5852,N_4285,N_4330);
and U5853 (N_5853,N_4129,N_4043);
nor U5854 (N_5854,N_4686,N_4783);
xnor U5855 (N_5855,N_4247,N_4824);
and U5856 (N_5856,N_4391,N_4282);
nand U5857 (N_5857,N_4560,N_4069);
nor U5858 (N_5858,N_4612,N_4223);
nor U5859 (N_5859,N_4052,N_4623);
nand U5860 (N_5860,N_4563,N_4388);
or U5861 (N_5861,N_4387,N_4628);
nand U5862 (N_5862,N_4114,N_4809);
nand U5863 (N_5863,N_4276,N_4117);
and U5864 (N_5864,N_4520,N_4230);
and U5865 (N_5865,N_4415,N_4621);
nor U5866 (N_5866,N_4818,N_4463);
or U5867 (N_5867,N_4748,N_4804);
and U5868 (N_5868,N_4513,N_4274);
nand U5869 (N_5869,N_4564,N_4118);
nand U5870 (N_5870,N_4180,N_4301);
and U5871 (N_5871,N_4462,N_4902);
or U5872 (N_5872,N_4810,N_4287);
and U5873 (N_5873,N_4878,N_4011);
nor U5874 (N_5874,N_4945,N_4959);
or U5875 (N_5875,N_4339,N_4701);
nand U5876 (N_5876,N_4355,N_4889);
nor U5877 (N_5877,N_4846,N_4986);
nand U5878 (N_5878,N_4126,N_4507);
and U5879 (N_5879,N_4326,N_4950);
nor U5880 (N_5880,N_4945,N_4501);
and U5881 (N_5881,N_4025,N_4935);
nor U5882 (N_5882,N_4272,N_4669);
nand U5883 (N_5883,N_4518,N_4284);
and U5884 (N_5884,N_4010,N_4067);
nor U5885 (N_5885,N_4210,N_4930);
and U5886 (N_5886,N_4917,N_4795);
nor U5887 (N_5887,N_4401,N_4809);
nor U5888 (N_5888,N_4976,N_4845);
nor U5889 (N_5889,N_4023,N_4586);
nand U5890 (N_5890,N_4530,N_4174);
nand U5891 (N_5891,N_4675,N_4019);
nor U5892 (N_5892,N_4902,N_4127);
nor U5893 (N_5893,N_4726,N_4957);
nand U5894 (N_5894,N_4419,N_4733);
and U5895 (N_5895,N_4856,N_4390);
and U5896 (N_5896,N_4536,N_4151);
nor U5897 (N_5897,N_4397,N_4954);
or U5898 (N_5898,N_4424,N_4266);
and U5899 (N_5899,N_4948,N_4771);
nand U5900 (N_5900,N_4752,N_4271);
and U5901 (N_5901,N_4880,N_4083);
and U5902 (N_5902,N_4257,N_4123);
or U5903 (N_5903,N_4446,N_4795);
nor U5904 (N_5904,N_4181,N_4555);
nand U5905 (N_5905,N_4576,N_4240);
nand U5906 (N_5906,N_4509,N_4479);
or U5907 (N_5907,N_4160,N_4202);
nand U5908 (N_5908,N_4707,N_4585);
and U5909 (N_5909,N_4507,N_4289);
nand U5910 (N_5910,N_4376,N_4076);
and U5911 (N_5911,N_4022,N_4209);
and U5912 (N_5912,N_4941,N_4190);
nor U5913 (N_5913,N_4022,N_4795);
and U5914 (N_5914,N_4045,N_4849);
and U5915 (N_5915,N_4223,N_4999);
nand U5916 (N_5916,N_4597,N_4225);
or U5917 (N_5917,N_4218,N_4595);
nand U5918 (N_5918,N_4374,N_4028);
or U5919 (N_5919,N_4100,N_4699);
and U5920 (N_5920,N_4044,N_4019);
or U5921 (N_5921,N_4296,N_4243);
or U5922 (N_5922,N_4217,N_4198);
or U5923 (N_5923,N_4352,N_4175);
and U5924 (N_5924,N_4300,N_4282);
and U5925 (N_5925,N_4054,N_4912);
nor U5926 (N_5926,N_4588,N_4178);
and U5927 (N_5927,N_4115,N_4390);
and U5928 (N_5928,N_4860,N_4821);
and U5929 (N_5929,N_4594,N_4125);
nand U5930 (N_5930,N_4445,N_4686);
nor U5931 (N_5931,N_4875,N_4971);
or U5932 (N_5932,N_4562,N_4767);
nand U5933 (N_5933,N_4583,N_4829);
nand U5934 (N_5934,N_4114,N_4290);
nand U5935 (N_5935,N_4455,N_4354);
or U5936 (N_5936,N_4818,N_4498);
xor U5937 (N_5937,N_4262,N_4199);
or U5938 (N_5938,N_4832,N_4218);
or U5939 (N_5939,N_4520,N_4606);
nor U5940 (N_5940,N_4669,N_4529);
or U5941 (N_5941,N_4505,N_4623);
nand U5942 (N_5942,N_4334,N_4911);
xor U5943 (N_5943,N_4256,N_4629);
xor U5944 (N_5944,N_4432,N_4384);
nand U5945 (N_5945,N_4674,N_4981);
nor U5946 (N_5946,N_4229,N_4018);
and U5947 (N_5947,N_4473,N_4341);
and U5948 (N_5948,N_4384,N_4198);
or U5949 (N_5949,N_4455,N_4195);
nand U5950 (N_5950,N_4590,N_4442);
nand U5951 (N_5951,N_4813,N_4084);
nand U5952 (N_5952,N_4510,N_4370);
nand U5953 (N_5953,N_4037,N_4872);
or U5954 (N_5954,N_4145,N_4846);
or U5955 (N_5955,N_4117,N_4352);
nor U5956 (N_5956,N_4633,N_4983);
nand U5957 (N_5957,N_4244,N_4770);
and U5958 (N_5958,N_4533,N_4408);
nor U5959 (N_5959,N_4376,N_4588);
and U5960 (N_5960,N_4981,N_4051);
nor U5961 (N_5961,N_4546,N_4451);
nor U5962 (N_5962,N_4097,N_4854);
nor U5963 (N_5963,N_4161,N_4519);
and U5964 (N_5964,N_4295,N_4553);
or U5965 (N_5965,N_4069,N_4612);
nand U5966 (N_5966,N_4036,N_4965);
and U5967 (N_5967,N_4322,N_4224);
and U5968 (N_5968,N_4486,N_4155);
nor U5969 (N_5969,N_4335,N_4421);
nor U5970 (N_5970,N_4656,N_4128);
or U5971 (N_5971,N_4893,N_4583);
nor U5972 (N_5972,N_4101,N_4187);
and U5973 (N_5973,N_4574,N_4066);
nor U5974 (N_5974,N_4439,N_4479);
nor U5975 (N_5975,N_4844,N_4723);
nand U5976 (N_5976,N_4732,N_4898);
or U5977 (N_5977,N_4256,N_4404);
nand U5978 (N_5978,N_4130,N_4070);
nor U5979 (N_5979,N_4674,N_4455);
nand U5980 (N_5980,N_4696,N_4616);
and U5981 (N_5981,N_4990,N_4745);
or U5982 (N_5982,N_4274,N_4415);
and U5983 (N_5983,N_4713,N_4870);
nand U5984 (N_5984,N_4773,N_4410);
nor U5985 (N_5985,N_4866,N_4529);
or U5986 (N_5986,N_4572,N_4935);
and U5987 (N_5987,N_4579,N_4680);
or U5988 (N_5988,N_4744,N_4285);
or U5989 (N_5989,N_4465,N_4109);
nor U5990 (N_5990,N_4359,N_4003);
nand U5991 (N_5991,N_4700,N_4680);
or U5992 (N_5992,N_4370,N_4894);
or U5993 (N_5993,N_4575,N_4337);
or U5994 (N_5994,N_4507,N_4641);
or U5995 (N_5995,N_4289,N_4913);
nor U5996 (N_5996,N_4389,N_4115);
nand U5997 (N_5997,N_4348,N_4929);
nand U5998 (N_5998,N_4682,N_4547);
and U5999 (N_5999,N_4939,N_4092);
xnor U6000 (N_6000,N_5733,N_5319);
or U6001 (N_6001,N_5502,N_5176);
and U6002 (N_6002,N_5623,N_5317);
xor U6003 (N_6003,N_5556,N_5025);
and U6004 (N_6004,N_5086,N_5645);
or U6005 (N_6005,N_5248,N_5706);
nor U6006 (N_6006,N_5607,N_5469);
and U6007 (N_6007,N_5386,N_5806);
nand U6008 (N_6008,N_5089,N_5701);
or U6009 (N_6009,N_5464,N_5493);
or U6010 (N_6010,N_5872,N_5841);
or U6011 (N_6011,N_5928,N_5059);
nand U6012 (N_6012,N_5141,N_5952);
or U6013 (N_6013,N_5293,N_5898);
nor U6014 (N_6014,N_5021,N_5605);
nand U6015 (N_6015,N_5267,N_5546);
and U6016 (N_6016,N_5221,N_5197);
nand U6017 (N_6017,N_5250,N_5174);
and U6018 (N_6018,N_5827,N_5439);
or U6019 (N_6019,N_5753,N_5316);
nor U6020 (N_6020,N_5273,N_5366);
nand U6021 (N_6021,N_5077,N_5178);
or U6022 (N_6022,N_5061,N_5673);
or U6023 (N_6023,N_5096,N_5635);
nor U6024 (N_6024,N_5318,N_5154);
or U6025 (N_6025,N_5644,N_5191);
nand U6026 (N_6026,N_5982,N_5474);
or U6027 (N_6027,N_5687,N_5545);
or U6028 (N_6028,N_5268,N_5093);
or U6029 (N_6029,N_5690,N_5716);
nor U6030 (N_6030,N_5901,N_5244);
and U6031 (N_6031,N_5906,N_5462);
or U6032 (N_6032,N_5185,N_5591);
and U6033 (N_6033,N_5146,N_5815);
nand U6034 (N_6034,N_5784,N_5411);
and U6035 (N_6035,N_5613,N_5981);
and U6036 (N_6036,N_5140,N_5242);
nand U6037 (N_6037,N_5942,N_5159);
nand U6038 (N_6038,N_5307,N_5105);
nand U6039 (N_6039,N_5557,N_5330);
or U6040 (N_6040,N_5947,N_5372);
and U6041 (N_6041,N_5786,N_5726);
and U6042 (N_6042,N_5322,N_5488);
and U6043 (N_6043,N_5589,N_5905);
and U6044 (N_6044,N_5683,N_5202);
or U6045 (N_6045,N_5357,N_5045);
or U6046 (N_6046,N_5422,N_5744);
xor U6047 (N_6047,N_5388,N_5199);
nand U6048 (N_6048,N_5720,N_5455);
or U6049 (N_6049,N_5731,N_5266);
nand U6050 (N_6050,N_5611,N_5642);
nor U6051 (N_6051,N_5741,N_5990);
and U6052 (N_6052,N_5704,N_5855);
or U6053 (N_6053,N_5926,N_5732);
or U6054 (N_6054,N_5848,N_5938);
nand U6055 (N_6055,N_5847,N_5115);
and U6056 (N_6056,N_5972,N_5810);
and U6057 (N_6057,N_5097,N_5088);
nand U6058 (N_6058,N_5854,N_5012);
nand U6059 (N_6059,N_5286,N_5845);
nor U6060 (N_6060,N_5308,N_5467);
or U6061 (N_6061,N_5575,N_5087);
xnor U6062 (N_6062,N_5281,N_5999);
nand U6063 (N_6063,N_5943,N_5352);
and U6064 (N_6064,N_5071,N_5864);
nand U6065 (N_6065,N_5337,N_5870);
and U6066 (N_6066,N_5037,N_5193);
or U6067 (N_6067,N_5759,N_5179);
nand U6068 (N_6068,N_5609,N_5064);
or U6069 (N_6069,N_5371,N_5006);
and U6070 (N_6070,N_5238,N_5158);
and U6071 (N_6071,N_5807,N_5124);
nand U6072 (N_6072,N_5479,N_5038);
xnor U6073 (N_6073,N_5151,N_5822);
nand U6074 (N_6074,N_5216,N_5656);
nand U6075 (N_6075,N_5785,N_5808);
xor U6076 (N_6076,N_5583,N_5769);
nor U6077 (N_6077,N_5194,N_5849);
or U6078 (N_6078,N_5376,N_5188);
nor U6079 (N_6079,N_5950,N_5887);
and U6080 (N_6080,N_5788,N_5498);
and U6081 (N_6081,N_5987,N_5358);
and U6082 (N_6082,N_5927,N_5994);
and U6083 (N_6083,N_5084,N_5101);
nor U6084 (N_6084,N_5228,N_5483);
nor U6085 (N_6085,N_5597,N_5306);
nand U6086 (N_6086,N_5857,N_5997);
nand U6087 (N_6087,N_5405,N_5108);
or U6088 (N_6088,N_5363,N_5936);
nor U6089 (N_6089,N_5402,N_5820);
and U6090 (N_6090,N_5552,N_5082);
or U6091 (N_6091,N_5787,N_5057);
nand U6092 (N_6092,N_5588,N_5183);
nor U6093 (N_6093,N_5230,N_5102);
or U6094 (N_6094,N_5996,N_5722);
and U6095 (N_6095,N_5914,N_5135);
nand U6096 (N_6096,N_5155,N_5336);
or U6097 (N_6097,N_5364,N_5576);
nor U6098 (N_6098,N_5619,N_5190);
or U6099 (N_6099,N_5328,N_5570);
and U6100 (N_6100,N_5668,N_5044);
nor U6101 (N_6101,N_5828,N_5241);
and U6102 (N_6102,N_5875,N_5166);
nor U6103 (N_6103,N_5959,N_5091);
or U6104 (N_6104,N_5068,N_5862);
or U6105 (N_6105,N_5470,N_5234);
nor U6106 (N_6106,N_5237,N_5516);
nand U6107 (N_6107,N_5117,N_5809);
or U6108 (N_6108,N_5829,N_5378);
or U6109 (N_6109,N_5508,N_5360);
and U6110 (N_6110,N_5893,N_5081);
nand U6111 (N_6111,N_5072,N_5220);
nor U6112 (N_6112,N_5646,N_5921);
nor U6113 (N_6113,N_5053,N_5180);
nand U6114 (N_6114,N_5023,N_5128);
nor U6115 (N_6115,N_5080,N_5450);
nor U6116 (N_6116,N_5367,N_5442);
and U6117 (N_6117,N_5975,N_5418);
or U6118 (N_6118,N_5675,N_5401);
nand U6119 (N_6119,N_5526,N_5587);
and U6120 (N_6120,N_5349,N_5647);
nand U6121 (N_6121,N_5963,N_5835);
and U6122 (N_6122,N_5399,N_5288);
nor U6123 (N_6123,N_5133,N_5377);
nor U6124 (N_6124,N_5487,N_5946);
nand U6125 (N_6125,N_5544,N_5648);
and U6126 (N_6126,N_5163,N_5004);
nor U6127 (N_6127,N_5627,N_5560);
or U6128 (N_6128,N_5079,N_5016);
nand U6129 (N_6129,N_5305,N_5908);
and U6130 (N_6130,N_5419,N_5655);
and U6131 (N_6131,N_5641,N_5172);
or U6132 (N_6132,N_5030,N_5505);
nor U6133 (N_6133,N_5264,N_5246);
xor U6134 (N_6134,N_5814,N_5734);
nor U6135 (N_6135,N_5276,N_5931);
nor U6136 (N_6136,N_5674,N_5076);
or U6137 (N_6137,N_5761,N_5348);
nor U6138 (N_6138,N_5111,N_5995);
nor U6139 (N_6139,N_5750,N_5177);
nand U6140 (N_6140,N_5684,N_5798);
nand U6141 (N_6141,N_5708,N_5599);
nor U6142 (N_6142,N_5555,N_5507);
nor U6143 (N_6143,N_5916,N_5280);
or U6144 (N_6144,N_5932,N_5430);
and U6145 (N_6145,N_5837,N_5586);
and U6146 (N_6146,N_5326,N_5638);
nor U6147 (N_6147,N_5412,N_5425);
or U6148 (N_6148,N_5533,N_5033);
and U6149 (N_6149,N_5491,N_5410);
nand U6150 (N_6150,N_5136,N_5781);
nor U6151 (N_6151,N_5413,N_5294);
or U6152 (N_6152,N_5964,N_5340);
or U6153 (N_6153,N_5098,N_5398);
nand U6154 (N_6154,N_5737,N_5390);
nand U6155 (N_6155,N_5940,N_5253);
or U6156 (N_6156,N_5368,N_5739);
nor U6157 (N_6157,N_5725,N_5011);
and U6158 (N_6158,N_5572,N_5070);
nor U6159 (N_6159,N_5486,N_5900);
and U6160 (N_6160,N_5937,N_5629);
and U6161 (N_6161,N_5275,N_5272);
and U6162 (N_6162,N_5126,N_5239);
nor U6163 (N_6163,N_5834,N_5303);
or U6164 (N_6164,N_5020,N_5351);
nand U6165 (N_6165,N_5974,N_5512);
or U6166 (N_6166,N_5354,N_5547);
nor U6167 (N_6167,N_5153,N_5078);
nand U6168 (N_6168,N_5417,N_5973);
and U6169 (N_6169,N_5649,N_5839);
and U6170 (N_6170,N_5407,N_5592);
nand U6171 (N_6171,N_5663,N_5658);
xnor U6172 (N_6172,N_5681,N_5876);
nand U6173 (N_6173,N_5760,N_5035);
nor U6174 (N_6174,N_5813,N_5953);
nor U6175 (N_6175,N_5500,N_5110);
nand U6176 (N_6176,N_5899,N_5224);
nor U6177 (N_6177,N_5453,N_5186);
nand U6178 (N_6178,N_5454,N_5618);
and U6179 (N_6179,N_5014,N_5149);
nor U6180 (N_6180,N_5143,N_5564);
or U6181 (N_6181,N_5332,N_5490);
nor U6182 (N_6182,N_5260,N_5338);
nand U6183 (N_6183,N_5888,N_5840);
nor U6184 (N_6184,N_5799,N_5327);
or U6185 (N_6185,N_5171,N_5593);
nand U6186 (N_6186,N_5740,N_5287);
or U6187 (N_6187,N_5812,N_5122);
and U6188 (N_6188,N_5831,N_5971);
xor U6189 (N_6189,N_5139,N_5047);
nand U6190 (N_6190,N_5615,N_5707);
nor U6191 (N_6191,N_5393,N_5604);
and U6192 (N_6192,N_5382,N_5883);
nor U6193 (N_6193,N_5823,N_5075);
nand U6194 (N_6194,N_5529,N_5521);
and U6195 (N_6195,N_5015,N_5951);
nor U6196 (N_6196,N_5119,N_5863);
or U6197 (N_6197,N_5198,N_5851);
nand U6198 (N_6198,N_5231,N_5825);
nor U6199 (N_6199,N_5571,N_5895);
or U6200 (N_6200,N_5107,N_5695);
nand U6201 (N_6201,N_5387,N_5596);
nor U6202 (N_6202,N_5046,N_5229);
or U6203 (N_6203,N_5423,N_5986);
nor U6204 (N_6204,N_5558,N_5144);
and U6205 (N_6205,N_5217,N_5438);
nand U6206 (N_6206,N_5456,N_5632);
and U6207 (N_6207,N_5309,N_5773);
nor U6208 (N_6208,N_5670,N_5243);
or U6209 (N_6209,N_5494,N_5770);
and U6210 (N_6210,N_5672,N_5636);
nor U6211 (N_6211,N_5775,N_5836);
nor U6212 (N_6212,N_5853,N_5295);
nor U6213 (N_6213,N_5099,N_5614);
nand U6214 (N_6214,N_5634,N_5257);
nand U6215 (N_6215,N_5189,N_5513);
nor U6216 (N_6216,N_5429,N_5125);
nand U6217 (N_6217,N_5944,N_5925);
and U6218 (N_6218,N_5594,N_5054);
or U6219 (N_6219,N_5067,N_5457);
nor U6220 (N_6220,N_5639,N_5603);
or U6221 (N_6221,N_5009,N_5279);
nand U6222 (N_6222,N_5039,N_5742);
or U6223 (N_6223,N_5542,N_5471);
nor U6224 (N_6224,N_5622,N_5550);
or U6225 (N_6225,N_5466,N_5050);
nand U6226 (N_6226,N_5458,N_5090);
and U6227 (N_6227,N_5522,N_5657);
or U6228 (N_6228,N_5728,N_5539);
nor U6229 (N_6229,N_5918,N_5528);
nand U6230 (N_6230,N_5441,N_5793);
or U6231 (N_6231,N_5283,N_5600);
xnor U6232 (N_6232,N_5738,N_5882);
and U6233 (N_6233,N_5427,N_5568);
nand U6234 (N_6234,N_5700,N_5421);
nor U6235 (N_6235,N_5381,N_5917);
or U6236 (N_6236,N_5637,N_5976);
nor U6237 (N_6237,N_5948,N_5109);
nor U6238 (N_6238,N_5169,N_5984);
nand U6239 (N_6239,N_5585,N_5150);
nor U6240 (N_6240,N_5310,N_5436);
and U6241 (N_6241,N_5343,N_5311);
and U6242 (N_6242,N_5561,N_5432);
nor U6243 (N_6243,N_5499,N_5271);
and U6244 (N_6244,N_5394,N_5284);
or U6245 (N_6245,N_5519,N_5207);
nor U6246 (N_6246,N_5132,N_5383);
and U6247 (N_6247,N_5566,N_5361);
nand U6248 (N_6248,N_5989,N_5447);
nor U6249 (N_6249,N_5475,N_5856);
nor U6250 (N_6250,N_5757,N_5858);
and U6251 (N_6251,N_5515,N_5939);
nor U6252 (N_6252,N_5958,N_5184);
nor U6253 (N_6253,N_5162,N_5850);
nand U6254 (N_6254,N_5106,N_5902);
and U6255 (N_6255,N_5800,N_5152);
and U6256 (N_6256,N_5551,N_5606);
nor U6257 (N_6257,N_5113,N_5960);
nor U6258 (N_6258,N_5320,N_5679);
or U6259 (N_6259,N_5127,N_5578);
and U6260 (N_6260,N_5736,N_5208);
and U6261 (N_6261,N_5659,N_5985);
or U6262 (N_6262,N_5711,N_5195);
or U6263 (N_6263,N_5751,N_5746);
nor U6264 (N_6264,N_5541,N_5608);
or U6265 (N_6265,N_5771,N_5204);
or U6266 (N_6266,N_5083,N_5392);
nor U6267 (N_6267,N_5440,N_5962);
nor U6268 (N_6268,N_5463,N_5000);
or U6269 (N_6269,N_5930,N_5910);
or U6270 (N_6270,N_5452,N_5365);
or U6271 (N_6271,N_5803,N_5331);
or U6272 (N_6272,N_5919,N_5215);
and U6273 (N_6273,N_5764,N_5852);
nand U6274 (N_6274,N_5844,N_5617);
nor U6275 (N_6275,N_5223,N_5804);
and U6276 (N_6276,N_5923,N_5278);
nand U6277 (N_6277,N_5353,N_5312);
nor U6278 (N_6278,N_5915,N_5433);
and U6279 (N_6279,N_5896,N_5660);
or U6280 (N_6280,N_5289,N_5678);
nor U6281 (N_6281,N_5029,N_5598);
nor U6282 (N_6282,N_5933,N_5395);
nand U6283 (N_6283,N_5580,N_5833);
or U6284 (N_6284,N_5993,N_5138);
or U6285 (N_6285,N_5693,N_5894);
or U6286 (N_6286,N_5790,N_5274);
nor U6287 (N_6287,N_5375,N_5718);
and U6288 (N_6288,N_5446,N_5247);
nand U6289 (N_6289,N_5665,N_5482);
nand U6290 (N_6290,N_5341,N_5263);
nand U6291 (N_6291,N_5160,N_5729);
nor U6292 (N_6292,N_5866,N_5026);
or U6293 (N_6293,N_5503,N_5801);
or U6294 (N_6294,N_5885,N_5983);
nand U6295 (N_6295,N_5104,N_5626);
or U6296 (N_6296,N_5966,N_5206);
nor U6297 (N_6297,N_5019,N_5772);
or U6298 (N_6298,N_5339,N_5886);
and U6299 (N_6299,N_5789,N_5233);
and U6300 (N_6300,N_5650,N_5724);
nand U6301 (N_6301,N_5333,N_5218);
nand U6302 (N_6302,N_5291,N_5802);
or U6303 (N_6303,N_5406,N_5369);
or U6304 (N_6304,N_5752,N_5671);
or U6305 (N_6305,N_5779,N_5041);
and U6306 (N_6306,N_5007,N_5414);
nor U6307 (N_6307,N_5285,N_5010);
xnor U6308 (N_6308,N_5969,N_5956);
nor U6309 (N_6309,N_5514,N_5721);
nand U6310 (N_6310,N_5201,N_5922);
and U6311 (N_6311,N_5967,N_5727);
nor U6312 (N_6312,N_5538,N_5350);
nor U6313 (N_6313,N_5868,N_5762);
nor U6314 (N_6314,N_5385,N_5095);
nand U6315 (N_6315,N_5584,N_5595);
nand U6316 (N_6316,N_5485,N_5473);
nand U6317 (N_6317,N_5434,N_5379);
nand U6318 (N_6318,N_5536,N_5878);
nand U6319 (N_6319,N_5409,N_5121);
or U6320 (N_6320,N_5692,N_5748);
nor U6321 (N_6321,N_5416,N_5055);
nor U6322 (N_6322,N_5017,N_5347);
nor U6323 (N_6323,N_5749,N_5874);
nor U6324 (N_6324,N_5296,N_5477);
nand U6325 (N_6325,N_5314,N_5062);
nor U6326 (N_6326,N_5662,N_5449);
or U6327 (N_6327,N_5270,N_5624);
nand U6328 (N_6328,N_5370,N_5256);
nand U6329 (N_6329,N_5811,N_5680);
nor U6330 (N_6330,N_5713,N_5181);
nand U6331 (N_6331,N_5408,N_5774);
nor U6332 (N_6332,N_5792,N_5818);
and U6333 (N_6333,N_5816,N_5142);
and U6334 (N_6334,N_5957,N_5344);
and U6335 (N_6335,N_5574,N_5460);
or U6336 (N_6336,N_5912,N_5001);
nand U6337 (N_6337,N_5805,N_5685);
and U6338 (N_6338,N_5060,N_5478);
or U6339 (N_6339,N_5445,N_5173);
and U6340 (N_6340,N_5213,N_5911);
nand U6341 (N_6341,N_5537,N_5297);
or U6342 (N_6342,N_5074,N_5052);
nand U6343 (N_6343,N_5028,N_5669);
and U6344 (N_6344,N_5832,N_5667);
or U6345 (N_6345,N_5058,N_5302);
and U6346 (N_6346,N_5255,N_5245);
nor U6347 (N_6347,N_5346,N_5676);
and U6348 (N_6348,N_5569,N_5559);
or U6349 (N_6349,N_5161,N_5384);
nor U6350 (N_6350,N_5509,N_5156);
nand U6351 (N_6351,N_5209,N_5165);
and U6352 (N_6352,N_5920,N_5032);
and U6353 (N_6353,N_5819,N_5396);
and U6354 (N_6354,N_5282,N_5970);
and U6355 (N_6355,N_5123,N_5022);
or U6356 (N_6356,N_5504,N_5730);
nor U6357 (N_6357,N_5003,N_5534);
nand U6358 (N_6358,N_5924,N_5373);
nor U6359 (N_6359,N_5100,N_5651);
and U6360 (N_6360,N_5698,N_5776);
or U6361 (N_6361,N_5324,N_5869);
or U6362 (N_6362,N_5525,N_5420);
nand U6363 (N_6363,N_5342,N_5535);
and U6364 (N_6364,N_5824,N_5147);
or U6365 (N_6365,N_5625,N_5826);
and U6366 (N_6366,N_5907,N_5991);
nand U6367 (N_6367,N_5315,N_5763);
nand U6368 (N_6368,N_5582,N_5640);
nand U6369 (N_6369,N_5531,N_5232);
nor U6370 (N_6370,N_5778,N_5168);
nor U6371 (N_6371,N_5380,N_5780);
nor U6372 (N_6372,N_5992,N_5867);
nand U6373 (N_6373,N_5065,N_5476);
nand U6374 (N_6374,N_5240,N_5715);
nand U6375 (N_6375,N_5871,N_5955);
nand U6376 (N_6376,N_5865,N_5049);
nor U6377 (N_6377,N_5404,N_5219);
nor U6378 (N_6378,N_5697,N_5484);
or U6379 (N_6379,N_5654,N_5520);
nor U6380 (N_6380,N_5540,N_5881);
nor U6381 (N_6381,N_5703,N_5628);
or U6382 (N_6382,N_5719,N_5563);
or U6383 (N_6383,N_5489,N_5465);
nand U6384 (N_6384,N_5590,N_5205);
and U6385 (N_6385,N_5492,N_5501);
and U6386 (N_6386,N_5548,N_5480);
and U6387 (N_6387,N_5114,N_5691);
nand U6388 (N_6388,N_5709,N_5222);
nand U6389 (N_6389,N_5170,N_5664);
nor U6390 (N_6390,N_5567,N_5334);
or U6391 (N_6391,N_5904,N_5130);
or U6392 (N_6392,N_5796,N_5036);
and U6393 (N_6393,N_5018,N_5325);
and U6394 (N_6394,N_5024,N_5259);
and U6395 (N_6395,N_5428,N_5323);
or U6396 (N_6396,N_5843,N_5689);
nand U6397 (N_6397,N_5998,N_5817);
nor U6398 (N_6398,N_5112,N_5251);
or U6399 (N_6399,N_5431,N_5211);
nor U6400 (N_6400,N_5167,N_5040);
nand U6401 (N_6401,N_5120,N_5860);
or U6402 (N_6402,N_5069,N_5300);
nor U6403 (N_6403,N_5362,N_5437);
nand U6404 (N_6404,N_5355,N_5510);
or U6405 (N_6405,N_5118,N_5002);
or U6406 (N_6406,N_5758,N_5415);
or U6407 (N_6407,N_5212,N_5745);
and U6408 (N_6408,N_5236,N_5301);
nor U6409 (N_6409,N_5777,N_5616);
nor U6410 (N_6410,N_5448,N_5652);
or U6411 (N_6411,N_5523,N_5157);
and U6412 (N_6412,N_5979,N_5830);
nand U6413 (N_6413,N_5506,N_5031);
or U6414 (N_6414,N_5903,N_5400);
nor U6415 (N_6415,N_5131,N_5227);
nor U6416 (N_6416,N_5666,N_5661);
nor U6417 (N_6417,N_5511,N_5553);
and U6418 (N_6418,N_5890,N_5426);
nor U6419 (N_6419,N_5092,N_5723);
xnor U6420 (N_6420,N_5610,N_5859);
or U6421 (N_6421,N_5934,N_5164);
nand U6422 (N_6422,N_5013,N_5027);
and U6423 (N_6423,N_5196,N_5497);
nor U6424 (N_6424,N_5148,N_5621);
nand U6425 (N_6425,N_5602,N_5889);
or U6426 (N_6426,N_5265,N_5980);
nand U6427 (N_6427,N_5743,N_5696);
nand U6428 (N_6428,N_5524,N_5735);
and U6429 (N_6429,N_5042,N_5389);
or U6430 (N_6430,N_5134,N_5633);
nor U6431 (N_6431,N_5717,N_5688);
or U6432 (N_6432,N_5794,N_5298);
nand U6433 (N_6433,N_5137,N_5226);
and U6434 (N_6434,N_5612,N_5329);
nor U6435 (N_6435,N_5043,N_5424);
and U6436 (N_6436,N_5277,N_5653);
nor U6437 (N_6437,N_5254,N_5435);
nor U6438 (N_6438,N_5968,N_5094);
and U6439 (N_6439,N_5913,N_5756);
or U6440 (N_6440,N_5496,N_5714);
or U6441 (N_6441,N_5877,N_5444);
nand U6442 (N_6442,N_5699,N_5949);
and U6443 (N_6443,N_5892,N_5403);
nor U6444 (N_6444,N_5397,N_5073);
nand U6445 (N_6445,N_5085,N_5063);
nor U6446 (N_6446,N_5356,N_5034);
nand U6447 (N_6447,N_5258,N_5880);
and U6448 (N_6448,N_5891,N_5766);
and U6449 (N_6449,N_5795,N_5182);
nor U6450 (N_6450,N_5783,N_5941);
nand U6451 (N_6451,N_5203,N_5945);
or U6452 (N_6452,N_5066,N_5269);
and U6453 (N_6453,N_5192,N_5056);
or U6454 (N_6454,N_5175,N_5677);
or U6455 (N_6455,N_5335,N_5518);
nand U6456 (N_6456,N_5187,N_5686);
nor U6457 (N_6457,N_5631,N_5359);
and U6458 (N_6458,N_5048,N_5755);
and U6459 (N_6459,N_5481,N_5782);
or U6460 (N_6460,N_5008,N_5601);
nand U6461 (N_6461,N_5235,N_5145);
and U6462 (N_6462,N_5821,N_5846);
nor U6463 (N_6463,N_5573,N_5005);
or U6464 (N_6464,N_5838,N_5530);
or U6465 (N_6465,N_5630,N_5051);
and U6466 (N_6466,N_5495,N_5643);
and U6467 (N_6467,N_5443,N_5129);
nor U6468 (N_6468,N_5954,N_5842);
nor U6469 (N_6469,N_5554,N_5581);
or U6470 (N_6470,N_5252,N_5747);
and U6471 (N_6471,N_5961,N_5527);
nand U6472 (N_6472,N_5292,N_5321);
and U6473 (N_6473,N_5214,N_5200);
and U6474 (N_6474,N_5225,N_5543);
nand U6475 (N_6475,N_5873,N_5929);
and U6476 (N_6476,N_5451,N_5532);
nand U6477 (N_6477,N_5935,N_5754);
nor U6478 (N_6478,N_5861,N_5577);
nor U6479 (N_6479,N_5468,N_5884);
nor U6480 (N_6480,N_5374,N_5694);
nand U6481 (N_6481,N_5879,N_5909);
nor U6482 (N_6482,N_5472,N_5988);
or U6483 (N_6483,N_5768,N_5620);
nand U6484 (N_6484,N_5705,N_5579);
or U6485 (N_6485,N_5562,N_5897);
nor U6486 (N_6486,N_5262,N_5461);
and U6487 (N_6487,N_5565,N_5313);
nand U6488 (N_6488,N_5978,N_5977);
and U6489 (N_6489,N_5299,N_5261);
and U6490 (N_6490,N_5797,N_5290);
nand U6491 (N_6491,N_5103,N_5517);
or U6492 (N_6492,N_5791,N_5345);
nand U6493 (N_6493,N_5116,N_5249);
or U6494 (N_6494,N_5549,N_5702);
and U6495 (N_6495,N_5712,N_5391);
nand U6496 (N_6496,N_5965,N_5767);
and U6497 (N_6497,N_5765,N_5304);
nor U6498 (N_6498,N_5459,N_5682);
or U6499 (N_6499,N_5710,N_5210);
and U6500 (N_6500,N_5332,N_5670);
nand U6501 (N_6501,N_5234,N_5837);
nand U6502 (N_6502,N_5265,N_5413);
nor U6503 (N_6503,N_5747,N_5926);
and U6504 (N_6504,N_5154,N_5532);
nand U6505 (N_6505,N_5703,N_5766);
and U6506 (N_6506,N_5533,N_5250);
and U6507 (N_6507,N_5205,N_5980);
xnor U6508 (N_6508,N_5230,N_5164);
nand U6509 (N_6509,N_5144,N_5809);
or U6510 (N_6510,N_5954,N_5431);
and U6511 (N_6511,N_5863,N_5581);
or U6512 (N_6512,N_5705,N_5197);
nand U6513 (N_6513,N_5868,N_5620);
nand U6514 (N_6514,N_5218,N_5043);
or U6515 (N_6515,N_5312,N_5962);
nor U6516 (N_6516,N_5690,N_5368);
or U6517 (N_6517,N_5936,N_5205);
nor U6518 (N_6518,N_5398,N_5023);
nand U6519 (N_6519,N_5368,N_5148);
and U6520 (N_6520,N_5343,N_5570);
and U6521 (N_6521,N_5171,N_5144);
nor U6522 (N_6522,N_5953,N_5088);
nand U6523 (N_6523,N_5778,N_5551);
or U6524 (N_6524,N_5338,N_5864);
nor U6525 (N_6525,N_5456,N_5175);
nor U6526 (N_6526,N_5082,N_5778);
xor U6527 (N_6527,N_5539,N_5315);
and U6528 (N_6528,N_5577,N_5191);
and U6529 (N_6529,N_5278,N_5266);
xor U6530 (N_6530,N_5662,N_5869);
xnor U6531 (N_6531,N_5756,N_5564);
nor U6532 (N_6532,N_5476,N_5810);
or U6533 (N_6533,N_5068,N_5509);
nand U6534 (N_6534,N_5412,N_5288);
and U6535 (N_6535,N_5913,N_5626);
xnor U6536 (N_6536,N_5220,N_5960);
or U6537 (N_6537,N_5909,N_5790);
or U6538 (N_6538,N_5766,N_5572);
or U6539 (N_6539,N_5420,N_5787);
and U6540 (N_6540,N_5146,N_5644);
or U6541 (N_6541,N_5514,N_5927);
and U6542 (N_6542,N_5493,N_5363);
or U6543 (N_6543,N_5363,N_5747);
and U6544 (N_6544,N_5622,N_5223);
and U6545 (N_6545,N_5057,N_5081);
and U6546 (N_6546,N_5384,N_5737);
nor U6547 (N_6547,N_5420,N_5609);
nor U6548 (N_6548,N_5185,N_5152);
nand U6549 (N_6549,N_5283,N_5413);
nand U6550 (N_6550,N_5657,N_5373);
nand U6551 (N_6551,N_5006,N_5316);
and U6552 (N_6552,N_5330,N_5231);
nor U6553 (N_6553,N_5786,N_5094);
or U6554 (N_6554,N_5552,N_5338);
nor U6555 (N_6555,N_5204,N_5143);
or U6556 (N_6556,N_5792,N_5163);
and U6557 (N_6557,N_5837,N_5067);
nor U6558 (N_6558,N_5580,N_5674);
or U6559 (N_6559,N_5313,N_5776);
or U6560 (N_6560,N_5434,N_5888);
or U6561 (N_6561,N_5207,N_5298);
or U6562 (N_6562,N_5804,N_5998);
nand U6563 (N_6563,N_5620,N_5874);
nor U6564 (N_6564,N_5687,N_5359);
nand U6565 (N_6565,N_5214,N_5713);
nor U6566 (N_6566,N_5918,N_5816);
or U6567 (N_6567,N_5064,N_5826);
nor U6568 (N_6568,N_5747,N_5431);
nand U6569 (N_6569,N_5557,N_5796);
or U6570 (N_6570,N_5945,N_5234);
nor U6571 (N_6571,N_5013,N_5591);
and U6572 (N_6572,N_5635,N_5923);
nand U6573 (N_6573,N_5203,N_5741);
and U6574 (N_6574,N_5968,N_5306);
nor U6575 (N_6575,N_5508,N_5180);
or U6576 (N_6576,N_5165,N_5814);
or U6577 (N_6577,N_5809,N_5554);
and U6578 (N_6578,N_5400,N_5739);
nand U6579 (N_6579,N_5481,N_5283);
nand U6580 (N_6580,N_5125,N_5210);
or U6581 (N_6581,N_5936,N_5717);
and U6582 (N_6582,N_5977,N_5264);
nand U6583 (N_6583,N_5518,N_5545);
nand U6584 (N_6584,N_5750,N_5149);
and U6585 (N_6585,N_5766,N_5221);
and U6586 (N_6586,N_5935,N_5233);
nand U6587 (N_6587,N_5473,N_5863);
nand U6588 (N_6588,N_5584,N_5326);
or U6589 (N_6589,N_5668,N_5729);
and U6590 (N_6590,N_5249,N_5772);
nor U6591 (N_6591,N_5098,N_5601);
nand U6592 (N_6592,N_5731,N_5776);
nand U6593 (N_6593,N_5295,N_5883);
nand U6594 (N_6594,N_5997,N_5495);
nand U6595 (N_6595,N_5597,N_5857);
nor U6596 (N_6596,N_5645,N_5060);
and U6597 (N_6597,N_5118,N_5979);
nand U6598 (N_6598,N_5851,N_5788);
nand U6599 (N_6599,N_5029,N_5872);
xor U6600 (N_6600,N_5721,N_5211);
or U6601 (N_6601,N_5828,N_5491);
and U6602 (N_6602,N_5608,N_5200);
and U6603 (N_6603,N_5909,N_5725);
or U6604 (N_6604,N_5238,N_5963);
and U6605 (N_6605,N_5521,N_5492);
nand U6606 (N_6606,N_5238,N_5290);
and U6607 (N_6607,N_5546,N_5301);
and U6608 (N_6608,N_5720,N_5177);
nor U6609 (N_6609,N_5847,N_5014);
nand U6610 (N_6610,N_5371,N_5805);
or U6611 (N_6611,N_5669,N_5242);
and U6612 (N_6612,N_5197,N_5430);
and U6613 (N_6613,N_5463,N_5944);
nand U6614 (N_6614,N_5731,N_5924);
or U6615 (N_6615,N_5828,N_5021);
or U6616 (N_6616,N_5860,N_5593);
nand U6617 (N_6617,N_5671,N_5230);
nor U6618 (N_6618,N_5950,N_5036);
nor U6619 (N_6619,N_5956,N_5749);
and U6620 (N_6620,N_5657,N_5953);
xor U6621 (N_6621,N_5103,N_5125);
nor U6622 (N_6622,N_5715,N_5296);
nor U6623 (N_6623,N_5251,N_5447);
or U6624 (N_6624,N_5298,N_5954);
nor U6625 (N_6625,N_5312,N_5340);
or U6626 (N_6626,N_5260,N_5463);
nor U6627 (N_6627,N_5182,N_5854);
nand U6628 (N_6628,N_5935,N_5987);
nor U6629 (N_6629,N_5446,N_5267);
or U6630 (N_6630,N_5287,N_5457);
nand U6631 (N_6631,N_5553,N_5363);
and U6632 (N_6632,N_5278,N_5430);
and U6633 (N_6633,N_5269,N_5719);
and U6634 (N_6634,N_5719,N_5983);
nand U6635 (N_6635,N_5388,N_5382);
nand U6636 (N_6636,N_5670,N_5756);
and U6637 (N_6637,N_5293,N_5699);
nand U6638 (N_6638,N_5121,N_5807);
or U6639 (N_6639,N_5575,N_5813);
nand U6640 (N_6640,N_5363,N_5556);
or U6641 (N_6641,N_5157,N_5591);
and U6642 (N_6642,N_5912,N_5272);
nand U6643 (N_6643,N_5312,N_5671);
and U6644 (N_6644,N_5856,N_5442);
nand U6645 (N_6645,N_5229,N_5642);
or U6646 (N_6646,N_5844,N_5471);
and U6647 (N_6647,N_5289,N_5370);
or U6648 (N_6648,N_5882,N_5642);
nor U6649 (N_6649,N_5376,N_5692);
or U6650 (N_6650,N_5677,N_5666);
and U6651 (N_6651,N_5157,N_5840);
nor U6652 (N_6652,N_5284,N_5305);
and U6653 (N_6653,N_5688,N_5784);
nor U6654 (N_6654,N_5205,N_5658);
or U6655 (N_6655,N_5730,N_5147);
nor U6656 (N_6656,N_5535,N_5690);
nor U6657 (N_6657,N_5171,N_5009);
and U6658 (N_6658,N_5662,N_5072);
and U6659 (N_6659,N_5591,N_5860);
and U6660 (N_6660,N_5549,N_5763);
nand U6661 (N_6661,N_5161,N_5418);
and U6662 (N_6662,N_5476,N_5873);
nand U6663 (N_6663,N_5978,N_5222);
nand U6664 (N_6664,N_5456,N_5961);
and U6665 (N_6665,N_5440,N_5242);
or U6666 (N_6666,N_5757,N_5783);
or U6667 (N_6667,N_5398,N_5576);
and U6668 (N_6668,N_5586,N_5609);
xnor U6669 (N_6669,N_5561,N_5321);
nor U6670 (N_6670,N_5346,N_5237);
nor U6671 (N_6671,N_5276,N_5344);
nor U6672 (N_6672,N_5322,N_5004);
nand U6673 (N_6673,N_5810,N_5929);
nor U6674 (N_6674,N_5708,N_5575);
nor U6675 (N_6675,N_5863,N_5232);
nand U6676 (N_6676,N_5366,N_5956);
nor U6677 (N_6677,N_5289,N_5905);
and U6678 (N_6678,N_5575,N_5414);
nand U6679 (N_6679,N_5265,N_5937);
and U6680 (N_6680,N_5133,N_5719);
nor U6681 (N_6681,N_5888,N_5677);
nor U6682 (N_6682,N_5903,N_5115);
and U6683 (N_6683,N_5579,N_5343);
nor U6684 (N_6684,N_5255,N_5384);
nand U6685 (N_6685,N_5492,N_5176);
and U6686 (N_6686,N_5216,N_5405);
and U6687 (N_6687,N_5953,N_5862);
and U6688 (N_6688,N_5376,N_5287);
and U6689 (N_6689,N_5655,N_5042);
or U6690 (N_6690,N_5877,N_5491);
nor U6691 (N_6691,N_5252,N_5676);
or U6692 (N_6692,N_5137,N_5495);
and U6693 (N_6693,N_5260,N_5526);
or U6694 (N_6694,N_5586,N_5106);
nand U6695 (N_6695,N_5895,N_5292);
nand U6696 (N_6696,N_5859,N_5807);
nor U6697 (N_6697,N_5369,N_5548);
nand U6698 (N_6698,N_5915,N_5014);
or U6699 (N_6699,N_5113,N_5466);
or U6700 (N_6700,N_5186,N_5006);
nor U6701 (N_6701,N_5423,N_5480);
and U6702 (N_6702,N_5680,N_5610);
and U6703 (N_6703,N_5711,N_5302);
and U6704 (N_6704,N_5311,N_5466);
nor U6705 (N_6705,N_5588,N_5496);
or U6706 (N_6706,N_5163,N_5469);
nor U6707 (N_6707,N_5807,N_5176);
and U6708 (N_6708,N_5017,N_5003);
and U6709 (N_6709,N_5283,N_5183);
and U6710 (N_6710,N_5394,N_5723);
and U6711 (N_6711,N_5775,N_5372);
and U6712 (N_6712,N_5900,N_5836);
xnor U6713 (N_6713,N_5470,N_5895);
nor U6714 (N_6714,N_5879,N_5629);
nor U6715 (N_6715,N_5199,N_5888);
and U6716 (N_6716,N_5485,N_5972);
or U6717 (N_6717,N_5927,N_5799);
or U6718 (N_6718,N_5966,N_5531);
or U6719 (N_6719,N_5092,N_5108);
nand U6720 (N_6720,N_5423,N_5017);
nand U6721 (N_6721,N_5348,N_5278);
nand U6722 (N_6722,N_5898,N_5298);
nor U6723 (N_6723,N_5923,N_5097);
nor U6724 (N_6724,N_5228,N_5068);
or U6725 (N_6725,N_5688,N_5202);
nor U6726 (N_6726,N_5993,N_5614);
nand U6727 (N_6727,N_5599,N_5445);
or U6728 (N_6728,N_5766,N_5362);
or U6729 (N_6729,N_5526,N_5515);
nor U6730 (N_6730,N_5939,N_5682);
nand U6731 (N_6731,N_5781,N_5378);
or U6732 (N_6732,N_5269,N_5372);
and U6733 (N_6733,N_5228,N_5852);
nand U6734 (N_6734,N_5310,N_5204);
nor U6735 (N_6735,N_5282,N_5226);
or U6736 (N_6736,N_5582,N_5801);
and U6737 (N_6737,N_5060,N_5157);
or U6738 (N_6738,N_5396,N_5718);
nand U6739 (N_6739,N_5795,N_5523);
nor U6740 (N_6740,N_5619,N_5996);
and U6741 (N_6741,N_5462,N_5714);
and U6742 (N_6742,N_5434,N_5551);
and U6743 (N_6743,N_5307,N_5081);
and U6744 (N_6744,N_5792,N_5667);
or U6745 (N_6745,N_5778,N_5457);
or U6746 (N_6746,N_5637,N_5902);
nand U6747 (N_6747,N_5587,N_5195);
nand U6748 (N_6748,N_5183,N_5905);
nor U6749 (N_6749,N_5970,N_5867);
and U6750 (N_6750,N_5542,N_5513);
and U6751 (N_6751,N_5964,N_5751);
nand U6752 (N_6752,N_5280,N_5909);
nand U6753 (N_6753,N_5305,N_5861);
nor U6754 (N_6754,N_5655,N_5623);
nor U6755 (N_6755,N_5164,N_5937);
and U6756 (N_6756,N_5336,N_5311);
or U6757 (N_6757,N_5685,N_5981);
and U6758 (N_6758,N_5438,N_5405);
and U6759 (N_6759,N_5257,N_5388);
and U6760 (N_6760,N_5936,N_5167);
or U6761 (N_6761,N_5723,N_5594);
nand U6762 (N_6762,N_5281,N_5417);
xnor U6763 (N_6763,N_5947,N_5520);
and U6764 (N_6764,N_5696,N_5387);
and U6765 (N_6765,N_5134,N_5316);
or U6766 (N_6766,N_5686,N_5669);
or U6767 (N_6767,N_5358,N_5530);
nor U6768 (N_6768,N_5240,N_5462);
nor U6769 (N_6769,N_5949,N_5698);
nand U6770 (N_6770,N_5435,N_5154);
nand U6771 (N_6771,N_5910,N_5060);
nand U6772 (N_6772,N_5779,N_5726);
nor U6773 (N_6773,N_5784,N_5110);
and U6774 (N_6774,N_5841,N_5460);
nand U6775 (N_6775,N_5941,N_5986);
and U6776 (N_6776,N_5429,N_5239);
or U6777 (N_6777,N_5564,N_5057);
and U6778 (N_6778,N_5088,N_5346);
nor U6779 (N_6779,N_5914,N_5808);
nor U6780 (N_6780,N_5272,N_5309);
nor U6781 (N_6781,N_5842,N_5653);
or U6782 (N_6782,N_5364,N_5745);
nor U6783 (N_6783,N_5601,N_5605);
nor U6784 (N_6784,N_5796,N_5620);
nor U6785 (N_6785,N_5684,N_5075);
or U6786 (N_6786,N_5364,N_5309);
nand U6787 (N_6787,N_5360,N_5257);
nand U6788 (N_6788,N_5144,N_5413);
nand U6789 (N_6789,N_5191,N_5844);
xor U6790 (N_6790,N_5715,N_5845);
and U6791 (N_6791,N_5698,N_5126);
nand U6792 (N_6792,N_5734,N_5678);
and U6793 (N_6793,N_5776,N_5330);
nor U6794 (N_6794,N_5097,N_5708);
and U6795 (N_6795,N_5023,N_5288);
nand U6796 (N_6796,N_5402,N_5963);
nor U6797 (N_6797,N_5519,N_5092);
and U6798 (N_6798,N_5397,N_5213);
nor U6799 (N_6799,N_5765,N_5008);
nor U6800 (N_6800,N_5126,N_5936);
and U6801 (N_6801,N_5798,N_5787);
nand U6802 (N_6802,N_5586,N_5590);
nand U6803 (N_6803,N_5909,N_5101);
or U6804 (N_6804,N_5223,N_5913);
nand U6805 (N_6805,N_5035,N_5355);
or U6806 (N_6806,N_5716,N_5259);
and U6807 (N_6807,N_5577,N_5215);
nand U6808 (N_6808,N_5507,N_5317);
nor U6809 (N_6809,N_5000,N_5983);
nor U6810 (N_6810,N_5185,N_5111);
nor U6811 (N_6811,N_5857,N_5559);
nand U6812 (N_6812,N_5279,N_5321);
and U6813 (N_6813,N_5030,N_5906);
nor U6814 (N_6814,N_5971,N_5275);
or U6815 (N_6815,N_5382,N_5688);
nand U6816 (N_6816,N_5066,N_5671);
or U6817 (N_6817,N_5476,N_5516);
nor U6818 (N_6818,N_5894,N_5455);
nand U6819 (N_6819,N_5634,N_5821);
or U6820 (N_6820,N_5599,N_5894);
nor U6821 (N_6821,N_5487,N_5149);
or U6822 (N_6822,N_5089,N_5136);
and U6823 (N_6823,N_5267,N_5214);
nor U6824 (N_6824,N_5125,N_5908);
nand U6825 (N_6825,N_5221,N_5495);
nand U6826 (N_6826,N_5035,N_5379);
nor U6827 (N_6827,N_5766,N_5504);
or U6828 (N_6828,N_5311,N_5160);
xnor U6829 (N_6829,N_5681,N_5405);
and U6830 (N_6830,N_5325,N_5227);
and U6831 (N_6831,N_5699,N_5925);
or U6832 (N_6832,N_5857,N_5232);
and U6833 (N_6833,N_5476,N_5767);
nand U6834 (N_6834,N_5355,N_5761);
nand U6835 (N_6835,N_5588,N_5961);
and U6836 (N_6836,N_5788,N_5689);
nand U6837 (N_6837,N_5917,N_5651);
nand U6838 (N_6838,N_5605,N_5655);
or U6839 (N_6839,N_5937,N_5960);
or U6840 (N_6840,N_5364,N_5647);
nor U6841 (N_6841,N_5467,N_5352);
xor U6842 (N_6842,N_5493,N_5642);
nor U6843 (N_6843,N_5082,N_5263);
nor U6844 (N_6844,N_5498,N_5574);
or U6845 (N_6845,N_5633,N_5503);
nor U6846 (N_6846,N_5306,N_5315);
and U6847 (N_6847,N_5840,N_5943);
nand U6848 (N_6848,N_5455,N_5247);
and U6849 (N_6849,N_5051,N_5110);
or U6850 (N_6850,N_5379,N_5549);
and U6851 (N_6851,N_5392,N_5944);
nand U6852 (N_6852,N_5953,N_5892);
and U6853 (N_6853,N_5497,N_5264);
nand U6854 (N_6854,N_5305,N_5699);
nand U6855 (N_6855,N_5265,N_5241);
or U6856 (N_6856,N_5164,N_5196);
or U6857 (N_6857,N_5232,N_5777);
nor U6858 (N_6858,N_5132,N_5150);
or U6859 (N_6859,N_5660,N_5912);
nand U6860 (N_6860,N_5713,N_5194);
nand U6861 (N_6861,N_5562,N_5795);
nand U6862 (N_6862,N_5899,N_5774);
and U6863 (N_6863,N_5458,N_5513);
and U6864 (N_6864,N_5390,N_5879);
nand U6865 (N_6865,N_5964,N_5314);
and U6866 (N_6866,N_5156,N_5784);
nand U6867 (N_6867,N_5126,N_5498);
nand U6868 (N_6868,N_5808,N_5766);
or U6869 (N_6869,N_5118,N_5397);
and U6870 (N_6870,N_5297,N_5538);
nand U6871 (N_6871,N_5377,N_5200);
nor U6872 (N_6872,N_5036,N_5593);
and U6873 (N_6873,N_5467,N_5707);
or U6874 (N_6874,N_5763,N_5985);
or U6875 (N_6875,N_5483,N_5867);
nor U6876 (N_6876,N_5955,N_5200);
or U6877 (N_6877,N_5010,N_5312);
nor U6878 (N_6878,N_5241,N_5133);
nand U6879 (N_6879,N_5730,N_5124);
and U6880 (N_6880,N_5707,N_5217);
nand U6881 (N_6881,N_5369,N_5441);
nor U6882 (N_6882,N_5087,N_5701);
nor U6883 (N_6883,N_5087,N_5638);
nor U6884 (N_6884,N_5051,N_5964);
and U6885 (N_6885,N_5133,N_5608);
and U6886 (N_6886,N_5228,N_5049);
nor U6887 (N_6887,N_5985,N_5337);
nor U6888 (N_6888,N_5876,N_5653);
nand U6889 (N_6889,N_5715,N_5449);
and U6890 (N_6890,N_5026,N_5655);
nor U6891 (N_6891,N_5312,N_5807);
and U6892 (N_6892,N_5794,N_5397);
nand U6893 (N_6893,N_5326,N_5525);
nand U6894 (N_6894,N_5668,N_5890);
or U6895 (N_6895,N_5356,N_5277);
and U6896 (N_6896,N_5254,N_5881);
or U6897 (N_6897,N_5635,N_5644);
or U6898 (N_6898,N_5091,N_5999);
and U6899 (N_6899,N_5765,N_5611);
and U6900 (N_6900,N_5759,N_5377);
and U6901 (N_6901,N_5267,N_5516);
or U6902 (N_6902,N_5867,N_5780);
nand U6903 (N_6903,N_5389,N_5832);
or U6904 (N_6904,N_5100,N_5623);
and U6905 (N_6905,N_5534,N_5260);
and U6906 (N_6906,N_5143,N_5408);
and U6907 (N_6907,N_5894,N_5218);
or U6908 (N_6908,N_5285,N_5949);
and U6909 (N_6909,N_5297,N_5755);
and U6910 (N_6910,N_5057,N_5339);
or U6911 (N_6911,N_5302,N_5017);
or U6912 (N_6912,N_5867,N_5354);
nand U6913 (N_6913,N_5201,N_5965);
nor U6914 (N_6914,N_5606,N_5856);
nor U6915 (N_6915,N_5558,N_5505);
xor U6916 (N_6916,N_5771,N_5612);
nand U6917 (N_6917,N_5206,N_5001);
nor U6918 (N_6918,N_5553,N_5420);
nor U6919 (N_6919,N_5147,N_5669);
nor U6920 (N_6920,N_5021,N_5142);
nand U6921 (N_6921,N_5485,N_5667);
nand U6922 (N_6922,N_5596,N_5119);
nand U6923 (N_6923,N_5541,N_5643);
nand U6924 (N_6924,N_5111,N_5184);
nand U6925 (N_6925,N_5545,N_5141);
nand U6926 (N_6926,N_5106,N_5516);
or U6927 (N_6927,N_5282,N_5275);
nor U6928 (N_6928,N_5706,N_5018);
or U6929 (N_6929,N_5953,N_5357);
or U6930 (N_6930,N_5934,N_5492);
nand U6931 (N_6931,N_5617,N_5760);
nand U6932 (N_6932,N_5756,N_5434);
or U6933 (N_6933,N_5734,N_5390);
and U6934 (N_6934,N_5979,N_5720);
or U6935 (N_6935,N_5863,N_5340);
or U6936 (N_6936,N_5148,N_5142);
nand U6937 (N_6937,N_5754,N_5583);
nor U6938 (N_6938,N_5584,N_5836);
or U6939 (N_6939,N_5237,N_5582);
and U6940 (N_6940,N_5623,N_5964);
or U6941 (N_6941,N_5169,N_5109);
and U6942 (N_6942,N_5013,N_5283);
and U6943 (N_6943,N_5388,N_5264);
nand U6944 (N_6944,N_5115,N_5937);
nand U6945 (N_6945,N_5658,N_5725);
and U6946 (N_6946,N_5638,N_5860);
or U6947 (N_6947,N_5377,N_5786);
and U6948 (N_6948,N_5668,N_5922);
and U6949 (N_6949,N_5075,N_5377);
or U6950 (N_6950,N_5115,N_5530);
and U6951 (N_6951,N_5658,N_5898);
nor U6952 (N_6952,N_5947,N_5558);
or U6953 (N_6953,N_5930,N_5987);
and U6954 (N_6954,N_5401,N_5726);
nor U6955 (N_6955,N_5409,N_5540);
nand U6956 (N_6956,N_5424,N_5114);
nor U6957 (N_6957,N_5490,N_5917);
and U6958 (N_6958,N_5183,N_5107);
xor U6959 (N_6959,N_5233,N_5469);
or U6960 (N_6960,N_5823,N_5712);
nand U6961 (N_6961,N_5615,N_5873);
and U6962 (N_6962,N_5407,N_5987);
or U6963 (N_6963,N_5915,N_5174);
or U6964 (N_6964,N_5431,N_5840);
and U6965 (N_6965,N_5507,N_5368);
nor U6966 (N_6966,N_5001,N_5036);
nand U6967 (N_6967,N_5757,N_5370);
or U6968 (N_6968,N_5003,N_5396);
nand U6969 (N_6969,N_5989,N_5617);
and U6970 (N_6970,N_5462,N_5097);
or U6971 (N_6971,N_5174,N_5236);
or U6972 (N_6972,N_5296,N_5331);
or U6973 (N_6973,N_5366,N_5578);
and U6974 (N_6974,N_5544,N_5207);
or U6975 (N_6975,N_5756,N_5910);
nor U6976 (N_6976,N_5753,N_5426);
nand U6977 (N_6977,N_5624,N_5758);
or U6978 (N_6978,N_5693,N_5600);
and U6979 (N_6979,N_5872,N_5998);
and U6980 (N_6980,N_5195,N_5396);
nand U6981 (N_6981,N_5233,N_5642);
nor U6982 (N_6982,N_5560,N_5323);
nand U6983 (N_6983,N_5535,N_5050);
nand U6984 (N_6984,N_5487,N_5754);
or U6985 (N_6985,N_5947,N_5799);
nor U6986 (N_6986,N_5271,N_5418);
or U6987 (N_6987,N_5118,N_5675);
and U6988 (N_6988,N_5888,N_5080);
nand U6989 (N_6989,N_5478,N_5350);
or U6990 (N_6990,N_5575,N_5875);
and U6991 (N_6991,N_5208,N_5964);
nor U6992 (N_6992,N_5826,N_5854);
nand U6993 (N_6993,N_5475,N_5344);
and U6994 (N_6994,N_5150,N_5462);
nand U6995 (N_6995,N_5056,N_5352);
or U6996 (N_6996,N_5763,N_5744);
and U6997 (N_6997,N_5754,N_5206);
or U6998 (N_6998,N_5727,N_5126);
nand U6999 (N_6999,N_5261,N_5846);
and U7000 (N_7000,N_6448,N_6904);
nor U7001 (N_7001,N_6557,N_6895);
nand U7002 (N_7002,N_6650,N_6391);
nand U7003 (N_7003,N_6819,N_6174);
or U7004 (N_7004,N_6794,N_6258);
and U7005 (N_7005,N_6899,N_6333);
nor U7006 (N_7006,N_6042,N_6300);
or U7007 (N_7007,N_6327,N_6640);
nand U7008 (N_7008,N_6198,N_6137);
nor U7009 (N_7009,N_6499,N_6750);
or U7010 (N_7010,N_6175,N_6921);
nor U7011 (N_7011,N_6562,N_6338);
nor U7012 (N_7012,N_6411,N_6808);
or U7013 (N_7013,N_6454,N_6044);
nand U7014 (N_7014,N_6236,N_6207);
or U7015 (N_7015,N_6951,N_6491);
or U7016 (N_7016,N_6708,N_6076);
or U7017 (N_7017,N_6464,N_6032);
nor U7018 (N_7018,N_6512,N_6288);
or U7019 (N_7019,N_6960,N_6201);
nand U7020 (N_7020,N_6219,N_6609);
nor U7021 (N_7021,N_6273,N_6013);
nand U7022 (N_7022,N_6551,N_6526);
nand U7023 (N_7023,N_6954,N_6837);
nor U7024 (N_7024,N_6395,N_6296);
nand U7025 (N_7025,N_6800,N_6286);
and U7026 (N_7026,N_6058,N_6432);
nand U7027 (N_7027,N_6340,N_6636);
nor U7028 (N_7028,N_6048,N_6759);
or U7029 (N_7029,N_6374,N_6457);
or U7030 (N_7030,N_6756,N_6582);
nor U7031 (N_7031,N_6572,N_6618);
and U7032 (N_7032,N_6278,N_6758);
xor U7033 (N_7033,N_6888,N_6369);
or U7034 (N_7034,N_6194,N_6620);
and U7035 (N_7035,N_6823,N_6372);
and U7036 (N_7036,N_6285,N_6178);
nand U7037 (N_7037,N_6601,N_6703);
nand U7038 (N_7038,N_6264,N_6927);
or U7039 (N_7039,N_6687,N_6188);
nand U7040 (N_7040,N_6295,N_6145);
or U7041 (N_7041,N_6734,N_6041);
or U7042 (N_7042,N_6458,N_6973);
or U7043 (N_7043,N_6284,N_6302);
nor U7044 (N_7044,N_6509,N_6698);
nand U7045 (N_7045,N_6939,N_6580);
or U7046 (N_7046,N_6518,N_6337);
and U7047 (N_7047,N_6057,N_6078);
nor U7048 (N_7048,N_6321,N_6896);
nor U7049 (N_7049,N_6067,N_6999);
and U7050 (N_7050,N_6567,N_6481);
nor U7051 (N_7051,N_6928,N_6073);
and U7052 (N_7052,N_6543,N_6328);
and U7053 (N_7053,N_6747,N_6035);
nor U7054 (N_7054,N_6453,N_6757);
nand U7055 (N_7055,N_6574,N_6094);
nand U7056 (N_7056,N_6045,N_6473);
nand U7057 (N_7057,N_6393,N_6246);
nor U7058 (N_7058,N_6446,N_6981);
nor U7059 (N_7059,N_6664,N_6922);
nor U7060 (N_7060,N_6782,N_6743);
or U7061 (N_7061,N_6280,N_6694);
or U7062 (N_7062,N_6052,N_6441);
nand U7063 (N_7063,N_6677,N_6482);
nor U7064 (N_7064,N_6005,N_6886);
nor U7065 (N_7065,N_6524,N_6406);
nand U7066 (N_7066,N_6519,N_6608);
nand U7067 (N_7067,N_6034,N_6294);
nand U7068 (N_7068,N_6874,N_6623);
nor U7069 (N_7069,N_6478,N_6730);
and U7070 (N_7070,N_6820,N_6413);
and U7071 (N_7071,N_6081,N_6143);
or U7072 (N_7072,N_6845,N_6495);
nand U7073 (N_7073,N_6365,N_6191);
nand U7074 (N_7074,N_6082,N_6079);
or U7075 (N_7075,N_6517,N_6317);
nand U7076 (N_7076,N_6434,N_6788);
nor U7077 (N_7077,N_6607,N_6549);
nand U7078 (N_7078,N_6570,N_6459);
and U7079 (N_7079,N_6087,N_6063);
and U7080 (N_7080,N_6371,N_6712);
nor U7081 (N_7081,N_6069,N_6672);
and U7082 (N_7082,N_6479,N_6293);
nand U7083 (N_7083,N_6646,N_6537);
nand U7084 (N_7084,N_6203,N_6304);
nand U7085 (N_7085,N_6552,N_6150);
or U7086 (N_7086,N_6802,N_6477);
or U7087 (N_7087,N_6059,N_6168);
nand U7088 (N_7088,N_6653,N_6056);
nand U7089 (N_7089,N_6472,N_6050);
nor U7090 (N_7090,N_6615,N_6866);
nor U7091 (N_7091,N_6471,N_6726);
nor U7092 (N_7092,N_6436,N_6941);
nand U7093 (N_7093,N_6792,N_6637);
nand U7094 (N_7094,N_6129,N_6256);
or U7095 (N_7095,N_6313,N_6786);
and U7096 (N_7096,N_6148,N_6844);
nor U7097 (N_7097,N_6311,N_6772);
nand U7098 (N_7098,N_6652,N_6947);
or U7099 (N_7099,N_6153,N_6513);
nand U7100 (N_7100,N_6323,N_6658);
and U7101 (N_7101,N_6944,N_6959);
and U7102 (N_7102,N_6504,N_6754);
or U7103 (N_7103,N_6775,N_6815);
and U7104 (N_7104,N_6319,N_6269);
and U7105 (N_7105,N_6848,N_6039);
nand U7106 (N_7106,N_6813,N_6696);
or U7107 (N_7107,N_6669,N_6538);
nor U7108 (N_7108,N_6809,N_6115);
nor U7109 (N_7109,N_6430,N_6165);
or U7110 (N_7110,N_6200,N_6721);
or U7111 (N_7111,N_6749,N_6354);
and U7112 (N_7112,N_6793,N_6437);
nor U7113 (N_7113,N_6399,N_6351);
or U7114 (N_7114,N_6155,N_6209);
or U7115 (N_7115,N_6587,N_6334);
nor U7116 (N_7116,N_6826,N_6007);
nand U7117 (N_7117,N_6455,N_6578);
or U7118 (N_7118,N_6733,N_6723);
nor U7119 (N_7119,N_6893,N_6841);
or U7120 (N_7120,N_6325,N_6979);
nor U7121 (N_7121,N_6215,N_6010);
and U7122 (N_7122,N_6225,N_6752);
nor U7123 (N_7123,N_6289,N_6767);
or U7124 (N_7124,N_6428,N_6342);
nand U7125 (N_7125,N_6142,N_6693);
nand U7126 (N_7126,N_6424,N_6965);
nand U7127 (N_7127,N_6638,N_6425);
and U7128 (N_7128,N_6860,N_6626);
or U7129 (N_7129,N_6508,N_6345);
and U7130 (N_7130,N_6510,N_6952);
nor U7131 (N_7131,N_6942,N_6261);
nor U7132 (N_7132,N_6544,N_6421);
and U7133 (N_7133,N_6697,N_6741);
or U7134 (N_7134,N_6326,N_6803);
nor U7135 (N_7135,N_6656,N_6167);
nand U7136 (N_7136,N_6072,N_6484);
and U7137 (N_7137,N_6908,N_6659);
nor U7138 (N_7138,N_6503,N_6379);
nor U7139 (N_7139,N_6925,N_6465);
and U7140 (N_7140,N_6276,N_6883);
or U7141 (N_7141,N_6777,N_6456);
nor U7142 (N_7142,N_6346,N_6699);
and U7143 (N_7143,N_6984,N_6382);
and U7144 (N_7144,N_6085,N_6426);
nor U7145 (N_7145,N_6830,N_6972);
nand U7146 (N_7146,N_6604,N_6239);
nand U7147 (N_7147,N_6870,N_6834);
nand U7148 (N_7148,N_6462,N_6431);
nand U7149 (N_7149,N_6114,N_6080);
nor U7150 (N_7150,N_6595,N_6935);
and U7151 (N_7151,N_6903,N_6689);
and U7152 (N_7152,N_6681,N_6980);
or U7153 (N_7153,N_6475,N_6166);
nand U7154 (N_7154,N_6238,N_6109);
and U7155 (N_7155,N_6711,N_6282);
nor U7156 (N_7156,N_6210,N_6695);
nand U7157 (N_7157,N_6790,N_6778);
or U7158 (N_7158,N_6255,N_6560);
and U7159 (N_7159,N_6597,N_6092);
nand U7160 (N_7160,N_6237,N_6214);
and U7161 (N_7161,N_6579,N_6546);
and U7162 (N_7162,N_6420,N_6678);
and U7163 (N_7163,N_6111,N_6516);
nand U7164 (N_7164,N_6520,N_6110);
and U7165 (N_7165,N_6611,N_6390);
and U7166 (N_7166,N_6684,N_6970);
nand U7167 (N_7167,N_6600,N_6212);
xor U7168 (N_7168,N_6071,N_6913);
nand U7169 (N_7169,N_6906,N_6344);
and U7170 (N_7170,N_6961,N_6132);
or U7171 (N_7171,N_6797,N_6829);
nand U7172 (N_7172,N_6159,N_6173);
nor U7173 (N_7173,N_6054,N_6850);
or U7174 (N_7174,N_6349,N_6522);
nand U7175 (N_7175,N_6853,N_6355);
or U7176 (N_7176,N_6134,N_6799);
nor U7177 (N_7177,N_6217,N_6907);
or U7178 (N_7178,N_6529,N_6417);
nand U7179 (N_7179,N_6969,N_6384);
nor U7180 (N_7180,N_6303,N_6176);
nand U7181 (N_7181,N_6451,N_6657);
and U7182 (N_7182,N_6226,N_6547);
and U7183 (N_7183,N_6314,N_6014);
nor U7184 (N_7184,N_6575,N_6683);
nand U7185 (N_7185,N_6704,N_6271);
nor U7186 (N_7186,N_6884,N_6305);
nand U7187 (N_7187,N_6184,N_6483);
nor U7188 (N_7188,N_6352,N_6070);
nand U7189 (N_7189,N_6610,N_6877);
and U7190 (N_7190,N_6192,N_6616);
or U7191 (N_7191,N_6397,N_6389);
nor U7192 (N_7192,N_6910,N_6242);
nand U7193 (N_7193,N_6388,N_6131);
xor U7194 (N_7194,N_6360,N_6842);
and U7195 (N_7195,N_6283,N_6891);
nor U7196 (N_7196,N_6967,N_6894);
nand U7197 (N_7197,N_6555,N_6583);
nand U7198 (N_7198,N_6245,N_6233);
and U7199 (N_7199,N_6049,N_6966);
nor U7200 (N_7200,N_6368,N_6710);
and U7201 (N_7201,N_6591,N_6051);
or U7202 (N_7202,N_6008,N_6852);
nor U7203 (N_7203,N_6009,N_6875);
nand U7204 (N_7204,N_6364,N_6146);
nand U7205 (N_7205,N_6702,N_6573);
nand U7206 (N_7206,N_6385,N_6651);
nand U7207 (N_7207,N_6097,N_6862);
nor U7208 (N_7208,N_6789,N_6090);
or U7209 (N_7209,N_6851,N_6229);
xor U7210 (N_7210,N_6539,N_6106);
nor U7211 (N_7211,N_6735,N_6810);
and U7212 (N_7212,N_6938,N_6997);
nor U7213 (N_7213,N_6632,N_6639);
nor U7214 (N_7214,N_6419,N_6996);
nand U7215 (N_7215,N_6634,N_6206);
and U7216 (N_7216,N_6202,N_6152);
nand U7217 (N_7217,N_6031,N_6665);
nand U7218 (N_7218,N_6140,N_6243);
and U7219 (N_7219,N_6274,N_6729);
nand U7220 (N_7220,N_6272,N_6102);
or U7221 (N_7221,N_6622,N_6962);
nand U7222 (N_7222,N_6765,N_6377);
nand U7223 (N_7223,N_6828,N_6847);
and U7224 (N_7224,N_6164,N_6002);
nor U7225 (N_7225,N_6900,N_6182);
nor U7226 (N_7226,N_6489,N_6946);
or U7227 (N_7227,N_6507,N_6811);
nand U7228 (N_7228,N_6817,N_6692);
nor U7229 (N_7229,N_6705,N_6861);
or U7230 (N_7230,N_6400,N_6252);
xor U7231 (N_7231,N_6037,N_6287);
or U7232 (N_7232,N_6849,N_6309);
nand U7233 (N_7233,N_6737,N_6668);
or U7234 (N_7234,N_6964,N_6447);
or U7235 (N_7235,N_6548,N_6026);
or U7236 (N_7236,N_6655,N_6854);
nand U7237 (N_7237,N_6412,N_6105);
or U7238 (N_7238,N_6588,N_6727);
and U7239 (N_7239,N_6408,N_6427);
and U7240 (N_7240,N_6745,N_6599);
xnor U7241 (N_7241,N_6675,N_6511);
nor U7242 (N_7242,N_6028,N_6831);
nor U7243 (N_7243,N_6401,N_6937);
xnor U7244 (N_7244,N_6121,N_6700);
nand U7245 (N_7245,N_6450,N_6801);
or U7246 (N_7246,N_6642,N_6889);
or U7247 (N_7247,N_6248,N_6119);
and U7248 (N_7248,N_6897,N_6949);
and U7249 (N_7249,N_6171,N_6130);
nor U7250 (N_7250,N_6047,N_6929);
nor U7251 (N_7251,N_6253,N_6918);
nand U7252 (N_7252,N_6486,N_6074);
nand U7253 (N_7253,N_6440,N_6713);
and U7254 (N_7254,N_6864,N_6066);
nand U7255 (N_7255,N_6322,N_6189);
nand U7256 (N_7256,N_6924,N_6240);
nor U7257 (N_7257,N_6628,N_6738);
nor U7258 (N_7258,N_6649,N_6885);
and U7259 (N_7259,N_6033,N_6987);
nand U7260 (N_7260,N_6958,N_6840);
and U7261 (N_7261,N_6805,N_6022);
nor U7262 (N_7262,N_6186,N_6666);
or U7263 (N_7263,N_6839,N_6645);
or U7264 (N_7264,N_6162,N_6863);
and U7265 (N_7265,N_6443,N_6662);
nor U7266 (N_7266,N_6621,N_6204);
nand U7267 (N_7267,N_6157,N_6541);
nor U7268 (N_7268,N_6075,N_6108);
and U7269 (N_7269,N_6163,N_6989);
nor U7270 (N_7270,N_6916,N_6373);
nor U7271 (N_7271,N_6501,N_6263);
nor U7272 (N_7272,N_6671,N_6732);
and U7273 (N_7273,N_6625,N_6414);
nand U7274 (N_7274,N_6227,N_6631);
nor U7275 (N_7275,N_6061,N_6107);
and U7276 (N_7276,N_6310,N_6348);
nand U7277 (N_7277,N_6977,N_6976);
and U7278 (N_7278,N_6912,N_6331);
and U7279 (N_7279,N_6667,N_6843);
and U7280 (N_7280,N_6846,N_6530);
and U7281 (N_7281,N_6423,N_6633);
or U7282 (N_7282,N_6525,N_6487);
or U7283 (N_7283,N_6876,N_6480);
xnor U7284 (N_7284,N_6521,N_6301);
nand U7285 (N_7285,N_6196,N_6466);
or U7286 (N_7286,N_6857,N_6407);
nor U7287 (N_7287,N_6553,N_6991);
nor U7288 (N_7288,N_6902,N_6596);
nand U7289 (N_7289,N_6545,N_6686);
nand U7290 (N_7290,N_6773,N_6235);
and U7291 (N_7291,N_6350,N_6617);
nand U7292 (N_7292,N_6474,N_6015);
and U7293 (N_7293,N_6012,N_6011);
and U7294 (N_7294,N_6267,N_6147);
and U7295 (N_7295,N_6905,N_6807);
or U7296 (N_7296,N_6559,N_6187);
or U7297 (N_7297,N_6470,N_6298);
and U7298 (N_7298,N_6785,N_6460);
and U7299 (N_7299,N_6324,N_6376);
xnor U7300 (N_7300,N_6394,N_6485);
and U7301 (N_7301,N_6315,N_6766);
nand U7302 (N_7302,N_6139,N_6234);
or U7303 (N_7303,N_6442,N_6030);
nand U7304 (N_7304,N_6502,N_6190);
or U7305 (N_7305,N_6709,N_6880);
and U7306 (N_7306,N_6154,N_6534);
nand U7307 (N_7307,N_6835,N_6911);
nor U7308 (N_7308,N_6956,N_6536);
nand U7309 (N_7309,N_6444,N_6701);
or U7310 (N_7310,N_6763,N_6133);
or U7311 (N_7311,N_6383,N_6359);
xor U7312 (N_7312,N_6714,N_6663);
or U7313 (N_7313,N_6161,N_6361);
nor U7314 (N_7314,N_6307,N_6629);
and U7315 (N_7315,N_6685,N_6812);
or U7316 (N_7316,N_6020,N_6254);
and U7317 (N_7317,N_6216,N_6781);
and U7318 (N_7318,N_6836,N_6527);
nand U7319 (N_7319,N_6872,N_6339);
or U7320 (N_7320,N_6392,N_6585);
nor U7321 (N_7321,N_6873,N_6490);
nand U7322 (N_7322,N_6855,N_6776);
and U7323 (N_7323,N_6493,N_6197);
or U7324 (N_7324,N_6332,N_6029);
nor U7325 (N_7325,N_6532,N_6290);
nand U7326 (N_7326,N_6306,N_6593);
nor U7327 (N_7327,N_6613,N_6004);
nand U7328 (N_7328,N_6416,N_6535);
or U7329 (N_7329,N_6122,N_6463);
nand U7330 (N_7330,N_6128,N_6387);
and U7331 (N_7331,N_6433,N_6644);
nand U7332 (N_7332,N_6099,N_6318);
nand U7333 (N_7333,N_6920,N_6748);
nor U7334 (N_7334,N_6124,N_6680);
and U7335 (N_7335,N_6279,N_6795);
and U7336 (N_7336,N_6584,N_6871);
or U7337 (N_7337,N_6312,N_6151);
nand U7338 (N_7338,N_6018,N_6577);
nand U7339 (N_7339,N_6127,N_6488);
nand U7340 (N_7340,N_6898,N_6783);
or U7341 (N_7341,N_6223,N_6764);
nand U7342 (N_7342,N_6833,N_6630);
nand U7343 (N_7343,N_6859,N_6770);
nand U7344 (N_7344,N_6992,N_6222);
xnor U7345 (N_7345,N_6016,N_6569);
nor U7346 (N_7346,N_6654,N_6768);
or U7347 (N_7347,N_6403,N_6021);
xnor U7348 (N_7348,N_6716,N_6402);
nor U7349 (N_7349,N_6291,N_6558);
nor U7350 (N_7350,N_6247,N_6936);
or U7351 (N_7351,N_6230,N_6760);
nor U7352 (N_7352,N_6586,N_6919);
nor U7353 (N_7353,N_6720,N_6761);
and U7354 (N_7354,N_6780,N_6590);
nand U7355 (N_7355,N_6878,N_6358);
or U7356 (N_7356,N_6265,N_6232);
nand U7357 (N_7357,N_6292,N_6112);
and U7358 (N_7358,N_6096,N_6753);
or U7359 (N_7359,N_6329,N_6975);
nor U7360 (N_7360,N_6260,N_6429);
or U7361 (N_7361,N_6978,N_6771);
nand U7362 (N_7362,N_6341,N_6804);
or U7363 (N_7363,N_6892,N_6561);
nor U7364 (N_7364,N_6755,N_6185);
xnor U7365 (N_7365,N_6118,N_6299);
or U7366 (N_7366,N_6277,N_6605);
nor U7367 (N_7367,N_6409,N_6439);
nand U7368 (N_7368,N_6858,N_6515);
nand U7369 (N_7369,N_6158,N_6715);
nor U7370 (N_7370,N_6452,N_6869);
nor U7371 (N_7371,N_6343,N_6744);
nor U7372 (N_7372,N_6868,N_6043);
nand U7373 (N_7373,N_6335,N_6065);
nor U7374 (N_7374,N_6241,N_6691);
nand U7375 (N_7375,N_6506,N_6957);
and U7376 (N_7376,N_6062,N_6867);
nor U7377 (N_7377,N_6576,N_6103);
nand U7378 (N_7378,N_6136,N_6719);
nor U7379 (N_7379,N_6986,N_6923);
or U7380 (N_7380,N_6149,N_6213);
nand U7381 (N_7381,N_6740,N_6231);
and U7382 (N_7382,N_6948,N_6375);
or U7383 (N_7383,N_6968,N_6467);
nand U7384 (N_7384,N_6926,N_6682);
nor U7385 (N_7385,N_6492,N_6268);
and U7386 (N_7386,N_6971,N_6040);
nor U7387 (N_7387,N_6931,N_6940);
nor U7388 (N_7388,N_6281,N_6101);
nor U7389 (N_7389,N_6019,N_6707);
nor U7390 (N_7390,N_6945,N_6024);
nor U7391 (N_7391,N_6542,N_6181);
nand U7392 (N_7392,N_6676,N_6670);
nor U7393 (N_7393,N_6528,N_6554);
or U7394 (N_7394,N_6160,N_6838);
nor U7395 (N_7395,N_6498,N_6170);
nor U7396 (N_7396,N_6468,N_6422);
or U7397 (N_7397,N_6641,N_6083);
nand U7398 (N_7398,N_6932,N_6179);
and U7399 (N_7399,N_6023,N_6717);
or U7400 (N_7400,N_6086,N_6674);
nand U7401 (N_7401,N_6779,N_6901);
and U7402 (N_7402,N_6461,N_6095);
nor U7403 (N_7403,N_6386,N_6126);
nor U7404 (N_7404,N_6221,N_6762);
and U7405 (N_7405,N_6093,N_6089);
and U7406 (N_7406,N_6881,N_6827);
or U7407 (N_7407,N_6398,N_6060);
nand U7408 (N_7408,N_6523,N_6550);
or U7409 (N_7409,N_6565,N_6378);
nor U7410 (N_7410,N_6953,N_6220);
nor U7411 (N_7411,N_6228,N_6224);
or U7412 (N_7412,N_6000,N_6627);
or U7413 (N_7413,N_6088,N_6784);
nor U7414 (N_7414,N_6619,N_6330);
and U7415 (N_7415,N_6614,N_6077);
and U7416 (N_7416,N_6993,N_6262);
and U7417 (N_7417,N_6722,N_6405);
and U7418 (N_7418,N_6943,N_6816);
or U7419 (N_7419,N_6068,N_6169);
nand U7420 (N_7420,N_6915,N_6193);
xor U7421 (N_7421,N_6120,N_6728);
and U7422 (N_7422,N_6098,N_6647);
nor U7423 (N_7423,N_6690,N_6125);
nor U7424 (N_7424,N_6914,N_6249);
and U7425 (N_7425,N_6564,N_6320);
or U7426 (N_7426,N_6890,N_6381);
nand U7427 (N_7427,N_6825,N_6606);
or U7428 (N_7428,N_6602,N_6100);
or U7429 (N_7429,N_6818,N_6824);
or U7430 (N_7430,N_6724,N_6211);
nand U7431 (N_7431,N_6275,N_6046);
nand U7432 (N_7432,N_6983,N_6367);
or U7433 (N_7433,N_6438,N_6449);
or U7434 (N_7434,N_6036,N_6308);
or U7435 (N_7435,N_6259,N_6718);
or U7436 (N_7436,N_6404,N_6950);
and U7437 (N_7437,N_6806,N_6251);
nor U7438 (N_7438,N_6396,N_6661);
and U7439 (N_7439,N_6363,N_6648);
nor U7440 (N_7440,N_6144,N_6739);
nor U7441 (N_7441,N_6917,N_6598);
and U7442 (N_7442,N_6205,N_6500);
and U7443 (N_7443,N_6113,N_6116);
or U7444 (N_7444,N_6250,N_6995);
and U7445 (N_7445,N_6679,N_6183);
and U7446 (N_7446,N_6974,N_6635);
nand U7447 (N_7447,N_6603,N_6380);
and U7448 (N_7448,N_6909,N_6347);
nand U7449 (N_7449,N_6643,N_6418);
and U7450 (N_7450,N_6257,N_6370);
nor U7451 (N_7451,N_6832,N_6496);
or U7452 (N_7452,N_6415,N_6821);
nor U7453 (N_7453,N_6336,N_6985);
and U7454 (N_7454,N_6027,N_6594);
and U7455 (N_7455,N_6297,N_6366);
and U7456 (N_7456,N_6660,N_6266);
nor U7457 (N_7457,N_6963,N_6353);
nor U7458 (N_7458,N_6879,N_6791);
and U7459 (N_7459,N_6362,N_6038);
nand U7460 (N_7460,N_6017,N_6933);
and U7461 (N_7461,N_6540,N_6934);
nand U7462 (N_7462,N_6796,N_6025);
nand U7463 (N_7463,N_6822,N_6568);
and U7464 (N_7464,N_6990,N_6357);
xnor U7465 (N_7465,N_6135,N_6856);
nor U7466 (N_7466,N_6172,N_6123);
and U7467 (N_7467,N_6787,N_6494);
and U7468 (N_7468,N_6930,N_6218);
or U7469 (N_7469,N_6865,N_6180);
and U7470 (N_7470,N_6581,N_6955);
nand U7471 (N_7471,N_6497,N_6731);
nand U7472 (N_7472,N_6117,N_6988);
nor U7473 (N_7473,N_6053,N_6505);
nand U7474 (N_7474,N_6531,N_6156);
or U7475 (N_7475,N_6199,N_6688);
nand U7476 (N_7476,N_6994,N_6141);
or U7477 (N_7477,N_6091,N_6725);
and U7478 (N_7478,N_6138,N_6742);
nor U7479 (N_7479,N_6673,N_6064);
or U7480 (N_7480,N_6055,N_6556);
nand U7481 (N_7481,N_6356,N_6887);
or U7482 (N_7482,N_6982,N_6769);
and U7483 (N_7483,N_6533,N_6798);
nor U7484 (N_7484,N_6469,N_6882);
and U7485 (N_7485,N_6195,N_6514);
xnor U7486 (N_7486,N_6998,N_6706);
nor U7487 (N_7487,N_6746,N_6006);
nand U7488 (N_7488,N_6736,N_6316);
or U7489 (N_7489,N_6177,N_6566);
nor U7490 (N_7490,N_6003,N_6624);
nand U7491 (N_7491,N_6104,N_6612);
and U7492 (N_7492,N_6244,N_6563);
or U7493 (N_7493,N_6589,N_6445);
and U7494 (N_7494,N_6476,N_6410);
nor U7495 (N_7495,N_6571,N_6592);
or U7496 (N_7496,N_6751,N_6001);
nand U7497 (N_7497,N_6814,N_6435);
nor U7498 (N_7498,N_6774,N_6208);
nor U7499 (N_7499,N_6270,N_6084);
and U7500 (N_7500,N_6190,N_6013);
or U7501 (N_7501,N_6101,N_6539);
or U7502 (N_7502,N_6269,N_6023);
nor U7503 (N_7503,N_6917,N_6591);
and U7504 (N_7504,N_6055,N_6497);
nand U7505 (N_7505,N_6150,N_6886);
nand U7506 (N_7506,N_6720,N_6899);
or U7507 (N_7507,N_6528,N_6772);
and U7508 (N_7508,N_6812,N_6290);
nor U7509 (N_7509,N_6990,N_6395);
or U7510 (N_7510,N_6219,N_6848);
or U7511 (N_7511,N_6725,N_6187);
or U7512 (N_7512,N_6138,N_6893);
and U7513 (N_7513,N_6266,N_6243);
nand U7514 (N_7514,N_6917,N_6656);
or U7515 (N_7515,N_6473,N_6247);
nand U7516 (N_7516,N_6900,N_6020);
nand U7517 (N_7517,N_6597,N_6300);
and U7518 (N_7518,N_6023,N_6515);
nand U7519 (N_7519,N_6190,N_6939);
and U7520 (N_7520,N_6318,N_6257);
nand U7521 (N_7521,N_6698,N_6456);
nand U7522 (N_7522,N_6715,N_6764);
nor U7523 (N_7523,N_6825,N_6745);
or U7524 (N_7524,N_6129,N_6405);
or U7525 (N_7525,N_6294,N_6612);
and U7526 (N_7526,N_6540,N_6894);
nor U7527 (N_7527,N_6171,N_6801);
or U7528 (N_7528,N_6372,N_6102);
or U7529 (N_7529,N_6522,N_6673);
nand U7530 (N_7530,N_6986,N_6829);
and U7531 (N_7531,N_6551,N_6758);
nor U7532 (N_7532,N_6604,N_6386);
and U7533 (N_7533,N_6652,N_6512);
or U7534 (N_7534,N_6140,N_6365);
nor U7535 (N_7535,N_6922,N_6690);
or U7536 (N_7536,N_6325,N_6433);
or U7537 (N_7537,N_6154,N_6638);
or U7538 (N_7538,N_6020,N_6814);
nor U7539 (N_7539,N_6212,N_6346);
or U7540 (N_7540,N_6279,N_6811);
or U7541 (N_7541,N_6438,N_6922);
and U7542 (N_7542,N_6388,N_6404);
nor U7543 (N_7543,N_6624,N_6554);
nand U7544 (N_7544,N_6355,N_6889);
and U7545 (N_7545,N_6391,N_6464);
nor U7546 (N_7546,N_6744,N_6906);
and U7547 (N_7547,N_6973,N_6014);
or U7548 (N_7548,N_6830,N_6410);
nor U7549 (N_7549,N_6310,N_6671);
nand U7550 (N_7550,N_6438,N_6480);
and U7551 (N_7551,N_6304,N_6155);
nand U7552 (N_7552,N_6125,N_6607);
and U7553 (N_7553,N_6099,N_6634);
and U7554 (N_7554,N_6038,N_6193);
or U7555 (N_7555,N_6554,N_6492);
nand U7556 (N_7556,N_6059,N_6751);
nor U7557 (N_7557,N_6743,N_6861);
and U7558 (N_7558,N_6179,N_6027);
nand U7559 (N_7559,N_6537,N_6209);
and U7560 (N_7560,N_6992,N_6178);
nor U7561 (N_7561,N_6429,N_6711);
and U7562 (N_7562,N_6063,N_6854);
or U7563 (N_7563,N_6310,N_6747);
nor U7564 (N_7564,N_6245,N_6878);
or U7565 (N_7565,N_6630,N_6321);
nor U7566 (N_7566,N_6425,N_6967);
xor U7567 (N_7567,N_6982,N_6170);
nor U7568 (N_7568,N_6337,N_6982);
nor U7569 (N_7569,N_6835,N_6469);
or U7570 (N_7570,N_6582,N_6745);
xnor U7571 (N_7571,N_6985,N_6379);
nand U7572 (N_7572,N_6426,N_6463);
and U7573 (N_7573,N_6365,N_6707);
or U7574 (N_7574,N_6948,N_6346);
nand U7575 (N_7575,N_6606,N_6022);
nor U7576 (N_7576,N_6244,N_6236);
nand U7577 (N_7577,N_6880,N_6254);
and U7578 (N_7578,N_6074,N_6987);
and U7579 (N_7579,N_6194,N_6092);
or U7580 (N_7580,N_6323,N_6867);
nor U7581 (N_7581,N_6786,N_6631);
nand U7582 (N_7582,N_6084,N_6994);
nand U7583 (N_7583,N_6501,N_6899);
nor U7584 (N_7584,N_6795,N_6664);
or U7585 (N_7585,N_6140,N_6691);
and U7586 (N_7586,N_6426,N_6527);
or U7587 (N_7587,N_6873,N_6368);
or U7588 (N_7588,N_6688,N_6320);
nor U7589 (N_7589,N_6827,N_6012);
nand U7590 (N_7590,N_6462,N_6642);
nand U7591 (N_7591,N_6064,N_6662);
xnor U7592 (N_7592,N_6734,N_6640);
and U7593 (N_7593,N_6449,N_6659);
or U7594 (N_7594,N_6833,N_6764);
nand U7595 (N_7595,N_6458,N_6103);
and U7596 (N_7596,N_6222,N_6437);
nor U7597 (N_7597,N_6696,N_6240);
xor U7598 (N_7598,N_6560,N_6083);
or U7599 (N_7599,N_6460,N_6225);
nor U7600 (N_7600,N_6739,N_6512);
nor U7601 (N_7601,N_6697,N_6521);
and U7602 (N_7602,N_6355,N_6979);
and U7603 (N_7603,N_6320,N_6180);
nor U7604 (N_7604,N_6397,N_6379);
and U7605 (N_7605,N_6209,N_6451);
nand U7606 (N_7606,N_6248,N_6040);
or U7607 (N_7607,N_6357,N_6468);
and U7608 (N_7608,N_6634,N_6092);
nor U7609 (N_7609,N_6321,N_6373);
nand U7610 (N_7610,N_6875,N_6520);
or U7611 (N_7611,N_6965,N_6358);
or U7612 (N_7612,N_6943,N_6913);
nand U7613 (N_7613,N_6079,N_6784);
or U7614 (N_7614,N_6722,N_6205);
nor U7615 (N_7615,N_6365,N_6145);
nand U7616 (N_7616,N_6881,N_6765);
nand U7617 (N_7617,N_6547,N_6512);
and U7618 (N_7618,N_6113,N_6755);
nor U7619 (N_7619,N_6905,N_6340);
nand U7620 (N_7620,N_6097,N_6311);
or U7621 (N_7621,N_6738,N_6344);
or U7622 (N_7622,N_6036,N_6580);
and U7623 (N_7623,N_6320,N_6961);
nor U7624 (N_7624,N_6884,N_6771);
nand U7625 (N_7625,N_6998,N_6484);
or U7626 (N_7626,N_6686,N_6157);
or U7627 (N_7627,N_6033,N_6339);
nor U7628 (N_7628,N_6938,N_6794);
and U7629 (N_7629,N_6454,N_6089);
nor U7630 (N_7630,N_6523,N_6237);
and U7631 (N_7631,N_6601,N_6559);
and U7632 (N_7632,N_6655,N_6042);
and U7633 (N_7633,N_6016,N_6942);
nor U7634 (N_7634,N_6862,N_6199);
and U7635 (N_7635,N_6799,N_6329);
or U7636 (N_7636,N_6686,N_6993);
nand U7637 (N_7637,N_6588,N_6824);
nor U7638 (N_7638,N_6800,N_6081);
nor U7639 (N_7639,N_6055,N_6358);
nand U7640 (N_7640,N_6190,N_6164);
and U7641 (N_7641,N_6471,N_6495);
nand U7642 (N_7642,N_6860,N_6880);
and U7643 (N_7643,N_6209,N_6131);
nor U7644 (N_7644,N_6345,N_6383);
nor U7645 (N_7645,N_6844,N_6335);
and U7646 (N_7646,N_6663,N_6845);
nor U7647 (N_7647,N_6915,N_6537);
nor U7648 (N_7648,N_6147,N_6343);
nand U7649 (N_7649,N_6324,N_6552);
and U7650 (N_7650,N_6284,N_6356);
or U7651 (N_7651,N_6733,N_6572);
or U7652 (N_7652,N_6301,N_6262);
nand U7653 (N_7653,N_6915,N_6309);
and U7654 (N_7654,N_6085,N_6180);
nand U7655 (N_7655,N_6168,N_6558);
nand U7656 (N_7656,N_6046,N_6577);
nand U7657 (N_7657,N_6707,N_6413);
or U7658 (N_7658,N_6475,N_6886);
or U7659 (N_7659,N_6212,N_6189);
and U7660 (N_7660,N_6131,N_6995);
nand U7661 (N_7661,N_6521,N_6763);
nand U7662 (N_7662,N_6858,N_6610);
nand U7663 (N_7663,N_6807,N_6198);
nand U7664 (N_7664,N_6668,N_6764);
or U7665 (N_7665,N_6992,N_6562);
and U7666 (N_7666,N_6569,N_6436);
nor U7667 (N_7667,N_6944,N_6111);
or U7668 (N_7668,N_6587,N_6572);
nand U7669 (N_7669,N_6032,N_6358);
nor U7670 (N_7670,N_6495,N_6932);
nor U7671 (N_7671,N_6686,N_6039);
or U7672 (N_7672,N_6090,N_6157);
or U7673 (N_7673,N_6260,N_6219);
nand U7674 (N_7674,N_6734,N_6443);
nand U7675 (N_7675,N_6100,N_6469);
and U7676 (N_7676,N_6342,N_6922);
nand U7677 (N_7677,N_6679,N_6059);
nor U7678 (N_7678,N_6431,N_6929);
nand U7679 (N_7679,N_6730,N_6280);
nand U7680 (N_7680,N_6700,N_6650);
nor U7681 (N_7681,N_6503,N_6631);
or U7682 (N_7682,N_6873,N_6031);
or U7683 (N_7683,N_6022,N_6691);
nor U7684 (N_7684,N_6306,N_6237);
and U7685 (N_7685,N_6804,N_6564);
or U7686 (N_7686,N_6331,N_6310);
and U7687 (N_7687,N_6605,N_6681);
nand U7688 (N_7688,N_6722,N_6953);
and U7689 (N_7689,N_6367,N_6834);
or U7690 (N_7690,N_6003,N_6807);
or U7691 (N_7691,N_6230,N_6000);
nand U7692 (N_7692,N_6701,N_6263);
and U7693 (N_7693,N_6553,N_6459);
nor U7694 (N_7694,N_6271,N_6685);
nand U7695 (N_7695,N_6115,N_6934);
or U7696 (N_7696,N_6270,N_6316);
nor U7697 (N_7697,N_6182,N_6828);
or U7698 (N_7698,N_6589,N_6075);
and U7699 (N_7699,N_6183,N_6363);
and U7700 (N_7700,N_6562,N_6601);
nor U7701 (N_7701,N_6278,N_6315);
nor U7702 (N_7702,N_6323,N_6364);
nor U7703 (N_7703,N_6522,N_6797);
nor U7704 (N_7704,N_6093,N_6560);
nand U7705 (N_7705,N_6481,N_6253);
and U7706 (N_7706,N_6889,N_6706);
nor U7707 (N_7707,N_6112,N_6965);
nor U7708 (N_7708,N_6421,N_6902);
or U7709 (N_7709,N_6701,N_6422);
or U7710 (N_7710,N_6014,N_6901);
and U7711 (N_7711,N_6685,N_6157);
nand U7712 (N_7712,N_6781,N_6300);
and U7713 (N_7713,N_6877,N_6344);
nor U7714 (N_7714,N_6328,N_6719);
or U7715 (N_7715,N_6855,N_6247);
nand U7716 (N_7716,N_6099,N_6090);
nand U7717 (N_7717,N_6028,N_6845);
or U7718 (N_7718,N_6780,N_6517);
nor U7719 (N_7719,N_6338,N_6058);
and U7720 (N_7720,N_6632,N_6101);
nand U7721 (N_7721,N_6959,N_6520);
nor U7722 (N_7722,N_6841,N_6137);
nand U7723 (N_7723,N_6865,N_6753);
nor U7724 (N_7724,N_6207,N_6810);
nand U7725 (N_7725,N_6322,N_6383);
or U7726 (N_7726,N_6296,N_6336);
or U7727 (N_7727,N_6321,N_6831);
or U7728 (N_7728,N_6915,N_6764);
nand U7729 (N_7729,N_6971,N_6366);
and U7730 (N_7730,N_6891,N_6667);
and U7731 (N_7731,N_6161,N_6280);
and U7732 (N_7732,N_6437,N_6324);
nand U7733 (N_7733,N_6685,N_6828);
or U7734 (N_7734,N_6835,N_6956);
or U7735 (N_7735,N_6981,N_6460);
xnor U7736 (N_7736,N_6922,N_6041);
or U7737 (N_7737,N_6540,N_6761);
xnor U7738 (N_7738,N_6123,N_6388);
nor U7739 (N_7739,N_6189,N_6168);
nand U7740 (N_7740,N_6071,N_6364);
nor U7741 (N_7741,N_6781,N_6160);
nor U7742 (N_7742,N_6885,N_6402);
or U7743 (N_7743,N_6816,N_6085);
nand U7744 (N_7744,N_6894,N_6987);
and U7745 (N_7745,N_6119,N_6468);
and U7746 (N_7746,N_6115,N_6223);
and U7747 (N_7747,N_6767,N_6608);
nor U7748 (N_7748,N_6503,N_6170);
and U7749 (N_7749,N_6743,N_6703);
nor U7750 (N_7750,N_6843,N_6770);
nand U7751 (N_7751,N_6930,N_6643);
nor U7752 (N_7752,N_6119,N_6611);
nor U7753 (N_7753,N_6079,N_6967);
nand U7754 (N_7754,N_6743,N_6209);
and U7755 (N_7755,N_6464,N_6075);
nor U7756 (N_7756,N_6936,N_6792);
nand U7757 (N_7757,N_6222,N_6512);
or U7758 (N_7758,N_6372,N_6920);
and U7759 (N_7759,N_6887,N_6871);
or U7760 (N_7760,N_6239,N_6536);
nor U7761 (N_7761,N_6268,N_6871);
or U7762 (N_7762,N_6937,N_6762);
nor U7763 (N_7763,N_6581,N_6858);
nand U7764 (N_7764,N_6911,N_6158);
and U7765 (N_7765,N_6407,N_6838);
nor U7766 (N_7766,N_6366,N_6392);
nor U7767 (N_7767,N_6804,N_6587);
and U7768 (N_7768,N_6424,N_6623);
nand U7769 (N_7769,N_6279,N_6295);
or U7770 (N_7770,N_6383,N_6269);
and U7771 (N_7771,N_6596,N_6165);
nand U7772 (N_7772,N_6492,N_6363);
or U7773 (N_7773,N_6706,N_6436);
or U7774 (N_7774,N_6844,N_6265);
nor U7775 (N_7775,N_6060,N_6259);
nor U7776 (N_7776,N_6988,N_6652);
and U7777 (N_7777,N_6361,N_6314);
nand U7778 (N_7778,N_6101,N_6028);
nand U7779 (N_7779,N_6520,N_6249);
nor U7780 (N_7780,N_6060,N_6062);
and U7781 (N_7781,N_6851,N_6863);
or U7782 (N_7782,N_6763,N_6442);
and U7783 (N_7783,N_6774,N_6575);
or U7784 (N_7784,N_6237,N_6561);
or U7785 (N_7785,N_6226,N_6248);
and U7786 (N_7786,N_6900,N_6259);
and U7787 (N_7787,N_6782,N_6769);
and U7788 (N_7788,N_6200,N_6404);
nor U7789 (N_7789,N_6754,N_6053);
and U7790 (N_7790,N_6175,N_6207);
nand U7791 (N_7791,N_6662,N_6938);
nor U7792 (N_7792,N_6340,N_6985);
nor U7793 (N_7793,N_6560,N_6233);
nand U7794 (N_7794,N_6627,N_6066);
nand U7795 (N_7795,N_6736,N_6145);
nand U7796 (N_7796,N_6411,N_6123);
xnor U7797 (N_7797,N_6785,N_6999);
nor U7798 (N_7798,N_6386,N_6240);
and U7799 (N_7799,N_6918,N_6503);
or U7800 (N_7800,N_6942,N_6287);
nor U7801 (N_7801,N_6615,N_6127);
and U7802 (N_7802,N_6234,N_6230);
or U7803 (N_7803,N_6569,N_6885);
or U7804 (N_7804,N_6669,N_6942);
nor U7805 (N_7805,N_6554,N_6116);
nand U7806 (N_7806,N_6077,N_6957);
nand U7807 (N_7807,N_6712,N_6160);
or U7808 (N_7808,N_6146,N_6944);
nand U7809 (N_7809,N_6016,N_6209);
or U7810 (N_7810,N_6329,N_6167);
nand U7811 (N_7811,N_6536,N_6173);
nand U7812 (N_7812,N_6599,N_6261);
nor U7813 (N_7813,N_6413,N_6608);
nand U7814 (N_7814,N_6075,N_6729);
nor U7815 (N_7815,N_6373,N_6779);
nand U7816 (N_7816,N_6478,N_6785);
nor U7817 (N_7817,N_6701,N_6656);
nand U7818 (N_7818,N_6774,N_6471);
nor U7819 (N_7819,N_6089,N_6534);
or U7820 (N_7820,N_6306,N_6997);
or U7821 (N_7821,N_6562,N_6994);
nand U7822 (N_7822,N_6789,N_6415);
and U7823 (N_7823,N_6054,N_6219);
and U7824 (N_7824,N_6368,N_6417);
or U7825 (N_7825,N_6137,N_6800);
nor U7826 (N_7826,N_6244,N_6707);
or U7827 (N_7827,N_6704,N_6431);
or U7828 (N_7828,N_6255,N_6616);
and U7829 (N_7829,N_6857,N_6182);
nor U7830 (N_7830,N_6570,N_6684);
nor U7831 (N_7831,N_6691,N_6579);
nand U7832 (N_7832,N_6730,N_6110);
or U7833 (N_7833,N_6888,N_6230);
nand U7834 (N_7834,N_6953,N_6474);
and U7835 (N_7835,N_6363,N_6140);
nand U7836 (N_7836,N_6223,N_6212);
or U7837 (N_7837,N_6422,N_6718);
nand U7838 (N_7838,N_6847,N_6435);
nand U7839 (N_7839,N_6547,N_6626);
or U7840 (N_7840,N_6307,N_6021);
nor U7841 (N_7841,N_6451,N_6536);
nand U7842 (N_7842,N_6272,N_6062);
or U7843 (N_7843,N_6116,N_6697);
and U7844 (N_7844,N_6748,N_6925);
or U7845 (N_7845,N_6369,N_6178);
and U7846 (N_7846,N_6799,N_6770);
nor U7847 (N_7847,N_6667,N_6409);
or U7848 (N_7848,N_6974,N_6594);
nor U7849 (N_7849,N_6377,N_6000);
or U7850 (N_7850,N_6933,N_6290);
nor U7851 (N_7851,N_6488,N_6332);
nor U7852 (N_7852,N_6714,N_6428);
or U7853 (N_7853,N_6707,N_6406);
nand U7854 (N_7854,N_6017,N_6743);
nor U7855 (N_7855,N_6970,N_6253);
nor U7856 (N_7856,N_6392,N_6295);
or U7857 (N_7857,N_6384,N_6142);
nand U7858 (N_7858,N_6915,N_6175);
nand U7859 (N_7859,N_6064,N_6922);
and U7860 (N_7860,N_6398,N_6647);
and U7861 (N_7861,N_6554,N_6060);
nor U7862 (N_7862,N_6507,N_6499);
and U7863 (N_7863,N_6369,N_6527);
and U7864 (N_7864,N_6262,N_6433);
nor U7865 (N_7865,N_6126,N_6892);
and U7866 (N_7866,N_6932,N_6734);
or U7867 (N_7867,N_6047,N_6488);
nor U7868 (N_7868,N_6650,N_6172);
nor U7869 (N_7869,N_6193,N_6513);
or U7870 (N_7870,N_6239,N_6240);
nand U7871 (N_7871,N_6598,N_6371);
nor U7872 (N_7872,N_6110,N_6857);
nor U7873 (N_7873,N_6860,N_6029);
nand U7874 (N_7874,N_6600,N_6614);
and U7875 (N_7875,N_6229,N_6601);
or U7876 (N_7876,N_6839,N_6924);
nor U7877 (N_7877,N_6615,N_6376);
or U7878 (N_7878,N_6754,N_6748);
nor U7879 (N_7879,N_6438,N_6692);
nand U7880 (N_7880,N_6939,N_6159);
nor U7881 (N_7881,N_6434,N_6601);
nor U7882 (N_7882,N_6866,N_6232);
or U7883 (N_7883,N_6673,N_6302);
nand U7884 (N_7884,N_6943,N_6042);
nor U7885 (N_7885,N_6074,N_6468);
nor U7886 (N_7886,N_6839,N_6497);
xnor U7887 (N_7887,N_6401,N_6319);
nand U7888 (N_7888,N_6164,N_6564);
and U7889 (N_7889,N_6666,N_6758);
nand U7890 (N_7890,N_6038,N_6647);
nor U7891 (N_7891,N_6172,N_6319);
and U7892 (N_7892,N_6586,N_6760);
nor U7893 (N_7893,N_6548,N_6107);
and U7894 (N_7894,N_6012,N_6448);
and U7895 (N_7895,N_6299,N_6920);
nand U7896 (N_7896,N_6080,N_6201);
nand U7897 (N_7897,N_6647,N_6547);
nor U7898 (N_7898,N_6883,N_6110);
nor U7899 (N_7899,N_6660,N_6421);
or U7900 (N_7900,N_6659,N_6328);
nor U7901 (N_7901,N_6563,N_6250);
or U7902 (N_7902,N_6095,N_6751);
or U7903 (N_7903,N_6128,N_6263);
and U7904 (N_7904,N_6210,N_6039);
nand U7905 (N_7905,N_6678,N_6954);
or U7906 (N_7906,N_6811,N_6938);
nand U7907 (N_7907,N_6571,N_6208);
nand U7908 (N_7908,N_6843,N_6574);
nor U7909 (N_7909,N_6141,N_6400);
or U7910 (N_7910,N_6526,N_6079);
or U7911 (N_7911,N_6753,N_6790);
and U7912 (N_7912,N_6689,N_6442);
nand U7913 (N_7913,N_6188,N_6926);
or U7914 (N_7914,N_6506,N_6766);
or U7915 (N_7915,N_6554,N_6093);
nand U7916 (N_7916,N_6957,N_6189);
or U7917 (N_7917,N_6163,N_6760);
and U7918 (N_7918,N_6668,N_6357);
nand U7919 (N_7919,N_6818,N_6498);
nand U7920 (N_7920,N_6362,N_6851);
nand U7921 (N_7921,N_6376,N_6149);
nand U7922 (N_7922,N_6904,N_6718);
nand U7923 (N_7923,N_6828,N_6692);
and U7924 (N_7924,N_6572,N_6204);
and U7925 (N_7925,N_6435,N_6120);
and U7926 (N_7926,N_6629,N_6640);
nor U7927 (N_7927,N_6718,N_6945);
and U7928 (N_7928,N_6822,N_6104);
and U7929 (N_7929,N_6716,N_6758);
nand U7930 (N_7930,N_6195,N_6358);
nor U7931 (N_7931,N_6349,N_6579);
and U7932 (N_7932,N_6598,N_6266);
or U7933 (N_7933,N_6130,N_6155);
nor U7934 (N_7934,N_6369,N_6206);
or U7935 (N_7935,N_6607,N_6344);
nor U7936 (N_7936,N_6082,N_6383);
nor U7937 (N_7937,N_6281,N_6156);
nor U7938 (N_7938,N_6400,N_6957);
and U7939 (N_7939,N_6054,N_6637);
nor U7940 (N_7940,N_6340,N_6335);
nor U7941 (N_7941,N_6942,N_6067);
or U7942 (N_7942,N_6298,N_6396);
nand U7943 (N_7943,N_6981,N_6045);
and U7944 (N_7944,N_6713,N_6755);
xnor U7945 (N_7945,N_6315,N_6625);
and U7946 (N_7946,N_6875,N_6051);
or U7947 (N_7947,N_6061,N_6185);
or U7948 (N_7948,N_6072,N_6385);
nand U7949 (N_7949,N_6763,N_6263);
and U7950 (N_7950,N_6400,N_6847);
nand U7951 (N_7951,N_6579,N_6623);
nor U7952 (N_7952,N_6550,N_6663);
or U7953 (N_7953,N_6464,N_6853);
nand U7954 (N_7954,N_6856,N_6378);
nand U7955 (N_7955,N_6655,N_6904);
or U7956 (N_7956,N_6533,N_6872);
nor U7957 (N_7957,N_6684,N_6495);
and U7958 (N_7958,N_6904,N_6645);
nand U7959 (N_7959,N_6496,N_6108);
nor U7960 (N_7960,N_6095,N_6153);
nor U7961 (N_7961,N_6072,N_6696);
nand U7962 (N_7962,N_6417,N_6184);
and U7963 (N_7963,N_6636,N_6940);
or U7964 (N_7964,N_6871,N_6025);
or U7965 (N_7965,N_6509,N_6593);
nand U7966 (N_7966,N_6023,N_6818);
nand U7967 (N_7967,N_6397,N_6480);
nor U7968 (N_7968,N_6165,N_6337);
or U7969 (N_7969,N_6780,N_6291);
nand U7970 (N_7970,N_6187,N_6024);
or U7971 (N_7971,N_6128,N_6666);
nand U7972 (N_7972,N_6960,N_6832);
and U7973 (N_7973,N_6271,N_6338);
and U7974 (N_7974,N_6834,N_6543);
or U7975 (N_7975,N_6249,N_6724);
nor U7976 (N_7976,N_6039,N_6638);
and U7977 (N_7977,N_6077,N_6822);
and U7978 (N_7978,N_6381,N_6948);
or U7979 (N_7979,N_6035,N_6354);
or U7980 (N_7980,N_6252,N_6024);
nand U7981 (N_7981,N_6052,N_6051);
nand U7982 (N_7982,N_6094,N_6521);
nor U7983 (N_7983,N_6923,N_6779);
and U7984 (N_7984,N_6835,N_6640);
and U7985 (N_7985,N_6452,N_6400);
nand U7986 (N_7986,N_6262,N_6364);
and U7987 (N_7987,N_6728,N_6025);
and U7988 (N_7988,N_6807,N_6185);
nand U7989 (N_7989,N_6339,N_6755);
or U7990 (N_7990,N_6924,N_6525);
and U7991 (N_7991,N_6541,N_6683);
nand U7992 (N_7992,N_6949,N_6630);
nand U7993 (N_7993,N_6111,N_6310);
nand U7994 (N_7994,N_6760,N_6728);
nand U7995 (N_7995,N_6851,N_6360);
nand U7996 (N_7996,N_6322,N_6857);
nor U7997 (N_7997,N_6112,N_6807);
nand U7998 (N_7998,N_6455,N_6309);
nand U7999 (N_7999,N_6375,N_6112);
or U8000 (N_8000,N_7451,N_7543);
nand U8001 (N_8001,N_7768,N_7994);
nand U8002 (N_8002,N_7252,N_7267);
or U8003 (N_8003,N_7036,N_7747);
or U8004 (N_8004,N_7726,N_7222);
nand U8005 (N_8005,N_7925,N_7044);
or U8006 (N_8006,N_7688,N_7496);
and U8007 (N_8007,N_7875,N_7559);
nand U8008 (N_8008,N_7235,N_7159);
and U8009 (N_8009,N_7492,N_7469);
nor U8010 (N_8010,N_7070,N_7961);
nand U8011 (N_8011,N_7184,N_7326);
nor U8012 (N_8012,N_7314,N_7274);
and U8013 (N_8013,N_7432,N_7756);
nand U8014 (N_8014,N_7748,N_7833);
nor U8015 (N_8015,N_7118,N_7531);
and U8016 (N_8016,N_7308,N_7862);
or U8017 (N_8017,N_7077,N_7124);
xor U8018 (N_8018,N_7318,N_7888);
nor U8019 (N_8019,N_7799,N_7444);
and U8020 (N_8020,N_7401,N_7761);
and U8021 (N_8021,N_7373,N_7105);
nand U8022 (N_8022,N_7494,N_7312);
or U8023 (N_8023,N_7995,N_7063);
and U8024 (N_8024,N_7157,N_7237);
nor U8025 (N_8025,N_7725,N_7233);
nand U8026 (N_8026,N_7632,N_7187);
or U8027 (N_8027,N_7651,N_7043);
nor U8028 (N_8028,N_7923,N_7589);
nand U8029 (N_8029,N_7853,N_7915);
or U8030 (N_8030,N_7269,N_7746);
or U8031 (N_8031,N_7145,N_7803);
nand U8032 (N_8032,N_7609,N_7041);
or U8033 (N_8033,N_7479,N_7968);
xnor U8034 (N_8034,N_7434,N_7565);
or U8035 (N_8035,N_7634,N_7734);
nand U8036 (N_8036,N_7765,N_7652);
and U8037 (N_8037,N_7016,N_7873);
xnor U8038 (N_8038,N_7592,N_7795);
and U8039 (N_8039,N_7655,N_7057);
nor U8040 (N_8040,N_7167,N_7593);
nor U8041 (N_8041,N_7840,N_7532);
and U8042 (N_8042,N_7520,N_7902);
nor U8043 (N_8043,N_7302,N_7100);
and U8044 (N_8044,N_7488,N_7028);
nor U8045 (N_8045,N_7505,N_7218);
and U8046 (N_8046,N_7396,N_7279);
nand U8047 (N_8047,N_7296,N_7564);
and U8048 (N_8048,N_7871,N_7273);
or U8049 (N_8049,N_7539,N_7483);
and U8050 (N_8050,N_7402,N_7838);
or U8051 (N_8051,N_7426,N_7107);
nand U8052 (N_8052,N_7851,N_7395);
nand U8053 (N_8053,N_7360,N_7775);
and U8054 (N_8054,N_7645,N_7439);
and U8055 (N_8055,N_7038,N_7416);
nor U8056 (N_8056,N_7605,N_7018);
nor U8057 (N_8057,N_7368,N_7876);
nor U8058 (N_8058,N_7507,N_7320);
or U8059 (N_8059,N_7717,N_7195);
and U8060 (N_8060,N_7811,N_7497);
or U8061 (N_8061,N_7354,N_7560);
nand U8062 (N_8062,N_7810,N_7990);
nand U8063 (N_8063,N_7653,N_7246);
or U8064 (N_8064,N_7343,N_7394);
nand U8065 (N_8065,N_7677,N_7192);
and U8066 (N_8066,N_7721,N_7827);
nand U8067 (N_8067,N_7856,N_7263);
nor U8068 (N_8068,N_7076,N_7963);
nand U8069 (N_8069,N_7621,N_7914);
or U8070 (N_8070,N_7842,N_7808);
nand U8071 (N_8071,N_7946,N_7309);
nor U8072 (N_8072,N_7051,N_7431);
or U8073 (N_8073,N_7045,N_7813);
or U8074 (N_8074,N_7170,N_7620);
nand U8075 (N_8075,N_7180,N_7919);
nand U8076 (N_8076,N_7174,N_7206);
nor U8077 (N_8077,N_7596,N_7011);
and U8078 (N_8078,N_7452,N_7513);
and U8079 (N_8079,N_7328,N_7903);
nand U8080 (N_8080,N_7511,N_7115);
or U8081 (N_8081,N_7224,N_7441);
and U8082 (N_8082,N_7874,N_7575);
and U8083 (N_8083,N_7739,N_7351);
nand U8084 (N_8084,N_7804,N_7232);
and U8085 (N_8085,N_7460,N_7936);
nor U8086 (N_8086,N_7568,N_7489);
nor U8087 (N_8087,N_7806,N_7937);
nor U8088 (N_8088,N_7147,N_7327);
or U8089 (N_8089,N_7816,N_7899);
nor U8090 (N_8090,N_7023,N_7099);
and U8091 (N_8091,N_7962,N_7997);
nand U8092 (N_8092,N_7472,N_7695);
nor U8093 (N_8093,N_7942,N_7209);
or U8094 (N_8094,N_7030,N_7841);
nand U8095 (N_8095,N_7163,N_7103);
or U8096 (N_8096,N_7084,N_7890);
and U8097 (N_8097,N_7817,N_7372);
nand U8098 (N_8098,N_7859,N_7540);
nand U8099 (N_8099,N_7334,N_7852);
or U8100 (N_8100,N_7188,N_7193);
and U8101 (N_8101,N_7713,N_7732);
nor U8102 (N_8102,N_7608,N_7606);
and U8103 (N_8103,N_7675,N_7125);
or U8104 (N_8104,N_7658,N_7300);
and U8105 (N_8105,N_7176,N_7034);
and U8106 (N_8106,N_7142,N_7219);
nor U8107 (N_8107,N_7735,N_7144);
nand U8108 (N_8108,N_7083,N_7399);
nor U8109 (N_8109,N_7307,N_7945);
nor U8110 (N_8110,N_7301,N_7501);
nand U8111 (N_8111,N_7085,N_7359);
or U8112 (N_8112,N_7283,N_7705);
or U8113 (N_8113,N_7009,N_7330);
nor U8114 (N_8114,N_7635,N_7284);
and U8115 (N_8115,N_7977,N_7064);
and U8116 (N_8116,N_7595,N_7173);
nand U8117 (N_8117,N_7892,N_7484);
nand U8118 (N_8118,N_7062,N_7440);
nand U8119 (N_8119,N_7391,N_7500);
and U8120 (N_8120,N_7162,N_7008);
and U8121 (N_8121,N_7628,N_7864);
or U8122 (N_8122,N_7528,N_7780);
nand U8123 (N_8123,N_7668,N_7268);
nor U8124 (N_8124,N_7525,N_7390);
nor U8125 (N_8125,N_7669,N_7427);
or U8126 (N_8126,N_7435,N_7029);
nand U8127 (N_8127,N_7133,N_7880);
and U8128 (N_8128,N_7638,N_7863);
and U8129 (N_8129,N_7707,N_7088);
or U8130 (N_8130,N_7000,N_7357);
and U8131 (N_8131,N_7371,N_7969);
or U8132 (N_8132,N_7438,N_7317);
nand U8133 (N_8133,N_7367,N_7220);
nand U8134 (N_8134,N_7911,N_7454);
and U8135 (N_8135,N_7680,N_7067);
nand U8136 (N_8136,N_7350,N_7690);
and U8137 (N_8137,N_7517,N_7987);
nor U8138 (N_8138,N_7455,N_7563);
and U8139 (N_8139,N_7214,N_7012);
and U8140 (N_8140,N_7625,N_7829);
or U8141 (N_8141,N_7792,N_7724);
and U8142 (N_8142,N_7666,N_7745);
nand U8143 (N_8143,N_7908,N_7490);
or U8144 (N_8144,N_7555,N_7927);
or U8145 (N_8145,N_7644,N_7823);
nand U8146 (N_8146,N_7904,N_7411);
or U8147 (N_8147,N_7633,N_7509);
nor U8148 (N_8148,N_7336,N_7763);
nand U8149 (N_8149,N_7897,N_7388);
and U8150 (N_8150,N_7230,N_7313);
nand U8151 (N_8151,N_7935,N_7749);
nand U8152 (N_8152,N_7831,N_7339);
and U8153 (N_8153,N_7461,N_7319);
nor U8154 (N_8154,N_7259,N_7442);
nor U8155 (N_8155,N_7380,N_7957);
and U8156 (N_8156,N_7169,N_7534);
and U8157 (N_8157,N_7253,N_7884);
or U8158 (N_8158,N_7861,N_7190);
and U8159 (N_8159,N_7211,N_7533);
nand U8160 (N_8160,N_7117,N_7930);
nand U8161 (N_8161,N_7938,N_7689);
nor U8162 (N_8162,N_7098,N_7171);
and U8163 (N_8163,N_7907,N_7346);
and U8164 (N_8164,N_7843,N_7983);
nand U8165 (N_8165,N_7421,N_7129);
or U8166 (N_8166,N_7132,N_7151);
and U8167 (N_8167,N_7600,N_7499);
and U8168 (N_8168,N_7583,N_7581);
or U8169 (N_8169,N_7264,N_7882);
and U8170 (N_8170,N_7976,N_7754);
nor U8171 (N_8171,N_7248,N_7039);
nand U8172 (N_8172,N_7877,N_7290);
nor U8173 (N_8173,N_7094,N_7771);
nand U8174 (N_8174,N_7671,N_7556);
or U8175 (N_8175,N_7139,N_7537);
or U8176 (N_8176,N_7090,N_7844);
nand U8177 (N_8177,N_7141,N_7185);
or U8178 (N_8178,N_7545,N_7299);
and U8179 (N_8179,N_7657,N_7755);
nor U8180 (N_8180,N_7213,N_7549);
nor U8181 (N_8181,N_7152,N_7052);
nand U8182 (N_8182,N_7566,N_7287);
or U8183 (N_8183,N_7934,N_7909);
nor U8184 (N_8184,N_7358,N_7203);
nor U8185 (N_8185,N_7325,N_7515);
nand U8186 (N_8186,N_7017,N_7991);
xnor U8187 (N_8187,N_7573,N_7065);
or U8188 (N_8188,N_7698,N_7392);
nand U8189 (N_8189,N_7424,N_7074);
nor U8190 (N_8190,N_7766,N_7538);
or U8191 (N_8191,N_7182,N_7998);
or U8192 (N_8192,N_7800,N_7604);
nand U8193 (N_8193,N_7413,N_7049);
nand U8194 (N_8194,N_7199,N_7767);
nor U8195 (N_8195,N_7356,N_7123);
nor U8196 (N_8196,N_7362,N_7068);
nand U8197 (N_8197,N_7420,N_7447);
or U8198 (N_8198,N_7542,N_7202);
and U8199 (N_8199,N_7751,N_7239);
nand U8200 (N_8200,N_7710,N_7985);
and U8201 (N_8201,N_7241,N_7275);
or U8202 (N_8202,N_7640,N_7126);
or U8203 (N_8203,N_7429,N_7082);
nor U8204 (N_8204,N_7629,N_7311);
or U8205 (N_8205,N_7055,N_7040);
and U8206 (N_8206,N_7281,N_7437);
nand U8207 (N_8207,N_7458,N_7574);
and U8208 (N_8208,N_7626,N_7929);
or U8209 (N_8209,N_7958,N_7854);
or U8210 (N_8210,N_7262,N_7329);
and U8211 (N_8211,N_7385,N_7616);
and U8212 (N_8212,N_7647,N_7485);
or U8213 (N_8213,N_7217,N_7673);
or U8214 (N_8214,N_7338,N_7196);
or U8215 (N_8215,N_7005,N_7097);
nand U8216 (N_8216,N_7430,N_7002);
or U8217 (N_8217,N_7631,N_7924);
nand U8218 (N_8218,N_7364,N_7014);
or U8219 (N_8219,N_7798,N_7603);
and U8220 (N_8220,N_7153,N_7069);
nand U8221 (N_8221,N_7205,N_7297);
and U8222 (N_8222,N_7042,N_7857);
nand U8223 (N_8223,N_7703,N_7114);
nand U8224 (N_8224,N_7266,N_7656);
and U8225 (N_8225,N_7720,N_7168);
and U8226 (N_8226,N_7591,N_7850);
and U8227 (N_8227,N_7419,N_7530);
nor U8228 (N_8228,N_7086,N_7932);
and U8229 (N_8229,N_7236,N_7245);
xor U8230 (N_8230,N_7331,N_7178);
nand U8231 (N_8231,N_7701,N_7601);
and U8232 (N_8232,N_7448,N_7744);
or U8233 (N_8233,N_7835,N_7477);
nand U8234 (N_8234,N_7481,N_7926);
nor U8235 (N_8235,N_7414,N_7917);
nand U8236 (N_8236,N_7304,N_7164);
or U8237 (N_8237,N_7053,N_7201);
or U8238 (N_8238,N_7900,N_7712);
and U8239 (N_8239,N_7750,N_7022);
or U8240 (N_8240,N_7112,N_7387);
or U8241 (N_8241,N_7369,N_7104);
nand U8242 (N_8242,N_7736,N_7887);
nor U8243 (N_8243,N_7582,N_7271);
or U8244 (N_8244,N_7407,N_7409);
nand U8245 (N_8245,N_7298,N_7665);
nand U8246 (N_8246,N_7825,N_7753);
nor U8247 (N_8247,N_7109,N_7594);
and U8248 (N_8248,N_7672,N_7954);
or U8249 (N_8249,N_7664,N_7860);
nand U8250 (N_8250,N_7940,N_7355);
nor U8251 (N_8251,N_7805,N_7138);
nor U8252 (N_8252,N_7198,N_7557);
nor U8253 (N_8253,N_7423,N_7941);
nor U8254 (N_8254,N_7686,N_7809);
and U8255 (N_8255,N_7648,N_7839);
nand U8256 (N_8256,N_7928,N_7374);
nand U8257 (N_8257,N_7378,N_7127);
or U8258 (N_8258,N_7377,N_7881);
nand U8259 (N_8259,N_7459,N_7986);
nor U8260 (N_8260,N_7847,N_7554);
nand U8261 (N_8261,N_7569,N_7580);
nand U8262 (N_8262,N_7349,N_7365);
nor U8263 (N_8263,N_7474,N_7704);
and U8264 (N_8264,N_7054,N_7512);
nor U8265 (N_8265,N_7812,N_7933);
nand U8266 (N_8266,N_7315,N_7687);
nand U8267 (N_8267,N_7150,N_7410);
or U8268 (N_8268,N_7973,N_7918);
nor U8269 (N_8269,N_7955,N_7495);
or U8270 (N_8270,N_7676,N_7031);
and U8271 (N_8271,N_7122,N_7649);
nor U8272 (N_8272,N_7674,N_7836);
or U8273 (N_8273,N_7119,N_7135);
and U8274 (N_8274,N_7212,N_7110);
and U8275 (N_8275,N_7571,N_7376);
and U8276 (N_8276,N_7337,N_7944);
or U8277 (N_8277,N_7551,N_7116);
nor U8278 (N_8278,N_7272,N_7280);
or U8279 (N_8279,N_7491,N_7790);
and U8280 (N_8280,N_7971,N_7793);
or U8281 (N_8281,N_7503,N_7161);
nand U8282 (N_8282,N_7026,N_7613);
or U8283 (N_8283,N_7037,N_7425);
or U8284 (N_8284,N_7916,N_7353);
nand U8285 (N_8285,N_7363,N_7967);
nor U8286 (N_8286,N_7743,N_7659);
or U8287 (N_8287,N_7684,N_7417);
nor U8288 (N_8288,N_7140,N_7047);
nor U8289 (N_8289,N_7694,N_7508);
and U8290 (N_8290,N_7291,N_7092);
nor U8291 (N_8291,N_7727,N_7693);
or U8292 (N_8292,N_7375,N_7821);
nand U8293 (N_8293,N_7579,N_7885);
nor U8294 (N_8294,N_7342,N_7519);
nand U8295 (N_8295,N_7059,N_7783);
or U8296 (N_8296,N_7641,N_7293);
nand U8297 (N_8297,N_7160,N_7443);
nand U8298 (N_8298,N_7324,N_7692);
nor U8299 (N_8299,N_7234,N_7516);
nand U8300 (N_8300,N_7678,N_7277);
or U8301 (N_8301,N_7699,N_7465);
or U8302 (N_8302,N_7247,N_7415);
and U8303 (N_8303,N_7316,N_7970);
nand U8304 (N_8304,N_7462,N_7518);
and U8305 (N_8305,N_7265,N_7013);
nor U8306 (N_8306,N_7521,N_7920);
nor U8307 (N_8307,N_7587,N_7471);
nor U8308 (N_8308,N_7614,N_7258);
nor U8309 (N_8309,N_7345,N_7397);
nand U8310 (N_8310,N_7959,N_7889);
or U8311 (N_8311,N_7956,N_7691);
xnor U8312 (N_8312,N_7215,N_7244);
nand U8313 (N_8313,N_7352,N_7001);
or U8314 (N_8314,N_7183,N_7384);
and U8315 (N_8315,N_7654,N_7586);
and U8316 (N_8316,N_7493,N_7642);
xor U8317 (N_8317,N_7544,N_7514);
nor U8318 (N_8318,N_7627,N_7607);
and U8319 (N_8319,N_7344,N_7989);
or U8320 (N_8320,N_7035,N_7663);
and U8321 (N_8321,N_7643,N_7361);
nand U8322 (N_8322,N_7577,N_7737);
nand U8323 (N_8323,N_7130,N_7951);
and U8324 (N_8324,N_7243,N_7254);
nand U8325 (N_8325,N_7033,N_7504);
and U8326 (N_8326,N_7788,N_7108);
or U8327 (N_8327,N_7091,N_7120);
nand U8328 (N_8328,N_7348,N_7733);
or U8329 (N_8329,N_7468,N_7335);
and U8330 (N_8330,N_7981,N_7572);
nor U8331 (N_8331,N_7470,N_7498);
nor U8332 (N_8332,N_7660,N_7696);
nand U8333 (N_8333,N_7146,N_7422);
nand U8334 (N_8334,N_7553,N_7370);
or U8335 (N_8335,N_7019,N_7791);
and U8336 (N_8336,N_7081,N_7463);
nor U8337 (N_8337,N_7984,N_7590);
or U8338 (N_8338,N_7585,N_7868);
or U8339 (N_8339,N_7408,N_7858);
and U8340 (N_8340,N_7867,N_7506);
or U8341 (N_8341,N_7166,N_7257);
nand U8342 (N_8342,N_7238,N_7295);
nand U8343 (N_8343,N_7848,N_7670);
or U8344 (N_8344,N_7714,N_7950);
or U8345 (N_8345,N_7898,N_7136);
nor U8346 (N_8346,N_7913,N_7403);
or U8347 (N_8347,N_7878,N_7612);
and U8348 (N_8348,N_7306,N_7131);
and U8349 (N_8349,N_7972,N_7548);
nor U8350 (N_8350,N_7286,N_7906);
nor U8351 (N_8351,N_7723,N_7834);
nor U8352 (N_8352,N_7637,N_7711);
or U8353 (N_8353,N_7901,N_7822);
and U8354 (N_8354,N_7718,N_7191);
or U8355 (N_8355,N_7197,N_7740);
or U8356 (N_8356,N_7412,N_7393);
or U8357 (N_8357,N_7781,N_7060);
nor U8358 (N_8358,N_7730,N_7667);
nand U8359 (N_8359,N_7570,N_7960);
and U8360 (N_8360,N_7027,N_7773);
nor U8361 (N_8361,N_7722,N_7288);
and U8362 (N_8362,N_7156,N_7895);
and U8363 (N_8363,N_7630,N_7386);
nor U8364 (N_8364,N_7204,N_7610);
or U8365 (N_8365,N_7870,N_7467);
nand U8366 (N_8366,N_7774,N_7294);
or U8367 (N_8367,N_7547,N_7075);
nand U8368 (N_8368,N_7679,N_7762);
and U8369 (N_8369,N_7786,N_7700);
nand U8370 (N_8370,N_7260,N_7025);
nand U8371 (N_8371,N_7993,N_7032);
or U8372 (N_8372,N_7400,N_7826);
and U8373 (N_8373,N_7524,N_7794);
nand U8374 (N_8374,N_7636,N_7787);
or U8375 (N_8375,N_7742,N_7289);
nand U8376 (N_8376,N_7475,N_7321);
or U8377 (N_8377,N_7210,N_7466);
nand U8378 (N_8378,N_7964,N_7073);
nand U8379 (N_8379,N_7883,N_7510);
or U8380 (N_8380,N_7615,N_7476);
nand U8381 (N_8381,N_7584,N_7179);
or U8382 (N_8382,N_7079,N_7276);
or U8383 (N_8383,N_7784,N_7979);
and U8384 (N_8384,N_7134,N_7341);
and U8385 (N_8385,N_7797,N_7550);
nand U8386 (N_8386,N_7228,N_7974);
and U8387 (N_8387,N_7869,N_7398);
nand U8388 (N_8388,N_7980,N_7121);
and U8389 (N_8389,N_7250,N_7200);
or U8390 (N_8390,N_7617,N_7802);
and U8391 (N_8391,N_7406,N_7966);
nand U8392 (N_8392,N_7820,N_7685);
and U8393 (N_8393,N_7061,N_7830);
or U8394 (N_8394,N_7865,N_7709);
nand U8395 (N_8395,N_7240,N_7261);
or U8396 (N_8396,N_7716,N_7155);
nand U8397 (N_8397,N_7292,N_7529);
or U8398 (N_8398,N_7681,N_7778);
nand U8399 (N_8399,N_7522,N_7251);
nand U8400 (N_8400,N_7552,N_7752);
nand U8401 (N_8401,N_7148,N_7482);
and U8402 (N_8402,N_7741,N_7846);
nor U8403 (N_8403,N_7772,N_7332);
and U8404 (N_8404,N_7223,N_7015);
nor U8405 (N_8405,N_7457,N_7845);
nor U8406 (N_8406,N_7093,N_7789);
nand U8407 (N_8407,N_7769,N_7922);
nand U8408 (N_8408,N_7891,N_7020);
nor U8409 (N_8409,N_7619,N_7270);
nand U8410 (N_8410,N_7988,N_7177);
and U8411 (N_8411,N_7562,N_7004);
nor U8412 (N_8412,N_7588,N_7894);
or U8413 (N_8413,N_7256,N_7999);
nand U8414 (N_8414,N_7096,N_7450);
or U8415 (N_8415,N_7087,N_7101);
and U8416 (N_8416,N_7828,N_7527);
or U8417 (N_8417,N_7389,N_7347);
and U8418 (N_8418,N_7611,N_7216);
or U8419 (N_8419,N_7661,N_7526);
nor U8420 (N_8420,N_7815,N_7080);
and U8421 (N_8421,N_7445,N_7078);
nor U8422 (N_8422,N_7728,N_7056);
nor U8423 (N_8423,N_7006,N_7186);
or U8424 (N_8424,N_7910,N_7282);
and U8425 (N_8425,N_7622,N_7486);
nor U8426 (N_8426,N_7058,N_7137);
or U8427 (N_8427,N_7650,N_7111);
nor U8428 (N_8428,N_7285,N_7921);
nand U8429 (N_8429,N_7456,N_7824);
nor U8430 (N_8430,N_7576,N_7436);
nand U8431 (N_8431,N_7879,N_7208);
nand U8432 (N_8432,N_7305,N_7702);
xor U8433 (N_8433,N_7165,N_7708);
and U8434 (N_8434,N_7639,N_7221);
nor U8435 (N_8435,N_7487,N_7623);
and U8436 (N_8436,N_7102,N_7523);
or U8437 (N_8437,N_7715,N_7567);
nand U8438 (N_8438,N_7478,N_7949);
and U8439 (N_8439,N_7738,N_7757);
or U8440 (N_8440,N_7535,N_7226);
nand U8441 (N_8441,N_7558,N_7646);
nor U8442 (N_8442,N_7449,N_7382);
xor U8443 (N_8443,N_7383,N_7189);
nand U8444 (N_8444,N_7578,N_7278);
or U8445 (N_8445,N_7379,N_7323);
nor U8446 (N_8446,N_7818,N_7807);
nand U8447 (N_8447,N_7003,N_7758);
and U8448 (N_8448,N_7837,N_7066);
and U8449 (N_8449,N_7149,N_7975);
nor U8450 (N_8450,N_7965,N_7175);
and U8451 (N_8451,N_7996,N_7089);
nor U8452 (N_8452,N_7255,N_7948);
or U8453 (N_8453,N_7207,N_7598);
nor U8454 (N_8454,N_7418,N_7095);
nor U8455 (N_8455,N_7814,N_7154);
nor U8456 (N_8456,N_7952,N_7599);
or U8457 (N_8457,N_7697,N_7682);
nor U8458 (N_8458,N_7464,N_7249);
or U8459 (N_8459,N_7007,N_7428);
nor U8460 (N_8460,N_7128,N_7801);
nor U8461 (N_8461,N_7143,N_7333);
and U8462 (N_8462,N_7106,N_7404);
nor U8463 (N_8463,N_7453,N_7480);
nor U8464 (N_8464,N_7158,N_7731);
nor U8465 (N_8465,N_7381,N_7340);
and U8466 (N_8466,N_7227,N_7194);
nor U8467 (N_8467,N_7785,N_7849);
nor U8468 (N_8468,N_7433,N_7764);
nand U8469 (N_8469,N_7473,N_7992);
and U8470 (N_8470,N_7546,N_7010);
nor U8471 (N_8471,N_7618,N_7048);
nand U8472 (N_8472,N_7310,N_7366);
or U8473 (N_8473,N_7978,N_7050);
or U8474 (N_8474,N_7624,N_7303);
or U8475 (N_8475,N_7072,N_7782);
and U8476 (N_8476,N_7683,N_7760);
and U8477 (N_8477,N_7242,N_7597);
nor U8478 (N_8478,N_7893,N_7536);
nor U8479 (N_8479,N_7021,N_7172);
nand U8480 (N_8480,N_7322,N_7502);
nand U8481 (N_8481,N_7819,N_7759);
nand U8482 (N_8482,N_7719,N_7446);
nor U8483 (N_8483,N_7231,N_7113);
nand U8484 (N_8484,N_7181,N_7939);
nand U8485 (N_8485,N_7024,N_7943);
nor U8486 (N_8486,N_7931,N_7729);
and U8487 (N_8487,N_7896,N_7561);
nand U8488 (N_8488,N_7886,N_7982);
and U8489 (N_8489,N_7953,N_7832);
xor U8490 (N_8490,N_7541,N_7662);
nand U8491 (N_8491,N_7872,N_7706);
or U8492 (N_8492,N_7776,N_7770);
nor U8493 (N_8493,N_7405,N_7779);
and U8494 (N_8494,N_7796,N_7046);
and U8495 (N_8495,N_7229,N_7905);
nand U8496 (N_8496,N_7071,N_7225);
and U8497 (N_8497,N_7912,N_7855);
or U8498 (N_8498,N_7602,N_7777);
nand U8499 (N_8499,N_7947,N_7866);
or U8500 (N_8500,N_7514,N_7749);
nand U8501 (N_8501,N_7407,N_7275);
nand U8502 (N_8502,N_7532,N_7342);
nor U8503 (N_8503,N_7560,N_7150);
and U8504 (N_8504,N_7295,N_7149);
nor U8505 (N_8505,N_7103,N_7808);
or U8506 (N_8506,N_7456,N_7586);
nand U8507 (N_8507,N_7877,N_7829);
or U8508 (N_8508,N_7431,N_7723);
or U8509 (N_8509,N_7912,N_7806);
nand U8510 (N_8510,N_7930,N_7936);
nand U8511 (N_8511,N_7420,N_7001);
or U8512 (N_8512,N_7990,N_7717);
or U8513 (N_8513,N_7141,N_7840);
and U8514 (N_8514,N_7430,N_7219);
nand U8515 (N_8515,N_7769,N_7503);
or U8516 (N_8516,N_7172,N_7327);
nand U8517 (N_8517,N_7618,N_7339);
nand U8518 (N_8518,N_7243,N_7400);
and U8519 (N_8519,N_7272,N_7246);
nand U8520 (N_8520,N_7452,N_7986);
nor U8521 (N_8521,N_7907,N_7427);
nor U8522 (N_8522,N_7875,N_7050);
and U8523 (N_8523,N_7295,N_7007);
or U8524 (N_8524,N_7103,N_7123);
nand U8525 (N_8525,N_7992,N_7640);
nor U8526 (N_8526,N_7019,N_7066);
and U8527 (N_8527,N_7769,N_7063);
or U8528 (N_8528,N_7033,N_7236);
nand U8529 (N_8529,N_7286,N_7615);
or U8530 (N_8530,N_7706,N_7993);
and U8531 (N_8531,N_7970,N_7709);
and U8532 (N_8532,N_7118,N_7265);
or U8533 (N_8533,N_7375,N_7923);
and U8534 (N_8534,N_7070,N_7111);
and U8535 (N_8535,N_7169,N_7033);
nand U8536 (N_8536,N_7168,N_7150);
or U8537 (N_8537,N_7655,N_7436);
and U8538 (N_8538,N_7254,N_7771);
nand U8539 (N_8539,N_7325,N_7916);
or U8540 (N_8540,N_7646,N_7437);
nor U8541 (N_8541,N_7827,N_7032);
nor U8542 (N_8542,N_7559,N_7058);
nand U8543 (N_8543,N_7435,N_7737);
or U8544 (N_8544,N_7452,N_7500);
nand U8545 (N_8545,N_7917,N_7837);
and U8546 (N_8546,N_7210,N_7495);
nand U8547 (N_8547,N_7774,N_7498);
and U8548 (N_8548,N_7597,N_7349);
nand U8549 (N_8549,N_7205,N_7304);
or U8550 (N_8550,N_7966,N_7265);
or U8551 (N_8551,N_7019,N_7241);
nand U8552 (N_8552,N_7691,N_7900);
nand U8553 (N_8553,N_7426,N_7968);
nand U8554 (N_8554,N_7964,N_7378);
and U8555 (N_8555,N_7258,N_7846);
or U8556 (N_8556,N_7087,N_7192);
or U8557 (N_8557,N_7614,N_7909);
nand U8558 (N_8558,N_7345,N_7739);
or U8559 (N_8559,N_7441,N_7444);
nand U8560 (N_8560,N_7663,N_7468);
nand U8561 (N_8561,N_7686,N_7884);
nand U8562 (N_8562,N_7376,N_7695);
or U8563 (N_8563,N_7893,N_7867);
or U8564 (N_8564,N_7437,N_7147);
nor U8565 (N_8565,N_7906,N_7165);
and U8566 (N_8566,N_7692,N_7135);
or U8567 (N_8567,N_7500,N_7914);
or U8568 (N_8568,N_7819,N_7250);
nor U8569 (N_8569,N_7475,N_7319);
and U8570 (N_8570,N_7249,N_7086);
or U8571 (N_8571,N_7273,N_7964);
nor U8572 (N_8572,N_7407,N_7552);
nor U8573 (N_8573,N_7690,N_7449);
or U8574 (N_8574,N_7773,N_7940);
or U8575 (N_8575,N_7995,N_7765);
nand U8576 (N_8576,N_7888,N_7997);
nand U8577 (N_8577,N_7839,N_7271);
nand U8578 (N_8578,N_7212,N_7927);
or U8579 (N_8579,N_7042,N_7050);
or U8580 (N_8580,N_7535,N_7189);
or U8581 (N_8581,N_7412,N_7751);
or U8582 (N_8582,N_7763,N_7250);
nand U8583 (N_8583,N_7674,N_7935);
or U8584 (N_8584,N_7315,N_7560);
or U8585 (N_8585,N_7460,N_7779);
or U8586 (N_8586,N_7938,N_7752);
or U8587 (N_8587,N_7969,N_7488);
or U8588 (N_8588,N_7737,N_7155);
nor U8589 (N_8589,N_7775,N_7002);
nand U8590 (N_8590,N_7691,N_7060);
and U8591 (N_8591,N_7873,N_7375);
and U8592 (N_8592,N_7376,N_7223);
nor U8593 (N_8593,N_7419,N_7668);
nor U8594 (N_8594,N_7718,N_7791);
nand U8595 (N_8595,N_7069,N_7175);
or U8596 (N_8596,N_7520,N_7437);
nand U8597 (N_8597,N_7244,N_7780);
and U8598 (N_8598,N_7806,N_7002);
or U8599 (N_8599,N_7500,N_7071);
and U8600 (N_8600,N_7931,N_7885);
nand U8601 (N_8601,N_7109,N_7057);
nand U8602 (N_8602,N_7515,N_7574);
or U8603 (N_8603,N_7932,N_7930);
or U8604 (N_8604,N_7802,N_7674);
or U8605 (N_8605,N_7614,N_7598);
and U8606 (N_8606,N_7963,N_7526);
or U8607 (N_8607,N_7959,N_7542);
and U8608 (N_8608,N_7905,N_7530);
or U8609 (N_8609,N_7706,N_7168);
nand U8610 (N_8610,N_7709,N_7449);
and U8611 (N_8611,N_7200,N_7513);
nor U8612 (N_8612,N_7841,N_7408);
nand U8613 (N_8613,N_7401,N_7185);
nand U8614 (N_8614,N_7694,N_7642);
and U8615 (N_8615,N_7132,N_7007);
nand U8616 (N_8616,N_7581,N_7903);
and U8617 (N_8617,N_7564,N_7804);
or U8618 (N_8618,N_7076,N_7326);
or U8619 (N_8619,N_7373,N_7473);
nand U8620 (N_8620,N_7571,N_7930);
and U8621 (N_8621,N_7517,N_7457);
nor U8622 (N_8622,N_7460,N_7588);
and U8623 (N_8623,N_7777,N_7872);
nor U8624 (N_8624,N_7486,N_7589);
and U8625 (N_8625,N_7087,N_7425);
and U8626 (N_8626,N_7767,N_7865);
nor U8627 (N_8627,N_7719,N_7265);
or U8628 (N_8628,N_7626,N_7608);
xnor U8629 (N_8629,N_7361,N_7167);
xnor U8630 (N_8630,N_7964,N_7131);
or U8631 (N_8631,N_7601,N_7923);
nor U8632 (N_8632,N_7602,N_7501);
nand U8633 (N_8633,N_7394,N_7823);
and U8634 (N_8634,N_7751,N_7543);
nand U8635 (N_8635,N_7466,N_7254);
nand U8636 (N_8636,N_7454,N_7801);
nand U8637 (N_8637,N_7882,N_7141);
nand U8638 (N_8638,N_7310,N_7100);
or U8639 (N_8639,N_7165,N_7497);
nor U8640 (N_8640,N_7446,N_7503);
nor U8641 (N_8641,N_7713,N_7240);
nand U8642 (N_8642,N_7638,N_7352);
nand U8643 (N_8643,N_7023,N_7699);
and U8644 (N_8644,N_7008,N_7694);
nor U8645 (N_8645,N_7824,N_7390);
or U8646 (N_8646,N_7615,N_7007);
nand U8647 (N_8647,N_7641,N_7569);
or U8648 (N_8648,N_7078,N_7171);
nor U8649 (N_8649,N_7342,N_7745);
nand U8650 (N_8650,N_7717,N_7242);
nand U8651 (N_8651,N_7604,N_7293);
or U8652 (N_8652,N_7249,N_7053);
and U8653 (N_8653,N_7727,N_7234);
nand U8654 (N_8654,N_7498,N_7023);
and U8655 (N_8655,N_7281,N_7653);
nor U8656 (N_8656,N_7344,N_7774);
or U8657 (N_8657,N_7527,N_7285);
nand U8658 (N_8658,N_7634,N_7810);
or U8659 (N_8659,N_7925,N_7945);
nand U8660 (N_8660,N_7800,N_7934);
and U8661 (N_8661,N_7083,N_7504);
xor U8662 (N_8662,N_7510,N_7006);
nor U8663 (N_8663,N_7057,N_7529);
nor U8664 (N_8664,N_7189,N_7624);
and U8665 (N_8665,N_7353,N_7377);
and U8666 (N_8666,N_7328,N_7224);
or U8667 (N_8667,N_7816,N_7642);
and U8668 (N_8668,N_7275,N_7550);
nand U8669 (N_8669,N_7135,N_7474);
and U8670 (N_8670,N_7585,N_7797);
and U8671 (N_8671,N_7965,N_7777);
or U8672 (N_8672,N_7528,N_7159);
and U8673 (N_8673,N_7491,N_7968);
or U8674 (N_8674,N_7356,N_7869);
nand U8675 (N_8675,N_7946,N_7663);
and U8676 (N_8676,N_7932,N_7366);
or U8677 (N_8677,N_7060,N_7895);
nand U8678 (N_8678,N_7173,N_7249);
xnor U8679 (N_8679,N_7554,N_7161);
and U8680 (N_8680,N_7005,N_7380);
nor U8681 (N_8681,N_7748,N_7736);
or U8682 (N_8682,N_7719,N_7095);
or U8683 (N_8683,N_7858,N_7955);
or U8684 (N_8684,N_7874,N_7536);
or U8685 (N_8685,N_7615,N_7226);
nor U8686 (N_8686,N_7953,N_7236);
or U8687 (N_8687,N_7141,N_7582);
nor U8688 (N_8688,N_7944,N_7217);
and U8689 (N_8689,N_7430,N_7126);
xnor U8690 (N_8690,N_7783,N_7798);
or U8691 (N_8691,N_7259,N_7242);
nand U8692 (N_8692,N_7621,N_7629);
nand U8693 (N_8693,N_7086,N_7377);
nor U8694 (N_8694,N_7873,N_7520);
and U8695 (N_8695,N_7570,N_7912);
or U8696 (N_8696,N_7163,N_7434);
and U8697 (N_8697,N_7071,N_7777);
nor U8698 (N_8698,N_7443,N_7004);
nand U8699 (N_8699,N_7474,N_7306);
nor U8700 (N_8700,N_7940,N_7738);
or U8701 (N_8701,N_7489,N_7552);
nand U8702 (N_8702,N_7225,N_7771);
nor U8703 (N_8703,N_7140,N_7210);
nor U8704 (N_8704,N_7647,N_7944);
or U8705 (N_8705,N_7836,N_7379);
and U8706 (N_8706,N_7674,N_7180);
xnor U8707 (N_8707,N_7114,N_7956);
and U8708 (N_8708,N_7196,N_7687);
nand U8709 (N_8709,N_7927,N_7989);
and U8710 (N_8710,N_7132,N_7145);
nand U8711 (N_8711,N_7071,N_7081);
and U8712 (N_8712,N_7472,N_7557);
and U8713 (N_8713,N_7407,N_7659);
nand U8714 (N_8714,N_7916,N_7718);
or U8715 (N_8715,N_7312,N_7368);
nor U8716 (N_8716,N_7826,N_7586);
nand U8717 (N_8717,N_7120,N_7972);
or U8718 (N_8718,N_7877,N_7985);
nand U8719 (N_8719,N_7831,N_7574);
or U8720 (N_8720,N_7777,N_7278);
nor U8721 (N_8721,N_7894,N_7213);
nand U8722 (N_8722,N_7115,N_7692);
xor U8723 (N_8723,N_7279,N_7588);
nand U8724 (N_8724,N_7620,N_7403);
and U8725 (N_8725,N_7526,N_7940);
and U8726 (N_8726,N_7523,N_7371);
and U8727 (N_8727,N_7902,N_7657);
and U8728 (N_8728,N_7927,N_7887);
nor U8729 (N_8729,N_7759,N_7826);
and U8730 (N_8730,N_7923,N_7667);
nand U8731 (N_8731,N_7206,N_7489);
or U8732 (N_8732,N_7588,N_7979);
and U8733 (N_8733,N_7103,N_7027);
or U8734 (N_8734,N_7551,N_7185);
nor U8735 (N_8735,N_7508,N_7313);
or U8736 (N_8736,N_7596,N_7602);
nand U8737 (N_8737,N_7333,N_7117);
and U8738 (N_8738,N_7066,N_7229);
nor U8739 (N_8739,N_7545,N_7867);
nor U8740 (N_8740,N_7001,N_7055);
nand U8741 (N_8741,N_7759,N_7004);
nor U8742 (N_8742,N_7692,N_7037);
nor U8743 (N_8743,N_7888,N_7152);
or U8744 (N_8744,N_7302,N_7355);
or U8745 (N_8745,N_7197,N_7671);
or U8746 (N_8746,N_7675,N_7426);
nand U8747 (N_8747,N_7642,N_7866);
nand U8748 (N_8748,N_7001,N_7675);
nand U8749 (N_8749,N_7455,N_7130);
or U8750 (N_8750,N_7380,N_7955);
or U8751 (N_8751,N_7661,N_7625);
nand U8752 (N_8752,N_7136,N_7572);
and U8753 (N_8753,N_7430,N_7859);
or U8754 (N_8754,N_7267,N_7231);
and U8755 (N_8755,N_7881,N_7332);
or U8756 (N_8756,N_7137,N_7321);
nor U8757 (N_8757,N_7518,N_7318);
nand U8758 (N_8758,N_7570,N_7231);
or U8759 (N_8759,N_7781,N_7408);
or U8760 (N_8760,N_7564,N_7158);
nor U8761 (N_8761,N_7875,N_7251);
or U8762 (N_8762,N_7413,N_7575);
nor U8763 (N_8763,N_7549,N_7540);
and U8764 (N_8764,N_7476,N_7063);
and U8765 (N_8765,N_7634,N_7579);
and U8766 (N_8766,N_7864,N_7588);
and U8767 (N_8767,N_7739,N_7259);
and U8768 (N_8768,N_7624,N_7920);
nor U8769 (N_8769,N_7507,N_7872);
and U8770 (N_8770,N_7731,N_7406);
nand U8771 (N_8771,N_7172,N_7200);
nor U8772 (N_8772,N_7628,N_7322);
nor U8773 (N_8773,N_7141,N_7135);
nor U8774 (N_8774,N_7079,N_7122);
and U8775 (N_8775,N_7346,N_7464);
nand U8776 (N_8776,N_7728,N_7973);
and U8777 (N_8777,N_7055,N_7131);
nand U8778 (N_8778,N_7080,N_7622);
nand U8779 (N_8779,N_7605,N_7561);
or U8780 (N_8780,N_7504,N_7638);
nor U8781 (N_8781,N_7585,N_7578);
and U8782 (N_8782,N_7815,N_7863);
xnor U8783 (N_8783,N_7517,N_7065);
nand U8784 (N_8784,N_7848,N_7010);
nor U8785 (N_8785,N_7262,N_7087);
or U8786 (N_8786,N_7757,N_7321);
and U8787 (N_8787,N_7183,N_7989);
and U8788 (N_8788,N_7640,N_7281);
nand U8789 (N_8789,N_7521,N_7240);
or U8790 (N_8790,N_7147,N_7238);
nand U8791 (N_8791,N_7014,N_7749);
nand U8792 (N_8792,N_7023,N_7861);
nor U8793 (N_8793,N_7450,N_7318);
nand U8794 (N_8794,N_7579,N_7529);
nor U8795 (N_8795,N_7406,N_7889);
or U8796 (N_8796,N_7138,N_7459);
nor U8797 (N_8797,N_7338,N_7322);
nor U8798 (N_8798,N_7486,N_7113);
nand U8799 (N_8799,N_7868,N_7309);
nor U8800 (N_8800,N_7164,N_7614);
or U8801 (N_8801,N_7351,N_7149);
and U8802 (N_8802,N_7832,N_7206);
nor U8803 (N_8803,N_7070,N_7896);
or U8804 (N_8804,N_7342,N_7833);
and U8805 (N_8805,N_7345,N_7457);
nand U8806 (N_8806,N_7357,N_7752);
nand U8807 (N_8807,N_7877,N_7025);
or U8808 (N_8808,N_7486,N_7071);
nor U8809 (N_8809,N_7521,N_7585);
nand U8810 (N_8810,N_7157,N_7473);
nor U8811 (N_8811,N_7074,N_7950);
nor U8812 (N_8812,N_7755,N_7142);
nor U8813 (N_8813,N_7661,N_7796);
or U8814 (N_8814,N_7124,N_7941);
nand U8815 (N_8815,N_7515,N_7848);
and U8816 (N_8816,N_7185,N_7188);
and U8817 (N_8817,N_7474,N_7600);
nor U8818 (N_8818,N_7714,N_7047);
nor U8819 (N_8819,N_7641,N_7148);
nand U8820 (N_8820,N_7258,N_7053);
nor U8821 (N_8821,N_7148,N_7653);
and U8822 (N_8822,N_7862,N_7515);
xor U8823 (N_8823,N_7970,N_7705);
or U8824 (N_8824,N_7690,N_7643);
and U8825 (N_8825,N_7699,N_7697);
or U8826 (N_8826,N_7201,N_7898);
nor U8827 (N_8827,N_7995,N_7894);
and U8828 (N_8828,N_7194,N_7639);
nor U8829 (N_8829,N_7094,N_7890);
nor U8830 (N_8830,N_7618,N_7405);
nand U8831 (N_8831,N_7772,N_7583);
or U8832 (N_8832,N_7254,N_7548);
and U8833 (N_8833,N_7615,N_7788);
nand U8834 (N_8834,N_7199,N_7877);
and U8835 (N_8835,N_7020,N_7888);
or U8836 (N_8836,N_7207,N_7515);
or U8837 (N_8837,N_7149,N_7177);
or U8838 (N_8838,N_7719,N_7057);
or U8839 (N_8839,N_7978,N_7177);
nor U8840 (N_8840,N_7966,N_7465);
or U8841 (N_8841,N_7872,N_7321);
nand U8842 (N_8842,N_7595,N_7356);
or U8843 (N_8843,N_7721,N_7379);
nor U8844 (N_8844,N_7285,N_7086);
and U8845 (N_8845,N_7968,N_7582);
and U8846 (N_8846,N_7844,N_7387);
nand U8847 (N_8847,N_7709,N_7286);
nand U8848 (N_8848,N_7251,N_7558);
and U8849 (N_8849,N_7315,N_7212);
nand U8850 (N_8850,N_7720,N_7963);
or U8851 (N_8851,N_7996,N_7327);
and U8852 (N_8852,N_7591,N_7273);
nor U8853 (N_8853,N_7740,N_7806);
nor U8854 (N_8854,N_7662,N_7202);
nand U8855 (N_8855,N_7964,N_7616);
or U8856 (N_8856,N_7258,N_7830);
and U8857 (N_8857,N_7030,N_7049);
nand U8858 (N_8858,N_7166,N_7223);
or U8859 (N_8859,N_7827,N_7208);
and U8860 (N_8860,N_7128,N_7831);
nand U8861 (N_8861,N_7071,N_7440);
and U8862 (N_8862,N_7233,N_7470);
and U8863 (N_8863,N_7548,N_7021);
and U8864 (N_8864,N_7454,N_7565);
and U8865 (N_8865,N_7086,N_7721);
or U8866 (N_8866,N_7463,N_7522);
and U8867 (N_8867,N_7314,N_7275);
nand U8868 (N_8868,N_7079,N_7605);
nand U8869 (N_8869,N_7424,N_7585);
or U8870 (N_8870,N_7845,N_7514);
nand U8871 (N_8871,N_7161,N_7625);
and U8872 (N_8872,N_7626,N_7781);
nor U8873 (N_8873,N_7027,N_7747);
nand U8874 (N_8874,N_7531,N_7173);
nor U8875 (N_8875,N_7569,N_7890);
nor U8876 (N_8876,N_7628,N_7165);
and U8877 (N_8877,N_7170,N_7723);
nand U8878 (N_8878,N_7136,N_7738);
or U8879 (N_8879,N_7726,N_7997);
and U8880 (N_8880,N_7292,N_7136);
nor U8881 (N_8881,N_7803,N_7516);
nand U8882 (N_8882,N_7373,N_7926);
nor U8883 (N_8883,N_7647,N_7663);
nor U8884 (N_8884,N_7224,N_7301);
nand U8885 (N_8885,N_7405,N_7581);
or U8886 (N_8886,N_7769,N_7026);
nor U8887 (N_8887,N_7586,N_7345);
nor U8888 (N_8888,N_7919,N_7494);
nor U8889 (N_8889,N_7627,N_7120);
or U8890 (N_8890,N_7635,N_7886);
nor U8891 (N_8891,N_7814,N_7585);
nor U8892 (N_8892,N_7227,N_7381);
or U8893 (N_8893,N_7762,N_7215);
or U8894 (N_8894,N_7662,N_7573);
nor U8895 (N_8895,N_7014,N_7726);
or U8896 (N_8896,N_7830,N_7412);
or U8897 (N_8897,N_7830,N_7692);
nor U8898 (N_8898,N_7052,N_7989);
or U8899 (N_8899,N_7461,N_7586);
nand U8900 (N_8900,N_7926,N_7102);
and U8901 (N_8901,N_7944,N_7440);
nand U8902 (N_8902,N_7746,N_7932);
and U8903 (N_8903,N_7390,N_7263);
and U8904 (N_8904,N_7210,N_7738);
nor U8905 (N_8905,N_7328,N_7705);
nor U8906 (N_8906,N_7917,N_7174);
or U8907 (N_8907,N_7090,N_7224);
and U8908 (N_8908,N_7046,N_7484);
and U8909 (N_8909,N_7147,N_7547);
nand U8910 (N_8910,N_7396,N_7246);
or U8911 (N_8911,N_7905,N_7131);
nand U8912 (N_8912,N_7714,N_7483);
nor U8913 (N_8913,N_7014,N_7152);
nand U8914 (N_8914,N_7975,N_7861);
or U8915 (N_8915,N_7040,N_7713);
nand U8916 (N_8916,N_7284,N_7380);
nor U8917 (N_8917,N_7785,N_7324);
nor U8918 (N_8918,N_7662,N_7825);
nand U8919 (N_8919,N_7245,N_7832);
nor U8920 (N_8920,N_7243,N_7609);
nand U8921 (N_8921,N_7554,N_7634);
nand U8922 (N_8922,N_7957,N_7421);
or U8923 (N_8923,N_7426,N_7456);
and U8924 (N_8924,N_7976,N_7446);
and U8925 (N_8925,N_7402,N_7636);
and U8926 (N_8926,N_7547,N_7409);
nor U8927 (N_8927,N_7639,N_7464);
and U8928 (N_8928,N_7442,N_7204);
or U8929 (N_8929,N_7223,N_7091);
nand U8930 (N_8930,N_7604,N_7921);
and U8931 (N_8931,N_7804,N_7021);
or U8932 (N_8932,N_7986,N_7465);
nand U8933 (N_8933,N_7737,N_7448);
nor U8934 (N_8934,N_7976,N_7874);
and U8935 (N_8935,N_7758,N_7543);
nor U8936 (N_8936,N_7501,N_7525);
and U8937 (N_8937,N_7206,N_7797);
nor U8938 (N_8938,N_7928,N_7598);
nor U8939 (N_8939,N_7470,N_7932);
nand U8940 (N_8940,N_7656,N_7045);
nand U8941 (N_8941,N_7082,N_7814);
or U8942 (N_8942,N_7663,N_7066);
or U8943 (N_8943,N_7001,N_7894);
and U8944 (N_8944,N_7642,N_7202);
or U8945 (N_8945,N_7858,N_7497);
and U8946 (N_8946,N_7005,N_7083);
nand U8947 (N_8947,N_7674,N_7781);
or U8948 (N_8948,N_7899,N_7777);
or U8949 (N_8949,N_7868,N_7645);
or U8950 (N_8950,N_7961,N_7463);
and U8951 (N_8951,N_7961,N_7053);
nor U8952 (N_8952,N_7447,N_7945);
nor U8953 (N_8953,N_7700,N_7119);
nor U8954 (N_8954,N_7096,N_7029);
nand U8955 (N_8955,N_7924,N_7648);
and U8956 (N_8956,N_7285,N_7786);
nand U8957 (N_8957,N_7233,N_7429);
and U8958 (N_8958,N_7550,N_7164);
or U8959 (N_8959,N_7741,N_7166);
or U8960 (N_8960,N_7180,N_7786);
or U8961 (N_8961,N_7491,N_7739);
nor U8962 (N_8962,N_7308,N_7363);
nor U8963 (N_8963,N_7430,N_7474);
and U8964 (N_8964,N_7544,N_7179);
and U8965 (N_8965,N_7142,N_7787);
nor U8966 (N_8966,N_7272,N_7814);
or U8967 (N_8967,N_7203,N_7640);
nor U8968 (N_8968,N_7138,N_7300);
and U8969 (N_8969,N_7209,N_7482);
nand U8970 (N_8970,N_7496,N_7300);
or U8971 (N_8971,N_7434,N_7675);
or U8972 (N_8972,N_7283,N_7152);
nand U8973 (N_8973,N_7799,N_7836);
nand U8974 (N_8974,N_7884,N_7304);
and U8975 (N_8975,N_7831,N_7006);
and U8976 (N_8976,N_7689,N_7035);
nor U8977 (N_8977,N_7319,N_7341);
nor U8978 (N_8978,N_7207,N_7401);
and U8979 (N_8979,N_7764,N_7523);
or U8980 (N_8980,N_7564,N_7846);
and U8981 (N_8981,N_7279,N_7128);
or U8982 (N_8982,N_7254,N_7327);
or U8983 (N_8983,N_7950,N_7566);
or U8984 (N_8984,N_7003,N_7417);
or U8985 (N_8985,N_7240,N_7844);
and U8986 (N_8986,N_7000,N_7254);
and U8987 (N_8987,N_7191,N_7056);
and U8988 (N_8988,N_7403,N_7465);
nor U8989 (N_8989,N_7710,N_7571);
and U8990 (N_8990,N_7372,N_7984);
or U8991 (N_8991,N_7194,N_7005);
nand U8992 (N_8992,N_7967,N_7949);
or U8993 (N_8993,N_7472,N_7596);
or U8994 (N_8994,N_7895,N_7766);
nand U8995 (N_8995,N_7014,N_7828);
nor U8996 (N_8996,N_7501,N_7857);
or U8997 (N_8997,N_7173,N_7369);
nor U8998 (N_8998,N_7038,N_7277);
nor U8999 (N_8999,N_7387,N_7775);
or U9000 (N_9000,N_8330,N_8417);
or U9001 (N_9001,N_8016,N_8618);
nand U9002 (N_9002,N_8190,N_8071);
nor U9003 (N_9003,N_8400,N_8283);
or U9004 (N_9004,N_8224,N_8165);
and U9005 (N_9005,N_8461,N_8835);
and U9006 (N_9006,N_8183,N_8667);
and U9007 (N_9007,N_8407,N_8264);
nand U9008 (N_9008,N_8997,N_8064);
nand U9009 (N_9009,N_8120,N_8536);
nor U9010 (N_9010,N_8669,N_8037);
and U9011 (N_9011,N_8068,N_8988);
and U9012 (N_9012,N_8313,N_8180);
or U9013 (N_9013,N_8854,N_8742);
and U9014 (N_9014,N_8754,N_8333);
nor U9015 (N_9015,N_8355,N_8289);
and U9016 (N_9016,N_8615,N_8307);
nand U9017 (N_9017,N_8746,N_8455);
and U9018 (N_9018,N_8665,N_8865);
or U9019 (N_9019,N_8427,N_8406);
and U9020 (N_9020,N_8714,N_8610);
or U9021 (N_9021,N_8537,N_8114);
or U9022 (N_9022,N_8431,N_8270);
and U9023 (N_9023,N_8682,N_8050);
and U9024 (N_9024,N_8998,N_8634);
nor U9025 (N_9025,N_8918,N_8317);
or U9026 (N_9026,N_8859,N_8823);
nand U9027 (N_9027,N_8477,N_8342);
nand U9028 (N_9028,N_8545,N_8240);
and U9029 (N_9029,N_8167,N_8077);
nand U9030 (N_9030,N_8948,N_8767);
or U9031 (N_9031,N_8853,N_8149);
or U9032 (N_9032,N_8848,N_8761);
nor U9033 (N_9033,N_8556,N_8834);
and U9034 (N_9034,N_8715,N_8907);
nor U9035 (N_9035,N_8097,N_8329);
or U9036 (N_9036,N_8412,N_8643);
nor U9037 (N_9037,N_8015,N_8124);
nor U9038 (N_9038,N_8301,N_8891);
or U9039 (N_9039,N_8992,N_8365);
nand U9040 (N_9040,N_8334,N_8182);
or U9041 (N_9041,N_8532,N_8815);
or U9042 (N_9042,N_8631,N_8135);
or U9043 (N_9043,N_8189,N_8011);
nand U9044 (N_9044,N_8936,N_8446);
or U9045 (N_9045,N_8248,N_8499);
nor U9046 (N_9046,N_8995,N_8121);
nor U9047 (N_9047,N_8625,N_8425);
or U9048 (N_9048,N_8193,N_8373);
nand U9049 (N_9049,N_8292,N_8328);
and U9050 (N_9050,N_8519,N_8405);
nor U9051 (N_9051,N_8977,N_8156);
nand U9052 (N_9052,N_8382,N_8402);
nand U9053 (N_9053,N_8842,N_8586);
or U9054 (N_9054,N_8778,N_8459);
nor U9055 (N_9055,N_8020,N_8900);
nor U9056 (N_9056,N_8582,N_8398);
nor U9057 (N_9057,N_8058,N_8086);
and U9058 (N_9058,N_8435,N_8639);
or U9059 (N_9059,N_8718,N_8901);
or U9060 (N_9060,N_8929,N_8876);
or U9061 (N_9061,N_8690,N_8249);
nand U9062 (N_9062,N_8739,N_8698);
and U9063 (N_9063,N_8055,N_8242);
and U9064 (N_9064,N_8560,N_8442);
nand U9065 (N_9065,N_8115,N_8934);
nor U9066 (N_9066,N_8557,N_8027);
nor U9067 (N_9067,N_8042,N_8724);
and U9068 (N_9068,N_8443,N_8561);
nor U9069 (N_9069,N_8388,N_8451);
nor U9070 (N_9070,N_8510,N_8445);
nand U9071 (N_9071,N_8155,N_8535);
or U9072 (N_9072,N_8655,N_8873);
nor U9073 (N_9073,N_8662,N_8187);
nand U9074 (N_9074,N_8090,N_8810);
or U9075 (N_9075,N_8401,N_8460);
or U9076 (N_9076,N_8512,N_8766);
xnor U9077 (N_9077,N_8757,N_8697);
or U9078 (N_9078,N_8544,N_8421);
nor U9079 (N_9079,N_8980,N_8983);
nor U9080 (N_9080,N_8214,N_8009);
nor U9081 (N_9081,N_8517,N_8701);
nand U9082 (N_9082,N_8311,N_8419);
nand U9083 (N_9083,N_8158,N_8202);
nor U9084 (N_9084,N_8483,N_8308);
and U9085 (N_9085,N_8890,N_8023);
nor U9086 (N_9086,N_8775,N_8740);
nor U9087 (N_9087,N_8881,N_8862);
or U9088 (N_9088,N_8833,N_8973);
nor U9089 (N_9089,N_8103,N_8143);
nor U9090 (N_9090,N_8604,N_8474);
nand U9091 (N_9091,N_8837,N_8237);
or U9092 (N_9092,N_8319,N_8347);
and U9093 (N_9093,N_8954,N_8142);
and U9094 (N_9094,N_8717,N_8014);
or U9095 (N_9095,N_8856,N_8990);
nor U9096 (N_9096,N_8392,N_8683);
nor U9097 (N_9097,N_8257,N_8993);
or U9098 (N_9098,N_8589,N_8246);
nor U9099 (N_9099,N_8112,N_8039);
nor U9100 (N_9100,N_8895,N_8432);
and U9101 (N_9101,N_8816,N_8469);
nand U9102 (N_9102,N_8032,N_8194);
and U9103 (N_9103,N_8503,N_8827);
or U9104 (N_9104,N_8148,N_8719);
nand U9105 (N_9105,N_8164,N_8747);
and U9106 (N_9106,N_8056,N_8256);
and U9107 (N_9107,N_8260,N_8236);
and U9108 (N_9108,N_8966,N_8919);
or U9109 (N_9109,N_8651,N_8234);
or U9110 (N_9110,N_8358,N_8386);
or U9111 (N_9111,N_8668,N_8571);
nand U9112 (N_9112,N_8024,N_8614);
nand U9113 (N_9113,N_8000,N_8538);
nand U9114 (N_9114,N_8576,N_8920);
or U9115 (N_9115,N_8291,N_8542);
nand U9116 (N_9116,N_8709,N_8626);
nor U9117 (N_9117,N_8134,N_8213);
nor U9118 (N_9118,N_8850,N_8838);
nor U9119 (N_9119,N_8822,N_8389);
or U9120 (N_9120,N_8422,N_8831);
nand U9121 (N_9121,N_8423,N_8953);
and U9122 (N_9122,N_8297,N_8686);
or U9123 (N_9123,N_8345,N_8010);
or U9124 (N_9124,N_8507,N_8984);
or U9125 (N_9125,N_8711,N_8905);
or U9126 (N_9126,N_8772,N_8795);
or U9127 (N_9127,N_8318,N_8628);
nor U9128 (N_9128,N_8416,N_8151);
nor U9129 (N_9129,N_8937,N_8551);
nand U9130 (N_9130,N_8339,N_8250);
nor U9131 (N_9131,N_8282,N_8813);
and U9132 (N_9132,N_8547,N_8391);
or U9133 (N_9133,N_8633,N_8241);
nand U9134 (N_9134,N_8267,N_8933);
nor U9135 (N_9135,N_8426,N_8684);
nand U9136 (N_9136,N_8284,N_8734);
nor U9137 (N_9137,N_8921,N_8758);
nand U9138 (N_9138,N_8553,N_8482);
or U9139 (N_9139,N_8844,N_8072);
nand U9140 (N_9140,N_8087,N_8521);
nand U9141 (N_9141,N_8916,N_8029);
xnor U9142 (N_9142,N_8206,N_8491);
and U9143 (N_9143,N_8229,N_8981);
or U9144 (N_9144,N_8368,N_8570);
and U9145 (N_9145,N_8679,N_8897);
or U9146 (N_9146,N_8587,N_8073);
nand U9147 (N_9147,N_8108,N_8777);
and U9148 (N_9148,N_8498,N_8550);
and U9149 (N_9149,N_8380,N_8192);
or U9150 (N_9150,N_8909,N_8958);
nand U9151 (N_9151,N_8475,N_8262);
nand U9152 (N_9152,N_8930,N_8565);
or U9153 (N_9153,N_8395,N_8473);
nor U9154 (N_9154,N_8776,N_8502);
or U9155 (N_9155,N_8809,N_8326);
and U9156 (N_9156,N_8244,N_8843);
or U9157 (N_9157,N_8573,N_8962);
nand U9158 (N_9158,N_8955,N_8152);
or U9159 (N_9159,N_8575,N_8659);
and U9160 (N_9160,N_8996,N_8741);
and U9161 (N_9161,N_8341,N_8799);
nand U9162 (N_9162,N_8638,N_8723);
and U9163 (N_9163,N_8803,N_8069);
nor U9164 (N_9164,N_8913,N_8526);
nor U9165 (N_9165,N_8172,N_8566);
or U9166 (N_9166,N_8923,N_8627);
nand U9167 (N_9167,N_8893,N_8336);
nor U9168 (N_9168,N_8774,N_8074);
nor U9169 (N_9169,N_8279,N_8525);
or U9170 (N_9170,N_8485,N_8140);
nor U9171 (N_9171,N_8075,N_8232);
nand U9172 (N_9172,N_8153,N_8971);
or U9173 (N_9173,N_8790,N_8581);
nand U9174 (N_9174,N_8527,N_8621);
nor U9175 (N_9175,N_8028,N_8607);
nor U9176 (N_9176,N_8814,N_8534);
nand U9177 (N_9177,N_8548,N_8195);
or U9178 (N_9178,N_8082,N_8888);
nor U9179 (N_9179,N_8511,N_8572);
nor U9180 (N_9180,N_8013,N_8820);
or U9181 (N_9181,N_8356,N_8044);
nor U9182 (N_9182,N_8902,N_8127);
or U9183 (N_9183,N_8314,N_8070);
nor U9184 (N_9184,N_8462,N_8784);
and U9185 (N_9185,N_8166,N_8418);
nor U9186 (N_9186,N_8749,N_8440);
nor U9187 (N_9187,N_8982,N_8706);
and U9188 (N_9188,N_8695,N_8825);
and U9189 (N_9189,N_8969,N_8611);
nand U9190 (N_9190,N_8231,N_8309);
or U9191 (N_9191,N_8600,N_8751);
and U9192 (N_9192,N_8605,N_8978);
nor U9193 (N_9193,N_8871,N_8340);
or U9194 (N_9194,N_8119,N_8145);
and U9195 (N_9195,N_8107,N_8179);
or U9196 (N_9196,N_8671,N_8131);
or U9197 (N_9197,N_8006,N_8062);
nand U9198 (N_9198,N_8692,N_8568);
or U9199 (N_9199,N_8926,N_8490);
or U9200 (N_9200,N_8084,N_8579);
and U9201 (N_9201,N_8051,N_8468);
or U9202 (N_9202,N_8259,N_8322);
nor U9203 (N_9203,N_8298,N_8209);
or U9204 (N_9204,N_8851,N_8805);
nor U9205 (N_9205,N_8922,N_8253);
and U9206 (N_9206,N_8606,N_8932);
nand U9207 (N_9207,N_8704,N_8592);
nand U9208 (N_9208,N_8663,N_8759);
and U9209 (N_9209,N_8176,N_8049);
nor U9210 (N_9210,N_8635,N_8360);
and U9211 (N_9211,N_8812,N_8808);
nor U9212 (N_9212,N_8530,N_8130);
and U9213 (N_9213,N_8904,N_8448);
and U9214 (N_9214,N_8046,N_8221);
or U9215 (N_9215,N_8273,N_8181);
or U9216 (N_9216,N_8867,N_8660);
nor U9217 (N_9217,N_8409,N_8162);
nor U9218 (N_9218,N_8100,N_8454);
nand U9219 (N_9219,N_8523,N_8546);
or U9220 (N_9220,N_8303,N_8396);
nor U9221 (N_9221,N_8722,N_8641);
nand U9222 (N_9222,N_8495,N_8122);
nor U9223 (N_9223,N_8590,N_8312);
nor U9224 (N_9224,N_8999,N_8238);
or U9225 (N_9225,N_8732,N_8911);
nand U9226 (N_9226,N_8057,N_8063);
and U9227 (N_9227,N_8949,N_8925);
and U9228 (N_9228,N_8346,N_8956);
and U9229 (N_9229,N_8497,N_8529);
or U9230 (N_9230,N_8293,N_8496);
and U9231 (N_9231,N_8840,N_8569);
nor U9232 (N_9232,N_8378,N_8593);
nand U9233 (N_9233,N_8894,N_8323);
nor U9234 (N_9234,N_8787,N_8185);
or U9235 (N_9235,N_8824,N_8096);
and U9236 (N_9236,N_8687,N_8332);
nor U9237 (N_9237,N_8296,N_8728);
nand U9238 (N_9238,N_8696,N_8136);
xor U9239 (N_9239,N_8559,N_8645);
nor U9240 (N_9240,N_8233,N_8744);
and U9241 (N_9241,N_8694,N_8059);
nand U9242 (N_9242,N_8337,N_8670);
nor U9243 (N_9243,N_8048,N_8258);
nor U9244 (N_9244,N_8830,N_8254);
or U9245 (N_9245,N_8963,N_8961);
and U9246 (N_9246,N_8678,N_8005);
nor U9247 (N_9247,N_8452,N_8630);
nand U9248 (N_9248,N_8101,N_8617);
and U9249 (N_9249,N_8225,N_8287);
nand U9250 (N_9250,N_8672,N_8047);
nand U9251 (N_9251,N_8272,N_8945);
nand U9252 (N_9252,N_8410,N_8492);
or U9253 (N_9253,N_8622,N_8624);
nor U9254 (N_9254,N_8789,N_8796);
or U9255 (N_9255,N_8792,N_8596);
nor U9256 (N_9256,N_8003,N_8434);
and U9257 (N_9257,N_8736,N_8354);
nand U9258 (N_9258,N_8616,N_8489);
nand U9259 (N_9259,N_8285,N_8125);
or U9260 (N_9260,N_8729,N_8102);
nand U9261 (N_9261,N_8163,N_8227);
and U9262 (N_9262,N_8889,N_8760);
nand U9263 (N_9263,N_8266,N_8699);
nor U9264 (N_9264,N_8737,N_8716);
or U9265 (N_9265,N_8745,N_8078);
nand U9266 (N_9266,N_8369,N_8243);
or U9267 (N_9267,N_8861,N_8201);
nand U9268 (N_9268,N_8217,N_8159);
and U9269 (N_9269,N_8880,N_8806);
or U9270 (N_9270,N_8801,N_8637);
nor U9271 (N_9271,N_8280,N_8769);
or U9272 (N_9272,N_8105,N_8450);
nand U9273 (N_9273,N_8478,N_8883);
nand U9274 (N_9274,N_8447,N_8677);
nor U9275 (N_9275,N_8268,N_8807);
nor U9276 (N_9276,N_8661,N_8199);
xnor U9277 (N_9277,N_8362,N_8457);
and U9278 (N_9278,N_8886,N_8642);
and U9279 (N_9279,N_8379,N_8174);
nor U9280 (N_9280,N_8390,N_8852);
or U9281 (N_9281,N_8403,N_8481);
and U9282 (N_9282,N_8088,N_8196);
nor U9283 (N_9283,N_8674,N_8353);
and U9284 (N_9284,N_8504,N_8821);
nand U9285 (N_9285,N_8691,N_8374);
nor U9286 (N_9286,N_8278,N_8411);
or U9287 (N_9287,N_8666,N_8035);
nor U9288 (N_9288,N_8066,N_8316);
or U9289 (N_9289,N_8574,N_8914);
nor U9290 (N_9290,N_8750,N_8549);
and U9291 (N_9291,N_8315,N_8212);
nor U9292 (N_9292,N_8493,N_8438);
nand U9293 (N_9293,N_8584,N_8466);
nor U9294 (N_9294,N_8397,N_8177);
or U9295 (N_9295,N_8869,N_8171);
nand U9296 (N_9296,N_8210,N_8974);
nand U9297 (N_9297,N_8205,N_8636);
and U9298 (N_9298,N_8271,N_8786);
nand U9299 (N_9299,N_8693,N_8522);
nor U9300 (N_9300,N_8743,N_8832);
and U9301 (N_9301,N_8783,N_8748);
nand U9302 (N_9302,N_8720,N_8846);
or U9303 (N_9303,N_8294,N_8092);
nand U9304 (N_9304,N_8884,N_8972);
and U9305 (N_9305,N_8619,N_8847);
or U9306 (N_9306,N_8300,N_8111);
and U9307 (N_9307,N_8408,N_8970);
or U9308 (N_9308,N_8026,N_8022);
nor U9309 (N_9309,N_8924,N_8877);
or U9310 (N_9310,N_8220,N_8351);
nand U9311 (N_9311,N_8518,N_8290);
or U9312 (N_9312,N_8175,N_8915);
nor U9313 (N_9313,N_8836,N_8531);
or U9314 (N_9314,N_8343,N_8735);
or U9315 (N_9315,N_8321,N_8083);
or U9316 (N_9316,N_8539,N_8726);
and U9317 (N_9317,N_8817,N_8857);
or U9318 (N_9318,N_8501,N_8415);
nand U9319 (N_9319,N_8479,N_8987);
nand U9320 (N_9320,N_8208,N_8506);
or U9321 (N_9321,N_8578,N_8960);
or U9322 (N_9322,N_8344,N_8331);
or U9323 (N_9323,N_8045,N_8053);
or U9324 (N_9324,N_8959,N_8874);
and U9325 (N_9325,N_8458,N_8826);
nor U9326 (N_9326,N_8819,N_8094);
and U9327 (N_9327,N_8223,N_8689);
or U9328 (N_9328,N_8128,N_8095);
and U9329 (N_9329,N_8520,N_8043);
or U9330 (N_9330,N_8038,N_8533);
nor U9331 (N_9331,N_8173,N_8839);
and U9332 (N_9332,N_8310,N_8912);
nand U9333 (N_9333,N_8899,N_8733);
and U9334 (N_9334,N_8146,N_8986);
nor U9335 (N_9335,N_8306,N_8387);
or U9336 (N_9336,N_8603,N_8444);
or U9337 (N_9337,N_8994,N_8991);
and U9338 (N_9338,N_8305,N_8878);
nand U9339 (N_9339,N_8335,N_8424);
nor U9340 (N_9340,N_8376,N_8942);
nor U9341 (N_9341,N_8935,N_8872);
nor U9342 (N_9342,N_8060,N_8941);
or U9343 (N_9343,N_8106,N_8648);
nor U9344 (N_9344,N_8773,N_8371);
nor U9345 (N_9345,N_8467,N_8255);
nor U9346 (N_9346,N_8203,N_8472);
or U9347 (N_9347,N_8800,N_8275);
nor U9348 (N_9348,N_8126,N_8765);
nand U9349 (N_9349,N_8791,N_8730);
and U9350 (N_9350,N_8989,N_8154);
or U9351 (N_9351,N_8613,N_8099);
or U9352 (N_9352,N_8178,N_8012);
or U9353 (N_9353,N_8656,N_8286);
nor U9354 (N_9354,N_8947,N_8967);
nand U9355 (N_9355,N_8110,N_8700);
and U9356 (N_9356,N_8067,N_8357);
and U9357 (N_9357,N_8802,N_8620);
nand U9358 (N_9358,N_8008,N_8609);
nand U9359 (N_9359,N_8041,N_8150);
or U9360 (N_9360,N_8864,N_8456);
nor U9361 (N_9361,N_8211,N_8104);
nand U9362 (N_9362,N_8384,N_8780);
nor U9363 (N_9363,N_8002,N_8144);
nor U9364 (N_9364,N_8160,N_8222);
nor U9365 (N_9365,N_8885,N_8430);
nand U9366 (N_9366,N_8429,N_8188);
and U9367 (N_9367,N_8191,N_8855);
or U9368 (N_9368,N_8752,N_8034);
and U9369 (N_9369,N_8261,N_8404);
and U9370 (N_9370,N_8602,N_8428);
or U9371 (N_9371,N_8361,N_8712);
nand U9372 (N_9372,N_8681,N_8580);
and U9373 (N_9373,N_8868,N_8950);
nand U9374 (N_9374,N_8509,N_8139);
nor U9375 (N_9375,N_8348,N_8327);
and U9376 (N_9376,N_8965,N_8299);
nor U9377 (N_9377,N_8653,N_8141);
or U9378 (N_9378,N_8702,N_8598);
or U9379 (N_9379,N_8705,N_8184);
or U9380 (N_9380,N_8594,N_8957);
nand U9381 (N_9381,N_8359,N_8505);
or U9382 (N_9382,N_8540,N_8230);
nor U9383 (N_9383,N_8710,N_8928);
and U9384 (N_9384,N_8599,N_8875);
or U9385 (N_9385,N_8870,N_8555);
nand U9386 (N_9386,N_8860,N_8463);
or U9387 (N_9387,N_8471,N_8938);
and U9388 (N_9388,N_8004,N_8516);
or U9389 (N_9389,N_8845,N_8943);
nor U9390 (N_9390,N_8033,N_8054);
and U9391 (N_9391,N_8138,N_8541);
and U9392 (N_9392,N_8393,N_8528);
and U9393 (N_9393,N_8436,N_8939);
nor U9394 (N_9394,N_8370,N_8325);
nand U9395 (N_9395,N_8975,N_8567);
and U9396 (N_9396,N_8324,N_8508);
or U9397 (N_9397,N_8768,N_8725);
and U9398 (N_9398,N_8779,N_8216);
nand U9399 (N_9399,N_8025,N_8274);
or U9400 (N_9400,N_8763,N_8887);
nor U9401 (N_9401,N_8065,N_8818);
nand U9402 (N_9402,N_8794,N_8277);
nor U9403 (N_9403,N_8788,N_8204);
nor U9404 (N_9404,N_8487,N_8964);
and U9405 (N_9405,N_8879,N_8713);
nand U9406 (N_9406,N_8021,N_8375);
or U9407 (N_9407,N_8931,N_8944);
and U9408 (N_9408,N_8811,N_8976);
and U9409 (N_9409,N_8755,N_8951);
or U9410 (N_9410,N_8771,N_8673);
nand U9411 (N_9411,N_8927,N_8654);
nand U9412 (N_9412,N_8018,N_8601);
and U9413 (N_9413,N_8782,N_8001);
nand U9414 (N_9414,N_8708,N_8030);
nor U9415 (N_9415,N_8168,N_8414);
nand U9416 (N_9416,N_8089,N_8500);
or U9417 (N_9417,N_8132,N_8770);
nand U9418 (N_9418,N_8437,N_8215);
or U9419 (N_9419,N_8762,N_8372);
nand U9420 (N_9420,N_8882,N_8363);
and U9421 (N_9421,N_8804,N_8169);
or U9422 (N_9422,N_8946,N_8513);
and U9423 (N_9423,N_8892,N_8383);
nand U9424 (N_9424,N_8465,N_8828);
and U9425 (N_9425,N_8595,N_8543);
nand U9426 (N_9426,N_8664,N_8798);
nand U9427 (N_9427,N_8198,N_8688);
and U9428 (N_9428,N_8113,N_8484);
or U9429 (N_9429,N_8652,N_8377);
nand U9430 (N_9430,N_8228,N_8583);
nand U9431 (N_9431,N_8197,N_8908);
nand U9432 (N_9432,N_8118,N_8076);
nor U9433 (N_9433,N_8186,N_8849);
nor U9434 (N_9434,N_8680,N_8764);
nor U9435 (N_9435,N_8281,N_8721);
and U9436 (N_9436,N_8480,N_8453);
nand U9437 (N_9437,N_8394,N_8170);
or U9438 (N_9438,N_8588,N_8133);
nor U9439 (N_9439,N_8439,N_8263);
nor U9440 (N_9440,N_8420,N_8036);
and U9441 (N_9441,N_8367,N_8081);
or U9442 (N_9442,N_8650,N_8200);
and U9443 (N_9443,N_8399,N_8226);
and U9444 (N_9444,N_8910,N_8563);
nor U9445 (N_9445,N_8629,N_8640);
nor U9446 (N_9446,N_8433,N_8207);
nand U9447 (N_9447,N_8269,N_8738);
nor U9448 (N_9448,N_8123,N_8157);
and U9449 (N_9449,N_8657,N_8320);
and U9450 (N_9450,N_8219,N_8829);
or U9451 (N_9451,N_8239,N_8117);
or U9452 (N_9452,N_8350,N_8903);
and U9453 (N_9453,N_8093,N_8441);
or U9454 (N_9454,N_8040,N_8952);
and U9455 (N_9455,N_8449,N_8476);
nor U9456 (N_9456,N_8288,N_8858);
nor U9457 (N_9457,N_8863,N_8302);
nand U9458 (N_9458,N_8797,N_8079);
or U9459 (N_9459,N_8098,N_8017);
nand U9460 (N_9460,N_8080,N_8753);
nand U9461 (N_9461,N_8304,N_8116);
nand U9462 (N_9462,N_8658,N_8649);
and U9463 (N_9463,N_8091,N_8514);
nand U9464 (N_9464,N_8245,N_8488);
nor U9465 (N_9465,N_8793,N_8413);
nor U9466 (N_9466,N_8727,N_8585);
or U9467 (N_9467,N_8486,N_8218);
or U9468 (N_9468,N_8917,N_8608);
nand U9469 (N_9469,N_8494,N_8338);
nand U9470 (N_9470,N_8464,N_8896);
nand U9471 (N_9471,N_8597,N_8554);
nor U9472 (N_9472,N_8676,N_8364);
nand U9473 (N_9473,N_8235,N_8979);
and U9474 (N_9474,N_8906,N_8781);
nand U9475 (N_9475,N_8756,N_8109);
nand U9476 (N_9476,N_8524,N_8558);
nand U9477 (N_9477,N_8612,N_8985);
nand U9478 (N_9478,N_8731,N_8940);
or U9479 (N_9479,N_8381,N_8675);
or U9480 (N_9480,N_8061,N_8552);
or U9481 (N_9481,N_8265,N_8515);
or U9482 (N_9482,N_8147,N_8785);
and U9483 (N_9483,N_8647,N_8385);
nor U9484 (N_9484,N_8685,N_8247);
nor U9485 (N_9485,N_8031,N_8644);
nand U9486 (N_9486,N_8707,N_8562);
or U9487 (N_9487,N_8968,N_8085);
nor U9488 (N_9488,N_8019,N_8646);
or U9489 (N_9489,N_8898,N_8295);
or U9490 (N_9490,N_8349,N_8252);
or U9491 (N_9491,N_8161,N_8841);
nor U9492 (N_9492,N_8577,N_8276);
nor U9493 (N_9493,N_8866,N_8470);
nand U9494 (N_9494,N_8591,N_8703);
nand U9495 (N_9495,N_8251,N_8007);
and U9496 (N_9496,N_8564,N_8052);
or U9497 (N_9497,N_8623,N_8137);
nor U9498 (N_9498,N_8366,N_8129);
nor U9499 (N_9499,N_8632,N_8352);
nor U9500 (N_9500,N_8920,N_8124);
xor U9501 (N_9501,N_8651,N_8615);
and U9502 (N_9502,N_8425,N_8088);
or U9503 (N_9503,N_8867,N_8269);
or U9504 (N_9504,N_8864,N_8221);
or U9505 (N_9505,N_8710,N_8230);
nand U9506 (N_9506,N_8826,N_8959);
nand U9507 (N_9507,N_8310,N_8751);
and U9508 (N_9508,N_8239,N_8747);
nand U9509 (N_9509,N_8331,N_8485);
or U9510 (N_9510,N_8768,N_8239);
nor U9511 (N_9511,N_8087,N_8992);
nand U9512 (N_9512,N_8121,N_8119);
nand U9513 (N_9513,N_8615,N_8325);
and U9514 (N_9514,N_8262,N_8973);
nand U9515 (N_9515,N_8957,N_8081);
nand U9516 (N_9516,N_8799,N_8390);
and U9517 (N_9517,N_8752,N_8021);
nor U9518 (N_9518,N_8537,N_8744);
or U9519 (N_9519,N_8741,N_8376);
or U9520 (N_9520,N_8742,N_8551);
and U9521 (N_9521,N_8922,N_8443);
nand U9522 (N_9522,N_8404,N_8883);
and U9523 (N_9523,N_8189,N_8621);
nand U9524 (N_9524,N_8269,N_8060);
nand U9525 (N_9525,N_8888,N_8680);
or U9526 (N_9526,N_8864,N_8091);
nand U9527 (N_9527,N_8166,N_8408);
or U9528 (N_9528,N_8287,N_8006);
nand U9529 (N_9529,N_8498,N_8975);
and U9530 (N_9530,N_8761,N_8272);
and U9531 (N_9531,N_8696,N_8836);
or U9532 (N_9532,N_8637,N_8286);
or U9533 (N_9533,N_8071,N_8240);
nor U9534 (N_9534,N_8339,N_8975);
and U9535 (N_9535,N_8131,N_8345);
nand U9536 (N_9536,N_8901,N_8848);
or U9537 (N_9537,N_8521,N_8726);
nand U9538 (N_9538,N_8752,N_8400);
nor U9539 (N_9539,N_8205,N_8425);
or U9540 (N_9540,N_8902,N_8045);
and U9541 (N_9541,N_8660,N_8107);
nor U9542 (N_9542,N_8822,N_8364);
nor U9543 (N_9543,N_8485,N_8458);
nand U9544 (N_9544,N_8685,N_8729);
nand U9545 (N_9545,N_8401,N_8619);
and U9546 (N_9546,N_8121,N_8036);
nand U9547 (N_9547,N_8104,N_8583);
nand U9548 (N_9548,N_8772,N_8594);
nand U9549 (N_9549,N_8877,N_8057);
nand U9550 (N_9550,N_8444,N_8014);
nand U9551 (N_9551,N_8918,N_8542);
or U9552 (N_9552,N_8360,N_8647);
nand U9553 (N_9553,N_8080,N_8891);
and U9554 (N_9554,N_8663,N_8797);
and U9555 (N_9555,N_8835,N_8173);
or U9556 (N_9556,N_8741,N_8666);
and U9557 (N_9557,N_8596,N_8605);
or U9558 (N_9558,N_8292,N_8287);
and U9559 (N_9559,N_8850,N_8805);
nor U9560 (N_9560,N_8412,N_8738);
and U9561 (N_9561,N_8551,N_8957);
nor U9562 (N_9562,N_8723,N_8034);
or U9563 (N_9563,N_8573,N_8946);
or U9564 (N_9564,N_8718,N_8174);
nor U9565 (N_9565,N_8467,N_8431);
nor U9566 (N_9566,N_8194,N_8388);
and U9567 (N_9567,N_8617,N_8484);
nand U9568 (N_9568,N_8481,N_8548);
nor U9569 (N_9569,N_8884,N_8153);
or U9570 (N_9570,N_8153,N_8234);
or U9571 (N_9571,N_8056,N_8534);
and U9572 (N_9572,N_8900,N_8492);
or U9573 (N_9573,N_8085,N_8227);
or U9574 (N_9574,N_8230,N_8250);
nand U9575 (N_9575,N_8563,N_8294);
nand U9576 (N_9576,N_8881,N_8753);
nand U9577 (N_9577,N_8837,N_8841);
nor U9578 (N_9578,N_8758,N_8167);
or U9579 (N_9579,N_8614,N_8090);
nand U9580 (N_9580,N_8706,N_8856);
and U9581 (N_9581,N_8039,N_8665);
nor U9582 (N_9582,N_8873,N_8907);
or U9583 (N_9583,N_8688,N_8594);
or U9584 (N_9584,N_8878,N_8564);
and U9585 (N_9585,N_8100,N_8599);
nand U9586 (N_9586,N_8822,N_8018);
or U9587 (N_9587,N_8788,N_8699);
nand U9588 (N_9588,N_8526,N_8784);
and U9589 (N_9589,N_8157,N_8848);
nand U9590 (N_9590,N_8072,N_8412);
and U9591 (N_9591,N_8107,N_8065);
nor U9592 (N_9592,N_8371,N_8586);
and U9593 (N_9593,N_8011,N_8111);
nand U9594 (N_9594,N_8005,N_8636);
or U9595 (N_9595,N_8036,N_8869);
nor U9596 (N_9596,N_8426,N_8768);
or U9597 (N_9597,N_8450,N_8487);
or U9598 (N_9598,N_8410,N_8185);
and U9599 (N_9599,N_8267,N_8603);
or U9600 (N_9600,N_8437,N_8658);
or U9601 (N_9601,N_8754,N_8029);
nor U9602 (N_9602,N_8108,N_8528);
nand U9603 (N_9603,N_8613,N_8892);
nor U9604 (N_9604,N_8651,N_8003);
nand U9605 (N_9605,N_8684,N_8594);
nand U9606 (N_9606,N_8033,N_8950);
and U9607 (N_9607,N_8958,N_8265);
or U9608 (N_9608,N_8894,N_8803);
nor U9609 (N_9609,N_8691,N_8883);
nand U9610 (N_9610,N_8455,N_8650);
nand U9611 (N_9611,N_8580,N_8101);
and U9612 (N_9612,N_8038,N_8785);
or U9613 (N_9613,N_8757,N_8632);
nor U9614 (N_9614,N_8445,N_8442);
nand U9615 (N_9615,N_8339,N_8212);
and U9616 (N_9616,N_8774,N_8499);
nor U9617 (N_9617,N_8017,N_8171);
nor U9618 (N_9618,N_8743,N_8578);
or U9619 (N_9619,N_8991,N_8975);
and U9620 (N_9620,N_8831,N_8605);
nor U9621 (N_9621,N_8935,N_8243);
nor U9622 (N_9622,N_8153,N_8801);
or U9623 (N_9623,N_8966,N_8373);
nand U9624 (N_9624,N_8205,N_8549);
or U9625 (N_9625,N_8405,N_8834);
nand U9626 (N_9626,N_8836,N_8200);
nand U9627 (N_9627,N_8580,N_8137);
nand U9628 (N_9628,N_8677,N_8146);
nand U9629 (N_9629,N_8109,N_8754);
and U9630 (N_9630,N_8672,N_8913);
and U9631 (N_9631,N_8130,N_8714);
or U9632 (N_9632,N_8057,N_8399);
and U9633 (N_9633,N_8302,N_8400);
nand U9634 (N_9634,N_8100,N_8203);
nand U9635 (N_9635,N_8831,N_8748);
nor U9636 (N_9636,N_8651,N_8518);
nor U9637 (N_9637,N_8334,N_8492);
and U9638 (N_9638,N_8360,N_8241);
nand U9639 (N_9639,N_8002,N_8689);
nor U9640 (N_9640,N_8175,N_8309);
or U9641 (N_9641,N_8622,N_8125);
or U9642 (N_9642,N_8179,N_8161);
nand U9643 (N_9643,N_8095,N_8438);
or U9644 (N_9644,N_8735,N_8671);
nor U9645 (N_9645,N_8438,N_8348);
nand U9646 (N_9646,N_8559,N_8910);
nor U9647 (N_9647,N_8688,N_8881);
or U9648 (N_9648,N_8519,N_8279);
nor U9649 (N_9649,N_8568,N_8318);
and U9650 (N_9650,N_8336,N_8962);
or U9651 (N_9651,N_8493,N_8225);
nand U9652 (N_9652,N_8358,N_8272);
or U9653 (N_9653,N_8663,N_8885);
nor U9654 (N_9654,N_8693,N_8410);
and U9655 (N_9655,N_8545,N_8914);
and U9656 (N_9656,N_8617,N_8127);
nor U9657 (N_9657,N_8068,N_8974);
nand U9658 (N_9658,N_8292,N_8140);
or U9659 (N_9659,N_8718,N_8748);
xnor U9660 (N_9660,N_8562,N_8306);
nor U9661 (N_9661,N_8296,N_8764);
or U9662 (N_9662,N_8408,N_8099);
and U9663 (N_9663,N_8674,N_8823);
and U9664 (N_9664,N_8060,N_8204);
nand U9665 (N_9665,N_8666,N_8445);
and U9666 (N_9666,N_8878,N_8883);
or U9667 (N_9667,N_8483,N_8122);
nor U9668 (N_9668,N_8400,N_8380);
nor U9669 (N_9669,N_8265,N_8946);
or U9670 (N_9670,N_8014,N_8589);
or U9671 (N_9671,N_8714,N_8178);
nand U9672 (N_9672,N_8696,N_8202);
or U9673 (N_9673,N_8056,N_8852);
nor U9674 (N_9674,N_8899,N_8563);
or U9675 (N_9675,N_8755,N_8040);
nand U9676 (N_9676,N_8874,N_8077);
nand U9677 (N_9677,N_8941,N_8545);
or U9678 (N_9678,N_8619,N_8635);
or U9679 (N_9679,N_8989,N_8530);
nor U9680 (N_9680,N_8946,N_8807);
and U9681 (N_9681,N_8365,N_8805);
nand U9682 (N_9682,N_8016,N_8632);
or U9683 (N_9683,N_8382,N_8250);
and U9684 (N_9684,N_8275,N_8802);
and U9685 (N_9685,N_8556,N_8745);
and U9686 (N_9686,N_8752,N_8479);
nor U9687 (N_9687,N_8683,N_8676);
nor U9688 (N_9688,N_8658,N_8490);
nand U9689 (N_9689,N_8127,N_8578);
nand U9690 (N_9690,N_8579,N_8364);
nor U9691 (N_9691,N_8856,N_8844);
nor U9692 (N_9692,N_8417,N_8386);
nand U9693 (N_9693,N_8344,N_8095);
nor U9694 (N_9694,N_8862,N_8308);
and U9695 (N_9695,N_8366,N_8103);
or U9696 (N_9696,N_8382,N_8128);
nor U9697 (N_9697,N_8254,N_8612);
nor U9698 (N_9698,N_8042,N_8542);
nor U9699 (N_9699,N_8070,N_8568);
nand U9700 (N_9700,N_8782,N_8817);
or U9701 (N_9701,N_8114,N_8026);
nand U9702 (N_9702,N_8254,N_8779);
and U9703 (N_9703,N_8562,N_8546);
and U9704 (N_9704,N_8017,N_8706);
and U9705 (N_9705,N_8924,N_8630);
and U9706 (N_9706,N_8400,N_8127);
or U9707 (N_9707,N_8657,N_8131);
nor U9708 (N_9708,N_8844,N_8279);
nand U9709 (N_9709,N_8540,N_8240);
and U9710 (N_9710,N_8475,N_8688);
nand U9711 (N_9711,N_8996,N_8038);
nand U9712 (N_9712,N_8600,N_8095);
and U9713 (N_9713,N_8004,N_8221);
or U9714 (N_9714,N_8017,N_8889);
nand U9715 (N_9715,N_8160,N_8784);
xnor U9716 (N_9716,N_8103,N_8529);
and U9717 (N_9717,N_8529,N_8458);
and U9718 (N_9718,N_8015,N_8775);
nand U9719 (N_9719,N_8217,N_8490);
and U9720 (N_9720,N_8095,N_8698);
nor U9721 (N_9721,N_8783,N_8409);
nor U9722 (N_9722,N_8692,N_8826);
nand U9723 (N_9723,N_8009,N_8207);
nor U9724 (N_9724,N_8974,N_8983);
nor U9725 (N_9725,N_8737,N_8401);
or U9726 (N_9726,N_8675,N_8438);
and U9727 (N_9727,N_8542,N_8606);
or U9728 (N_9728,N_8555,N_8284);
nor U9729 (N_9729,N_8739,N_8488);
nand U9730 (N_9730,N_8745,N_8817);
xnor U9731 (N_9731,N_8942,N_8731);
nor U9732 (N_9732,N_8977,N_8295);
nand U9733 (N_9733,N_8957,N_8903);
nor U9734 (N_9734,N_8327,N_8049);
nand U9735 (N_9735,N_8045,N_8331);
or U9736 (N_9736,N_8627,N_8321);
xor U9737 (N_9737,N_8983,N_8161);
nor U9738 (N_9738,N_8370,N_8704);
or U9739 (N_9739,N_8016,N_8750);
nor U9740 (N_9740,N_8341,N_8834);
nor U9741 (N_9741,N_8349,N_8676);
nor U9742 (N_9742,N_8632,N_8390);
nor U9743 (N_9743,N_8827,N_8094);
nand U9744 (N_9744,N_8729,N_8514);
nor U9745 (N_9745,N_8571,N_8029);
or U9746 (N_9746,N_8354,N_8486);
nor U9747 (N_9747,N_8077,N_8204);
nand U9748 (N_9748,N_8949,N_8722);
or U9749 (N_9749,N_8585,N_8469);
or U9750 (N_9750,N_8641,N_8782);
nor U9751 (N_9751,N_8419,N_8084);
or U9752 (N_9752,N_8111,N_8949);
nand U9753 (N_9753,N_8566,N_8041);
nand U9754 (N_9754,N_8495,N_8660);
nor U9755 (N_9755,N_8618,N_8574);
or U9756 (N_9756,N_8440,N_8894);
nor U9757 (N_9757,N_8115,N_8772);
nand U9758 (N_9758,N_8702,N_8448);
or U9759 (N_9759,N_8130,N_8467);
or U9760 (N_9760,N_8931,N_8929);
or U9761 (N_9761,N_8284,N_8480);
nand U9762 (N_9762,N_8710,N_8404);
nand U9763 (N_9763,N_8897,N_8477);
nand U9764 (N_9764,N_8616,N_8771);
or U9765 (N_9765,N_8847,N_8564);
nor U9766 (N_9766,N_8400,N_8686);
and U9767 (N_9767,N_8890,N_8671);
and U9768 (N_9768,N_8846,N_8172);
or U9769 (N_9769,N_8688,N_8318);
and U9770 (N_9770,N_8841,N_8610);
nand U9771 (N_9771,N_8365,N_8600);
nand U9772 (N_9772,N_8941,N_8576);
or U9773 (N_9773,N_8405,N_8979);
or U9774 (N_9774,N_8751,N_8464);
nand U9775 (N_9775,N_8853,N_8102);
and U9776 (N_9776,N_8555,N_8803);
and U9777 (N_9777,N_8933,N_8048);
and U9778 (N_9778,N_8402,N_8971);
or U9779 (N_9779,N_8659,N_8062);
or U9780 (N_9780,N_8626,N_8960);
nand U9781 (N_9781,N_8114,N_8366);
nand U9782 (N_9782,N_8696,N_8183);
nand U9783 (N_9783,N_8449,N_8646);
nor U9784 (N_9784,N_8296,N_8558);
nand U9785 (N_9785,N_8376,N_8256);
nor U9786 (N_9786,N_8309,N_8227);
nor U9787 (N_9787,N_8764,N_8780);
and U9788 (N_9788,N_8549,N_8584);
or U9789 (N_9789,N_8172,N_8556);
nor U9790 (N_9790,N_8912,N_8669);
nor U9791 (N_9791,N_8414,N_8618);
and U9792 (N_9792,N_8314,N_8960);
and U9793 (N_9793,N_8449,N_8185);
or U9794 (N_9794,N_8132,N_8052);
and U9795 (N_9795,N_8668,N_8258);
nand U9796 (N_9796,N_8218,N_8290);
and U9797 (N_9797,N_8084,N_8746);
nand U9798 (N_9798,N_8595,N_8291);
nand U9799 (N_9799,N_8429,N_8617);
and U9800 (N_9800,N_8062,N_8788);
and U9801 (N_9801,N_8363,N_8148);
nor U9802 (N_9802,N_8756,N_8403);
or U9803 (N_9803,N_8202,N_8710);
and U9804 (N_9804,N_8468,N_8293);
and U9805 (N_9805,N_8062,N_8397);
and U9806 (N_9806,N_8896,N_8348);
nor U9807 (N_9807,N_8939,N_8961);
or U9808 (N_9808,N_8402,N_8895);
and U9809 (N_9809,N_8629,N_8083);
and U9810 (N_9810,N_8986,N_8438);
nand U9811 (N_9811,N_8745,N_8471);
and U9812 (N_9812,N_8573,N_8175);
or U9813 (N_9813,N_8961,N_8735);
nor U9814 (N_9814,N_8430,N_8565);
nor U9815 (N_9815,N_8100,N_8079);
nand U9816 (N_9816,N_8388,N_8539);
nor U9817 (N_9817,N_8603,N_8350);
or U9818 (N_9818,N_8283,N_8782);
nand U9819 (N_9819,N_8090,N_8783);
and U9820 (N_9820,N_8802,N_8405);
nand U9821 (N_9821,N_8204,N_8569);
or U9822 (N_9822,N_8991,N_8254);
or U9823 (N_9823,N_8577,N_8916);
nor U9824 (N_9824,N_8297,N_8897);
or U9825 (N_9825,N_8837,N_8152);
nand U9826 (N_9826,N_8140,N_8452);
nand U9827 (N_9827,N_8122,N_8694);
or U9828 (N_9828,N_8579,N_8233);
nor U9829 (N_9829,N_8671,N_8833);
and U9830 (N_9830,N_8889,N_8129);
and U9831 (N_9831,N_8260,N_8038);
or U9832 (N_9832,N_8378,N_8980);
or U9833 (N_9833,N_8743,N_8475);
and U9834 (N_9834,N_8901,N_8509);
nor U9835 (N_9835,N_8844,N_8096);
nor U9836 (N_9836,N_8721,N_8879);
or U9837 (N_9837,N_8563,N_8504);
and U9838 (N_9838,N_8675,N_8625);
and U9839 (N_9839,N_8767,N_8838);
and U9840 (N_9840,N_8213,N_8119);
nor U9841 (N_9841,N_8740,N_8219);
and U9842 (N_9842,N_8233,N_8889);
nand U9843 (N_9843,N_8594,N_8976);
nor U9844 (N_9844,N_8380,N_8952);
and U9845 (N_9845,N_8192,N_8779);
nand U9846 (N_9846,N_8122,N_8904);
and U9847 (N_9847,N_8145,N_8814);
or U9848 (N_9848,N_8574,N_8474);
nor U9849 (N_9849,N_8962,N_8803);
or U9850 (N_9850,N_8658,N_8172);
and U9851 (N_9851,N_8029,N_8085);
and U9852 (N_9852,N_8205,N_8554);
nand U9853 (N_9853,N_8835,N_8266);
or U9854 (N_9854,N_8873,N_8214);
or U9855 (N_9855,N_8374,N_8979);
and U9856 (N_9856,N_8831,N_8595);
nand U9857 (N_9857,N_8752,N_8312);
nor U9858 (N_9858,N_8361,N_8038);
nand U9859 (N_9859,N_8539,N_8719);
and U9860 (N_9860,N_8744,N_8508);
nand U9861 (N_9861,N_8448,N_8360);
nor U9862 (N_9862,N_8081,N_8784);
or U9863 (N_9863,N_8684,N_8713);
or U9864 (N_9864,N_8940,N_8853);
and U9865 (N_9865,N_8171,N_8813);
xnor U9866 (N_9866,N_8094,N_8084);
nor U9867 (N_9867,N_8792,N_8165);
or U9868 (N_9868,N_8394,N_8563);
or U9869 (N_9869,N_8184,N_8429);
and U9870 (N_9870,N_8789,N_8804);
nand U9871 (N_9871,N_8141,N_8043);
nand U9872 (N_9872,N_8564,N_8966);
and U9873 (N_9873,N_8787,N_8344);
or U9874 (N_9874,N_8321,N_8194);
and U9875 (N_9875,N_8488,N_8635);
nor U9876 (N_9876,N_8074,N_8389);
and U9877 (N_9877,N_8999,N_8567);
or U9878 (N_9878,N_8508,N_8963);
nand U9879 (N_9879,N_8022,N_8655);
nor U9880 (N_9880,N_8485,N_8309);
nand U9881 (N_9881,N_8516,N_8344);
nand U9882 (N_9882,N_8562,N_8563);
nor U9883 (N_9883,N_8719,N_8100);
nor U9884 (N_9884,N_8467,N_8656);
or U9885 (N_9885,N_8427,N_8309);
nand U9886 (N_9886,N_8527,N_8731);
xnor U9887 (N_9887,N_8467,N_8321);
nand U9888 (N_9888,N_8172,N_8093);
or U9889 (N_9889,N_8673,N_8254);
nand U9890 (N_9890,N_8683,N_8621);
nand U9891 (N_9891,N_8609,N_8287);
or U9892 (N_9892,N_8564,N_8664);
nor U9893 (N_9893,N_8710,N_8998);
nand U9894 (N_9894,N_8912,N_8477);
and U9895 (N_9895,N_8993,N_8457);
and U9896 (N_9896,N_8091,N_8723);
nand U9897 (N_9897,N_8248,N_8795);
and U9898 (N_9898,N_8279,N_8190);
or U9899 (N_9899,N_8271,N_8593);
nand U9900 (N_9900,N_8058,N_8280);
or U9901 (N_9901,N_8062,N_8719);
or U9902 (N_9902,N_8754,N_8050);
nor U9903 (N_9903,N_8525,N_8843);
or U9904 (N_9904,N_8071,N_8128);
nand U9905 (N_9905,N_8940,N_8673);
or U9906 (N_9906,N_8768,N_8686);
or U9907 (N_9907,N_8483,N_8017);
and U9908 (N_9908,N_8618,N_8395);
nand U9909 (N_9909,N_8293,N_8736);
and U9910 (N_9910,N_8500,N_8948);
or U9911 (N_9911,N_8842,N_8332);
and U9912 (N_9912,N_8469,N_8917);
and U9913 (N_9913,N_8675,N_8552);
or U9914 (N_9914,N_8024,N_8847);
and U9915 (N_9915,N_8007,N_8084);
or U9916 (N_9916,N_8754,N_8145);
or U9917 (N_9917,N_8100,N_8445);
nor U9918 (N_9918,N_8243,N_8222);
or U9919 (N_9919,N_8220,N_8108);
nand U9920 (N_9920,N_8108,N_8242);
and U9921 (N_9921,N_8420,N_8762);
nor U9922 (N_9922,N_8908,N_8622);
and U9923 (N_9923,N_8084,N_8936);
nor U9924 (N_9924,N_8179,N_8869);
nand U9925 (N_9925,N_8380,N_8018);
nor U9926 (N_9926,N_8302,N_8738);
nor U9927 (N_9927,N_8419,N_8781);
nor U9928 (N_9928,N_8875,N_8464);
or U9929 (N_9929,N_8156,N_8587);
or U9930 (N_9930,N_8164,N_8808);
nor U9931 (N_9931,N_8675,N_8269);
nor U9932 (N_9932,N_8006,N_8956);
xor U9933 (N_9933,N_8152,N_8338);
or U9934 (N_9934,N_8452,N_8085);
nor U9935 (N_9935,N_8162,N_8685);
nand U9936 (N_9936,N_8793,N_8207);
nor U9937 (N_9937,N_8230,N_8411);
and U9938 (N_9938,N_8794,N_8409);
nand U9939 (N_9939,N_8455,N_8367);
and U9940 (N_9940,N_8768,N_8944);
nand U9941 (N_9941,N_8022,N_8873);
and U9942 (N_9942,N_8704,N_8809);
nand U9943 (N_9943,N_8462,N_8838);
nor U9944 (N_9944,N_8710,N_8676);
nor U9945 (N_9945,N_8422,N_8519);
nand U9946 (N_9946,N_8165,N_8343);
nand U9947 (N_9947,N_8892,N_8154);
nor U9948 (N_9948,N_8767,N_8956);
and U9949 (N_9949,N_8094,N_8353);
or U9950 (N_9950,N_8983,N_8250);
nor U9951 (N_9951,N_8248,N_8755);
nor U9952 (N_9952,N_8836,N_8227);
nor U9953 (N_9953,N_8149,N_8549);
nor U9954 (N_9954,N_8585,N_8148);
and U9955 (N_9955,N_8929,N_8973);
and U9956 (N_9956,N_8416,N_8715);
nand U9957 (N_9957,N_8348,N_8168);
or U9958 (N_9958,N_8572,N_8177);
and U9959 (N_9959,N_8230,N_8611);
and U9960 (N_9960,N_8315,N_8894);
nand U9961 (N_9961,N_8754,N_8390);
nor U9962 (N_9962,N_8571,N_8915);
nor U9963 (N_9963,N_8953,N_8949);
nor U9964 (N_9964,N_8875,N_8737);
and U9965 (N_9965,N_8572,N_8776);
or U9966 (N_9966,N_8072,N_8210);
and U9967 (N_9967,N_8264,N_8511);
nor U9968 (N_9968,N_8756,N_8155);
and U9969 (N_9969,N_8186,N_8311);
or U9970 (N_9970,N_8424,N_8340);
nand U9971 (N_9971,N_8486,N_8084);
or U9972 (N_9972,N_8658,N_8488);
nor U9973 (N_9973,N_8013,N_8842);
nand U9974 (N_9974,N_8436,N_8671);
and U9975 (N_9975,N_8532,N_8649);
nor U9976 (N_9976,N_8252,N_8424);
and U9977 (N_9977,N_8413,N_8041);
nand U9978 (N_9978,N_8506,N_8012);
nor U9979 (N_9979,N_8872,N_8470);
or U9980 (N_9980,N_8218,N_8213);
nand U9981 (N_9981,N_8762,N_8304);
or U9982 (N_9982,N_8236,N_8559);
and U9983 (N_9983,N_8047,N_8152);
or U9984 (N_9984,N_8877,N_8407);
nand U9985 (N_9985,N_8296,N_8114);
or U9986 (N_9986,N_8804,N_8935);
or U9987 (N_9987,N_8721,N_8928);
nand U9988 (N_9988,N_8486,N_8439);
or U9989 (N_9989,N_8222,N_8773);
and U9990 (N_9990,N_8144,N_8711);
nor U9991 (N_9991,N_8589,N_8503);
nand U9992 (N_9992,N_8352,N_8007);
or U9993 (N_9993,N_8762,N_8725);
or U9994 (N_9994,N_8824,N_8346);
or U9995 (N_9995,N_8145,N_8094);
or U9996 (N_9996,N_8110,N_8493);
or U9997 (N_9997,N_8270,N_8803);
or U9998 (N_9998,N_8213,N_8235);
xnor U9999 (N_9999,N_8211,N_8655);
nor UO_0 (O_0,N_9056,N_9229);
nor UO_1 (O_1,N_9869,N_9738);
nand UO_2 (O_2,N_9401,N_9148);
or UO_3 (O_3,N_9486,N_9980);
nor UO_4 (O_4,N_9429,N_9447);
nor UO_5 (O_5,N_9457,N_9638);
nand UO_6 (O_6,N_9513,N_9078);
and UO_7 (O_7,N_9102,N_9350);
nand UO_8 (O_8,N_9245,N_9271);
nor UO_9 (O_9,N_9130,N_9297);
or UO_10 (O_10,N_9131,N_9410);
nor UO_11 (O_11,N_9799,N_9007);
nand UO_12 (O_12,N_9592,N_9988);
and UO_13 (O_13,N_9241,N_9963);
nand UO_14 (O_14,N_9335,N_9969);
and UO_15 (O_15,N_9087,N_9491);
nor UO_16 (O_16,N_9525,N_9284);
or UO_17 (O_17,N_9158,N_9202);
nor UO_18 (O_18,N_9762,N_9997);
nand UO_19 (O_19,N_9938,N_9309);
nand UO_20 (O_20,N_9181,N_9793);
or UO_21 (O_21,N_9450,N_9892);
or UO_22 (O_22,N_9016,N_9675);
and UO_23 (O_23,N_9701,N_9783);
nand UO_24 (O_24,N_9746,N_9755);
nor UO_25 (O_25,N_9665,N_9159);
or UO_26 (O_26,N_9975,N_9239);
or UO_27 (O_27,N_9461,N_9802);
nand UO_28 (O_28,N_9015,N_9797);
nand UO_29 (O_29,N_9246,N_9176);
and UO_30 (O_30,N_9786,N_9702);
or UO_31 (O_31,N_9994,N_9961);
and UO_32 (O_32,N_9707,N_9343);
xor UO_33 (O_33,N_9691,N_9101);
nand UO_34 (O_34,N_9222,N_9062);
or UO_35 (O_35,N_9020,N_9359);
and UO_36 (O_36,N_9921,N_9948);
or UO_37 (O_37,N_9185,N_9908);
or UO_38 (O_38,N_9647,N_9315);
or UO_39 (O_39,N_9937,N_9911);
and UO_40 (O_40,N_9737,N_9423);
or UO_41 (O_41,N_9837,N_9870);
nand UO_42 (O_42,N_9803,N_9372);
nand UO_43 (O_43,N_9956,N_9289);
or UO_44 (O_44,N_9273,N_9575);
nor UO_45 (O_45,N_9085,N_9337);
nand UO_46 (O_46,N_9281,N_9195);
nand UO_47 (O_47,N_9238,N_9287);
nand UO_48 (O_48,N_9864,N_9563);
nand UO_49 (O_49,N_9024,N_9778);
and UO_50 (O_50,N_9127,N_9221);
or UO_51 (O_51,N_9951,N_9192);
nor UO_52 (O_52,N_9568,N_9674);
or UO_53 (O_53,N_9259,N_9520);
and UO_54 (O_54,N_9144,N_9099);
or UO_55 (O_55,N_9001,N_9371);
and UO_56 (O_56,N_9818,N_9605);
nor UO_57 (O_57,N_9157,N_9698);
or UO_58 (O_58,N_9295,N_9889);
and UO_59 (O_59,N_9953,N_9950);
and UO_60 (O_60,N_9489,N_9827);
nor UO_61 (O_61,N_9266,N_9523);
and UO_62 (O_62,N_9111,N_9730);
nand UO_63 (O_63,N_9595,N_9881);
nor UO_64 (O_64,N_9077,N_9606);
or UO_65 (O_65,N_9143,N_9532);
nand UO_66 (O_66,N_9808,N_9692);
or UO_67 (O_67,N_9381,N_9645);
nand UO_68 (O_68,N_9634,N_9118);
or UO_69 (O_69,N_9231,N_9824);
nor UO_70 (O_70,N_9046,N_9557);
and UO_71 (O_71,N_9455,N_9546);
nand UO_72 (O_72,N_9188,N_9472);
and UO_73 (O_73,N_9353,N_9326);
xor UO_74 (O_74,N_9017,N_9213);
or UO_75 (O_75,N_9421,N_9871);
or UO_76 (O_76,N_9025,N_9739);
nand UO_77 (O_77,N_9415,N_9112);
nor UO_78 (O_78,N_9223,N_9706);
or UO_79 (O_79,N_9976,N_9654);
and UO_80 (O_80,N_9227,N_9646);
and UO_81 (O_81,N_9097,N_9957);
nor UO_82 (O_82,N_9933,N_9960);
or UO_83 (O_83,N_9280,N_9141);
nand UO_84 (O_84,N_9735,N_9392);
nand UO_85 (O_85,N_9906,N_9296);
and UO_86 (O_86,N_9795,N_9901);
or UO_87 (O_87,N_9219,N_9039);
and UO_88 (O_88,N_9140,N_9442);
nand UO_89 (O_89,N_9201,N_9791);
xnor UO_90 (O_90,N_9465,N_9368);
nor UO_91 (O_91,N_9715,N_9531);
and UO_92 (O_92,N_9059,N_9844);
or UO_93 (O_93,N_9731,N_9688);
and UO_94 (O_94,N_9362,N_9603);
and UO_95 (O_95,N_9828,N_9435);
or UO_96 (O_96,N_9409,N_9596);
nand UO_97 (O_97,N_9651,N_9612);
nand UO_98 (O_98,N_9434,N_9240);
and UO_99 (O_99,N_9011,N_9339);
nand UO_100 (O_100,N_9940,N_9218);
and UO_101 (O_101,N_9294,N_9175);
nand UO_102 (O_102,N_9466,N_9173);
or UO_103 (O_103,N_9153,N_9915);
and UO_104 (O_104,N_9913,N_9560);
xor UO_105 (O_105,N_9398,N_9801);
nand UO_106 (O_106,N_9866,N_9064);
or UO_107 (O_107,N_9449,N_9251);
and UO_108 (O_108,N_9577,N_9248);
and UO_109 (O_109,N_9189,N_9752);
nand UO_110 (O_110,N_9564,N_9652);
nand UO_111 (O_111,N_9865,N_9619);
or UO_112 (O_112,N_9321,N_9057);
nor UO_113 (O_113,N_9399,N_9905);
and UO_114 (O_114,N_9637,N_9724);
nand UO_115 (O_115,N_9781,N_9269);
or UO_116 (O_116,N_9314,N_9138);
nor UO_117 (O_117,N_9258,N_9813);
or UO_118 (O_118,N_9700,N_9829);
nand UO_119 (O_119,N_9225,N_9427);
or UO_120 (O_120,N_9740,N_9045);
nand UO_121 (O_121,N_9215,N_9501);
or UO_122 (O_122,N_9839,N_9726);
and UO_123 (O_123,N_9385,N_9649);
nand UO_124 (O_124,N_9894,N_9552);
nand UO_125 (O_125,N_9317,N_9877);
and UO_126 (O_126,N_9216,N_9556);
or UO_127 (O_127,N_9858,N_9172);
nand UO_128 (O_128,N_9260,N_9203);
and UO_129 (O_129,N_9842,N_9363);
or UO_130 (O_130,N_9884,N_9747);
and UO_131 (O_131,N_9500,N_9060);
nor UO_132 (O_132,N_9413,N_9763);
nand UO_133 (O_133,N_9150,N_9040);
and UO_134 (O_134,N_9787,N_9096);
or UO_135 (O_135,N_9920,N_9268);
nand UO_136 (O_136,N_9636,N_9806);
and UO_137 (O_137,N_9506,N_9947);
and UO_138 (O_138,N_9614,N_9855);
or UO_139 (O_139,N_9917,N_9609);
nand UO_140 (O_140,N_9772,N_9151);
or UO_141 (O_141,N_9643,N_9263);
or UO_142 (O_142,N_9689,N_9356);
and UO_143 (O_143,N_9162,N_9375);
nor UO_144 (O_144,N_9854,N_9374);
or UO_145 (O_145,N_9492,N_9623);
nor UO_146 (O_146,N_9699,N_9745);
or UO_147 (O_147,N_9305,N_9186);
and UO_148 (O_148,N_9760,N_9400);
nor UO_149 (O_149,N_9332,N_9931);
nand UO_150 (O_150,N_9285,N_9431);
and UO_151 (O_151,N_9872,N_9272);
nand UO_152 (O_152,N_9032,N_9822);
and UO_153 (O_153,N_9805,N_9416);
nor UO_154 (O_154,N_9704,N_9678);
and UO_155 (O_155,N_9562,N_9845);
or UO_156 (O_156,N_9515,N_9464);
nand UO_157 (O_157,N_9662,N_9926);
and UO_158 (O_158,N_9900,N_9946);
nor UO_159 (O_159,N_9279,N_9644);
and UO_160 (O_160,N_9544,N_9955);
nand UO_161 (O_161,N_9261,N_9528);
and UO_162 (O_162,N_9773,N_9211);
or UO_163 (O_163,N_9934,N_9511);
and UO_164 (O_164,N_9081,N_9054);
and UO_165 (O_165,N_9843,N_9384);
nor UO_166 (O_166,N_9110,N_9771);
or UO_167 (O_167,N_9481,N_9566);
nand UO_168 (O_168,N_9601,N_9454);
nand UO_169 (O_169,N_9168,N_9549);
and UO_170 (O_170,N_9657,N_9658);
nand UO_171 (O_171,N_9114,N_9659);
nor UO_172 (O_172,N_9536,N_9504);
and UO_173 (O_173,N_9846,N_9456);
and UO_174 (O_174,N_9696,N_9070);
nand UO_175 (O_175,N_9732,N_9517);
nand UO_176 (O_176,N_9952,N_9618);
or UO_177 (O_177,N_9256,N_9891);
nand UO_178 (O_178,N_9403,N_9578);
nor UO_179 (O_179,N_9918,N_9565);
nor UO_180 (O_180,N_9928,N_9503);
or UO_181 (O_181,N_9655,N_9323);
or UO_182 (O_182,N_9255,N_9460);
nand UO_183 (O_183,N_9545,N_9676);
or UO_184 (O_184,N_9823,N_9620);
and UO_185 (O_185,N_9290,N_9220);
nand UO_186 (O_186,N_9076,N_9518);
nor UO_187 (O_187,N_9572,N_9333);
nor UO_188 (O_188,N_9995,N_9320);
nor UO_189 (O_189,N_9812,N_9425);
and UO_190 (O_190,N_9733,N_9382);
and UO_191 (O_191,N_9448,N_9708);
or UO_192 (O_192,N_9792,N_9686);
or UO_193 (O_193,N_9370,N_9569);
xor UO_194 (O_194,N_9819,N_9117);
nand UO_195 (O_195,N_9169,N_9971);
nor UO_196 (O_196,N_9825,N_9932);
nor UO_197 (O_197,N_9554,N_9648);
nand UO_198 (O_198,N_9207,N_9710);
or UO_199 (O_199,N_9003,N_9499);
nand UO_200 (O_200,N_9301,N_9669);
nor UO_201 (O_201,N_9880,N_9196);
and UO_202 (O_202,N_9198,N_9452);
nor UO_203 (O_203,N_9814,N_9205);
or UO_204 (O_204,N_9217,N_9067);
nand UO_205 (O_205,N_9693,N_9182);
nor UO_206 (O_206,N_9018,N_9073);
and UO_207 (O_207,N_9847,N_9474);
nand UO_208 (O_208,N_9841,N_9958);
nand UO_209 (O_209,N_9863,N_9991);
or UO_210 (O_210,N_9179,N_9083);
nand UO_211 (O_211,N_9899,N_9929);
and UO_212 (O_212,N_9132,N_9754);
or UO_213 (O_213,N_9625,N_9613);
nor UO_214 (O_214,N_9538,N_9012);
nand UO_215 (O_215,N_9589,N_9071);
and UO_216 (O_216,N_9584,N_9631);
and UO_217 (O_217,N_9903,N_9981);
nand UO_218 (O_218,N_9809,N_9660);
or UO_219 (O_219,N_9488,N_9530);
nor UO_220 (O_220,N_9044,N_9681);
nor UO_221 (O_221,N_9909,N_9300);
or UO_222 (O_222,N_9264,N_9149);
nor UO_223 (O_223,N_9935,N_9789);
or UO_224 (O_224,N_9089,N_9622);
or UO_225 (O_225,N_9498,N_9019);
nor UO_226 (O_226,N_9318,N_9432);
or UO_227 (O_227,N_9079,N_9656);
nor UO_228 (O_228,N_9387,N_9088);
nor UO_229 (O_229,N_9850,N_9590);
or UO_230 (O_230,N_9887,N_9838);
and UO_231 (O_231,N_9687,N_9364);
or UO_232 (O_232,N_9242,N_9109);
nor UO_233 (O_233,N_9862,N_9133);
and UO_234 (O_234,N_9344,N_9650);
or UO_235 (O_235,N_9581,N_9237);
or UO_236 (O_236,N_9537,N_9848);
nand UO_237 (O_237,N_9360,N_9567);
nand UO_238 (O_238,N_9286,N_9541);
or UO_239 (O_239,N_9445,N_9526);
and UO_240 (O_240,N_9758,N_9635);
nand UO_241 (O_241,N_9725,N_9288);
and UO_242 (O_242,N_9598,N_9204);
or UO_243 (O_243,N_9741,N_9191);
or UO_244 (O_244,N_9502,N_9723);
and UO_245 (O_245,N_9630,N_9766);
nand UO_246 (O_246,N_9058,N_9555);
nor UO_247 (O_247,N_9734,N_9036);
nor UO_248 (O_248,N_9306,N_9916);
or UO_249 (O_249,N_9853,N_9482);
xnor UO_250 (O_250,N_9031,N_9411);
nand UO_251 (O_251,N_9230,N_9769);
or UO_252 (O_252,N_9234,N_9208);
nand UO_253 (O_253,N_9756,N_9507);
and UO_254 (O_254,N_9800,N_9604);
nand UO_255 (O_255,N_9147,N_9840);
nor UO_256 (O_256,N_9104,N_9583);
or UO_257 (O_257,N_9042,N_9653);
and UO_258 (O_258,N_9142,N_9856);
nor UO_259 (O_259,N_9100,N_9422);
nor UO_260 (O_260,N_9119,N_9599);
or UO_261 (O_261,N_9341,N_9436);
or UO_262 (O_262,N_9558,N_9441);
or UO_263 (O_263,N_9121,N_9875);
and UO_264 (O_264,N_9551,N_9668);
nand UO_265 (O_265,N_9402,N_9395);
nand UO_266 (O_266,N_9386,N_9868);
nor UO_267 (O_267,N_9171,N_9535);
nand UO_268 (O_268,N_9270,N_9559);
or UO_269 (O_269,N_9051,N_9600);
nor UO_270 (O_270,N_9125,N_9721);
nor UO_271 (O_271,N_9209,N_9084);
nand UO_272 (O_272,N_9233,N_9005);
nand UO_273 (O_273,N_9593,N_9210);
nand UO_274 (O_274,N_9468,N_9890);
and UO_275 (O_275,N_9508,N_9826);
and UO_276 (O_276,N_9964,N_9327);
or UO_277 (O_277,N_9907,N_9165);
or UO_278 (O_278,N_9419,N_9770);
or UO_279 (O_279,N_9945,N_9462);
and UO_280 (O_280,N_9529,N_9072);
nand UO_281 (O_281,N_9357,N_9383);
or UO_282 (O_282,N_9106,N_9055);
or UO_283 (O_283,N_9896,N_9002);
nor UO_284 (O_284,N_9155,N_9053);
and UO_285 (O_285,N_9103,N_9594);
or UO_286 (O_286,N_9912,N_9094);
and UO_287 (O_287,N_9616,N_9459);
or UO_288 (O_288,N_9524,N_9553);
nor UO_289 (O_289,N_9744,N_9408);
xnor UO_290 (O_290,N_9876,N_9033);
or UO_291 (O_291,N_9407,N_9883);
nand UO_292 (O_292,N_9428,N_9671);
or UO_293 (O_293,N_9048,N_9161);
and UO_294 (O_294,N_9663,N_9322);
and UO_295 (O_295,N_9919,N_9576);
and UO_296 (O_296,N_9331,N_9999);
nand UO_297 (O_297,N_9722,N_9831);
nand UO_298 (O_298,N_9080,N_9063);
nor UO_299 (O_299,N_9780,N_9610);
and UO_300 (O_300,N_9135,N_9629);
and UO_301 (O_301,N_9750,N_9910);
nand UO_302 (O_302,N_9214,N_9939);
nand UO_303 (O_303,N_9369,N_9661);
nor UO_304 (O_304,N_9519,N_9404);
or UO_305 (O_305,N_9683,N_9206);
or UO_306 (O_306,N_9979,N_9299);
and UO_307 (O_307,N_9376,N_9340);
and UO_308 (O_308,N_9712,N_9521);
nor UO_309 (O_309,N_9685,N_9949);
or UO_310 (O_310,N_9505,N_9128);
or UO_311 (O_311,N_9550,N_9160);
or UO_312 (O_312,N_9393,N_9120);
or UO_313 (O_313,N_9304,N_9542);
or UO_314 (O_314,N_9561,N_9471);
nor UO_315 (O_315,N_9418,N_9930);
or UO_316 (O_316,N_9137,N_9467);
nand UO_317 (O_317,N_9742,N_9998);
nor UO_318 (O_318,N_9989,N_9509);
and UO_319 (O_319,N_9815,N_9004);
xor UO_320 (O_320,N_9882,N_9310);
nand UO_321 (O_321,N_9052,N_9439);
nand UO_322 (O_322,N_9212,N_9113);
and UO_323 (O_323,N_9720,N_9859);
nand UO_324 (O_324,N_9897,N_9366);
nor UO_325 (O_325,N_9275,N_9389);
nand UO_326 (O_326,N_9817,N_9904);
nor UO_327 (O_327,N_9420,N_9570);
or UO_328 (O_328,N_9463,N_9035);
nand UO_329 (O_329,N_9718,N_9777);
nor UO_330 (O_330,N_9785,N_9338);
nor UO_331 (O_331,N_9412,N_9954);
nand UO_332 (O_332,N_9167,N_9727);
nor UO_333 (O_333,N_9832,N_9573);
and UO_334 (O_334,N_9095,N_9197);
or UO_335 (O_335,N_9252,N_9247);
and UO_336 (O_336,N_9249,N_9968);
nand UO_337 (O_337,N_9962,N_9522);
and UO_338 (O_338,N_9487,N_9367);
nor UO_339 (O_339,N_9354,N_9586);
nand UO_340 (O_340,N_9199,N_9302);
or UO_341 (O_341,N_9276,N_9378);
nand UO_342 (O_342,N_9074,N_9713);
and UO_343 (O_343,N_9090,N_9782);
and UO_344 (O_344,N_9026,N_9834);
nand UO_345 (O_345,N_9621,N_9765);
and UO_346 (O_346,N_9512,N_9878);
nor UO_347 (O_347,N_9022,N_9451);
or UO_348 (O_348,N_9679,N_9667);
and UO_349 (O_349,N_9334,N_9107);
nand UO_350 (O_350,N_9123,N_9974);
nand UO_351 (O_351,N_9642,N_9611);
nor UO_352 (O_352,N_9682,N_9146);
and UO_353 (O_353,N_9193,N_9602);
and UO_354 (O_354,N_9226,N_9034);
nand UO_355 (O_355,N_9177,N_9029);
nand UO_356 (O_356,N_9821,N_9027);
nand UO_357 (O_357,N_9547,N_9888);
and UO_358 (O_358,N_9835,N_9478);
and UO_359 (O_359,N_9497,N_9494);
nand UO_360 (O_360,N_9579,N_9068);
and UO_361 (O_361,N_9010,N_9986);
and UO_362 (O_362,N_9440,N_9849);
nand UO_363 (O_363,N_9666,N_9925);
or UO_364 (O_364,N_9993,N_9485);
or UO_365 (O_365,N_9830,N_9810);
nor UO_366 (O_366,N_9358,N_9942);
or UO_367 (O_367,N_9607,N_9365);
and UO_368 (O_368,N_9743,N_9043);
or UO_369 (O_369,N_9493,N_9548);
nand UO_370 (O_370,N_9328,N_9154);
or UO_371 (O_371,N_9041,N_9761);
nor UO_372 (O_372,N_9970,N_9139);
or UO_373 (O_373,N_9458,N_9394);
nor UO_374 (O_374,N_9639,N_9291);
and UO_375 (O_375,N_9807,N_9977);
xor UO_376 (O_376,N_9278,N_9923);
nor UO_377 (O_377,N_9927,N_9187);
or UO_378 (O_378,N_9990,N_9673);
nand UO_379 (O_379,N_9779,N_9776);
xor UO_380 (O_380,N_9316,N_9379);
nand UO_381 (O_381,N_9775,N_9265);
nand UO_382 (O_382,N_9388,N_9174);
or UO_383 (O_383,N_9943,N_9967);
and UO_384 (O_384,N_9470,N_9075);
and UO_385 (O_385,N_9250,N_9093);
nor UO_386 (O_386,N_9361,N_9628);
or UO_387 (O_387,N_9262,N_9941);
and UO_388 (O_388,N_9082,N_9617);
nand UO_389 (O_389,N_9574,N_9684);
nand UO_390 (O_390,N_9116,N_9764);
nor UO_391 (O_391,N_9000,N_9200);
nand UO_392 (O_392,N_9597,N_9345);
nor UO_393 (O_393,N_9030,N_9023);
nand UO_394 (O_394,N_9728,N_9228);
or UO_395 (O_395,N_9352,N_9473);
or UO_396 (O_396,N_9061,N_9978);
nand UO_397 (O_397,N_9640,N_9914);
nor UO_398 (O_398,N_9895,N_9426);
nor UO_399 (O_399,N_9163,N_9527);
nor UO_400 (O_400,N_9373,N_9588);
nor UO_401 (O_401,N_9697,N_9820);
and UO_402 (O_402,N_9008,N_9983);
and UO_403 (O_403,N_9253,N_9633);
nand UO_404 (O_404,N_9312,N_9736);
and UO_405 (O_405,N_9982,N_9798);
nor UO_406 (O_406,N_9816,N_9936);
nand UO_407 (O_407,N_9047,N_9292);
or UO_408 (O_408,N_9719,N_9924);
nand UO_409 (O_409,N_9893,N_9351);
nor UO_410 (O_410,N_9711,N_9748);
and UO_411 (O_411,N_9484,N_9313);
and UO_412 (O_412,N_9224,N_9283);
or UO_413 (O_413,N_9277,N_9009);
nor UO_414 (O_414,N_9319,N_9757);
nand UO_415 (O_415,N_9444,N_9126);
nand UO_416 (O_416,N_9170,N_9184);
nand UO_417 (O_417,N_9886,N_9066);
and UO_418 (O_418,N_9804,N_9811);
or UO_419 (O_419,N_9615,N_9790);
and UO_420 (O_420,N_9703,N_9180);
nor UO_421 (O_421,N_9324,N_9129);
nand UO_422 (O_422,N_9479,N_9329);
nand UO_423 (O_423,N_9580,N_9396);
and UO_424 (O_424,N_9627,N_9380);
or UO_425 (O_425,N_9759,N_9244);
nor UO_426 (O_426,N_9134,N_9751);
nor UO_427 (O_427,N_9086,N_9694);
nand UO_428 (O_428,N_9695,N_9879);
nor UO_429 (O_429,N_9680,N_9985);
and UO_430 (O_430,N_9774,N_9236);
or UO_431 (O_431,N_9543,N_9833);
and UO_432 (O_432,N_9414,N_9232);
nand UO_433 (O_433,N_9050,N_9235);
nand UO_434 (O_434,N_9965,N_9514);
nand UO_435 (O_435,N_9105,N_9788);
nor UO_436 (O_436,N_9496,N_9349);
or UO_437 (O_437,N_9677,N_9307);
nand UO_438 (O_438,N_9347,N_9857);
nand UO_439 (O_439,N_9902,N_9705);
nor UO_440 (O_440,N_9124,N_9495);
nand UO_441 (O_441,N_9443,N_9267);
or UO_442 (O_442,N_9664,N_9984);
or UO_443 (O_443,N_9406,N_9405);
nand UO_444 (O_444,N_9014,N_9303);
nand UO_445 (O_445,N_9959,N_9476);
or UO_446 (O_446,N_9377,N_9115);
or UO_447 (O_447,N_9626,N_9641);
nor UO_448 (O_448,N_9298,N_9717);
nand UO_449 (O_449,N_9391,N_9397);
nand UO_450 (O_450,N_9156,N_9308);
nor UO_451 (O_451,N_9346,N_9768);
and UO_452 (O_452,N_9475,N_9417);
and UO_453 (O_453,N_9145,N_9274);
or UO_454 (O_454,N_9898,N_9992);
and UO_455 (O_455,N_9867,N_9178);
and UO_456 (O_456,N_9293,N_9885);
and UO_457 (O_457,N_9021,N_9477);
nand UO_458 (O_458,N_9582,N_9571);
and UO_459 (O_459,N_9510,N_9430);
nor UO_460 (O_460,N_9852,N_9091);
nand UO_461 (O_461,N_9183,N_9972);
and UO_462 (O_462,N_9098,N_9330);
and UO_463 (O_463,N_9092,N_9446);
nor UO_464 (O_464,N_9608,N_9767);
and UO_465 (O_465,N_9716,N_9714);
or UO_466 (O_466,N_9585,N_9516);
nand UO_467 (O_467,N_9006,N_9973);
or UO_468 (O_468,N_9670,N_9996);
nand UO_469 (O_469,N_9028,N_9672);
nor UO_470 (O_470,N_9194,N_9860);
nor UO_471 (O_471,N_9257,N_9038);
nand UO_472 (O_472,N_9049,N_9152);
nor UO_473 (O_473,N_9690,N_9749);
and UO_474 (O_474,N_9490,N_9874);
nor UO_475 (O_475,N_9437,N_9311);
nor UO_476 (O_476,N_9013,N_9166);
and UO_477 (O_477,N_9390,N_9944);
and UO_478 (O_478,N_9122,N_9453);
and UO_479 (O_479,N_9784,N_9729);
nor UO_480 (O_480,N_9108,N_9438);
nor UO_481 (O_481,N_9483,N_9480);
nor UO_482 (O_482,N_9851,N_9433);
nor UO_483 (O_483,N_9587,N_9190);
nor UO_484 (O_484,N_9540,N_9533);
and UO_485 (O_485,N_9796,N_9861);
nor UO_486 (O_486,N_9709,N_9534);
and UO_487 (O_487,N_9243,N_9065);
nand UO_488 (O_488,N_9922,N_9632);
or UO_489 (O_489,N_9069,N_9469);
nor UO_490 (O_490,N_9282,N_9794);
nand UO_491 (O_491,N_9355,N_9539);
or UO_492 (O_492,N_9336,N_9254);
nand UO_493 (O_493,N_9164,N_9037);
or UO_494 (O_494,N_9987,N_9325);
and UO_495 (O_495,N_9348,N_9342);
and UO_496 (O_496,N_9836,N_9591);
or UO_497 (O_497,N_9966,N_9424);
and UO_498 (O_498,N_9624,N_9753);
nand UO_499 (O_499,N_9873,N_9136);
nor UO_500 (O_500,N_9163,N_9974);
nor UO_501 (O_501,N_9955,N_9670);
or UO_502 (O_502,N_9644,N_9544);
or UO_503 (O_503,N_9696,N_9755);
or UO_504 (O_504,N_9920,N_9369);
nor UO_505 (O_505,N_9891,N_9536);
nand UO_506 (O_506,N_9491,N_9357);
nor UO_507 (O_507,N_9145,N_9697);
nor UO_508 (O_508,N_9498,N_9998);
or UO_509 (O_509,N_9195,N_9754);
nor UO_510 (O_510,N_9893,N_9223);
nand UO_511 (O_511,N_9607,N_9804);
or UO_512 (O_512,N_9383,N_9496);
nor UO_513 (O_513,N_9809,N_9194);
nor UO_514 (O_514,N_9718,N_9412);
or UO_515 (O_515,N_9483,N_9672);
and UO_516 (O_516,N_9887,N_9538);
and UO_517 (O_517,N_9466,N_9410);
or UO_518 (O_518,N_9535,N_9359);
and UO_519 (O_519,N_9019,N_9386);
nand UO_520 (O_520,N_9248,N_9763);
nor UO_521 (O_521,N_9039,N_9255);
nand UO_522 (O_522,N_9470,N_9115);
or UO_523 (O_523,N_9501,N_9195);
or UO_524 (O_524,N_9470,N_9589);
nor UO_525 (O_525,N_9207,N_9995);
and UO_526 (O_526,N_9493,N_9242);
nand UO_527 (O_527,N_9747,N_9827);
or UO_528 (O_528,N_9146,N_9773);
or UO_529 (O_529,N_9854,N_9582);
and UO_530 (O_530,N_9059,N_9968);
and UO_531 (O_531,N_9381,N_9158);
and UO_532 (O_532,N_9329,N_9091);
nand UO_533 (O_533,N_9716,N_9291);
or UO_534 (O_534,N_9635,N_9023);
and UO_535 (O_535,N_9214,N_9434);
nor UO_536 (O_536,N_9223,N_9196);
nand UO_537 (O_537,N_9947,N_9468);
or UO_538 (O_538,N_9806,N_9975);
nand UO_539 (O_539,N_9075,N_9594);
nand UO_540 (O_540,N_9220,N_9760);
or UO_541 (O_541,N_9349,N_9631);
or UO_542 (O_542,N_9908,N_9694);
nand UO_543 (O_543,N_9955,N_9782);
and UO_544 (O_544,N_9221,N_9826);
nand UO_545 (O_545,N_9708,N_9359);
and UO_546 (O_546,N_9152,N_9975);
or UO_547 (O_547,N_9966,N_9388);
or UO_548 (O_548,N_9447,N_9069);
nand UO_549 (O_549,N_9377,N_9884);
or UO_550 (O_550,N_9632,N_9054);
and UO_551 (O_551,N_9185,N_9620);
nor UO_552 (O_552,N_9094,N_9636);
nand UO_553 (O_553,N_9352,N_9249);
and UO_554 (O_554,N_9891,N_9551);
or UO_555 (O_555,N_9704,N_9883);
nor UO_556 (O_556,N_9939,N_9900);
or UO_557 (O_557,N_9889,N_9121);
and UO_558 (O_558,N_9342,N_9534);
nand UO_559 (O_559,N_9754,N_9079);
nand UO_560 (O_560,N_9611,N_9415);
nor UO_561 (O_561,N_9351,N_9842);
or UO_562 (O_562,N_9808,N_9689);
or UO_563 (O_563,N_9455,N_9805);
and UO_564 (O_564,N_9440,N_9579);
or UO_565 (O_565,N_9534,N_9391);
xor UO_566 (O_566,N_9406,N_9323);
nor UO_567 (O_567,N_9732,N_9349);
nor UO_568 (O_568,N_9847,N_9119);
nand UO_569 (O_569,N_9636,N_9277);
nor UO_570 (O_570,N_9875,N_9625);
or UO_571 (O_571,N_9899,N_9391);
nor UO_572 (O_572,N_9957,N_9131);
nand UO_573 (O_573,N_9917,N_9569);
or UO_574 (O_574,N_9175,N_9837);
nor UO_575 (O_575,N_9303,N_9225);
and UO_576 (O_576,N_9172,N_9728);
nor UO_577 (O_577,N_9022,N_9741);
or UO_578 (O_578,N_9893,N_9182);
and UO_579 (O_579,N_9980,N_9178);
nand UO_580 (O_580,N_9426,N_9334);
nand UO_581 (O_581,N_9415,N_9637);
nand UO_582 (O_582,N_9109,N_9222);
nor UO_583 (O_583,N_9319,N_9560);
nand UO_584 (O_584,N_9540,N_9664);
nor UO_585 (O_585,N_9053,N_9507);
nand UO_586 (O_586,N_9718,N_9955);
and UO_587 (O_587,N_9372,N_9183);
and UO_588 (O_588,N_9221,N_9474);
or UO_589 (O_589,N_9608,N_9606);
and UO_590 (O_590,N_9899,N_9230);
and UO_591 (O_591,N_9843,N_9202);
nand UO_592 (O_592,N_9885,N_9758);
nand UO_593 (O_593,N_9293,N_9433);
or UO_594 (O_594,N_9902,N_9229);
nor UO_595 (O_595,N_9463,N_9661);
nor UO_596 (O_596,N_9468,N_9712);
and UO_597 (O_597,N_9624,N_9315);
or UO_598 (O_598,N_9192,N_9408);
nand UO_599 (O_599,N_9394,N_9190);
or UO_600 (O_600,N_9873,N_9861);
nor UO_601 (O_601,N_9627,N_9126);
and UO_602 (O_602,N_9369,N_9933);
and UO_603 (O_603,N_9932,N_9495);
or UO_604 (O_604,N_9457,N_9853);
and UO_605 (O_605,N_9348,N_9914);
nor UO_606 (O_606,N_9846,N_9861);
nor UO_607 (O_607,N_9209,N_9749);
nor UO_608 (O_608,N_9878,N_9346);
nor UO_609 (O_609,N_9157,N_9303);
nand UO_610 (O_610,N_9899,N_9002);
nor UO_611 (O_611,N_9098,N_9540);
nand UO_612 (O_612,N_9733,N_9738);
nor UO_613 (O_613,N_9282,N_9174);
or UO_614 (O_614,N_9873,N_9767);
or UO_615 (O_615,N_9916,N_9508);
nor UO_616 (O_616,N_9133,N_9003);
nor UO_617 (O_617,N_9621,N_9365);
or UO_618 (O_618,N_9619,N_9838);
and UO_619 (O_619,N_9262,N_9646);
and UO_620 (O_620,N_9086,N_9430);
nor UO_621 (O_621,N_9276,N_9302);
nand UO_622 (O_622,N_9620,N_9994);
and UO_623 (O_623,N_9155,N_9274);
or UO_624 (O_624,N_9684,N_9094);
or UO_625 (O_625,N_9389,N_9426);
or UO_626 (O_626,N_9811,N_9897);
nand UO_627 (O_627,N_9148,N_9992);
and UO_628 (O_628,N_9963,N_9440);
or UO_629 (O_629,N_9556,N_9454);
xor UO_630 (O_630,N_9797,N_9207);
and UO_631 (O_631,N_9643,N_9099);
nor UO_632 (O_632,N_9019,N_9655);
nor UO_633 (O_633,N_9274,N_9353);
nand UO_634 (O_634,N_9593,N_9170);
nand UO_635 (O_635,N_9911,N_9026);
or UO_636 (O_636,N_9783,N_9985);
and UO_637 (O_637,N_9807,N_9287);
nor UO_638 (O_638,N_9551,N_9600);
nand UO_639 (O_639,N_9210,N_9710);
and UO_640 (O_640,N_9152,N_9488);
and UO_641 (O_641,N_9309,N_9871);
or UO_642 (O_642,N_9137,N_9901);
or UO_643 (O_643,N_9882,N_9873);
or UO_644 (O_644,N_9707,N_9406);
or UO_645 (O_645,N_9159,N_9329);
or UO_646 (O_646,N_9653,N_9595);
or UO_647 (O_647,N_9936,N_9266);
nor UO_648 (O_648,N_9625,N_9240);
nand UO_649 (O_649,N_9342,N_9502);
or UO_650 (O_650,N_9394,N_9843);
nand UO_651 (O_651,N_9027,N_9819);
nor UO_652 (O_652,N_9649,N_9359);
nor UO_653 (O_653,N_9945,N_9285);
nor UO_654 (O_654,N_9369,N_9352);
nand UO_655 (O_655,N_9418,N_9859);
nor UO_656 (O_656,N_9588,N_9099);
and UO_657 (O_657,N_9313,N_9327);
nor UO_658 (O_658,N_9747,N_9924);
nand UO_659 (O_659,N_9290,N_9674);
nand UO_660 (O_660,N_9259,N_9438);
nor UO_661 (O_661,N_9268,N_9445);
xnor UO_662 (O_662,N_9306,N_9907);
nand UO_663 (O_663,N_9509,N_9582);
or UO_664 (O_664,N_9467,N_9812);
nor UO_665 (O_665,N_9697,N_9828);
nand UO_666 (O_666,N_9521,N_9210);
nor UO_667 (O_667,N_9498,N_9301);
nor UO_668 (O_668,N_9575,N_9669);
or UO_669 (O_669,N_9567,N_9475);
nor UO_670 (O_670,N_9441,N_9762);
or UO_671 (O_671,N_9264,N_9609);
and UO_672 (O_672,N_9386,N_9524);
and UO_673 (O_673,N_9550,N_9674);
or UO_674 (O_674,N_9309,N_9168);
nor UO_675 (O_675,N_9477,N_9009);
nor UO_676 (O_676,N_9368,N_9914);
and UO_677 (O_677,N_9730,N_9698);
or UO_678 (O_678,N_9985,N_9099);
and UO_679 (O_679,N_9235,N_9686);
or UO_680 (O_680,N_9897,N_9207);
and UO_681 (O_681,N_9062,N_9177);
nor UO_682 (O_682,N_9431,N_9281);
or UO_683 (O_683,N_9348,N_9164);
nor UO_684 (O_684,N_9255,N_9268);
and UO_685 (O_685,N_9161,N_9968);
nor UO_686 (O_686,N_9060,N_9553);
or UO_687 (O_687,N_9286,N_9940);
nor UO_688 (O_688,N_9524,N_9319);
xor UO_689 (O_689,N_9146,N_9590);
nor UO_690 (O_690,N_9628,N_9050);
nand UO_691 (O_691,N_9371,N_9953);
nand UO_692 (O_692,N_9933,N_9717);
nand UO_693 (O_693,N_9985,N_9915);
nand UO_694 (O_694,N_9164,N_9825);
or UO_695 (O_695,N_9141,N_9305);
and UO_696 (O_696,N_9495,N_9694);
or UO_697 (O_697,N_9023,N_9799);
or UO_698 (O_698,N_9277,N_9629);
or UO_699 (O_699,N_9906,N_9449);
xor UO_700 (O_700,N_9291,N_9723);
nand UO_701 (O_701,N_9333,N_9164);
and UO_702 (O_702,N_9415,N_9412);
or UO_703 (O_703,N_9833,N_9283);
or UO_704 (O_704,N_9639,N_9212);
nand UO_705 (O_705,N_9619,N_9330);
nor UO_706 (O_706,N_9860,N_9936);
nand UO_707 (O_707,N_9457,N_9554);
nand UO_708 (O_708,N_9445,N_9239);
and UO_709 (O_709,N_9461,N_9495);
or UO_710 (O_710,N_9028,N_9886);
nand UO_711 (O_711,N_9414,N_9763);
nand UO_712 (O_712,N_9289,N_9181);
nand UO_713 (O_713,N_9618,N_9669);
nor UO_714 (O_714,N_9892,N_9607);
nor UO_715 (O_715,N_9626,N_9746);
nor UO_716 (O_716,N_9216,N_9043);
nand UO_717 (O_717,N_9272,N_9666);
nor UO_718 (O_718,N_9796,N_9716);
nand UO_719 (O_719,N_9562,N_9616);
nand UO_720 (O_720,N_9130,N_9870);
nand UO_721 (O_721,N_9700,N_9392);
or UO_722 (O_722,N_9794,N_9291);
nand UO_723 (O_723,N_9648,N_9827);
or UO_724 (O_724,N_9832,N_9148);
nor UO_725 (O_725,N_9860,N_9176);
and UO_726 (O_726,N_9408,N_9476);
nand UO_727 (O_727,N_9114,N_9819);
nor UO_728 (O_728,N_9722,N_9077);
nand UO_729 (O_729,N_9143,N_9513);
or UO_730 (O_730,N_9514,N_9085);
nor UO_731 (O_731,N_9433,N_9290);
and UO_732 (O_732,N_9393,N_9762);
and UO_733 (O_733,N_9763,N_9502);
nor UO_734 (O_734,N_9551,N_9220);
nor UO_735 (O_735,N_9613,N_9063);
or UO_736 (O_736,N_9774,N_9964);
or UO_737 (O_737,N_9259,N_9572);
nand UO_738 (O_738,N_9984,N_9012);
nor UO_739 (O_739,N_9788,N_9862);
nand UO_740 (O_740,N_9317,N_9024);
and UO_741 (O_741,N_9807,N_9069);
nand UO_742 (O_742,N_9956,N_9846);
nor UO_743 (O_743,N_9692,N_9242);
nand UO_744 (O_744,N_9144,N_9362);
nand UO_745 (O_745,N_9372,N_9234);
nand UO_746 (O_746,N_9720,N_9834);
nand UO_747 (O_747,N_9347,N_9513);
and UO_748 (O_748,N_9150,N_9472);
xnor UO_749 (O_749,N_9375,N_9376);
and UO_750 (O_750,N_9472,N_9912);
or UO_751 (O_751,N_9530,N_9649);
nand UO_752 (O_752,N_9980,N_9807);
and UO_753 (O_753,N_9893,N_9834);
or UO_754 (O_754,N_9284,N_9873);
nor UO_755 (O_755,N_9929,N_9885);
nor UO_756 (O_756,N_9002,N_9720);
or UO_757 (O_757,N_9575,N_9362);
and UO_758 (O_758,N_9401,N_9714);
nand UO_759 (O_759,N_9751,N_9532);
and UO_760 (O_760,N_9928,N_9474);
or UO_761 (O_761,N_9278,N_9379);
and UO_762 (O_762,N_9397,N_9327);
nand UO_763 (O_763,N_9944,N_9799);
or UO_764 (O_764,N_9481,N_9134);
nor UO_765 (O_765,N_9208,N_9217);
or UO_766 (O_766,N_9017,N_9915);
nor UO_767 (O_767,N_9908,N_9884);
nand UO_768 (O_768,N_9266,N_9814);
nand UO_769 (O_769,N_9550,N_9492);
and UO_770 (O_770,N_9840,N_9689);
or UO_771 (O_771,N_9264,N_9401);
and UO_772 (O_772,N_9117,N_9984);
nor UO_773 (O_773,N_9682,N_9139);
or UO_774 (O_774,N_9073,N_9786);
or UO_775 (O_775,N_9434,N_9128);
and UO_776 (O_776,N_9568,N_9706);
nand UO_777 (O_777,N_9999,N_9707);
nand UO_778 (O_778,N_9979,N_9911);
and UO_779 (O_779,N_9490,N_9557);
and UO_780 (O_780,N_9054,N_9408);
nand UO_781 (O_781,N_9835,N_9263);
and UO_782 (O_782,N_9400,N_9348);
nor UO_783 (O_783,N_9931,N_9284);
nor UO_784 (O_784,N_9879,N_9779);
nand UO_785 (O_785,N_9345,N_9587);
and UO_786 (O_786,N_9357,N_9813);
or UO_787 (O_787,N_9668,N_9495);
and UO_788 (O_788,N_9519,N_9021);
or UO_789 (O_789,N_9794,N_9491);
and UO_790 (O_790,N_9865,N_9572);
and UO_791 (O_791,N_9634,N_9268);
and UO_792 (O_792,N_9760,N_9858);
and UO_793 (O_793,N_9524,N_9348);
nand UO_794 (O_794,N_9337,N_9208);
nand UO_795 (O_795,N_9624,N_9658);
or UO_796 (O_796,N_9564,N_9094);
nand UO_797 (O_797,N_9173,N_9270);
and UO_798 (O_798,N_9467,N_9547);
nor UO_799 (O_799,N_9477,N_9090);
nand UO_800 (O_800,N_9394,N_9870);
nor UO_801 (O_801,N_9171,N_9480);
nor UO_802 (O_802,N_9146,N_9884);
nor UO_803 (O_803,N_9693,N_9828);
nand UO_804 (O_804,N_9768,N_9243);
nor UO_805 (O_805,N_9330,N_9747);
nor UO_806 (O_806,N_9439,N_9923);
or UO_807 (O_807,N_9027,N_9092);
nor UO_808 (O_808,N_9491,N_9095);
nor UO_809 (O_809,N_9387,N_9787);
or UO_810 (O_810,N_9312,N_9835);
or UO_811 (O_811,N_9980,N_9498);
and UO_812 (O_812,N_9246,N_9831);
nor UO_813 (O_813,N_9744,N_9496);
nand UO_814 (O_814,N_9360,N_9817);
and UO_815 (O_815,N_9175,N_9961);
nor UO_816 (O_816,N_9285,N_9559);
nor UO_817 (O_817,N_9626,N_9839);
or UO_818 (O_818,N_9122,N_9092);
nor UO_819 (O_819,N_9577,N_9553);
nand UO_820 (O_820,N_9818,N_9749);
and UO_821 (O_821,N_9559,N_9737);
and UO_822 (O_822,N_9729,N_9477);
nand UO_823 (O_823,N_9031,N_9135);
nor UO_824 (O_824,N_9266,N_9612);
nor UO_825 (O_825,N_9036,N_9051);
nand UO_826 (O_826,N_9895,N_9893);
or UO_827 (O_827,N_9721,N_9980);
nor UO_828 (O_828,N_9998,N_9878);
or UO_829 (O_829,N_9642,N_9783);
nand UO_830 (O_830,N_9414,N_9323);
nor UO_831 (O_831,N_9532,N_9734);
and UO_832 (O_832,N_9474,N_9037);
and UO_833 (O_833,N_9963,N_9314);
nand UO_834 (O_834,N_9980,N_9217);
and UO_835 (O_835,N_9905,N_9394);
or UO_836 (O_836,N_9961,N_9026);
and UO_837 (O_837,N_9054,N_9262);
and UO_838 (O_838,N_9334,N_9116);
nor UO_839 (O_839,N_9784,N_9514);
nand UO_840 (O_840,N_9267,N_9897);
nor UO_841 (O_841,N_9023,N_9672);
nor UO_842 (O_842,N_9778,N_9086);
nor UO_843 (O_843,N_9929,N_9764);
or UO_844 (O_844,N_9797,N_9118);
or UO_845 (O_845,N_9266,N_9762);
nor UO_846 (O_846,N_9923,N_9628);
nor UO_847 (O_847,N_9915,N_9059);
and UO_848 (O_848,N_9989,N_9375);
and UO_849 (O_849,N_9838,N_9179);
and UO_850 (O_850,N_9248,N_9915);
nand UO_851 (O_851,N_9402,N_9139);
or UO_852 (O_852,N_9906,N_9029);
nand UO_853 (O_853,N_9398,N_9141);
or UO_854 (O_854,N_9539,N_9963);
xor UO_855 (O_855,N_9013,N_9409);
or UO_856 (O_856,N_9627,N_9068);
or UO_857 (O_857,N_9198,N_9992);
xor UO_858 (O_858,N_9070,N_9246);
nand UO_859 (O_859,N_9511,N_9663);
nand UO_860 (O_860,N_9519,N_9602);
or UO_861 (O_861,N_9523,N_9414);
nand UO_862 (O_862,N_9183,N_9546);
nand UO_863 (O_863,N_9444,N_9538);
and UO_864 (O_864,N_9258,N_9604);
or UO_865 (O_865,N_9503,N_9980);
nor UO_866 (O_866,N_9861,N_9217);
nand UO_867 (O_867,N_9353,N_9391);
nor UO_868 (O_868,N_9472,N_9335);
nand UO_869 (O_869,N_9081,N_9762);
and UO_870 (O_870,N_9415,N_9341);
nand UO_871 (O_871,N_9914,N_9323);
nand UO_872 (O_872,N_9135,N_9745);
nand UO_873 (O_873,N_9322,N_9021);
nor UO_874 (O_874,N_9333,N_9141);
nor UO_875 (O_875,N_9824,N_9640);
and UO_876 (O_876,N_9231,N_9127);
nand UO_877 (O_877,N_9804,N_9932);
and UO_878 (O_878,N_9964,N_9110);
and UO_879 (O_879,N_9852,N_9740);
nor UO_880 (O_880,N_9544,N_9693);
and UO_881 (O_881,N_9811,N_9399);
and UO_882 (O_882,N_9360,N_9684);
nand UO_883 (O_883,N_9228,N_9463);
or UO_884 (O_884,N_9820,N_9897);
or UO_885 (O_885,N_9081,N_9905);
and UO_886 (O_886,N_9283,N_9519);
nand UO_887 (O_887,N_9312,N_9791);
and UO_888 (O_888,N_9724,N_9122);
nand UO_889 (O_889,N_9688,N_9279);
and UO_890 (O_890,N_9987,N_9906);
and UO_891 (O_891,N_9212,N_9650);
or UO_892 (O_892,N_9304,N_9700);
nand UO_893 (O_893,N_9963,N_9723);
nand UO_894 (O_894,N_9665,N_9768);
or UO_895 (O_895,N_9478,N_9515);
nand UO_896 (O_896,N_9778,N_9235);
or UO_897 (O_897,N_9948,N_9904);
nor UO_898 (O_898,N_9300,N_9513);
nand UO_899 (O_899,N_9950,N_9384);
and UO_900 (O_900,N_9110,N_9838);
or UO_901 (O_901,N_9700,N_9744);
nor UO_902 (O_902,N_9564,N_9008);
nand UO_903 (O_903,N_9767,N_9281);
and UO_904 (O_904,N_9596,N_9570);
nand UO_905 (O_905,N_9594,N_9658);
or UO_906 (O_906,N_9768,N_9803);
nor UO_907 (O_907,N_9540,N_9145);
and UO_908 (O_908,N_9058,N_9907);
and UO_909 (O_909,N_9986,N_9192);
or UO_910 (O_910,N_9393,N_9547);
nand UO_911 (O_911,N_9361,N_9330);
nor UO_912 (O_912,N_9916,N_9471);
nand UO_913 (O_913,N_9297,N_9134);
or UO_914 (O_914,N_9848,N_9346);
or UO_915 (O_915,N_9163,N_9446);
nor UO_916 (O_916,N_9059,N_9305);
or UO_917 (O_917,N_9437,N_9529);
and UO_918 (O_918,N_9924,N_9338);
nand UO_919 (O_919,N_9554,N_9441);
nor UO_920 (O_920,N_9528,N_9098);
and UO_921 (O_921,N_9807,N_9976);
or UO_922 (O_922,N_9000,N_9168);
and UO_923 (O_923,N_9155,N_9089);
nand UO_924 (O_924,N_9907,N_9609);
nor UO_925 (O_925,N_9022,N_9121);
nor UO_926 (O_926,N_9188,N_9759);
or UO_927 (O_927,N_9150,N_9741);
and UO_928 (O_928,N_9733,N_9249);
and UO_929 (O_929,N_9240,N_9897);
xnor UO_930 (O_930,N_9372,N_9674);
or UO_931 (O_931,N_9272,N_9922);
or UO_932 (O_932,N_9059,N_9251);
nand UO_933 (O_933,N_9520,N_9679);
and UO_934 (O_934,N_9422,N_9725);
or UO_935 (O_935,N_9345,N_9399);
nor UO_936 (O_936,N_9633,N_9111);
and UO_937 (O_937,N_9557,N_9987);
or UO_938 (O_938,N_9370,N_9389);
and UO_939 (O_939,N_9902,N_9691);
or UO_940 (O_940,N_9953,N_9903);
or UO_941 (O_941,N_9474,N_9890);
nand UO_942 (O_942,N_9272,N_9933);
nand UO_943 (O_943,N_9956,N_9676);
nand UO_944 (O_944,N_9520,N_9246);
or UO_945 (O_945,N_9410,N_9467);
and UO_946 (O_946,N_9773,N_9760);
and UO_947 (O_947,N_9547,N_9142);
nand UO_948 (O_948,N_9610,N_9519);
and UO_949 (O_949,N_9498,N_9673);
and UO_950 (O_950,N_9642,N_9505);
and UO_951 (O_951,N_9939,N_9532);
nor UO_952 (O_952,N_9676,N_9992);
or UO_953 (O_953,N_9753,N_9868);
nand UO_954 (O_954,N_9306,N_9122);
or UO_955 (O_955,N_9898,N_9063);
nand UO_956 (O_956,N_9286,N_9454);
nor UO_957 (O_957,N_9430,N_9610);
and UO_958 (O_958,N_9309,N_9850);
nor UO_959 (O_959,N_9329,N_9170);
or UO_960 (O_960,N_9846,N_9047);
and UO_961 (O_961,N_9866,N_9683);
nand UO_962 (O_962,N_9029,N_9278);
and UO_963 (O_963,N_9841,N_9866);
and UO_964 (O_964,N_9582,N_9826);
and UO_965 (O_965,N_9991,N_9537);
and UO_966 (O_966,N_9372,N_9147);
nor UO_967 (O_967,N_9560,N_9671);
nor UO_968 (O_968,N_9054,N_9456);
nor UO_969 (O_969,N_9461,N_9358);
and UO_970 (O_970,N_9858,N_9419);
and UO_971 (O_971,N_9288,N_9080);
and UO_972 (O_972,N_9296,N_9821);
and UO_973 (O_973,N_9135,N_9336);
xor UO_974 (O_974,N_9330,N_9425);
nand UO_975 (O_975,N_9525,N_9031);
and UO_976 (O_976,N_9777,N_9231);
and UO_977 (O_977,N_9336,N_9830);
or UO_978 (O_978,N_9892,N_9449);
nand UO_979 (O_979,N_9429,N_9545);
nand UO_980 (O_980,N_9147,N_9355);
nor UO_981 (O_981,N_9330,N_9953);
and UO_982 (O_982,N_9897,N_9615);
nand UO_983 (O_983,N_9870,N_9338);
and UO_984 (O_984,N_9644,N_9353);
nor UO_985 (O_985,N_9962,N_9617);
nand UO_986 (O_986,N_9806,N_9389);
nor UO_987 (O_987,N_9247,N_9143);
or UO_988 (O_988,N_9817,N_9170);
nor UO_989 (O_989,N_9263,N_9219);
nor UO_990 (O_990,N_9764,N_9308);
nand UO_991 (O_991,N_9246,N_9227);
nor UO_992 (O_992,N_9333,N_9625);
and UO_993 (O_993,N_9825,N_9407);
or UO_994 (O_994,N_9630,N_9467);
nor UO_995 (O_995,N_9165,N_9427);
or UO_996 (O_996,N_9041,N_9755);
nor UO_997 (O_997,N_9415,N_9205);
nor UO_998 (O_998,N_9279,N_9487);
nor UO_999 (O_999,N_9349,N_9873);
nand UO_1000 (O_1000,N_9367,N_9346);
nand UO_1001 (O_1001,N_9622,N_9576);
nor UO_1002 (O_1002,N_9144,N_9344);
nand UO_1003 (O_1003,N_9169,N_9801);
or UO_1004 (O_1004,N_9470,N_9709);
nand UO_1005 (O_1005,N_9510,N_9620);
nor UO_1006 (O_1006,N_9171,N_9864);
nand UO_1007 (O_1007,N_9517,N_9543);
nand UO_1008 (O_1008,N_9096,N_9243);
or UO_1009 (O_1009,N_9109,N_9666);
nor UO_1010 (O_1010,N_9437,N_9912);
nand UO_1011 (O_1011,N_9268,N_9981);
nand UO_1012 (O_1012,N_9786,N_9356);
or UO_1013 (O_1013,N_9367,N_9774);
nand UO_1014 (O_1014,N_9669,N_9864);
nor UO_1015 (O_1015,N_9884,N_9173);
nand UO_1016 (O_1016,N_9321,N_9428);
and UO_1017 (O_1017,N_9115,N_9153);
nor UO_1018 (O_1018,N_9093,N_9797);
nand UO_1019 (O_1019,N_9992,N_9527);
nor UO_1020 (O_1020,N_9182,N_9734);
and UO_1021 (O_1021,N_9861,N_9441);
nand UO_1022 (O_1022,N_9971,N_9569);
nor UO_1023 (O_1023,N_9547,N_9863);
nand UO_1024 (O_1024,N_9338,N_9013);
nor UO_1025 (O_1025,N_9326,N_9698);
and UO_1026 (O_1026,N_9285,N_9950);
nor UO_1027 (O_1027,N_9355,N_9180);
nor UO_1028 (O_1028,N_9293,N_9283);
and UO_1029 (O_1029,N_9398,N_9004);
nor UO_1030 (O_1030,N_9071,N_9800);
and UO_1031 (O_1031,N_9215,N_9716);
nand UO_1032 (O_1032,N_9899,N_9802);
nor UO_1033 (O_1033,N_9467,N_9457);
nand UO_1034 (O_1034,N_9196,N_9555);
nand UO_1035 (O_1035,N_9994,N_9755);
nor UO_1036 (O_1036,N_9204,N_9657);
or UO_1037 (O_1037,N_9588,N_9026);
nor UO_1038 (O_1038,N_9828,N_9405);
or UO_1039 (O_1039,N_9184,N_9875);
and UO_1040 (O_1040,N_9529,N_9491);
nand UO_1041 (O_1041,N_9981,N_9134);
nand UO_1042 (O_1042,N_9331,N_9035);
nand UO_1043 (O_1043,N_9299,N_9400);
nor UO_1044 (O_1044,N_9506,N_9369);
nand UO_1045 (O_1045,N_9116,N_9144);
and UO_1046 (O_1046,N_9287,N_9246);
nand UO_1047 (O_1047,N_9087,N_9339);
and UO_1048 (O_1048,N_9877,N_9324);
nand UO_1049 (O_1049,N_9747,N_9671);
nand UO_1050 (O_1050,N_9004,N_9322);
xor UO_1051 (O_1051,N_9640,N_9136);
nand UO_1052 (O_1052,N_9313,N_9634);
nor UO_1053 (O_1053,N_9224,N_9940);
nor UO_1054 (O_1054,N_9277,N_9826);
nor UO_1055 (O_1055,N_9891,N_9310);
nand UO_1056 (O_1056,N_9323,N_9851);
nand UO_1057 (O_1057,N_9373,N_9239);
and UO_1058 (O_1058,N_9739,N_9620);
nand UO_1059 (O_1059,N_9750,N_9648);
nand UO_1060 (O_1060,N_9399,N_9271);
or UO_1061 (O_1061,N_9468,N_9170);
or UO_1062 (O_1062,N_9342,N_9567);
nand UO_1063 (O_1063,N_9665,N_9239);
nor UO_1064 (O_1064,N_9023,N_9590);
nor UO_1065 (O_1065,N_9017,N_9953);
or UO_1066 (O_1066,N_9387,N_9545);
or UO_1067 (O_1067,N_9205,N_9595);
nor UO_1068 (O_1068,N_9049,N_9084);
nor UO_1069 (O_1069,N_9682,N_9119);
nand UO_1070 (O_1070,N_9632,N_9144);
or UO_1071 (O_1071,N_9675,N_9588);
and UO_1072 (O_1072,N_9975,N_9995);
and UO_1073 (O_1073,N_9399,N_9403);
nand UO_1074 (O_1074,N_9441,N_9382);
or UO_1075 (O_1075,N_9596,N_9215);
nand UO_1076 (O_1076,N_9760,N_9501);
or UO_1077 (O_1077,N_9166,N_9252);
nand UO_1078 (O_1078,N_9433,N_9704);
nor UO_1079 (O_1079,N_9928,N_9480);
and UO_1080 (O_1080,N_9726,N_9472);
nor UO_1081 (O_1081,N_9468,N_9197);
and UO_1082 (O_1082,N_9414,N_9403);
nor UO_1083 (O_1083,N_9160,N_9439);
and UO_1084 (O_1084,N_9520,N_9373);
and UO_1085 (O_1085,N_9588,N_9387);
xor UO_1086 (O_1086,N_9856,N_9602);
nor UO_1087 (O_1087,N_9531,N_9662);
nor UO_1088 (O_1088,N_9431,N_9352);
or UO_1089 (O_1089,N_9511,N_9433);
and UO_1090 (O_1090,N_9478,N_9069);
xnor UO_1091 (O_1091,N_9599,N_9124);
nor UO_1092 (O_1092,N_9651,N_9874);
and UO_1093 (O_1093,N_9400,N_9272);
or UO_1094 (O_1094,N_9794,N_9677);
nand UO_1095 (O_1095,N_9781,N_9607);
nand UO_1096 (O_1096,N_9562,N_9486);
nand UO_1097 (O_1097,N_9170,N_9002);
and UO_1098 (O_1098,N_9215,N_9317);
and UO_1099 (O_1099,N_9199,N_9310);
and UO_1100 (O_1100,N_9993,N_9291);
nor UO_1101 (O_1101,N_9081,N_9372);
nor UO_1102 (O_1102,N_9238,N_9750);
or UO_1103 (O_1103,N_9559,N_9415);
and UO_1104 (O_1104,N_9353,N_9277);
nand UO_1105 (O_1105,N_9582,N_9950);
or UO_1106 (O_1106,N_9001,N_9260);
nand UO_1107 (O_1107,N_9155,N_9983);
and UO_1108 (O_1108,N_9169,N_9104);
and UO_1109 (O_1109,N_9783,N_9071);
nor UO_1110 (O_1110,N_9099,N_9145);
nand UO_1111 (O_1111,N_9294,N_9130);
and UO_1112 (O_1112,N_9080,N_9090);
and UO_1113 (O_1113,N_9675,N_9509);
and UO_1114 (O_1114,N_9798,N_9874);
nand UO_1115 (O_1115,N_9200,N_9067);
nand UO_1116 (O_1116,N_9683,N_9481);
or UO_1117 (O_1117,N_9175,N_9166);
nand UO_1118 (O_1118,N_9632,N_9336);
or UO_1119 (O_1119,N_9643,N_9219);
nand UO_1120 (O_1120,N_9750,N_9710);
or UO_1121 (O_1121,N_9209,N_9810);
or UO_1122 (O_1122,N_9902,N_9341);
nor UO_1123 (O_1123,N_9483,N_9945);
and UO_1124 (O_1124,N_9633,N_9295);
and UO_1125 (O_1125,N_9988,N_9956);
and UO_1126 (O_1126,N_9764,N_9619);
or UO_1127 (O_1127,N_9370,N_9230);
nand UO_1128 (O_1128,N_9780,N_9096);
and UO_1129 (O_1129,N_9115,N_9992);
nand UO_1130 (O_1130,N_9086,N_9690);
and UO_1131 (O_1131,N_9746,N_9177);
nand UO_1132 (O_1132,N_9087,N_9529);
nand UO_1133 (O_1133,N_9642,N_9272);
nand UO_1134 (O_1134,N_9282,N_9436);
xnor UO_1135 (O_1135,N_9113,N_9075);
or UO_1136 (O_1136,N_9747,N_9684);
nand UO_1137 (O_1137,N_9244,N_9343);
and UO_1138 (O_1138,N_9804,N_9796);
or UO_1139 (O_1139,N_9326,N_9763);
nor UO_1140 (O_1140,N_9698,N_9728);
or UO_1141 (O_1141,N_9531,N_9005);
and UO_1142 (O_1142,N_9911,N_9706);
nor UO_1143 (O_1143,N_9074,N_9503);
nor UO_1144 (O_1144,N_9216,N_9153);
or UO_1145 (O_1145,N_9475,N_9810);
nor UO_1146 (O_1146,N_9195,N_9778);
nor UO_1147 (O_1147,N_9186,N_9306);
nand UO_1148 (O_1148,N_9334,N_9070);
nand UO_1149 (O_1149,N_9285,N_9250);
nand UO_1150 (O_1150,N_9896,N_9973);
nor UO_1151 (O_1151,N_9000,N_9995);
or UO_1152 (O_1152,N_9695,N_9245);
or UO_1153 (O_1153,N_9645,N_9677);
and UO_1154 (O_1154,N_9635,N_9582);
nand UO_1155 (O_1155,N_9968,N_9673);
and UO_1156 (O_1156,N_9483,N_9436);
nand UO_1157 (O_1157,N_9512,N_9731);
and UO_1158 (O_1158,N_9423,N_9537);
nor UO_1159 (O_1159,N_9133,N_9688);
nor UO_1160 (O_1160,N_9084,N_9911);
or UO_1161 (O_1161,N_9823,N_9930);
nand UO_1162 (O_1162,N_9737,N_9992);
or UO_1163 (O_1163,N_9691,N_9580);
nand UO_1164 (O_1164,N_9678,N_9402);
nor UO_1165 (O_1165,N_9554,N_9377);
nand UO_1166 (O_1166,N_9233,N_9400);
or UO_1167 (O_1167,N_9966,N_9440);
nor UO_1168 (O_1168,N_9742,N_9156);
or UO_1169 (O_1169,N_9623,N_9811);
nand UO_1170 (O_1170,N_9897,N_9623);
nor UO_1171 (O_1171,N_9503,N_9213);
or UO_1172 (O_1172,N_9806,N_9418);
nand UO_1173 (O_1173,N_9591,N_9114);
nor UO_1174 (O_1174,N_9896,N_9648);
and UO_1175 (O_1175,N_9298,N_9182);
nand UO_1176 (O_1176,N_9289,N_9920);
and UO_1177 (O_1177,N_9100,N_9917);
nand UO_1178 (O_1178,N_9599,N_9781);
and UO_1179 (O_1179,N_9759,N_9342);
and UO_1180 (O_1180,N_9401,N_9520);
or UO_1181 (O_1181,N_9996,N_9224);
and UO_1182 (O_1182,N_9585,N_9207);
nor UO_1183 (O_1183,N_9280,N_9576);
and UO_1184 (O_1184,N_9499,N_9998);
or UO_1185 (O_1185,N_9364,N_9321);
or UO_1186 (O_1186,N_9176,N_9350);
and UO_1187 (O_1187,N_9545,N_9895);
nand UO_1188 (O_1188,N_9545,N_9945);
nand UO_1189 (O_1189,N_9986,N_9782);
and UO_1190 (O_1190,N_9675,N_9898);
nand UO_1191 (O_1191,N_9772,N_9598);
nand UO_1192 (O_1192,N_9408,N_9933);
or UO_1193 (O_1193,N_9924,N_9072);
or UO_1194 (O_1194,N_9627,N_9180);
nor UO_1195 (O_1195,N_9187,N_9204);
nor UO_1196 (O_1196,N_9147,N_9586);
nor UO_1197 (O_1197,N_9859,N_9691);
and UO_1198 (O_1198,N_9647,N_9691);
or UO_1199 (O_1199,N_9618,N_9795);
nor UO_1200 (O_1200,N_9620,N_9816);
or UO_1201 (O_1201,N_9579,N_9546);
or UO_1202 (O_1202,N_9291,N_9655);
nor UO_1203 (O_1203,N_9314,N_9215);
or UO_1204 (O_1204,N_9389,N_9009);
nand UO_1205 (O_1205,N_9868,N_9403);
nor UO_1206 (O_1206,N_9855,N_9683);
or UO_1207 (O_1207,N_9698,N_9045);
nor UO_1208 (O_1208,N_9946,N_9299);
nand UO_1209 (O_1209,N_9389,N_9639);
xnor UO_1210 (O_1210,N_9376,N_9118);
nor UO_1211 (O_1211,N_9910,N_9641);
and UO_1212 (O_1212,N_9214,N_9315);
and UO_1213 (O_1213,N_9491,N_9653);
nand UO_1214 (O_1214,N_9942,N_9470);
and UO_1215 (O_1215,N_9945,N_9655);
nand UO_1216 (O_1216,N_9554,N_9805);
or UO_1217 (O_1217,N_9299,N_9801);
nand UO_1218 (O_1218,N_9701,N_9760);
and UO_1219 (O_1219,N_9095,N_9739);
or UO_1220 (O_1220,N_9273,N_9859);
and UO_1221 (O_1221,N_9689,N_9824);
or UO_1222 (O_1222,N_9044,N_9102);
or UO_1223 (O_1223,N_9976,N_9333);
nor UO_1224 (O_1224,N_9693,N_9758);
or UO_1225 (O_1225,N_9692,N_9991);
nand UO_1226 (O_1226,N_9461,N_9163);
nand UO_1227 (O_1227,N_9074,N_9396);
or UO_1228 (O_1228,N_9199,N_9315);
and UO_1229 (O_1229,N_9476,N_9877);
nor UO_1230 (O_1230,N_9198,N_9487);
or UO_1231 (O_1231,N_9862,N_9410);
nand UO_1232 (O_1232,N_9789,N_9031);
or UO_1233 (O_1233,N_9648,N_9050);
nand UO_1234 (O_1234,N_9829,N_9974);
and UO_1235 (O_1235,N_9630,N_9545);
nor UO_1236 (O_1236,N_9572,N_9220);
nor UO_1237 (O_1237,N_9142,N_9110);
and UO_1238 (O_1238,N_9513,N_9455);
nor UO_1239 (O_1239,N_9917,N_9815);
nand UO_1240 (O_1240,N_9341,N_9777);
nand UO_1241 (O_1241,N_9655,N_9523);
nand UO_1242 (O_1242,N_9509,N_9855);
or UO_1243 (O_1243,N_9590,N_9393);
xnor UO_1244 (O_1244,N_9600,N_9768);
nor UO_1245 (O_1245,N_9287,N_9839);
nor UO_1246 (O_1246,N_9280,N_9263);
or UO_1247 (O_1247,N_9891,N_9692);
or UO_1248 (O_1248,N_9694,N_9238);
nor UO_1249 (O_1249,N_9600,N_9013);
or UO_1250 (O_1250,N_9347,N_9555);
or UO_1251 (O_1251,N_9156,N_9291);
nand UO_1252 (O_1252,N_9895,N_9148);
nand UO_1253 (O_1253,N_9772,N_9500);
or UO_1254 (O_1254,N_9339,N_9282);
nand UO_1255 (O_1255,N_9538,N_9144);
nand UO_1256 (O_1256,N_9100,N_9585);
nor UO_1257 (O_1257,N_9331,N_9884);
and UO_1258 (O_1258,N_9373,N_9138);
nor UO_1259 (O_1259,N_9065,N_9147);
nand UO_1260 (O_1260,N_9316,N_9472);
and UO_1261 (O_1261,N_9020,N_9180);
nor UO_1262 (O_1262,N_9221,N_9886);
nand UO_1263 (O_1263,N_9662,N_9569);
nor UO_1264 (O_1264,N_9000,N_9656);
and UO_1265 (O_1265,N_9430,N_9271);
nor UO_1266 (O_1266,N_9199,N_9375);
or UO_1267 (O_1267,N_9541,N_9127);
nand UO_1268 (O_1268,N_9179,N_9170);
nor UO_1269 (O_1269,N_9523,N_9347);
and UO_1270 (O_1270,N_9244,N_9162);
and UO_1271 (O_1271,N_9635,N_9497);
and UO_1272 (O_1272,N_9388,N_9476);
or UO_1273 (O_1273,N_9656,N_9034);
nand UO_1274 (O_1274,N_9154,N_9529);
nand UO_1275 (O_1275,N_9037,N_9945);
and UO_1276 (O_1276,N_9303,N_9287);
nand UO_1277 (O_1277,N_9259,N_9021);
nor UO_1278 (O_1278,N_9761,N_9754);
nor UO_1279 (O_1279,N_9105,N_9972);
and UO_1280 (O_1280,N_9114,N_9430);
nand UO_1281 (O_1281,N_9105,N_9027);
nand UO_1282 (O_1282,N_9389,N_9376);
nor UO_1283 (O_1283,N_9203,N_9554);
nand UO_1284 (O_1284,N_9325,N_9367);
nand UO_1285 (O_1285,N_9829,N_9668);
or UO_1286 (O_1286,N_9447,N_9513);
and UO_1287 (O_1287,N_9992,N_9827);
or UO_1288 (O_1288,N_9704,N_9015);
nor UO_1289 (O_1289,N_9524,N_9760);
nand UO_1290 (O_1290,N_9897,N_9922);
or UO_1291 (O_1291,N_9564,N_9322);
and UO_1292 (O_1292,N_9901,N_9319);
nor UO_1293 (O_1293,N_9102,N_9012);
nand UO_1294 (O_1294,N_9641,N_9251);
nor UO_1295 (O_1295,N_9181,N_9958);
nor UO_1296 (O_1296,N_9276,N_9358);
nor UO_1297 (O_1297,N_9576,N_9187);
nor UO_1298 (O_1298,N_9381,N_9287);
or UO_1299 (O_1299,N_9536,N_9016);
nor UO_1300 (O_1300,N_9553,N_9586);
nor UO_1301 (O_1301,N_9176,N_9487);
nor UO_1302 (O_1302,N_9445,N_9527);
or UO_1303 (O_1303,N_9733,N_9385);
or UO_1304 (O_1304,N_9879,N_9381);
or UO_1305 (O_1305,N_9320,N_9605);
and UO_1306 (O_1306,N_9086,N_9885);
and UO_1307 (O_1307,N_9523,N_9402);
and UO_1308 (O_1308,N_9226,N_9936);
nand UO_1309 (O_1309,N_9381,N_9980);
or UO_1310 (O_1310,N_9340,N_9513);
and UO_1311 (O_1311,N_9635,N_9779);
nor UO_1312 (O_1312,N_9894,N_9347);
nor UO_1313 (O_1313,N_9539,N_9175);
or UO_1314 (O_1314,N_9884,N_9095);
nand UO_1315 (O_1315,N_9895,N_9316);
nor UO_1316 (O_1316,N_9810,N_9753);
or UO_1317 (O_1317,N_9581,N_9208);
nand UO_1318 (O_1318,N_9165,N_9131);
or UO_1319 (O_1319,N_9262,N_9355);
nor UO_1320 (O_1320,N_9377,N_9357);
and UO_1321 (O_1321,N_9993,N_9452);
and UO_1322 (O_1322,N_9121,N_9958);
or UO_1323 (O_1323,N_9634,N_9266);
or UO_1324 (O_1324,N_9103,N_9881);
nor UO_1325 (O_1325,N_9642,N_9985);
or UO_1326 (O_1326,N_9018,N_9282);
and UO_1327 (O_1327,N_9147,N_9302);
nand UO_1328 (O_1328,N_9498,N_9000);
nand UO_1329 (O_1329,N_9796,N_9831);
nand UO_1330 (O_1330,N_9014,N_9585);
or UO_1331 (O_1331,N_9840,N_9228);
and UO_1332 (O_1332,N_9327,N_9093);
or UO_1333 (O_1333,N_9494,N_9310);
nand UO_1334 (O_1334,N_9196,N_9409);
and UO_1335 (O_1335,N_9814,N_9716);
or UO_1336 (O_1336,N_9969,N_9981);
or UO_1337 (O_1337,N_9965,N_9765);
nor UO_1338 (O_1338,N_9496,N_9158);
nand UO_1339 (O_1339,N_9354,N_9080);
nor UO_1340 (O_1340,N_9419,N_9898);
or UO_1341 (O_1341,N_9369,N_9291);
nor UO_1342 (O_1342,N_9161,N_9083);
nor UO_1343 (O_1343,N_9759,N_9120);
nand UO_1344 (O_1344,N_9345,N_9907);
nor UO_1345 (O_1345,N_9466,N_9604);
nand UO_1346 (O_1346,N_9462,N_9939);
nor UO_1347 (O_1347,N_9449,N_9613);
or UO_1348 (O_1348,N_9809,N_9211);
or UO_1349 (O_1349,N_9678,N_9030);
and UO_1350 (O_1350,N_9079,N_9033);
nand UO_1351 (O_1351,N_9200,N_9874);
and UO_1352 (O_1352,N_9215,N_9105);
and UO_1353 (O_1353,N_9998,N_9352);
and UO_1354 (O_1354,N_9690,N_9563);
or UO_1355 (O_1355,N_9291,N_9763);
nor UO_1356 (O_1356,N_9237,N_9115);
nand UO_1357 (O_1357,N_9683,N_9188);
or UO_1358 (O_1358,N_9811,N_9159);
nor UO_1359 (O_1359,N_9581,N_9288);
nand UO_1360 (O_1360,N_9447,N_9592);
and UO_1361 (O_1361,N_9345,N_9377);
and UO_1362 (O_1362,N_9074,N_9790);
nand UO_1363 (O_1363,N_9873,N_9689);
nor UO_1364 (O_1364,N_9435,N_9464);
or UO_1365 (O_1365,N_9604,N_9320);
nor UO_1366 (O_1366,N_9413,N_9521);
and UO_1367 (O_1367,N_9338,N_9098);
or UO_1368 (O_1368,N_9426,N_9342);
nand UO_1369 (O_1369,N_9413,N_9075);
nand UO_1370 (O_1370,N_9055,N_9457);
nor UO_1371 (O_1371,N_9904,N_9369);
or UO_1372 (O_1372,N_9031,N_9330);
and UO_1373 (O_1373,N_9634,N_9283);
nor UO_1374 (O_1374,N_9444,N_9863);
nand UO_1375 (O_1375,N_9090,N_9847);
and UO_1376 (O_1376,N_9226,N_9501);
and UO_1377 (O_1377,N_9781,N_9582);
and UO_1378 (O_1378,N_9384,N_9235);
nand UO_1379 (O_1379,N_9383,N_9621);
nor UO_1380 (O_1380,N_9952,N_9671);
or UO_1381 (O_1381,N_9446,N_9356);
nand UO_1382 (O_1382,N_9165,N_9579);
nand UO_1383 (O_1383,N_9235,N_9600);
and UO_1384 (O_1384,N_9847,N_9825);
nand UO_1385 (O_1385,N_9506,N_9412);
and UO_1386 (O_1386,N_9571,N_9655);
nand UO_1387 (O_1387,N_9086,N_9662);
and UO_1388 (O_1388,N_9600,N_9537);
nor UO_1389 (O_1389,N_9650,N_9599);
and UO_1390 (O_1390,N_9833,N_9214);
and UO_1391 (O_1391,N_9986,N_9068);
nor UO_1392 (O_1392,N_9123,N_9987);
nand UO_1393 (O_1393,N_9237,N_9879);
or UO_1394 (O_1394,N_9605,N_9757);
nor UO_1395 (O_1395,N_9472,N_9721);
or UO_1396 (O_1396,N_9503,N_9645);
and UO_1397 (O_1397,N_9453,N_9297);
and UO_1398 (O_1398,N_9035,N_9736);
nand UO_1399 (O_1399,N_9241,N_9343);
nand UO_1400 (O_1400,N_9412,N_9771);
nor UO_1401 (O_1401,N_9343,N_9035);
nand UO_1402 (O_1402,N_9761,N_9627);
nand UO_1403 (O_1403,N_9316,N_9858);
and UO_1404 (O_1404,N_9002,N_9856);
nor UO_1405 (O_1405,N_9711,N_9369);
and UO_1406 (O_1406,N_9413,N_9934);
nand UO_1407 (O_1407,N_9865,N_9411);
and UO_1408 (O_1408,N_9492,N_9856);
and UO_1409 (O_1409,N_9109,N_9081);
and UO_1410 (O_1410,N_9411,N_9325);
and UO_1411 (O_1411,N_9234,N_9859);
nor UO_1412 (O_1412,N_9675,N_9656);
and UO_1413 (O_1413,N_9678,N_9676);
nand UO_1414 (O_1414,N_9193,N_9854);
or UO_1415 (O_1415,N_9039,N_9885);
or UO_1416 (O_1416,N_9004,N_9407);
or UO_1417 (O_1417,N_9747,N_9833);
or UO_1418 (O_1418,N_9858,N_9462);
or UO_1419 (O_1419,N_9429,N_9760);
nor UO_1420 (O_1420,N_9932,N_9035);
or UO_1421 (O_1421,N_9526,N_9310);
and UO_1422 (O_1422,N_9030,N_9448);
xnor UO_1423 (O_1423,N_9617,N_9329);
or UO_1424 (O_1424,N_9040,N_9745);
or UO_1425 (O_1425,N_9483,N_9680);
or UO_1426 (O_1426,N_9546,N_9523);
nand UO_1427 (O_1427,N_9805,N_9049);
nor UO_1428 (O_1428,N_9144,N_9015);
or UO_1429 (O_1429,N_9576,N_9193);
nor UO_1430 (O_1430,N_9494,N_9161);
nand UO_1431 (O_1431,N_9342,N_9799);
or UO_1432 (O_1432,N_9839,N_9932);
and UO_1433 (O_1433,N_9482,N_9676);
nor UO_1434 (O_1434,N_9810,N_9173);
or UO_1435 (O_1435,N_9683,N_9203);
or UO_1436 (O_1436,N_9633,N_9748);
and UO_1437 (O_1437,N_9340,N_9306);
nand UO_1438 (O_1438,N_9683,N_9404);
or UO_1439 (O_1439,N_9551,N_9122);
or UO_1440 (O_1440,N_9446,N_9271);
nor UO_1441 (O_1441,N_9990,N_9726);
and UO_1442 (O_1442,N_9178,N_9620);
or UO_1443 (O_1443,N_9606,N_9366);
or UO_1444 (O_1444,N_9891,N_9189);
and UO_1445 (O_1445,N_9575,N_9721);
and UO_1446 (O_1446,N_9074,N_9368);
nand UO_1447 (O_1447,N_9958,N_9842);
nand UO_1448 (O_1448,N_9912,N_9069);
nor UO_1449 (O_1449,N_9654,N_9055);
or UO_1450 (O_1450,N_9344,N_9289);
nand UO_1451 (O_1451,N_9775,N_9939);
and UO_1452 (O_1452,N_9936,N_9134);
and UO_1453 (O_1453,N_9445,N_9104);
nor UO_1454 (O_1454,N_9648,N_9727);
and UO_1455 (O_1455,N_9885,N_9819);
nand UO_1456 (O_1456,N_9259,N_9451);
nand UO_1457 (O_1457,N_9024,N_9553);
or UO_1458 (O_1458,N_9483,N_9332);
nor UO_1459 (O_1459,N_9134,N_9945);
nor UO_1460 (O_1460,N_9071,N_9211);
or UO_1461 (O_1461,N_9330,N_9963);
and UO_1462 (O_1462,N_9425,N_9316);
or UO_1463 (O_1463,N_9000,N_9539);
nor UO_1464 (O_1464,N_9702,N_9545);
nor UO_1465 (O_1465,N_9558,N_9902);
or UO_1466 (O_1466,N_9442,N_9394);
and UO_1467 (O_1467,N_9585,N_9154);
nor UO_1468 (O_1468,N_9665,N_9031);
nor UO_1469 (O_1469,N_9190,N_9096);
nand UO_1470 (O_1470,N_9545,N_9001);
or UO_1471 (O_1471,N_9148,N_9793);
nand UO_1472 (O_1472,N_9570,N_9261);
or UO_1473 (O_1473,N_9432,N_9382);
nor UO_1474 (O_1474,N_9585,N_9912);
nor UO_1475 (O_1475,N_9743,N_9039);
and UO_1476 (O_1476,N_9642,N_9972);
nor UO_1477 (O_1477,N_9709,N_9479);
nor UO_1478 (O_1478,N_9274,N_9354);
nand UO_1479 (O_1479,N_9333,N_9462);
or UO_1480 (O_1480,N_9177,N_9610);
or UO_1481 (O_1481,N_9765,N_9966);
nand UO_1482 (O_1482,N_9587,N_9576);
nor UO_1483 (O_1483,N_9679,N_9791);
and UO_1484 (O_1484,N_9159,N_9891);
or UO_1485 (O_1485,N_9166,N_9504);
and UO_1486 (O_1486,N_9712,N_9745);
and UO_1487 (O_1487,N_9671,N_9261);
nor UO_1488 (O_1488,N_9492,N_9823);
nor UO_1489 (O_1489,N_9072,N_9069);
and UO_1490 (O_1490,N_9545,N_9440);
and UO_1491 (O_1491,N_9798,N_9934);
nor UO_1492 (O_1492,N_9180,N_9787);
or UO_1493 (O_1493,N_9039,N_9488);
or UO_1494 (O_1494,N_9931,N_9656);
nand UO_1495 (O_1495,N_9706,N_9563);
and UO_1496 (O_1496,N_9474,N_9253);
or UO_1497 (O_1497,N_9735,N_9216);
and UO_1498 (O_1498,N_9640,N_9602);
and UO_1499 (O_1499,N_9298,N_9171);
endmodule