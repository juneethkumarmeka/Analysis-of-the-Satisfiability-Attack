module basic_750_5000_1000_5_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_730,In_308);
nand U1 (N_1,In_437,In_131);
and U2 (N_2,In_524,In_438);
nand U3 (N_3,In_707,In_386);
or U4 (N_4,In_255,In_412);
or U5 (N_5,In_679,In_64);
nor U6 (N_6,In_315,In_740);
nor U7 (N_7,In_461,In_464);
nand U8 (N_8,In_112,In_663);
nor U9 (N_9,In_535,In_288);
nor U10 (N_10,In_132,In_682);
xor U11 (N_11,In_674,In_130);
nand U12 (N_12,In_257,In_172);
and U13 (N_13,In_743,In_459);
and U14 (N_14,In_676,In_606);
or U15 (N_15,In_741,In_197);
nand U16 (N_16,In_443,In_7);
or U17 (N_17,In_310,In_258);
nor U18 (N_18,In_168,In_700);
nand U19 (N_19,In_235,In_173);
or U20 (N_20,In_403,In_605);
nand U21 (N_21,In_693,In_244);
or U22 (N_22,In_346,In_328);
or U23 (N_23,In_721,In_465);
or U24 (N_24,In_436,In_242);
nand U25 (N_25,In_440,In_297);
nor U26 (N_26,In_542,In_594);
nor U27 (N_27,In_311,In_445);
nor U28 (N_28,In_14,In_336);
and U29 (N_29,In_17,In_215);
and U30 (N_30,In_536,In_234);
nor U31 (N_31,In_52,In_656);
and U32 (N_32,In_673,In_614);
and U33 (N_33,In_636,In_260);
or U34 (N_34,In_245,In_563);
nand U35 (N_35,In_141,In_347);
xor U36 (N_36,In_217,In_304);
nor U37 (N_37,In_98,In_302);
nor U38 (N_38,In_156,In_24);
nor U39 (N_39,In_632,In_425);
nor U40 (N_40,In_675,In_520);
nand U41 (N_41,In_314,In_405);
xnor U42 (N_42,In_121,In_239);
and U43 (N_43,In_249,In_195);
and U44 (N_44,In_36,In_610);
or U45 (N_45,In_192,In_163);
xnor U46 (N_46,In_56,In_486);
or U47 (N_47,In_479,In_62);
xnor U48 (N_48,In_724,In_313);
xor U49 (N_49,In_106,In_564);
or U50 (N_50,In_576,In_517);
and U51 (N_51,In_294,In_529);
nand U52 (N_52,In_541,In_96);
xor U53 (N_53,In_570,In_312);
xor U54 (N_54,In_387,In_414);
nand U55 (N_55,In_410,In_198);
or U56 (N_56,In_203,In_609);
nor U57 (N_57,In_122,In_621);
nor U58 (N_58,In_522,In_77);
nor U59 (N_59,In_363,In_646);
nand U60 (N_60,In_696,In_38);
nand U61 (N_61,In_635,In_76);
nor U62 (N_62,In_667,In_75);
and U63 (N_63,In_323,In_688);
nand U64 (N_64,In_366,In_429);
and U65 (N_65,In_644,In_589);
nor U66 (N_66,In_345,In_449);
or U67 (N_67,In_413,In_701);
and U68 (N_68,In_149,In_394);
and U69 (N_69,In_321,In_108);
or U70 (N_70,In_322,In_583);
xnor U71 (N_71,In_409,In_422);
xor U72 (N_72,In_109,In_680);
nand U73 (N_73,In_598,In_165);
and U74 (N_74,In_509,In_44);
and U75 (N_75,In_82,In_558);
xor U76 (N_76,In_400,In_418);
nand U77 (N_77,In_254,In_97);
nand U78 (N_78,In_483,In_556);
or U79 (N_79,In_424,In_608);
nor U80 (N_80,In_467,In_23);
xnor U81 (N_81,In_351,In_274);
and U82 (N_82,In_485,In_319);
xor U83 (N_83,In_379,In_247);
and U84 (N_84,In_538,In_451);
and U85 (N_85,In_9,In_175);
and U86 (N_86,In_284,In_374);
nor U87 (N_87,In_63,In_722);
xor U88 (N_88,In_623,In_123);
or U89 (N_89,In_665,In_531);
or U90 (N_90,In_708,In_706);
nor U91 (N_91,In_169,In_159);
or U92 (N_92,In_300,In_320);
nor U93 (N_93,In_388,In_177);
or U94 (N_94,In_602,In_162);
nor U95 (N_95,In_362,In_478);
or U96 (N_96,In_349,In_597);
xnor U97 (N_97,In_432,In_199);
or U98 (N_98,In_584,In_746);
or U99 (N_99,In_411,In_627);
or U100 (N_100,In_607,In_19);
nor U101 (N_101,In_715,In_678);
nand U102 (N_102,In_622,In_580);
nand U103 (N_103,In_89,In_246);
xor U104 (N_104,In_396,In_113);
xnor U105 (N_105,In_470,In_342);
nor U106 (N_106,In_37,In_657);
nand U107 (N_107,In_110,In_219);
or U108 (N_108,In_74,In_725);
or U109 (N_109,In_380,In_442);
or U110 (N_110,In_480,In_10);
and U111 (N_111,In_214,In_93);
or U112 (N_112,In_160,In_629);
and U113 (N_113,In_572,In_6);
xor U114 (N_114,In_80,In_732);
nor U115 (N_115,In_226,In_67);
nor U116 (N_116,In_184,In_687);
nor U117 (N_117,In_174,In_595);
nor U118 (N_118,In_381,In_651);
nor U119 (N_119,In_309,In_466);
nand U120 (N_120,In_3,In_684);
and U121 (N_121,In_279,In_428);
or U122 (N_122,In_474,In_265);
nand U123 (N_123,In_238,In_333);
or U124 (N_124,In_637,In_317);
or U125 (N_125,In_638,In_650);
and U126 (N_126,In_86,In_12);
nor U127 (N_127,In_664,In_454);
or U128 (N_128,In_143,In_277);
or U129 (N_129,In_115,In_747);
nor U130 (N_130,In_293,In_699);
nand U131 (N_131,In_117,In_554);
xor U132 (N_132,In_427,In_213);
nor U133 (N_133,In_551,In_545);
nand U134 (N_134,In_139,In_72);
nand U135 (N_135,In_138,In_25);
or U136 (N_136,In_625,In_224);
and U137 (N_137,In_515,In_187);
nand U138 (N_138,In_393,In_530);
and U139 (N_139,In_568,In_230);
nor U140 (N_140,In_45,In_201);
xor U141 (N_141,In_221,In_473);
nand U142 (N_142,In_434,In_167);
xnor U143 (N_143,In_471,In_487);
nand U144 (N_144,In_733,In_189);
xor U145 (N_145,In_671,In_736);
nand U146 (N_146,In_326,In_469);
and U147 (N_147,In_298,In_592);
nor U148 (N_148,In_516,In_497);
nor U149 (N_149,In_40,In_618);
or U150 (N_150,In_280,In_292);
nor U151 (N_151,In_291,In_276);
and U152 (N_152,In_70,In_237);
or U153 (N_153,In_419,In_344);
and U154 (N_154,In_301,In_401);
or U155 (N_155,In_670,In_513);
xnor U156 (N_156,In_719,In_227);
or U157 (N_157,In_502,In_229);
nor U158 (N_158,In_4,In_423);
or U159 (N_159,In_188,In_218);
or U160 (N_160,In_640,In_271);
nand U161 (N_161,In_18,In_689);
and U162 (N_162,In_281,In_233);
nor U163 (N_163,In_28,In_200);
or U164 (N_164,In_452,In_735);
xor U165 (N_165,In_361,In_5);
nand U166 (N_166,In_532,In_99);
nand U167 (N_167,In_518,In_335);
nor U168 (N_168,In_431,In_601);
and U169 (N_169,In_626,In_243);
xor U170 (N_170,In_713,In_241);
or U171 (N_171,In_153,In_661);
or U172 (N_172,In_140,In_78);
or U173 (N_173,In_225,In_378);
xor U174 (N_174,In_103,In_739);
nor U175 (N_175,In_508,In_357);
or U176 (N_176,In_496,In_107);
nor U177 (N_177,In_116,In_698);
and U178 (N_178,In_142,In_718);
nor U179 (N_179,In_441,In_41);
nor U180 (N_180,In_430,In_204);
and U181 (N_181,In_211,In_426);
and U182 (N_182,In_631,In_539);
nor U183 (N_183,In_543,In_416);
nor U184 (N_184,In_561,In_223);
or U185 (N_185,In_332,In_494);
nand U186 (N_186,In_642,In_446);
or U187 (N_187,In_668,In_194);
and U188 (N_188,In_182,In_34);
and U189 (N_189,In_49,In_578);
and U190 (N_190,In_190,In_295);
nand U191 (N_191,In_47,In_73);
or U192 (N_192,In_240,In_666);
nand U193 (N_193,In_95,In_591);
nor U194 (N_194,In_8,In_712);
and U195 (N_195,In_559,In_620);
nand U196 (N_196,In_514,In_385);
or U197 (N_197,In_544,In_653);
nor U198 (N_198,In_358,In_392);
and U199 (N_199,In_398,In_2);
nand U200 (N_200,In_397,In_453);
xor U201 (N_201,In_161,In_286);
nor U202 (N_202,In_519,In_35);
or U203 (N_203,In_571,In_283);
and U204 (N_204,In_596,In_216);
or U205 (N_205,In_402,In_526);
or U206 (N_206,In_185,In_261);
xnor U207 (N_207,In_340,In_58);
or U208 (N_208,In_649,In_354);
xnor U209 (N_209,In_127,In_222);
nor U210 (N_210,In_586,In_683);
nand U211 (N_211,In_125,In_692);
nand U212 (N_212,In_81,In_590);
and U213 (N_213,In_90,In_84);
or U214 (N_214,In_703,In_92);
and U215 (N_215,In_528,In_507);
nand U216 (N_216,In_726,In_250);
or U217 (N_217,In_417,In_33);
nand U218 (N_218,In_266,In_376);
and U219 (N_219,In_369,In_579);
nand U220 (N_220,In_390,In_498);
and U221 (N_221,In_729,In_348);
nand U222 (N_222,In_71,In_421);
and U223 (N_223,In_171,In_150);
or U224 (N_224,In_499,In_15);
or U225 (N_225,In_124,In_263);
or U226 (N_226,In_482,In_491);
nand U227 (N_227,In_85,In_359);
nor U228 (N_228,In_435,In_654);
and U229 (N_229,In_748,In_450);
or U230 (N_230,In_555,In_329);
nor U231 (N_231,In_296,In_709);
and U232 (N_232,In_61,In_617);
or U233 (N_233,In_737,In_447);
xnor U234 (N_234,In_433,In_476);
nand U235 (N_235,In_128,In_324);
xor U236 (N_236,In_231,In_119);
nor U237 (N_237,In_253,In_59);
or U238 (N_238,In_460,In_270);
nor U239 (N_239,In_521,In_547);
nor U240 (N_240,In_269,In_339);
nand U241 (N_241,In_285,In_180);
or U242 (N_242,In_133,In_745);
nor U243 (N_243,In_147,In_305);
nand U244 (N_244,In_151,In_193);
or U245 (N_245,In_65,In_196);
and U246 (N_246,In_236,In_337);
and U247 (N_247,In_456,In_749);
nor U248 (N_248,In_484,In_100);
nor U249 (N_249,In_399,In_22);
or U250 (N_250,In_669,In_704);
and U251 (N_251,In_207,In_290);
nand U252 (N_252,In_697,In_723);
and U253 (N_253,In_364,In_251);
or U254 (N_254,In_365,In_599);
or U255 (N_255,In_183,In_510);
nand U256 (N_256,In_384,In_129);
and U257 (N_257,In_645,In_206);
and U258 (N_258,In_686,In_501);
and U259 (N_259,In_1,In_604);
or U260 (N_260,In_367,In_615);
nand U261 (N_261,In_330,In_391);
nand U262 (N_262,In_372,In_463);
and U263 (N_263,In_118,In_155);
or U264 (N_264,In_659,In_630);
or U265 (N_265,In_21,In_220);
and U266 (N_266,In_135,In_264);
and U267 (N_267,In_611,In_720);
and U268 (N_268,In_550,In_560);
and U269 (N_269,In_439,In_619);
nand U270 (N_270,In_420,In_742);
and U271 (N_271,In_16,In_111);
or U272 (N_272,In_690,In_574);
nor U273 (N_273,In_643,In_355);
or U274 (N_274,In_278,In_91);
or U275 (N_275,In_101,In_154);
or U276 (N_276,In_641,In_731);
or U277 (N_277,In_338,In_694);
nand U278 (N_278,In_573,In_711);
nand U279 (N_279,In_705,In_506);
nor U280 (N_280,In_152,In_587);
and U281 (N_281,In_639,In_710);
nand U282 (N_282,In_389,In_503);
xnor U283 (N_283,In_157,In_672);
or U284 (N_284,In_565,In_120);
nor U285 (N_285,In_566,In_575);
or U286 (N_286,In_68,In_468);
or U287 (N_287,In_228,In_490);
nor U288 (N_288,In_395,In_633);
xor U289 (N_289,In_69,In_210);
nor U290 (N_290,In_647,In_569);
nand U291 (N_291,In_655,In_408);
or U292 (N_292,In_48,In_318);
or U293 (N_293,In_179,In_593);
xnor U294 (N_294,In_26,In_613);
or U295 (N_295,In_612,In_448);
or U296 (N_296,In_83,In_585);
or U297 (N_297,In_137,In_375);
nand U298 (N_298,In_170,In_272);
xor U299 (N_299,In_504,In_46);
xnor U300 (N_300,In_102,In_209);
nor U301 (N_301,In_42,In_353);
nor U302 (N_302,In_208,In_145);
nand U303 (N_303,In_356,In_552);
xor U304 (N_304,In_267,In_415);
or U305 (N_305,In_50,In_352);
nor U306 (N_306,In_289,In_136);
nor U307 (N_307,In_648,In_60);
or U308 (N_308,In_444,In_158);
nor U309 (N_309,In_31,In_186);
nand U310 (N_310,In_534,In_382);
nor U311 (N_311,In_325,In_727);
nor U312 (N_312,In_126,In_178);
xor U313 (N_313,In_368,In_702);
or U314 (N_314,In_104,In_734);
and U315 (N_315,In_523,In_248);
and U316 (N_316,In_681,In_29);
nand U317 (N_317,In_695,In_232);
and U318 (N_318,In_53,In_275);
nand U319 (N_319,In_677,In_166);
and U320 (N_320,In_134,In_331);
or U321 (N_321,In_88,In_477);
or U322 (N_322,In_455,In_282);
nor U323 (N_323,In_252,In_406);
nand U324 (N_324,In_546,In_662);
and U325 (N_325,In_341,In_43);
nor U326 (N_326,In_588,In_658);
nor U327 (N_327,In_32,In_205);
nor U328 (N_328,In_383,In_327);
nor U329 (N_329,In_495,In_262);
and U330 (N_330,In_377,In_525);
nand U331 (N_331,In_407,In_268);
xor U332 (N_332,In_624,In_567);
nor U333 (N_333,In_0,In_30);
xor U334 (N_334,In_511,In_79);
or U335 (N_335,In_94,In_370);
or U336 (N_336,In_481,In_148);
nor U337 (N_337,In_728,In_316);
nand U338 (N_338,In_212,In_492);
or U339 (N_339,In_373,In_489);
xnor U340 (N_340,In_628,In_634);
nor U341 (N_341,In_176,In_57);
nand U342 (N_342,In_738,In_744);
and U343 (N_343,In_259,In_256);
or U344 (N_344,In_191,In_714);
nor U345 (N_345,In_11,In_105);
nor U346 (N_346,In_472,In_27);
and U347 (N_347,In_691,In_616);
nor U348 (N_348,In_512,In_540);
or U349 (N_349,In_146,In_685);
xnor U350 (N_350,In_13,In_533);
nand U351 (N_351,In_537,In_202);
and U352 (N_352,In_144,In_716);
nand U353 (N_353,In_287,In_39);
or U354 (N_354,In_549,In_660);
xor U355 (N_355,In_371,In_562);
and U356 (N_356,In_20,In_581);
nor U357 (N_357,In_307,In_306);
nor U358 (N_358,In_181,In_505);
or U359 (N_359,In_553,In_303);
or U360 (N_360,In_500,In_717);
or U361 (N_361,In_577,In_54);
nor U362 (N_362,In_488,In_557);
nand U363 (N_363,In_527,In_66);
or U364 (N_364,In_458,In_360);
nand U365 (N_365,In_404,In_652);
nor U366 (N_366,In_457,In_51);
nor U367 (N_367,In_55,In_462);
nor U368 (N_368,In_548,In_600);
and U369 (N_369,In_299,In_493);
nor U370 (N_370,In_475,In_582);
nor U371 (N_371,In_87,In_334);
nor U372 (N_372,In_273,In_114);
and U373 (N_373,In_603,In_164);
and U374 (N_374,In_350,In_343);
nand U375 (N_375,In_553,In_323);
or U376 (N_376,In_364,In_550);
nand U377 (N_377,In_52,In_688);
nand U378 (N_378,In_678,In_89);
and U379 (N_379,In_667,In_347);
and U380 (N_380,In_133,In_705);
or U381 (N_381,In_615,In_412);
nand U382 (N_382,In_459,In_493);
or U383 (N_383,In_339,In_557);
nor U384 (N_384,In_102,In_94);
and U385 (N_385,In_623,In_418);
and U386 (N_386,In_44,In_79);
or U387 (N_387,In_595,In_290);
xnor U388 (N_388,In_374,In_106);
nor U389 (N_389,In_199,In_677);
nand U390 (N_390,In_266,In_605);
and U391 (N_391,In_629,In_626);
or U392 (N_392,In_501,In_0);
xnor U393 (N_393,In_717,In_152);
nor U394 (N_394,In_669,In_471);
or U395 (N_395,In_537,In_408);
or U396 (N_396,In_547,In_41);
nor U397 (N_397,In_192,In_640);
nand U398 (N_398,In_362,In_162);
and U399 (N_399,In_685,In_80);
and U400 (N_400,In_254,In_566);
xnor U401 (N_401,In_610,In_261);
and U402 (N_402,In_299,In_110);
or U403 (N_403,In_143,In_50);
and U404 (N_404,In_20,In_162);
nand U405 (N_405,In_128,In_589);
nor U406 (N_406,In_366,In_339);
and U407 (N_407,In_551,In_325);
and U408 (N_408,In_6,In_543);
nand U409 (N_409,In_332,In_65);
and U410 (N_410,In_513,In_481);
and U411 (N_411,In_608,In_596);
nand U412 (N_412,In_390,In_247);
or U413 (N_413,In_481,In_693);
or U414 (N_414,In_42,In_332);
nor U415 (N_415,In_30,In_204);
and U416 (N_416,In_98,In_713);
xnor U417 (N_417,In_306,In_216);
nor U418 (N_418,In_575,In_256);
xor U419 (N_419,In_733,In_70);
or U420 (N_420,In_35,In_93);
and U421 (N_421,In_63,In_59);
nor U422 (N_422,In_72,In_354);
nand U423 (N_423,In_679,In_729);
or U424 (N_424,In_487,In_240);
and U425 (N_425,In_338,In_672);
nor U426 (N_426,In_583,In_118);
nand U427 (N_427,In_91,In_556);
or U428 (N_428,In_474,In_538);
nand U429 (N_429,In_742,In_428);
and U430 (N_430,In_219,In_310);
nor U431 (N_431,In_120,In_562);
nor U432 (N_432,In_286,In_190);
nand U433 (N_433,In_688,In_650);
nand U434 (N_434,In_517,In_362);
nor U435 (N_435,In_353,In_579);
nor U436 (N_436,In_213,In_34);
xor U437 (N_437,In_617,In_687);
nand U438 (N_438,In_397,In_165);
or U439 (N_439,In_141,In_659);
or U440 (N_440,In_402,In_367);
nand U441 (N_441,In_387,In_200);
or U442 (N_442,In_276,In_161);
and U443 (N_443,In_189,In_233);
nor U444 (N_444,In_457,In_37);
and U445 (N_445,In_569,In_79);
xor U446 (N_446,In_621,In_209);
and U447 (N_447,In_235,In_89);
nand U448 (N_448,In_258,In_590);
or U449 (N_449,In_299,In_178);
and U450 (N_450,In_416,In_26);
or U451 (N_451,In_600,In_61);
or U452 (N_452,In_604,In_192);
or U453 (N_453,In_16,In_533);
nor U454 (N_454,In_143,In_234);
nand U455 (N_455,In_351,In_392);
nor U456 (N_456,In_422,In_357);
or U457 (N_457,In_657,In_712);
nor U458 (N_458,In_547,In_272);
or U459 (N_459,In_280,In_106);
and U460 (N_460,In_327,In_725);
and U461 (N_461,In_717,In_587);
or U462 (N_462,In_696,In_17);
and U463 (N_463,In_534,In_651);
nor U464 (N_464,In_290,In_461);
nand U465 (N_465,In_327,In_397);
or U466 (N_466,In_210,In_458);
and U467 (N_467,In_649,In_676);
nor U468 (N_468,In_10,In_235);
nor U469 (N_469,In_44,In_399);
nand U470 (N_470,In_512,In_253);
nand U471 (N_471,In_56,In_496);
nor U472 (N_472,In_14,In_87);
nand U473 (N_473,In_741,In_386);
nor U474 (N_474,In_346,In_456);
nand U475 (N_475,In_677,In_60);
nor U476 (N_476,In_6,In_84);
nor U477 (N_477,In_259,In_242);
or U478 (N_478,In_2,In_671);
nor U479 (N_479,In_598,In_148);
nor U480 (N_480,In_643,In_35);
and U481 (N_481,In_315,In_104);
nand U482 (N_482,In_217,In_234);
nand U483 (N_483,In_600,In_314);
nor U484 (N_484,In_363,In_153);
and U485 (N_485,In_45,In_104);
and U486 (N_486,In_461,In_428);
and U487 (N_487,In_554,In_632);
xor U488 (N_488,In_284,In_34);
and U489 (N_489,In_220,In_528);
or U490 (N_490,In_123,In_572);
nand U491 (N_491,In_125,In_284);
nor U492 (N_492,In_660,In_668);
and U493 (N_493,In_655,In_743);
xnor U494 (N_494,In_569,In_6);
nand U495 (N_495,In_513,In_610);
nand U496 (N_496,In_749,In_70);
nor U497 (N_497,In_585,In_457);
and U498 (N_498,In_118,In_157);
nand U499 (N_499,In_63,In_451);
nand U500 (N_500,In_493,In_309);
or U501 (N_501,In_172,In_102);
nand U502 (N_502,In_250,In_266);
or U503 (N_503,In_129,In_662);
or U504 (N_504,In_548,In_730);
and U505 (N_505,In_735,In_170);
nand U506 (N_506,In_549,In_425);
and U507 (N_507,In_693,In_315);
nor U508 (N_508,In_492,In_173);
nor U509 (N_509,In_600,In_6);
xnor U510 (N_510,In_522,In_235);
and U511 (N_511,In_402,In_228);
or U512 (N_512,In_603,In_503);
nor U513 (N_513,In_582,In_708);
nor U514 (N_514,In_404,In_723);
nand U515 (N_515,In_403,In_714);
and U516 (N_516,In_470,In_701);
and U517 (N_517,In_744,In_638);
and U518 (N_518,In_463,In_279);
nor U519 (N_519,In_572,In_334);
nor U520 (N_520,In_215,In_8);
or U521 (N_521,In_198,In_260);
or U522 (N_522,In_501,In_169);
nand U523 (N_523,In_453,In_710);
and U524 (N_524,In_499,In_337);
xnor U525 (N_525,In_442,In_10);
or U526 (N_526,In_404,In_372);
nand U527 (N_527,In_395,In_224);
nor U528 (N_528,In_371,In_608);
or U529 (N_529,In_288,In_358);
or U530 (N_530,In_667,In_688);
nand U531 (N_531,In_205,In_584);
and U532 (N_532,In_284,In_93);
nor U533 (N_533,In_141,In_538);
nand U534 (N_534,In_181,In_709);
or U535 (N_535,In_618,In_149);
nor U536 (N_536,In_8,In_267);
and U537 (N_537,In_246,In_548);
nor U538 (N_538,In_691,In_27);
and U539 (N_539,In_632,In_204);
nand U540 (N_540,In_324,In_198);
or U541 (N_541,In_286,In_604);
nand U542 (N_542,In_703,In_181);
nand U543 (N_543,In_108,In_402);
nand U544 (N_544,In_627,In_224);
or U545 (N_545,In_441,In_319);
or U546 (N_546,In_492,In_245);
and U547 (N_547,In_33,In_706);
and U548 (N_548,In_665,In_14);
nor U549 (N_549,In_366,In_235);
nand U550 (N_550,In_104,In_428);
nand U551 (N_551,In_182,In_144);
or U552 (N_552,In_40,In_312);
and U553 (N_553,In_213,In_743);
nor U554 (N_554,In_81,In_140);
nand U555 (N_555,In_668,In_146);
or U556 (N_556,In_712,In_698);
and U557 (N_557,In_70,In_687);
or U558 (N_558,In_561,In_74);
nor U559 (N_559,In_285,In_373);
and U560 (N_560,In_718,In_216);
nand U561 (N_561,In_448,In_748);
nand U562 (N_562,In_638,In_553);
or U563 (N_563,In_310,In_417);
nand U564 (N_564,In_618,In_598);
and U565 (N_565,In_210,In_453);
and U566 (N_566,In_524,In_207);
or U567 (N_567,In_467,In_71);
and U568 (N_568,In_125,In_616);
xnor U569 (N_569,In_167,In_740);
nor U570 (N_570,In_667,In_517);
nor U571 (N_571,In_649,In_239);
nor U572 (N_572,In_171,In_60);
nand U573 (N_573,In_248,In_146);
and U574 (N_574,In_232,In_710);
or U575 (N_575,In_372,In_91);
xnor U576 (N_576,In_181,In_521);
or U577 (N_577,In_59,In_43);
or U578 (N_578,In_67,In_677);
xnor U579 (N_579,In_89,In_337);
and U580 (N_580,In_626,In_458);
nor U581 (N_581,In_24,In_330);
or U582 (N_582,In_113,In_3);
and U583 (N_583,In_503,In_0);
or U584 (N_584,In_19,In_260);
and U585 (N_585,In_30,In_735);
nor U586 (N_586,In_457,In_170);
and U587 (N_587,In_642,In_242);
or U588 (N_588,In_640,In_180);
nand U589 (N_589,In_556,In_31);
nor U590 (N_590,In_302,In_37);
nor U591 (N_591,In_26,In_79);
nand U592 (N_592,In_613,In_22);
nand U593 (N_593,In_60,In_74);
and U594 (N_594,In_46,In_346);
nand U595 (N_595,In_346,In_336);
and U596 (N_596,In_413,In_272);
or U597 (N_597,In_649,In_14);
nor U598 (N_598,In_247,In_200);
nand U599 (N_599,In_626,In_686);
or U600 (N_600,In_389,In_361);
or U601 (N_601,In_243,In_389);
or U602 (N_602,In_488,In_622);
nand U603 (N_603,In_1,In_329);
and U604 (N_604,In_244,In_436);
or U605 (N_605,In_208,In_275);
and U606 (N_606,In_690,In_656);
nor U607 (N_607,In_423,In_5);
nor U608 (N_608,In_556,In_645);
nor U609 (N_609,In_210,In_252);
nand U610 (N_610,In_260,In_152);
nand U611 (N_611,In_505,In_508);
nand U612 (N_612,In_109,In_123);
nand U613 (N_613,In_467,In_679);
nand U614 (N_614,In_353,In_653);
nand U615 (N_615,In_332,In_425);
or U616 (N_616,In_605,In_52);
and U617 (N_617,In_581,In_125);
xnor U618 (N_618,In_96,In_152);
or U619 (N_619,In_355,In_748);
and U620 (N_620,In_3,In_65);
or U621 (N_621,In_551,In_361);
nand U622 (N_622,In_481,In_572);
nand U623 (N_623,In_394,In_399);
nor U624 (N_624,In_310,In_633);
nor U625 (N_625,In_179,In_704);
nor U626 (N_626,In_151,In_517);
or U627 (N_627,In_513,In_696);
and U628 (N_628,In_213,In_81);
nor U629 (N_629,In_532,In_98);
and U630 (N_630,In_128,In_557);
and U631 (N_631,In_536,In_118);
or U632 (N_632,In_679,In_701);
and U633 (N_633,In_648,In_702);
nand U634 (N_634,In_182,In_489);
and U635 (N_635,In_405,In_114);
or U636 (N_636,In_414,In_697);
or U637 (N_637,In_265,In_398);
and U638 (N_638,In_494,In_604);
nand U639 (N_639,In_86,In_28);
nand U640 (N_640,In_360,In_402);
and U641 (N_641,In_683,In_342);
nor U642 (N_642,In_4,In_520);
nor U643 (N_643,In_437,In_504);
xnor U644 (N_644,In_514,In_343);
nand U645 (N_645,In_342,In_702);
and U646 (N_646,In_455,In_218);
or U647 (N_647,In_518,In_123);
xor U648 (N_648,In_592,In_96);
nand U649 (N_649,In_546,In_130);
or U650 (N_650,In_420,In_186);
or U651 (N_651,In_663,In_522);
nor U652 (N_652,In_567,In_75);
or U653 (N_653,In_97,In_618);
xor U654 (N_654,In_532,In_531);
nand U655 (N_655,In_483,In_263);
and U656 (N_656,In_351,In_630);
or U657 (N_657,In_100,In_168);
and U658 (N_658,In_178,In_511);
and U659 (N_659,In_277,In_388);
and U660 (N_660,In_31,In_165);
and U661 (N_661,In_199,In_651);
and U662 (N_662,In_144,In_14);
or U663 (N_663,In_453,In_549);
nand U664 (N_664,In_264,In_745);
nand U665 (N_665,In_429,In_692);
and U666 (N_666,In_513,In_360);
xor U667 (N_667,In_269,In_246);
nor U668 (N_668,In_678,In_721);
or U669 (N_669,In_40,In_508);
and U670 (N_670,In_474,In_64);
or U671 (N_671,In_498,In_733);
nand U672 (N_672,In_92,In_234);
nor U673 (N_673,In_262,In_287);
or U674 (N_674,In_321,In_555);
and U675 (N_675,In_316,In_218);
and U676 (N_676,In_515,In_411);
nor U677 (N_677,In_503,In_735);
or U678 (N_678,In_84,In_520);
and U679 (N_679,In_314,In_5);
nor U680 (N_680,In_365,In_433);
nor U681 (N_681,In_653,In_0);
and U682 (N_682,In_413,In_670);
and U683 (N_683,In_401,In_240);
nand U684 (N_684,In_363,In_737);
nand U685 (N_685,In_177,In_677);
or U686 (N_686,In_56,In_355);
nand U687 (N_687,In_745,In_408);
or U688 (N_688,In_322,In_633);
nor U689 (N_689,In_189,In_724);
nand U690 (N_690,In_359,In_350);
nand U691 (N_691,In_599,In_185);
and U692 (N_692,In_309,In_89);
or U693 (N_693,In_327,In_530);
nor U694 (N_694,In_200,In_439);
nor U695 (N_695,In_57,In_548);
nor U696 (N_696,In_415,In_538);
nor U697 (N_697,In_199,In_492);
or U698 (N_698,In_654,In_476);
nand U699 (N_699,In_40,In_116);
nand U700 (N_700,In_361,In_305);
and U701 (N_701,In_274,In_268);
nor U702 (N_702,In_697,In_675);
nand U703 (N_703,In_748,In_613);
and U704 (N_704,In_102,In_682);
xnor U705 (N_705,In_263,In_333);
or U706 (N_706,In_67,In_223);
nor U707 (N_707,In_224,In_443);
nor U708 (N_708,In_662,In_291);
and U709 (N_709,In_186,In_639);
nand U710 (N_710,In_25,In_460);
nand U711 (N_711,In_35,In_198);
and U712 (N_712,In_516,In_216);
and U713 (N_713,In_267,In_370);
xor U714 (N_714,In_620,In_173);
and U715 (N_715,In_69,In_458);
xnor U716 (N_716,In_339,In_674);
nor U717 (N_717,In_38,In_434);
nand U718 (N_718,In_637,In_533);
nor U719 (N_719,In_83,In_45);
nor U720 (N_720,In_435,In_224);
or U721 (N_721,In_667,In_294);
or U722 (N_722,In_585,In_313);
xnor U723 (N_723,In_76,In_196);
or U724 (N_724,In_269,In_166);
or U725 (N_725,In_486,In_590);
or U726 (N_726,In_109,In_244);
nand U727 (N_727,In_287,In_206);
and U728 (N_728,In_509,In_270);
nand U729 (N_729,In_392,In_111);
nor U730 (N_730,In_504,In_546);
nand U731 (N_731,In_374,In_390);
or U732 (N_732,In_470,In_672);
and U733 (N_733,In_89,In_25);
and U734 (N_734,In_490,In_378);
nand U735 (N_735,In_591,In_277);
nor U736 (N_736,In_297,In_166);
and U737 (N_737,In_283,In_681);
nand U738 (N_738,In_21,In_739);
xnor U739 (N_739,In_278,In_433);
and U740 (N_740,In_37,In_384);
and U741 (N_741,In_520,In_17);
or U742 (N_742,In_477,In_73);
and U743 (N_743,In_632,In_478);
or U744 (N_744,In_412,In_324);
nand U745 (N_745,In_410,In_247);
nand U746 (N_746,In_484,In_224);
or U747 (N_747,In_44,In_492);
nor U748 (N_748,In_467,In_672);
nand U749 (N_749,In_612,In_171);
nand U750 (N_750,In_624,In_389);
nor U751 (N_751,In_627,In_591);
xor U752 (N_752,In_127,In_691);
nor U753 (N_753,In_553,In_1);
or U754 (N_754,In_284,In_375);
and U755 (N_755,In_98,In_197);
nand U756 (N_756,In_269,In_390);
xnor U757 (N_757,In_616,In_295);
nor U758 (N_758,In_197,In_208);
and U759 (N_759,In_682,In_217);
and U760 (N_760,In_304,In_514);
and U761 (N_761,In_515,In_83);
and U762 (N_762,In_706,In_169);
and U763 (N_763,In_186,In_190);
or U764 (N_764,In_518,In_113);
nand U765 (N_765,In_618,In_360);
nand U766 (N_766,In_53,In_248);
xnor U767 (N_767,In_76,In_703);
nor U768 (N_768,In_382,In_309);
and U769 (N_769,In_668,In_243);
or U770 (N_770,In_719,In_655);
and U771 (N_771,In_48,In_205);
xnor U772 (N_772,In_188,In_190);
and U773 (N_773,In_591,In_110);
nand U774 (N_774,In_672,In_86);
nand U775 (N_775,In_39,In_328);
and U776 (N_776,In_715,In_325);
nand U777 (N_777,In_604,In_606);
xnor U778 (N_778,In_649,In_687);
or U779 (N_779,In_563,In_35);
xor U780 (N_780,In_678,In_598);
nand U781 (N_781,In_332,In_339);
nand U782 (N_782,In_570,In_384);
nor U783 (N_783,In_555,In_430);
or U784 (N_784,In_496,In_621);
or U785 (N_785,In_322,In_320);
or U786 (N_786,In_673,In_348);
nor U787 (N_787,In_484,In_246);
nand U788 (N_788,In_654,In_456);
nand U789 (N_789,In_694,In_622);
nor U790 (N_790,In_137,In_433);
and U791 (N_791,In_215,In_559);
nand U792 (N_792,In_393,In_585);
and U793 (N_793,In_258,In_27);
nand U794 (N_794,In_131,In_561);
or U795 (N_795,In_588,In_181);
or U796 (N_796,In_150,In_388);
nand U797 (N_797,In_614,In_731);
and U798 (N_798,In_746,In_550);
or U799 (N_799,In_450,In_407);
nand U800 (N_800,In_550,In_370);
and U801 (N_801,In_635,In_496);
nor U802 (N_802,In_348,In_430);
nand U803 (N_803,In_375,In_94);
or U804 (N_804,In_114,In_103);
nor U805 (N_805,In_108,In_284);
xor U806 (N_806,In_313,In_424);
and U807 (N_807,In_717,In_746);
nor U808 (N_808,In_711,In_168);
nand U809 (N_809,In_746,In_286);
and U810 (N_810,In_598,In_396);
and U811 (N_811,In_224,In_103);
and U812 (N_812,In_105,In_619);
and U813 (N_813,In_648,In_164);
nor U814 (N_814,In_560,In_269);
xor U815 (N_815,In_90,In_326);
nand U816 (N_816,In_466,In_164);
xnor U817 (N_817,In_49,In_1);
nor U818 (N_818,In_452,In_503);
and U819 (N_819,In_206,In_470);
and U820 (N_820,In_680,In_20);
nand U821 (N_821,In_474,In_601);
nor U822 (N_822,In_502,In_224);
and U823 (N_823,In_633,In_355);
or U824 (N_824,In_19,In_737);
nor U825 (N_825,In_117,In_561);
nor U826 (N_826,In_264,In_438);
nand U827 (N_827,In_425,In_17);
xor U828 (N_828,In_659,In_638);
or U829 (N_829,In_279,In_439);
or U830 (N_830,In_419,In_6);
nor U831 (N_831,In_535,In_47);
nand U832 (N_832,In_317,In_409);
nor U833 (N_833,In_233,In_320);
nand U834 (N_834,In_624,In_299);
nor U835 (N_835,In_2,In_108);
nor U836 (N_836,In_357,In_311);
xor U837 (N_837,In_243,In_667);
nand U838 (N_838,In_537,In_261);
nor U839 (N_839,In_142,In_580);
or U840 (N_840,In_234,In_580);
or U841 (N_841,In_689,In_162);
and U842 (N_842,In_62,In_400);
xnor U843 (N_843,In_587,In_209);
and U844 (N_844,In_474,In_218);
nor U845 (N_845,In_469,In_256);
xor U846 (N_846,In_22,In_663);
nand U847 (N_847,In_247,In_224);
nand U848 (N_848,In_378,In_34);
xnor U849 (N_849,In_626,In_663);
nand U850 (N_850,In_369,In_590);
or U851 (N_851,In_357,In_736);
and U852 (N_852,In_681,In_345);
nand U853 (N_853,In_641,In_195);
xnor U854 (N_854,In_541,In_511);
xnor U855 (N_855,In_538,In_682);
or U856 (N_856,In_219,In_164);
or U857 (N_857,In_669,In_210);
or U858 (N_858,In_734,In_155);
and U859 (N_859,In_379,In_190);
xnor U860 (N_860,In_40,In_381);
or U861 (N_861,In_509,In_555);
nand U862 (N_862,In_383,In_146);
nand U863 (N_863,In_526,In_212);
nand U864 (N_864,In_132,In_122);
or U865 (N_865,In_498,In_654);
or U866 (N_866,In_417,In_467);
or U867 (N_867,In_360,In_124);
nand U868 (N_868,In_390,In_403);
nand U869 (N_869,In_303,In_682);
or U870 (N_870,In_130,In_731);
or U871 (N_871,In_183,In_154);
nand U872 (N_872,In_283,In_675);
and U873 (N_873,In_319,In_12);
or U874 (N_874,In_719,In_730);
or U875 (N_875,In_577,In_352);
nor U876 (N_876,In_103,In_678);
and U877 (N_877,In_389,In_491);
nor U878 (N_878,In_68,In_410);
and U879 (N_879,In_619,In_154);
nor U880 (N_880,In_308,In_40);
nand U881 (N_881,In_163,In_718);
and U882 (N_882,In_56,In_28);
nor U883 (N_883,In_383,In_216);
or U884 (N_884,In_705,In_647);
xor U885 (N_885,In_75,In_152);
and U886 (N_886,In_673,In_138);
or U887 (N_887,In_195,In_68);
nand U888 (N_888,In_228,In_412);
or U889 (N_889,In_690,In_539);
or U890 (N_890,In_631,In_398);
xnor U891 (N_891,In_457,In_32);
nand U892 (N_892,In_191,In_672);
nand U893 (N_893,In_415,In_83);
nand U894 (N_894,In_398,In_374);
nor U895 (N_895,In_737,In_620);
nor U896 (N_896,In_585,In_643);
and U897 (N_897,In_447,In_538);
nor U898 (N_898,In_410,In_541);
nor U899 (N_899,In_87,In_715);
and U900 (N_900,In_617,In_44);
and U901 (N_901,In_349,In_743);
nor U902 (N_902,In_499,In_33);
or U903 (N_903,In_112,In_381);
nor U904 (N_904,In_712,In_62);
nand U905 (N_905,In_429,In_563);
nor U906 (N_906,In_180,In_298);
xor U907 (N_907,In_255,In_210);
nand U908 (N_908,In_141,In_275);
nor U909 (N_909,In_304,In_120);
nand U910 (N_910,In_338,In_359);
nand U911 (N_911,In_146,In_597);
or U912 (N_912,In_149,In_445);
nand U913 (N_913,In_464,In_49);
nor U914 (N_914,In_139,In_338);
or U915 (N_915,In_295,In_391);
and U916 (N_916,In_68,In_145);
nand U917 (N_917,In_347,In_460);
xnor U918 (N_918,In_241,In_740);
nand U919 (N_919,In_317,In_165);
and U920 (N_920,In_518,In_377);
nor U921 (N_921,In_713,In_575);
or U922 (N_922,In_207,In_497);
xor U923 (N_923,In_401,In_226);
or U924 (N_924,In_715,In_712);
nand U925 (N_925,In_240,In_522);
nor U926 (N_926,In_737,In_491);
and U927 (N_927,In_604,In_599);
or U928 (N_928,In_125,In_184);
and U929 (N_929,In_647,In_197);
or U930 (N_930,In_92,In_619);
xor U931 (N_931,In_267,In_312);
or U932 (N_932,In_460,In_115);
or U933 (N_933,In_317,In_618);
or U934 (N_934,In_730,In_18);
and U935 (N_935,In_654,In_108);
or U936 (N_936,In_470,In_152);
nand U937 (N_937,In_543,In_157);
xnor U938 (N_938,In_53,In_254);
and U939 (N_939,In_246,In_270);
nand U940 (N_940,In_240,In_708);
nand U941 (N_941,In_598,In_345);
nand U942 (N_942,In_17,In_412);
or U943 (N_943,In_648,In_508);
nor U944 (N_944,In_678,In_43);
xnor U945 (N_945,In_678,In_297);
and U946 (N_946,In_525,In_318);
nor U947 (N_947,In_71,In_657);
and U948 (N_948,In_541,In_39);
nor U949 (N_949,In_500,In_666);
nand U950 (N_950,In_288,In_230);
nand U951 (N_951,In_661,In_592);
or U952 (N_952,In_165,In_94);
or U953 (N_953,In_390,In_283);
nand U954 (N_954,In_278,In_293);
nor U955 (N_955,In_123,In_136);
or U956 (N_956,In_157,In_302);
nor U957 (N_957,In_590,In_723);
nor U958 (N_958,In_228,In_746);
or U959 (N_959,In_82,In_47);
and U960 (N_960,In_13,In_707);
nor U961 (N_961,In_132,In_72);
nor U962 (N_962,In_361,In_132);
nand U963 (N_963,In_738,In_357);
or U964 (N_964,In_175,In_540);
and U965 (N_965,In_70,In_301);
and U966 (N_966,In_29,In_339);
nor U967 (N_967,In_531,In_614);
and U968 (N_968,In_45,In_186);
nor U969 (N_969,In_374,In_178);
and U970 (N_970,In_737,In_584);
or U971 (N_971,In_341,In_261);
nand U972 (N_972,In_302,In_405);
nor U973 (N_973,In_403,In_658);
nand U974 (N_974,In_635,In_34);
and U975 (N_975,In_55,In_327);
nand U976 (N_976,In_588,In_480);
xor U977 (N_977,In_511,In_654);
nor U978 (N_978,In_726,In_138);
or U979 (N_979,In_140,In_68);
nand U980 (N_980,In_389,In_482);
nand U981 (N_981,In_365,In_109);
and U982 (N_982,In_42,In_179);
xor U983 (N_983,In_438,In_540);
nand U984 (N_984,In_474,In_34);
nor U985 (N_985,In_670,In_726);
nor U986 (N_986,In_511,In_217);
xor U987 (N_987,In_691,In_487);
or U988 (N_988,In_544,In_467);
and U989 (N_989,In_450,In_476);
xnor U990 (N_990,In_747,In_46);
nor U991 (N_991,In_550,In_318);
or U992 (N_992,In_538,In_239);
or U993 (N_993,In_255,In_96);
xor U994 (N_994,In_679,In_629);
or U995 (N_995,In_209,In_96);
nor U996 (N_996,In_106,In_176);
or U997 (N_997,In_501,In_728);
and U998 (N_998,In_28,In_242);
nand U999 (N_999,In_457,In_563);
nor U1000 (N_1000,N_913,N_909);
xnor U1001 (N_1001,N_619,N_56);
nand U1002 (N_1002,N_60,N_222);
xnor U1003 (N_1003,N_151,N_706);
nor U1004 (N_1004,N_745,N_639);
and U1005 (N_1005,N_699,N_38);
nand U1006 (N_1006,N_622,N_727);
nand U1007 (N_1007,N_442,N_251);
nand U1008 (N_1008,N_968,N_778);
and U1009 (N_1009,N_363,N_184);
or U1010 (N_1010,N_289,N_101);
and U1011 (N_1011,N_32,N_624);
nor U1012 (N_1012,N_634,N_200);
and U1013 (N_1013,N_541,N_29);
and U1014 (N_1014,N_237,N_343);
xnor U1015 (N_1015,N_938,N_471);
or U1016 (N_1016,N_886,N_589);
xnor U1017 (N_1017,N_862,N_204);
or U1018 (N_1018,N_721,N_24);
nor U1019 (N_1019,N_605,N_796);
nand U1020 (N_1020,N_395,N_677);
nand U1021 (N_1021,N_493,N_660);
xnor U1022 (N_1022,N_537,N_689);
and U1023 (N_1023,N_974,N_997);
nor U1024 (N_1024,N_335,N_275);
nor U1025 (N_1025,N_262,N_172);
and U1026 (N_1026,N_636,N_318);
nor U1027 (N_1027,N_531,N_765);
or U1028 (N_1028,N_181,N_146);
nor U1029 (N_1029,N_351,N_517);
or U1030 (N_1030,N_243,N_413);
xnor U1031 (N_1031,N_91,N_818);
and U1032 (N_1032,N_231,N_789);
nor U1033 (N_1033,N_255,N_452);
or U1034 (N_1034,N_337,N_885);
nor U1035 (N_1035,N_577,N_540);
and U1036 (N_1036,N_404,N_238);
or U1037 (N_1037,N_871,N_903);
or U1038 (N_1038,N_529,N_406);
nand U1039 (N_1039,N_436,N_908);
or U1040 (N_1040,N_368,N_787);
nand U1041 (N_1041,N_614,N_739);
nor U1042 (N_1042,N_393,N_349);
xnor U1043 (N_1043,N_941,N_336);
or U1044 (N_1044,N_595,N_365);
and U1045 (N_1045,N_379,N_784);
and U1046 (N_1046,N_836,N_8);
nand U1047 (N_1047,N_266,N_165);
and U1048 (N_1048,N_302,N_800);
nand U1049 (N_1049,N_664,N_82);
xnor U1050 (N_1050,N_196,N_117);
nor U1051 (N_1051,N_408,N_307);
and U1052 (N_1052,N_297,N_369);
nor U1053 (N_1053,N_681,N_444);
nand U1054 (N_1054,N_330,N_194);
nor U1055 (N_1055,N_767,N_338);
nor U1056 (N_1056,N_135,N_348);
nor U1057 (N_1057,N_278,N_157);
and U1058 (N_1058,N_575,N_567);
xor U1059 (N_1059,N_928,N_661);
or U1060 (N_1060,N_17,N_362);
or U1061 (N_1061,N_392,N_848);
nor U1062 (N_1062,N_870,N_596);
nor U1063 (N_1063,N_426,N_169);
or U1064 (N_1064,N_560,N_586);
nand U1065 (N_1065,N_667,N_371);
nor U1066 (N_1066,N_116,N_785);
nor U1067 (N_1067,N_829,N_858);
and U1068 (N_1068,N_579,N_118);
nor U1069 (N_1069,N_719,N_613);
and U1070 (N_1070,N_90,N_949);
or U1071 (N_1071,N_300,N_821);
nand U1072 (N_1072,N_924,N_731);
and U1073 (N_1073,N_378,N_84);
and U1074 (N_1074,N_1,N_290);
or U1075 (N_1075,N_475,N_612);
nand U1076 (N_1076,N_156,N_602);
nand U1077 (N_1077,N_0,N_686);
and U1078 (N_1078,N_902,N_367);
nor U1079 (N_1079,N_547,N_31);
and U1080 (N_1080,N_995,N_876);
or U1081 (N_1081,N_69,N_357);
or U1082 (N_1082,N_621,N_158);
and U1083 (N_1083,N_234,N_269);
nand U1084 (N_1084,N_865,N_833);
nand U1085 (N_1085,N_897,N_466);
or U1086 (N_1086,N_482,N_512);
and U1087 (N_1087,N_143,N_199);
or U1088 (N_1088,N_80,N_182);
or U1089 (N_1089,N_376,N_201);
and U1090 (N_1090,N_542,N_643);
nand U1091 (N_1091,N_180,N_525);
or U1092 (N_1092,N_5,N_259);
and U1093 (N_1093,N_301,N_810);
or U1094 (N_1094,N_286,N_45);
and U1095 (N_1095,N_528,N_861);
or U1096 (N_1096,N_191,N_421);
nand U1097 (N_1097,N_7,N_54);
or U1098 (N_1098,N_957,N_98);
or U1099 (N_1099,N_919,N_630);
nand U1100 (N_1100,N_933,N_625);
xnor U1101 (N_1101,N_744,N_457);
or U1102 (N_1102,N_795,N_960);
and U1103 (N_1103,N_561,N_685);
nand U1104 (N_1104,N_854,N_332);
nor U1105 (N_1105,N_455,N_202);
nand U1106 (N_1106,N_61,N_986);
nor U1107 (N_1107,N_57,N_543);
nand U1108 (N_1108,N_533,N_164);
or U1109 (N_1109,N_14,N_887);
nor U1110 (N_1110,N_137,N_971);
nor U1111 (N_1111,N_414,N_948);
nand U1112 (N_1112,N_170,N_581);
nand U1113 (N_1113,N_92,N_284);
and U1114 (N_1114,N_983,N_68);
xor U1115 (N_1115,N_174,N_9);
nor U1116 (N_1116,N_979,N_709);
or U1117 (N_1117,N_945,N_272);
and U1118 (N_1118,N_549,N_808);
or U1119 (N_1119,N_217,N_279);
nand U1120 (N_1120,N_726,N_776);
or U1121 (N_1121,N_891,N_568);
xor U1122 (N_1122,N_947,N_768);
and U1123 (N_1123,N_959,N_698);
or U1124 (N_1124,N_915,N_49);
or U1125 (N_1125,N_304,N_884);
and U1126 (N_1126,N_823,N_213);
nand U1127 (N_1127,N_877,N_741);
nand U1128 (N_1128,N_822,N_433);
and U1129 (N_1129,N_780,N_690);
and U1130 (N_1130,N_831,N_964);
nand U1131 (N_1131,N_694,N_749);
nor U1132 (N_1132,N_400,N_782);
nand U1133 (N_1133,N_611,N_773);
and U1134 (N_1134,N_696,N_669);
xor U1135 (N_1135,N_256,N_626);
nand U1136 (N_1136,N_849,N_50);
xor U1137 (N_1137,N_292,N_935);
nor U1138 (N_1138,N_880,N_932);
nand U1139 (N_1139,N_334,N_942);
or U1140 (N_1140,N_448,N_769);
and U1141 (N_1141,N_429,N_454);
or U1142 (N_1142,N_930,N_852);
xnor U1143 (N_1143,N_963,N_546);
nor U1144 (N_1144,N_265,N_844);
xor U1145 (N_1145,N_663,N_791);
xnor U1146 (N_1146,N_710,N_853);
and U1147 (N_1147,N_261,N_381);
and U1148 (N_1148,N_513,N_820);
xor U1149 (N_1149,N_480,N_564);
or U1150 (N_1150,N_270,N_972);
nand U1151 (N_1151,N_779,N_310);
and U1152 (N_1152,N_940,N_962);
or U1153 (N_1153,N_592,N_651);
nor U1154 (N_1154,N_377,N_642);
xor U1155 (N_1155,N_520,N_641);
or U1156 (N_1156,N_841,N_329);
xnor U1157 (N_1157,N_764,N_133);
and U1158 (N_1158,N_760,N_670);
nor U1159 (N_1159,N_497,N_139);
nor U1160 (N_1160,N_927,N_42);
nand U1161 (N_1161,N_285,N_490);
nor U1162 (N_1162,N_834,N_427);
xnor U1163 (N_1163,N_460,N_94);
nor U1164 (N_1164,N_811,N_389);
nor U1165 (N_1165,N_291,N_4);
nor U1166 (N_1166,N_922,N_314);
or U1167 (N_1167,N_30,N_345);
or U1168 (N_1168,N_572,N_762);
nand U1169 (N_1169,N_804,N_28);
nor U1170 (N_1170,N_197,N_226);
nor U1171 (N_1171,N_210,N_701);
nand U1172 (N_1172,N_505,N_140);
and U1173 (N_1173,N_481,N_929);
nor U1174 (N_1174,N_840,N_236);
xnor U1175 (N_1175,N_206,N_125);
nor U1176 (N_1176,N_35,N_874);
and U1177 (N_1177,N_847,N_273);
and U1178 (N_1178,N_341,N_346);
nor U1179 (N_1179,N_325,N_958);
or U1180 (N_1180,N_674,N_216);
nand U1181 (N_1181,N_716,N_43);
nor U1182 (N_1182,N_228,N_248);
and U1183 (N_1183,N_323,N_123);
nand U1184 (N_1184,N_652,N_827);
nor U1185 (N_1185,N_729,N_737);
and U1186 (N_1186,N_707,N_714);
nand U1187 (N_1187,N_772,N_514);
nor U1188 (N_1188,N_851,N_85);
nor U1189 (N_1189,N_387,N_649);
or U1190 (N_1190,N_750,N_249);
and U1191 (N_1191,N_824,N_551);
or U1192 (N_1192,N_501,N_11);
and U1193 (N_1193,N_524,N_743);
or U1194 (N_1194,N_188,N_440);
nor U1195 (N_1195,N_280,N_676);
and U1196 (N_1196,N_458,N_89);
nand U1197 (N_1197,N_583,N_794);
and U1198 (N_1198,N_423,N_921);
and U1199 (N_1199,N_244,N_905);
and U1200 (N_1200,N_679,N_488);
nand U1201 (N_1201,N_618,N_678);
or U1202 (N_1202,N_430,N_771);
and U1203 (N_1203,N_189,N_288);
or U1204 (N_1204,N_609,N_766);
xor U1205 (N_1205,N_671,N_246);
nor U1206 (N_1206,N_186,N_746);
and U1207 (N_1207,N_81,N_584);
and U1208 (N_1208,N_889,N_580);
nand U1209 (N_1209,N_263,N_364);
nor U1210 (N_1210,N_461,N_386);
and U1211 (N_1211,N_814,N_375);
xnor U1212 (N_1212,N_845,N_692);
or U1213 (N_1213,N_370,N_797);
xor U1214 (N_1214,N_372,N_405);
and U1215 (N_1215,N_629,N_893);
nand U1216 (N_1216,N_985,N_920);
and U1217 (N_1217,N_813,N_740);
or U1218 (N_1218,N_224,N_937);
nor U1219 (N_1219,N_906,N_700);
nor U1220 (N_1220,N_955,N_593);
or U1221 (N_1221,N_144,N_817);
nand U1222 (N_1222,N_391,N_462);
nor U1223 (N_1223,N_100,N_485);
nor U1224 (N_1224,N_645,N_121);
or U1225 (N_1225,N_309,N_875);
and U1226 (N_1226,N_313,N_126);
nand U1227 (N_1227,N_354,N_153);
nor U1228 (N_1228,N_635,N_359);
and U1229 (N_1229,N_16,N_617);
and U1230 (N_1230,N_896,N_59);
or U1231 (N_1231,N_107,N_783);
nor U1232 (N_1232,N_658,N_235);
nand U1233 (N_1233,N_682,N_742);
or U1234 (N_1234,N_904,N_478);
nor U1235 (N_1235,N_825,N_590);
nand U1236 (N_1236,N_350,N_770);
xor U1237 (N_1237,N_758,N_425);
nor U1238 (N_1238,N_434,N_240);
nor U1239 (N_1239,N_250,N_177);
nand U1240 (N_1240,N_805,N_912);
nand U1241 (N_1241,N_138,N_171);
xor U1242 (N_1242,N_214,N_258);
and U1243 (N_1243,N_360,N_601);
or U1244 (N_1244,N_717,N_230);
nor U1245 (N_1245,N_420,N_147);
and U1246 (N_1246,N_576,N_253);
and U1247 (N_1247,N_438,N_419);
nand U1248 (N_1248,N_755,N_691);
nor U1249 (N_1249,N_130,N_606);
and U1250 (N_1250,N_931,N_276);
and U1251 (N_1251,N_382,N_93);
nor U1252 (N_1252,N_215,N_657);
or U1253 (N_1253,N_450,N_989);
nor U1254 (N_1254,N_907,N_315);
and U1255 (N_1255,N_102,N_342);
and U1256 (N_1256,N_648,N_868);
or U1257 (N_1257,N_688,N_668);
or U1258 (N_1258,N_132,N_788);
nand U1259 (N_1259,N_515,N_724);
nor U1260 (N_1260,N_155,N_675);
and U1261 (N_1261,N_208,N_632);
or U1262 (N_1262,N_449,N_843);
and U1263 (N_1263,N_71,N_873);
xnor U1264 (N_1264,N_558,N_603);
and U1265 (N_1265,N_75,N_287);
and U1266 (N_1266,N_383,N_394);
and U1267 (N_1267,N_422,N_299);
or U1268 (N_1268,N_507,N_806);
or U1269 (N_1269,N_161,N_111);
and U1270 (N_1270,N_523,N_185);
nand U1271 (N_1271,N_168,N_761);
xor U1272 (N_1272,N_129,N_134);
and U1273 (N_1273,N_18,N_910);
nor U1274 (N_1274,N_646,N_864);
nor U1275 (N_1275,N_535,N_939);
and U1276 (N_1276,N_693,N_64);
nor U1277 (N_1277,N_347,N_899);
and U1278 (N_1278,N_491,N_977);
and U1279 (N_1279,N_976,N_77);
or U1280 (N_1280,N_916,N_555);
xnor U1281 (N_1281,N_982,N_926);
xor U1282 (N_1282,N_409,N_736);
or U1283 (N_1283,N_339,N_402);
nand U1284 (N_1284,N_588,N_655);
nor U1285 (N_1285,N_355,N_439);
or U1286 (N_1286,N_839,N_892);
or U1287 (N_1287,N_136,N_860);
or U1288 (N_1288,N_159,N_863);
and U1289 (N_1289,N_494,N_306);
and U1290 (N_1290,N_837,N_66);
nor U1291 (N_1291,N_211,N_410);
xnor U1292 (N_1292,N_176,N_428);
xnor U1293 (N_1293,N_511,N_954);
or U1294 (N_1294,N_242,N_120);
nor U1295 (N_1295,N_6,N_397);
and U1296 (N_1296,N_503,N_119);
nor U1297 (N_1297,N_311,N_544);
or U1298 (N_1298,N_160,N_152);
xor U1299 (N_1299,N_987,N_998);
nor U1300 (N_1300,N_190,N_103);
or U1301 (N_1301,N_239,N_990);
and U1302 (N_1302,N_633,N_319);
or U1303 (N_1303,N_775,N_563);
nand U1304 (N_1304,N_78,N_322);
or U1305 (N_1305,N_192,N_145);
or U1306 (N_1306,N_162,N_527);
or U1307 (N_1307,N_747,N_838);
nand U1308 (N_1308,N_925,N_803);
or U1309 (N_1309,N_594,N_321);
nand U1310 (N_1310,N_79,N_356);
and U1311 (N_1311,N_95,N_502);
nand U1312 (N_1312,N_640,N_819);
and U1313 (N_1313,N_366,N_385);
nor U1314 (N_1314,N_388,N_665);
nand U1315 (N_1315,N_777,N_631);
nand U1316 (N_1316,N_759,N_553);
nand U1317 (N_1317,N_277,N_953);
nor U1318 (N_1318,N_711,N_241);
nand U1319 (N_1319,N_122,N_801);
nor U1320 (N_1320,N_735,N_399);
nand U1321 (N_1321,N_712,N_697);
or U1322 (N_1322,N_713,N_738);
and U1323 (N_1323,N_21,N_472);
nor U1324 (N_1324,N_569,N_282);
nand U1325 (N_1325,N_358,N_476);
nor U1326 (N_1326,N_879,N_295);
or U1327 (N_1327,N_390,N_150);
or U1328 (N_1328,N_331,N_229);
and U1329 (N_1329,N_294,N_991);
or U1330 (N_1330,N_195,N_994);
nor U1331 (N_1331,N_274,N_148);
xor U1332 (N_1332,N_856,N_46);
nand U1333 (N_1333,N_373,N_857);
nand U1334 (N_1334,N_934,N_374);
and U1335 (N_1335,N_27,N_914);
or U1336 (N_1336,N_654,N_396);
nor U1337 (N_1337,N_883,N_895);
and U1338 (N_1338,N_509,N_967);
or U1339 (N_1339,N_308,N_548);
or U1340 (N_1340,N_984,N_401);
and U1341 (N_1341,N_600,N_970);
nor U1342 (N_1342,N_112,N_114);
or U1343 (N_1343,N_585,N_944);
nand U1344 (N_1344,N_344,N_183);
xnor U1345 (N_1345,N_62,N_550);
xor U1346 (N_1346,N_424,N_504);
or U1347 (N_1347,N_257,N_219);
or U1348 (N_1348,N_793,N_530);
nor U1349 (N_1349,N_598,N_757);
and U1350 (N_1350,N_687,N_812);
nor U1351 (N_1351,N_751,N_469);
or U1352 (N_1352,N_483,N_850);
nor U1353 (N_1353,N_702,N_254);
nor U1354 (N_1354,N_781,N_468);
nand U1355 (N_1355,N_882,N_105);
or U1356 (N_1356,N_521,N_36);
or U1357 (N_1357,N_956,N_486);
nand U1358 (N_1358,N_859,N_470);
or U1359 (N_1359,N_437,N_495);
and U1360 (N_1360,N_799,N_141);
nor U1361 (N_1361,N_264,N_19);
or U1362 (N_1362,N_220,N_443);
nor U1363 (N_1363,N_763,N_999);
or U1364 (N_1364,N_901,N_774);
and U1365 (N_1365,N_888,N_510);
and U1366 (N_1366,N_407,N_487);
nor U1367 (N_1367,N_48,N_225);
or U1368 (N_1368,N_317,N_898);
or U1369 (N_1369,N_104,N_13);
or U1370 (N_1370,N_536,N_203);
nor U1371 (N_1371,N_975,N_936);
nor U1372 (N_1372,N_672,N_918);
nand U1373 (N_1373,N_418,N_988);
xor U1374 (N_1374,N_207,N_53);
nand U1375 (N_1375,N_39,N_894);
and U1376 (N_1376,N_432,N_51);
or U1377 (N_1377,N_96,N_247);
nor U1378 (N_1378,N_492,N_464);
or U1379 (N_1379,N_545,N_554);
xnor U1380 (N_1380,N_384,N_445);
or U1381 (N_1381,N_733,N_534);
and U1382 (N_1382,N_22,N_127);
xor U1383 (N_1383,N_966,N_175);
xnor U1384 (N_1384,N_526,N_587);
and U1385 (N_1385,N_506,N_538);
nand U1386 (N_1386,N_106,N_212);
and U1387 (N_1387,N_271,N_26);
or U1388 (N_1388,N_644,N_832);
nor U1389 (N_1389,N_403,N_218);
nand U1390 (N_1390,N_980,N_518);
and U1391 (N_1391,N_58,N_380);
and U1392 (N_1392,N_752,N_695);
and U1393 (N_1393,N_33,N_684);
nand U1394 (N_1394,N_435,N_604);
xor U1395 (N_1395,N_993,N_232);
and U1396 (N_1396,N_683,N_303);
xor U1397 (N_1397,N_615,N_245);
or U1398 (N_1398,N_173,N_115);
or U1399 (N_1399,N_978,N_969);
nor U1400 (N_1400,N_166,N_108);
and U1401 (N_1401,N_890,N_704);
nor U1402 (N_1402,N_867,N_835);
nand U1403 (N_1403,N_489,N_99);
nand U1404 (N_1404,N_72,N_87);
or U1405 (N_1405,N_656,N_881);
xor U1406 (N_1406,N_946,N_312);
and U1407 (N_1407,N_221,N_477);
and U1408 (N_1408,N_131,N_109);
nand U1409 (N_1409,N_163,N_519);
nand U1410 (N_1410,N_412,N_637);
or U1411 (N_1411,N_573,N_283);
and U1412 (N_1412,N_281,N_623);
nor U1413 (N_1413,N_878,N_950);
and U1414 (N_1414,N_798,N_730);
or U1415 (N_1415,N_725,N_474);
nor U1416 (N_1416,N_463,N_522);
nor U1417 (N_1417,N_37,N_578);
nand U1418 (N_1418,N_532,N_830);
and U1419 (N_1419,N_340,N_320);
and U1420 (N_1420,N_571,N_25);
nand U1421 (N_1421,N_708,N_842);
nor U1422 (N_1422,N_63,N_599);
xor U1423 (N_1423,N_923,N_943);
nor U1424 (N_1424,N_500,N_268);
or U1425 (N_1425,N_662,N_508);
nor U1426 (N_1426,N_328,N_198);
or U1427 (N_1427,N_179,N_792);
and U1428 (N_1428,N_193,N_666);
or U1429 (N_1429,N_673,N_209);
or U1430 (N_1430,N_83,N_446);
and U1431 (N_1431,N_86,N_327);
nor U1432 (N_1432,N_566,N_260);
nor U1433 (N_1433,N_574,N_516);
or U1434 (N_1434,N_65,N_911);
nor U1435 (N_1435,N_802,N_73);
or U1436 (N_1436,N_233,N_456);
nand U1437 (N_1437,N_479,N_659);
and U1438 (N_1438,N_167,N_223);
nor U1439 (N_1439,N_298,N_992);
nand U1440 (N_1440,N_23,N_40);
or U1441 (N_1441,N_110,N_556);
nand U1442 (N_1442,N_415,N_41);
and U1443 (N_1443,N_398,N_178);
and U1444 (N_1444,N_539,N_411);
or U1445 (N_1445,N_754,N_705);
xor U1446 (N_1446,N_15,N_149);
and U1447 (N_1447,N_753,N_496);
nand U1448 (N_1448,N_570,N_55);
or U1449 (N_1449,N_723,N_498);
or U1450 (N_1450,N_20,N_296);
or U1451 (N_1451,N_459,N_353);
or U1452 (N_1452,N_205,N_465);
or U1453 (N_1453,N_416,N_756);
xnor U1454 (N_1454,N_638,N_869);
and U1455 (N_1455,N_720,N_52);
xnor U1456 (N_1456,N_607,N_562);
nand U1457 (N_1457,N_627,N_267);
nor U1458 (N_1458,N_154,N_790);
and U1459 (N_1459,N_34,N_67);
nand U1460 (N_1460,N_97,N_872);
or U1461 (N_1461,N_728,N_855);
or U1462 (N_1462,N_917,N_361);
and U1463 (N_1463,N_142,N_961);
or U1464 (N_1464,N_952,N_352);
nor U1465 (N_1465,N_333,N_499);
or U1466 (N_1466,N_326,N_866);
nand U1467 (N_1467,N_473,N_815);
or U1468 (N_1468,N_951,N_715);
and U1469 (N_1469,N_680,N_441);
nand U1470 (N_1470,N_74,N_2);
or U1471 (N_1471,N_597,N_807);
or U1472 (N_1472,N_417,N_718);
nor U1473 (N_1473,N_981,N_965);
nand U1474 (N_1474,N_565,N_324);
nor U1475 (N_1475,N_653,N_76);
nand U1476 (N_1476,N_451,N_3);
nand U1477 (N_1477,N_10,N_559);
nor U1478 (N_1478,N_316,N_431);
and U1479 (N_1479,N_620,N_453);
nand U1480 (N_1480,N_826,N_70);
or U1481 (N_1481,N_591,N_484);
xor U1482 (N_1482,N_722,N_293);
or U1483 (N_1483,N_557,N_734);
nor U1484 (N_1484,N_12,N_703);
nand U1485 (N_1485,N_610,N_608);
nor U1486 (N_1486,N_187,N_305);
nor U1487 (N_1487,N_227,N_650);
and U1488 (N_1488,N_900,N_828);
nand U1489 (N_1489,N_628,N_88);
and U1490 (N_1490,N_816,N_996);
xor U1491 (N_1491,N_786,N_552);
nand U1492 (N_1492,N_252,N_113);
and U1493 (N_1493,N_732,N_467);
nand U1494 (N_1494,N_748,N_582);
nand U1495 (N_1495,N_124,N_647);
and U1496 (N_1496,N_809,N_128);
or U1497 (N_1497,N_846,N_973);
nand U1498 (N_1498,N_616,N_47);
or U1499 (N_1499,N_447,N_44);
and U1500 (N_1500,N_539,N_850);
nand U1501 (N_1501,N_223,N_591);
nor U1502 (N_1502,N_108,N_707);
nor U1503 (N_1503,N_973,N_458);
nand U1504 (N_1504,N_896,N_709);
nor U1505 (N_1505,N_345,N_375);
and U1506 (N_1506,N_867,N_116);
and U1507 (N_1507,N_604,N_580);
nor U1508 (N_1508,N_74,N_825);
nand U1509 (N_1509,N_196,N_786);
nor U1510 (N_1510,N_749,N_207);
nor U1511 (N_1511,N_312,N_688);
nor U1512 (N_1512,N_588,N_739);
nand U1513 (N_1513,N_271,N_908);
and U1514 (N_1514,N_966,N_652);
nor U1515 (N_1515,N_851,N_27);
and U1516 (N_1516,N_212,N_799);
or U1517 (N_1517,N_985,N_511);
nor U1518 (N_1518,N_484,N_990);
or U1519 (N_1519,N_663,N_923);
nor U1520 (N_1520,N_259,N_451);
nand U1521 (N_1521,N_853,N_840);
nand U1522 (N_1522,N_675,N_669);
and U1523 (N_1523,N_721,N_571);
and U1524 (N_1524,N_243,N_252);
or U1525 (N_1525,N_696,N_371);
nand U1526 (N_1526,N_395,N_754);
nor U1527 (N_1527,N_882,N_36);
or U1528 (N_1528,N_317,N_640);
xnor U1529 (N_1529,N_690,N_810);
and U1530 (N_1530,N_131,N_890);
xnor U1531 (N_1531,N_71,N_423);
nor U1532 (N_1532,N_892,N_835);
and U1533 (N_1533,N_397,N_589);
nor U1534 (N_1534,N_12,N_553);
and U1535 (N_1535,N_752,N_580);
nor U1536 (N_1536,N_290,N_496);
and U1537 (N_1537,N_568,N_592);
xnor U1538 (N_1538,N_327,N_121);
nand U1539 (N_1539,N_203,N_496);
nand U1540 (N_1540,N_443,N_927);
nand U1541 (N_1541,N_674,N_57);
nand U1542 (N_1542,N_888,N_673);
and U1543 (N_1543,N_372,N_309);
and U1544 (N_1544,N_50,N_736);
and U1545 (N_1545,N_532,N_883);
nand U1546 (N_1546,N_593,N_499);
nor U1547 (N_1547,N_303,N_467);
and U1548 (N_1548,N_315,N_196);
nor U1549 (N_1549,N_425,N_446);
nor U1550 (N_1550,N_715,N_742);
and U1551 (N_1551,N_606,N_991);
or U1552 (N_1552,N_970,N_247);
nor U1553 (N_1553,N_639,N_50);
and U1554 (N_1554,N_391,N_330);
nand U1555 (N_1555,N_442,N_880);
or U1556 (N_1556,N_673,N_485);
nand U1557 (N_1557,N_46,N_928);
and U1558 (N_1558,N_6,N_794);
or U1559 (N_1559,N_473,N_311);
and U1560 (N_1560,N_164,N_199);
nor U1561 (N_1561,N_780,N_167);
nand U1562 (N_1562,N_475,N_56);
nand U1563 (N_1563,N_446,N_172);
and U1564 (N_1564,N_745,N_579);
or U1565 (N_1565,N_937,N_695);
nor U1566 (N_1566,N_810,N_825);
and U1567 (N_1567,N_349,N_640);
and U1568 (N_1568,N_926,N_64);
nor U1569 (N_1569,N_509,N_214);
nor U1570 (N_1570,N_652,N_997);
and U1571 (N_1571,N_975,N_65);
and U1572 (N_1572,N_165,N_608);
or U1573 (N_1573,N_845,N_38);
nor U1574 (N_1574,N_808,N_949);
xor U1575 (N_1575,N_531,N_729);
nor U1576 (N_1576,N_629,N_651);
nand U1577 (N_1577,N_310,N_109);
nand U1578 (N_1578,N_879,N_103);
nor U1579 (N_1579,N_629,N_864);
and U1580 (N_1580,N_392,N_910);
nand U1581 (N_1581,N_1,N_259);
xnor U1582 (N_1582,N_119,N_939);
nand U1583 (N_1583,N_578,N_506);
nand U1584 (N_1584,N_287,N_776);
and U1585 (N_1585,N_931,N_829);
nor U1586 (N_1586,N_192,N_800);
nand U1587 (N_1587,N_791,N_170);
nand U1588 (N_1588,N_680,N_719);
xor U1589 (N_1589,N_654,N_330);
or U1590 (N_1590,N_651,N_29);
xnor U1591 (N_1591,N_660,N_791);
and U1592 (N_1592,N_279,N_411);
nor U1593 (N_1593,N_204,N_925);
or U1594 (N_1594,N_645,N_595);
nor U1595 (N_1595,N_137,N_127);
and U1596 (N_1596,N_741,N_981);
nand U1597 (N_1597,N_668,N_875);
or U1598 (N_1598,N_925,N_532);
or U1599 (N_1599,N_730,N_321);
nand U1600 (N_1600,N_83,N_894);
nor U1601 (N_1601,N_292,N_314);
and U1602 (N_1602,N_185,N_8);
nor U1603 (N_1603,N_943,N_473);
or U1604 (N_1604,N_659,N_930);
nand U1605 (N_1605,N_865,N_565);
nand U1606 (N_1606,N_331,N_657);
nand U1607 (N_1607,N_385,N_282);
xor U1608 (N_1608,N_992,N_941);
or U1609 (N_1609,N_382,N_670);
and U1610 (N_1610,N_757,N_773);
xnor U1611 (N_1611,N_35,N_785);
nor U1612 (N_1612,N_916,N_589);
nand U1613 (N_1613,N_718,N_879);
or U1614 (N_1614,N_397,N_667);
or U1615 (N_1615,N_689,N_846);
or U1616 (N_1616,N_336,N_631);
nand U1617 (N_1617,N_730,N_752);
nor U1618 (N_1618,N_928,N_841);
nor U1619 (N_1619,N_181,N_781);
nor U1620 (N_1620,N_344,N_74);
nor U1621 (N_1621,N_199,N_181);
nand U1622 (N_1622,N_737,N_864);
nand U1623 (N_1623,N_119,N_537);
or U1624 (N_1624,N_61,N_145);
and U1625 (N_1625,N_763,N_234);
or U1626 (N_1626,N_360,N_324);
xnor U1627 (N_1627,N_407,N_416);
xor U1628 (N_1628,N_216,N_284);
and U1629 (N_1629,N_667,N_610);
or U1630 (N_1630,N_213,N_331);
xnor U1631 (N_1631,N_476,N_501);
nand U1632 (N_1632,N_491,N_952);
nand U1633 (N_1633,N_341,N_206);
nor U1634 (N_1634,N_594,N_723);
nor U1635 (N_1635,N_961,N_797);
and U1636 (N_1636,N_829,N_504);
and U1637 (N_1637,N_857,N_919);
nand U1638 (N_1638,N_147,N_829);
nand U1639 (N_1639,N_192,N_518);
nor U1640 (N_1640,N_576,N_942);
nand U1641 (N_1641,N_203,N_458);
xnor U1642 (N_1642,N_321,N_906);
and U1643 (N_1643,N_581,N_237);
nand U1644 (N_1644,N_540,N_488);
or U1645 (N_1645,N_983,N_328);
xnor U1646 (N_1646,N_135,N_711);
or U1647 (N_1647,N_195,N_789);
nor U1648 (N_1648,N_38,N_312);
xor U1649 (N_1649,N_772,N_319);
or U1650 (N_1650,N_150,N_715);
and U1651 (N_1651,N_920,N_313);
or U1652 (N_1652,N_109,N_709);
nand U1653 (N_1653,N_544,N_51);
and U1654 (N_1654,N_812,N_940);
and U1655 (N_1655,N_190,N_258);
and U1656 (N_1656,N_336,N_210);
or U1657 (N_1657,N_705,N_893);
xor U1658 (N_1658,N_283,N_669);
and U1659 (N_1659,N_20,N_628);
and U1660 (N_1660,N_320,N_941);
or U1661 (N_1661,N_538,N_6);
and U1662 (N_1662,N_557,N_883);
nand U1663 (N_1663,N_265,N_521);
and U1664 (N_1664,N_521,N_871);
and U1665 (N_1665,N_131,N_403);
nor U1666 (N_1666,N_564,N_353);
xor U1667 (N_1667,N_349,N_812);
nand U1668 (N_1668,N_208,N_352);
or U1669 (N_1669,N_77,N_362);
or U1670 (N_1670,N_624,N_109);
or U1671 (N_1671,N_258,N_82);
nor U1672 (N_1672,N_200,N_531);
and U1673 (N_1673,N_411,N_727);
or U1674 (N_1674,N_795,N_527);
nor U1675 (N_1675,N_614,N_999);
and U1676 (N_1676,N_738,N_137);
and U1677 (N_1677,N_403,N_175);
or U1678 (N_1678,N_275,N_533);
nand U1679 (N_1679,N_914,N_799);
and U1680 (N_1680,N_917,N_567);
nand U1681 (N_1681,N_9,N_548);
or U1682 (N_1682,N_70,N_915);
or U1683 (N_1683,N_838,N_507);
and U1684 (N_1684,N_840,N_861);
nor U1685 (N_1685,N_38,N_259);
or U1686 (N_1686,N_362,N_512);
nand U1687 (N_1687,N_764,N_33);
or U1688 (N_1688,N_28,N_78);
nor U1689 (N_1689,N_678,N_428);
xnor U1690 (N_1690,N_108,N_685);
nor U1691 (N_1691,N_146,N_511);
nor U1692 (N_1692,N_952,N_165);
nor U1693 (N_1693,N_835,N_382);
nor U1694 (N_1694,N_171,N_181);
nand U1695 (N_1695,N_902,N_81);
xnor U1696 (N_1696,N_247,N_324);
nand U1697 (N_1697,N_813,N_595);
nor U1698 (N_1698,N_547,N_94);
nand U1699 (N_1699,N_690,N_109);
and U1700 (N_1700,N_703,N_624);
nand U1701 (N_1701,N_330,N_238);
and U1702 (N_1702,N_734,N_189);
or U1703 (N_1703,N_605,N_296);
and U1704 (N_1704,N_858,N_282);
nor U1705 (N_1705,N_678,N_974);
xor U1706 (N_1706,N_748,N_679);
and U1707 (N_1707,N_507,N_237);
nor U1708 (N_1708,N_534,N_204);
and U1709 (N_1709,N_867,N_83);
and U1710 (N_1710,N_341,N_286);
nor U1711 (N_1711,N_700,N_73);
xor U1712 (N_1712,N_615,N_45);
or U1713 (N_1713,N_235,N_723);
or U1714 (N_1714,N_168,N_369);
and U1715 (N_1715,N_20,N_232);
or U1716 (N_1716,N_386,N_193);
nand U1717 (N_1717,N_985,N_688);
or U1718 (N_1718,N_474,N_352);
nand U1719 (N_1719,N_176,N_873);
and U1720 (N_1720,N_0,N_249);
or U1721 (N_1721,N_919,N_259);
xnor U1722 (N_1722,N_477,N_152);
nand U1723 (N_1723,N_774,N_135);
nand U1724 (N_1724,N_558,N_562);
and U1725 (N_1725,N_980,N_575);
or U1726 (N_1726,N_437,N_709);
or U1727 (N_1727,N_330,N_257);
xnor U1728 (N_1728,N_337,N_417);
or U1729 (N_1729,N_840,N_769);
and U1730 (N_1730,N_804,N_378);
nor U1731 (N_1731,N_869,N_967);
nor U1732 (N_1732,N_930,N_717);
or U1733 (N_1733,N_675,N_335);
nand U1734 (N_1734,N_62,N_863);
nor U1735 (N_1735,N_675,N_467);
nor U1736 (N_1736,N_119,N_312);
and U1737 (N_1737,N_746,N_468);
or U1738 (N_1738,N_112,N_856);
or U1739 (N_1739,N_364,N_367);
nand U1740 (N_1740,N_615,N_96);
or U1741 (N_1741,N_381,N_814);
and U1742 (N_1742,N_362,N_150);
or U1743 (N_1743,N_806,N_497);
xor U1744 (N_1744,N_405,N_344);
or U1745 (N_1745,N_435,N_658);
nor U1746 (N_1746,N_883,N_993);
nand U1747 (N_1747,N_842,N_435);
nor U1748 (N_1748,N_398,N_570);
and U1749 (N_1749,N_957,N_39);
nand U1750 (N_1750,N_933,N_158);
xor U1751 (N_1751,N_161,N_663);
xor U1752 (N_1752,N_177,N_524);
or U1753 (N_1753,N_561,N_498);
nor U1754 (N_1754,N_311,N_657);
or U1755 (N_1755,N_603,N_661);
and U1756 (N_1756,N_847,N_503);
nand U1757 (N_1757,N_672,N_483);
nand U1758 (N_1758,N_827,N_723);
nor U1759 (N_1759,N_115,N_543);
xnor U1760 (N_1760,N_71,N_280);
nor U1761 (N_1761,N_856,N_940);
xor U1762 (N_1762,N_696,N_269);
xor U1763 (N_1763,N_935,N_543);
and U1764 (N_1764,N_417,N_317);
xor U1765 (N_1765,N_851,N_682);
nor U1766 (N_1766,N_762,N_277);
and U1767 (N_1767,N_297,N_17);
and U1768 (N_1768,N_37,N_796);
or U1769 (N_1769,N_79,N_909);
and U1770 (N_1770,N_384,N_60);
nor U1771 (N_1771,N_214,N_419);
xnor U1772 (N_1772,N_825,N_327);
nand U1773 (N_1773,N_979,N_574);
xor U1774 (N_1774,N_963,N_157);
xnor U1775 (N_1775,N_663,N_408);
or U1776 (N_1776,N_665,N_842);
nand U1777 (N_1777,N_694,N_484);
and U1778 (N_1778,N_580,N_382);
nor U1779 (N_1779,N_440,N_900);
nand U1780 (N_1780,N_835,N_836);
or U1781 (N_1781,N_459,N_776);
xor U1782 (N_1782,N_192,N_506);
nand U1783 (N_1783,N_260,N_33);
and U1784 (N_1784,N_495,N_458);
and U1785 (N_1785,N_621,N_44);
nor U1786 (N_1786,N_129,N_752);
or U1787 (N_1787,N_438,N_116);
or U1788 (N_1788,N_748,N_295);
nor U1789 (N_1789,N_607,N_702);
nor U1790 (N_1790,N_205,N_293);
nor U1791 (N_1791,N_595,N_173);
and U1792 (N_1792,N_190,N_59);
or U1793 (N_1793,N_139,N_859);
or U1794 (N_1794,N_124,N_50);
nor U1795 (N_1795,N_674,N_779);
and U1796 (N_1796,N_720,N_492);
nor U1797 (N_1797,N_454,N_562);
or U1798 (N_1798,N_854,N_133);
nand U1799 (N_1799,N_399,N_58);
nor U1800 (N_1800,N_370,N_314);
nand U1801 (N_1801,N_249,N_534);
xnor U1802 (N_1802,N_71,N_261);
nand U1803 (N_1803,N_533,N_737);
nand U1804 (N_1804,N_10,N_853);
or U1805 (N_1805,N_437,N_480);
or U1806 (N_1806,N_639,N_869);
and U1807 (N_1807,N_563,N_140);
xor U1808 (N_1808,N_168,N_754);
nor U1809 (N_1809,N_98,N_155);
and U1810 (N_1810,N_83,N_833);
and U1811 (N_1811,N_76,N_104);
nor U1812 (N_1812,N_79,N_805);
nor U1813 (N_1813,N_666,N_437);
nor U1814 (N_1814,N_163,N_542);
nor U1815 (N_1815,N_429,N_552);
xnor U1816 (N_1816,N_860,N_998);
xnor U1817 (N_1817,N_454,N_923);
nor U1818 (N_1818,N_321,N_890);
and U1819 (N_1819,N_606,N_204);
or U1820 (N_1820,N_578,N_467);
or U1821 (N_1821,N_774,N_837);
xor U1822 (N_1822,N_523,N_348);
or U1823 (N_1823,N_706,N_900);
xor U1824 (N_1824,N_876,N_822);
or U1825 (N_1825,N_910,N_404);
and U1826 (N_1826,N_842,N_749);
nor U1827 (N_1827,N_140,N_915);
nand U1828 (N_1828,N_295,N_460);
or U1829 (N_1829,N_212,N_894);
or U1830 (N_1830,N_399,N_177);
nor U1831 (N_1831,N_401,N_259);
and U1832 (N_1832,N_463,N_613);
xnor U1833 (N_1833,N_428,N_114);
or U1834 (N_1834,N_24,N_92);
and U1835 (N_1835,N_184,N_233);
xnor U1836 (N_1836,N_924,N_91);
nor U1837 (N_1837,N_892,N_384);
or U1838 (N_1838,N_760,N_753);
or U1839 (N_1839,N_333,N_326);
nand U1840 (N_1840,N_651,N_8);
nand U1841 (N_1841,N_53,N_684);
nor U1842 (N_1842,N_914,N_434);
nor U1843 (N_1843,N_846,N_680);
or U1844 (N_1844,N_820,N_836);
and U1845 (N_1845,N_483,N_980);
or U1846 (N_1846,N_482,N_455);
nor U1847 (N_1847,N_544,N_873);
nand U1848 (N_1848,N_935,N_598);
or U1849 (N_1849,N_435,N_791);
and U1850 (N_1850,N_340,N_198);
nand U1851 (N_1851,N_482,N_213);
nand U1852 (N_1852,N_902,N_943);
nor U1853 (N_1853,N_983,N_533);
and U1854 (N_1854,N_534,N_941);
or U1855 (N_1855,N_222,N_828);
xor U1856 (N_1856,N_88,N_983);
xnor U1857 (N_1857,N_293,N_911);
xnor U1858 (N_1858,N_786,N_263);
and U1859 (N_1859,N_461,N_941);
nor U1860 (N_1860,N_495,N_118);
xor U1861 (N_1861,N_725,N_30);
nor U1862 (N_1862,N_275,N_410);
nand U1863 (N_1863,N_286,N_754);
or U1864 (N_1864,N_590,N_441);
nor U1865 (N_1865,N_88,N_568);
nor U1866 (N_1866,N_833,N_743);
or U1867 (N_1867,N_525,N_865);
and U1868 (N_1868,N_874,N_539);
nand U1869 (N_1869,N_584,N_870);
and U1870 (N_1870,N_916,N_365);
nor U1871 (N_1871,N_437,N_881);
or U1872 (N_1872,N_804,N_21);
nand U1873 (N_1873,N_723,N_221);
or U1874 (N_1874,N_776,N_437);
nor U1875 (N_1875,N_874,N_117);
xnor U1876 (N_1876,N_829,N_440);
and U1877 (N_1877,N_475,N_500);
nor U1878 (N_1878,N_520,N_539);
and U1879 (N_1879,N_305,N_442);
and U1880 (N_1880,N_943,N_931);
and U1881 (N_1881,N_615,N_756);
xnor U1882 (N_1882,N_523,N_878);
nor U1883 (N_1883,N_943,N_151);
nor U1884 (N_1884,N_312,N_622);
xnor U1885 (N_1885,N_458,N_910);
nand U1886 (N_1886,N_536,N_685);
and U1887 (N_1887,N_872,N_331);
and U1888 (N_1888,N_772,N_922);
and U1889 (N_1889,N_316,N_985);
nand U1890 (N_1890,N_893,N_900);
nor U1891 (N_1891,N_251,N_411);
and U1892 (N_1892,N_440,N_101);
nor U1893 (N_1893,N_585,N_860);
nand U1894 (N_1894,N_115,N_755);
or U1895 (N_1895,N_190,N_74);
and U1896 (N_1896,N_761,N_61);
xor U1897 (N_1897,N_658,N_169);
and U1898 (N_1898,N_550,N_726);
nor U1899 (N_1899,N_797,N_853);
or U1900 (N_1900,N_208,N_651);
nand U1901 (N_1901,N_123,N_999);
nand U1902 (N_1902,N_954,N_684);
and U1903 (N_1903,N_361,N_105);
or U1904 (N_1904,N_858,N_592);
and U1905 (N_1905,N_246,N_680);
and U1906 (N_1906,N_355,N_965);
nand U1907 (N_1907,N_939,N_559);
nor U1908 (N_1908,N_783,N_263);
nor U1909 (N_1909,N_534,N_49);
and U1910 (N_1910,N_362,N_159);
nor U1911 (N_1911,N_298,N_491);
nand U1912 (N_1912,N_413,N_311);
nor U1913 (N_1913,N_640,N_702);
nand U1914 (N_1914,N_486,N_131);
or U1915 (N_1915,N_35,N_388);
and U1916 (N_1916,N_452,N_460);
or U1917 (N_1917,N_386,N_204);
and U1918 (N_1918,N_859,N_662);
nand U1919 (N_1919,N_29,N_567);
or U1920 (N_1920,N_945,N_325);
xor U1921 (N_1921,N_919,N_304);
xor U1922 (N_1922,N_728,N_59);
nand U1923 (N_1923,N_342,N_79);
nand U1924 (N_1924,N_743,N_518);
nand U1925 (N_1925,N_994,N_884);
and U1926 (N_1926,N_706,N_478);
and U1927 (N_1927,N_166,N_993);
and U1928 (N_1928,N_996,N_185);
and U1929 (N_1929,N_130,N_958);
or U1930 (N_1930,N_707,N_265);
or U1931 (N_1931,N_183,N_476);
and U1932 (N_1932,N_36,N_796);
xnor U1933 (N_1933,N_515,N_657);
nand U1934 (N_1934,N_736,N_428);
nor U1935 (N_1935,N_562,N_22);
xnor U1936 (N_1936,N_487,N_165);
or U1937 (N_1937,N_695,N_930);
nor U1938 (N_1938,N_702,N_121);
nor U1939 (N_1939,N_162,N_93);
xnor U1940 (N_1940,N_241,N_174);
nor U1941 (N_1941,N_321,N_683);
and U1942 (N_1942,N_713,N_819);
nor U1943 (N_1943,N_830,N_104);
nor U1944 (N_1944,N_297,N_508);
nand U1945 (N_1945,N_703,N_997);
nand U1946 (N_1946,N_332,N_612);
and U1947 (N_1947,N_770,N_363);
xnor U1948 (N_1948,N_282,N_643);
nor U1949 (N_1949,N_265,N_535);
nor U1950 (N_1950,N_944,N_306);
or U1951 (N_1951,N_277,N_70);
nor U1952 (N_1952,N_843,N_143);
xnor U1953 (N_1953,N_170,N_294);
nor U1954 (N_1954,N_185,N_725);
nand U1955 (N_1955,N_461,N_276);
or U1956 (N_1956,N_545,N_462);
nand U1957 (N_1957,N_393,N_490);
or U1958 (N_1958,N_325,N_501);
and U1959 (N_1959,N_712,N_637);
and U1960 (N_1960,N_10,N_653);
and U1961 (N_1961,N_38,N_399);
xor U1962 (N_1962,N_971,N_772);
nor U1963 (N_1963,N_53,N_356);
or U1964 (N_1964,N_544,N_989);
and U1965 (N_1965,N_993,N_507);
and U1966 (N_1966,N_542,N_383);
nor U1967 (N_1967,N_612,N_0);
and U1968 (N_1968,N_44,N_896);
nor U1969 (N_1969,N_571,N_924);
or U1970 (N_1970,N_842,N_867);
or U1971 (N_1971,N_529,N_989);
or U1972 (N_1972,N_598,N_633);
or U1973 (N_1973,N_190,N_921);
and U1974 (N_1974,N_26,N_457);
and U1975 (N_1975,N_957,N_235);
xor U1976 (N_1976,N_863,N_607);
nor U1977 (N_1977,N_898,N_974);
and U1978 (N_1978,N_701,N_0);
nand U1979 (N_1979,N_630,N_55);
or U1980 (N_1980,N_490,N_893);
nor U1981 (N_1981,N_858,N_218);
or U1982 (N_1982,N_222,N_701);
xnor U1983 (N_1983,N_876,N_239);
nor U1984 (N_1984,N_154,N_486);
nor U1985 (N_1985,N_812,N_586);
nand U1986 (N_1986,N_586,N_273);
nand U1987 (N_1987,N_362,N_261);
and U1988 (N_1988,N_752,N_453);
nor U1989 (N_1989,N_451,N_777);
or U1990 (N_1990,N_594,N_620);
nor U1991 (N_1991,N_673,N_817);
or U1992 (N_1992,N_933,N_193);
or U1993 (N_1993,N_58,N_391);
and U1994 (N_1994,N_553,N_461);
or U1995 (N_1995,N_11,N_254);
nor U1996 (N_1996,N_152,N_951);
and U1997 (N_1997,N_621,N_841);
and U1998 (N_1998,N_581,N_864);
and U1999 (N_1999,N_34,N_746);
and U2000 (N_2000,N_1838,N_1957);
nand U2001 (N_2001,N_1932,N_1877);
nand U2002 (N_2002,N_1496,N_1105);
nor U2003 (N_2003,N_1761,N_1835);
nand U2004 (N_2004,N_1902,N_1941);
nor U2005 (N_2005,N_1412,N_1491);
nor U2006 (N_2006,N_1899,N_1148);
and U2007 (N_2007,N_1219,N_1182);
and U2008 (N_2008,N_1828,N_1458);
and U2009 (N_2009,N_1631,N_1717);
or U2010 (N_2010,N_1951,N_1041);
or U2011 (N_2011,N_1548,N_1969);
nand U2012 (N_2012,N_1664,N_1065);
nand U2013 (N_2013,N_1366,N_1968);
or U2014 (N_2014,N_1830,N_1947);
xor U2015 (N_2015,N_1441,N_1840);
nand U2016 (N_2016,N_1422,N_1111);
nor U2017 (N_2017,N_1874,N_1134);
and U2018 (N_2018,N_1284,N_1628);
nand U2019 (N_2019,N_1948,N_1497);
and U2020 (N_2020,N_1652,N_1019);
nor U2021 (N_2021,N_1925,N_1586);
nor U2022 (N_2022,N_1821,N_1788);
nor U2023 (N_2023,N_1097,N_1248);
xnor U2024 (N_2024,N_1391,N_1725);
nand U2025 (N_2025,N_1171,N_1075);
nor U2026 (N_2026,N_1605,N_1343);
or U2027 (N_2027,N_1876,N_1591);
xor U2028 (N_2028,N_1678,N_1798);
or U2029 (N_2029,N_1519,N_1723);
nor U2030 (N_2030,N_1047,N_1989);
and U2031 (N_2031,N_1571,N_1885);
and U2032 (N_2032,N_1595,N_1699);
and U2033 (N_2033,N_1118,N_1375);
nor U2034 (N_2034,N_1260,N_1855);
and U2035 (N_2035,N_1800,N_1220);
and U2036 (N_2036,N_1641,N_1367);
nand U2037 (N_2037,N_1898,N_1238);
and U2038 (N_2038,N_1977,N_1550);
and U2039 (N_2039,N_1241,N_1671);
xor U2040 (N_2040,N_1311,N_1890);
nor U2041 (N_2041,N_1377,N_1214);
xnor U2042 (N_2042,N_1648,N_1132);
and U2043 (N_2043,N_1013,N_1954);
nor U2044 (N_2044,N_1558,N_1848);
and U2045 (N_2045,N_1833,N_1263);
and U2046 (N_2046,N_1368,N_1727);
nand U2047 (N_2047,N_1089,N_1495);
nor U2048 (N_2048,N_1435,N_1991);
or U2049 (N_2049,N_1690,N_1625);
and U2050 (N_2050,N_1084,N_1135);
nand U2051 (N_2051,N_1577,N_1726);
nor U2052 (N_2052,N_1396,N_1159);
xnor U2053 (N_2053,N_1384,N_1862);
or U2054 (N_2054,N_1466,N_1538);
nand U2055 (N_2055,N_1554,N_1745);
and U2056 (N_2056,N_1479,N_1144);
or U2057 (N_2057,N_1967,N_1270);
and U2058 (N_2058,N_1101,N_1108);
or U2059 (N_2059,N_1752,N_1303);
nand U2060 (N_2060,N_1277,N_1295);
or U2061 (N_2061,N_1252,N_1770);
nand U2062 (N_2062,N_1975,N_1354);
nand U2063 (N_2063,N_1156,N_1693);
nand U2064 (N_2064,N_1506,N_1326);
xor U2065 (N_2065,N_1468,N_1846);
nor U2066 (N_2066,N_1228,N_1331);
and U2067 (N_2067,N_1492,N_1184);
and U2068 (N_2068,N_1891,N_1288);
or U2069 (N_2069,N_1024,N_1121);
nor U2070 (N_2070,N_1669,N_1404);
nand U2071 (N_2071,N_1981,N_1516);
or U2072 (N_2072,N_1837,N_1470);
xor U2073 (N_2073,N_1610,N_1552);
nor U2074 (N_2074,N_1361,N_1759);
nand U2075 (N_2075,N_1087,N_1204);
and U2076 (N_2076,N_1411,N_1455);
nor U2077 (N_2077,N_1477,N_1449);
and U2078 (N_2078,N_1243,N_1341);
or U2079 (N_2079,N_1911,N_1762);
and U2080 (N_2080,N_1253,N_1863);
or U2081 (N_2081,N_1465,N_1250);
or U2082 (N_2082,N_1199,N_1600);
nor U2083 (N_2083,N_1426,N_1212);
and U2084 (N_2084,N_1692,N_1149);
nor U2085 (N_2085,N_1033,N_1741);
and U2086 (N_2086,N_1390,N_1884);
or U2087 (N_2087,N_1486,N_1645);
or U2088 (N_2088,N_1432,N_1684);
or U2089 (N_2089,N_1680,N_1417);
nor U2090 (N_2090,N_1498,N_1882);
or U2091 (N_2091,N_1824,N_1859);
or U2092 (N_2092,N_1142,N_1870);
and U2093 (N_2093,N_1106,N_1454);
and U2094 (N_2094,N_1842,N_1461);
nor U2095 (N_2095,N_1520,N_1494);
and U2096 (N_2096,N_1999,N_1198);
xor U2097 (N_2097,N_1040,N_1609);
nor U2098 (N_2098,N_1191,N_1606);
xor U2099 (N_2099,N_1298,N_1488);
and U2100 (N_2100,N_1534,N_1124);
or U2101 (N_2101,N_1382,N_1537);
nand U2102 (N_2102,N_1236,N_1261);
nor U2103 (N_2103,N_1569,N_1061);
nor U2104 (N_2104,N_1005,N_1036);
nand U2105 (N_2105,N_1918,N_1383);
nand U2106 (N_2106,N_1878,N_1566);
and U2107 (N_2107,N_1100,N_1493);
nand U2108 (N_2108,N_1565,N_1173);
xnor U2109 (N_2109,N_1076,N_1117);
nand U2110 (N_2110,N_1827,N_1110);
and U2111 (N_2111,N_1147,N_1694);
nand U2112 (N_2112,N_1808,N_1414);
and U2113 (N_2113,N_1599,N_1549);
nor U2114 (N_2114,N_1953,N_1376);
nor U2115 (N_2115,N_1944,N_1809);
or U2116 (N_2116,N_1467,N_1203);
or U2117 (N_2117,N_1507,N_1419);
nor U2118 (N_2118,N_1096,N_1803);
nand U2119 (N_2119,N_1114,N_1524);
nor U2120 (N_2120,N_1000,N_1767);
nand U2121 (N_2121,N_1700,N_1528);
or U2122 (N_2122,N_1958,N_1518);
or U2123 (N_2123,N_1020,N_1563);
and U2124 (N_2124,N_1141,N_1854);
nand U2125 (N_2125,N_1643,N_1272);
or U2126 (N_2126,N_1875,N_1302);
or U2127 (N_2127,N_1457,N_1342);
and U2128 (N_2128,N_1370,N_1309);
nand U2129 (N_2129,N_1564,N_1940);
nand U2130 (N_2130,N_1093,N_1713);
nand U2131 (N_2131,N_1598,N_1845);
nand U2132 (N_2132,N_1615,N_1894);
xor U2133 (N_2133,N_1380,N_1650);
nor U2134 (N_2134,N_1621,N_1781);
or U2135 (N_2135,N_1195,N_1102);
nand U2136 (N_2136,N_1900,N_1997);
nor U2137 (N_2137,N_1234,N_1668);
and U2138 (N_2138,N_1751,N_1073);
and U2139 (N_2139,N_1133,N_1805);
nor U2140 (N_2140,N_1464,N_1052);
and U2141 (N_2141,N_1233,N_1672);
nand U2142 (N_2142,N_1682,N_1965);
and U2143 (N_2143,N_1649,N_1592);
and U2144 (N_2144,N_1131,N_1796);
nor U2145 (N_2145,N_1766,N_1231);
xor U2146 (N_2146,N_1374,N_1490);
or U2147 (N_2147,N_1627,N_1398);
or U2148 (N_2148,N_1579,N_1974);
or U2149 (N_2149,N_1748,N_1852);
xor U2150 (N_2150,N_1437,N_1697);
or U2151 (N_2151,N_1945,N_1378);
and U2152 (N_2152,N_1626,N_1088);
nor U2153 (N_2153,N_1060,N_1813);
xnor U2154 (N_2154,N_1596,N_1879);
xor U2155 (N_2155,N_1551,N_1613);
or U2156 (N_2156,N_1415,N_1581);
or U2157 (N_2157,N_1765,N_1371);
or U2158 (N_2158,N_1804,N_1624);
nor U2159 (N_2159,N_1916,N_1224);
nor U2160 (N_2160,N_1286,N_1531);
nand U2161 (N_2161,N_1602,N_1720);
nor U2162 (N_2162,N_1312,N_1667);
and U2163 (N_2163,N_1436,N_1934);
nor U2164 (N_2164,N_1880,N_1753);
nor U2165 (N_2165,N_1499,N_1608);
xnor U2166 (N_2166,N_1080,N_1305);
and U2167 (N_2167,N_1434,N_1815);
nand U2168 (N_2168,N_1698,N_1976);
nor U2169 (N_2169,N_1973,N_1883);
and U2170 (N_2170,N_1607,N_1381);
nand U2171 (N_2171,N_1795,N_1618);
and U2172 (N_2172,N_1308,N_1868);
nor U2173 (N_2173,N_1984,N_1174);
or U2174 (N_2174,N_1794,N_1201);
nand U2175 (N_2175,N_1410,N_1433);
nor U2176 (N_2176,N_1632,N_1511);
nand U2177 (N_2177,N_1369,N_1450);
or U2178 (N_2178,N_1737,N_1924);
xor U2179 (N_2179,N_1315,N_1829);
nand U2180 (N_2180,N_1249,N_1092);
nand U2181 (N_2181,N_1448,N_1055);
or U2182 (N_2182,N_1688,N_1439);
or U2183 (N_2183,N_1193,N_1601);
xor U2184 (N_2184,N_1162,N_1362);
or U2185 (N_2185,N_1614,N_1843);
nor U2186 (N_2186,N_1786,N_1273);
nand U2187 (N_2187,N_1027,N_1285);
or U2188 (N_2188,N_1379,N_1861);
or U2189 (N_2189,N_1107,N_1675);
or U2190 (N_2190,N_1982,N_1530);
nand U2191 (N_2191,N_1903,N_1557);
or U2192 (N_2192,N_1801,N_1319);
nand U2193 (N_2193,N_1094,N_1860);
xor U2194 (N_2194,N_1771,N_1853);
nand U2195 (N_2195,N_1635,N_1502);
nand U2196 (N_2196,N_1578,N_1017);
and U2197 (N_2197,N_1764,N_1194);
and U2198 (N_2198,N_1773,N_1267);
nor U2199 (N_2199,N_1744,N_1138);
and U2200 (N_2200,N_1685,N_1812);
nand U2201 (N_2201,N_1081,N_1474);
and U2202 (N_2202,N_1429,N_1015);
nand U2203 (N_2203,N_1749,N_1012);
xnor U2204 (N_2204,N_1481,N_1639);
or U2205 (N_2205,N_1119,N_1059);
nand U2206 (N_2206,N_1588,N_1045);
nand U2207 (N_2207,N_1992,N_1594);
or U2208 (N_2208,N_1562,N_1583);
and U2209 (N_2209,N_1401,N_1157);
and U2210 (N_2210,N_1345,N_1418);
nand U2211 (N_2211,N_1996,N_1556);
or U2212 (N_2212,N_1078,N_1116);
xor U2213 (N_2213,N_1559,N_1560);
or U2214 (N_2214,N_1320,N_1510);
nand U2215 (N_2215,N_1128,N_1109);
or U2216 (N_2216,N_1640,N_1127);
and U2217 (N_2217,N_1790,N_1349);
or U2218 (N_2218,N_1258,N_1168);
nand U2219 (N_2219,N_1789,N_1471);
and U2220 (N_2220,N_1251,N_1508);
nand U2221 (N_2221,N_1963,N_1955);
nor U2222 (N_2222,N_1754,N_1930);
and U2223 (N_2223,N_1068,N_1637);
and U2224 (N_2224,N_1653,N_1083);
or U2225 (N_2225,N_1120,N_1057);
nand U2226 (N_2226,N_1905,N_1509);
nor U2227 (N_2227,N_1904,N_1453);
and U2228 (N_2228,N_1028,N_1070);
and U2229 (N_2229,N_1048,N_1163);
nor U2230 (N_2230,N_1523,N_1095);
nand U2231 (N_2231,N_1501,N_1176);
and U2232 (N_2232,N_1225,N_1832);
nor U2233 (N_2233,N_1950,N_1318);
nor U2234 (N_2234,N_1420,N_1504);
and U2235 (N_2235,N_1023,N_1540);
nand U2236 (N_2236,N_1513,N_1164);
nor U2237 (N_2237,N_1255,N_1259);
or U2238 (N_2238,N_1844,N_1907);
nand U2239 (N_2239,N_1515,N_1405);
or U2240 (N_2240,N_1780,N_1185);
nand U2241 (N_2241,N_1597,N_1254);
nand U2242 (N_2242,N_1711,N_1889);
nand U2243 (N_2243,N_1756,N_1221);
or U2244 (N_2244,N_1049,N_1031);
nand U2245 (N_2245,N_1561,N_1099);
or U2246 (N_2246,N_1011,N_1262);
nor U2247 (N_2247,N_1352,N_1689);
and U2248 (N_2248,N_1145,N_1871);
nand U2249 (N_2249,N_1856,N_1926);
nor U2250 (N_2250,N_1503,N_1665);
nand U2251 (N_2251,N_1483,N_1460);
nand U2252 (N_2252,N_1043,N_1189);
nand U2253 (N_2253,N_1008,N_1399);
xor U2254 (N_2254,N_1864,N_1553);
or U2255 (N_2255,N_1687,N_1358);
or U2256 (N_2256,N_1962,N_1304);
and U2257 (N_2257,N_1927,N_1659);
or U2258 (N_2258,N_1881,N_1517);
nor U2259 (N_2259,N_1799,N_1541);
nor U2260 (N_2260,N_1006,N_1187);
or U2261 (N_2261,N_1196,N_1351);
nand U2262 (N_2262,N_1683,N_1686);
nand U2263 (N_2263,N_1539,N_1938);
nor U2264 (N_2264,N_1256,N_1575);
xor U2265 (N_2265,N_1629,N_1291);
nor U2266 (N_2266,N_1154,N_1293);
nand U2267 (N_2267,N_1445,N_1032);
or U2268 (N_2268,N_1489,N_1359);
and U2269 (N_2269,N_1910,N_1505);
nor U2270 (N_2270,N_1775,N_1177);
nor U2271 (N_2271,N_1806,N_1215);
or U2272 (N_2272,N_1933,N_1086);
xor U2273 (N_2273,N_1816,N_1617);
nor U2274 (N_2274,N_1527,N_1660);
xnor U2275 (N_2275,N_1703,N_1662);
nor U2276 (N_2276,N_1733,N_1873);
nor U2277 (N_2277,N_1067,N_1280);
or U2278 (N_2278,N_1758,N_1300);
or U2279 (N_2279,N_1642,N_1986);
or U2280 (N_2280,N_1555,N_1229);
and U2281 (N_2281,N_1360,N_1661);
nand U2282 (N_2282,N_1545,N_1181);
and U2283 (N_2283,N_1014,N_1750);
and U2284 (N_2284,N_1535,N_1747);
nand U2285 (N_2285,N_1834,N_1819);
and U2286 (N_2286,N_1423,N_1869);
or U2287 (N_2287,N_1993,N_1529);
nor U2288 (N_2288,N_1484,N_1995);
or U2289 (N_2289,N_1783,N_1072);
and U2290 (N_2290,N_1329,N_1646);
or U2291 (N_2291,N_1666,N_1339);
or U2292 (N_2292,N_1676,N_1334);
xnor U2293 (N_2293,N_1915,N_1777);
and U2294 (N_2294,N_1322,N_1021);
or U2295 (N_2295,N_1392,N_1257);
nand U2296 (N_2296,N_1153,N_1851);
nor U2297 (N_2297,N_1939,N_1230);
and U2298 (N_2298,N_1406,N_1026);
and U2299 (N_2299,N_1179,N_1901);
nor U2300 (N_2300,N_1636,N_1317);
nor U2301 (N_2301,N_1402,N_1161);
and U2302 (N_2302,N_1867,N_1935);
nand U2303 (N_2303,N_1395,N_1393);
and U2304 (N_2304,N_1327,N_1943);
and U2305 (N_2305,N_1872,N_1892);
and U2306 (N_2306,N_1244,N_1409);
and U2307 (N_2307,N_1447,N_1472);
and U2308 (N_2308,N_1839,N_1348);
nand U2309 (N_2309,N_1292,N_1324);
nand U2310 (N_2310,N_1207,N_1811);
nand U2311 (N_2311,N_1357,N_1914);
nand U2312 (N_2312,N_1002,N_1774);
xnor U2313 (N_2313,N_1886,N_1030);
and U2314 (N_2314,N_1707,N_1887);
nand U2315 (N_2315,N_1408,N_1054);
xor U2316 (N_2316,N_1323,N_1307);
and U2317 (N_2317,N_1695,N_1546);
xnor U2318 (N_2318,N_1140,N_1792);
xnor U2319 (N_2319,N_1010,N_1544);
and U2320 (N_2320,N_1928,N_1480);
nand U2321 (N_2321,N_1919,N_1029);
and U2322 (N_2322,N_1485,N_1647);
or U2323 (N_2323,N_1922,N_1912);
and U2324 (N_2324,N_1038,N_1651);
xor U2325 (N_2325,N_1743,N_1478);
or U2326 (N_2326,N_1604,N_1514);
nor U2327 (N_2327,N_1739,N_1287);
nand U2328 (N_2328,N_1018,N_1574);
or U2329 (N_2329,N_1572,N_1053);
or U2330 (N_2330,N_1909,N_1722);
nand U2331 (N_2331,N_1442,N_1158);
and U2332 (N_2332,N_1670,N_1619);
xnor U2333 (N_2333,N_1746,N_1130);
nand U2334 (N_2334,N_1825,N_1736);
nand U2335 (N_2335,N_1730,N_1178);
nor U2336 (N_2336,N_1797,N_1966);
xor U2337 (N_2337,N_1582,N_1742);
and U2338 (N_2338,N_1208,N_1681);
and U2339 (N_2339,N_1718,N_1372);
nand U2340 (N_2340,N_1269,N_1009);
and U2341 (N_2341,N_1160,N_1264);
nor U2342 (N_2342,N_1146,N_1724);
nand U2343 (N_2343,N_1778,N_1897);
xnor U2344 (N_2344,N_1644,N_1353);
nor U2345 (N_2345,N_1473,N_1482);
and U2346 (N_2346,N_1363,N_1663);
or U2347 (N_2347,N_1533,N_1321);
nor U2348 (N_2348,N_1657,N_1622);
and U2349 (N_2349,N_1712,N_1979);
nand U2350 (N_2350,N_1350,N_1281);
or U2351 (N_2351,N_1956,N_1866);
or U2352 (N_2352,N_1908,N_1587);
or U2353 (N_2353,N_1823,N_1701);
nor U2354 (N_2354,N_1278,N_1656);
or U2355 (N_2355,N_1172,N_1271);
nor U2356 (N_2356,N_1696,N_1355);
xor U2357 (N_2357,N_1016,N_1200);
nand U2358 (N_2358,N_1734,N_1475);
or U2359 (N_2359,N_1959,N_1568);
or U2360 (N_2360,N_1235,N_1056);
nand U2361 (N_2361,N_1451,N_1136);
nor U2362 (N_2362,N_1385,N_1103);
and U2363 (N_2363,N_1763,N_1785);
or U2364 (N_2364,N_1988,N_1266);
nand U2365 (N_2365,N_1223,N_1186);
nor U2366 (N_2366,N_1276,N_1137);
nand U2367 (N_2367,N_1630,N_1782);
and U2368 (N_2368,N_1570,N_1407);
and U2369 (N_2369,N_1791,N_1113);
or U2370 (N_2370,N_1025,N_1990);
xnor U2371 (N_2371,N_1705,N_1603);
or U2372 (N_2372,N_1768,N_1463);
nand U2373 (N_2373,N_1034,N_1972);
nor U2374 (N_2374,N_1400,N_1294);
and U2375 (N_2375,N_1090,N_1165);
nand U2376 (N_2376,N_1740,N_1738);
nor U2377 (N_2377,N_1547,N_1337);
and U2378 (N_2378,N_1857,N_1003);
nor U2379 (N_2379,N_1227,N_1330);
nor U2380 (N_2380,N_1386,N_1893);
and U2381 (N_2381,N_1784,N_1242);
and U2382 (N_2382,N_1268,N_1704);
or U2383 (N_2383,N_1850,N_1542);
nand U2384 (N_2384,N_1336,N_1929);
and U2385 (N_2385,N_1807,N_1325);
or U2386 (N_2386,N_1456,N_1237);
or U2387 (N_2387,N_1274,N_1937);
nand U2388 (N_2388,N_1998,N_1139);
or U2389 (N_2389,N_1802,N_1206);
or U2390 (N_2390,N_1942,N_1462);
nand U2391 (N_2391,N_1122,N_1388);
nand U2392 (N_2392,N_1567,N_1283);
and U2393 (N_2393,N_1469,N_1978);
or U2394 (N_2394,N_1190,N_1074);
or U2395 (N_2395,N_1772,N_1521);
nor U2396 (N_2396,N_1987,N_1123);
nand U2397 (N_2397,N_1818,N_1757);
and U2398 (N_2398,N_1169,N_1062);
and U2399 (N_2399,N_1431,N_1888);
or U2400 (N_2400,N_1715,N_1338);
and U2401 (N_2401,N_1188,N_1779);
nand U2402 (N_2402,N_1446,N_1590);
and U2403 (N_2403,N_1776,N_1580);
or U2404 (N_2404,N_1443,N_1906);
and U2405 (N_2405,N_1655,N_1896);
or U2406 (N_2406,N_1151,N_1769);
nor U2407 (N_2407,N_1732,N_1787);
and U2408 (N_2408,N_1197,N_1129);
nand U2409 (N_2409,N_1344,N_1051);
nand U2410 (N_2410,N_1373,N_1822);
nand U2411 (N_2411,N_1211,N_1192);
or U2412 (N_2412,N_1522,N_1332);
or U2413 (N_2413,N_1427,N_1536);
or U2414 (N_2414,N_1440,N_1623);
and U2415 (N_2415,N_1007,N_1082);
and U2416 (N_2416,N_1525,N_1612);
nor U2417 (N_2417,N_1444,N_1346);
xor U2418 (N_2418,N_1616,N_1708);
or U2419 (N_2419,N_1714,N_1296);
or U2420 (N_2420,N_1039,N_1282);
xnor U2421 (N_2421,N_1593,N_1275);
nor U2422 (N_2422,N_1239,N_1091);
nand U2423 (N_2423,N_1611,N_1333);
and U2424 (N_2424,N_1170,N_1299);
and U2425 (N_2425,N_1487,N_1971);
or U2426 (N_2426,N_1222,N_1397);
nand U2427 (N_2427,N_1952,N_1064);
or U2428 (N_2428,N_1265,N_1674);
nand U2429 (N_2429,N_1865,N_1297);
nand U2430 (N_2430,N_1328,N_1983);
nand U2431 (N_2431,N_1970,N_1980);
nor U2432 (N_2432,N_1183,N_1917);
or U2433 (N_2433,N_1077,N_1512);
or U2434 (N_2434,N_1576,N_1793);
nand U2435 (N_2435,N_1702,N_1585);
nand U2436 (N_2436,N_1246,N_1155);
and U2437 (N_2437,N_1584,N_1633);
nand U2438 (N_2438,N_1335,N_1403);
or U2439 (N_2439,N_1066,N_1961);
xnor U2440 (N_2440,N_1301,N_1425);
and U2441 (N_2441,N_1001,N_1735);
and U2442 (N_2442,N_1532,N_1217);
nor U2443 (N_2443,N_1210,N_1213);
or U2444 (N_2444,N_1205,N_1389);
and U2445 (N_2445,N_1104,N_1071);
xnor U2446 (N_2446,N_1037,N_1573);
and U2447 (N_2447,N_1895,N_1313);
nand U2448 (N_2448,N_1710,N_1365);
or U2449 (N_2449,N_1430,N_1050);
and U2450 (N_2450,N_1654,N_1716);
nor U2451 (N_2451,N_1589,N_1279);
nor U2452 (N_2452,N_1706,N_1413);
nand U2453 (N_2453,N_1152,N_1731);
nor U2454 (N_2454,N_1836,N_1310);
and U2455 (N_2455,N_1459,N_1526);
nand U2456 (N_2456,N_1143,N_1387);
or U2457 (N_2457,N_1340,N_1035);
nand U2458 (N_2458,N_1949,N_1946);
and U2459 (N_2459,N_1126,N_1638);
nor U2460 (N_2460,N_1673,N_1810);
or U2461 (N_2461,N_1175,N_1180);
nor U2462 (N_2462,N_1069,N_1438);
and U2463 (N_2463,N_1046,N_1316);
nor U2464 (N_2464,N_1931,N_1921);
nor U2465 (N_2465,N_1209,N_1247);
xnor U2466 (N_2466,N_1079,N_1760);
nand U2467 (N_2467,N_1920,N_1817);
nor U2468 (N_2468,N_1936,N_1452);
nand U2469 (N_2469,N_1634,N_1202);
and U2470 (N_2470,N_1913,N_1500);
or U2471 (N_2471,N_1364,N_1112);
or U2472 (N_2472,N_1306,N_1394);
nand U2473 (N_2473,N_1232,N_1985);
and U2474 (N_2474,N_1421,N_1923);
nor U2475 (N_2475,N_1167,N_1826);
nor U2476 (N_2476,N_1166,N_1841);
nand U2477 (N_2477,N_1125,N_1964);
nor U2478 (N_2478,N_1847,N_1755);
xnor U2479 (N_2479,N_1719,N_1314);
nand U2480 (N_2480,N_1218,N_1831);
nand U2481 (N_2481,N_1424,N_1960);
nor U2482 (N_2482,N_1814,N_1022);
and U2483 (N_2483,N_1994,N_1849);
nand U2484 (N_2484,N_1728,N_1115);
nand U2485 (N_2485,N_1691,N_1004);
nor U2486 (N_2486,N_1042,N_1245);
and U2487 (N_2487,N_1063,N_1085);
xor U2488 (N_2488,N_1347,N_1150);
nand U2489 (N_2489,N_1820,N_1240);
nor U2490 (N_2490,N_1729,N_1356);
and U2491 (N_2491,N_1858,N_1416);
xor U2492 (N_2492,N_1428,N_1290);
nor U2493 (N_2493,N_1677,N_1289);
nand U2494 (N_2494,N_1216,N_1679);
nand U2495 (N_2495,N_1044,N_1543);
nor U2496 (N_2496,N_1098,N_1476);
or U2497 (N_2497,N_1709,N_1226);
nor U2498 (N_2498,N_1620,N_1658);
or U2499 (N_2499,N_1721,N_1058);
and U2500 (N_2500,N_1824,N_1847);
and U2501 (N_2501,N_1373,N_1029);
nor U2502 (N_2502,N_1135,N_1094);
and U2503 (N_2503,N_1873,N_1144);
nand U2504 (N_2504,N_1301,N_1498);
and U2505 (N_2505,N_1235,N_1124);
and U2506 (N_2506,N_1415,N_1395);
nor U2507 (N_2507,N_1456,N_1309);
xnor U2508 (N_2508,N_1185,N_1449);
nand U2509 (N_2509,N_1942,N_1649);
nor U2510 (N_2510,N_1651,N_1869);
nor U2511 (N_2511,N_1738,N_1442);
nor U2512 (N_2512,N_1855,N_1367);
and U2513 (N_2513,N_1639,N_1468);
or U2514 (N_2514,N_1594,N_1651);
nand U2515 (N_2515,N_1049,N_1972);
and U2516 (N_2516,N_1550,N_1336);
and U2517 (N_2517,N_1351,N_1117);
nor U2518 (N_2518,N_1119,N_1127);
nand U2519 (N_2519,N_1816,N_1513);
xor U2520 (N_2520,N_1040,N_1570);
nor U2521 (N_2521,N_1891,N_1418);
and U2522 (N_2522,N_1015,N_1501);
nor U2523 (N_2523,N_1064,N_1218);
nor U2524 (N_2524,N_1015,N_1621);
xnor U2525 (N_2525,N_1421,N_1502);
nand U2526 (N_2526,N_1307,N_1436);
nand U2527 (N_2527,N_1780,N_1357);
xnor U2528 (N_2528,N_1512,N_1462);
nand U2529 (N_2529,N_1736,N_1184);
nor U2530 (N_2530,N_1026,N_1387);
nor U2531 (N_2531,N_1965,N_1638);
and U2532 (N_2532,N_1886,N_1239);
xnor U2533 (N_2533,N_1189,N_1695);
nor U2534 (N_2534,N_1238,N_1014);
nand U2535 (N_2535,N_1376,N_1381);
nor U2536 (N_2536,N_1171,N_1013);
xnor U2537 (N_2537,N_1485,N_1228);
nand U2538 (N_2538,N_1489,N_1864);
or U2539 (N_2539,N_1700,N_1451);
nor U2540 (N_2540,N_1994,N_1632);
nor U2541 (N_2541,N_1554,N_1849);
and U2542 (N_2542,N_1537,N_1464);
nor U2543 (N_2543,N_1331,N_1134);
nand U2544 (N_2544,N_1998,N_1069);
xnor U2545 (N_2545,N_1204,N_1009);
nand U2546 (N_2546,N_1672,N_1842);
or U2547 (N_2547,N_1595,N_1161);
or U2548 (N_2548,N_1887,N_1849);
and U2549 (N_2549,N_1065,N_1632);
nand U2550 (N_2550,N_1840,N_1036);
and U2551 (N_2551,N_1540,N_1013);
and U2552 (N_2552,N_1503,N_1477);
nor U2553 (N_2553,N_1183,N_1441);
nor U2554 (N_2554,N_1956,N_1269);
and U2555 (N_2555,N_1380,N_1715);
nor U2556 (N_2556,N_1925,N_1860);
and U2557 (N_2557,N_1821,N_1836);
and U2558 (N_2558,N_1878,N_1455);
and U2559 (N_2559,N_1940,N_1328);
and U2560 (N_2560,N_1124,N_1098);
xnor U2561 (N_2561,N_1193,N_1239);
xnor U2562 (N_2562,N_1754,N_1994);
nand U2563 (N_2563,N_1287,N_1973);
nor U2564 (N_2564,N_1817,N_1219);
and U2565 (N_2565,N_1148,N_1794);
or U2566 (N_2566,N_1059,N_1071);
or U2567 (N_2567,N_1045,N_1031);
or U2568 (N_2568,N_1884,N_1542);
nand U2569 (N_2569,N_1798,N_1839);
or U2570 (N_2570,N_1024,N_1974);
xor U2571 (N_2571,N_1174,N_1456);
nand U2572 (N_2572,N_1149,N_1887);
or U2573 (N_2573,N_1589,N_1094);
xnor U2574 (N_2574,N_1774,N_1854);
or U2575 (N_2575,N_1764,N_1071);
nor U2576 (N_2576,N_1825,N_1217);
or U2577 (N_2577,N_1683,N_1737);
and U2578 (N_2578,N_1004,N_1176);
nor U2579 (N_2579,N_1038,N_1252);
nor U2580 (N_2580,N_1084,N_1711);
nand U2581 (N_2581,N_1516,N_1866);
nor U2582 (N_2582,N_1660,N_1024);
nand U2583 (N_2583,N_1875,N_1481);
or U2584 (N_2584,N_1120,N_1502);
nor U2585 (N_2585,N_1230,N_1583);
nand U2586 (N_2586,N_1915,N_1207);
nand U2587 (N_2587,N_1671,N_1814);
and U2588 (N_2588,N_1191,N_1737);
xnor U2589 (N_2589,N_1389,N_1871);
nor U2590 (N_2590,N_1817,N_1261);
or U2591 (N_2591,N_1824,N_1474);
and U2592 (N_2592,N_1406,N_1699);
nand U2593 (N_2593,N_1508,N_1710);
nand U2594 (N_2594,N_1592,N_1961);
nand U2595 (N_2595,N_1507,N_1019);
and U2596 (N_2596,N_1427,N_1399);
and U2597 (N_2597,N_1268,N_1318);
nand U2598 (N_2598,N_1292,N_1707);
nor U2599 (N_2599,N_1490,N_1821);
nand U2600 (N_2600,N_1197,N_1641);
and U2601 (N_2601,N_1870,N_1517);
and U2602 (N_2602,N_1497,N_1391);
and U2603 (N_2603,N_1201,N_1733);
nand U2604 (N_2604,N_1071,N_1929);
nor U2605 (N_2605,N_1071,N_1088);
nand U2606 (N_2606,N_1323,N_1754);
and U2607 (N_2607,N_1904,N_1282);
nor U2608 (N_2608,N_1602,N_1289);
and U2609 (N_2609,N_1824,N_1720);
nand U2610 (N_2610,N_1031,N_1978);
or U2611 (N_2611,N_1454,N_1674);
nand U2612 (N_2612,N_1289,N_1878);
or U2613 (N_2613,N_1861,N_1746);
xor U2614 (N_2614,N_1919,N_1936);
nand U2615 (N_2615,N_1584,N_1512);
nand U2616 (N_2616,N_1844,N_1366);
nand U2617 (N_2617,N_1846,N_1153);
or U2618 (N_2618,N_1257,N_1743);
or U2619 (N_2619,N_1725,N_1289);
or U2620 (N_2620,N_1059,N_1565);
and U2621 (N_2621,N_1936,N_1018);
or U2622 (N_2622,N_1664,N_1302);
and U2623 (N_2623,N_1661,N_1338);
and U2624 (N_2624,N_1846,N_1892);
or U2625 (N_2625,N_1083,N_1679);
or U2626 (N_2626,N_1264,N_1204);
and U2627 (N_2627,N_1960,N_1600);
or U2628 (N_2628,N_1591,N_1618);
nor U2629 (N_2629,N_1299,N_1780);
xor U2630 (N_2630,N_1566,N_1792);
nor U2631 (N_2631,N_1005,N_1650);
xor U2632 (N_2632,N_1987,N_1695);
and U2633 (N_2633,N_1189,N_1036);
nor U2634 (N_2634,N_1615,N_1856);
nor U2635 (N_2635,N_1855,N_1033);
and U2636 (N_2636,N_1854,N_1153);
or U2637 (N_2637,N_1102,N_1280);
nand U2638 (N_2638,N_1967,N_1882);
nor U2639 (N_2639,N_1972,N_1756);
or U2640 (N_2640,N_1821,N_1319);
nand U2641 (N_2641,N_1338,N_1937);
or U2642 (N_2642,N_1466,N_1675);
or U2643 (N_2643,N_1490,N_1942);
nor U2644 (N_2644,N_1069,N_1056);
nor U2645 (N_2645,N_1695,N_1355);
xor U2646 (N_2646,N_1373,N_1685);
nand U2647 (N_2647,N_1495,N_1019);
and U2648 (N_2648,N_1908,N_1026);
nand U2649 (N_2649,N_1786,N_1340);
nand U2650 (N_2650,N_1049,N_1845);
nor U2651 (N_2651,N_1181,N_1883);
or U2652 (N_2652,N_1451,N_1406);
nand U2653 (N_2653,N_1645,N_1667);
nand U2654 (N_2654,N_1168,N_1613);
or U2655 (N_2655,N_1577,N_1178);
nand U2656 (N_2656,N_1424,N_1174);
nand U2657 (N_2657,N_1708,N_1317);
nand U2658 (N_2658,N_1162,N_1294);
nor U2659 (N_2659,N_1423,N_1891);
and U2660 (N_2660,N_1350,N_1876);
or U2661 (N_2661,N_1553,N_1397);
nand U2662 (N_2662,N_1342,N_1340);
or U2663 (N_2663,N_1832,N_1040);
or U2664 (N_2664,N_1414,N_1583);
and U2665 (N_2665,N_1330,N_1773);
nor U2666 (N_2666,N_1601,N_1666);
or U2667 (N_2667,N_1965,N_1486);
and U2668 (N_2668,N_1349,N_1655);
or U2669 (N_2669,N_1632,N_1414);
nand U2670 (N_2670,N_1938,N_1747);
and U2671 (N_2671,N_1899,N_1881);
nor U2672 (N_2672,N_1355,N_1194);
nor U2673 (N_2673,N_1144,N_1309);
or U2674 (N_2674,N_1954,N_1335);
nor U2675 (N_2675,N_1020,N_1375);
nor U2676 (N_2676,N_1126,N_1096);
nand U2677 (N_2677,N_1359,N_1029);
or U2678 (N_2678,N_1059,N_1852);
nand U2679 (N_2679,N_1461,N_1566);
and U2680 (N_2680,N_1397,N_1941);
nor U2681 (N_2681,N_1033,N_1716);
nor U2682 (N_2682,N_1426,N_1210);
nor U2683 (N_2683,N_1691,N_1834);
and U2684 (N_2684,N_1179,N_1743);
nand U2685 (N_2685,N_1285,N_1051);
and U2686 (N_2686,N_1775,N_1345);
nand U2687 (N_2687,N_1198,N_1534);
or U2688 (N_2688,N_1110,N_1118);
nor U2689 (N_2689,N_1999,N_1958);
or U2690 (N_2690,N_1026,N_1106);
nand U2691 (N_2691,N_1917,N_1230);
nand U2692 (N_2692,N_1454,N_1460);
and U2693 (N_2693,N_1436,N_1988);
nand U2694 (N_2694,N_1091,N_1056);
nand U2695 (N_2695,N_1333,N_1156);
and U2696 (N_2696,N_1325,N_1708);
or U2697 (N_2697,N_1152,N_1832);
nor U2698 (N_2698,N_1543,N_1681);
or U2699 (N_2699,N_1393,N_1535);
nor U2700 (N_2700,N_1159,N_1025);
and U2701 (N_2701,N_1204,N_1230);
nand U2702 (N_2702,N_1216,N_1071);
nand U2703 (N_2703,N_1119,N_1850);
or U2704 (N_2704,N_1220,N_1201);
and U2705 (N_2705,N_1470,N_1811);
or U2706 (N_2706,N_1608,N_1197);
or U2707 (N_2707,N_1419,N_1114);
nor U2708 (N_2708,N_1280,N_1335);
and U2709 (N_2709,N_1804,N_1435);
or U2710 (N_2710,N_1352,N_1326);
nor U2711 (N_2711,N_1253,N_1828);
nand U2712 (N_2712,N_1398,N_1385);
and U2713 (N_2713,N_1284,N_1789);
and U2714 (N_2714,N_1496,N_1369);
nor U2715 (N_2715,N_1855,N_1280);
nor U2716 (N_2716,N_1124,N_1643);
or U2717 (N_2717,N_1951,N_1962);
or U2718 (N_2718,N_1112,N_1664);
nor U2719 (N_2719,N_1142,N_1775);
nand U2720 (N_2720,N_1471,N_1586);
nor U2721 (N_2721,N_1476,N_1633);
or U2722 (N_2722,N_1962,N_1089);
or U2723 (N_2723,N_1607,N_1493);
or U2724 (N_2724,N_1024,N_1858);
nand U2725 (N_2725,N_1738,N_1170);
nand U2726 (N_2726,N_1281,N_1453);
and U2727 (N_2727,N_1826,N_1672);
nor U2728 (N_2728,N_1805,N_1406);
nor U2729 (N_2729,N_1541,N_1481);
and U2730 (N_2730,N_1871,N_1039);
nand U2731 (N_2731,N_1878,N_1214);
or U2732 (N_2732,N_1392,N_1885);
nor U2733 (N_2733,N_1388,N_1334);
nand U2734 (N_2734,N_1572,N_1594);
or U2735 (N_2735,N_1129,N_1887);
or U2736 (N_2736,N_1431,N_1448);
or U2737 (N_2737,N_1898,N_1505);
nand U2738 (N_2738,N_1350,N_1821);
xor U2739 (N_2739,N_1900,N_1347);
or U2740 (N_2740,N_1055,N_1833);
nand U2741 (N_2741,N_1174,N_1104);
or U2742 (N_2742,N_1130,N_1291);
or U2743 (N_2743,N_1019,N_1777);
and U2744 (N_2744,N_1566,N_1830);
nor U2745 (N_2745,N_1302,N_1286);
nor U2746 (N_2746,N_1050,N_1561);
nor U2747 (N_2747,N_1295,N_1533);
or U2748 (N_2748,N_1892,N_1093);
nor U2749 (N_2749,N_1006,N_1295);
or U2750 (N_2750,N_1230,N_1617);
nor U2751 (N_2751,N_1456,N_1976);
or U2752 (N_2752,N_1290,N_1867);
and U2753 (N_2753,N_1029,N_1710);
or U2754 (N_2754,N_1151,N_1090);
and U2755 (N_2755,N_1424,N_1573);
or U2756 (N_2756,N_1430,N_1258);
or U2757 (N_2757,N_1730,N_1616);
and U2758 (N_2758,N_1576,N_1201);
nand U2759 (N_2759,N_1639,N_1426);
nand U2760 (N_2760,N_1752,N_1691);
nor U2761 (N_2761,N_1393,N_1135);
nand U2762 (N_2762,N_1855,N_1602);
or U2763 (N_2763,N_1872,N_1177);
or U2764 (N_2764,N_1160,N_1038);
and U2765 (N_2765,N_1504,N_1460);
nor U2766 (N_2766,N_1381,N_1608);
and U2767 (N_2767,N_1510,N_1102);
and U2768 (N_2768,N_1253,N_1069);
xnor U2769 (N_2769,N_1237,N_1329);
xnor U2770 (N_2770,N_1564,N_1154);
nand U2771 (N_2771,N_1738,N_1332);
nor U2772 (N_2772,N_1388,N_1637);
or U2773 (N_2773,N_1101,N_1802);
and U2774 (N_2774,N_1608,N_1744);
or U2775 (N_2775,N_1867,N_1178);
or U2776 (N_2776,N_1223,N_1780);
and U2777 (N_2777,N_1864,N_1497);
or U2778 (N_2778,N_1294,N_1966);
xor U2779 (N_2779,N_1097,N_1290);
nor U2780 (N_2780,N_1022,N_1597);
nand U2781 (N_2781,N_1242,N_1983);
and U2782 (N_2782,N_1983,N_1410);
and U2783 (N_2783,N_1897,N_1968);
nor U2784 (N_2784,N_1898,N_1033);
nand U2785 (N_2785,N_1489,N_1398);
nor U2786 (N_2786,N_1911,N_1185);
nand U2787 (N_2787,N_1857,N_1416);
or U2788 (N_2788,N_1178,N_1222);
nor U2789 (N_2789,N_1790,N_1293);
or U2790 (N_2790,N_1918,N_1530);
xnor U2791 (N_2791,N_1502,N_1640);
xnor U2792 (N_2792,N_1467,N_1388);
nand U2793 (N_2793,N_1998,N_1375);
nor U2794 (N_2794,N_1037,N_1443);
and U2795 (N_2795,N_1470,N_1219);
xor U2796 (N_2796,N_1936,N_1883);
or U2797 (N_2797,N_1649,N_1409);
xor U2798 (N_2798,N_1925,N_1273);
nand U2799 (N_2799,N_1707,N_1800);
or U2800 (N_2800,N_1972,N_1697);
nor U2801 (N_2801,N_1708,N_1466);
nor U2802 (N_2802,N_1277,N_1396);
nand U2803 (N_2803,N_1174,N_1105);
and U2804 (N_2804,N_1396,N_1374);
and U2805 (N_2805,N_1849,N_1530);
or U2806 (N_2806,N_1102,N_1045);
nand U2807 (N_2807,N_1054,N_1987);
xnor U2808 (N_2808,N_1001,N_1482);
or U2809 (N_2809,N_1682,N_1117);
and U2810 (N_2810,N_1248,N_1518);
nand U2811 (N_2811,N_1382,N_1568);
or U2812 (N_2812,N_1749,N_1452);
nand U2813 (N_2813,N_1967,N_1264);
and U2814 (N_2814,N_1786,N_1861);
and U2815 (N_2815,N_1101,N_1569);
or U2816 (N_2816,N_1532,N_1861);
nand U2817 (N_2817,N_1785,N_1350);
and U2818 (N_2818,N_1882,N_1501);
and U2819 (N_2819,N_1705,N_1478);
or U2820 (N_2820,N_1899,N_1822);
and U2821 (N_2821,N_1253,N_1143);
nor U2822 (N_2822,N_1955,N_1841);
and U2823 (N_2823,N_1090,N_1718);
or U2824 (N_2824,N_1263,N_1630);
nand U2825 (N_2825,N_1513,N_1248);
or U2826 (N_2826,N_1812,N_1660);
nand U2827 (N_2827,N_1312,N_1491);
or U2828 (N_2828,N_1770,N_1798);
nand U2829 (N_2829,N_1013,N_1423);
nand U2830 (N_2830,N_1686,N_1455);
or U2831 (N_2831,N_1424,N_1719);
and U2832 (N_2832,N_1806,N_1544);
nor U2833 (N_2833,N_1854,N_1161);
or U2834 (N_2834,N_1925,N_1086);
nor U2835 (N_2835,N_1920,N_1391);
and U2836 (N_2836,N_1035,N_1066);
and U2837 (N_2837,N_1253,N_1610);
nand U2838 (N_2838,N_1844,N_1415);
nor U2839 (N_2839,N_1394,N_1703);
or U2840 (N_2840,N_1914,N_1082);
and U2841 (N_2841,N_1969,N_1783);
or U2842 (N_2842,N_1793,N_1438);
nand U2843 (N_2843,N_1468,N_1647);
nand U2844 (N_2844,N_1712,N_1749);
xor U2845 (N_2845,N_1105,N_1122);
xor U2846 (N_2846,N_1040,N_1619);
nor U2847 (N_2847,N_1899,N_1944);
nand U2848 (N_2848,N_1779,N_1385);
nand U2849 (N_2849,N_1118,N_1926);
and U2850 (N_2850,N_1497,N_1265);
or U2851 (N_2851,N_1269,N_1317);
and U2852 (N_2852,N_1440,N_1007);
nand U2853 (N_2853,N_1759,N_1386);
nor U2854 (N_2854,N_1599,N_1979);
and U2855 (N_2855,N_1066,N_1644);
xor U2856 (N_2856,N_1008,N_1451);
or U2857 (N_2857,N_1695,N_1660);
nand U2858 (N_2858,N_1923,N_1579);
and U2859 (N_2859,N_1921,N_1697);
nor U2860 (N_2860,N_1708,N_1414);
nor U2861 (N_2861,N_1399,N_1813);
xnor U2862 (N_2862,N_1582,N_1338);
or U2863 (N_2863,N_1017,N_1173);
nor U2864 (N_2864,N_1617,N_1090);
and U2865 (N_2865,N_1145,N_1920);
or U2866 (N_2866,N_1255,N_1293);
and U2867 (N_2867,N_1345,N_1321);
or U2868 (N_2868,N_1093,N_1198);
and U2869 (N_2869,N_1585,N_1221);
nor U2870 (N_2870,N_1371,N_1920);
or U2871 (N_2871,N_1072,N_1069);
xnor U2872 (N_2872,N_1084,N_1344);
nor U2873 (N_2873,N_1551,N_1939);
xor U2874 (N_2874,N_1176,N_1116);
or U2875 (N_2875,N_1185,N_1610);
and U2876 (N_2876,N_1763,N_1277);
or U2877 (N_2877,N_1007,N_1680);
nand U2878 (N_2878,N_1928,N_1312);
nor U2879 (N_2879,N_1556,N_1790);
or U2880 (N_2880,N_1177,N_1252);
nand U2881 (N_2881,N_1491,N_1090);
and U2882 (N_2882,N_1266,N_1511);
and U2883 (N_2883,N_1530,N_1850);
or U2884 (N_2884,N_1360,N_1269);
xnor U2885 (N_2885,N_1971,N_1622);
or U2886 (N_2886,N_1937,N_1035);
or U2887 (N_2887,N_1620,N_1105);
nor U2888 (N_2888,N_1383,N_1961);
or U2889 (N_2889,N_1914,N_1750);
nand U2890 (N_2890,N_1343,N_1079);
nor U2891 (N_2891,N_1311,N_1162);
and U2892 (N_2892,N_1032,N_1619);
and U2893 (N_2893,N_1409,N_1603);
xor U2894 (N_2894,N_1565,N_1794);
nor U2895 (N_2895,N_1136,N_1770);
or U2896 (N_2896,N_1556,N_1647);
and U2897 (N_2897,N_1991,N_1740);
or U2898 (N_2898,N_1780,N_1186);
nand U2899 (N_2899,N_1049,N_1588);
nand U2900 (N_2900,N_1492,N_1888);
and U2901 (N_2901,N_1322,N_1986);
nor U2902 (N_2902,N_1249,N_1435);
and U2903 (N_2903,N_1799,N_1726);
nor U2904 (N_2904,N_1302,N_1794);
or U2905 (N_2905,N_1691,N_1810);
or U2906 (N_2906,N_1380,N_1084);
or U2907 (N_2907,N_1252,N_1622);
or U2908 (N_2908,N_1251,N_1540);
or U2909 (N_2909,N_1987,N_1653);
nor U2910 (N_2910,N_1112,N_1261);
nand U2911 (N_2911,N_1186,N_1163);
or U2912 (N_2912,N_1226,N_1356);
nand U2913 (N_2913,N_1779,N_1937);
nor U2914 (N_2914,N_1256,N_1553);
or U2915 (N_2915,N_1465,N_1220);
or U2916 (N_2916,N_1411,N_1973);
or U2917 (N_2917,N_1209,N_1116);
and U2918 (N_2918,N_1973,N_1398);
nor U2919 (N_2919,N_1715,N_1248);
nor U2920 (N_2920,N_1527,N_1810);
and U2921 (N_2921,N_1466,N_1540);
nor U2922 (N_2922,N_1567,N_1580);
nand U2923 (N_2923,N_1235,N_1010);
xor U2924 (N_2924,N_1262,N_1296);
nand U2925 (N_2925,N_1420,N_1389);
or U2926 (N_2926,N_1986,N_1453);
and U2927 (N_2927,N_1961,N_1431);
and U2928 (N_2928,N_1193,N_1061);
and U2929 (N_2929,N_1818,N_1211);
or U2930 (N_2930,N_1226,N_1221);
nor U2931 (N_2931,N_1368,N_1585);
nand U2932 (N_2932,N_1830,N_1891);
xnor U2933 (N_2933,N_1164,N_1041);
nor U2934 (N_2934,N_1739,N_1136);
nand U2935 (N_2935,N_1729,N_1872);
nand U2936 (N_2936,N_1188,N_1033);
and U2937 (N_2937,N_1217,N_1856);
or U2938 (N_2938,N_1728,N_1833);
or U2939 (N_2939,N_1398,N_1476);
nor U2940 (N_2940,N_1262,N_1422);
and U2941 (N_2941,N_1931,N_1670);
or U2942 (N_2942,N_1653,N_1227);
or U2943 (N_2943,N_1062,N_1552);
and U2944 (N_2944,N_1853,N_1080);
nor U2945 (N_2945,N_1835,N_1171);
or U2946 (N_2946,N_1526,N_1617);
nand U2947 (N_2947,N_1274,N_1840);
and U2948 (N_2948,N_1571,N_1615);
nand U2949 (N_2949,N_1459,N_1325);
nand U2950 (N_2950,N_1646,N_1260);
nand U2951 (N_2951,N_1829,N_1373);
and U2952 (N_2952,N_1119,N_1140);
nor U2953 (N_2953,N_1740,N_1002);
xnor U2954 (N_2954,N_1681,N_1610);
or U2955 (N_2955,N_1089,N_1396);
nand U2956 (N_2956,N_1748,N_1496);
nand U2957 (N_2957,N_1805,N_1180);
and U2958 (N_2958,N_1325,N_1485);
and U2959 (N_2959,N_1487,N_1957);
or U2960 (N_2960,N_1605,N_1809);
nand U2961 (N_2961,N_1011,N_1741);
nand U2962 (N_2962,N_1087,N_1453);
or U2963 (N_2963,N_1026,N_1381);
nand U2964 (N_2964,N_1356,N_1162);
nand U2965 (N_2965,N_1149,N_1557);
nor U2966 (N_2966,N_1587,N_1944);
nand U2967 (N_2967,N_1311,N_1991);
nand U2968 (N_2968,N_1152,N_1604);
or U2969 (N_2969,N_1738,N_1179);
or U2970 (N_2970,N_1686,N_1179);
and U2971 (N_2971,N_1516,N_1941);
xnor U2972 (N_2972,N_1355,N_1292);
nor U2973 (N_2973,N_1981,N_1064);
nor U2974 (N_2974,N_1262,N_1940);
nor U2975 (N_2975,N_1936,N_1969);
nor U2976 (N_2976,N_1749,N_1694);
nand U2977 (N_2977,N_1427,N_1049);
and U2978 (N_2978,N_1015,N_1078);
or U2979 (N_2979,N_1776,N_1598);
and U2980 (N_2980,N_1521,N_1105);
nor U2981 (N_2981,N_1979,N_1751);
nor U2982 (N_2982,N_1005,N_1262);
and U2983 (N_2983,N_1454,N_1334);
xnor U2984 (N_2984,N_1843,N_1523);
nand U2985 (N_2985,N_1490,N_1486);
and U2986 (N_2986,N_1872,N_1877);
xnor U2987 (N_2987,N_1916,N_1319);
nor U2988 (N_2988,N_1025,N_1871);
nand U2989 (N_2989,N_1400,N_1507);
and U2990 (N_2990,N_1986,N_1267);
nor U2991 (N_2991,N_1379,N_1674);
nor U2992 (N_2992,N_1973,N_1650);
and U2993 (N_2993,N_1334,N_1655);
nor U2994 (N_2994,N_1949,N_1242);
and U2995 (N_2995,N_1740,N_1316);
nor U2996 (N_2996,N_1493,N_1902);
or U2997 (N_2997,N_1593,N_1310);
or U2998 (N_2998,N_1582,N_1241);
nand U2999 (N_2999,N_1478,N_1651);
and U3000 (N_3000,N_2613,N_2397);
and U3001 (N_3001,N_2718,N_2874);
nor U3002 (N_3002,N_2914,N_2941);
nor U3003 (N_3003,N_2125,N_2631);
nor U3004 (N_3004,N_2781,N_2357);
or U3005 (N_3005,N_2623,N_2383);
and U3006 (N_3006,N_2855,N_2198);
or U3007 (N_3007,N_2528,N_2949);
nor U3008 (N_3008,N_2745,N_2680);
nor U3009 (N_3009,N_2689,N_2759);
or U3010 (N_3010,N_2495,N_2346);
nor U3011 (N_3011,N_2318,N_2922);
xor U3012 (N_3012,N_2811,N_2575);
or U3013 (N_3013,N_2925,N_2684);
xor U3014 (N_3014,N_2656,N_2070);
nand U3015 (N_3015,N_2334,N_2446);
nand U3016 (N_3016,N_2124,N_2892);
and U3017 (N_3017,N_2886,N_2064);
and U3018 (N_3018,N_2821,N_2844);
nand U3019 (N_3019,N_2061,N_2907);
nor U3020 (N_3020,N_2433,N_2894);
nand U3021 (N_3021,N_2443,N_2931);
nor U3022 (N_3022,N_2839,N_2724);
nor U3023 (N_3023,N_2675,N_2521);
xnor U3024 (N_3024,N_2214,N_2598);
nand U3025 (N_3025,N_2592,N_2254);
xnor U3026 (N_3026,N_2002,N_2104);
and U3027 (N_3027,N_2135,N_2524);
and U3028 (N_3028,N_2935,N_2704);
and U3029 (N_3029,N_2976,N_2576);
nand U3030 (N_3030,N_2556,N_2748);
nand U3031 (N_3031,N_2022,N_2450);
or U3032 (N_3032,N_2175,N_2060);
xnor U3033 (N_3033,N_2978,N_2614);
or U3034 (N_3034,N_2234,N_2325);
or U3035 (N_3035,N_2414,N_2813);
nor U3036 (N_3036,N_2908,N_2226);
or U3037 (N_3037,N_2227,N_2469);
nor U3038 (N_3038,N_2764,N_2952);
or U3039 (N_3039,N_2785,N_2902);
or U3040 (N_3040,N_2452,N_2842);
or U3041 (N_3041,N_2906,N_2196);
and U3042 (N_3042,N_2496,N_2507);
and U3043 (N_3043,N_2557,N_2676);
nor U3044 (N_3044,N_2702,N_2158);
or U3045 (N_3045,N_2942,N_2281);
nor U3046 (N_3046,N_2585,N_2996);
nand U3047 (N_3047,N_2619,N_2426);
and U3048 (N_3048,N_2927,N_2462);
xor U3049 (N_3049,N_2787,N_2572);
nand U3050 (N_3050,N_2627,N_2683);
nor U3051 (N_3051,N_2869,N_2019);
and U3052 (N_3052,N_2622,N_2505);
xor U3053 (N_3053,N_2593,N_2312);
nand U3054 (N_3054,N_2531,N_2403);
nor U3055 (N_3055,N_2539,N_2330);
or U3056 (N_3056,N_2673,N_2932);
and U3057 (N_3057,N_2344,N_2999);
nor U3058 (N_3058,N_2968,N_2668);
nor U3059 (N_3059,N_2563,N_2177);
nor U3060 (N_3060,N_2962,N_2244);
or U3061 (N_3061,N_2895,N_2805);
or U3062 (N_3062,N_2584,N_2909);
or U3063 (N_3063,N_2766,N_2480);
and U3064 (N_3064,N_2100,N_2213);
or U3065 (N_3065,N_2231,N_2917);
nor U3066 (N_3066,N_2065,N_2834);
xnor U3067 (N_3067,N_2247,N_2295);
or U3068 (N_3068,N_2966,N_2694);
nand U3069 (N_3069,N_2473,N_2536);
or U3070 (N_3070,N_2690,N_2432);
and U3071 (N_3071,N_2845,N_2775);
xnor U3072 (N_3072,N_2406,N_2918);
nand U3073 (N_3073,N_2245,N_2195);
nand U3074 (N_3074,N_2977,N_2930);
or U3075 (N_3075,N_2385,N_2629);
nand U3076 (N_3076,N_2075,N_2970);
or U3077 (N_3077,N_2358,N_2736);
nand U3078 (N_3078,N_2508,N_2569);
and U3079 (N_3079,N_2985,N_2147);
and U3080 (N_3080,N_2487,N_2905);
or U3081 (N_3081,N_2898,N_2023);
xnor U3082 (N_3082,N_2589,N_2605);
or U3083 (N_3083,N_2550,N_2818);
and U3084 (N_3084,N_2677,N_2340);
or U3085 (N_3085,N_2415,N_2276);
or U3086 (N_3086,N_2581,N_2225);
nor U3087 (N_3087,N_2934,N_2936);
or U3088 (N_3088,N_2559,N_2519);
and U3089 (N_3089,N_2612,N_2848);
or U3090 (N_3090,N_2296,N_2482);
nand U3091 (N_3091,N_2392,N_2271);
nand U3092 (N_3092,N_2850,N_2355);
or U3093 (N_3093,N_2365,N_2756);
or U3094 (N_3094,N_2458,N_2826);
or U3095 (N_3095,N_2753,N_2875);
or U3096 (N_3096,N_2535,N_2882);
and U3097 (N_3097,N_2489,N_2719);
and U3098 (N_3098,N_2279,N_2698);
and U3099 (N_3099,N_2972,N_2001);
and U3100 (N_3100,N_2199,N_2721);
and U3101 (N_3101,N_2530,N_2049);
or U3102 (N_3102,N_2393,N_2747);
nor U3103 (N_3103,N_2373,N_2817);
nor U3104 (N_3104,N_2588,N_2161);
nand U3105 (N_3105,N_2693,N_2003);
xnor U3106 (N_3106,N_2143,N_2094);
and U3107 (N_3107,N_2448,N_2309);
nand U3108 (N_3108,N_2034,N_2411);
or U3109 (N_3109,N_2101,N_2464);
xor U3110 (N_3110,N_2933,N_2016);
nand U3111 (N_3111,N_2278,N_2425);
nand U3112 (N_3112,N_2682,N_2633);
or U3113 (N_3113,N_2568,N_2408);
nand U3114 (N_3114,N_2460,N_2144);
and U3115 (N_3115,N_2351,N_2995);
or U3116 (N_3116,N_2251,N_2709);
or U3117 (N_3117,N_2582,N_2797);
nor U3118 (N_3118,N_2802,N_2771);
nand U3119 (N_3119,N_2789,N_2072);
or U3120 (N_3120,N_2246,N_2730);
nand U3121 (N_3121,N_2692,N_2728);
xor U3122 (N_3122,N_2017,N_2549);
nor U3123 (N_3123,N_2428,N_2274);
and U3124 (N_3124,N_2218,N_2435);
or U3125 (N_3125,N_2722,N_2678);
or U3126 (N_3126,N_2504,N_2142);
or U3127 (N_3127,N_2674,N_2663);
or U3128 (N_3128,N_2066,N_2937);
xnor U3129 (N_3129,N_2751,N_2300);
nand U3130 (N_3130,N_2378,N_2434);
nor U3131 (N_3131,N_2777,N_2029);
or U3132 (N_3132,N_2595,N_2205);
nor U3133 (N_3133,N_2628,N_2329);
and U3134 (N_3134,N_2621,N_2288);
xnor U3135 (N_3135,N_2538,N_2043);
nor U3136 (N_3136,N_2243,N_2103);
and U3137 (N_3137,N_2824,N_2832);
nor U3138 (N_3138,N_2285,N_2252);
or U3139 (N_3139,N_2697,N_2294);
and U3140 (N_3140,N_2742,N_2599);
and U3141 (N_3141,N_2857,N_2222);
nand U3142 (N_3142,N_2794,N_2367);
nand U3143 (N_3143,N_2642,N_2041);
nor U3144 (N_3144,N_2963,N_2838);
or U3145 (N_3145,N_2345,N_2913);
nor U3146 (N_3146,N_2801,N_2547);
nand U3147 (N_3147,N_2988,N_2938);
xnor U3148 (N_3148,N_2980,N_2189);
or U3149 (N_3149,N_2455,N_2998);
and U3150 (N_3150,N_2302,N_2239);
nor U3151 (N_3151,N_2501,N_2961);
and U3152 (N_3152,N_2077,N_2868);
nand U3153 (N_3153,N_2308,N_2493);
nor U3154 (N_3154,N_2228,N_2743);
nor U3155 (N_3155,N_2282,N_2085);
or U3156 (N_3156,N_2200,N_2000);
or U3157 (N_3157,N_2497,N_2368);
nand U3158 (N_3158,N_2752,N_2151);
and U3159 (N_3159,N_2876,N_2732);
or U3160 (N_3160,N_2229,N_2384);
or U3161 (N_3161,N_2658,N_2639);
nand U3162 (N_3162,N_2040,N_2640);
nor U3163 (N_3163,N_2799,N_2184);
or U3164 (N_3164,N_2945,N_2780);
or U3165 (N_3165,N_2587,N_2140);
and U3166 (N_3166,N_2565,N_2873);
nand U3167 (N_3167,N_2871,N_2352);
or U3168 (N_3168,N_2989,N_2864);
or U3169 (N_3169,N_2526,N_2422);
nand U3170 (N_3170,N_2960,N_2790);
nor U3171 (N_3171,N_2207,N_2812);
and U3172 (N_3172,N_2560,N_2669);
and U3173 (N_3173,N_2417,N_2610);
nand U3174 (N_3174,N_2074,N_2632);
nand U3175 (N_3175,N_2044,N_2662);
nand U3176 (N_3176,N_2418,N_2471);
or U3177 (N_3177,N_2134,N_2518);
and U3178 (N_3178,N_2659,N_2242);
nor U3179 (N_3179,N_2891,N_2727);
or U3180 (N_3180,N_2139,N_2136);
or U3181 (N_3181,N_2903,N_2990);
or U3182 (N_3182,N_2843,N_2603);
and U3183 (N_3183,N_2160,N_2532);
nor U3184 (N_3184,N_2670,N_2087);
nor U3185 (N_3185,N_2374,N_2541);
xor U3186 (N_3186,N_2950,N_2884);
nor U3187 (N_3187,N_2354,N_2561);
nand U3188 (N_3188,N_2900,N_2091);
nand U3189 (N_3189,N_2401,N_2410);
xnor U3190 (N_3190,N_2080,N_2763);
and U3191 (N_3191,N_2203,N_2304);
nand U3192 (N_3192,N_2024,N_2258);
nand U3193 (N_3193,N_2007,N_2943);
nand U3194 (N_3194,N_2853,N_2131);
and U3195 (N_3195,N_2117,N_2264);
nor U3196 (N_3196,N_2110,N_2755);
nor U3197 (N_3197,N_2540,N_2808);
or U3198 (N_3198,N_2767,N_2267);
nand U3199 (N_3199,N_2310,N_2170);
nand U3200 (N_3200,N_2316,N_2154);
xor U3201 (N_3201,N_2716,N_2923);
nand U3202 (N_3202,N_2237,N_2904);
nor U3203 (N_3203,N_2638,N_2216);
xor U3204 (N_3204,N_2885,N_2498);
and U3205 (N_3205,N_2953,N_2653);
nand U3206 (N_3206,N_2293,N_2944);
or U3207 (N_3207,N_2825,N_2577);
xor U3208 (N_3208,N_2283,N_2940);
nor U3209 (N_3209,N_2277,N_2512);
nand U3210 (N_3210,N_2861,N_2375);
nor U3211 (N_3211,N_2706,N_2153);
or U3212 (N_3212,N_2607,N_2602);
nor U3213 (N_3213,N_2350,N_2037);
nand U3214 (N_3214,N_2798,N_2708);
or U3215 (N_3215,N_2109,N_2793);
nor U3216 (N_3216,N_2046,N_2510);
xnor U3217 (N_3217,N_2377,N_2888);
nor U3218 (N_3218,N_2533,N_2695);
xnor U3219 (N_3219,N_2899,N_2809);
xor U3220 (N_3220,N_2858,N_2849);
and U3221 (N_3221,N_2618,N_2955);
nor U3222 (N_3222,N_2356,N_2782);
or U3223 (N_3223,N_2646,N_2431);
or U3224 (N_3224,N_2167,N_2166);
and U3225 (N_3225,N_2219,N_2987);
xor U3226 (N_3226,N_2685,N_2454);
and U3227 (N_3227,N_2776,N_2475);
xor U3228 (N_3228,N_2067,N_2720);
xnor U3229 (N_3229,N_2055,N_2726);
and U3230 (N_3230,N_2652,N_2836);
or U3231 (N_3231,N_2847,N_2298);
nor U3232 (N_3232,N_2654,N_2820);
or U3233 (N_3233,N_2707,N_2947);
nor U3234 (N_3234,N_2113,N_2145);
or U3235 (N_3235,N_2339,N_2215);
nand U3236 (N_3236,N_2086,N_2118);
and U3237 (N_3237,N_2542,N_2926);
or U3238 (N_3238,N_2486,N_2725);
nand U3239 (N_3239,N_2097,N_2407);
nor U3240 (N_3240,N_2758,N_2290);
nor U3241 (N_3241,N_2047,N_2173);
xor U3242 (N_3242,N_2664,N_2974);
and U3243 (N_3243,N_2786,N_2106);
nor U3244 (N_3244,N_2341,N_2604);
or U3245 (N_3245,N_2901,N_2093);
and U3246 (N_3246,N_2833,N_2361);
nand U3247 (N_3247,N_2208,N_2197);
and U3248 (N_3248,N_2870,N_2039);
nor U3249 (N_3249,N_2359,N_2360);
nor U3250 (N_3250,N_2863,N_2171);
and U3251 (N_3251,N_2608,N_2620);
and U3252 (N_3252,N_2223,N_2624);
and U3253 (N_3253,N_2409,N_2430);
or U3254 (N_3254,N_2739,N_2399);
and U3255 (N_3255,N_2112,N_2691);
nand U3256 (N_3256,N_2583,N_2919);
or U3257 (N_3257,N_2212,N_2194);
and U3258 (N_3258,N_2650,N_2566);
nor U3259 (N_3259,N_2018,N_2567);
or U3260 (N_3260,N_2301,N_2911);
nor U3261 (N_3261,N_2564,N_2307);
nor U3262 (N_3262,N_2051,N_2461);
xnor U3263 (N_3263,N_2265,N_2703);
nor U3264 (N_3264,N_2823,N_2405);
xnor U3265 (N_3265,N_2262,N_2969);
and U3266 (N_3266,N_2157,N_2463);
xnor U3267 (N_3267,N_2474,N_2073);
nand U3268 (N_3268,N_2616,N_2322);
nor U3269 (N_3269,N_2983,N_2630);
nand U3270 (N_3270,N_2335,N_2026);
or U3271 (N_3271,N_2386,N_2590);
nand U3272 (N_3272,N_2317,N_2814);
or U3273 (N_3273,N_2313,N_2163);
and U3274 (N_3274,N_2444,N_2558);
nand U3275 (N_3275,N_2636,N_2159);
nor U3276 (N_3276,N_2773,N_2353);
or U3277 (N_3277,N_2879,N_2148);
and U3278 (N_3278,N_2079,N_2467);
nor U3279 (N_3279,N_2372,N_2829);
and U3280 (N_3280,N_2762,N_2068);
and U3281 (N_3281,N_2735,N_2394);
xor U3282 (N_3282,N_2058,N_2390);
nand U3283 (N_3283,N_2315,N_2439);
nand U3284 (N_3284,N_2164,N_2948);
and U3285 (N_3285,N_2544,N_2169);
nor U3286 (N_3286,N_2021,N_2421);
nand U3287 (N_3287,N_2500,N_2625);
and U3288 (N_3288,N_2027,N_2712);
xnor U3289 (N_3289,N_2248,N_2666);
nand U3290 (N_3290,N_2973,N_2032);
or U3291 (N_3291,N_2741,N_2445);
or U3292 (N_3292,N_2398,N_2319);
or U3293 (N_3293,N_2553,N_2562);
nand U3294 (N_3294,N_2116,N_2573);
nor U3295 (N_3295,N_2644,N_2520);
xnor U3296 (N_3296,N_2701,N_2641);
nand U3297 (N_3297,N_2715,N_2880);
and U3298 (N_3298,N_2548,N_2803);
or U3299 (N_3299,N_2362,N_2783);
or U3300 (N_3300,N_2438,N_2321);
and U3301 (N_3301,N_2182,N_2956);
xnor U3302 (N_3302,N_2483,N_2993);
nor U3303 (N_3303,N_2059,N_2511);
nor U3304 (N_3304,N_2738,N_2651);
or U3305 (N_3305,N_2297,N_2209);
nor U3306 (N_3306,N_2975,N_2889);
and U3307 (N_3307,N_2057,N_2178);
and U3308 (N_3308,N_2342,N_2806);
or U3309 (N_3309,N_2048,N_2615);
nand U3310 (N_3310,N_2015,N_2111);
and U3311 (N_3311,N_2141,N_2760);
or U3312 (N_3312,N_2854,N_2096);
nand U3313 (N_3313,N_2380,N_2671);
or U3314 (N_3314,N_2492,N_2009);
xor U3315 (N_3315,N_2946,N_2050);
nor U3316 (N_3316,N_2133,N_2366);
nor U3317 (N_3317,N_2082,N_2594);
nor U3318 (N_3318,N_2750,N_2071);
nand U3319 (N_3319,N_2069,N_2179);
or U3320 (N_3320,N_2083,N_2052);
xor U3321 (N_3321,N_2089,N_2757);
xnor U3322 (N_3322,N_2449,N_2025);
or U3323 (N_3323,N_2437,N_2191);
nand U3324 (N_3324,N_2490,N_2174);
nand U3325 (N_3325,N_2423,N_2115);
and U3326 (N_3326,N_2172,N_2273);
or U3327 (N_3327,N_2723,N_2201);
nand U3328 (N_3328,N_2447,N_2056);
nor U3329 (N_3329,N_2791,N_2081);
nor U3330 (N_3330,N_2700,N_2349);
or U3331 (N_3331,N_2146,N_2102);
xor U3332 (N_3332,N_2287,N_2600);
or U3333 (N_3333,N_2517,N_2261);
nor U3334 (N_3334,N_2872,N_2127);
xor U3335 (N_3335,N_2788,N_2749);
and U3336 (N_3336,N_2303,N_2617);
and U3337 (N_3337,N_2665,N_2570);
nand U3338 (N_3338,N_2688,N_2816);
or U3339 (N_3339,N_2921,N_2020);
xnor U3340 (N_3340,N_2867,N_2714);
or U3341 (N_3341,N_2328,N_2181);
or U3342 (N_3342,N_2597,N_2381);
and U3343 (N_3343,N_2859,N_2591);
nand U3344 (N_3344,N_2457,N_2660);
or U3345 (N_3345,N_2013,N_2466);
or U3346 (N_3346,N_2250,N_2571);
and U3347 (N_3347,N_2484,N_2442);
nand U3348 (N_3348,N_2233,N_2994);
nand U3349 (N_3349,N_2337,N_2982);
or U3350 (N_3350,N_2920,N_2655);
nand U3351 (N_3351,N_2130,N_2292);
nand U3352 (N_3352,N_2150,N_2388);
xor U3353 (N_3353,N_2132,N_2717);
nand U3354 (N_3354,N_2270,N_2054);
or U3355 (N_3355,N_2740,N_2552);
or U3356 (N_3356,N_2984,N_2031);
and U3357 (N_3357,N_2256,N_2126);
nand U3358 (N_3358,N_2796,N_2551);
nor U3359 (N_3359,N_2137,N_2778);
or U3360 (N_3360,N_2635,N_2515);
and U3361 (N_3361,N_2453,N_2795);
or U3362 (N_3362,N_2601,N_2611);
nand U3363 (N_3363,N_2865,N_2187);
or U3364 (N_3364,N_2259,N_2509);
or U3365 (N_3365,N_2860,N_2772);
xor U3366 (N_3366,N_2770,N_2331);
nor U3367 (N_3367,N_2815,N_2733);
or U3368 (N_3368,N_2221,N_2238);
or U3369 (N_3369,N_2107,N_2657);
xor U3370 (N_3370,N_2241,N_2371);
nand U3371 (N_3371,N_2291,N_2395);
nor U3372 (N_3372,N_2468,N_2958);
nand U3373 (N_3373,N_2912,N_2333);
or U3374 (N_3374,N_2729,N_2516);
nor U3375 (N_3375,N_2255,N_2606);
and U3376 (N_3376,N_2545,N_2681);
nor U3377 (N_3377,N_2327,N_2396);
and U3378 (N_3378,N_2416,N_2176);
or U3379 (N_3379,N_2578,N_2846);
xnor U3380 (N_3380,N_2138,N_2687);
xnor U3381 (N_3381,N_2128,N_2579);
nor U3382 (N_3382,N_2165,N_2004);
nand U3383 (N_3383,N_2014,N_2499);
or U3384 (N_3384,N_2376,N_2078);
or U3385 (N_3385,N_2090,N_2391);
and U3386 (N_3386,N_2710,N_2555);
nor U3387 (N_3387,N_2643,N_2705);
and U3388 (N_3388,N_2413,N_2284);
and U3389 (N_3389,N_2609,N_2476);
and U3390 (N_3390,N_2306,N_2971);
and U3391 (N_3391,N_2554,N_2045);
or U3392 (N_3392,N_2939,N_2035);
or U3393 (N_3393,N_2810,N_2204);
or U3394 (N_3394,N_2008,N_2964);
nor U3395 (N_3395,N_2456,N_2311);
nor U3396 (N_3396,N_2389,N_2099);
xor U3397 (N_3397,N_2230,N_2711);
nand U3398 (N_3398,N_2382,N_2180);
nand U3399 (N_3399,N_2765,N_2036);
nand U3400 (N_3400,N_2896,N_2831);
or U3401 (N_3401,N_2183,N_2011);
or U3402 (N_3402,N_2890,N_2929);
xnor U3403 (N_3403,N_2852,N_2866);
or U3404 (N_3404,N_2320,N_2830);
nor U3405 (N_3405,N_2686,N_2105);
nand U3406 (N_3406,N_2924,N_2525);
and U3407 (N_3407,N_2959,N_2667);
and U3408 (N_3408,N_2472,N_2451);
or U3409 (N_3409,N_2827,N_2586);
or U3410 (N_3410,N_2400,N_2897);
or U3411 (N_3411,N_2877,N_2835);
nand U3412 (N_3412,N_2063,N_2211);
and U3413 (N_3413,N_2746,N_2114);
nand U3414 (N_3414,N_2910,N_2272);
and U3415 (N_3415,N_2162,N_2030);
and U3416 (N_3416,N_2338,N_2465);
nor U3417 (N_3417,N_2263,N_2289);
or U3418 (N_3418,N_2120,N_2220);
nor U3419 (N_3419,N_2343,N_2095);
or U3420 (N_3420,N_2347,N_2420);
or U3421 (N_3421,N_2240,N_2062);
nand U3422 (N_3422,N_2928,N_2696);
nor U3423 (N_3423,N_2915,N_2186);
nor U3424 (N_3424,N_2440,N_2232);
or U3425 (N_3425,N_2485,N_2206);
nor U3426 (N_3426,N_2957,N_2774);
nand U3427 (N_3427,N_2991,N_2737);
nand U3428 (N_3428,N_2369,N_2076);
or U3429 (N_3429,N_2190,N_2266);
xor U3430 (N_3430,N_2280,N_2427);
nand U3431 (N_3431,N_2779,N_2807);
nor U3432 (N_3432,N_2479,N_2992);
nor U3433 (N_3433,N_2005,N_2862);
nor U3434 (N_3434,N_2537,N_2168);
and U3435 (N_3435,N_2012,N_2084);
nand U3436 (N_3436,N_2053,N_2580);
xnor U3437 (N_3437,N_2314,N_2543);
nand U3438 (N_3438,N_2481,N_2441);
nor U3439 (N_3439,N_2954,N_2477);
and U3440 (N_3440,N_2513,N_2332);
nand U3441 (N_3441,N_2503,N_2488);
and U3442 (N_3442,N_2412,N_2522);
nand U3443 (N_3443,N_2840,N_2149);
xnor U3444 (N_3444,N_2249,N_2878);
nand U3445 (N_3445,N_2260,N_2236);
xnor U3446 (N_3446,N_2965,N_2202);
nor U3447 (N_3447,N_2661,N_2713);
nor U3448 (N_3448,N_2470,N_2224);
or U3449 (N_3449,N_2647,N_2634);
nand U3450 (N_3450,N_2527,N_2419);
nand U3451 (N_3451,N_2192,N_2038);
or U3452 (N_3452,N_2364,N_2828);
or U3453 (N_3453,N_2851,N_2387);
nor U3454 (N_3454,N_2323,N_2546);
nor U3455 (N_3455,N_2092,N_2257);
or U3456 (N_3456,N_2152,N_2856);
or U3457 (N_3457,N_2370,N_2253);
or U3458 (N_3458,N_2269,N_2506);
nand U3459 (N_3459,N_2649,N_2819);
nor U3460 (N_3460,N_2010,N_2042);
nor U3461 (N_3461,N_2672,N_2981);
nand U3462 (N_3462,N_2596,N_2028);
or U3463 (N_3463,N_2837,N_2123);
or U3464 (N_3464,N_2491,N_2429);
and U3465 (N_3465,N_2699,N_2534);
nor U3466 (N_3466,N_2424,N_2402);
and U3467 (N_3467,N_2324,N_2404);
nand U3468 (N_3468,N_2185,N_2305);
and U3469 (N_3469,N_2626,N_2379);
nand U3470 (N_3470,N_2119,N_2754);
nand U3471 (N_3471,N_2893,N_2822);
or U3472 (N_3472,N_2744,N_2502);
nor U3473 (N_3473,N_2523,N_2648);
and U3474 (N_3474,N_2235,N_2768);
nand U3475 (N_3475,N_2436,N_2129);
and U3476 (N_3476,N_2679,N_2210);
or U3477 (N_3477,N_2193,N_2336);
nand U3478 (N_3478,N_2188,N_2883);
nand U3479 (N_3479,N_2514,N_2217);
nor U3480 (N_3480,N_2088,N_2761);
and U3481 (N_3481,N_2156,N_2784);
nand U3482 (N_3482,N_2979,N_2951);
nor U3483 (N_3483,N_2734,N_2033);
or U3484 (N_3484,N_2363,N_2800);
and U3485 (N_3485,N_2098,N_2459);
nor U3486 (N_3486,N_2121,N_2108);
or U3487 (N_3487,N_2299,N_2769);
xor U3488 (N_3488,N_2804,N_2348);
or U3489 (N_3489,N_2268,N_2478);
nor U3490 (N_3490,N_2006,N_2286);
nor U3491 (N_3491,N_2529,N_2841);
nor U3492 (N_3492,N_2637,N_2494);
nand U3493 (N_3493,N_2997,N_2326);
and U3494 (N_3494,N_2645,N_2967);
nand U3495 (N_3495,N_2731,N_2986);
xor U3496 (N_3496,N_2881,N_2122);
or U3497 (N_3497,N_2916,N_2887);
nor U3498 (N_3498,N_2155,N_2574);
or U3499 (N_3499,N_2275,N_2792);
nand U3500 (N_3500,N_2370,N_2369);
or U3501 (N_3501,N_2485,N_2355);
nand U3502 (N_3502,N_2855,N_2904);
or U3503 (N_3503,N_2006,N_2694);
nand U3504 (N_3504,N_2305,N_2959);
and U3505 (N_3505,N_2781,N_2722);
nand U3506 (N_3506,N_2899,N_2274);
nor U3507 (N_3507,N_2658,N_2064);
and U3508 (N_3508,N_2973,N_2294);
nor U3509 (N_3509,N_2371,N_2549);
and U3510 (N_3510,N_2979,N_2045);
nand U3511 (N_3511,N_2898,N_2376);
nor U3512 (N_3512,N_2188,N_2725);
nor U3513 (N_3513,N_2607,N_2395);
and U3514 (N_3514,N_2166,N_2477);
and U3515 (N_3515,N_2297,N_2509);
nand U3516 (N_3516,N_2009,N_2726);
xor U3517 (N_3517,N_2388,N_2309);
or U3518 (N_3518,N_2808,N_2867);
xnor U3519 (N_3519,N_2409,N_2384);
nand U3520 (N_3520,N_2273,N_2524);
nand U3521 (N_3521,N_2024,N_2737);
nand U3522 (N_3522,N_2533,N_2993);
and U3523 (N_3523,N_2894,N_2036);
or U3524 (N_3524,N_2422,N_2991);
xnor U3525 (N_3525,N_2789,N_2272);
nand U3526 (N_3526,N_2277,N_2580);
and U3527 (N_3527,N_2108,N_2341);
nand U3528 (N_3528,N_2429,N_2620);
or U3529 (N_3529,N_2458,N_2609);
nand U3530 (N_3530,N_2793,N_2483);
nand U3531 (N_3531,N_2508,N_2650);
nor U3532 (N_3532,N_2718,N_2133);
xor U3533 (N_3533,N_2945,N_2353);
xor U3534 (N_3534,N_2252,N_2063);
nor U3535 (N_3535,N_2005,N_2376);
or U3536 (N_3536,N_2133,N_2370);
xnor U3537 (N_3537,N_2255,N_2293);
xnor U3538 (N_3538,N_2469,N_2466);
or U3539 (N_3539,N_2162,N_2417);
nand U3540 (N_3540,N_2484,N_2904);
or U3541 (N_3541,N_2011,N_2231);
and U3542 (N_3542,N_2603,N_2633);
nor U3543 (N_3543,N_2355,N_2780);
xor U3544 (N_3544,N_2464,N_2617);
nor U3545 (N_3545,N_2187,N_2952);
nor U3546 (N_3546,N_2780,N_2639);
nor U3547 (N_3547,N_2995,N_2934);
and U3548 (N_3548,N_2219,N_2356);
or U3549 (N_3549,N_2469,N_2515);
nand U3550 (N_3550,N_2292,N_2461);
xnor U3551 (N_3551,N_2882,N_2045);
nor U3552 (N_3552,N_2690,N_2435);
and U3553 (N_3553,N_2465,N_2014);
xor U3554 (N_3554,N_2519,N_2151);
and U3555 (N_3555,N_2721,N_2575);
and U3556 (N_3556,N_2896,N_2856);
nor U3557 (N_3557,N_2535,N_2926);
or U3558 (N_3558,N_2517,N_2800);
nor U3559 (N_3559,N_2304,N_2255);
nand U3560 (N_3560,N_2589,N_2707);
xnor U3561 (N_3561,N_2750,N_2727);
or U3562 (N_3562,N_2350,N_2516);
and U3563 (N_3563,N_2497,N_2971);
and U3564 (N_3564,N_2274,N_2506);
nor U3565 (N_3565,N_2405,N_2004);
nor U3566 (N_3566,N_2199,N_2246);
or U3567 (N_3567,N_2752,N_2727);
nand U3568 (N_3568,N_2940,N_2974);
nor U3569 (N_3569,N_2128,N_2097);
nor U3570 (N_3570,N_2675,N_2045);
nor U3571 (N_3571,N_2767,N_2666);
or U3572 (N_3572,N_2426,N_2065);
nor U3573 (N_3573,N_2411,N_2210);
xor U3574 (N_3574,N_2802,N_2060);
and U3575 (N_3575,N_2828,N_2847);
xor U3576 (N_3576,N_2243,N_2170);
nor U3577 (N_3577,N_2674,N_2999);
or U3578 (N_3578,N_2258,N_2781);
or U3579 (N_3579,N_2815,N_2858);
and U3580 (N_3580,N_2306,N_2353);
nor U3581 (N_3581,N_2912,N_2473);
or U3582 (N_3582,N_2920,N_2391);
or U3583 (N_3583,N_2278,N_2213);
xnor U3584 (N_3584,N_2827,N_2965);
and U3585 (N_3585,N_2112,N_2256);
nor U3586 (N_3586,N_2466,N_2597);
nand U3587 (N_3587,N_2488,N_2352);
and U3588 (N_3588,N_2734,N_2930);
nand U3589 (N_3589,N_2750,N_2747);
or U3590 (N_3590,N_2924,N_2178);
nor U3591 (N_3591,N_2213,N_2131);
nor U3592 (N_3592,N_2370,N_2986);
or U3593 (N_3593,N_2777,N_2860);
and U3594 (N_3594,N_2661,N_2849);
nor U3595 (N_3595,N_2545,N_2760);
nand U3596 (N_3596,N_2991,N_2897);
or U3597 (N_3597,N_2823,N_2007);
and U3598 (N_3598,N_2322,N_2258);
and U3599 (N_3599,N_2751,N_2282);
and U3600 (N_3600,N_2012,N_2752);
nand U3601 (N_3601,N_2932,N_2172);
nand U3602 (N_3602,N_2019,N_2232);
xor U3603 (N_3603,N_2039,N_2372);
xor U3604 (N_3604,N_2162,N_2632);
nor U3605 (N_3605,N_2205,N_2070);
nor U3606 (N_3606,N_2454,N_2551);
or U3607 (N_3607,N_2711,N_2411);
and U3608 (N_3608,N_2048,N_2968);
nand U3609 (N_3609,N_2773,N_2177);
and U3610 (N_3610,N_2716,N_2903);
or U3611 (N_3611,N_2505,N_2902);
or U3612 (N_3612,N_2918,N_2542);
nor U3613 (N_3613,N_2596,N_2429);
or U3614 (N_3614,N_2810,N_2194);
and U3615 (N_3615,N_2856,N_2396);
nor U3616 (N_3616,N_2530,N_2286);
or U3617 (N_3617,N_2774,N_2581);
or U3618 (N_3618,N_2853,N_2278);
xor U3619 (N_3619,N_2251,N_2644);
xnor U3620 (N_3620,N_2633,N_2545);
nand U3621 (N_3621,N_2716,N_2994);
nor U3622 (N_3622,N_2159,N_2391);
and U3623 (N_3623,N_2425,N_2237);
nand U3624 (N_3624,N_2104,N_2248);
or U3625 (N_3625,N_2792,N_2661);
and U3626 (N_3626,N_2567,N_2416);
nand U3627 (N_3627,N_2370,N_2010);
and U3628 (N_3628,N_2946,N_2188);
or U3629 (N_3629,N_2467,N_2489);
nand U3630 (N_3630,N_2568,N_2043);
nand U3631 (N_3631,N_2502,N_2147);
xnor U3632 (N_3632,N_2817,N_2207);
or U3633 (N_3633,N_2258,N_2912);
nor U3634 (N_3634,N_2854,N_2498);
xor U3635 (N_3635,N_2410,N_2791);
and U3636 (N_3636,N_2339,N_2856);
nand U3637 (N_3637,N_2118,N_2874);
nor U3638 (N_3638,N_2308,N_2701);
nor U3639 (N_3639,N_2657,N_2642);
xor U3640 (N_3640,N_2907,N_2575);
nor U3641 (N_3641,N_2991,N_2009);
xnor U3642 (N_3642,N_2145,N_2732);
and U3643 (N_3643,N_2426,N_2852);
and U3644 (N_3644,N_2084,N_2105);
xnor U3645 (N_3645,N_2289,N_2882);
or U3646 (N_3646,N_2105,N_2211);
and U3647 (N_3647,N_2711,N_2104);
or U3648 (N_3648,N_2474,N_2403);
or U3649 (N_3649,N_2414,N_2569);
xnor U3650 (N_3650,N_2295,N_2246);
or U3651 (N_3651,N_2687,N_2755);
xnor U3652 (N_3652,N_2062,N_2090);
xor U3653 (N_3653,N_2294,N_2577);
nand U3654 (N_3654,N_2681,N_2188);
or U3655 (N_3655,N_2640,N_2750);
nor U3656 (N_3656,N_2087,N_2860);
nor U3657 (N_3657,N_2453,N_2184);
nor U3658 (N_3658,N_2454,N_2853);
nand U3659 (N_3659,N_2178,N_2672);
or U3660 (N_3660,N_2558,N_2760);
nand U3661 (N_3661,N_2177,N_2081);
nand U3662 (N_3662,N_2384,N_2909);
and U3663 (N_3663,N_2275,N_2925);
or U3664 (N_3664,N_2483,N_2741);
nor U3665 (N_3665,N_2043,N_2593);
nand U3666 (N_3666,N_2781,N_2290);
and U3667 (N_3667,N_2239,N_2427);
or U3668 (N_3668,N_2345,N_2594);
or U3669 (N_3669,N_2647,N_2133);
nand U3670 (N_3670,N_2506,N_2933);
and U3671 (N_3671,N_2174,N_2310);
and U3672 (N_3672,N_2411,N_2816);
or U3673 (N_3673,N_2286,N_2446);
or U3674 (N_3674,N_2391,N_2453);
nand U3675 (N_3675,N_2265,N_2049);
or U3676 (N_3676,N_2636,N_2461);
xor U3677 (N_3677,N_2641,N_2511);
nor U3678 (N_3678,N_2782,N_2521);
or U3679 (N_3679,N_2447,N_2581);
nand U3680 (N_3680,N_2085,N_2259);
nor U3681 (N_3681,N_2639,N_2826);
and U3682 (N_3682,N_2986,N_2773);
or U3683 (N_3683,N_2127,N_2193);
nor U3684 (N_3684,N_2002,N_2136);
nor U3685 (N_3685,N_2989,N_2458);
or U3686 (N_3686,N_2623,N_2059);
and U3687 (N_3687,N_2594,N_2078);
or U3688 (N_3688,N_2283,N_2092);
nor U3689 (N_3689,N_2762,N_2134);
nor U3690 (N_3690,N_2752,N_2172);
nor U3691 (N_3691,N_2348,N_2085);
or U3692 (N_3692,N_2764,N_2437);
nand U3693 (N_3693,N_2945,N_2611);
nand U3694 (N_3694,N_2000,N_2656);
nor U3695 (N_3695,N_2681,N_2324);
nand U3696 (N_3696,N_2720,N_2979);
or U3697 (N_3697,N_2002,N_2214);
and U3698 (N_3698,N_2212,N_2845);
or U3699 (N_3699,N_2065,N_2597);
nand U3700 (N_3700,N_2106,N_2128);
nand U3701 (N_3701,N_2267,N_2261);
and U3702 (N_3702,N_2051,N_2868);
xnor U3703 (N_3703,N_2966,N_2179);
nand U3704 (N_3704,N_2438,N_2917);
nand U3705 (N_3705,N_2707,N_2474);
nor U3706 (N_3706,N_2807,N_2623);
or U3707 (N_3707,N_2260,N_2882);
nand U3708 (N_3708,N_2762,N_2392);
and U3709 (N_3709,N_2243,N_2697);
nand U3710 (N_3710,N_2912,N_2117);
xnor U3711 (N_3711,N_2687,N_2739);
nor U3712 (N_3712,N_2047,N_2528);
or U3713 (N_3713,N_2588,N_2725);
nor U3714 (N_3714,N_2381,N_2876);
nor U3715 (N_3715,N_2564,N_2544);
nor U3716 (N_3716,N_2812,N_2293);
xnor U3717 (N_3717,N_2733,N_2105);
nor U3718 (N_3718,N_2377,N_2581);
or U3719 (N_3719,N_2703,N_2114);
nand U3720 (N_3720,N_2482,N_2950);
nor U3721 (N_3721,N_2969,N_2960);
nand U3722 (N_3722,N_2390,N_2911);
nor U3723 (N_3723,N_2789,N_2240);
nor U3724 (N_3724,N_2545,N_2060);
or U3725 (N_3725,N_2585,N_2958);
and U3726 (N_3726,N_2846,N_2092);
or U3727 (N_3727,N_2463,N_2910);
and U3728 (N_3728,N_2410,N_2489);
or U3729 (N_3729,N_2278,N_2962);
nand U3730 (N_3730,N_2283,N_2258);
nor U3731 (N_3731,N_2475,N_2364);
nor U3732 (N_3732,N_2722,N_2612);
nand U3733 (N_3733,N_2395,N_2705);
xor U3734 (N_3734,N_2534,N_2423);
and U3735 (N_3735,N_2583,N_2484);
and U3736 (N_3736,N_2676,N_2916);
and U3737 (N_3737,N_2035,N_2695);
nor U3738 (N_3738,N_2422,N_2174);
and U3739 (N_3739,N_2258,N_2687);
nand U3740 (N_3740,N_2729,N_2236);
nor U3741 (N_3741,N_2712,N_2171);
nand U3742 (N_3742,N_2791,N_2436);
nand U3743 (N_3743,N_2495,N_2038);
nand U3744 (N_3744,N_2253,N_2584);
nor U3745 (N_3745,N_2345,N_2649);
nand U3746 (N_3746,N_2429,N_2858);
and U3747 (N_3747,N_2529,N_2392);
nor U3748 (N_3748,N_2846,N_2812);
nor U3749 (N_3749,N_2482,N_2661);
xnor U3750 (N_3750,N_2028,N_2944);
nor U3751 (N_3751,N_2779,N_2899);
nand U3752 (N_3752,N_2467,N_2304);
or U3753 (N_3753,N_2380,N_2226);
nor U3754 (N_3754,N_2276,N_2039);
or U3755 (N_3755,N_2051,N_2302);
nor U3756 (N_3756,N_2449,N_2907);
nand U3757 (N_3757,N_2883,N_2871);
or U3758 (N_3758,N_2427,N_2164);
and U3759 (N_3759,N_2462,N_2907);
or U3760 (N_3760,N_2724,N_2072);
and U3761 (N_3761,N_2223,N_2004);
nor U3762 (N_3762,N_2419,N_2560);
and U3763 (N_3763,N_2734,N_2421);
nand U3764 (N_3764,N_2349,N_2863);
and U3765 (N_3765,N_2684,N_2119);
nand U3766 (N_3766,N_2284,N_2814);
nand U3767 (N_3767,N_2690,N_2152);
and U3768 (N_3768,N_2440,N_2310);
or U3769 (N_3769,N_2546,N_2397);
nand U3770 (N_3770,N_2782,N_2911);
and U3771 (N_3771,N_2805,N_2051);
nor U3772 (N_3772,N_2923,N_2282);
nor U3773 (N_3773,N_2541,N_2870);
or U3774 (N_3774,N_2623,N_2507);
and U3775 (N_3775,N_2540,N_2990);
xor U3776 (N_3776,N_2098,N_2400);
nand U3777 (N_3777,N_2280,N_2060);
and U3778 (N_3778,N_2033,N_2812);
and U3779 (N_3779,N_2674,N_2368);
nand U3780 (N_3780,N_2928,N_2750);
and U3781 (N_3781,N_2385,N_2530);
nand U3782 (N_3782,N_2581,N_2701);
nor U3783 (N_3783,N_2103,N_2222);
and U3784 (N_3784,N_2488,N_2121);
and U3785 (N_3785,N_2796,N_2897);
nor U3786 (N_3786,N_2749,N_2114);
nor U3787 (N_3787,N_2198,N_2515);
nor U3788 (N_3788,N_2928,N_2689);
and U3789 (N_3789,N_2809,N_2486);
and U3790 (N_3790,N_2531,N_2821);
and U3791 (N_3791,N_2028,N_2817);
and U3792 (N_3792,N_2319,N_2761);
or U3793 (N_3793,N_2165,N_2776);
nand U3794 (N_3794,N_2777,N_2616);
xnor U3795 (N_3795,N_2695,N_2559);
xor U3796 (N_3796,N_2700,N_2523);
and U3797 (N_3797,N_2744,N_2018);
and U3798 (N_3798,N_2733,N_2244);
nand U3799 (N_3799,N_2753,N_2568);
and U3800 (N_3800,N_2521,N_2915);
or U3801 (N_3801,N_2157,N_2016);
and U3802 (N_3802,N_2899,N_2095);
or U3803 (N_3803,N_2342,N_2362);
nor U3804 (N_3804,N_2561,N_2352);
and U3805 (N_3805,N_2047,N_2966);
and U3806 (N_3806,N_2668,N_2594);
and U3807 (N_3807,N_2123,N_2357);
or U3808 (N_3808,N_2161,N_2119);
and U3809 (N_3809,N_2366,N_2031);
or U3810 (N_3810,N_2116,N_2928);
nand U3811 (N_3811,N_2670,N_2292);
and U3812 (N_3812,N_2293,N_2653);
nor U3813 (N_3813,N_2750,N_2133);
and U3814 (N_3814,N_2319,N_2201);
or U3815 (N_3815,N_2239,N_2277);
nand U3816 (N_3816,N_2817,N_2219);
or U3817 (N_3817,N_2879,N_2637);
nand U3818 (N_3818,N_2262,N_2291);
nand U3819 (N_3819,N_2395,N_2919);
and U3820 (N_3820,N_2841,N_2226);
and U3821 (N_3821,N_2643,N_2311);
or U3822 (N_3822,N_2593,N_2222);
nor U3823 (N_3823,N_2004,N_2356);
or U3824 (N_3824,N_2259,N_2800);
xor U3825 (N_3825,N_2397,N_2179);
nor U3826 (N_3826,N_2309,N_2506);
xor U3827 (N_3827,N_2940,N_2852);
or U3828 (N_3828,N_2402,N_2008);
nand U3829 (N_3829,N_2834,N_2392);
and U3830 (N_3830,N_2956,N_2534);
nor U3831 (N_3831,N_2907,N_2465);
nor U3832 (N_3832,N_2844,N_2842);
or U3833 (N_3833,N_2040,N_2530);
or U3834 (N_3834,N_2984,N_2600);
and U3835 (N_3835,N_2360,N_2354);
nor U3836 (N_3836,N_2805,N_2511);
nor U3837 (N_3837,N_2039,N_2247);
nand U3838 (N_3838,N_2836,N_2041);
nand U3839 (N_3839,N_2440,N_2940);
nand U3840 (N_3840,N_2187,N_2182);
or U3841 (N_3841,N_2403,N_2232);
and U3842 (N_3842,N_2321,N_2236);
or U3843 (N_3843,N_2535,N_2190);
nand U3844 (N_3844,N_2096,N_2284);
nand U3845 (N_3845,N_2672,N_2179);
nor U3846 (N_3846,N_2337,N_2037);
nand U3847 (N_3847,N_2823,N_2002);
or U3848 (N_3848,N_2346,N_2658);
nand U3849 (N_3849,N_2102,N_2879);
nor U3850 (N_3850,N_2149,N_2931);
and U3851 (N_3851,N_2223,N_2390);
nor U3852 (N_3852,N_2300,N_2062);
and U3853 (N_3853,N_2420,N_2405);
nor U3854 (N_3854,N_2659,N_2566);
nand U3855 (N_3855,N_2213,N_2711);
or U3856 (N_3856,N_2502,N_2811);
or U3857 (N_3857,N_2161,N_2085);
and U3858 (N_3858,N_2981,N_2369);
nor U3859 (N_3859,N_2162,N_2344);
nor U3860 (N_3860,N_2531,N_2726);
nand U3861 (N_3861,N_2963,N_2381);
or U3862 (N_3862,N_2786,N_2701);
or U3863 (N_3863,N_2640,N_2707);
and U3864 (N_3864,N_2430,N_2088);
nand U3865 (N_3865,N_2902,N_2850);
nand U3866 (N_3866,N_2984,N_2233);
and U3867 (N_3867,N_2777,N_2003);
and U3868 (N_3868,N_2179,N_2139);
nand U3869 (N_3869,N_2261,N_2034);
or U3870 (N_3870,N_2889,N_2114);
and U3871 (N_3871,N_2257,N_2517);
and U3872 (N_3872,N_2066,N_2842);
and U3873 (N_3873,N_2040,N_2633);
nor U3874 (N_3874,N_2262,N_2251);
nand U3875 (N_3875,N_2638,N_2372);
or U3876 (N_3876,N_2126,N_2065);
nor U3877 (N_3877,N_2896,N_2580);
or U3878 (N_3878,N_2355,N_2374);
or U3879 (N_3879,N_2972,N_2684);
nor U3880 (N_3880,N_2988,N_2202);
or U3881 (N_3881,N_2167,N_2795);
or U3882 (N_3882,N_2588,N_2005);
or U3883 (N_3883,N_2008,N_2653);
or U3884 (N_3884,N_2505,N_2891);
nand U3885 (N_3885,N_2035,N_2602);
nor U3886 (N_3886,N_2773,N_2524);
and U3887 (N_3887,N_2682,N_2680);
and U3888 (N_3888,N_2690,N_2700);
and U3889 (N_3889,N_2808,N_2352);
nand U3890 (N_3890,N_2649,N_2365);
nor U3891 (N_3891,N_2508,N_2872);
or U3892 (N_3892,N_2275,N_2949);
nor U3893 (N_3893,N_2881,N_2977);
nor U3894 (N_3894,N_2103,N_2261);
nand U3895 (N_3895,N_2718,N_2865);
nor U3896 (N_3896,N_2102,N_2639);
and U3897 (N_3897,N_2842,N_2783);
and U3898 (N_3898,N_2472,N_2722);
and U3899 (N_3899,N_2282,N_2223);
nor U3900 (N_3900,N_2841,N_2757);
or U3901 (N_3901,N_2365,N_2595);
and U3902 (N_3902,N_2426,N_2419);
xnor U3903 (N_3903,N_2363,N_2964);
or U3904 (N_3904,N_2509,N_2678);
and U3905 (N_3905,N_2413,N_2712);
nand U3906 (N_3906,N_2057,N_2355);
nand U3907 (N_3907,N_2489,N_2336);
or U3908 (N_3908,N_2834,N_2458);
and U3909 (N_3909,N_2038,N_2928);
or U3910 (N_3910,N_2348,N_2035);
and U3911 (N_3911,N_2803,N_2713);
and U3912 (N_3912,N_2214,N_2006);
nand U3913 (N_3913,N_2466,N_2912);
nand U3914 (N_3914,N_2971,N_2085);
xor U3915 (N_3915,N_2204,N_2041);
nand U3916 (N_3916,N_2133,N_2448);
nor U3917 (N_3917,N_2848,N_2802);
nand U3918 (N_3918,N_2214,N_2290);
nor U3919 (N_3919,N_2500,N_2201);
or U3920 (N_3920,N_2861,N_2673);
or U3921 (N_3921,N_2794,N_2850);
xor U3922 (N_3922,N_2840,N_2447);
nor U3923 (N_3923,N_2013,N_2286);
xor U3924 (N_3924,N_2113,N_2347);
nand U3925 (N_3925,N_2099,N_2285);
nor U3926 (N_3926,N_2071,N_2845);
or U3927 (N_3927,N_2660,N_2479);
or U3928 (N_3928,N_2885,N_2374);
nand U3929 (N_3929,N_2255,N_2992);
nand U3930 (N_3930,N_2786,N_2599);
nor U3931 (N_3931,N_2309,N_2959);
nor U3932 (N_3932,N_2836,N_2385);
or U3933 (N_3933,N_2941,N_2531);
nor U3934 (N_3934,N_2854,N_2556);
nand U3935 (N_3935,N_2472,N_2290);
xnor U3936 (N_3936,N_2749,N_2427);
and U3937 (N_3937,N_2408,N_2192);
nor U3938 (N_3938,N_2021,N_2125);
nor U3939 (N_3939,N_2948,N_2807);
xnor U3940 (N_3940,N_2910,N_2858);
nor U3941 (N_3941,N_2500,N_2975);
or U3942 (N_3942,N_2818,N_2194);
nor U3943 (N_3943,N_2807,N_2915);
nand U3944 (N_3944,N_2029,N_2341);
and U3945 (N_3945,N_2839,N_2637);
and U3946 (N_3946,N_2224,N_2323);
or U3947 (N_3947,N_2450,N_2363);
or U3948 (N_3948,N_2450,N_2721);
or U3949 (N_3949,N_2231,N_2646);
and U3950 (N_3950,N_2971,N_2273);
nand U3951 (N_3951,N_2420,N_2593);
and U3952 (N_3952,N_2277,N_2739);
xor U3953 (N_3953,N_2508,N_2193);
nand U3954 (N_3954,N_2080,N_2847);
and U3955 (N_3955,N_2790,N_2636);
and U3956 (N_3956,N_2406,N_2429);
nand U3957 (N_3957,N_2252,N_2090);
nand U3958 (N_3958,N_2764,N_2413);
xor U3959 (N_3959,N_2786,N_2519);
or U3960 (N_3960,N_2459,N_2090);
nor U3961 (N_3961,N_2081,N_2688);
and U3962 (N_3962,N_2666,N_2021);
and U3963 (N_3963,N_2920,N_2661);
nor U3964 (N_3964,N_2699,N_2669);
xnor U3965 (N_3965,N_2597,N_2859);
or U3966 (N_3966,N_2160,N_2719);
nor U3967 (N_3967,N_2001,N_2909);
or U3968 (N_3968,N_2535,N_2240);
or U3969 (N_3969,N_2274,N_2510);
nand U3970 (N_3970,N_2502,N_2289);
nand U3971 (N_3971,N_2186,N_2136);
or U3972 (N_3972,N_2777,N_2188);
nand U3973 (N_3973,N_2154,N_2870);
or U3974 (N_3974,N_2549,N_2583);
nor U3975 (N_3975,N_2492,N_2618);
nand U3976 (N_3976,N_2605,N_2990);
nor U3977 (N_3977,N_2662,N_2560);
and U3978 (N_3978,N_2725,N_2491);
or U3979 (N_3979,N_2218,N_2920);
or U3980 (N_3980,N_2388,N_2379);
nand U3981 (N_3981,N_2578,N_2860);
or U3982 (N_3982,N_2092,N_2130);
and U3983 (N_3983,N_2948,N_2277);
and U3984 (N_3984,N_2055,N_2529);
nor U3985 (N_3985,N_2528,N_2469);
or U3986 (N_3986,N_2941,N_2930);
nor U3987 (N_3987,N_2517,N_2526);
nor U3988 (N_3988,N_2592,N_2856);
and U3989 (N_3989,N_2691,N_2349);
or U3990 (N_3990,N_2111,N_2855);
nand U3991 (N_3991,N_2007,N_2244);
or U3992 (N_3992,N_2930,N_2412);
or U3993 (N_3993,N_2452,N_2755);
nand U3994 (N_3994,N_2736,N_2945);
nor U3995 (N_3995,N_2678,N_2534);
xor U3996 (N_3996,N_2091,N_2534);
xor U3997 (N_3997,N_2999,N_2821);
and U3998 (N_3998,N_2570,N_2110);
nand U3999 (N_3999,N_2853,N_2988);
nor U4000 (N_4000,N_3920,N_3867);
xor U4001 (N_4001,N_3218,N_3880);
or U4002 (N_4002,N_3862,N_3709);
nand U4003 (N_4003,N_3843,N_3447);
xnor U4004 (N_4004,N_3342,N_3759);
and U4005 (N_4005,N_3388,N_3486);
nor U4006 (N_4006,N_3762,N_3414);
and U4007 (N_4007,N_3804,N_3153);
xnor U4008 (N_4008,N_3972,N_3010);
or U4009 (N_4009,N_3555,N_3874);
nor U4010 (N_4010,N_3864,N_3608);
or U4011 (N_4011,N_3537,N_3931);
xnor U4012 (N_4012,N_3358,N_3444);
or U4013 (N_4013,N_3875,N_3522);
or U4014 (N_4014,N_3248,N_3210);
and U4015 (N_4015,N_3623,N_3487);
xor U4016 (N_4016,N_3283,N_3127);
nand U4017 (N_4017,N_3377,N_3661);
and U4018 (N_4018,N_3173,N_3566);
or U4019 (N_4019,N_3273,N_3230);
or U4020 (N_4020,N_3686,N_3446);
nor U4021 (N_4021,N_3160,N_3036);
or U4022 (N_4022,N_3368,N_3390);
or U4023 (N_4023,N_3224,N_3202);
or U4024 (N_4024,N_3723,N_3016);
and U4025 (N_4025,N_3611,N_3459);
and U4026 (N_4026,N_3167,N_3635);
nand U4027 (N_4027,N_3883,N_3485);
and U4028 (N_4028,N_3062,N_3268);
or U4029 (N_4029,N_3278,N_3775);
nor U4030 (N_4030,N_3474,N_3691);
nand U4031 (N_4031,N_3831,N_3114);
and U4032 (N_4032,N_3734,N_3135);
or U4033 (N_4033,N_3174,N_3809);
xor U4034 (N_4034,N_3535,N_3333);
or U4035 (N_4035,N_3648,N_3760);
or U4036 (N_4036,N_3392,N_3212);
or U4037 (N_4037,N_3871,N_3011);
xnor U4038 (N_4038,N_3288,N_3764);
nor U4039 (N_4039,N_3823,N_3860);
nor U4040 (N_4040,N_3621,N_3731);
xnor U4041 (N_4041,N_3163,N_3196);
nand U4042 (N_4042,N_3583,N_3585);
xor U4043 (N_4043,N_3440,N_3742);
nand U4044 (N_4044,N_3622,N_3391);
or U4045 (N_4045,N_3798,N_3477);
nor U4046 (N_4046,N_3292,N_3675);
nor U4047 (N_4047,N_3293,N_3887);
nor U4048 (N_4048,N_3554,N_3647);
nor U4049 (N_4049,N_3665,N_3143);
or U4050 (N_4050,N_3311,N_3393);
nor U4051 (N_4051,N_3467,N_3480);
nand U4052 (N_4052,N_3145,N_3028);
or U4053 (N_4053,N_3296,N_3873);
or U4054 (N_4054,N_3136,N_3992);
and U4055 (N_4055,N_3654,N_3866);
nand U4056 (N_4056,N_3024,N_3352);
or U4057 (N_4057,N_3948,N_3420);
and U4058 (N_4058,N_3921,N_3934);
nor U4059 (N_4059,N_3568,N_3175);
nor U4060 (N_4060,N_3814,N_3200);
and U4061 (N_4061,N_3400,N_3189);
or U4062 (N_4062,N_3641,N_3501);
nand U4063 (N_4063,N_3952,N_3735);
nor U4064 (N_4064,N_3490,N_3262);
nor U4065 (N_4065,N_3989,N_3194);
nor U4066 (N_4066,N_3861,N_3591);
nor U4067 (N_4067,N_3243,N_3969);
and U4068 (N_4068,N_3544,N_3386);
or U4069 (N_4069,N_3106,N_3778);
nor U4070 (N_4070,N_3201,N_3916);
nor U4071 (N_4071,N_3048,N_3567);
and U4072 (N_4072,N_3780,N_3550);
xor U4073 (N_4073,N_3813,N_3919);
or U4074 (N_4074,N_3402,N_3154);
or U4075 (N_4075,N_3499,N_3721);
nor U4076 (N_4076,N_3796,N_3897);
xor U4077 (N_4077,N_3833,N_3557);
nand U4078 (N_4078,N_3614,N_3679);
nand U4079 (N_4079,N_3081,N_3882);
xor U4080 (N_4080,N_3363,N_3624);
or U4081 (N_4081,N_3133,N_3620);
or U4082 (N_4082,N_3807,N_3411);
nand U4083 (N_4083,N_3784,N_3337);
nand U4084 (N_4084,N_3852,N_3085);
and U4085 (N_4085,N_3455,N_3445);
nor U4086 (N_4086,N_3284,N_3443);
or U4087 (N_4087,N_3839,N_3435);
nand U4088 (N_4088,N_3877,N_3034);
or U4089 (N_4089,N_3859,N_3000);
or U4090 (N_4090,N_3613,N_3604);
nand U4091 (N_4091,N_3941,N_3587);
or U4092 (N_4092,N_3628,N_3131);
or U4093 (N_4093,N_3602,N_3714);
and U4094 (N_4094,N_3379,N_3090);
or U4095 (N_4095,N_3161,N_3682);
nand U4096 (N_4096,N_3002,N_3067);
nand U4097 (N_4097,N_3932,N_3380);
or U4098 (N_4098,N_3494,N_3412);
or U4099 (N_4099,N_3222,N_3704);
nor U4100 (N_4100,N_3336,N_3851);
and U4101 (N_4101,N_3774,N_3598);
nand U4102 (N_4102,N_3270,N_3732);
nor U4103 (N_4103,N_3961,N_3801);
nor U4104 (N_4104,N_3410,N_3779);
and U4105 (N_4105,N_3895,N_3018);
or U4106 (N_4106,N_3508,N_3898);
or U4107 (N_4107,N_3902,N_3981);
nand U4108 (N_4108,N_3592,N_3536);
nand U4109 (N_4109,N_3318,N_3773);
and U4110 (N_4110,N_3226,N_3022);
or U4111 (N_4111,N_3538,N_3936);
and U4112 (N_4112,N_3188,N_3103);
nor U4113 (N_4113,N_3097,N_3206);
xor U4114 (N_4114,N_3346,N_3396);
nand U4115 (N_4115,N_3893,N_3975);
nor U4116 (N_4116,N_3247,N_3818);
nand U4117 (N_4117,N_3542,N_3965);
nand U4118 (N_4118,N_3905,N_3700);
nand U4119 (N_4119,N_3706,N_3511);
and U4120 (N_4120,N_3289,N_3539);
nor U4121 (N_4121,N_3607,N_3806);
and U4122 (N_4122,N_3245,N_3171);
or U4123 (N_4123,N_3427,N_3408);
nand U4124 (N_4124,N_3345,N_3821);
and U4125 (N_4125,N_3279,N_3110);
or U4126 (N_4126,N_3159,N_3914);
and U4127 (N_4127,N_3701,N_3122);
nand U4128 (N_4128,N_3302,N_3421);
nand U4129 (N_4129,N_3979,N_3316);
nor U4130 (N_4130,N_3484,N_3261);
xnor U4131 (N_4131,N_3238,N_3193);
nand U4132 (N_4132,N_3586,N_3083);
and U4133 (N_4133,N_3930,N_3693);
nor U4134 (N_4134,N_3102,N_3357);
and U4135 (N_4135,N_3810,N_3208);
nand U4136 (N_4136,N_3182,N_3929);
nand U4137 (N_4137,N_3609,N_3560);
nand U4138 (N_4138,N_3974,N_3475);
and U4139 (N_4139,N_3255,N_3741);
or U4140 (N_4140,N_3448,N_3190);
nand U4141 (N_4141,N_3514,N_3678);
nand U4142 (N_4142,N_3186,N_3012);
nand U4143 (N_4143,N_3978,N_3533);
and U4144 (N_4144,N_3319,N_3359);
nor U4145 (N_4145,N_3770,N_3053);
and U4146 (N_4146,N_3640,N_3235);
nor U4147 (N_4147,N_3394,N_3505);
nand U4148 (N_4148,N_3783,N_3324);
nand U4149 (N_4149,N_3968,N_3372);
and U4150 (N_4150,N_3951,N_3170);
nand U4151 (N_4151,N_3439,N_3680);
nand U4152 (N_4152,N_3498,N_3457);
or U4153 (N_4153,N_3808,N_3828);
and U4154 (N_4154,N_3939,N_3483);
nand U4155 (N_4155,N_3325,N_3373);
and U4156 (N_4156,N_3959,N_3451);
or U4157 (N_4157,N_3672,N_3387);
nand U4158 (N_4158,N_3223,N_3531);
xor U4159 (N_4159,N_3777,N_3631);
nand U4160 (N_4160,N_3184,N_3082);
nor U4161 (N_4161,N_3558,N_3313);
and U4162 (N_4162,N_3076,N_3872);
nor U4163 (N_4163,N_3479,N_3954);
nor U4164 (N_4164,N_3967,N_3216);
and U4165 (N_4165,N_3697,N_3579);
and U4166 (N_4166,N_3304,N_3219);
nand U4167 (N_4167,N_3633,N_3320);
xnor U4168 (N_4168,N_3306,N_3128);
nand U4169 (N_4169,N_3149,N_3695);
nor U4170 (N_4170,N_3619,N_3785);
nor U4171 (N_4171,N_3684,N_3205);
nand U4172 (N_4172,N_3037,N_3546);
and U4173 (N_4173,N_3792,N_3815);
or U4174 (N_4174,N_3855,N_3429);
and U4175 (N_4175,N_3793,N_3722);
or U4176 (N_4176,N_3917,N_3718);
nand U4177 (N_4177,N_3049,N_3995);
nand U4178 (N_4178,N_3822,N_3087);
nand U4179 (N_4179,N_3099,N_3572);
xor U4180 (N_4180,N_3924,N_3158);
nor U4181 (N_4181,N_3891,N_3213);
or U4182 (N_4182,N_3234,N_3364);
nand U4183 (N_4183,N_3039,N_3079);
and U4184 (N_4184,N_3653,N_3799);
and U4185 (N_4185,N_3669,N_3582);
nand U4186 (N_4186,N_3056,N_3847);
or U4187 (N_4187,N_3908,N_3378);
or U4188 (N_4188,N_3603,N_3006);
or U4189 (N_4189,N_3254,N_3155);
nand U4190 (N_4190,N_3528,N_3842);
or U4191 (N_4191,N_3834,N_3267);
or U4192 (N_4192,N_3468,N_3856);
and U4193 (N_4193,N_3740,N_3549);
nand U4194 (N_4194,N_3524,N_3589);
nand U4195 (N_4195,N_3698,N_3343);
or U4196 (N_4196,N_3026,N_3331);
or U4197 (N_4197,N_3300,N_3502);
nor U4198 (N_4198,N_3559,N_3575);
or U4199 (N_4199,N_3187,N_3976);
or U4200 (N_4200,N_3009,N_3064);
nand U4201 (N_4201,N_3705,N_3627);
or U4202 (N_4202,N_3973,N_3600);
nor U4203 (N_4203,N_3172,N_3599);
and U4204 (N_4204,N_3199,N_3264);
nand U4205 (N_4205,N_3984,N_3144);
nand U4206 (N_4206,N_3465,N_3356);
nor U4207 (N_4207,N_3758,N_3258);
nor U4208 (N_4208,N_3738,N_3957);
and U4209 (N_4209,N_3383,N_3339);
nor U4210 (N_4210,N_3460,N_3947);
and U4211 (N_4211,N_3168,N_3795);
nor U4212 (N_4212,N_3417,N_3482);
nor U4213 (N_4213,N_3694,N_3894);
nor U4214 (N_4214,N_3727,N_3282);
xnor U4215 (N_4215,N_3040,N_3636);
or U4216 (N_4216,N_3632,N_3362);
nor U4217 (N_4217,N_3398,N_3577);
nand U4218 (N_4218,N_3327,N_3500);
and U4219 (N_4219,N_3433,N_3826);
and U4220 (N_4220,N_3370,N_3491);
xnor U4221 (N_4221,N_3518,N_3148);
nand U4222 (N_4222,N_3658,N_3432);
or U4223 (N_4223,N_3013,N_3584);
xnor U4224 (N_4224,N_3928,N_3719);
and U4225 (N_4225,N_3660,N_3985);
nor U4226 (N_4226,N_3115,N_3425);
xor U4227 (N_4227,N_3285,N_3495);
and U4228 (N_4228,N_3117,N_3492);
nand U4229 (N_4229,N_3938,N_3138);
nand U4230 (N_4230,N_3074,N_3747);
or U4231 (N_4231,N_3771,N_3310);
and U4232 (N_4232,N_3113,N_3280);
and U4233 (N_4233,N_3574,N_3980);
nor U4234 (N_4234,N_3848,N_3207);
or U4235 (N_4235,N_3032,N_3845);
nor U4236 (N_4236,N_3098,N_3183);
or U4237 (N_4237,N_3015,N_3580);
nor U4238 (N_4238,N_3260,N_3922);
nand U4239 (N_4239,N_3050,N_3753);
xnor U4240 (N_4240,N_3696,N_3228);
nor U4241 (N_4241,N_3305,N_3096);
nor U4242 (N_4242,N_3545,N_3365);
and U4243 (N_4243,N_3382,N_3712);
nand U4244 (N_4244,N_3715,N_3047);
and U4245 (N_4245,N_3752,N_3519);
and U4246 (N_4246,N_3178,N_3236);
or U4247 (N_4247,N_3366,N_3787);
or U4248 (N_4248,N_3926,N_3552);
nand U4249 (N_4249,N_3576,N_3233);
or U4250 (N_4250,N_3430,N_3878);
and U4251 (N_4251,N_3949,N_3720);
nand U4252 (N_4252,N_3021,N_3676);
nand U4253 (N_4253,N_3225,N_3058);
xnor U4254 (N_4254,N_3563,N_3125);
nor U4255 (N_4255,N_3166,N_3068);
nand U4256 (N_4256,N_3541,N_3340);
or U4257 (N_4257,N_3211,N_3060);
and U4258 (N_4258,N_3458,N_3130);
and U4259 (N_4259,N_3999,N_3835);
nor U4260 (N_4260,N_3923,N_3892);
nor U4261 (N_4261,N_3562,N_3863);
xor U4262 (N_4262,N_3204,N_3084);
xnor U4263 (N_4263,N_3092,N_3825);
nand U4264 (N_4264,N_3088,N_3523);
nor U4265 (N_4265,N_3497,N_3739);
and U4266 (N_4266,N_3755,N_3464);
nand U4267 (N_4267,N_3666,N_3297);
or U4268 (N_4268,N_3901,N_3385);
and U4269 (N_4269,N_3059,N_3504);
or U4270 (N_4270,N_3516,N_3470);
nor U4271 (N_4271,N_3038,N_3244);
nor U4272 (N_4272,N_3045,N_3513);
or U4273 (N_4273,N_3904,N_3071);
nor U4274 (N_4274,N_3360,N_3745);
or U4275 (N_4275,N_3315,N_3215);
nand U4276 (N_4276,N_3790,N_3532);
nand U4277 (N_4277,N_3118,N_3942);
xnor U4278 (N_4278,N_3104,N_3423);
nand U4279 (N_4279,N_3652,N_3935);
nor U4280 (N_4280,N_3570,N_3111);
nor U4281 (N_4281,N_3351,N_3257);
nor U4282 (N_4282,N_3334,N_3918);
and U4283 (N_4283,N_3716,N_3865);
and U4284 (N_4284,N_3132,N_3946);
nand U4285 (N_4285,N_3332,N_3330);
or U4286 (N_4286,N_3618,N_3997);
or U4287 (N_4287,N_3900,N_3030);
nand U4288 (N_4288,N_3890,N_3830);
nand U4289 (N_4289,N_3548,N_3181);
and U4290 (N_4290,N_3072,N_3454);
nor U4291 (N_4291,N_3593,N_3404);
nand U4292 (N_4292,N_3141,N_3736);
nand U4293 (N_4293,N_3927,N_3525);
xor U4294 (N_4294,N_3564,N_3191);
or U4295 (N_4295,N_3303,N_3765);
and U4296 (N_4296,N_3766,N_3512);
and U4297 (N_4297,N_3126,N_3077);
or U4298 (N_4298,N_3651,N_3868);
or U4299 (N_4299,N_3517,N_3431);
or U4300 (N_4300,N_3031,N_3750);
and U4301 (N_4301,N_3744,N_3990);
or U4302 (N_4302,N_3051,N_3556);
xor U4303 (N_4303,N_3349,N_3017);
and U4304 (N_4304,N_3462,N_3657);
or U4305 (N_4305,N_3322,N_3070);
and U4306 (N_4306,N_3998,N_3699);
xor U4307 (N_4307,N_3019,N_3291);
nor U4308 (N_4308,N_3381,N_3768);
nor U4309 (N_4309,N_3348,N_3471);
or U4310 (N_4310,N_3646,N_3913);
nor U4311 (N_4311,N_3023,N_3043);
nand U4312 (N_4312,N_3341,N_3945);
xnor U4313 (N_4313,N_3662,N_3725);
or U4314 (N_4314,N_3256,N_3272);
or U4315 (N_4315,N_3249,N_3637);
and U4316 (N_4316,N_3616,N_3452);
and U4317 (N_4317,N_3674,N_3659);
and U4318 (N_4318,N_3655,N_3061);
nor U4319 (N_4319,N_3726,N_3899);
nor U4320 (N_4320,N_3724,N_3020);
and U4321 (N_4321,N_3885,N_3673);
or U4322 (N_4322,N_3046,N_3746);
nor U4323 (N_4323,N_3326,N_3237);
or U4324 (N_4324,N_3395,N_3473);
nand U4325 (N_4325,N_3150,N_3095);
or U4326 (N_4326,N_3710,N_3418);
nor U4327 (N_4327,N_3137,N_3376);
or U4328 (N_4328,N_3271,N_3052);
and U4329 (N_4329,N_3123,N_3925);
xor U4330 (N_4330,N_3817,N_3287);
nor U4331 (N_4331,N_3625,N_3642);
and U4332 (N_4332,N_3849,N_3933);
nor U4333 (N_4333,N_3434,N_3107);
xnor U4334 (N_4334,N_3756,N_3966);
or U4335 (N_4335,N_3910,N_3496);
or U4336 (N_4336,N_3707,N_3685);
and U4337 (N_4337,N_3754,N_3422);
nor U4338 (N_4338,N_3645,N_3007);
nor U4339 (N_4339,N_3854,N_3140);
nand U4340 (N_4340,N_3605,N_3829);
or U4341 (N_4341,N_3789,N_3595);
xor U4342 (N_4342,N_3129,N_3403);
and U4343 (N_4343,N_3108,N_3708);
nand U4344 (N_4344,N_3438,N_3717);
nand U4345 (N_4345,N_3503,N_3819);
or U4346 (N_4346,N_3761,N_3769);
nor U4347 (N_4347,N_3361,N_3231);
nor U4348 (N_4348,N_3008,N_3065);
and U4349 (N_4349,N_3240,N_3767);
nand U4350 (N_4350,N_3937,N_3419);
nand U4351 (N_4351,N_3275,N_3266);
nand U4352 (N_4352,N_3307,N_3399);
nand U4353 (N_4353,N_3005,N_3820);
and U4354 (N_4354,N_3197,N_3711);
xnor U4355 (N_4355,N_3165,N_3469);
nor U4356 (N_4356,N_3347,N_3800);
and U4357 (N_4357,N_3335,N_3232);
nor U4358 (N_4358,N_3080,N_3146);
or U4359 (N_4359,N_3786,N_3994);
nand U4360 (N_4360,N_3903,N_3838);
or U4361 (N_4361,N_3488,N_3220);
or U4362 (N_4362,N_3543,N_3229);
xor U4363 (N_4363,N_3269,N_3987);
and U4364 (N_4364,N_3827,N_3578);
nand U4365 (N_4365,N_3367,N_3463);
or U4366 (N_4366,N_3242,N_3489);
or U4367 (N_4367,N_3014,N_3003);
nand U4368 (N_4368,N_3671,N_3328);
nand U4369 (N_4369,N_3837,N_3639);
or U4370 (N_4370,N_3035,N_3251);
nand U4371 (N_4371,N_3870,N_3677);
or U4372 (N_4372,N_3853,N_3437);
nor U4373 (N_4373,N_3915,N_3176);
or U4374 (N_4374,N_3086,N_3594);
xor U4375 (N_4375,N_3250,N_3986);
nor U4376 (N_4376,N_3944,N_3629);
xnor U4377 (N_4377,N_3953,N_3389);
nor U4378 (N_4378,N_3301,N_3909);
and U4379 (N_4379,N_3044,N_3879);
or U4380 (N_4380,N_3198,N_3824);
or U4381 (N_4381,N_3940,N_3956);
xnor U4382 (N_4382,N_3991,N_3042);
nor U4383 (N_4383,N_3329,N_3263);
nor U4384 (N_4384,N_3656,N_3371);
nand U4385 (N_4385,N_3209,N_3962);
or U4386 (N_4386,N_3643,N_3791);
or U4387 (N_4387,N_3441,N_3630);
nand U4388 (N_4388,N_3521,N_3912);
and U4389 (N_4389,N_3781,N_3907);
nor U4390 (N_4390,N_3529,N_3109);
and U4391 (N_4391,N_3478,N_3763);
nand U4392 (N_4392,N_3350,N_3450);
xnor U4393 (N_4393,N_3314,N_3298);
and U4394 (N_4394,N_3606,N_3416);
nor U4395 (N_4395,N_3157,N_3743);
nand U4396 (N_4396,N_3409,N_3663);
nand U4397 (N_4397,N_3241,N_3993);
or U4398 (N_4398,N_3840,N_3055);
and U4399 (N_4399,N_3520,N_3526);
xor U4400 (N_4400,N_3075,N_3375);
nand U4401 (N_4401,N_3142,N_3025);
nand U4402 (N_4402,N_3832,N_3453);
nand U4403 (N_4403,N_3221,N_3274);
nand U4404 (N_4404,N_3527,N_3461);
and U4405 (N_4405,N_3803,N_3507);
or U4406 (N_4406,N_3596,N_3041);
and U4407 (N_4407,N_3355,N_3958);
or U4408 (N_4408,N_3185,N_3515);
nand U4409 (N_4409,N_3428,N_3737);
xnor U4410 (N_4410,N_3290,N_3876);
nand U4411 (N_4411,N_3812,N_3858);
nand U4412 (N_4412,N_3689,N_3571);
nand U4413 (N_4413,N_3312,N_3857);
nor U4414 (N_4414,N_3177,N_3323);
nor U4415 (N_4415,N_3259,N_3749);
nor U4416 (N_4416,N_3405,N_3751);
nand U4417 (N_4417,N_3836,N_3317);
or U4418 (N_4418,N_3195,N_3124);
nand U4419 (N_4419,N_3816,N_3029);
and U4420 (N_4420,N_3553,N_3281);
nor U4421 (N_4421,N_3702,N_3309);
nor U4422 (N_4422,N_3276,N_3493);
nor U4423 (N_4423,N_3971,N_3590);
nor U4424 (N_4424,N_3733,N_3415);
or U4425 (N_4425,N_3179,N_3089);
nand U4426 (N_4426,N_3573,N_3729);
or U4427 (N_4427,N_3788,N_3681);
and U4428 (N_4428,N_3565,N_3466);
or U4429 (N_4429,N_3413,N_3794);
nor U4430 (N_4430,N_3227,N_3308);
nand U4431 (N_4431,N_3192,N_3561);
nand U4432 (N_4432,N_3407,N_3510);
nand U4433 (N_4433,N_3506,N_3286);
nand U4434 (N_4434,N_3551,N_3277);
nand U4435 (N_4435,N_3321,N_3802);
nand U4436 (N_4436,N_3692,N_3977);
or U4437 (N_4437,N_3094,N_3950);
nand U4438 (N_4438,N_3601,N_3569);
and U4439 (N_4439,N_3456,N_3449);
xor U4440 (N_4440,N_3846,N_3690);
or U4441 (N_4441,N_3509,N_3436);
or U4442 (N_4442,N_3299,N_3811);
nand U4443 (N_4443,N_3772,N_3782);
and U4444 (N_4444,N_3713,N_3147);
nor U4445 (N_4445,N_3246,N_3112);
xor U4446 (N_4446,N_3384,N_3442);
and U4447 (N_4447,N_3397,N_3748);
and U4448 (N_4448,N_3472,N_3001);
nor U4449 (N_4449,N_3884,N_3105);
nor U4450 (N_4450,N_3688,N_3649);
and U4451 (N_4451,N_3481,N_3063);
nor U4452 (N_4452,N_3805,N_3728);
or U4453 (N_4453,N_3374,N_3896);
xnor U4454 (N_4454,N_3121,N_3963);
and U4455 (N_4455,N_3588,N_3638);
nor U4456 (N_4456,N_3239,N_3888);
nor U4457 (N_4457,N_3906,N_3151);
nor U4458 (N_4458,N_3612,N_3369);
xor U4459 (N_4459,N_3850,N_3091);
nand U4460 (N_4460,N_3644,N_3911);
nand U4461 (N_4461,N_3164,N_3027);
or U4462 (N_4462,N_3615,N_3581);
nand U4463 (N_4463,N_3667,N_3597);
or U4464 (N_4464,N_3344,N_3547);
nor U4465 (N_4465,N_3703,N_3295);
and U4466 (N_4466,N_3530,N_3730);
nand U4467 (N_4467,N_3169,N_3162);
or U4468 (N_4468,N_3476,N_3626);
and U4469 (N_4469,N_3970,N_3116);
nor U4470 (N_4470,N_3101,N_3426);
and U4471 (N_4471,N_3943,N_3354);
nand U4472 (N_4472,N_3294,N_3217);
and U4473 (N_4473,N_3886,N_3253);
and U4474 (N_4474,N_3424,N_3668);
and U4475 (N_4475,N_3776,N_3634);
or U4476 (N_4476,N_3139,N_3033);
and U4477 (N_4477,N_3687,N_3797);
nor U4478 (N_4478,N_3881,N_3214);
nand U4479 (N_4479,N_3066,N_3996);
nor U4480 (N_4480,N_3338,N_3100);
nand U4481 (N_4481,N_3983,N_3844);
nor U4482 (N_4482,N_3757,N_3203);
nor U4483 (N_4483,N_3540,N_3988);
nand U4484 (N_4484,N_3134,N_3534);
xnor U4485 (N_4485,N_3057,N_3955);
nand U4486 (N_4486,N_3252,N_3960);
xor U4487 (N_4487,N_3180,N_3119);
xnor U4488 (N_4488,N_3004,N_3841);
nor U4489 (N_4489,N_3869,N_3156);
nand U4490 (N_4490,N_3353,N_3650);
xor U4491 (N_4491,N_3617,N_3610);
nor U4492 (N_4492,N_3078,N_3964);
xor U4493 (N_4493,N_3401,N_3120);
and U4494 (N_4494,N_3054,N_3093);
or U4495 (N_4495,N_3152,N_3406);
nor U4496 (N_4496,N_3265,N_3073);
nor U4497 (N_4497,N_3683,N_3982);
nor U4498 (N_4498,N_3069,N_3889);
and U4499 (N_4499,N_3670,N_3664);
xnor U4500 (N_4500,N_3006,N_3794);
nor U4501 (N_4501,N_3769,N_3692);
or U4502 (N_4502,N_3358,N_3496);
xnor U4503 (N_4503,N_3592,N_3079);
or U4504 (N_4504,N_3135,N_3001);
nand U4505 (N_4505,N_3099,N_3773);
or U4506 (N_4506,N_3481,N_3632);
or U4507 (N_4507,N_3163,N_3001);
nand U4508 (N_4508,N_3009,N_3526);
nand U4509 (N_4509,N_3038,N_3920);
nor U4510 (N_4510,N_3407,N_3213);
nand U4511 (N_4511,N_3579,N_3931);
nor U4512 (N_4512,N_3936,N_3515);
nor U4513 (N_4513,N_3864,N_3632);
nor U4514 (N_4514,N_3624,N_3761);
nor U4515 (N_4515,N_3700,N_3455);
nor U4516 (N_4516,N_3958,N_3475);
xnor U4517 (N_4517,N_3553,N_3029);
xnor U4518 (N_4518,N_3923,N_3791);
nand U4519 (N_4519,N_3141,N_3386);
or U4520 (N_4520,N_3782,N_3753);
and U4521 (N_4521,N_3004,N_3096);
nor U4522 (N_4522,N_3508,N_3464);
and U4523 (N_4523,N_3871,N_3037);
or U4524 (N_4524,N_3488,N_3502);
or U4525 (N_4525,N_3725,N_3339);
nor U4526 (N_4526,N_3694,N_3692);
nor U4527 (N_4527,N_3428,N_3968);
or U4528 (N_4528,N_3464,N_3144);
nor U4529 (N_4529,N_3750,N_3889);
nor U4530 (N_4530,N_3551,N_3791);
nor U4531 (N_4531,N_3687,N_3903);
or U4532 (N_4532,N_3408,N_3467);
nor U4533 (N_4533,N_3899,N_3938);
nand U4534 (N_4534,N_3661,N_3495);
or U4535 (N_4535,N_3618,N_3799);
or U4536 (N_4536,N_3206,N_3330);
nand U4537 (N_4537,N_3855,N_3025);
and U4538 (N_4538,N_3264,N_3027);
nor U4539 (N_4539,N_3149,N_3117);
nand U4540 (N_4540,N_3191,N_3219);
and U4541 (N_4541,N_3153,N_3362);
nor U4542 (N_4542,N_3832,N_3328);
or U4543 (N_4543,N_3484,N_3214);
and U4544 (N_4544,N_3649,N_3198);
or U4545 (N_4545,N_3385,N_3021);
and U4546 (N_4546,N_3628,N_3824);
or U4547 (N_4547,N_3218,N_3586);
and U4548 (N_4548,N_3620,N_3097);
nor U4549 (N_4549,N_3499,N_3492);
nor U4550 (N_4550,N_3370,N_3093);
and U4551 (N_4551,N_3412,N_3327);
xnor U4552 (N_4552,N_3052,N_3657);
xnor U4553 (N_4553,N_3626,N_3201);
nor U4554 (N_4554,N_3523,N_3403);
nor U4555 (N_4555,N_3058,N_3159);
xnor U4556 (N_4556,N_3075,N_3049);
nand U4557 (N_4557,N_3742,N_3617);
nor U4558 (N_4558,N_3733,N_3162);
xnor U4559 (N_4559,N_3917,N_3391);
and U4560 (N_4560,N_3543,N_3186);
and U4561 (N_4561,N_3251,N_3183);
and U4562 (N_4562,N_3168,N_3824);
nor U4563 (N_4563,N_3680,N_3444);
nand U4564 (N_4564,N_3727,N_3327);
or U4565 (N_4565,N_3173,N_3773);
or U4566 (N_4566,N_3413,N_3464);
or U4567 (N_4567,N_3680,N_3689);
nand U4568 (N_4568,N_3973,N_3552);
xnor U4569 (N_4569,N_3903,N_3720);
nor U4570 (N_4570,N_3609,N_3679);
nor U4571 (N_4571,N_3513,N_3052);
nor U4572 (N_4572,N_3765,N_3115);
or U4573 (N_4573,N_3907,N_3026);
xor U4574 (N_4574,N_3623,N_3225);
or U4575 (N_4575,N_3528,N_3688);
nand U4576 (N_4576,N_3794,N_3645);
xnor U4577 (N_4577,N_3313,N_3404);
and U4578 (N_4578,N_3824,N_3325);
and U4579 (N_4579,N_3766,N_3821);
nand U4580 (N_4580,N_3169,N_3530);
nand U4581 (N_4581,N_3275,N_3868);
nand U4582 (N_4582,N_3075,N_3265);
xnor U4583 (N_4583,N_3733,N_3251);
or U4584 (N_4584,N_3748,N_3269);
or U4585 (N_4585,N_3613,N_3679);
nand U4586 (N_4586,N_3940,N_3380);
xor U4587 (N_4587,N_3203,N_3736);
nand U4588 (N_4588,N_3437,N_3169);
and U4589 (N_4589,N_3373,N_3614);
and U4590 (N_4590,N_3834,N_3899);
and U4591 (N_4591,N_3652,N_3902);
nand U4592 (N_4592,N_3013,N_3284);
xnor U4593 (N_4593,N_3153,N_3585);
and U4594 (N_4594,N_3268,N_3207);
nor U4595 (N_4595,N_3432,N_3155);
or U4596 (N_4596,N_3254,N_3544);
and U4597 (N_4597,N_3386,N_3613);
nand U4598 (N_4598,N_3789,N_3567);
and U4599 (N_4599,N_3108,N_3650);
or U4600 (N_4600,N_3790,N_3097);
and U4601 (N_4601,N_3085,N_3804);
nor U4602 (N_4602,N_3150,N_3091);
nand U4603 (N_4603,N_3000,N_3584);
nor U4604 (N_4604,N_3672,N_3611);
and U4605 (N_4605,N_3363,N_3264);
or U4606 (N_4606,N_3508,N_3308);
or U4607 (N_4607,N_3082,N_3168);
nor U4608 (N_4608,N_3789,N_3644);
nor U4609 (N_4609,N_3791,N_3602);
nand U4610 (N_4610,N_3475,N_3035);
nor U4611 (N_4611,N_3858,N_3484);
nand U4612 (N_4612,N_3688,N_3076);
or U4613 (N_4613,N_3544,N_3346);
nand U4614 (N_4614,N_3056,N_3232);
or U4615 (N_4615,N_3915,N_3083);
and U4616 (N_4616,N_3176,N_3214);
nor U4617 (N_4617,N_3547,N_3900);
or U4618 (N_4618,N_3529,N_3070);
and U4619 (N_4619,N_3284,N_3939);
nand U4620 (N_4620,N_3332,N_3473);
and U4621 (N_4621,N_3268,N_3035);
nor U4622 (N_4622,N_3595,N_3755);
or U4623 (N_4623,N_3939,N_3918);
and U4624 (N_4624,N_3570,N_3430);
and U4625 (N_4625,N_3308,N_3609);
nand U4626 (N_4626,N_3654,N_3851);
nand U4627 (N_4627,N_3968,N_3422);
nor U4628 (N_4628,N_3047,N_3560);
and U4629 (N_4629,N_3977,N_3795);
or U4630 (N_4630,N_3232,N_3880);
nand U4631 (N_4631,N_3778,N_3650);
nand U4632 (N_4632,N_3621,N_3130);
nor U4633 (N_4633,N_3020,N_3264);
nand U4634 (N_4634,N_3245,N_3252);
nor U4635 (N_4635,N_3606,N_3953);
nand U4636 (N_4636,N_3996,N_3246);
and U4637 (N_4637,N_3738,N_3782);
and U4638 (N_4638,N_3510,N_3499);
and U4639 (N_4639,N_3816,N_3227);
nor U4640 (N_4640,N_3612,N_3143);
and U4641 (N_4641,N_3189,N_3208);
nand U4642 (N_4642,N_3835,N_3203);
or U4643 (N_4643,N_3908,N_3482);
and U4644 (N_4644,N_3793,N_3352);
xor U4645 (N_4645,N_3640,N_3004);
nand U4646 (N_4646,N_3068,N_3025);
or U4647 (N_4647,N_3939,N_3055);
and U4648 (N_4648,N_3389,N_3249);
nand U4649 (N_4649,N_3139,N_3829);
nor U4650 (N_4650,N_3865,N_3313);
nor U4651 (N_4651,N_3828,N_3729);
or U4652 (N_4652,N_3313,N_3725);
xnor U4653 (N_4653,N_3016,N_3518);
and U4654 (N_4654,N_3852,N_3251);
nor U4655 (N_4655,N_3722,N_3434);
nor U4656 (N_4656,N_3816,N_3850);
or U4657 (N_4657,N_3539,N_3128);
nand U4658 (N_4658,N_3326,N_3018);
nand U4659 (N_4659,N_3459,N_3513);
and U4660 (N_4660,N_3747,N_3728);
nand U4661 (N_4661,N_3122,N_3921);
nand U4662 (N_4662,N_3489,N_3146);
and U4663 (N_4663,N_3852,N_3762);
nor U4664 (N_4664,N_3131,N_3407);
and U4665 (N_4665,N_3260,N_3165);
nor U4666 (N_4666,N_3320,N_3438);
nor U4667 (N_4667,N_3979,N_3624);
nand U4668 (N_4668,N_3074,N_3490);
nand U4669 (N_4669,N_3202,N_3611);
nor U4670 (N_4670,N_3799,N_3453);
or U4671 (N_4671,N_3927,N_3266);
nand U4672 (N_4672,N_3938,N_3019);
nor U4673 (N_4673,N_3133,N_3818);
nand U4674 (N_4674,N_3114,N_3483);
nand U4675 (N_4675,N_3253,N_3831);
nand U4676 (N_4676,N_3665,N_3789);
nand U4677 (N_4677,N_3848,N_3969);
xnor U4678 (N_4678,N_3918,N_3138);
nor U4679 (N_4679,N_3702,N_3202);
nand U4680 (N_4680,N_3233,N_3616);
nor U4681 (N_4681,N_3595,N_3116);
and U4682 (N_4682,N_3096,N_3037);
and U4683 (N_4683,N_3716,N_3336);
or U4684 (N_4684,N_3089,N_3687);
nor U4685 (N_4685,N_3174,N_3798);
nor U4686 (N_4686,N_3858,N_3396);
nor U4687 (N_4687,N_3473,N_3047);
nor U4688 (N_4688,N_3726,N_3896);
and U4689 (N_4689,N_3467,N_3327);
or U4690 (N_4690,N_3486,N_3299);
and U4691 (N_4691,N_3142,N_3395);
or U4692 (N_4692,N_3742,N_3804);
nor U4693 (N_4693,N_3924,N_3256);
and U4694 (N_4694,N_3505,N_3468);
nor U4695 (N_4695,N_3830,N_3926);
xnor U4696 (N_4696,N_3651,N_3653);
and U4697 (N_4697,N_3760,N_3442);
nor U4698 (N_4698,N_3717,N_3212);
and U4699 (N_4699,N_3856,N_3771);
nand U4700 (N_4700,N_3863,N_3418);
nor U4701 (N_4701,N_3016,N_3230);
nand U4702 (N_4702,N_3280,N_3073);
nor U4703 (N_4703,N_3106,N_3772);
nor U4704 (N_4704,N_3167,N_3263);
or U4705 (N_4705,N_3126,N_3562);
and U4706 (N_4706,N_3384,N_3573);
and U4707 (N_4707,N_3085,N_3221);
and U4708 (N_4708,N_3119,N_3560);
or U4709 (N_4709,N_3223,N_3446);
nand U4710 (N_4710,N_3270,N_3694);
and U4711 (N_4711,N_3141,N_3435);
nand U4712 (N_4712,N_3517,N_3788);
nand U4713 (N_4713,N_3438,N_3927);
or U4714 (N_4714,N_3423,N_3867);
and U4715 (N_4715,N_3818,N_3427);
nor U4716 (N_4716,N_3700,N_3005);
nor U4717 (N_4717,N_3681,N_3319);
xor U4718 (N_4718,N_3570,N_3184);
and U4719 (N_4719,N_3096,N_3440);
and U4720 (N_4720,N_3215,N_3509);
nand U4721 (N_4721,N_3512,N_3151);
or U4722 (N_4722,N_3200,N_3497);
and U4723 (N_4723,N_3252,N_3888);
and U4724 (N_4724,N_3371,N_3905);
or U4725 (N_4725,N_3235,N_3475);
nand U4726 (N_4726,N_3448,N_3422);
or U4727 (N_4727,N_3656,N_3609);
and U4728 (N_4728,N_3697,N_3165);
and U4729 (N_4729,N_3457,N_3906);
or U4730 (N_4730,N_3091,N_3474);
nand U4731 (N_4731,N_3897,N_3523);
nor U4732 (N_4732,N_3028,N_3944);
nor U4733 (N_4733,N_3002,N_3674);
nand U4734 (N_4734,N_3233,N_3857);
nor U4735 (N_4735,N_3086,N_3026);
nor U4736 (N_4736,N_3341,N_3049);
or U4737 (N_4737,N_3998,N_3520);
nor U4738 (N_4738,N_3119,N_3809);
or U4739 (N_4739,N_3365,N_3636);
nand U4740 (N_4740,N_3171,N_3309);
nand U4741 (N_4741,N_3046,N_3213);
xnor U4742 (N_4742,N_3823,N_3831);
and U4743 (N_4743,N_3274,N_3715);
nor U4744 (N_4744,N_3576,N_3524);
xor U4745 (N_4745,N_3566,N_3526);
nand U4746 (N_4746,N_3836,N_3982);
and U4747 (N_4747,N_3633,N_3323);
nand U4748 (N_4748,N_3060,N_3964);
and U4749 (N_4749,N_3603,N_3168);
or U4750 (N_4750,N_3466,N_3768);
nor U4751 (N_4751,N_3244,N_3619);
and U4752 (N_4752,N_3485,N_3797);
nand U4753 (N_4753,N_3311,N_3041);
nor U4754 (N_4754,N_3536,N_3634);
or U4755 (N_4755,N_3083,N_3511);
nor U4756 (N_4756,N_3698,N_3232);
xnor U4757 (N_4757,N_3584,N_3469);
nor U4758 (N_4758,N_3284,N_3753);
and U4759 (N_4759,N_3866,N_3063);
nand U4760 (N_4760,N_3941,N_3369);
or U4761 (N_4761,N_3323,N_3643);
and U4762 (N_4762,N_3998,N_3985);
nand U4763 (N_4763,N_3950,N_3662);
or U4764 (N_4764,N_3371,N_3311);
xnor U4765 (N_4765,N_3627,N_3899);
nor U4766 (N_4766,N_3029,N_3374);
and U4767 (N_4767,N_3274,N_3168);
xor U4768 (N_4768,N_3244,N_3938);
nand U4769 (N_4769,N_3659,N_3908);
nor U4770 (N_4770,N_3265,N_3661);
nor U4771 (N_4771,N_3015,N_3076);
or U4772 (N_4772,N_3392,N_3520);
nand U4773 (N_4773,N_3095,N_3703);
nand U4774 (N_4774,N_3874,N_3461);
xor U4775 (N_4775,N_3014,N_3965);
or U4776 (N_4776,N_3762,N_3945);
xor U4777 (N_4777,N_3422,N_3854);
or U4778 (N_4778,N_3537,N_3892);
or U4779 (N_4779,N_3520,N_3336);
or U4780 (N_4780,N_3954,N_3346);
nor U4781 (N_4781,N_3821,N_3944);
nor U4782 (N_4782,N_3065,N_3462);
nand U4783 (N_4783,N_3076,N_3293);
or U4784 (N_4784,N_3450,N_3612);
xor U4785 (N_4785,N_3623,N_3834);
and U4786 (N_4786,N_3377,N_3885);
and U4787 (N_4787,N_3121,N_3049);
and U4788 (N_4788,N_3684,N_3071);
nor U4789 (N_4789,N_3846,N_3029);
nor U4790 (N_4790,N_3127,N_3072);
and U4791 (N_4791,N_3770,N_3664);
xor U4792 (N_4792,N_3065,N_3987);
or U4793 (N_4793,N_3690,N_3132);
and U4794 (N_4794,N_3018,N_3467);
or U4795 (N_4795,N_3134,N_3326);
and U4796 (N_4796,N_3019,N_3652);
and U4797 (N_4797,N_3551,N_3080);
and U4798 (N_4798,N_3637,N_3578);
nor U4799 (N_4799,N_3282,N_3426);
or U4800 (N_4800,N_3615,N_3464);
nor U4801 (N_4801,N_3735,N_3860);
nand U4802 (N_4802,N_3038,N_3897);
and U4803 (N_4803,N_3520,N_3346);
xor U4804 (N_4804,N_3751,N_3757);
xor U4805 (N_4805,N_3160,N_3422);
or U4806 (N_4806,N_3464,N_3111);
xnor U4807 (N_4807,N_3934,N_3478);
nand U4808 (N_4808,N_3425,N_3331);
or U4809 (N_4809,N_3533,N_3573);
or U4810 (N_4810,N_3437,N_3841);
nand U4811 (N_4811,N_3304,N_3379);
or U4812 (N_4812,N_3545,N_3382);
xor U4813 (N_4813,N_3731,N_3683);
nor U4814 (N_4814,N_3485,N_3185);
nor U4815 (N_4815,N_3816,N_3452);
and U4816 (N_4816,N_3936,N_3020);
nor U4817 (N_4817,N_3420,N_3362);
nor U4818 (N_4818,N_3656,N_3280);
or U4819 (N_4819,N_3244,N_3892);
and U4820 (N_4820,N_3094,N_3960);
xnor U4821 (N_4821,N_3782,N_3597);
nand U4822 (N_4822,N_3223,N_3992);
and U4823 (N_4823,N_3430,N_3823);
or U4824 (N_4824,N_3542,N_3252);
or U4825 (N_4825,N_3958,N_3802);
nand U4826 (N_4826,N_3718,N_3569);
nor U4827 (N_4827,N_3156,N_3703);
nand U4828 (N_4828,N_3656,N_3130);
nor U4829 (N_4829,N_3723,N_3786);
or U4830 (N_4830,N_3064,N_3861);
nor U4831 (N_4831,N_3116,N_3657);
nor U4832 (N_4832,N_3666,N_3195);
and U4833 (N_4833,N_3637,N_3383);
nor U4834 (N_4834,N_3392,N_3930);
and U4835 (N_4835,N_3680,N_3289);
xnor U4836 (N_4836,N_3669,N_3560);
nor U4837 (N_4837,N_3080,N_3278);
nor U4838 (N_4838,N_3674,N_3489);
nor U4839 (N_4839,N_3756,N_3340);
and U4840 (N_4840,N_3164,N_3393);
nor U4841 (N_4841,N_3163,N_3324);
or U4842 (N_4842,N_3672,N_3631);
or U4843 (N_4843,N_3466,N_3341);
and U4844 (N_4844,N_3063,N_3654);
nand U4845 (N_4845,N_3993,N_3142);
or U4846 (N_4846,N_3648,N_3797);
nand U4847 (N_4847,N_3452,N_3508);
nor U4848 (N_4848,N_3478,N_3246);
nor U4849 (N_4849,N_3960,N_3649);
nor U4850 (N_4850,N_3770,N_3008);
nand U4851 (N_4851,N_3600,N_3729);
nand U4852 (N_4852,N_3590,N_3563);
nand U4853 (N_4853,N_3766,N_3333);
and U4854 (N_4854,N_3937,N_3734);
nor U4855 (N_4855,N_3789,N_3016);
and U4856 (N_4856,N_3766,N_3689);
nand U4857 (N_4857,N_3357,N_3643);
or U4858 (N_4858,N_3681,N_3421);
nand U4859 (N_4859,N_3573,N_3138);
nor U4860 (N_4860,N_3503,N_3611);
or U4861 (N_4861,N_3836,N_3418);
and U4862 (N_4862,N_3950,N_3885);
nor U4863 (N_4863,N_3656,N_3273);
nor U4864 (N_4864,N_3143,N_3274);
nor U4865 (N_4865,N_3564,N_3274);
nor U4866 (N_4866,N_3287,N_3417);
or U4867 (N_4867,N_3422,N_3289);
nor U4868 (N_4868,N_3199,N_3661);
and U4869 (N_4869,N_3042,N_3918);
or U4870 (N_4870,N_3552,N_3068);
xor U4871 (N_4871,N_3540,N_3877);
and U4872 (N_4872,N_3152,N_3270);
nand U4873 (N_4873,N_3751,N_3019);
or U4874 (N_4874,N_3545,N_3103);
nand U4875 (N_4875,N_3210,N_3331);
nor U4876 (N_4876,N_3057,N_3558);
nand U4877 (N_4877,N_3359,N_3764);
nand U4878 (N_4878,N_3424,N_3284);
nor U4879 (N_4879,N_3803,N_3791);
xor U4880 (N_4880,N_3978,N_3824);
nor U4881 (N_4881,N_3564,N_3093);
or U4882 (N_4882,N_3227,N_3418);
and U4883 (N_4883,N_3809,N_3721);
nand U4884 (N_4884,N_3340,N_3871);
nor U4885 (N_4885,N_3544,N_3484);
xor U4886 (N_4886,N_3310,N_3840);
xnor U4887 (N_4887,N_3337,N_3343);
and U4888 (N_4888,N_3416,N_3809);
nand U4889 (N_4889,N_3766,N_3831);
nor U4890 (N_4890,N_3950,N_3629);
nand U4891 (N_4891,N_3612,N_3913);
and U4892 (N_4892,N_3574,N_3965);
nand U4893 (N_4893,N_3906,N_3676);
and U4894 (N_4894,N_3969,N_3544);
and U4895 (N_4895,N_3669,N_3205);
xnor U4896 (N_4896,N_3288,N_3608);
xnor U4897 (N_4897,N_3347,N_3283);
nor U4898 (N_4898,N_3404,N_3645);
xnor U4899 (N_4899,N_3847,N_3505);
or U4900 (N_4900,N_3134,N_3985);
and U4901 (N_4901,N_3284,N_3987);
nor U4902 (N_4902,N_3323,N_3276);
nor U4903 (N_4903,N_3457,N_3044);
nand U4904 (N_4904,N_3874,N_3566);
or U4905 (N_4905,N_3672,N_3401);
nor U4906 (N_4906,N_3249,N_3489);
nor U4907 (N_4907,N_3025,N_3620);
and U4908 (N_4908,N_3867,N_3313);
nor U4909 (N_4909,N_3889,N_3064);
or U4910 (N_4910,N_3017,N_3690);
xor U4911 (N_4911,N_3146,N_3954);
nand U4912 (N_4912,N_3827,N_3190);
xnor U4913 (N_4913,N_3573,N_3388);
xor U4914 (N_4914,N_3323,N_3521);
nor U4915 (N_4915,N_3214,N_3788);
and U4916 (N_4916,N_3491,N_3353);
or U4917 (N_4917,N_3311,N_3045);
nand U4918 (N_4918,N_3268,N_3982);
xnor U4919 (N_4919,N_3244,N_3558);
nand U4920 (N_4920,N_3569,N_3855);
nand U4921 (N_4921,N_3215,N_3603);
and U4922 (N_4922,N_3184,N_3146);
or U4923 (N_4923,N_3136,N_3909);
or U4924 (N_4924,N_3360,N_3963);
and U4925 (N_4925,N_3943,N_3651);
or U4926 (N_4926,N_3357,N_3814);
and U4927 (N_4927,N_3086,N_3297);
nor U4928 (N_4928,N_3512,N_3524);
nor U4929 (N_4929,N_3118,N_3499);
and U4930 (N_4930,N_3640,N_3422);
nor U4931 (N_4931,N_3501,N_3116);
nand U4932 (N_4932,N_3007,N_3430);
nand U4933 (N_4933,N_3103,N_3160);
xor U4934 (N_4934,N_3557,N_3834);
nor U4935 (N_4935,N_3102,N_3795);
nand U4936 (N_4936,N_3350,N_3381);
and U4937 (N_4937,N_3874,N_3650);
xor U4938 (N_4938,N_3249,N_3604);
nand U4939 (N_4939,N_3987,N_3561);
nor U4940 (N_4940,N_3931,N_3745);
and U4941 (N_4941,N_3699,N_3480);
nor U4942 (N_4942,N_3054,N_3444);
nand U4943 (N_4943,N_3618,N_3562);
nand U4944 (N_4944,N_3176,N_3797);
or U4945 (N_4945,N_3792,N_3835);
or U4946 (N_4946,N_3734,N_3221);
or U4947 (N_4947,N_3089,N_3288);
and U4948 (N_4948,N_3016,N_3348);
or U4949 (N_4949,N_3831,N_3829);
and U4950 (N_4950,N_3990,N_3589);
nor U4951 (N_4951,N_3259,N_3356);
nor U4952 (N_4952,N_3639,N_3382);
and U4953 (N_4953,N_3703,N_3506);
and U4954 (N_4954,N_3704,N_3093);
nand U4955 (N_4955,N_3763,N_3484);
or U4956 (N_4956,N_3181,N_3443);
nor U4957 (N_4957,N_3755,N_3810);
and U4958 (N_4958,N_3079,N_3078);
and U4959 (N_4959,N_3348,N_3518);
and U4960 (N_4960,N_3696,N_3152);
and U4961 (N_4961,N_3671,N_3634);
nand U4962 (N_4962,N_3205,N_3039);
nor U4963 (N_4963,N_3130,N_3240);
nand U4964 (N_4964,N_3789,N_3687);
or U4965 (N_4965,N_3422,N_3294);
or U4966 (N_4966,N_3519,N_3133);
nor U4967 (N_4967,N_3519,N_3624);
nand U4968 (N_4968,N_3237,N_3858);
nor U4969 (N_4969,N_3849,N_3609);
nand U4970 (N_4970,N_3670,N_3346);
nor U4971 (N_4971,N_3810,N_3775);
and U4972 (N_4972,N_3547,N_3971);
nand U4973 (N_4973,N_3803,N_3024);
and U4974 (N_4974,N_3509,N_3000);
and U4975 (N_4975,N_3447,N_3354);
nor U4976 (N_4976,N_3326,N_3594);
and U4977 (N_4977,N_3733,N_3158);
or U4978 (N_4978,N_3134,N_3879);
or U4979 (N_4979,N_3722,N_3702);
or U4980 (N_4980,N_3568,N_3065);
or U4981 (N_4981,N_3171,N_3497);
and U4982 (N_4982,N_3789,N_3420);
nand U4983 (N_4983,N_3848,N_3697);
nor U4984 (N_4984,N_3747,N_3448);
xnor U4985 (N_4985,N_3772,N_3111);
and U4986 (N_4986,N_3234,N_3929);
or U4987 (N_4987,N_3517,N_3388);
or U4988 (N_4988,N_3841,N_3784);
xor U4989 (N_4989,N_3334,N_3032);
xnor U4990 (N_4990,N_3491,N_3191);
nor U4991 (N_4991,N_3041,N_3717);
nand U4992 (N_4992,N_3909,N_3302);
and U4993 (N_4993,N_3817,N_3148);
nand U4994 (N_4994,N_3084,N_3338);
and U4995 (N_4995,N_3930,N_3781);
or U4996 (N_4996,N_3805,N_3355);
nand U4997 (N_4997,N_3810,N_3087);
or U4998 (N_4998,N_3886,N_3511);
xor U4999 (N_4999,N_3870,N_3806);
and UO_0 (O_0,N_4903,N_4108);
nand UO_1 (O_1,N_4436,N_4761);
or UO_2 (O_2,N_4719,N_4043);
or UO_3 (O_3,N_4412,N_4075);
and UO_4 (O_4,N_4435,N_4013);
nor UO_5 (O_5,N_4994,N_4393);
and UO_6 (O_6,N_4301,N_4225);
and UO_7 (O_7,N_4609,N_4327);
or UO_8 (O_8,N_4593,N_4131);
xnor UO_9 (O_9,N_4129,N_4190);
nand UO_10 (O_10,N_4360,N_4828);
nand UO_11 (O_11,N_4857,N_4434);
and UO_12 (O_12,N_4232,N_4291);
nand UO_13 (O_13,N_4637,N_4362);
and UO_14 (O_14,N_4069,N_4230);
or UO_15 (O_15,N_4364,N_4368);
and UO_16 (O_16,N_4711,N_4862);
or UO_17 (O_17,N_4428,N_4749);
nand UO_18 (O_18,N_4779,N_4509);
xor UO_19 (O_19,N_4197,N_4198);
or UO_20 (O_20,N_4625,N_4841);
nor UO_21 (O_21,N_4599,N_4475);
or UO_22 (O_22,N_4326,N_4164);
or UO_23 (O_23,N_4872,N_4924);
and UO_24 (O_24,N_4552,N_4682);
nor UO_25 (O_25,N_4695,N_4688);
nor UO_26 (O_26,N_4864,N_4910);
or UO_27 (O_27,N_4624,N_4716);
or UO_28 (O_28,N_4135,N_4298);
nand UO_29 (O_29,N_4212,N_4259);
or UO_30 (O_30,N_4242,N_4406);
nor UO_31 (O_31,N_4904,N_4105);
or UO_32 (O_32,N_4549,N_4087);
or UO_33 (O_33,N_4438,N_4827);
nor UO_34 (O_34,N_4618,N_4104);
nand UO_35 (O_35,N_4751,N_4600);
nor UO_36 (O_36,N_4034,N_4630);
nand UO_37 (O_37,N_4317,N_4532);
nand UO_38 (O_38,N_4037,N_4257);
or UO_39 (O_39,N_4134,N_4830);
nor UO_40 (O_40,N_4781,N_4112);
xor UO_41 (O_41,N_4268,N_4589);
and UO_42 (O_42,N_4775,N_4491);
nand UO_43 (O_43,N_4742,N_4014);
or UO_44 (O_44,N_4502,N_4889);
or UO_45 (O_45,N_4739,N_4539);
nor UO_46 (O_46,N_4359,N_4165);
xnor UO_47 (O_47,N_4080,N_4656);
nand UO_48 (O_48,N_4991,N_4885);
and UO_49 (O_49,N_4495,N_4420);
xor UO_50 (O_50,N_4223,N_4640);
nor UO_51 (O_51,N_4469,N_4285);
nand UO_52 (O_52,N_4768,N_4005);
and UO_53 (O_53,N_4059,N_4896);
nand UO_54 (O_54,N_4562,N_4633);
nand UO_55 (O_55,N_4363,N_4806);
and UO_56 (O_56,N_4934,N_4559);
xor UO_57 (O_57,N_4295,N_4673);
nand UO_58 (O_58,N_4990,N_4208);
nand UO_59 (O_59,N_4842,N_4708);
and UO_60 (O_60,N_4173,N_4721);
nor UO_61 (O_61,N_4747,N_4477);
and UO_62 (O_62,N_4323,N_4400);
nor UO_63 (O_63,N_4905,N_4643);
nor UO_64 (O_64,N_4329,N_4355);
and UO_65 (O_65,N_4963,N_4535);
nor UO_66 (O_66,N_4047,N_4764);
nand UO_67 (O_67,N_4382,N_4531);
or UO_68 (O_68,N_4856,N_4750);
and UO_69 (O_69,N_4098,N_4283);
and UO_70 (O_70,N_4540,N_4243);
and UO_71 (O_71,N_4703,N_4201);
nor UO_72 (O_72,N_4163,N_4100);
or UO_73 (O_73,N_4451,N_4151);
nand UO_74 (O_74,N_4762,N_4726);
nand UO_75 (O_75,N_4691,N_4858);
nand UO_76 (O_76,N_4456,N_4648);
nor UO_77 (O_77,N_4012,N_4373);
or UO_78 (O_78,N_4962,N_4709);
nand UO_79 (O_79,N_4217,N_4187);
and UO_80 (O_80,N_4063,N_4122);
or UO_81 (O_81,N_4769,N_4686);
nor UO_82 (O_82,N_4678,N_4140);
or UO_83 (O_83,N_4398,N_4838);
nor UO_84 (O_84,N_4950,N_4661);
nand UO_85 (O_85,N_4748,N_4229);
or UO_86 (O_86,N_4483,N_4818);
or UO_87 (O_87,N_4040,N_4000);
nor UO_88 (O_88,N_4794,N_4632);
nand UO_89 (O_89,N_4979,N_4580);
nor UO_90 (O_90,N_4961,N_4426);
nand UO_91 (O_91,N_4654,N_4055);
nand UO_92 (O_92,N_4044,N_4925);
or UO_93 (O_93,N_4732,N_4567);
nand UO_94 (O_94,N_4563,N_4556);
nor UO_95 (O_95,N_4999,N_4003);
nor UO_96 (O_96,N_4763,N_4579);
xnor UO_97 (O_97,N_4124,N_4333);
or UO_98 (O_98,N_4976,N_4227);
or UO_99 (O_99,N_4465,N_4349);
nor UO_100 (O_100,N_4597,N_4578);
nand UO_101 (O_101,N_4353,N_4148);
xor UO_102 (O_102,N_4615,N_4712);
nand UO_103 (O_103,N_4136,N_4078);
nand UO_104 (O_104,N_4448,N_4462);
or UO_105 (O_105,N_4265,N_4161);
and UO_106 (O_106,N_4753,N_4536);
and UO_107 (O_107,N_4146,N_4141);
or UO_108 (O_108,N_4162,N_4029);
nor UO_109 (O_109,N_4541,N_4423);
xor UO_110 (O_110,N_4236,N_4452);
nor UO_111 (O_111,N_4667,N_4743);
or UO_112 (O_112,N_4677,N_4613);
and UO_113 (O_113,N_4083,N_4304);
and UO_114 (O_114,N_4402,N_4320);
and UO_115 (O_115,N_4530,N_4825);
nand UO_116 (O_116,N_4193,N_4226);
nand UO_117 (O_117,N_4516,N_4346);
nor UO_118 (O_118,N_4777,N_4394);
nand UO_119 (O_119,N_4693,N_4370);
and UO_120 (O_120,N_4094,N_4901);
and UO_121 (O_121,N_4981,N_4812);
nand UO_122 (O_122,N_4046,N_4590);
or UO_123 (O_123,N_4286,N_4453);
and UO_124 (O_124,N_4879,N_4202);
nand UO_125 (O_125,N_4365,N_4045);
xnor UO_126 (O_126,N_4287,N_4916);
nand UO_127 (O_127,N_4868,N_4391);
and UO_128 (O_128,N_4154,N_4074);
nor UO_129 (O_129,N_4143,N_4185);
and UO_130 (O_130,N_4690,N_4417);
nand UO_131 (O_131,N_4321,N_4472);
nand UO_132 (O_132,N_4199,N_4132);
nor UO_133 (O_133,N_4808,N_4622);
xor UO_134 (O_134,N_4289,N_4432);
or UO_135 (O_135,N_4527,N_4926);
nand UO_136 (O_136,N_4238,N_4011);
or UO_137 (O_137,N_4819,N_4987);
nand UO_138 (O_138,N_4036,N_4966);
or UO_139 (O_139,N_4324,N_4817);
or UO_140 (O_140,N_4514,N_4120);
nand UO_141 (O_141,N_4026,N_4731);
nor UO_142 (O_142,N_4487,N_4687);
and UO_143 (O_143,N_4008,N_4115);
and UO_144 (O_144,N_4486,N_4325);
xor UO_145 (O_145,N_4805,N_4672);
and UO_146 (O_146,N_4574,N_4490);
and UO_147 (O_147,N_4376,N_4262);
or UO_148 (O_148,N_4809,N_4922);
or UO_149 (O_149,N_4255,N_4454);
and UO_150 (O_150,N_4529,N_4065);
nand UO_151 (O_151,N_4607,N_4671);
nor UO_152 (O_152,N_4821,N_4947);
or UO_153 (O_153,N_4499,N_4788);
nand UO_154 (O_154,N_4085,N_4553);
nor UO_155 (O_155,N_4783,N_4109);
xnor UO_156 (O_156,N_4649,N_4839);
and UO_157 (O_157,N_4224,N_4663);
xor UO_158 (O_158,N_4016,N_4829);
and UO_159 (O_159,N_4389,N_4729);
and UO_160 (O_160,N_4538,N_4493);
xor UO_161 (O_161,N_4873,N_4284);
nor UO_162 (O_162,N_4964,N_4342);
nor UO_163 (O_163,N_4117,N_4049);
or UO_164 (O_164,N_4652,N_4585);
or UO_165 (O_165,N_4082,N_4347);
nand UO_166 (O_166,N_4513,N_4666);
nand UO_167 (O_167,N_4431,N_4089);
and UO_168 (O_168,N_4754,N_4179);
or UO_169 (O_169,N_4339,N_4644);
and UO_170 (O_170,N_4523,N_4852);
or UO_171 (O_171,N_4031,N_4911);
or UO_172 (O_172,N_4820,N_4378);
or UO_173 (O_173,N_4586,N_4997);
and UO_174 (O_174,N_4114,N_4528);
and UO_175 (O_175,N_4815,N_4623);
and UO_176 (O_176,N_4066,N_4292);
xnor UO_177 (O_177,N_4883,N_4791);
nand UO_178 (O_178,N_4878,N_4930);
nand UO_179 (O_179,N_4650,N_4366);
nor UO_180 (O_180,N_4959,N_4077);
and UO_181 (O_181,N_4471,N_4575);
nor UO_182 (O_182,N_4282,N_4494);
or UO_183 (O_183,N_4641,N_4955);
and UO_184 (O_184,N_4273,N_4890);
nor UO_185 (O_185,N_4315,N_4773);
and UO_186 (O_186,N_4480,N_4511);
nand UO_187 (O_187,N_4522,N_4311);
or UO_188 (O_188,N_4091,N_4935);
and UO_189 (O_189,N_4568,N_4174);
and UO_190 (O_190,N_4070,N_4944);
nand UO_191 (O_191,N_4679,N_4107);
nor UO_192 (O_192,N_4694,N_4081);
or UO_193 (O_193,N_4537,N_4032);
and UO_194 (O_194,N_4022,N_4621);
nand UO_195 (O_195,N_4172,N_4571);
nand UO_196 (O_196,N_4488,N_4847);
nand UO_197 (O_197,N_4388,N_4209);
nor UO_198 (O_198,N_4759,N_4334);
nand UO_199 (O_199,N_4440,N_4021);
nor UO_200 (O_200,N_4980,N_4802);
nand UO_201 (O_201,N_4598,N_4772);
or UO_202 (O_202,N_4738,N_4581);
or UO_203 (O_203,N_4845,N_4949);
nor UO_204 (O_204,N_4627,N_4237);
nor UO_205 (O_205,N_4848,N_4205);
or UO_206 (O_206,N_4241,N_4125);
or UO_207 (O_207,N_4737,N_4655);
nor UO_208 (O_208,N_4002,N_4051);
nor UO_209 (O_209,N_4908,N_4181);
and UO_210 (O_210,N_4390,N_4042);
or UO_211 (O_211,N_4776,N_4706);
nand UO_212 (O_212,N_4826,N_4533);
and UO_213 (O_213,N_4720,N_4084);
nand UO_214 (O_214,N_4657,N_4584);
nor UO_215 (O_215,N_4337,N_4024);
nand UO_216 (O_216,N_4459,N_4573);
xnor UO_217 (O_217,N_4191,N_4534);
and UO_218 (O_218,N_4468,N_4372);
nand UO_219 (O_219,N_4504,N_4269);
and UO_220 (O_220,N_4127,N_4917);
or UO_221 (O_221,N_4741,N_4492);
and UO_222 (O_222,N_4410,N_4211);
xnor UO_223 (O_223,N_4204,N_4860);
nor UO_224 (O_224,N_4796,N_4811);
and UO_225 (O_225,N_4369,N_4119);
and UO_226 (O_226,N_4923,N_4875);
nor UO_227 (O_227,N_4668,N_4272);
nand UO_228 (O_228,N_4893,N_4007);
xor UO_229 (O_229,N_4906,N_4251);
nor UO_230 (O_230,N_4415,N_4614);
nand UO_231 (O_231,N_4702,N_4548);
or UO_232 (O_232,N_4921,N_4318);
and UO_233 (O_233,N_4439,N_4728);
and UO_234 (O_234,N_4348,N_4116);
nor UO_235 (O_235,N_4912,N_4833);
or UO_236 (O_236,N_4167,N_4096);
nand UO_237 (O_237,N_4130,N_4744);
or UO_238 (O_238,N_4060,N_4928);
xor UO_239 (O_239,N_4079,N_4027);
or UO_240 (O_240,N_4258,N_4458);
nand UO_241 (O_241,N_4009,N_4793);
and UO_242 (O_242,N_4447,N_4631);
xnor UO_243 (O_243,N_4700,N_4658);
or UO_244 (O_244,N_4110,N_4416);
and UO_245 (O_245,N_4968,N_4379);
or UO_246 (O_246,N_4844,N_4300);
xnor UO_247 (O_247,N_4951,N_4445);
and UO_248 (O_248,N_4954,N_4888);
and UO_249 (O_249,N_4970,N_4816);
nor UO_250 (O_250,N_4725,N_4218);
xor UO_251 (O_251,N_4629,N_4061);
nor UO_252 (O_252,N_4028,N_4771);
or UO_253 (O_253,N_4113,N_4484);
nand UO_254 (O_254,N_4545,N_4992);
nand UO_255 (O_255,N_4352,N_4433);
nor UO_256 (O_256,N_4152,N_4313);
nor UO_257 (O_257,N_4354,N_4149);
nand UO_258 (O_258,N_4290,N_4869);
nor UO_259 (O_259,N_4233,N_4299);
or UO_260 (O_260,N_4813,N_4746);
xor UO_261 (O_261,N_4635,N_4408);
and UO_262 (O_262,N_4264,N_4038);
nor UO_263 (O_263,N_4787,N_4025);
or UO_264 (O_264,N_4399,N_4336);
and UO_265 (O_265,N_4437,N_4798);
nand UO_266 (O_266,N_4250,N_4215);
nand UO_267 (O_267,N_4177,N_4517);
nor UO_268 (O_268,N_4249,N_4111);
nor UO_269 (O_269,N_4166,N_4405);
or UO_270 (O_270,N_4497,N_4778);
or UO_271 (O_271,N_4642,N_4128);
nand UO_272 (O_272,N_4698,N_4697);
and UO_273 (O_273,N_4064,N_4785);
or UO_274 (O_274,N_4422,N_4594);
or UO_275 (O_275,N_4424,N_4804);
and UO_276 (O_276,N_4756,N_4518);
nand UO_277 (O_277,N_4971,N_4974);
xnor UO_278 (O_278,N_4170,N_4526);
nand UO_279 (O_279,N_4474,N_4881);
or UO_280 (O_280,N_4095,N_4919);
nand UO_281 (O_281,N_4381,N_4160);
or UO_282 (O_282,N_4073,N_4482);
xor UO_283 (O_283,N_4118,N_4404);
or UO_284 (O_284,N_4430,N_4306);
nor UO_285 (O_285,N_4587,N_4035);
nor UO_286 (O_286,N_4245,N_4797);
and UO_287 (O_287,N_4986,N_4234);
nor UO_288 (O_288,N_4973,N_4260);
and UO_289 (O_289,N_4183,N_4510);
and UO_290 (O_290,N_4853,N_4267);
or UO_291 (O_291,N_4015,N_4280);
and UO_292 (O_292,N_4865,N_4570);
xor UO_293 (O_293,N_4039,N_4832);
xor UO_294 (O_294,N_4216,N_4837);
xnor UO_295 (O_295,N_4566,N_4933);
nor UO_296 (O_296,N_4929,N_4880);
or UO_297 (O_297,N_4975,N_4569);
and UO_298 (O_298,N_4619,N_4616);
and UO_299 (O_299,N_4106,N_4121);
nand UO_300 (O_300,N_4409,N_4425);
xnor UO_301 (O_301,N_4996,N_4358);
nand UO_302 (O_302,N_4942,N_4638);
or UO_303 (O_303,N_4591,N_4240);
or UO_304 (O_304,N_4675,N_4429);
or UO_305 (O_305,N_4155,N_4740);
and UO_306 (O_306,N_4086,N_4194);
or UO_307 (O_307,N_4512,N_4386);
nor UO_308 (O_308,N_4139,N_4450);
nor UO_309 (O_309,N_4972,N_4309);
or UO_310 (O_310,N_4401,N_4344);
nor UO_311 (O_311,N_4093,N_4196);
nand UO_312 (O_312,N_4302,N_4153);
and UO_313 (O_313,N_4831,N_4395);
nor UO_314 (O_314,N_4989,N_4943);
and UO_315 (O_315,N_4247,N_4646);
and UO_316 (O_316,N_4020,N_4056);
nand UO_317 (O_317,N_4998,N_4018);
or UO_318 (O_318,N_4601,N_4861);
nor UO_319 (O_319,N_4956,N_4351);
nand UO_320 (O_320,N_4696,N_4544);
or UO_321 (O_321,N_4988,N_4479);
or UO_322 (O_322,N_4863,N_4898);
and UO_323 (O_323,N_4192,N_4374);
nand UO_324 (O_324,N_4789,N_4909);
nor UO_325 (O_325,N_4953,N_4705);
nand UO_326 (O_326,N_4920,N_4684);
or UO_327 (O_327,N_4887,N_4945);
or UO_328 (O_328,N_4017,N_4071);
nor UO_329 (O_329,N_4758,N_4602);
nand UO_330 (O_330,N_4851,N_4946);
nor UO_331 (O_331,N_4846,N_4496);
or UO_332 (O_332,N_4214,N_4939);
xnor UO_333 (O_333,N_4076,N_4727);
nand UO_334 (O_334,N_4322,N_4206);
nand UO_335 (O_335,N_4557,N_4766);
and UO_336 (O_336,N_4780,N_4874);
and UO_337 (O_337,N_4169,N_4692);
or UO_338 (O_338,N_4010,N_4288);
and UO_339 (O_339,N_4396,N_4332);
or UO_340 (O_340,N_4801,N_4357);
or UO_341 (O_341,N_4561,N_4639);
or UO_342 (O_342,N_4701,N_4713);
nand UO_343 (O_343,N_4498,N_4220);
nor UO_344 (O_344,N_4680,N_4807);
xor UO_345 (O_345,N_4931,N_4271);
nand UO_346 (O_346,N_4244,N_4123);
and UO_347 (O_347,N_4411,N_4297);
nand UO_348 (O_348,N_4222,N_4895);
and UO_349 (O_349,N_4982,N_4156);
and UO_350 (O_350,N_4276,N_4519);
nand UO_351 (O_351,N_4554,N_4606);
or UO_352 (O_352,N_4913,N_4275);
or UO_353 (O_353,N_4328,N_4004);
xnor UO_354 (O_354,N_4984,N_4551);
nor UO_355 (O_355,N_4836,N_4350);
nand UO_356 (O_356,N_4467,N_4446);
nand UO_357 (O_357,N_4543,N_4266);
or UO_358 (O_358,N_4605,N_4707);
or UO_359 (O_359,N_4305,N_4665);
or UO_360 (O_360,N_4733,N_4608);
nand UO_361 (O_361,N_4023,N_4470);
nor UO_362 (O_362,N_4231,N_4239);
nor UO_363 (O_363,N_4765,N_4824);
and UO_364 (O_364,N_4653,N_4176);
and UO_365 (O_365,N_4834,N_4660);
nor UO_366 (O_366,N_4810,N_4722);
and UO_367 (O_367,N_4546,N_4341);
nor UO_368 (O_368,N_4500,N_4186);
xnor UO_369 (O_369,N_4375,N_4604);
nor UO_370 (O_370,N_4281,N_4256);
nand UO_371 (O_371,N_4054,N_4877);
and UO_372 (O_372,N_4356,N_4221);
xnor UO_373 (O_373,N_4978,N_4520);
nand UO_374 (O_374,N_4476,N_4795);
nand UO_375 (O_375,N_4188,N_4361);
and UO_376 (O_376,N_4294,N_4048);
and UO_377 (O_377,N_4582,N_4147);
and UO_378 (O_378,N_4884,N_4455);
nand UO_379 (O_379,N_4101,N_4891);
or UO_380 (O_380,N_4558,N_4755);
nor UO_381 (O_381,N_4620,N_4867);
or UO_382 (O_382,N_4588,N_4715);
or UO_383 (O_383,N_4068,N_4899);
nor UO_384 (O_384,N_4371,N_4914);
nor UO_385 (O_385,N_4723,N_4345);
or UO_386 (O_386,N_4983,N_4158);
and UO_387 (O_387,N_4489,N_4030);
nor UO_388 (O_388,N_4803,N_4142);
or UO_389 (O_389,N_4659,N_4444);
nor UO_390 (O_390,N_4506,N_4270);
xnor UO_391 (O_391,N_4126,N_4463);
xnor UO_392 (O_392,N_4246,N_4335);
xor UO_393 (O_393,N_4413,N_4547);
nor UO_394 (O_394,N_4823,N_4800);
or UO_395 (O_395,N_4213,N_4178);
nor UO_396 (O_396,N_4550,N_4952);
nor UO_397 (O_397,N_4235,N_4714);
nor UO_398 (O_398,N_4441,N_4752);
or UO_399 (O_399,N_4138,N_4274);
or UO_400 (O_400,N_4850,N_4481);
and UO_401 (O_401,N_4681,N_4228);
nor UO_402 (O_402,N_4699,N_4184);
or UO_403 (O_403,N_4067,N_4219);
nand UO_404 (O_404,N_4717,N_4210);
nand UO_405 (O_405,N_4849,N_4611);
and UO_406 (O_406,N_4457,N_4958);
nor UO_407 (O_407,N_4343,N_4907);
and UO_408 (O_408,N_4383,N_4050);
nor UO_409 (O_409,N_4145,N_4835);
and UO_410 (O_410,N_4886,N_4617);
or UO_411 (O_411,N_4674,N_4293);
nand UO_412 (O_412,N_4403,N_4427);
nor UO_413 (O_413,N_4203,N_4876);
nor UO_414 (O_414,N_4932,N_4133);
xnor UO_415 (O_415,N_4710,N_4577);
xor UO_416 (O_416,N_4736,N_4261);
nor UO_417 (O_417,N_4053,N_4757);
nor UO_418 (O_418,N_4006,N_4894);
nor UO_419 (O_419,N_4576,N_4248);
or UO_420 (O_420,N_4685,N_4969);
and UO_421 (O_421,N_4689,N_4995);
or UO_422 (O_422,N_4927,N_4760);
or UO_423 (O_423,N_4967,N_4180);
or UO_424 (O_424,N_4936,N_4735);
and UO_425 (O_425,N_4515,N_4840);
or UO_426 (O_426,N_4505,N_4307);
and UO_427 (O_427,N_4985,N_4384);
nand UO_428 (O_428,N_4308,N_4770);
nand UO_429 (O_429,N_4279,N_4871);
nor UO_430 (O_430,N_4310,N_4421);
nand UO_431 (O_431,N_4965,N_4189);
nor UO_432 (O_432,N_4419,N_4277);
and UO_433 (O_433,N_4612,N_4088);
and UO_434 (O_434,N_4102,N_4157);
nor UO_435 (O_435,N_4501,N_4312);
and UO_436 (O_436,N_4168,N_4767);
xor UO_437 (O_437,N_4397,N_4418);
or UO_438 (O_438,N_4814,N_4159);
nand UO_439 (O_439,N_4724,N_4651);
nor UO_440 (O_440,N_4200,N_4670);
and UO_441 (O_441,N_4001,N_4057);
nand UO_442 (O_442,N_4900,N_4782);
and UO_443 (O_443,N_4303,N_4957);
nor UO_444 (O_444,N_4610,N_4380);
nor UO_445 (O_445,N_4175,N_4892);
and UO_446 (O_446,N_4704,N_4525);
or UO_447 (O_447,N_4799,N_4443);
or UO_448 (O_448,N_4626,N_4253);
xnor UO_449 (O_449,N_4676,N_4508);
xor UO_450 (O_450,N_4019,N_4664);
or UO_451 (O_451,N_4822,N_4466);
or UO_452 (O_452,N_4137,N_4866);
or UO_453 (O_453,N_4790,N_4592);
nor UO_454 (O_454,N_4171,N_4784);
nand UO_455 (O_455,N_4948,N_4150);
or UO_456 (O_456,N_4263,N_4542);
nor UO_457 (O_457,N_4385,N_4977);
and UO_458 (O_458,N_4052,N_4792);
nand UO_459 (O_459,N_4882,N_4734);
or UO_460 (O_460,N_4182,N_4854);
nor UO_461 (O_461,N_4072,N_4033);
or UO_462 (O_462,N_4316,N_4565);
xor UO_463 (O_463,N_4786,N_4859);
and UO_464 (O_464,N_4897,N_4855);
nand UO_465 (O_465,N_4478,N_4340);
and UO_466 (O_466,N_4774,N_4560);
or UO_467 (O_467,N_4993,N_4058);
and UO_468 (O_468,N_4902,N_4097);
nand UO_469 (O_469,N_4603,N_4092);
and UO_470 (O_470,N_4414,N_4103);
nor UO_471 (O_471,N_4662,N_4367);
or UO_472 (O_472,N_4683,N_4392);
or UO_473 (O_473,N_4460,N_4041);
and UO_474 (O_474,N_4572,N_4252);
nor UO_475 (O_475,N_4843,N_4503);
nand UO_476 (O_476,N_4730,N_4645);
or UO_477 (O_477,N_4937,N_4464);
and UO_478 (O_478,N_4596,N_4507);
nor UO_479 (O_479,N_4485,N_4938);
nor UO_480 (O_480,N_4583,N_4195);
and UO_481 (O_481,N_4461,N_4555);
nand UO_482 (O_482,N_4099,N_4144);
xnor UO_483 (O_483,N_4377,N_4628);
and UO_484 (O_484,N_4473,N_4278);
nor UO_485 (O_485,N_4331,N_4870);
nor UO_486 (O_486,N_4564,N_4207);
nand UO_487 (O_487,N_4595,N_4647);
and UO_488 (O_488,N_4296,N_4941);
nor UO_489 (O_489,N_4918,N_4449);
nand UO_490 (O_490,N_4718,N_4442);
nand UO_491 (O_491,N_4669,N_4745);
and UO_492 (O_492,N_4314,N_4062);
nor UO_493 (O_493,N_4524,N_4407);
and UO_494 (O_494,N_4338,N_4960);
and UO_495 (O_495,N_4521,N_4387);
xnor UO_496 (O_496,N_4634,N_4940);
or UO_497 (O_497,N_4636,N_4330);
nor UO_498 (O_498,N_4915,N_4319);
and UO_499 (O_499,N_4090,N_4254);
and UO_500 (O_500,N_4649,N_4884);
or UO_501 (O_501,N_4268,N_4398);
and UO_502 (O_502,N_4391,N_4078);
or UO_503 (O_503,N_4989,N_4325);
nand UO_504 (O_504,N_4484,N_4516);
nor UO_505 (O_505,N_4950,N_4644);
nand UO_506 (O_506,N_4519,N_4857);
nand UO_507 (O_507,N_4833,N_4054);
nand UO_508 (O_508,N_4399,N_4104);
nand UO_509 (O_509,N_4297,N_4831);
nor UO_510 (O_510,N_4467,N_4196);
nand UO_511 (O_511,N_4620,N_4274);
and UO_512 (O_512,N_4469,N_4063);
or UO_513 (O_513,N_4108,N_4243);
nand UO_514 (O_514,N_4099,N_4688);
nand UO_515 (O_515,N_4796,N_4383);
nand UO_516 (O_516,N_4216,N_4905);
xor UO_517 (O_517,N_4103,N_4088);
and UO_518 (O_518,N_4239,N_4706);
or UO_519 (O_519,N_4820,N_4954);
and UO_520 (O_520,N_4845,N_4510);
or UO_521 (O_521,N_4520,N_4944);
or UO_522 (O_522,N_4828,N_4890);
nand UO_523 (O_523,N_4453,N_4802);
xnor UO_524 (O_524,N_4388,N_4852);
or UO_525 (O_525,N_4411,N_4130);
nor UO_526 (O_526,N_4992,N_4575);
and UO_527 (O_527,N_4733,N_4453);
nor UO_528 (O_528,N_4439,N_4032);
nor UO_529 (O_529,N_4167,N_4352);
and UO_530 (O_530,N_4289,N_4057);
or UO_531 (O_531,N_4388,N_4171);
or UO_532 (O_532,N_4154,N_4011);
nor UO_533 (O_533,N_4503,N_4257);
xnor UO_534 (O_534,N_4375,N_4971);
nor UO_535 (O_535,N_4691,N_4334);
nand UO_536 (O_536,N_4912,N_4433);
nand UO_537 (O_537,N_4436,N_4026);
or UO_538 (O_538,N_4789,N_4300);
nand UO_539 (O_539,N_4198,N_4135);
or UO_540 (O_540,N_4084,N_4609);
nand UO_541 (O_541,N_4899,N_4948);
nor UO_542 (O_542,N_4974,N_4420);
and UO_543 (O_543,N_4473,N_4350);
nand UO_544 (O_544,N_4208,N_4299);
and UO_545 (O_545,N_4745,N_4680);
nand UO_546 (O_546,N_4554,N_4281);
and UO_547 (O_547,N_4029,N_4009);
or UO_548 (O_548,N_4016,N_4604);
or UO_549 (O_549,N_4935,N_4744);
and UO_550 (O_550,N_4485,N_4673);
and UO_551 (O_551,N_4411,N_4889);
and UO_552 (O_552,N_4626,N_4406);
and UO_553 (O_553,N_4835,N_4538);
and UO_554 (O_554,N_4038,N_4945);
or UO_555 (O_555,N_4407,N_4180);
or UO_556 (O_556,N_4471,N_4847);
xnor UO_557 (O_557,N_4213,N_4171);
xor UO_558 (O_558,N_4810,N_4485);
and UO_559 (O_559,N_4607,N_4182);
nor UO_560 (O_560,N_4098,N_4498);
nand UO_561 (O_561,N_4960,N_4345);
nor UO_562 (O_562,N_4707,N_4402);
nand UO_563 (O_563,N_4659,N_4883);
xnor UO_564 (O_564,N_4391,N_4608);
and UO_565 (O_565,N_4304,N_4154);
nor UO_566 (O_566,N_4469,N_4869);
or UO_567 (O_567,N_4382,N_4791);
nand UO_568 (O_568,N_4636,N_4633);
and UO_569 (O_569,N_4057,N_4820);
nand UO_570 (O_570,N_4644,N_4565);
nand UO_571 (O_571,N_4054,N_4019);
or UO_572 (O_572,N_4806,N_4817);
nor UO_573 (O_573,N_4760,N_4555);
nor UO_574 (O_574,N_4334,N_4432);
xnor UO_575 (O_575,N_4124,N_4369);
or UO_576 (O_576,N_4673,N_4205);
nand UO_577 (O_577,N_4134,N_4199);
or UO_578 (O_578,N_4934,N_4883);
nand UO_579 (O_579,N_4571,N_4223);
or UO_580 (O_580,N_4025,N_4299);
nand UO_581 (O_581,N_4189,N_4741);
nor UO_582 (O_582,N_4501,N_4788);
nand UO_583 (O_583,N_4466,N_4874);
nor UO_584 (O_584,N_4556,N_4254);
nor UO_585 (O_585,N_4709,N_4103);
and UO_586 (O_586,N_4091,N_4418);
or UO_587 (O_587,N_4140,N_4508);
or UO_588 (O_588,N_4217,N_4559);
or UO_589 (O_589,N_4206,N_4859);
nand UO_590 (O_590,N_4047,N_4994);
nand UO_591 (O_591,N_4551,N_4814);
or UO_592 (O_592,N_4088,N_4648);
and UO_593 (O_593,N_4197,N_4684);
nor UO_594 (O_594,N_4527,N_4577);
and UO_595 (O_595,N_4283,N_4160);
or UO_596 (O_596,N_4941,N_4822);
nor UO_597 (O_597,N_4759,N_4827);
and UO_598 (O_598,N_4808,N_4847);
xor UO_599 (O_599,N_4290,N_4196);
nand UO_600 (O_600,N_4708,N_4696);
nand UO_601 (O_601,N_4731,N_4200);
and UO_602 (O_602,N_4519,N_4566);
nor UO_603 (O_603,N_4482,N_4636);
nor UO_604 (O_604,N_4880,N_4636);
xor UO_605 (O_605,N_4207,N_4781);
nand UO_606 (O_606,N_4924,N_4820);
nor UO_607 (O_607,N_4772,N_4473);
and UO_608 (O_608,N_4683,N_4207);
or UO_609 (O_609,N_4199,N_4742);
nor UO_610 (O_610,N_4159,N_4754);
nand UO_611 (O_611,N_4564,N_4342);
and UO_612 (O_612,N_4190,N_4474);
or UO_613 (O_613,N_4982,N_4821);
or UO_614 (O_614,N_4611,N_4205);
and UO_615 (O_615,N_4044,N_4459);
nor UO_616 (O_616,N_4750,N_4087);
and UO_617 (O_617,N_4099,N_4766);
nor UO_618 (O_618,N_4005,N_4152);
and UO_619 (O_619,N_4971,N_4639);
nand UO_620 (O_620,N_4847,N_4604);
and UO_621 (O_621,N_4584,N_4327);
nor UO_622 (O_622,N_4874,N_4687);
nand UO_623 (O_623,N_4610,N_4148);
or UO_624 (O_624,N_4116,N_4313);
or UO_625 (O_625,N_4893,N_4635);
nand UO_626 (O_626,N_4127,N_4501);
and UO_627 (O_627,N_4917,N_4329);
nand UO_628 (O_628,N_4554,N_4433);
or UO_629 (O_629,N_4873,N_4550);
and UO_630 (O_630,N_4828,N_4774);
nor UO_631 (O_631,N_4867,N_4141);
nand UO_632 (O_632,N_4928,N_4481);
or UO_633 (O_633,N_4229,N_4178);
nor UO_634 (O_634,N_4792,N_4394);
nand UO_635 (O_635,N_4540,N_4254);
nand UO_636 (O_636,N_4472,N_4626);
nor UO_637 (O_637,N_4783,N_4409);
nor UO_638 (O_638,N_4933,N_4114);
or UO_639 (O_639,N_4571,N_4965);
and UO_640 (O_640,N_4798,N_4576);
xnor UO_641 (O_641,N_4842,N_4845);
nand UO_642 (O_642,N_4468,N_4449);
xor UO_643 (O_643,N_4577,N_4621);
nor UO_644 (O_644,N_4763,N_4673);
nor UO_645 (O_645,N_4613,N_4374);
nand UO_646 (O_646,N_4778,N_4139);
or UO_647 (O_647,N_4046,N_4736);
and UO_648 (O_648,N_4409,N_4308);
or UO_649 (O_649,N_4207,N_4188);
and UO_650 (O_650,N_4060,N_4985);
and UO_651 (O_651,N_4802,N_4046);
and UO_652 (O_652,N_4304,N_4632);
nand UO_653 (O_653,N_4480,N_4910);
nand UO_654 (O_654,N_4281,N_4542);
nand UO_655 (O_655,N_4269,N_4068);
nand UO_656 (O_656,N_4309,N_4408);
or UO_657 (O_657,N_4526,N_4441);
xor UO_658 (O_658,N_4971,N_4550);
and UO_659 (O_659,N_4284,N_4680);
nor UO_660 (O_660,N_4710,N_4647);
or UO_661 (O_661,N_4668,N_4078);
and UO_662 (O_662,N_4797,N_4863);
and UO_663 (O_663,N_4208,N_4423);
xnor UO_664 (O_664,N_4778,N_4107);
nand UO_665 (O_665,N_4423,N_4440);
nand UO_666 (O_666,N_4669,N_4044);
nand UO_667 (O_667,N_4661,N_4619);
or UO_668 (O_668,N_4604,N_4209);
or UO_669 (O_669,N_4263,N_4254);
xnor UO_670 (O_670,N_4541,N_4635);
nand UO_671 (O_671,N_4545,N_4507);
and UO_672 (O_672,N_4877,N_4141);
nor UO_673 (O_673,N_4910,N_4881);
nor UO_674 (O_674,N_4877,N_4852);
and UO_675 (O_675,N_4511,N_4502);
nand UO_676 (O_676,N_4087,N_4152);
or UO_677 (O_677,N_4919,N_4554);
or UO_678 (O_678,N_4191,N_4814);
or UO_679 (O_679,N_4579,N_4213);
or UO_680 (O_680,N_4246,N_4844);
or UO_681 (O_681,N_4415,N_4205);
and UO_682 (O_682,N_4608,N_4819);
and UO_683 (O_683,N_4595,N_4747);
xor UO_684 (O_684,N_4726,N_4051);
nand UO_685 (O_685,N_4990,N_4558);
and UO_686 (O_686,N_4413,N_4434);
and UO_687 (O_687,N_4545,N_4156);
nor UO_688 (O_688,N_4948,N_4666);
and UO_689 (O_689,N_4049,N_4513);
xor UO_690 (O_690,N_4163,N_4515);
or UO_691 (O_691,N_4305,N_4050);
and UO_692 (O_692,N_4217,N_4715);
nand UO_693 (O_693,N_4569,N_4931);
and UO_694 (O_694,N_4823,N_4845);
or UO_695 (O_695,N_4628,N_4819);
and UO_696 (O_696,N_4786,N_4422);
and UO_697 (O_697,N_4449,N_4893);
xor UO_698 (O_698,N_4805,N_4199);
xnor UO_699 (O_699,N_4308,N_4080);
nor UO_700 (O_700,N_4887,N_4188);
nand UO_701 (O_701,N_4913,N_4395);
or UO_702 (O_702,N_4679,N_4939);
and UO_703 (O_703,N_4941,N_4792);
nand UO_704 (O_704,N_4476,N_4044);
nor UO_705 (O_705,N_4970,N_4431);
nor UO_706 (O_706,N_4279,N_4230);
xnor UO_707 (O_707,N_4205,N_4023);
and UO_708 (O_708,N_4823,N_4428);
nor UO_709 (O_709,N_4316,N_4952);
nor UO_710 (O_710,N_4625,N_4387);
nor UO_711 (O_711,N_4916,N_4145);
nand UO_712 (O_712,N_4613,N_4088);
and UO_713 (O_713,N_4676,N_4382);
nand UO_714 (O_714,N_4123,N_4833);
and UO_715 (O_715,N_4351,N_4558);
nand UO_716 (O_716,N_4765,N_4344);
nand UO_717 (O_717,N_4434,N_4981);
nand UO_718 (O_718,N_4813,N_4732);
and UO_719 (O_719,N_4526,N_4542);
nor UO_720 (O_720,N_4365,N_4545);
and UO_721 (O_721,N_4503,N_4612);
nand UO_722 (O_722,N_4313,N_4163);
and UO_723 (O_723,N_4126,N_4490);
nor UO_724 (O_724,N_4970,N_4080);
or UO_725 (O_725,N_4592,N_4533);
nor UO_726 (O_726,N_4787,N_4430);
nor UO_727 (O_727,N_4578,N_4892);
or UO_728 (O_728,N_4625,N_4536);
and UO_729 (O_729,N_4593,N_4894);
nor UO_730 (O_730,N_4150,N_4857);
nor UO_731 (O_731,N_4685,N_4799);
and UO_732 (O_732,N_4570,N_4141);
nand UO_733 (O_733,N_4928,N_4366);
nor UO_734 (O_734,N_4582,N_4492);
nand UO_735 (O_735,N_4447,N_4935);
nand UO_736 (O_736,N_4439,N_4207);
nand UO_737 (O_737,N_4799,N_4300);
nor UO_738 (O_738,N_4019,N_4247);
nor UO_739 (O_739,N_4319,N_4185);
nor UO_740 (O_740,N_4666,N_4461);
or UO_741 (O_741,N_4275,N_4409);
xnor UO_742 (O_742,N_4639,N_4754);
xor UO_743 (O_743,N_4277,N_4003);
nor UO_744 (O_744,N_4583,N_4135);
nand UO_745 (O_745,N_4877,N_4327);
nor UO_746 (O_746,N_4955,N_4693);
xnor UO_747 (O_747,N_4758,N_4206);
and UO_748 (O_748,N_4763,N_4899);
nor UO_749 (O_749,N_4925,N_4887);
or UO_750 (O_750,N_4636,N_4515);
xnor UO_751 (O_751,N_4545,N_4048);
and UO_752 (O_752,N_4961,N_4933);
or UO_753 (O_753,N_4967,N_4578);
and UO_754 (O_754,N_4175,N_4447);
or UO_755 (O_755,N_4248,N_4763);
nor UO_756 (O_756,N_4907,N_4174);
or UO_757 (O_757,N_4903,N_4308);
nor UO_758 (O_758,N_4524,N_4301);
nand UO_759 (O_759,N_4960,N_4257);
nor UO_760 (O_760,N_4385,N_4423);
xor UO_761 (O_761,N_4559,N_4448);
nor UO_762 (O_762,N_4626,N_4751);
or UO_763 (O_763,N_4964,N_4008);
and UO_764 (O_764,N_4601,N_4925);
nor UO_765 (O_765,N_4860,N_4100);
nor UO_766 (O_766,N_4521,N_4096);
nand UO_767 (O_767,N_4909,N_4058);
and UO_768 (O_768,N_4723,N_4437);
or UO_769 (O_769,N_4695,N_4769);
or UO_770 (O_770,N_4580,N_4701);
nor UO_771 (O_771,N_4307,N_4237);
nor UO_772 (O_772,N_4018,N_4327);
nor UO_773 (O_773,N_4624,N_4067);
or UO_774 (O_774,N_4176,N_4404);
nor UO_775 (O_775,N_4761,N_4822);
nor UO_776 (O_776,N_4360,N_4546);
and UO_777 (O_777,N_4258,N_4416);
nor UO_778 (O_778,N_4458,N_4993);
or UO_779 (O_779,N_4726,N_4116);
nor UO_780 (O_780,N_4018,N_4069);
xnor UO_781 (O_781,N_4325,N_4448);
nor UO_782 (O_782,N_4297,N_4001);
and UO_783 (O_783,N_4533,N_4899);
or UO_784 (O_784,N_4364,N_4219);
or UO_785 (O_785,N_4164,N_4411);
nor UO_786 (O_786,N_4665,N_4974);
nor UO_787 (O_787,N_4580,N_4266);
xor UO_788 (O_788,N_4434,N_4520);
nor UO_789 (O_789,N_4347,N_4637);
or UO_790 (O_790,N_4451,N_4575);
or UO_791 (O_791,N_4580,N_4325);
xnor UO_792 (O_792,N_4825,N_4858);
or UO_793 (O_793,N_4361,N_4061);
nand UO_794 (O_794,N_4037,N_4214);
nand UO_795 (O_795,N_4621,N_4273);
nor UO_796 (O_796,N_4589,N_4722);
or UO_797 (O_797,N_4257,N_4545);
nor UO_798 (O_798,N_4404,N_4659);
and UO_799 (O_799,N_4769,N_4005);
or UO_800 (O_800,N_4535,N_4218);
nand UO_801 (O_801,N_4740,N_4121);
nand UO_802 (O_802,N_4509,N_4202);
nor UO_803 (O_803,N_4090,N_4188);
nor UO_804 (O_804,N_4039,N_4338);
nor UO_805 (O_805,N_4339,N_4529);
nor UO_806 (O_806,N_4711,N_4169);
nor UO_807 (O_807,N_4883,N_4168);
nand UO_808 (O_808,N_4483,N_4115);
nor UO_809 (O_809,N_4463,N_4150);
and UO_810 (O_810,N_4931,N_4444);
nand UO_811 (O_811,N_4489,N_4549);
nor UO_812 (O_812,N_4672,N_4668);
nand UO_813 (O_813,N_4135,N_4294);
and UO_814 (O_814,N_4750,N_4268);
xnor UO_815 (O_815,N_4914,N_4975);
xor UO_816 (O_816,N_4435,N_4245);
and UO_817 (O_817,N_4352,N_4833);
nor UO_818 (O_818,N_4907,N_4578);
nor UO_819 (O_819,N_4669,N_4706);
nor UO_820 (O_820,N_4450,N_4941);
nor UO_821 (O_821,N_4881,N_4583);
nand UO_822 (O_822,N_4105,N_4255);
or UO_823 (O_823,N_4639,N_4428);
or UO_824 (O_824,N_4337,N_4117);
and UO_825 (O_825,N_4655,N_4526);
or UO_826 (O_826,N_4264,N_4115);
nor UO_827 (O_827,N_4145,N_4617);
xor UO_828 (O_828,N_4102,N_4768);
nand UO_829 (O_829,N_4363,N_4111);
or UO_830 (O_830,N_4716,N_4469);
nand UO_831 (O_831,N_4542,N_4552);
or UO_832 (O_832,N_4237,N_4094);
nor UO_833 (O_833,N_4364,N_4540);
nand UO_834 (O_834,N_4599,N_4783);
nor UO_835 (O_835,N_4474,N_4166);
or UO_836 (O_836,N_4605,N_4143);
nor UO_837 (O_837,N_4913,N_4379);
xor UO_838 (O_838,N_4822,N_4123);
or UO_839 (O_839,N_4124,N_4292);
and UO_840 (O_840,N_4747,N_4505);
xnor UO_841 (O_841,N_4397,N_4073);
nand UO_842 (O_842,N_4032,N_4860);
or UO_843 (O_843,N_4938,N_4839);
and UO_844 (O_844,N_4511,N_4160);
xor UO_845 (O_845,N_4945,N_4913);
or UO_846 (O_846,N_4307,N_4066);
nand UO_847 (O_847,N_4580,N_4529);
and UO_848 (O_848,N_4311,N_4934);
nand UO_849 (O_849,N_4894,N_4378);
nor UO_850 (O_850,N_4050,N_4873);
or UO_851 (O_851,N_4331,N_4818);
nor UO_852 (O_852,N_4397,N_4055);
and UO_853 (O_853,N_4363,N_4467);
and UO_854 (O_854,N_4855,N_4509);
and UO_855 (O_855,N_4412,N_4541);
nand UO_856 (O_856,N_4064,N_4040);
and UO_857 (O_857,N_4789,N_4795);
or UO_858 (O_858,N_4393,N_4241);
nor UO_859 (O_859,N_4793,N_4658);
or UO_860 (O_860,N_4159,N_4150);
or UO_861 (O_861,N_4345,N_4187);
and UO_862 (O_862,N_4736,N_4118);
nand UO_863 (O_863,N_4329,N_4533);
or UO_864 (O_864,N_4146,N_4453);
nor UO_865 (O_865,N_4859,N_4617);
nand UO_866 (O_866,N_4395,N_4861);
nand UO_867 (O_867,N_4299,N_4017);
nand UO_868 (O_868,N_4806,N_4915);
and UO_869 (O_869,N_4697,N_4042);
xnor UO_870 (O_870,N_4186,N_4528);
and UO_871 (O_871,N_4553,N_4597);
nand UO_872 (O_872,N_4424,N_4637);
and UO_873 (O_873,N_4486,N_4975);
nand UO_874 (O_874,N_4787,N_4819);
or UO_875 (O_875,N_4710,N_4139);
xor UO_876 (O_876,N_4133,N_4876);
or UO_877 (O_877,N_4767,N_4303);
nor UO_878 (O_878,N_4380,N_4709);
nand UO_879 (O_879,N_4954,N_4330);
nand UO_880 (O_880,N_4914,N_4799);
or UO_881 (O_881,N_4574,N_4268);
or UO_882 (O_882,N_4853,N_4579);
and UO_883 (O_883,N_4802,N_4184);
nor UO_884 (O_884,N_4361,N_4857);
nor UO_885 (O_885,N_4192,N_4235);
nor UO_886 (O_886,N_4460,N_4712);
nand UO_887 (O_887,N_4199,N_4557);
nand UO_888 (O_888,N_4759,N_4256);
nor UO_889 (O_889,N_4251,N_4421);
nand UO_890 (O_890,N_4137,N_4168);
and UO_891 (O_891,N_4929,N_4256);
nor UO_892 (O_892,N_4581,N_4266);
nor UO_893 (O_893,N_4789,N_4035);
nor UO_894 (O_894,N_4162,N_4362);
xnor UO_895 (O_895,N_4012,N_4712);
or UO_896 (O_896,N_4413,N_4623);
nor UO_897 (O_897,N_4767,N_4713);
and UO_898 (O_898,N_4876,N_4139);
nor UO_899 (O_899,N_4156,N_4321);
nand UO_900 (O_900,N_4063,N_4204);
and UO_901 (O_901,N_4246,N_4784);
and UO_902 (O_902,N_4586,N_4750);
and UO_903 (O_903,N_4187,N_4173);
nor UO_904 (O_904,N_4230,N_4053);
nor UO_905 (O_905,N_4302,N_4397);
and UO_906 (O_906,N_4011,N_4897);
nor UO_907 (O_907,N_4806,N_4088);
and UO_908 (O_908,N_4960,N_4673);
nand UO_909 (O_909,N_4606,N_4400);
and UO_910 (O_910,N_4876,N_4734);
nor UO_911 (O_911,N_4959,N_4940);
xnor UO_912 (O_912,N_4046,N_4990);
and UO_913 (O_913,N_4675,N_4717);
and UO_914 (O_914,N_4564,N_4400);
and UO_915 (O_915,N_4191,N_4370);
or UO_916 (O_916,N_4423,N_4222);
or UO_917 (O_917,N_4979,N_4625);
nand UO_918 (O_918,N_4931,N_4454);
and UO_919 (O_919,N_4314,N_4986);
or UO_920 (O_920,N_4759,N_4230);
nand UO_921 (O_921,N_4571,N_4698);
nand UO_922 (O_922,N_4179,N_4762);
and UO_923 (O_923,N_4394,N_4757);
xnor UO_924 (O_924,N_4918,N_4223);
and UO_925 (O_925,N_4897,N_4972);
nor UO_926 (O_926,N_4075,N_4220);
nand UO_927 (O_927,N_4928,N_4397);
nor UO_928 (O_928,N_4356,N_4838);
nor UO_929 (O_929,N_4448,N_4474);
and UO_930 (O_930,N_4499,N_4288);
nor UO_931 (O_931,N_4431,N_4305);
nand UO_932 (O_932,N_4628,N_4765);
or UO_933 (O_933,N_4919,N_4096);
nand UO_934 (O_934,N_4700,N_4473);
and UO_935 (O_935,N_4702,N_4510);
or UO_936 (O_936,N_4766,N_4511);
nor UO_937 (O_937,N_4241,N_4892);
xnor UO_938 (O_938,N_4173,N_4009);
nor UO_939 (O_939,N_4827,N_4347);
and UO_940 (O_940,N_4748,N_4621);
nand UO_941 (O_941,N_4568,N_4551);
nor UO_942 (O_942,N_4409,N_4834);
xor UO_943 (O_943,N_4842,N_4600);
or UO_944 (O_944,N_4534,N_4837);
or UO_945 (O_945,N_4897,N_4375);
nor UO_946 (O_946,N_4467,N_4739);
nand UO_947 (O_947,N_4176,N_4088);
or UO_948 (O_948,N_4443,N_4990);
nor UO_949 (O_949,N_4099,N_4328);
and UO_950 (O_950,N_4598,N_4965);
nand UO_951 (O_951,N_4865,N_4027);
nor UO_952 (O_952,N_4493,N_4166);
and UO_953 (O_953,N_4277,N_4616);
xor UO_954 (O_954,N_4041,N_4715);
or UO_955 (O_955,N_4315,N_4595);
xnor UO_956 (O_956,N_4204,N_4574);
and UO_957 (O_957,N_4598,N_4368);
nand UO_958 (O_958,N_4622,N_4178);
or UO_959 (O_959,N_4566,N_4448);
nand UO_960 (O_960,N_4801,N_4334);
nand UO_961 (O_961,N_4369,N_4018);
or UO_962 (O_962,N_4709,N_4222);
and UO_963 (O_963,N_4703,N_4044);
or UO_964 (O_964,N_4690,N_4264);
or UO_965 (O_965,N_4319,N_4853);
or UO_966 (O_966,N_4775,N_4967);
or UO_967 (O_967,N_4410,N_4521);
nand UO_968 (O_968,N_4587,N_4343);
nand UO_969 (O_969,N_4876,N_4616);
nor UO_970 (O_970,N_4170,N_4166);
nor UO_971 (O_971,N_4138,N_4162);
nand UO_972 (O_972,N_4756,N_4654);
and UO_973 (O_973,N_4475,N_4923);
nor UO_974 (O_974,N_4830,N_4691);
nand UO_975 (O_975,N_4401,N_4584);
or UO_976 (O_976,N_4670,N_4649);
nand UO_977 (O_977,N_4165,N_4704);
nor UO_978 (O_978,N_4287,N_4979);
and UO_979 (O_979,N_4413,N_4349);
nor UO_980 (O_980,N_4783,N_4873);
nor UO_981 (O_981,N_4914,N_4380);
nor UO_982 (O_982,N_4017,N_4796);
nand UO_983 (O_983,N_4797,N_4109);
nor UO_984 (O_984,N_4454,N_4016);
and UO_985 (O_985,N_4162,N_4675);
nor UO_986 (O_986,N_4651,N_4828);
nand UO_987 (O_987,N_4071,N_4937);
nand UO_988 (O_988,N_4395,N_4709);
nor UO_989 (O_989,N_4326,N_4938);
nor UO_990 (O_990,N_4141,N_4636);
and UO_991 (O_991,N_4984,N_4331);
nand UO_992 (O_992,N_4127,N_4172);
and UO_993 (O_993,N_4650,N_4914);
xnor UO_994 (O_994,N_4209,N_4813);
or UO_995 (O_995,N_4882,N_4456);
and UO_996 (O_996,N_4196,N_4079);
and UO_997 (O_997,N_4386,N_4154);
xor UO_998 (O_998,N_4086,N_4119);
or UO_999 (O_999,N_4369,N_4546);
endmodule