module basic_2000_20000_2500_10_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1695,In_834);
or U1 (N_1,In_610,In_970);
or U2 (N_2,In_1018,In_370);
nor U3 (N_3,In_1882,In_1232);
xor U4 (N_4,In_1535,In_318);
or U5 (N_5,In_206,In_1488);
and U6 (N_6,In_708,In_347);
and U7 (N_7,In_321,In_338);
nand U8 (N_8,In_1682,In_634);
nand U9 (N_9,In_1323,In_1979);
or U10 (N_10,In_1898,In_1280);
nor U11 (N_11,In_1799,In_1177);
nor U12 (N_12,In_1199,In_1723);
nand U13 (N_13,In_393,In_1539);
nand U14 (N_14,In_1374,In_574);
nor U15 (N_15,In_343,In_312);
or U16 (N_16,In_1759,In_1709);
nor U17 (N_17,In_995,In_1163);
or U18 (N_18,In_1890,In_1640);
and U19 (N_19,In_55,In_128);
nand U20 (N_20,In_1333,In_1254);
and U21 (N_21,In_407,In_739);
or U22 (N_22,In_894,In_1997);
nand U23 (N_23,In_1827,In_322);
and U24 (N_24,In_1495,In_53);
nor U25 (N_25,In_123,In_924);
xnor U26 (N_26,In_399,In_444);
nand U27 (N_27,In_942,In_199);
or U28 (N_28,In_1390,In_358);
nor U29 (N_29,In_909,In_1393);
nor U30 (N_30,In_1010,In_458);
xor U31 (N_31,In_583,In_654);
or U32 (N_32,In_1097,In_177);
nor U33 (N_33,In_682,In_1472);
and U34 (N_34,In_964,In_1897);
and U35 (N_35,In_716,In_1895);
or U36 (N_36,In_895,In_556);
nand U37 (N_37,In_1060,In_74);
xor U38 (N_38,In_421,In_1514);
nand U39 (N_39,In_1080,In_1491);
or U40 (N_40,In_723,In_1557);
or U41 (N_41,In_1204,In_33);
and U42 (N_42,In_819,In_516);
and U43 (N_43,In_744,In_1612);
xor U44 (N_44,In_481,In_1774);
and U45 (N_45,In_1515,In_1518);
and U46 (N_46,In_1486,In_267);
and U47 (N_47,In_1257,In_1470);
or U48 (N_48,In_455,In_673);
nor U49 (N_49,In_196,In_1490);
and U50 (N_50,In_911,In_1685);
nand U51 (N_51,In_777,In_807);
xor U52 (N_52,In_1580,In_527);
nor U53 (N_53,In_701,In_1626);
and U54 (N_54,In_724,In_1193);
or U55 (N_55,In_1386,In_1952);
xor U56 (N_56,In_1639,In_1595);
nand U57 (N_57,In_1290,In_1750);
and U58 (N_58,In_1127,In_468);
or U59 (N_59,In_19,In_1594);
nor U60 (N_60,In_400,In_905);
nand U61 (N_61,In_222,In_1752);
nand U62 (N_62,In_820,In_1237);
nand U63 (N_63,In_586,In_502);
and U64 (N_64,In_687,In_1591);
nor U65 (N_65,In_757,In_355);
nand U66 (N_66,In_404,In_725);
or U67 (N_67,In_329,In_1305);
nand U68 (N_68,In_1468,In_1522);
and U69 (N_69,In_917,In_1065);
nor U70 (N_70,In_1854,In_1441);
or U71 (N_71,In_1085,In_1231);
and U72 (N_72,In_867,In_1094);
or U73 (N_73,In_122,In_1943);
and U74 (N_74,In_1637,In_1106);
or U75 (N_75,In_1415,In_562);
and U76 (N_76,In_1316,In_1928);
and U77 (N_77,In_389,In_1630);
and U78 (N_78,In_180,In_939);
nand U79 (N_79,In_97,In_838);
nor U80 (N_80,In_1966,In_1235);
nor U81 (N_81,In_362,In_1540);
nor U82 (N_82,In_1781,In_402);
and U83 (N_83,In_1961,In_1315);
or U84 (N_84,In_1383,In_361);
and U85 (N_85,In_498,In_1);
or U86 (N_86,In_1924,In_156);
or U87 (N_87,In_1593,In_472);
xnor U88 (N_88,In_1796,In_1657);
nand U89 (N_89,In_657,In_398);
or U90 (N_90,In_1615,In_885);
nand U91 (N_91,In_533,In_800);
nand U92 (N_92,In_1355,In_1766);
nor U93 (N_93,In_636,In_1465);
nand U94 (N_94,In_1104,In_1680);
nand U95 (N_95,In_1800,In_1443);
nor U96 (N_96,In_875,In_1746);
nor U97 (N_97,In_469,In_1099);
and U98 (N_98,In_855,In_396);
nor U99 (N_99,In_44,In_1608);
nand U100 (N_100,In_990,In_535);
nor U101 (N_101,In_1824,In_1831);
and U102 (N_102,In_549,In_390);
and U103 (N_103,In_1963,In_114);
nor U104 (N_104,In_286,In_83);
nor U105 (N_105,In_1132,In_1817);
nor U106 (N_106,In_703,In_577);
and U107 (N_107,In_1716,In_1707);
or U108 (N_108,In_1131,In_1138);
and U109 (N_109,In_1652,In_581);
or U110 (N_110,In_1967,In_1789);
and U111 (N_111,In_137,In_1100);
nand U112 (N_112,In_1842,In_426);
nand U113 (N_113,In_1263,In_296);
and U114 (N_114,In_1675,In_1696);
xor U115 (N_115,In_1338,In_1407);
and U116 (N_116,In_208,In_949);
and U117 (N_117,In_1722,In_1201);
nor U118 (N_118,In_1000,In_89);
and U119 (N_119,In_873,In_135);
and U120 (N_120,In_899,In_1194);
nand U121 (N_121,In_1041,In_524);
xnor U122 (N_122,In_350,In_1371);
and U123 (N_123,In_1860,In_1401);
xor U124 (N_124,In_1769,In_1359);
nor U125 (N_125,In_377,In_1025);
nand U126 (N_126,In_1372,In_1845);
nor U127 (N_127,In_1439,In_417);
and U128 (N_128,In_730,In_1052);
and U129 (N_129,In_1627,In_1334);
nor U130 (N_130,In_1363,In_82);
xor U131 (N_131,In_87,In_1108);
xor U132 (N_132,In_649,In_1932);
or U133 (N_133,In_997,In_1075);
nand U134 (N_134,In_454,In_1662);
or U135 (N_135,In_102,In_1007);
nor U136 (N_136,In_259,In_954);
or U137 (N_137,In_1275,In_1466);
nor U138 (N_138,In_963,In_521);
nor U139 (N_139,In_1724,In_299);
nand U140 (N_140,In_1298,In_1061);
or U141 (N_141,In_314,In_1843);
nor U142 (N_142,In_422,In_1159);
and U143 (N_143,In_613,In_275);
or U144 (N_144,In_814,In_1480);
and U145 (N_145,In_879,In_31);
and U146 (N_146,In_1717,In_1278);
or U147 (N_147,In_1471,In_606);
or U148 (N_148,In_1478,In_552);
nor U149 (N_149,In_754,In_983);
or U150 (N_150,In_1647,In_1764);
and U151 (N_151,In_1366,In_929);
or U152 (N_152,In_1973,In_1208);
or U153 (N_153,In_642,In_1534);
and U154 (N_154,In_143,In_912);
nand U155 (N_155,In_496,In_1483);
or U156 (N_156,In_445,In_862);
or U157 (N_157,In_134,In_795);
or U158 (N_158,In_796,In_202);
xor U159 (N_159,In_29,In_695);
and U160 (N_160,In_1510,In_1765);
xnor U161 (N_161,In_414,In_1563);
and U162 (N_162,In_1909,In_1325);
or U163 (N_163,In_637,In_538);
and U164 (N_164,In_914,In_225);
or U165 (N_165,In_993,In_1572);
or U166 (N_166,In_648,In_652);
or U167 (N_167,In_497,In_1327);
or U168 (N_168,In_1806,In_1020);
and U169 (N_169,In_697,In_843);
or U170 (N_170,In_1741,In_1993);
nor U171 (N_171,In_623,In_1590);
nor U172 (N_172,In_1644,In_1566);
nand U173 (N_173,In_856,In_1803);
nor U174 (N_174,In_752,In_1708);
nor U175 (N_175,In_1346,In_848);
or U176 (N_176,In_976,In_798);
nand U177 (N_177,In_269,In_1006);
or U178 (N_178,In_488,In_268);
nand U179 (N_179,In_1576,In_785);
nand U180 (N_180,In_1711,In_1602);
xor U181 (N_181,In_566,In_1757);
nor U182 (N_182,In_385,In_1669);
and U183 (N_183,In_354,In_959);
or U184 (N_184,In_1040,In_1674);
nand U185 (N_185,In_1115,In_1846);
nor U186 (N_186,In_302,In_424);
and U187 (N_187,In_434,In_631);
nor U188 (N_188,In_508,In_1035);
nand U189 (N_189,In_768,In_570);
and U190 (N_190,In_947,In_1192);
nand U191 (N_191,In_906,In_72);
xor U192 (N_192,In_242,In_678);
nand U193 (N_193,In_1788,In_844);
and U194 (N_194,In_1421,In_1376);
nand U195 (N_195,In_77,In_1819);
nand U196 (N_196,In_237,In_1400);
or U197 (N_197,In_726,In_387);
nand U198 (N_198,In_153,In_335);
nand U199 (N_199,In_553,In_1999);
xnor U200 (N_200,In_1760,In_258);
or U201 (N_201,In_943,In_741);
and U202 (N_202,In_1779,In_1504);
and U203 (N_203,In_1880,In_471);
xor U204 (N_204,In_1673,In_337);
nor U205 (N_205,In_26,In_841);
nor U206 (N_206,In_81,In_786);
nand U207 (N_207,In_1903,In_1452);
nor U208 (N_208,In_1700,In_1833);
nand U209 (N_209,In_1918,In_889);
nand U210 (N_210,In_1509,In_1888);
nand U211 (N_211,In_647,In_1336);
and U212 (N_212,In_1445,In_828);
or U213 (N_213,In_1288,In_1936);
nor U214 (N_214,In_1092,In_791);
nor U215 (N_215,In_1461,In_893);
and U216 (N_216,In_568,In_1927);
or U217 (N_217,In_1137,In_213);
and U218 (N_218,In_4,In_863);
nor U219 (N_219,In_28,In_59);
or U220 (N_220,In_480,In_1073);
xor U221 (N_221,In_1917,In_835);
or U222 (N_222,In_1907,In_672);
nand U223 (N_223,In_1823,In_1002);
and U224 (N_224,In_324,In_325);
and U225 (N_225,In_1229,In_1243);
nor U226 (N_226,In_1031,In_1250);
nor U227 (N_227,In_1024,In_640);
nand U228 (N_228,In_1067,In_901);
and U229 (N_229,In_375,In_1384);
or U230 (N_230,In_94,In_790);
and U231 (N_231,In_860,In_1929);
nor U232 (N_232,In_1428,In_282);
nand U233 (N_233,In_223,In_628);
nand U234 (N_234,In_994,In_1962);
or U235 (N_235,In_712,In_859);
nand U236 (N_236,In_490,In_1349);
nand U237 (N_237,In_295,In_69);
nor U238 (N_238,In_512,In_1311);
and U239 (N_239,In_32,In_1683);
xnor U240 (N_240,In_1658,In_1926);
or U241 (N_241,In_840,In_1482);
xor U242 (N_242,In_1151,In_1772);
or U243 (N_243,In_1030,In_1487);
or U244 (N_244,In_1588,In_985);
nand U245 (N_245,In_1981,In_428);
nor U246 (N_246,In_1844,In_987);
xor U247 (N_247,In_593,In_185);
and U248 (N_248,In_1751,In_369);
nor U249 (N_249,In_1840,In_1871);
and U250 (N_250,In_450,In_1265);
nand U251 (N_251,In_1735,In_381);
or U252 (N_252,In_147,In_729);
or U253 (N_253,In_965,In_962);
nor U254 (N_254,In_780,In_951);
nand U255 (N_255,In_1352,In_1744);
and U256 (N_256,In_1200,In_35);
nor U257 (N_257,In_1719,In_1889);
nor U258 (N_258,In_1167,In_1168);
or U259 (N_259,In_833,In_98);
nor U260 (N_260,In_772,In_509);
xor U261 (N_261,In_207,In_1426);
nand U262 (N_262,In_1337,In_1185);
nand U263 (N_263,In_1834,In_1432);
or U264 (N_264,In_60,In_1596);
and U265 (N_265,In_812,In_1331);
nor U266 (N_266,In_1302,In_443);
or U267 (N_267,In_1435,In_234);
or U268 (N_268,In_1982,In_832);
nand U269 (N_269,In_1899,In_289);
nand U270 (N_270,In_1162,In_249);
nor U271 (N_271,In_1164,In_626);
nor U272 (N_272,In_316,In_715);
and U273 (N_273,In_684,In_698);
nand U274 (N_274,In_67,In_204);
nand U275 (N_275,In_861,In_974);
nand U276 (N_276,In_1687,In_1036);
nand U277 (N_277,In_892,In_534);
nor U278 (N_278,In_565,In_868);
nor U279 (N_279,In_1732,In_493);
and U280 (N_280,In_1783,In_1727);
nor U281 (N_281,In_1793,In_717);
and U282 (N_282,In_430,In_330);
nor U283 (N_283,In_736,In_1965);
nor U284 (N_284,In_176,In_960);
or U285 (N_285,In_501,In_1663);
nor U286 (N_286,In_1190,In_588);
and U287 (N_287,In_1004,In_1297);
and U288 (N_288,In_447,In_526);
and U289 (N_289,In_92,In_1826);
nand U290 (N_290,In_139,In_218);
or U291 (N_291,In_671,In_183);
xor U292 (N_292,In_1919,In_1610);
and U293 (N_293,In_68,In_1560);
and U294 (N_294,In_1958,In_1385);
and U295 (N_295,In_1987,In_1354);
and U296 (N_296,In_981,In_1976);
nor U297 (N_297,In_1144,In_1546);
and U298 (N_298,In_1043,In_1592);
nand U299 (N_299,In_705,In_129);
nand U300 (N_300,In_1447,In_1370);
and U301 (N_301,In_1207,In_1887);
or U302 (N_302,In_591,In_1545);
and U303 (N_303,In_1214,In_1614);
nor U304 (N_304,In_884,In_563);
or U305 (N_305,In_233,In_1812);
nor U306 (N_306,In_1524,In_690);
nor U307 (N_307,In_1058,In_240);
nor U308 (N_308,In_1770,In_1046);
nor U309 (N_309,In_1442,In_1537);
and U310 (N_310,In_1628,In_1205);
nor U311 (N_311,In_602,In_1664);
nand U312 (N_312,In_557,In_476);
nand U313 (N_313,In_992,In_6);
or U314 (N_314,In_1496,In_276);
nand U315 (N_315,In_448,In_190);
xor U316 (N_316,In_1145,In_1475);
nor U317 (N_317,In_425,In_1113);
nor U318 (N_318,In_1996,In_622);
nand U319 (N_319,In_931,In_881);
nor U320 (N_320,In_11,In_70);
nor U321 (N_321,In_110,In_95);
xnor U322 (N_322,In_283,In_519);
nor U323 (N_323,In_853,In_125);
nor U324 (N_324,In_320,In_1931);
or U325 (N_325,In_1666,In_543);
nor U326 (N_326,In_507,In_1105);
nor U327 (N_327,In_1285,In_301);
nor U328 (N_328,In_457,In_745);
nand U329 (N_329,In_198,In_1222);
and U330 (N_330,In_1702,In_1011);
nor U331 (N_331,In_874,In_595);
xor U332 (N_332,In_1176,In_646);
nand U333 (N_333,In_64,In_1513);
xor U334 (N_334,In_1577,In_513);
nand U335 (N_335,In_163,In_550);
or U336 (N_336,In_617,In_1611);
xnor U337 (N_337,In_1125,In_93);
and U338 (N_338,In_1992,In_1665);
and U339 (N_339,In_1429,In_872);
nor U340 (N_340,In_1601,In_181);
nand U341 (N_341,In_88,In_1438);
nand U342 (N_342,In_406,In_559);
nor U343 (N_343,In_1550,In_40);
nand U344 (N_344,In_1940,In_397);
nor U345 (N_345,In_1409,In_1989);
or U346 (N_346,In_1239,In_1066);
or U347 (N_347,In_1597,In_162);
and U348 (N_348,In_75,In_132);
and U349 (N_349,In_529,In_781);
nor U350 (N_350,In_184,In_1877);
and U351 (N_351,In_39,In_1473);
nand U352 (N_352,In_1985,In_284);
and U353 (N_353,In_1905,In_187);
nand U354 (N_354,In_285,In_1624);
nor U355 (N_355,In_482,In_1348);
or U356 (N_356,In_1233,In_720);
nor U357 (N_357,In_1506,In_499);
and U358 (N_358,In_1520,In_643);
nand U359 (N_359,In_1286,In_1156);
nand U360 (N_360,In_341,In_531);
and U361 (N_361,In_1287,In_1253);
nor U362 (N_362,In_200,In_1911);
nand U363 (N_363,In_688,In_1629);
nor U364 (N_364,In_522,In_821);
nor U365 (N_365,In_449,In_13);
nor U366 (N_366,In_1867,In_1303);
or U367 (N_367,In_262,In_696);
nor U368 (N_368,In_174,In_1956);
xnor U369 (N_369,In_1489,In_704);
nand U370 (N_370,In_1948,In_336);
and U371 (N_371,In_1692,In_1218);
nor U372 (N_372,In_46,In_1247);
xnor U373 (N_373,In_311,In_1153);
and U374 (N_374,In_727,In_359);
and U375 (N_375,In_131,In_1693);
and U376 (N_376,In_1015,In_1848);
and U377 (N_377,In_1815,In_1836);
or U378 (N_378,In_380,In_1883);
nor U379 (N_379,In_773,In_418);
and U380 (N_380,In_733,In_251);
nand U381 (N_381,In_1146,In_1643);
xnor U382 (N_382,In_1706,In_603);
or U383 (N_383,In_344,In_813);
and U384 (N_384,In_916,In_1259);
and U385 (N_385,In_464,In_572);
nor U386 (N_386,In_334,In_1368);
or U387 (N_387,In_818,In_264);
nor U388 (N_388,In_749,In_1782);
and U389 (N_389,In_1391,In_332);
or U390 (N_390,In_1567,In_1555);
and U391 (N_391,In_323,In_632);
nor U392 (N_392,In_1310,In_1736);
and U393 (N_393,In_483,In_1276);
xor U394 (N_394,In_645,In_1837);
nor U395 (N_395,In_1017,In_1802);
or U396 (N_396,In_157,In_1878);
nand U397 (N_397,In_575,In_857);
and U398 (N_398,In_165,In_824);
nand U399 (N_399,In_1460,In_79);
nor U400 (N_400,In_429,In_510);
nand U401 (N_401,In_1345,In_1925);
nor U402 (N_402,In_927,In_1057);
nor U403 (N_403,In_104,In_300);
nand U404 (N_404,In_1032,In_273);
nand U405 (N_405,In_718,In_378);
nor U406 (N_406,In_1568,In_221);
nand U407 (N_407,In_142,In_1778);
nor U408 (N_408,In_1330,In_664);
and U409 (N_409,In_1688,In_1668);
and U410 (N_410,In_339,In_1530);
nor U411 (N_411,In_50,In_470);
nand U412 (N_412,In_787,In_1485);
nor U413 (N_413,In_1324,In_36);
xor U414 (N_414,In_217,In_1456);
nand U415 (N_415,In_1110,In_854);
xor U416 (N_416,In_1619,In_1851);
nor U417 (N_417,In_327,In_614);
nand U418 (N_418,In_817,In_1063);
or U419 (N_419,In_1904,In_544);
nand U420 (N_420,In_532,In_1304);
xor U421 (N_421,In_352,In_85);
and U422 (N_422,In_1676,In_303);
or U423 (N_423,In_1394,In_520);
nand U424 (N_424,In_353,In_761);
and U425 (N_425,In_902,In_1920);
or U426 (N_426,In_261,In_1016);
or U427 (N_427,In_548,In_63);
or U428 (N_428,In_956,In_30);
and U429 (N_429,In_1402,In_1689);
and U430 (N_430,In_105,In_864);
and U431 (N_431,In_740,In_317);
and U432 (N_432,In_598,In_279);
nand U433 (N_433,In_1014,In_232);
xnor U434 (N_434,In_1150,In_1344);
and U435 (N_435,In_427,In_1559);
or U436 (N_436,In_1809,In_260);
and U437 (N_437,In_1852,In_439);
nor U438 (N_438,In_113,In_1342);
nand U439 (N_439,In_1951,In_395);
nor U440 (N_440,In_629,In_277);
nor U441 (N_441,In_620,In_1885);
and U442 (N_442,In_1224,In_627);
nand U443 (N_443,In_918,In_41);
and U444 (N_444,In_111,In_1938);
or U445 (N_445,In_608,In_45);
or U446 (N_446,In_762,In_1584);
and U447 (N_447,In_751,In_201);
nand U448 (N_448,In_1217,In_1264);
nor U449 (N_449,In_1726,In_528);
and U450 (N_450,In_890,In_106);
or U451 (N_451,In_1990,In_789);
or U452 (N_452,In_1955,In_1140);
nand U453 (N_453,In_1822,In_920);
xor U454 (N_454,In_989,In_1396);
nor U455 (N_455,In_433,In_656);
or U456 (N_456,In_1281,In_517);
and U457 (N_457,In_319,In_1913);
nor U458 (N_458,In_1620,In_1120);
nor U459 (N_459,In_1431,In_883);
nor U460 (N_460,In_1398,In_978);
xor U461 (N_461,In_1147,In_689);
and U462 (N_462,In_1656,In_1564);
and U463 (N_463,In_1451,In_1771);
or U464 (N_464,In_1134,In_1818);
or U465 (N_465,In_551,In_1335);
nand U466 (N_466,In_1725,In_1154);
and U467 (N_467,In_1047,In_419);
or U468 (N_468,In_1607,In_760);
or U469 (N_469,In_1915,In_1070);
nand U470 (N_470,In_765,In_1273);
nand U471 (N_471,In_121,In_1126);
or U472 (N_472,In_1314,In_1076);
nor U473 (N_473,In_1569,In_525);
nor U474 (N_474,In_500,In_1552);
or U475 (N_475,In_1849,In_919);
and U476 (N_476,In_721,In_1245);
nor U477 (N_477,In_1223,In_1101);
or U478 (N_478,In_411,In_413);
nand U479 (N_479,In_96,In_1300);
or U480 (N_480,In_408,In_17);
nand U481 (N_481,In_410,In_830);
and U482 (N_482,In_1458,In_1859);
nor U483 (N_483,In_230,In_766);
nor U484 (N_484,In_1605,In_1875);
nand U485 (N_485,In_1021,In_1554);
and U486 (N_486,In_1516,In_368);
nand U487 (N_487,In_366,In_1672);
nand U488 (N_488,In_364,In_1599);
or U489 (N_489,In_1112,In_907);
xor U490 (N_490,In_1148,In_837);
nor U491 (N_491,In_1309,In_799);
or U492 (N_492,In_197,In_10);
xor U493 (N_493,In_1804,In_1399);
nor U494 (N_494,In_936,In_1197);
or U495 (N_495,In_120,In_1704);
xnor U496 (N_496,In_118,In_37);
xor U497 (N_497,In_792,In_644);
nor U498 (N_498,In_1318,In_850);
or U499 (N_499,In_1271,In_270);
or U500 (N_500,In_71,In_1455);
and U501 (N_501,In_858,In_1241);
or U502 (N_502,In_1733,In_1847);
nor U503 (N_503,In_677,In_349);
nor U504 (N_504,In_1679,In_108);
nor U505 (N_505,In_374,In_25);
or U506 (N_506,In_1169,In_1141);
and U507 (N_507,In_661,In_803);
nor U508 (N_508,In_152,In_783);
nor U509 (N_509,In_980,In_1681);
xor U510 (N_510,In_1444,In_882);
nand U511 (N_511,In_188,In_1525);
nand U512 (N_512,In_933,In_1828);
or U513 (N_513,In_1701,In_1282);
nand U514 (N_514,In_1841,In_1616);
or U515 (N_515,In_1949,In_244);
nand U516 (N_516,In_80,In_54);
or U517 (N_517,In_1196,In_1414);
or U518 (N_518,In_1494,In_1763);
or U519 (N_519,In_463,In_1969);
and U520 (N_520,In_112,In_437);
nand U521 (N_521,In_576,In_1013);
nor U522 (N_522,In_659,In_579);
nand U523 (N_523,In_38,In_1795);
or U524 (N_524,In_567,In_383);
xor U525 (N_525,In_166,In_241);
and U526 (N_526,In_76,In_1450);
nand U527 (N_527,In_771,In_126);
and U528 (N_528,In_144,In_1881);
nor U529 (N_529,In_307,In_1536);
nor U530 (N_530,In_272,In_1754);
nand U531 (N_531,In_435,In_865);
or U532 (N_532,In_391,In_1661);
nor U533 (N_533,In_1157,In_1258);
nand U534 (N_534,In_934,In_1329);
or U535 (N_535,In_5,In_1306);
or U536 (N_536,In_573,In_801);
and U537 (N_537,In_540,In_371);
or U538 (N_538,In_1074,In_554);
nand U539 (N_539,In_292,In_1573);
nor U540 (N_540,In_1691,In_1503);
or U541 (N_541,In_903,In_1019);
or U542 (N_542,In_887,In_913);
xnor U543 (N_543,In_1978,In_891);
nand U544 (N_544,In_1645,In_904);
nand U545 (N_545,In_247,In_748);
and U546 (N_546,In_494,In_1195);
nand U547 (N_547,In_1178,In_764);
or U548 (N_548,In_148,In_1755);
and U549 (N_549,In_1872,In_1638);
nor U550 (N_550,In_466,In_831);
nand U551 (N_551,In_1625,In_62);
nor U552 (N_552,In_1382,In_1728);
and U553 (N_553,In_172,In_1051);
xor U554 (N_554,In_1553,In_119);
or U555 (N_555,In_287,In_1642);
nand U556 (N_556,In_1622,In_1857);
or U557 (N_557,In_685,In_811);
nor U558 (N_558,In_991,In_1747);
nand U559 (N_559,In_1252,In_839);
nor U560 (N_560,In_298,In_589);
or U561 (N_561,In_1776,In_146);
xnor U562 (N_562,In_758,In_1916);
nor U563 (N_563,In_1561,In_1079);
nand U564 (N_564,In_1361,In_823);
nor U565 (N_565,In_1089,In_1587);
nor U566 (N_566,In_216,In_1216);
nor U567 (N_567,In_601,In_1260);
and U568 (N_568,In_367,In_1033);
or U569 (N_569,In_639,In_186);
nor U570 (N_570,In_1972,In_1418);
and U571 (N_571,In_1320,In_1448);
or U572 (N_572,In_56,In_1215);
nand U573 (N_573,In_1910,In_1810);
nand U574 (N_574,In_1677,In_1180);
or U575 (N_575,In_1527,In_1044);
and U576 (N_576,In_161,In_238);
or U577 (N_577,In_487,In_797);
and U578 (N_578,In_34,In_485);
nor U579 (N_579,In_115,In_1405);
and U580 (N_580,In_141,In_281);
and U581 (N_581,In_1165,In_722);
nand U582 (N_582,In_189,In_1825);
or U583 (N_583,In_984,In_1121);
xor U584 (N_584,In_280,In_609);
xnor U585 (N_585,In_713,In_1968);
xnor U586 (N_586,In_655,In_1873);
nand U587 (N_587,In_1449,In_1856);
nor U588 (N_588,In_1266,In_999);
and U589 (N_589,In_806,In_779);
nand U590 (N_590,In_1558,In_898);
nand U591 (N_591,In_1179,In_1039);
nand U592 (N_592,In_775,In_145);
nand U593 (N_593,In_1173,In_1977);
nor U594 (N_594,In_1053,In_1617);
nand U595 (N_595,In_1313,In_1050);
or U596 (N_596,In_1971,In_1172);
and U597 (N_597,In_211,In_1914);
nor U598 (N_598,In_735,In_518);
nand U599 (N_599,In_1753,In_1246);
xnor U600 (N_600,In_328,In_309);
nand U601 (N_601,In_1791,In_746);
nor U602 (N_602,In_1133,In_1984);
nor U603 (N_603,In_1369,In_1446);
nand U604 (N_604,In_1773,In_1532);
or U605 (N_605,In_91,In_1158);
and U606 (N_606,In_1533,In_1474);
xnor U607 (N_607,In_226,In_1549);
or U608 (N_608,In_1538,In_243);
nand U609 (N_609,In_702,In_1511);
and U610 (N_610,In_409,In_674);
xnor U611 (N_611,In_456,In_248);
or U612 (N_612,In_1523,In_254);
xor U613 (N_613,In_246,In_1321);
and U614 (N_614,In_505,In_1143);
nor U615 (N_615,In_1377,In_1284);
or U616 (N_616,In_1921,In_220);
nand U617 (N_617,In_1730,In_1453);
nor U618 (N_618,In_971,In_401);
and U619 (N_619,In_24,In_660);
and U620 (N_620,In_1139,In_1720);
and U621 (N_621,In_1797,In_1182);
nand U622 (N_622,In_616,In_676);
and U623 (N_623,In_810,In_1667);
or U624 (N_624,In_1332,In_1835);
or U625 (N_625,In_1886,In_1242);
nor U626 (N_626,In_1174,In_388);
and U627 (N_627,In_1269,In_955);
nand U628 (N_628,In_742,In_1970);
or U629 (N_629,In_605,In_988);
or U630 (N_630,In_460,In_1798);
nand U631 (N_631,In_996,In_1378);
xnor U632 (N_632,In_666,In_1780);
and U633 (N_633,In_1210,In_1268);
and U634 (N_634,In_851,In_1206);
and U635 (N_635,In_1713,In_1430);
nand U636 (N_636,In_558,In_1578);
nand U637 (N_637,In_306,In_1671);
nor U638 (N_638,In_1526,In_537);
or U639 (N_639,In_1768,In_376);
or U640 (N_640,In_966,In_1586);
nand U641 (N_641,In_1551,In_578);
xor U642 (N_642,In_641,In_78);
and U643 (N_643,In_1123,In_523);
or U644 (N_644,In_826,In_8);
and U645 (N_645,In_1467,In_382);
and U646 (N_646,In_683,In_547);
or U647 (N_647,In_293,In_1186);
nand U648 (N_648,In_681,In_969);
nand U649 (N_649,In_753,In_239);
nor U650 (N_650,In_486,In_66);
or U651 (N_651,In_594,In_1425);
nand U652 (N_652,In_1493,In_1562);
nand U653 (N_653,In_596,In_679);
nor U654 (N_654,In_42,In_998);
nor U655 (N_655,In_1481,In_155);
or U656 (N_656,In_191,In_15);
or U657 (N_657,In_515,In_808);
or U658 (N_658,In_192,In_441);
nand U659 (N_659,In_236,In_1109);
and U660 (N_660,In_1699,In_1312);
nor U661 (N_661,In_506,In_1544);
or U662 (N_662,In_9,In_227);
and U663 (N_663,In_1262,In_1777);
or U664 (N_664,In_1389,In_1362);
or U665 (N_665,In_290,In_86);
nand U666 (N_666,In_256,In_1272);
and U667 (N_667,In_816,In_73);
or U668 (N_668,In_1756,In_1069);
nand U669 (N_669,In_1048,In_1411);
nand U670 (N_670,In_1440,In_1705);
nand U671 (N_671,In_847,In_150);
and U672 (N_672,In_804,In_1497);
nor U673 (N_673,In_1930,In_1423);
or U674 (N_674,In_1901,In_580);
nand U675 (N_675,In_346,In_1476);
nor U676 (N_676,In_1994,In_1049);
and U677 (N_677,In_1404,In_1570);
nand U678 (N_678,In_1062,In_937);
and U679 (N_679,In_1009,In_265);
or U680 (N_680,In_154,In_1270);
or U681 (N_681,In_1130,In_910);
or U682 (N_682,In_194,In_467);
nand U683 (N_683,In_763,In_18);
and U684 (N_684,In_802,In_1945);
and U685 (N_685,In_1589,In_630);
xnor U686 (N_686,In_1319,In_1801);
nand U687 (N_687,In_1900,In_585);
nor U688 (N_688,In_305,In_896);
or U689 (N_689,In_1037,In_728);
nand U690 (N_690,In_1738,In_1381);
nand U691 (N_691,In_961,In_1034);
nor U692 (N_692,In_979,In_1054);
xnor U693 (N_693,In_587,In_109);
nand U694 (N_694,In_212,In_1603);
nand U695 (N_695,In_1419,In_1459);
and U696 (N_696,In_1161,In_612);
nand U697 (N_697,In_1807,In_957);
nand U698 (N_698,In_432,In_229);
xnor U699 (N_699,In_1698,In_12);
nor U700 (N_700,In_1874,In_1684);
and U701 (N_701,In_1301,In_250);
or U702 (N_702,In_1947,In_171);
nand U703 (N_703,In_542,In_1142);
nor U704 (N_704,In_877,In_541);
or U705 (N_705,In_946,In_1119);
and U706 (N_706,In_1829,In_228);
nor U707 (N_707,In_478,In_1814);
and U708 (N_708,In_1980,In_1582);
nor U709 (N_709,In_1519,In_459);
xnor U710 (N_710,In_900,In_1811);
or U711 (N_711,In_1071,In_1427);
nand U712 (N_712,In_351,In_1865);
nand U713 (N_713,In_1028,In_1499);
nand U714 (N_714,In_22,In_1234);
nand U715 (N_715,In_908,In_977);
xor U716 (N_716,In_737,In_1283);
nand U717 (N_717,In_1618,In_1068);
xor U718 (N_718,In_1209,In_175);
nor U719 (N_719,In_1879,In_1230);
nand U720 (N_720,In_1029,In_357);
or U721 (N_721,In_1715,In_635);
and U722 (N_722,In_1358,In_1651);
nor U723 (N_723,In_1081,In_356);
or U724 (N_724,In_1322,In_1864);
and U725 (N_725,In_842,In_1556);
or U726 (N_726,In_274,In_1858);
and U727 (N_727,In_1547,In_1118);
and U728 (N_728,In_1340,In_1103);
nand U729 (N_729,In_90,In_930);
nor U730 (N_730,In_1923,In_1739);
and U731 (N_731,In_921,In_1655);
and U732 (N_732,In_1373,In_1541);
nand U733 (N_733,In_484,In_1542);
or U734 (N_734,In_1128,In_599);
and U735 (N_735,In_950,In_815);
nor U736 (N_736,In_1585,In_1116);
or U737 (N_737,In_278,In_489);
and U738 (N_738,In_224,In_1360);
nor U739 (N_739,In_1745,In_982);
nand U740 (N_740,In_836,In_767);
or U741 (N_741,In_340,In_294);
nand U742 (N_742,In_140,In_1416);
nand U743 (N_743,In_710,In_1896);
nor U744 (N_744,In_1678,In_179);
xor U745 (N_745,In_461,In_668);
and U746 (N_746,In_1003,In_313);
xor U747 (N_747,In_928,In_1056);
or U748 (N_748,In_1392,In_784);
or U749 (N_749,In_1220,In_1307);
nor U750 (N_750,In_348,In_1649);
xnor U751 (N_751,In_203,In_1934);
and U752 (N_752,In_1623,In_1529);
and U753 (N_753,In_1986,In_829);
or U754 (N_754,In_310,In_124);
xnor U755 (N_755,In_1964,In_1351);
nor U756 (N_756,In_1027,In_127);
nor U757 (N_757,In_1379,In_164);
and U758 (N_758,In_707,In_876);
nor U759 (N_759,In_1479,In_1022);
nor U760 (N_760,In_1077,In_1339);
nand U761 (N_761,In_412,In_536);
nand U762 (N_762,In_967,In_1654);
and U763 (N_763,In_1633,In_1740);
or U764 (N_764,In_100,In_1203);
or U765 (N_765,In_1437,In_1785);
xnor U766 (N_766,In_1225,In_1933);
and U767 (N_767,In_1543,In_1502);
xor U768 (N_768,In_1078,In_379);
and U769 (N_769,In_1498,In_747);
nand U770 (N_770,In_1694,In_291);
or U771 (N_771,In_416,In_938);
or U772 (N_772,In_1279,In_675);
nand U773 (N_773,In_1045,In_1038);
and U774 (N_774,In_1600,In_326);
and U775 (N_775,In_1609,In_193);
nor U776 (N_776,In_1876,In_1221);
nand U777 (N_777,In_1082,In_886);
or U778 (N_778,In_436,In_1023);
and U779 (N_779,In_1387,In_1512);
and U780 (N_780,In_1659,In_1187);
nor U781 (N_781,In_1171,In_827);
or U782 (N_782,In_1294,In_209);
nand U783 (N_783,In_1853,In_849);
and U784 (N_784,In_866,In_1507);
and U785 (N_785,In_607,In_1251);
nor U786 (N_786,In_1238,In_170);
or U787 (N_787,In_776,In_1868);
nor U788 (N_788,In_363,In_1129);
nor U789 (N_789,In_1477,In_1299);
nor U790 (N_790,In_870,In_271);
nor U791 (N_791,In_231,In_345);
and U792 (N_792,In_1734,In_590);
nor U793 (N_793,In_1749,In_1198);
or U794 (N_794,In_1202,In_1891);
and U795 (N_795,In_1417,In_952);
nand U796 (N_796,In_597,In_1462);
and U797 (N_797,In_584,In_1718);
and U798 (N_798,In_600,In_948);
or U799 (N_799,In_1784,In_477);
nand U800 (N_800,In_138,In_245);
xnor U801 (N_801,In_1292,In_304);
or U802 (N_802,In_1660,In_1821);
nor U803 (N_803,In_691,In_1787);
nor U804 (N_804,In_1571,In_922);
nand U805 (N_805,In_1839,In_530);
nor U806 (N_806,In_219,In_1884);
and U807 (N_807,In_923,In_1714);
or U808 (N_808,In_65,In_1721);
nand U809 (N_809,In_451,In_20);
or U810 (N_810,In_1184,In_1181);
and U811 (N_811,In_475,In_1114);
xnor U812 (N_812,In_1892,In_372);
and U813 (N_813,In_592,In_1998);
nor U814 (N_814,In_794,In_805);
or U815 (N_815,In_263,In_1341);
nand U816 (N_816,In_719,In_159);
and U817 (N_817,In_869,In_1422);
or U818 (N_818,In_1974,In_1767);
nand U819 (N_819,In_1598,In_738);
nor U820 (N_820,In_1122,In_1228);
nor U821 (N_821,In_1517,In_1219);
nand U822 (N_822,In_1731,In_1244);
nor U823 (N_823,In_1775,In_1861);
and U824 (N_824,In_1975,In_7);
and U825 (N_825,In_0,In_1991);
and U826 (N_826,In_23,In_1454);
or U827 (N_827,In_1650,In_1894);
nor U828 (N_828,In_205,In_699);
xnor U829 (N_829,In_1820,In_1059);
and U830 (N_830,In_845,In_774);
nand U831 (N_831,In_788,In_871);
or U832 (N_832,In_1255,In_958);
or U833 (N_833,In_1166,In_1838);
xnor U834 (N_834,In_1347,In_373);
nor U835 (N_835,In_1098,In_940);
nor U836 (N_836,In_288,In_420);
or U837 (N_837,In_897,In_1621);
nor U838 (N_838,In_1343,In_474);
xor U839 (N_839,In_178,In_1531);
nand U840 (N_840,In_173,In_1941);
xor U841 (N_841,In_1950,In_1632);
nand U842 (N_842,In_167,In_669);
and U843 (N_843,In_1703,In_1248);
nand U844 (N_844,In_778,In_1191);
nor U845 (N_845,In_1183,In_43);
and U846 (N_846,In_670,In_732);
nand U847 (N_847,In_27,In_555);
and U848 (N_848,In_1636,In_1583);
nand U849 (N_849,In_769,In_453);
nand U850 (N_850,In_878,In_1606);
and U851 (N_851,In_1869,In_1001);
and U852 (N_852,In_195,In_638);
nor U853 (N_853,In_1521,In_1906);
and U854 (N_854,In_342,In_1729);
nand U855 (N_855,In_495,In_667);
xor U856 (N_856,In_571,In_1748);
or U857 (N_857,In_1086,In_2);
nor U858 (N_858,In_663,In_255);
nor U859 (N_859,In_405,In_1505);
xnor U860 (N_860,In_658,In_169);
nor U861 (N_861,In_822,In_1758);
nor U862 (N_862,In_1912,In_650);
and U863 (N_863,In_182,In_168);
nor U864 (N_864,In_1160,In_58);
nor U865 (N_865,In_926,In_582);
or U866 (N_866,In_1710,In_1813);
or U867 (N_867,In_1055,In_1855);
or U868 (N_868,In_1960,In_1267);
or U869 (N_869,In_1635,In_1935);
or U870 (N_870,In_101,In_1367);
nor U871 (N_871,In_693,In_504);
nand U872 (N_872,In_941,In_423);
or U873 (N_873,In_1424,In_945);
nor U874 (N_874,In_1102,In_1226);
xor U875 (N_875,In_1395,In_440);
or U876 (N_876,In_266,In_1189);
and U877 (N_877,In_1026,In_52);
or U878 (N_878,In_1096,In_1743);
nor U879 (N_879,In_103,In_1357);
and U880 (N_880,In_1648,In_1175);
and U881 (N_881,In_846,In_1816);
or U882 (N_882,In_1953,In_782);
xnor U883 (N_883,In_1742,In_546);
nand U884 (N_884,In_539,In_1170);
and U885 (N_885,In_1866,In_1634);
and U886 (N_886,In_1289,In_1922);
and U887 (N_887,In_1084,In_706);
nand U888 (N_888,In_1090,In_1805);
or U889 (N_889,In_662,In_1604);
nor U890 (N_890,In_446,In_1211);
and U891 (N_891,In_915,In_651);
nand U892 (N_892,In_503,In_160);
and U893 (N_893,In_1093,In_1484);
and U894 (N_894,In_653,In_624);
nand U895 (N_895,In_1291,In_1408);
xor U896 (N_896,In_1641,In_1249);
and U897 (N_897,In_1328,In_365);
nand U898 (N_898,In_1508,In_442);
nand U899 (N_899,In_880,In_1850);
xnor U900 (N_900,In_431,In_1954);
or U901 (N_901,In_714,In_1613);
or U902 (N_902,In_1274,In_1792);
or U903 (N_903,In_1501,In_1712);
and U904 (N_904,In_759,In_16);
and U905 (N_905,In_99,In_1944);
or U906 (N_906,In_756,In_1117);
xnor U907 (N_907,In_1830,In_210);
nor U908 (N_908,In_1111,In_386);
nor U909 (N_909,In_1293,In_257);
nor U910 (N_910,In_1670,In_360);
or U911 (N_911,In_333,In_545);
nor U912 (N_912,In_394,In_1212);
nor U913 (N_913,In_694,In_1296);
nor U914 (N_914,In_133,In_1939);
and U915 (N_915,In_1317,In_252);
and U916 (N_916,In_1434,In_1902);
or U917 (N_917,In_1697,In_1995);
or U918 (N_918,In_743,In_315);
nor U919 (N_919,In_621,In_1403);
or U920 (N_920,In_1365,In_1072);
nor U921 (N_921,In_569,In_331);
and U922 (N_922,In_1575,In_809);
nand U923 (N_923,In_1528,In_1008);
nand U924 (N_924,In_1469,In_1463);
and U925 (N_925,In_953,In_793);
xnor U926 (N_926,In_61,In_514);
nand U927 (N_927,In_1690,In_1420);
nand U928 (N_928,In_1353,In_1832);
nor U929 (N_929,In_935,In_1410);
and U930 (N_930,In_1227,In_665);
nand U931 (N_931,In_130,In_1213);
nand U932 (N_932,In_1124,In_1295);
nor U933 (N_933,In_107,In_1152);
and U934 (N_934,In_1862,In_1893);
or U935 (N_935,In_618,In_1350);
and U936 (N_936,In_1863,In_1412);
or U937 (N_937,In_1433,In_633);
nand U938 (N_938,In_1762,In_491);
nand U939 (N_939,In_973,In_1761);
and U940 (N_940,In_253,In_158);
and U941 (N_941,In_48,In_1326);
or U942 (N_942,In_561,In_235);
xnor U943 (N_943,In_852,In_975);
nand U944 (N_944,In_1492,In_709);
nor U945 (N_945,In_1565,In_151);
or U946 (N_946,In_1500,In_731);
and U947 (N_947,In_1579,In_1686);
and U948 (N_948,In_21,In_1087);
and U949 (N_949,In_1786,In_1413);
or U950 (N_950,In_473,In_1149);
xor U951 (N_951,In_968,In_611);
xor U952 (N_952,In_452,In_564);
xor U953 (N_953,In_51,In_932);
nor U954 (N_954,In_384,In_392);
nor U955 (N_955,In_1983,In_492);
xor U956 (N_956,In_49,In_986);
and U957 (N_957,In_560,In_1397);
nor U958 (N_958,In_1808,In_925);
or U959 (N_959,In_1988,In_3);
xnor U960 (N_960,In_625,In_1870);
or U961 (N_961,In_1107,In_1646);
or U962 (N_962,In_1794,In_750);
nor U963 (N_963,In_1464,In_462);
nor U964 (N_964,In_1581,In_308);
or U965 (N_965,In_1937,In_1364);
xnor U966 (N_966,In_136,In_825);
or U967 (N_967,In_1236,In_1088);
nand U968 (N_968,In_944,In_1308);
or U969 (N_969,In_149,In_711);
nand U970 (N_970,In_1240,In_84);
nor U971 (N_971,In_734,In_692);
nand U972 (N_972,In_47,In_1091);
nor U973 (N_973,In_1574,In_1790);
or U974 (N_974,In_215,In_615);
nor U975 (N_975,In_1653,In_888);
nor U976 (N_976,In_1959,In_1631);
and U977 (N_977,In_1135,In_1005);
nand U978 (N_978,In_1064,In_438);
nor U979 (N_979,In_214,In_770);
or U980 (N_980,In_1737,In_680);
xnor U981 (N_981,In_1256,In_1042);
xor U982 (N_982,In_1095,In_117);
or U983 (N_983,In_1908,In_972);
nand U984 (N_984,In_1375,In_700);
nand U985 (N_985,In_604,In_1388);
nor U986 (N_986,In_1136,In_116);
nor U987 (N_987,In_465,In_619);
or U988 (N_988,In_511,In_1946);
and U989 (N_989,In_1548,In_1436);
or U990 (N_990,In_1957,In_1188);
nand U991 (N_991,In_1380,In_1356);
or U992 (N_992,In_297,In_1083);
xor U993 (N_993,In_1942,In_1406);
xnor U994 (N_994,In_686,In_1012);
nand U995 (N_995,In_57,In_415);
and U996 (N_996,In_14,In_1155);
nand U997 (N_997,In_1457,In_479);
nand U998 (N_998,In_1261,In_755);
or U999 (N_999,In_1277,In_403);
xnor U1000 (N_1000,In_758,In_1729);
or U1001 (N_1001,In_1935,In_1373);
and U1002 (N_1002,In_634,In_1960);
nor U1003 (N_1003,In_91,In_727);
nor U1004 (N_1004,In_525,In_1655);
nand U1005 (N_1005,In_533,In_1111);
nand U1006 (N_1006,In_929,In_1927);
nand U1007 (N_1007,In_901,In_1769);
or U1008 (N_1008,In_1243,In_1267);
or U1009 (N_1009,In_1447,In_1410);
and U1010 (N_1010,In_1796,In_1692);
nand U1011 (N_1011,In_851,In_1192);
and U1012 (N_1012,In_695,In_1068);
or U1013 (N_1013,In_845,In_266);
or U1014 (N_1014,In_592,In_94);
nand U1015 (N_1015,In_242,In_146);
and U1016 (N_1016,In_1689,In_268);
nor U1017 (N_1017,In_983,In_1778);
and U1018 (N_1018,In_1398,In_750);
and U1019 (N_1019,In_1354,In_1115);
or U1020 (N_1020,In_757,In_242);
nand U1021 (N_1021,In_1137,In_108);
or U1022 (N_1022,In_531,In_105);
or U1023 (N_1023,In_1941,In_1107);
and U1024 (N_1024,In_349,In_674);
xnor U1025 (N_1025,In_1744,In_843);
and U1026 (N_1026,In_1632,In_817);
xor U1027 (N_1027,In_190,In_578);
nand U1028 (N_1028,In_831,In_1421);
or U1029 (N_1029,In_707,In_67);
nor U1030 (N_1030,In_571,In_173);
xnor U1031 (N_1031,In_27,In_1066);
and U1032 (N_1032,In_691,In_647);
nor U1033 (N_1033,In_1366,In_1887);
and U1034 (N_1034,In_1719,In_661);
nor U1035 (N_1035,In_516,In_1294);
or U1036 (N_1036,In_1376,In_1308);
nor U1037 (N_1037,In_170,In_672);
or U1038 (N_1038,In_1455,In_583);
nand U1039 (N_1039,In_717,In_1135);
nand U1040 (N_1040,In_1580,In_1988);
or U1041 (N_1041,In_786,In_657);
and U1042 (N_1042,In_1860,In_257);
nor U1043 (N_1043,In_1094,In_1210);
nor U1044 (N_1044,In_1834,In_1468);
and U1045 (N_1045,In_6,In_263);
nor U1046 (N_1046,In_323,In_154);
or U1047 (N_1047,In_1910,In_1557);
nor U1048 (N_1048,In_874,In_754);
xor U1049 (N_1049,In_1528,In_567);
and U1050 (N_1050,In_5,In_866);
or U1051 (N_1051,In_240,In_1863);
nor U1052 (N_1052,In_1476,In_1244);
and U1053 (N_1053,In_1819,In_1781);
nor U1054 (N_1054,In_514,In_1706);
nor U1055 (N_1055,In_34,In_1894);
or U1056 (N_1056,In_1249,In_1114);
xor U1057 (N_1057,In_679,In_240);
or U1058 (N_1058,In_1566,In_110);
nand U1059 (N_1059,In_1727,In_1065);
nor U1060 (N_1060,In_602,In_1224);
or U1061 (N_1061,In_1565,In_976);
or U1062 (N_1062,In_517,In_1156);
nor U1063 (N_1063,In_1311,In_1483);
nand U1064 (N_1064,In_1058,In_1303);
nor U1065 (N_1065,In_1685,In_1027);
or U1066 (N_1066,In_1452,In_1588);
nand U1067 (N_1067,In_1164,In_192);
nand U1068 (N_1068,In_689,In_1963);
xor U1069 (N_1069,In_1806,In_571);
nand U1070 (N_1070,In_1789,In_1586);
nor U1071 (N_1071,In_793,In_966);
and U1072 (N_1072,In_1255,In_272);
nand U1073 (N_1073,In_1033,In_1091);
nand U1074 (N_1074,In_1507,In_1420);
or U1075 (N_1075,In_151,In_651);
nor U1076 (N_1076,In_382,In_710);
and U1077 (N_1077,In_711,In_1589);
nand U1078 (N_1078,In_1391,In_690);
nor U1079 (N_1079,In_398,In_418);
and U1080 (N_1080,In_1638,In_294);
nor U1081 (N_1081,In_1544,In_1115);
nor U1082 (N_1082,In_1641,In_1728);
and U1083 (N_1083,In_52,In_506);
or U1084 (N_1084,In_1537,In_41);
and U1085 (N_1085,In_172,In_1820);
nor U1086 (N_1086,In_1842,In_1313);
nand U1087 (N_1087,In_480,In_26);
nor U1088 (N_1088,In_1586,In_265);
or U1089 (N_1089,In_1632,In_712);
and U1090 (N_1090,In_565,In_1071);
nor U1091 (N_1091,In_419,In_1286);
nor U1092 (N_1092,In_598,In_336);
nor U1093 (N_1093,In_1714,In_1088);
nand U1094 (N_1094,In_649,In_1887);
or U1095 (N_1095,In_1106,In_1873);
and U1096 (N_1096,In_709,In_272);
or U1097 (N_1097,In_1994,In_13);
or U1098 (N_1098,In_1341,In_357);
nor U1099 (N_1099,In_1103,In_1268);
nand U1100 (N_1100,In_1805,In_1308);
or U1101 (N_1101,In_1743,In_1627);
or U1102 (N_1102,In_407,In_1444);
nand U1103 (N_1103,In_1371,In_220);
nor U1104 (N_1104,In_448,In_1566);
nand U1105 (N_1105,In_998,In_1204);
or U1106 (N_1106,In_1259,In_313);
or U1107 (N_1107,In_1614,In_868);
or U1108 (N_1108,In_587,In_1205);
and U1109 (N_1109,In_172,In_1943);
nand U1110 (N_1110,In_1111,In_1390);
and U1111 (N_1111,In_380,In_1823);
and U1112 (N_1112,In_84,In_457);
and U1113 (N_1113,In_628,In_1345);
and U1114 (N_1114,In_1976,In_1732);
nor U1115 (N_1115,In_945,In_1583);
nand U1116 (N_1116,In_1821,In_333);
nand U1117 (N_1117,In_799,In_1786);
nand U1118 (N_1118,In_88,In_1987);
or U1119 (N_1119,In_1972,In_558);
nand U1120 (N_1120,In_1362,In_1764);
and U1121 (N_1121,In_109,In_524);
nand U1122 (N_1122,In_1899,In_591);
or U1123 (N_1123,In_1521,In_1193);
nor U1124 (N_1124,In_669,In_1988);
xnor U1125 (N_1125,In_1915,In_682);
and U1126 (N_1126,In_1204,In_1141);
nand U1127 (N_1127,In_1385,In_1909);
or U1128 (N_1128,In_648,In_1305);
or U1129 (N_1129,In_702,In_1554);
nor U1130 (N_1130,In_669,In_1335);
xor U1131 (N_1131,In_251,In_596);
nor U1132 (N_1132,In_1123,In_433);
nor U1133 (N_1133,In_617,In_711);
nand U1134 (N_1134,In_782,In_584);
nor U1135 (N_1135,In_1055,In_1411);
nand U1136 (N_1136,In_29,In_306);
nand U1137 (N_1137,In_1718,In_548);
and U1138 (N_1138,In_1346,In_1883);
nand U1139 (N_1139,In_1219,In_1594);
and U1140 (N_1140,In_532,In_502);
and U1141 (N_1141,In_1600,In_1035);
nand U1142 (N_1142,In_1684,In_109);
nor U1143 (N_1143,In_1618,In_602);
and U1144 (N_1144,In_667,In_516);
nor U1145 (N_1145,In_409,In_1721);
or U1146 (N_1146,In_1659,In_438);
nor U1147 (N_1147,In_892,In_1948);
or U1148 (N_1148,In_1561,In_214);
and U1149 (N_1149,In_312,In_1557);
or U1150 (N_1150,In_216,In_436);
or U1151 (N_1151,In_1438,In_298);
or U1152 (N_1152,In_105,In_917);
or U1153 (N_1153,In_1606,In_655);
or U1154 (N_1154,In_1364,In_1834);
nor U1155 (N_1155,In_72,In_1390);
nor U1156 (N_1156,In_261,In_638);
nor U1157 (N_1157,In_1473,In_947);
xnor U1158 (N_1158,In_1516,In_1784);
nor U1159 (N_1159,In_94,In_882);
nor U1160 (N_1160,In_1564,In_1676);
or U1161 (N_1161,In_849,In_259);
nor U1162 (N_1162,In_1497,In_902);
or U1163 (N_1163,In_1496,In_1324);
nand U1164 (N_1164,In_421,In_60);
nand U1165 (N_1165,In_1877,In_792);
nor U1166 (N_1166,In_1444,In_684);
and U1167 (N_1167,In_344,In_1194);
xor U1168 (N_1168,In_1096,In_958);
and U1169 (N_1169,In_34,In_1099);
or U1170 (N_1170,In_269,In_747);
nand U1171 (N_1171,In_815,In_243);
nand U1172 (N_1172,In_336,In_1326);
or U1173 (N_1173,In_82,In_519);
nor U1174 (N_1174,In_1614,In_1723);
or U1175 (N_1175,In_778,In_1466);
and U1176 (N_1176,In_1379,In_1393);
nand U1177 (N_1177,In_652,In_201);
and U1178 (N_1178,In_1585,In_328);
or U1179 (N_1179,In_623,In_1374);
nor U1180 (N_1180,In_831,In_1818);
nand U1181 (N_1181,In_755,In_381);
nand U1182 (N_1182,In_25,In_1076);
nor U1183 (N_1183,In_1145,In_331);
nand U1184 (N_1184,In_464,In_363);
nand U1185 (N_1185,In_1934,In_9);
nand U1186 (N_1186,In_1414,In_828);
or U1187 (N_1187,In_1835,In_1739);
nor U1188 (N_1188,In_600,In_1062);
and U1189 (N_1189,In_1957,In_3);
and U1190 (N_1190,In_1170,In_433);
nor U1191 (N_1191,In_874,In_1580);
nor U1192 (N_1192,In_620,In_1685);
nor U1193 (N_1193,In_1377,In_584);
and U1194 (N_1194,In_576,In_432);
and U1195 (N_1195,In_888,In_869);
or U1196 (N_1196,In_845,In_710);
xnor U1197 (N_1197,In_1512,In_999);
or U1198 (N_1198,In_169,In_1109);
nand U1199 (N_1199,In_85,In_1977);
nand U1200 (N_1200,In_1596,In_1163);
or U1201 (N_1201,In_1933,In_252);
or U1202 (N_1202,In_438,In_1389);
and U1203 (N_1203,In_1459,In_450);
and U1204 (N_1204,In_1210,In_94);
xnor U1205 (N_1205,In_100,In_1340);
and U1206 (N_1206,In_873,In_64);
and U1207 (N_1207,In_1707,In_1952);
and U1208 (N_1208,In_1693,In_1315);
and U1209 (N_1209,In_1956,In_253);
xnor U1210 (N_1210,In_1376,In_875);
xor U1211 (N_1211,In_1373,In_1942);
nor U1212 (N_1212,In_88,In_1719);
and U1213 (N_1213,In_1364,In_796);
nor U1214 (N_1214,In_1588,In_1160);
or U1215 (N_1215,In_1516,In_1045);
xor U1216 (N_1216,In_1189,In_1353);
and U1217 (N_1217,In_93,In_571);
and U1218 (N_1218,In_1842,In_1476);
or U1219 (N_1219,In_928,In_872);
nand U1220 (N_1220,In_931,In_1588);
and U1221 (N_1221,In_1670,In_1104);
or U1222 (N_1222,In_279,In_208);
nand U1223 (N_1223,In_1477,In_1544);
nor U1224 (N_1224,In_1679,In_321);
nand U1225 (N_1225,In_282,In_880);
and U1226 (N_1226,In_1132,In_1957);
and U1227 (N_1227,In_1491,In_688);
xnor U1228 (N_1228,In_1761,In_862);
nand U1229 (N_1229,In_1563,In_30);
and U1230 (N_1230,In_1092,In_544);
nor U1231 (N_1231,In_1870,In_775);
nor U1232 (N_1232,In_1109,In_623);
and U1233 (N_1233,In_375,In_1045);
or U1234 (N_1234,In_1519,In_1052);
nor U1235 (N_1235,In_49,In_1221);
xor U1236 (N_1236,In_1267,In_1177);
or U1237 (N_1237,In_704,In_1638);
or U1238 (N_1238,In_609,In_1819);
xnor U1239 (N_1239,In_497,In_1167);
and U1240 (N_1240,In_1188,In_1706);
nor U1241 (N_1241,In_645,In_502);
nor U1242 (N_1242,In_86,In_1587);
nor U1243 (N_1243,In_1185,In_545);
or U1244 (N_1244,In_1192,In_837);
and U1245 (N_1245,In_869,In_95);
xnor U1246 (N_1246,In_1970,In_1612);
nor U1247 (N_1247,In_1244,In_882);
or U1248 (N_1248,In_761,In_748);
nand U1249 (N_1249,In_985,In_1558);
nand U1250 (N_1250,In_1288,In_265);
or U1251 (N_1251,In_793,In_725);
nand U1252 (N_1252,In_1398,In_1443);
nor U1253 (N_1253,In_675,In_816);
or U1254 (N_1254,In_816,In_78);
nand U1255 (N_1255,In_1692,In_1452);
nand U1256 (N_1256,In_1641,In_1868);
or U1257 (N_1257,In_1667,In_1250);
or U1258 (N_1258,In_1491,In_790);
nand U1259 (N_1259,In_1223,In_1498);
nor U1260 (N_1260,In_557,In_18);
and U1261 (N_1261,In_50,In_1397);
nor U1262 (N_1262,In_968,In_1112);
or U1263 (N_1263,In_1059,In_611);
and U1264 (N_1264,In_520,In_1863);
or U1265 (N_1265,In_1391,In_1771);
nand U1266 (N_1266,In_447,In_1602);
and U1267 (N_1267,In_153,In_1022);
or U1268 (N_1268,In_859,In_599);
nand U1269 (N_1269,In_1997,In_719);
xor U1270 (N_1270,In_320,In_386);
and U1271 (N_1271,In_469,In_1671);
nand U1272 (N_1272,In_1433,In_1760);
and U1273 (N_1273,In_324,In_624);
or U1274 (N_1274,In_53,In_541);
or U1275 (N_1275,In_1260,In_15);
nand U1276 (N_1276,In_1156,In_928);
nor U1277 (N_1277,In_1,In_1654);
nor U1278 (N_1278,In_1791,In_215);
and U1279 (N_1279,In_438,In_32);
nor U1280 (N_1280,In_1043,In_1028);
nand U1281 (N_1281,In_442,In_635);
nor U1282 (N_1282,In_1964,In_1667);
and U1283 (N_1283,In_60,In_1318);
and U1284 (N_1284,In_420,In_202);
nor U1285 (N_1285,In_1316,In_1449);
or U1286 (N_1286,In_1216,In_1038);
or U1287 (N_1287,In_579,In_1354);
or U1288 (N_1288,In_1813,In_823);
or U1289 (N_1289,In_956,In_1459);
or U1290 (N_1290,In_169,In_1468);
and U1291 (N_1291,In_1422,In_1878);
or U1292 (N_1292,In_1600,In_787);
xnor U1293 (N_1293,In_1652,In_870);
nor U1294 (N_1294,In_221,In_1249);
and U1295 (N_1295,In_457,In_105);
and U1296 (N_1296,In_298,In_714);
xnor U1297 (N_1297,In_1082,In_857);
nand U1298 (N_1298,In_494,In_1762);
or U1299 (N_1299,In_856,In_1580);
and U1300 (N_1300,In_451,In_1423);
nand U1301 (N_1301,In_1907,In_729);
and U1302 (N_1302,In_868,In_1477);
or U1303 (N_1303,In_627,In_543);
and U1304 (N_1304,In_868,In_1139);
and U1305 (N_1305,In_1015,In_1446);
nor U1306 (N_1306,In_1903,In_1247);
or U1307 (N_1307,In_1886,In_294);
nand U1308 (N_1308,In_1935,In_1677);
nand U1309 (N_1309,In_539,In_890);
nand U1310 (N_1310,In_1618,In_1824);
or U1311 (N_1311,In_257,In_1167);
or U1312 (N_1312,In_1094,In_1623);
or U1313 (N_1313,In_1207,In_41);
or U1314 (N_1314,In_1358,In_584);
and U1315 (N_1315,In_1683,In_1348);
and U1316 (N_1316,In_1175,In_1205);
or U1317 (N_1317,In_1269,In_1198);
nor U1318 (N_1318,In_575,In_914);
xor U1319 (N_1319,In_1917,In_1912);
and U1320 (N_1320,In_1174,In_209);
xor U1321 (N_1321,In_632,In_908);
nor U1322 (N_1322,In_1568,In_1708);
or U1323 (N_1323,In_1043,In_794);
or U1324 (N_1324,In_1739,In_490);
or U1325 (N_1325,In_1128,In_1798);
or U1326 (N_1326,In_20,In_606);
nand U1327 (N_1327,In_291,In_740);
xor U1328 (N_1328,In_751,In_52);
or U1329 (N_1329,In_1026,In_1778);
or U1330 (N_1330,In_1263,In_821);
xnor U1331 (N_1331,In_820,In_1759);
nor U1332 (N_1332,In_939,In_1800);
nand U1333 (N_1333,In_151,In_373);
or U1334 (N_1334,In_784,In_1179);
or U1335 (N_1335,In_1496,In_1923);
nor U1336 (N_1336,In_1632,In_1107);
or U1337 (N_1337,In_1866,In_96);
nor U1338 (N_1338,In_1537,In_1168);
nand U1339 (N_1339,In_463,In_727);
nand U1340 (N_1340,In_1536,In_1359);
and U1341 (N_1341,In_937,In_814);
nand U1342 (N_1342,In_1228,In_1988);
or U1343 (N_1343,In_1842,In_753);
xnor U1344 (N_1344,In_1664,In_78);
xnor U1345 (N_1345,In_206,In_1214);
nor U1346 (N_1346,In_391,In_306);
xor U1347 (N_1347,In_1559,In_1921);
or U1348 (N_1348,In_145,In_821);
nor U1349 (N_1349,In_102,In_487);
nand U1350 (N_1350,In_412,In_753);
or U1351 (N_1351,In_444,In_402);
and U1352 (N_1352,In_1299,In_178);
or U1353 (N_1353,In_228,In_446);
nor U1354 (N_1354,In_1858,In_431);
nor U1355 (N_1355,In_216,In_1981);
or U1356 (N_1356,In_1423,In_1085);
xor U1357 (N_1357,In_1462,In_1233);
or U1358 (N_1358,In_1051,In_358);
and U1359 (N_1359,In_1083,In_943);
or U1360 (N_1360,In_1273,In_847);
or U1361 (N_1361,In_1355,In_124);
nand U1362 (N_1362,In_1537,In_918);
and U1363 (N_1363,In_1220,In_1051);
nor U1364 (N_1364,In_1218,In_1971);
nand U1365 (N_1365,In_1352,In_131);
nor U1366 (N_1366,In_1283,In_1351);
and U1367 (N_1367,In_1972,In_806);
nand U1368 (N_1368,In_66,In_457);
nand U1369 (N_1369,In_425,In_1972);
nor U1370 (N_1370,In_202,In_162);
or U1371 (N_1371,In_64,In_1484);
or U1372 (N_1372,In_11,In_118);
or U1373 (N_1373,In_501,In_734);
nand U1374 (N_1374,In_1457,In_14);
nor U1375 (N_1375,In_970,In_664);
nand U1376 (N_1376,In_527,In_1441);
or U1377 (N_1377,In_1665,In_1258);
nand U1378 (N_1378,In_987,In_725);
xor U1379 (N_1379,In_1539,In_461);
and U1380 (N_1380,In_1152,In_541);
nor U1381 (N_1381,In_1290,In_480);
nor U1382 (N_1382,In_1375,In_60);
xor U1383 (N_1383,In_181,In_382);
or U1384 (N_1384,In_1535,In_661);
nand U1385 (N_1385,In_1371,In_817);
nor U1386 (N_1386,In_467,In_293);
or U1387 (N_1387,In_1959,In_393);
nand U1388 (N_1388,In_1013,In_193);
xnor U1389 (N_1389,In_1594,In_1323);
nor U1390 (N_1390,In_1827,In_1309);
nor U1391 (N_1391,In_1996,In_536);
nand U1392 (N_1392,In_7,In_634);
or U1393 (N_1393,In_702,In_1562);
or U1394 (N_1394,In_1966,In_1425);
nor U1395 (N_1395,In_1418,In_630);
xor U1396 (N_1396,In_1891,In_1104);
nand U1397 (N_1397,In_57,In_1597);
nand U1398 (N_1398,In_1942,In_1615);
or U1399 (N_1399,In_724,In_795);
or U1400 (N_1400,In_1734,In_376);
and U1401 (N_1401,In_1452,In_1798);
or U1402 (N_1402,In_1680,In_1212);
or U1403 (N_1403,In_1359,In_895);
nand U1404 (N_1404,In_525,In_1789);
nor U1405 (N_1405,In_1078,In_63);
xnor U1406 (N_1406,In_1048,In_988);
nor U1407 (N_1407,In_401,In_1259);
nor U1408 (N_1408,In_508,In_1802);
nor U1409 (N_1409,In_170,In_189);
nor U1410 (N_1410,In_131,In_603);
or U1411 (N_1411,In_637,In_688);
and U1412 (N_1412,In_1492,In_265);
nor U1413 (N_1413,In_1287,In_1923);
or U1414 (N_1414,In_269,In_1470);
nor U1415 (N_1415,In_30,In_976);
and U1416 (N_1416,In_775,In_957);
xor U1417 (N_1417,In_1157,In_824);
nor U1418 (N_1418,In_634,In_1923);
and U1419 (N_1419,In_340,In_419);
or U1420 (N_1420,In_85,In_1427);
or U1421 (N_1421,In_1266,In_1677);
and U1422 (N_1422,In_1765,In_625);
nor U1423 (N_1423,In_1471,In_65);
nor U1424 (N_1424,In_509,In_869);
nor U1425 (N_1425,In_1599,In_1728);
and U1426 (N_1426,In_158,In_1327);
and U1427 (N_1427,In_819,In_1479);
and U1428 (N_1428,In_1998,In_385);
nor U1429 (N_1429,In_1936,In_876);
or U1430 (N_1430,In_1432,In_1460);
and U1431 (N_1431,In_1280,In_585);
or U1432 (N_1432,In_298,In_1216);
and U1433 (N_1433,In_1384,In_953);
and U1434 (N_1434,In_1261,In_1076);
nor U1435 (N_1435,In_1376,In_358);
or U1436 (N_1436,In_37,In_689);
and U1437 (N_1437,In_1415,In_1693);
xnor U1438 (N_1438,In_734,In_1285);
or U1439 (N_1439,In_787,In_81);
nor U1440 (N_1440,In_439,In_1803);
and U1441 (N_1441,In_1959,In_1245);
nor U1442 (N_1442,In_1057,In_704);
nand U1443 (N_1443,In_1017,In_1634);
or U1444 (N_1444,In_1339,In_1709);
or U1445 (N_1445,In_35,In_530);
and U1446 (N_1446,In_871,In_181);
and U1447 (N_1447,In_173,In_1065);
or U1448 (N_1448,In_1255,In_1030);
or U1449 (N_1449,In_1329,In_825);
or U1450 (N_1450,In_571,In_1289);
or U1451 (N_1451,In_1353,In_1973);
nand U1452 (N_1452,In_1184,In_1844);
or U1453 (N_1453,In_242,In_115);
and U1454 (N_1454,In_1763,In_1307);
nor U1455 (N_1455,In_914,In_568);
nor U1456 (N_1456,In_1857,In_1096);
nor U1457 (N_1457,In_1311,In_1127);
nor U1458 (N_1458,In_431,In_277);
nand U1459 (N_1459,In_1135,In_1188);
nor U1460 (N_1460,In_1645,In_518);
nand U1461 (N_1461,In_1149,In_15);
xor U1462 (N_1462,In_335,In_1017);
or U1463 (N_1463,In_1382,In_620);
and U1464 (N_1464,In_1758,In_1127);
or U1465 (N_1465,In_1995,In_1072);
nand U1466 (N_1466,In_815,In_1367);
nor U1467 (N_1467,In_730,In_462);
or U1468 (N_1468,In_1801,In_220);
and U1469 (N_1469,In_16,In_237);
xnor U1470 (N_1470,In_1663,In_1375);
and U1471 (N_1471,In_1450,In_1464);
xor U1472 (N_1472,In_1799,In_1991);
nand U1473 (N_1473,In_1422,In_1881);
nand U1474 (N_1474,In_159,In_1335);
or U1475 (N_1475,In_418,In_1042);
nor U1476 (N_1476,In_623,In_1118);
xnor U1477 (N_1477,In_1279,In_1636);
or U1478 (N_1478,In_869,In_1872);
or U1479 (N_1479,In_601,In_1123);
or U1480 (N_1480,In_1887,In_1535);
xor U1481 (N_1481,In_295,In_908);
nand U1482 (N_1482,In_349,In_1010);
nand U1483 (N_1483,In_705,In_38);
nand U1484 (N_1484,In_1215,In_768);
nor U1485 (N_1485,In_1527,In_157);
nor U1486 (N_1486,In_655,In_256);
nor U1487 (N_1487,In_997,In_901);
and U1488 (N_1488,In_526,In_1685);
or U1489 (N_1489,In_1349,In_972);
xor U1490 (N_1490,In_84,In_478);
xnor U1491 (N_1491,In_1433,In_545);
nand U1492 (N_1492,In_1660,In_1050);
nand U1493 (N_1493,In_844,In_1343);
nor U1494 (N_1494,In_273,In_1087);
or U1495 (N_1495,In_178,In_1212);
and U1496 (N_1496,In_54,In_832);
xor U1497 (N_1497,In_447,In_1461);
xnor U1498 (N_1498,In_1839,In_1999);
or U1499 (N_1499,In_1109,In_368);
xnor U1500 (N_1500,In_173,In_1693);
nor U1501 (N_1501,In_304,In_156);
or U1502 (N_1502,In_1533,In_1920);
xor U1503 (N_1503,In_370,In_1535);
and U1504 (N_1504,In_1682,In_282);
nor U1505 (N_1505,In_1528,In_1841);
or U1506 (N_1506,In_108,In_1770);
nand U1507 (N_1507,In_845,In_687);
nor U1508 (N_1508,In_1305,In_1556);
nand U1509 (N_1509,In_1929,In_406);
nor U1510 (N_1510,In_1592,In_700);
nor U1511 (N_1511,In_346,In_1445);
or U1512 (N_1512,In_1693,In_769);
nand U1513 (N_1513,In_186,In_982);
nor U1514 (N_1514,In_957,In_317);
and U1515 (N_1515,In_792,In_1982);
or U1516 (N_1516,In_300,In_1262);
or U1517 (N_1517,In_462,In_1763);
xor U1518 (N_1518,In_111,In_741);
or U1519 (N_1519,In_6,In_991);
or U1520 (N_1520,In_1506,In_1021);
and U1521 (N_1521,In_1239,In_1747);
xnor U1522 (N_1522,In_1825,In_1611);
xnor U1523 (N_1523,In_1110,In_277);
and U1524 (N_1524,In_1488,In_1744);
xor U1525 (N_1525,In_1138,In_134);
nor U1526 (N_1526,In_1168,In_1304);
nand U1527 (N_1527,In_1459,In_1680);
or U1528 (N_1528,In_614,In_845);
nor U1529 (N_1529,In_152,In_687);
nand U1530 (N_1530,In_66,In_39);
or U1531 (N_1531,In_1134,In_1602);
and U1532 (N_1532,In_171,In_936);
xor U1533 (N_1533,In_445,In_1484);
nand U1534 (N_1534,In_75,In_37);
or U1535 (N_1535,In_1419,In_1104);
nor U1536 (N_1536,In_1040,In_1114);
nand U1537 (N_1537,In_56,In_1835);
nor U1538 (N_1538,In_229,In_1049);
or U1539 (N_1539,In_944,In_1472);
and U1540 (N_1540,In_1879,In_1270);
nor U1541 (N_1541,In_231,In_820);
or U1542 (N_1542,In_970,In_1904);
xor U1543 (N_1543,In_566,In_131);
or U1544 (N_1544,In_1398,In_1080);
nor U1545 (N_1545,In_383,In_1368);
xnor U1546 (N_1546,In_323,In_1604);
and U1547 (N_1547,In_965,In_629);
or U1548 (N_1548,In_667,In_123);
or U1549 (N_1549,In_670,In_1352);
or U1550 (N_1550,In_680,In_1583);
nor U1551 (N_1551,In_797,In_67);
nand U1552 (N_1552,In_395,In_349);
or U1553 (N_1553,In_765,In_245);
nand U1554 (N_1554,In_847,In_1783);
nor U1555 (N_1555,In_1172,In_1059);
or U1556 (N_1556,In_1018,In_255);
nor U1557 (N_1557,In_1007,In_1001);
or U1558 (N_1558,In_1383,In_900);
nand U1559 (N_1559,In_784,In_109);
nand U1560 (N_1560,In_546,In_415);
nand U1561 (N_1561,In_1370,In_657);
or U1562 (N_1562,In_305,In_1921);
nor U1563 (N_1563,In_1130,In_367);
or U1564 (N_1564,In_1489,In_982);
nor U1565 (N_1565,In_1266,In_6);
nor U1566 (N_1566,In_1281,In_1878);
or U1567 (N_1567,In_1292,In_119);
nor U1568 (N_1568,In_359,In_737);
nor U1569 (N_1569,In_1160,In_941);
nand U1570 (N_1570,In_1763,In_545);
nor U1571 (N_1571,In_1474,In_570);
and U1572 (N_1572,In_409,In_1995);
xnor U1573 (N_1573,In_1176,In_1440);
nand U1574 (N_1574,In_768,In_629);
or U1575 (N_1575,In_1257,In_1792);
or U1576 (N_1576,In_1907,In_442);
xor U1577 (N_1577,In_381,In_1389);
nand U1578 (N_1578,In_1318,In_1709);
nand U1579 (N_1579,In_1875,In_812);
nand U1580 (N_1580,In_1114,In_82);
and U1581 (N_1581,In_1152,In_1076);
or U1582 (N_1582,In_1739,In_15);
nor U1583 (N_1583,In_1790,In_694);
nand U1584 (N_1584,In_242,In_1219);
xnor U1585 (N_1585,In_1368,In_485);
nor U1586 (N_1586,In_1969,In_738);
and U1587 (N_1587,In_1258,In_1814);
or U1588 (N_1588,In_853,In_437);
and U1589 (N_1589,In_1792,In_634);
xor U1590 (N_1590,In_1369,In_738);
nand U1591 (N_1591,In_961,In_267);
nor U1592 (N_1592,In_1190,In_758);
xnor U1593 (N_1593,In_353,In_1466);
or U1594 (N_1594,In_1297,In_565);
or U1595 (N_1595,In_678,In_277);
xnor U1596 (N_1596,In_1323,In_1474);
xnor U1597 (N_1597,In_1202,In_1773);
xor U1598 (N_1598,In_593,In_1487);
and U1599 (N_1599,In_1015,In_1344);
or U1600 (N_1600,In_1777,In_1773);
nor U1601 (N_1601,In_895,In_874);
or U1602 (N_1602,In_854,In_590);
nor U1603 (N_1603,In_1413,In_1954);
or U1604 (N_1604,In_1277,In_1106);
and U1605 (N_1605,In_119,In_1796);
and U1606 (N_1606,In_1163,In_122);
or U1607 (N_1607,In_1416,In_62);
or U1608 (N_1608,In_1774,In_199);
or U1609 (N_1609,In_1395,In_1044);
or U1610 (N_1610,In_1019,In_1015);
nand U1611 (N_1611,In_1180,In_579);
xor U1612 (N_1612,In_1797,In_471);
nand U1613 (N_1613,In_790,In_542);
nand U1614 (N_1614,In_50,In_1654);
nor U1615 (N_1615,In_1796,In_1986);
nand U1616 (N_1616,In_131,In_521);
and U1617 (N_1617,In_1686,In_124);
and U1618 (N_1618,In_1919,In_1840);
and U1619 (N_1619,In_144,In_422);
and U1620 (N_1620,In_882,In_1559);
or U1621 (N_1621,In_1308,In_427);
and U1622 (N_1622,In_1498,In_974);
nor U1623 (N_1623,In_1042,In_1231);
and U1624 (N_1624,In_946,In_1647);
nand U1625 (N_1625,In_1458,In_687);
nand U1626 (N_1626,In_194,In_772);
nand U1627 (N_1627,In_442,In_865);
nand U1628 (N_1628,In_180,In_336);
nand U1629 (N_1629,In_826,In_261);
and U1630 (N_1630,In_458,In_1526);
nand U1631 (N_1631,In_1854,In_468);
nand U1632 (N_1632,In_1409,In_51);
nor U1633 (N_1633,In_1817,In_1770);
nor U1634 (N_1634,In_375,In_1615);
nor U1635 (N_1635,In_1046,In_1680);
and U1636 (N_1636,In_392,In_1157);
nand U1637 (N_1637,In_526,In_690);
nand U1638 (N_1638,In_220,In_1565);
nand U1639 (N_1639,In_642,In_88);
nor U1640 (N_1640,In_1516,In_1427);
and U1641 (N_1641,In_1334,In_197);
and U1642 (N_1642,In_803,In_8);
and U1643 (N_1643,In_839,In_941);
nor U1644 (N_1644,In_246,In_1736);
nand U1645 (N_1645,In_536,In_762);
and U1646 (N_1646,In_1264,In_1037);
nand U1647 (N_1647,In_1816,In_1132);
nor U1648 (N_1648,In_44,In_360);
or U1649 (N_1649,In_197,In_451);
or U1650 (N_1650,In_307,In_1321);
nand U1651 (N_1651,In_1427,In_648);
and U1652 (N_1652,In_938,In_1966);
and U1653 (N_1653,In_679,In_947);
nor U1654 (N_1654,In_1055,In_1929);
or U1655 (N_1655,In_259,In_1142);
nor U1656 (N_1656,In_153,In_270);
and U1657 (N_1657,In_1343,In_1710);
and U1658 (N_1658,In_1172,In_225);
xnor U1659 (N_1659,In_1061,In_1789);
nor U1660 (N_1660,In_456,In_679);
nor U1661 (N_1661,In_1658,In_1036);
or U1662 (N_1662,In_864,In_635);
nand U1663 (N_1663,In_1010,In_1437);
xor U1664 (N_1664,In_1559,In_275);
or U1665 (N_1665,In_1102,In_1601);
or U1666 (N_1666,In_1283,In_1717);
nor U1667 (N_1667,In_63,In_1492);
nor U1668 (N_1668,In_505,In_1527);
and U1669 (N_1669,In_875,In_1958);
nand U1670 (N_1670,In_1064,In_839);
and U1671 (N_1671,In_1292,In_1218);
nor U1672 (N_1672,In_1350,In_269);
nor U1673 (N_1673,In_872,In_1469);
xnor U1674 (N_1674,In_1470,In_116);
nand U1675 (N_1675,In_1965,In_1831);
xnor U1676 (N_1676,In_1854,In_909);
or U1677 (N_1677,In_550,In_1983);
and U1678 (N_1678,In_1512,In_600);
or U1679 (N_1679,In_152,In_993);
nor U1680 (N_1680,In_1626,In_911);
nand U1681 (N_1681,In_1301,In_746);
nor U1682 (N_1682,In_102,In_1221);
nor U1683 (N_1683,In_674,In_864);
and U1684 (N_1684,In_1130,In_1805);
and U1685 (N_1685,In_461,In_598);
xnor U1686 (N_1686,In_70,In_340);
xor U1687 (N_1687,In_449,In_1385);
nor U1688 (N_1688,In_543,In_1783);
nand U1689 (N_1689,In_238,In_1423);
nor U1690 (N_1690,In_1568,In_461);
and U1691 (N_1691,In_474,In_1828);
xnor U1692 (N_1692,In_182,In_208);
or U1693 (N_1693,In_1021,In_1265);
nor U1694 (N_1694,In_852,In_1108);
nor U1695 (N_1695,In_1563,In_811);
nand U1696 (N_1696,In_1362,In_185);
or U1697 (N_1697,In_581,In_661);
nand U1698 (N_1698,In_1005,In_1433);
and U1699 (N_1699,In_911,In_840);
or U1700 (N_1700,In_882,In_1390);
and U1701 (N_1701,In_1305,In_756);
and U1702 (N_1702,In_1670,In_1339);
and U1703 (N_1703,In_543,In_1770);
nor U1704 (N_1704,In_756,In_201);
and U1705 (N_1705,In_667,In_862);
nand U1706 (N_1706,In_1470,In_1618);
and U1707 (N_1707,In_1643,In_393);
and U1708 (N_1708,In_874,In_1809);
and U1709 (N_1709,In_1112,In_1974);
or U1710 (N_1710,In_1668,In_1299);
and U1711 (N_1711,In_1070,In_424);
nand U1712 (N_1712,In_1561,In_1971);
nand U1713 (N_1713,In_1402,In_1398);
or U1714 (N_1714,In_466,In_439);
nand U1715 (N_1715,In_1909,In_418);
nand U1716 (N_1716,In_1913,In_856);
nor U1717 (N_1717,In_1964,In_15);
and U1718 (N_1718,In_634,In_58);
nand U1719 (N_1719,In_576,In_48);
nand U1720 (N_1720,In_1029,In_857);
xnor U1721 (N_1721,In_569,In_1526);
nor U1722 (N_1722,In_1380,In_1147);
or U1723 (N_1723,In_1313,In_804);
or U1724 (N_1724,In_1517,In_646);
or U1725 (N_1725,In_1970,In_815);
or U1726 (N_1726,In_1105,In_1921);
nand U1727 (N_1727,In_1303,In_1326);
nand U1728 (N_1728,In_1362,In_14);
xnor U1729 (N_1729,In_235,In_997);
nand U1730 (N_1730,In_1150,In_648);
nand U1731 (N_1731,In_761,In_1851);
and U1732 (N_1732,In_607,In_1849);
and U1733 (N_1733,In_916,In_1736);
and U1734 (N_1734,In_1036,In_1980);
nor U1735 (N_1735,In_1978,In_1274);
nor U1736 (N_1736,In_755,In_1220);
nand U1737 (N_1737,In_1478,In_1965);
and U1738 (N_1738,In_1671,In_1676);
and U1739 (N_1739,In_1164,In_1557);
or U1740 (N_1740,In_1056,In_897);
or U1741 (N_1741,In_495,In_597);
or U1742 (N_1742,In_1807,In_610);
nand U1743 (N_1743,In_687,In_344);
xnor U1744 (N_1744,In_623,In_785);
and U1745 (N_1745,In_1082,In_1338);
xor U1746 (N_1746,In_1217,In_525);
and U1747 (N_1747,In_1349,In_513);
or U1748 (N_1748,In_1039,In_1004);
or U1749 (N_1749,In_1071,In_219);
and U1750 (N_1750,In_1629,In_1576);
nand U1751 (N_1751,In_332,In_147);
and U1752 (N_1752,In_880,In_1707);
nand U1753 (N_1753,In_1873,In_383);
or U1754 (N_1754,In_490,In_25);
xor U1755 (N_1755,In_1088,In_897);
nand U1756 (N_1756,In_1934,In_1801);
and U1757 (N_1757,In_1924,In_1365);
nand U1758 (N_1758,In_303,In_919);
nor U1759 (N_1759,In_109,In_150);
nand U1760 (N_1760,In_346,In_396);
nor U1761 (N_1761,In_1817,In_1593);
and U1762 (N_1762,In_1408,In_1074);
xnor U1763 (N_1763,In_1863,In_1705);
and U1764 (N_1764,In_1644,In_1022);
nand U1765 (N_1765,In_81,In_1510);
nand U1766 (N_1766,In_901,In_218);
or U1767 (N_1767,In_171,In_439);
nand U1768 (N_1768,In_1720,In_1025);
or U1769 (N_1769,In_919,In_704);
and U1770 (N_1770,In_1100,In_1045);
and U1771 (N_1771,In_210,In_929);
nand U1772 (N_1772,In_1626,In_454);
nor U1773 (N_1773,In_596,In_1783);
and U1774 (N_1774,In_149,In_1765);
xnor U1775 (N_1775,In_879,In_236);
nand U1776 (N_1776,In_1345,In_34);
nand U1777 (N_1777,In_188,In_1419);
nor U1778 (N_1778,In_665,In_1409);
and U1779 (N_1779,In_210,In_1309);
nor U1780 (N_1780,In_165,In_1155);
xnor U1781 (N_1781,In_55,In_1179);
nor U1782 (N_1782,In_1283,In_795);
nand U1783 (N_1783,In_810,In_1244);
xnor U1784 (N_1784,In_202,In_1260);
or U1785 (N_1785,In_718,In_545);
or U1786 (N_1786,In_320,In_943);
or U1787 (N_1787,In_323,In_1831);
or U1788 (N_1788,In_1531,In_652);
or U1789 (N_1789,In_1783,In_538);
nand U1790 (N_1790,In_878,In_1577);
and U1791 (N_1791,In_1265,In_120);
and U1792 (N_1792,In_1307,In_930);
or U1793 (N_1793,In_943,In_29);
xor U1794 (N_1794,In_1630,In_25);
nor U1795 (N_1795,In_1309,In_791);
nand U1796 (N_1796,In_1847,In_598);
and U1797 (N_1797,In_842,In_378);
and U1798 (N_1798,In_1445,In_1696);
or U1799 (N_1799,In_49,In_305);
and U1800 (N_1800,In_880,In_1580);
nor U1801 (N_1801,In_78,In_102);
and U1802 (N_1802,In_964,In_1456);
nand U1803 (N_1803,In_1677,In_1243);
xnor U1804 (N_1804,In_1836,In_1046);
and U1805 (N_1805,In_1146,In_1281);
nor U1806 (N_1806,In_606,In_1637);
or U1807 (N_1807,In_1089,In_961);
or U1808 (N_1808,In_230,In_650);
xnor U1809 (N_1809,In_1356,In_275);
nor U1810 (N_1810,In_1376,In_1173);
xnor U1811 (N_1811,In_1158,In_1594);
and U1812 (N_1812,In_370,In_1510);
xnor U1813 (N_1813,In_314,In_937);
or U1814 (N_1814,In_209,In_1659);
nand U1815 (N_1815,In_474,In_576);
nand U1816 (N_1816,In_1634,In_1599);
xnor U1817 (N_1817,In_803,In_956);
or U1818 (N_1818,In_342,In_1340);
and U1819 (N_1819,In_1196,In_904);
or U1820 (N_1820,In_707,In_64);
xor U1821 (N_1821,In_866,In_120);
xor U1822 (N_1822,In_993,In_1730);
nand U1823 (N_1823,In_1284,In_528);
nand U1824 (N_1824,In_736,In_857);
nor U1825 (N_1825,In_1974,In_1219);
or U1826 (N_1826,In_295,In_1377);
nor U1827 (N_1827,In_635,In_248);
or U1828 (N_1828,In_1591,In_1929);
or U1829 (N_1829,In_28,In_1722);
nand U1830 (N_1830,In_1319,In_711);
xnor U1831 (N_1831,In_722,In_1768);
or U1832 (N_1832,In_1305,In_761);
xor U1833 (N_1833,In_264,In_676);
or U1834 (N_1834,In_898,In_72);
xor U1835 (N_1835,In_125,In_5);
xnor U1836 (N_1836,In_1965,In_1334);
nand U1837 (N_1837,In_1993,In_339);
nor U1838 (N_1838,In_734,In_721);
xnor U1839 (N_1839,In_116,In_226);
and U1840 (N_1840,In_578,In_1860);
xnor U1841 (N_1841,In_175,In_1167);
and U1842 (N_1842,In_1331,In_1865);
or U1843 (N_1843,In_1400,In_1459);
nand U1844 (N_1844,In_1840,In_1991);
and U1845 (N_1845,In_206,In_1136);
nand U1846 (N_1846,In_350,In_1883);
and U1847 (N_1847,In_864,In_1541);
or U1848 (N_1848,In_1947,In_1745);
or U1849 (N_1849,In_752,In_1628);
nor U1850 (N_1850,In_449,In_1558);
and U1851 (N_1851,In_1559,In_89);
nor U1852 (N_1852,In_1439,In_441);
nand U1853 (N_1853,In_676,In_398);
nand U1854 (N_1854,In_411,In_165);
and U1855 (N_1855,In_1994,In_546);
nor U1856 (N_1856,In_1053,In_1771);
nor U1857 (N_1857,In_1495,In_1815);
or U1858 (N_1858,In_1508,In_303);
and U1859 (N_1859,In_588,In_1915);
nor U1860 (N_1860,In_983,In_1664);
nand U1861 (N_1861,In_490,In_1782);
and U1862 (N_1862,In_1421,In_1941);
nand U1863 (N_1863,In_703,In_1776);
nor U1864 (N_1864,In_126,In_991);
nand U1865 (N_1865,In_282,In_815);
nor U1866 (N_1866,In_1124,In_998);
nor U1867 (N_1867,In_240,In_1127);
nor U1868 (N_1868,In_1203,In_347);
nor U1869 (N_1869,In_861,In_1949);
or U1870 (N_1870,In_1274,In_549);
or U1871 (N_1871,In_219,In_439);
xor U1872 (N_1872,In_730,In_1589);
xor U1873 (N_1873,In_1745,In_1830);
or U1874 (N_1874,In_1976,In_412);
nor U1875 (N_1875,In_1282,In_274);
or U1876 (N_1876,In_487,In_667);
nand U1877 (N_1877,In_1355,In_128);
nor U1878 (N_1878,In_160,In_1030);
nor U1879 (N_1879,In_495,In_425);
nand U1880 (N_1880,In_1709,In_1026);
nand U1881 (N_1881,In_355,In_1477);
nor U1882 (N_1882,In_1513,In_702);
nand U1883 (N_1883,In_1154,In_98);
and U1884 (N_1884,In_259,In_951);
or U1885 (N_1885,In_161,In_6);
and U1886 (N_1886,In_242,In_1824);
and U1887 (N_1887,In_6,In_105);
nand U1888 (N_1888,In_1143,In_1846);
and U1889 (N_1889,In_255,In_810);
or U1890 (N_1890,In_1753,In_1434);
xnor U1891 (N_1891,In_1476,In_486);
nor U1892 (N_1892,In_447,In_1341);
or U1893 (N_1893,In_221,In_1624);
nand U1894 (N_1894,In_1695,In_1637);
and U1895 (N_1895,In_1134,In_1027);
or U1896 (N_1896,In_795,In_622);
xnor U1897 (N_1897,In_1658,In_389);
nor U1898 (N_1898,In_1911,In_1421);
nand U1899 (N_1899,In_265,In_350);
nand U1900 (N_1900,In_1400,In_1814);
xor U1901 (N_1901,In_1257,In_699);
or U1902 (N_1902,In_632,In_707);
and U1903 (N_1903,In_549,In_284);
and U1904 (N_1904,In_94,In_360);
and U1905 (N_1905,In_362,In_1748);
nor U1906 (N_1906,In_772,In_1150);
and U1907 (N_1907,In_610,In_806);
nand U1908 (N_1908,In_494,In_1798);
nand U1909 (N_1909,In_1230,In_1550);
and U1910 (N_1910,In_1898,In_1216);
nor U1911 (N_1911,In_490,In_1335);
nand U1912 (N_1912,In_191,In_1405);
nor U1913 (N_1913,In_1166,In_547);
xnor U1914 (N_1914,In_1916,In_564);
xnor U1915 (N_1915,In_1654,In_1082);
xnor U1916 (N_1916,In_914,In_1740);
nor U1917 (N_1917,In_1045,In_1601);
nor U1918 (N_1918,In_744,In_1398);
and U1919 (N_1919,In_543,In_1444);
and U1920 (N_1920,In_1293,In_1846);
and U1921 (N_1921,In_351,In_399);
nand U1922 (N_1922,In_45,In_260);
or U1923 (N_1923,In_1004,In_1985);
xor U1924 (N_1924,In_834,In_645);
xor U1925 (N_1925,In_222,In_1101);
and U1926 (N_1926,In_1849,In_1835);
or U1927 (N_1927,In_1854,In_1634);
nand U1928 (N_1928,In_449,In_416);
nand U1929 (N_1929,In_1140,In_1585);
nand U1930 (N_1930,In_574,In_1350);
nand U1931 (N_1931,In_608,In_736);
and U1932 (N_1932,In_214,In_1602);
and U1933 (N_1933,In_604,In_843);
nor U1934 (N_1934,In_1171,In_1680);
nand U1935 (N_1935,In_918,In_940);
nand U1936 (N_1936,In_1631,In_1297);
nand U1937 (N_1937,In_1557,In_1395);
or U1938 (N_1938,In_1880,In_1352);
nand U1939 (N_1939,In_1582,In_678);
or U1940 (N_1940,In_967,In_1699);
xor U1941 (N_1941,In_1892,In_731);
and U1942 (N_1942,In_349,In_1821);
or U1943 (N_1943,In_812,In_1771);
and U1944 (N_1944,In_916,In_140);
and U1945 (N_1945,In_284,In_1982);
or U1946 (N_1946,In_971,In_1197);
nand U1947 (N_1947,In_1953,In_1957);
nand U1948 (N_1948,In_467,In_1159);
nor U1949 (N_1949,In_970,In_938);
or U1950 (N_1950,In_944,In_1747);
nand U1951 (N_1951,In_1482,In_1760);
nand U1952 (N_1952,In_224,In_957);
and U1953 (N_1953,In_1521,In_1746);
and U1954 (N_1954,In_828,In_544);
nor U1955 (N_1955,In_242,In_52);
and U1956 (N_1956,In_1547,In_1262);
nand U1957 (N_1957,In_1680,In_61);
nor U1958 (N_1958,In_1993,In_1397);
or U1959 (N_1959,In_1689,In_144);
nor U1960 (N_1960,In_1827,In_1647);
nor U1961 (N_1961,In_582,In_438);
nand U1962 (N_1962,In_1699,In_1885);
nand U1963 (N_1963,In_1312,In_1216);
nand U1964 (N_1964,In_1367,In_1900);
or U1965 (N_1965,In_1134,In_1313);
xor U1966 (N_1966,In_1395,In_545);
nor U1967 (N_1967,In_1552,In_391);
xnor U1968 (N_1968,In_1485,In_52);
xor U1969 (N_1969,In_243,In_1693);
nand U1970 (N_1970,In_492,In_1567);
nand U1971 (N_1971,In_1377,In_358);
nand U1972 (N_1972,In_245,In_1229);
nand U1973 (N_1973,In_627,In_352);
or U1974 (N_1974,In_939,In_509);
xnor U1975 (N_1975,In_1031,In_1734);
nand U1976 (N_1976,In_1932,In_655);
or U1977 (N_1977,In_1759,In_1117);
nor U1978 (N_1978,In_443,In_1103);
and U1979 (N_1979,In_545,In_1759);
xor U1980 (N_1980,In_1613,In_151);
and U1981 (N_1981,In_1411,In_1690);
nor U1982 (N_1982,In_1968,In_888);
nor U1983 (N_1983,In_868,In_708);
nor U1984 (N_1984,In_590,In_249);
xor U1985 (N_1985,In_1705,In_491);
nor U1986 (N_1986,In_427,In_971);
and U1987 (N_1987,In_1132,In_535);
or U1988 (N_1988,In_340,In_159);
xnor U1989 (N_1989,In_378,In_444);
and U1990 (N_1990,In_192,In_858);
nor U1991 (N_1991,In_1859,In_1608);
or U1992 (N_1992,In_61,In_1386);
nor U1993 (N_1993,In_1393,In_365);
and U1994 (N_1994,In_292,In_137);
or U1995 (N_1995,In_503,In_475);
nor U1996 (N_1996,In_811,In_1337);
nor U1997 (N_1997,In_307,In_1695);
or U1998 (N_1998,In_1796,In_1423);
or U1999 (N_1999,In_1732,In_1530);
or U2000 (N_2000,N_1400,N_1878);
nand U2001 (N_2001,N_1782,N_139);
nand U2002 (N_2002,N_1234,N_677);
or U2003 (N_2003,N_976,N_1806);
or U2004 (N_2004,N_701,N_1100);
nand U2005 (N_2005,N_1921,N_913);
nand U2006 (N_2006,N_1999,N_1395);
nor U2007 (N_2007,N_1777,N_1338);
or U2008 (N_2008,N_972,N_1841);
xor U2009 (N_2009,N_1232,N_1358);
and U2010 (N_2010,N_1656,N_1866);
xor U2011 (N_2011,N_1821,N_339);
and U2012 (N_2012,N_504,N_719);
nor U2013 (N_2013,N_1096,N_1886);
nand U2014 (N_2014,N_1910,N_830);
or U2015 (N_2015,N_163,N_200);
xnor U2016 (N_2016,N_818,N_410);
nor U2017 (N_2017,N_458,N_375);
nand U2018 (N_2018,N_693,N_1581);
and U2019 (N_2019,N_977,N_1000);
and U2020 (N_2020,N_1922,N_1290);
or U2021 (N_2021,N_166,N_1480);
nor U2022 (N_2022,N_1090,N_1650);
nor U2023 (N_2023,N_270,N_153);
nor U2024 (N_2024,N_577,N_679);
or U2025 (N_2025,N_545,N_459);
xnor U2026 (N_2026,N_204,N_1964);
nor U2027 (N_2027,N_1768,N_58);
nand U2028 (N_2028,N_1792,N_1304);
nor U2029 (N_2029,N_1692,N_801);
or U2030 (N_2030,N_1439,N_670);
nor U2031 (N_2031,N_543,N_919);
or U2032 (N_2032,N_1824,N_1775);
nand U2033 (N_2033,N_1823,N_1546);
nor U2034 (N_2034,N_338,N_5);
nor U2035 (N_2035,N_1278,N_1276);
or U2036 (N_2036,N_1231,N_42);
nand U2037 (N_2037,N_198,N_579);
or U2038 (N_2038,N_321,N_615);
or U2039 (N_2039,N_1671,N_1519);
xnor U2040 (N_2040,N_1206,N_825);
or U2041 (N_2041,N_308,N_1780);
xnor U2042 (N_2042,N_1805,N_887);
nand U2043 (N_2043,N_981,N_1509);
or U2044 (N_2044,N_186,N_666);
xor U2045 (N_2045,N_790,N_609);
or U2046 (N_2046,N_1596,N_691);
nor U2047 (N_2047,N_39,N_625);
nand U2048 (N_2048,N_1004,N_1958);
and U2049 (N_2049,N_1372,N_189);
nand U2050 (N_2050,N_1109,N_792);
nor U2051 (N_2051,N_1474,N_353);
nand U2052 (N_2052,N_1376,N_512);
nor U2053 (N_2053,N_728,N_1467);
nand U2054 (N_2054,N_1407,N_448);
nand U2055 (N_2055,N_1471,N_1737);
nand U2056 (N_2056,N_982,N_92);
and U2057 (N_2057,N_1210,N_909);
and U2058 (N_2058,N_1040,N_262);
nand U2059 (N_2059,N_1417,N_494);
and U2060 (N_2060,N_1747,N_1923);
nor U2061 (N_2061,N_1184,N_793);
and U2062 (N_2062,N_1944,N_1660);
or U2063 (N_2063,N_1038,N_869);
and U2064 (N_2064,N_242,N_740);
nand U2065 (N_2065,N_6,N_889);
and U2066 (N_2066,N_829,N_1077);
and U2067 (N_2067,N_925,N_638);
or U2068 (N_2068,N_1148,N_1788);
or U2069 (N_2069,N_523,N_1243);
or U2070 (N_2070,N_271,N_1366);
or U2071 (N_2071,N_1716,N_574);
or U2072 (N_2072,N_483,N_462);
and U2073 (N_2073,N_383,N_9);
nand U2074 (N_2074,N_1666,N_155);
and U2075 (N_2075,N_1079,N_469);
and U2076 (N_2076,N_115,N_752);
nor U2077 (N_2077,N_687,N_108);
or U2078 (N_2078,N_1024,N_1108);
nand U2079 (N_2079,N_1569,N_1473);
xor U2080 (N_2080,N_33,N_1204);
and U2081 (N_2081,N_1507,N_1504);
xnor U2082 (N_2082,N_1355,N_152);
or U2083 (N_2083,N_1379,N_589);
nand U2084 (N_2084,N_284,N_559);
nor U2085 (N_2085,N_1979,N_429);
or U2086 (N_2086,N_1734,N_1216);
xor U2087 (N_2087,N_965,N_1237);
or U2088 (N_2088,N_1350,N_944);
or U2089 (N_2089,N_630,N_1811);
or U2090 (N_2090,N_1085,N_767);
and U2091 (N_2091,N_1399,N_88);
and U2092 (N_2092,N_1689,N_934);
nand U2093 (N_2093,N_46,N_1430);
or U2094 (N_2094,N_17,N_888);
nor U2095 (N_2095,N_309,N_403);
nand U2096 (N_2096,N_1822,N_629);
and U2097 (N_2097,N_1270,N_1104);
and U2098 (N_2098,N_116,N_287);
nand U2099 (N_2099,N_717,N_59);
or U2100 (N_2100,N_1492,N_1076);
nand U2101 (N_2101,N_1817,N_835);
and U2102 (N_2102,N_521,N_1906);
and U2103 (N_2103,N_1297,N_297);
nand U2104 (N_2104,N_1371,N_503);
nand U2105 (N_2105,N_351,N_1037);
and U2106 (N_2106,N_1592,N_1807);
nor U2107 (N_2107,N_1868,N_1753);
xnor U2108 (N_2108,N_335,N_1629);
and U2109 (N_2109,N_1043,N_1075);
nand U2110 (N_2110,N_884,N_1559);
or U2111 (N_2111,N_1778,N_566);
and U2112 (N_2112,N_1696,N_864);
nand U2113 (N_2113,N_1580,N_26);
or U2114 (N_2114,N_385,N_60);
nor U2115 (N_2115,N_648,N_724);
or U2116 (N_2116,N_959,N_182);
or U2117 (N_2117,N_1847,N_237);
or U2118 (N_2118,N_506,N_768);
nor U2119 (N_2119,N_703,N_1706);
and U2120 (N_2120,N_1762,N_998);
or U2121 (N_2121,N_813,N_1042);
and U2122 (N_2122,N_70,N_553);
nor U2123 (N_2123,N_1437,N_450);
nor U2124 (N_2124,N_1050,N_1987);
nand U2125 (N_2125,N_190,N_267);
nand U2126 (N_2126,N_1320,N_211);
or U2127 (N_2127,N_427,N_1908);
and U2128 (N_2128,N_1203,N_1272);
and U2129 (N_2129,N_1251,N_1902);
nand U2130 (N_2130,N_1134,N_1387);
nor U2131 (N_2131,N_1449,N_285);
and U2132 (N_2132,N_1548,N_1292);
nor U2133 (N_2133,N_248,N_149);
nand U2134 (N_2134,N_1489,N_336);
and U2135 (N_2135,N_1324,N_1208);
nor U2136 (N_2136,N_45,N_244);
nor U2137 (N_2137,N_519,N_973);
nand U2138 (N_2138,N_1432,N_72);
nor U2139 (N_2139,N_305,N_537);
nor U2140 (N_2140,N_1725,N_1728);
and U2141 (N_2141,N_1609,N_402);
or U2142 (N_2142,N_866,N_774);
and U2143 (N_2143,N_808,N_834);
nor U2144 (N_2144,N_809,N_632);
nand U2145 (N_2145,N_1053,N_389);
and U2146 (N_2146,N_1026,N_1326);
or U2147 (N_2147,N_228,N_302);
or U2148 (N_2148,N_1732,N_1284);
and U2149 (N_2149,N_358,N_949);
and U2150 (N_2150,N_507,N_1630);
or U2151 (N_2151,N_1651,N_897);
nand U2152 (N_2152,N_1832,N_764);
nor U2153 (N_2153,N_656,N_454);
xnor U2154 (N_2154,N_1286,N_1469);
or U2155 (N_2155,N_205,N_757);
or U2156 (N_2156,N_1460,N_644);
nand U2157 (N_2157,N_453,N_1887);
nor U2158 (N_2158,N_709,N_1834);
nor U2159 (N_2159,N_1563,N_1317);
and U2160 (N_2160,N_291,N_1645);
or U2161 (N_2161,N_990,N_995);
or U2162 (N_2162,N_1122,N_129);
nor U2163 (N_2163,N_931,N_730);
or U2164 (N_2164,N_1089,N_1901);
xnor U2165 (N_2165,N_23,N_343);
nand U2166 (N_2166,N_903,N_1176);
nor U2167 (N_2167,N_434,N_1566);
nand U2168 (N_2168,N_777,N_1200);
or U2169 (N_2169,N_127,N_1954);
or U2170 (N_2170,N_1647,N_422);
xnor U2171 (N_2171,N_256,N_1594);
or U2172 (N_2172,N_247,N_456);
nor U2173 (N_2173,N_775,N_63);
nor U2174 (N_2174,N_1328,N_664);
nand U2175 (N_2175,N_431,N_1720);
nor U2176 (N_2176,N_1508,N_1179);
or U2177 (N_2177,N_803,N_1045);
or U2178 (N_2178,N_1541,N_1533);
nand U2179 (N_2179,N_616,N_1194);
and U2180 (N_2180,N_804,N_858);
and U2181 (N_2181,N_1345,N_1325);
or U2182 (N_2182,N_999,N_821);
and U2183 (N_2183,N_1312,N_1107);
xnor U2184 (N_2184,N_1662,N_1105);
or U2185 (N_2185,N_1894,N_220);
nor U2186 (N_2186,N_1983,N_1828);
or U2187 (N_2187,N_178,N_570);
and U2188 (N_2188,N_432,N_1937);
nor U2189 (N_2189,N_334,N_86);
nand U2190 (N_2190,N_463,N_1146);
nand U2191 (N_2191,N_320,N_412);
nand U2192 (N_2192,N_1360,N_1313);
or U2193 (N_2193,N_1262,N_1362);
and U2194 (N_2194,N_327,N_706);
nand U2195 (N_2195,N_568,N_816);
and U2196 (N_2196,N_891,N_1061);
nor U2197 (N_2197,N_120,N_143);
nor U2198 (N_2198,N_1956,N_295);
nand U2199 (N_2199,N_1731,N_759);
and U2200 (N_2200,N_1468,N_544);
nor U2201 (N_2201,N_168,N_832);
or U2202 (N_2202,N_592,N_868);
and U2203 (N_2203,N_561,N_1938);
and U2204 (N_2204,N_1556,N_784);
xnor U2205 (N_2205,N_468,N_621);
nand U2206 (N_2206,N_489,N_1315);
nand U2207 (N_2207,N_109,N_1744);
and U2208 (N_2208,N_896,N_1282);
nor U2209 (N_2209,N_1438,N_1733);
nor U2210 (N_2210,N_1554,N_1907);
xnor U2211 (N_2211,N_1703,N_377);
nand U2212 (N_2212,N_1485,N_700);
nor U2213 (N_2213,N_94,N_1225);
or U2214 (N_2214,N_1205,N_647);
nand U2215 (N_2215,N_781,N_1642);
or U2216 (N_2216,N_435,N_760);
nor U2217 (N_2217,N_1535,N_927);
xnor U2218 (N_2218,N_48,N_179);
or U2219 (N_2219,N_1881,N_1751);
nand U2220 (N_2220,N_942,N_824);
or U2221 (N_2221,N_1565,N_1578);
nand U2222 (N_2222,N_350,N_333);
nand U2223 (N_2223,N_400,N_1403);
nor U2224 (N_2224,N_1771,N_1189);
xor U2225 (N_2225,N_352,N_837);
and U2226 (N_2226,N_1346,N_599);
nor U2227 (N_2227,N_895,N_1029);
nor U2228 (N_2228,N_1895,N_1941);
nand U2229 (N_2229,N_1041,N_1653);
and U2230 (N_2230,N_538,N_649);
or U2231 (N_2231,N_1606,N_1712);
and U2232 (N_2232,N_1008,N_1641);
and U2233 (N_2233,N_1446,N_1914);
nor U2234 (N_2234,N_37,N_645);
nand U2235 (N_2235,N_1248,N_1668);
or U2236 (N_2236,N_1856,N_201);
nand U2237 (N_2237,N_1572,N_484);
nand U2238 (N_2238,N_405,N_549);
and U2239 (N_2239,N_902,N_480);
and U2240 (N_2240,N_417,N_1974);
or U2241 (N_2241,N_1305,N_1143);
or U2242 (N_2242,N_967,N_1318);
or U2243 (N_2243,N_720,N_1212);
or U2244 (N_2244,N_683,N_732);
nand U2245 (N_2245,N_1110,N_373);
xnor U2246 (N_2246,N_240,N_1567);
xnor U2247 (N_2247,N_1961,N_388);
and U2248 (N_2248,N_38,N_1028);
nand U2249 (N_2249,N_1871,N_381);
and U2250 (N_2250,N_755,N_114);
nand U2251 (N_2251,N_1670,N_922);
nand U2252 (N_2252,N_257,N_745);
nand U2253 (N_2253,N_1831,N_328);
and U2254 (N_2254,N_430,N_340);
nor U2255 (N_2255,N_1537,N_1835);
and U2256 (N_2256,N_935,N_1685);
or U2257 (N_2257,N_1281,N_1560);
xor U2258 (N_2258,N_472,N_214);
nor U2259 (N_2259,N_1590,N_123);
or U2260 (N_2260,N_160,N_1269);
nand U2261 (N_2261,N_765,N_145);
and U2262 (N_2262,N_963,N_747);
or U2263 (N_2263,N_1975,N_122);
or U2264 (N_2264,N_1497,N_624);
nand U2265 (N_2265,N_1957,N_562);
nand U2266 (N_2266,N_289,N_565);
xnor U2267 (N_2267,N_1680,N_1499);
nor U2268 (N_2268,N_344,N_1215);
nand U2269 (N_2269,N_655,N_1101);
or U2270 (N_2270,N_1496,N_1260);
and U2271 (N_2271,N_319,N_1693);
nand U2272 (N_2272,N_1640,N_1800);
nand U2273 (N_2273,N_1551,N_1538);
nor U2274 (N_2274,N_1447,N_1681);
xnor U2275 (N_2275,N_1661,N_342);
and U2276 (N_2276,N_82,N_246);
nand U2277 (N_2277,N_95,N_234);
and U2278 (N_2278,N_174,N_1151);
and U2279 (N_2279,N_478,N_1749);
nor U2280 (N_2280,N_1611,N_1993);
nor U2281 (N_2281,N_660,N_32);
or U2282 (N_2282,N_1843,N_101);
and U2283 (N_2283,N_1764,N_1950);
and U2284 (N_2284,N_928,N_571);
nor U2285 (N_2285,N_726,N_1410);
nor U2286 (N_2286,N_1942,N_223);
xnor U2287 (N_2287,N_1664,N_1967);
nand U2288 (N_2288,N_1691,N_80);
nor U2289 (N_2289,N_159,N_67);
nor U2290 (N_2290,N_1391,N_1912);
nand U2291 (N_2291,N_1849,N_1013);
nor U2292 (N_2292,N_1465,N_266);
xor U2293 (N_2293,N_953,N_1652);
nor U2294 (N_2294,N_1099,N_419);
nand U2295 (N_2295,N_1406,N_1549);
nor U2296 (N_2296,N_477,N_1752);
or U2297 (N_2297,N_1054,N_1963);
and U2298 (N_2298,N_1339,N_1130);
and U2299 (N_2299,N_1699,N_1915);
or U2300 (N_2300,N_192,N_265);
xor U2301 (N_2301,N_508,N_1978);
nor U2302 (N_2302,N_1955,N_1126);
xnor U2303 (N_2303,N_1289,N_1718);
xor U2304 (N_2304,N_1758,N_886);
or U2305 (N_2305,N_161,N_1599);
nand U2306 (N_2306,N_1511,N_1619);
nand U2307 (N_2307,N_1991,N_197);
and U2308 (N_2308,N_511,N_1530);
nor U2309 (N_2309,N_355,N_1202);
nand U2310 (N_2310,N_294,N_1715);
nand U2311 (N_2311,N_641,N_1150);
xor U2312 (N_2312,N_1925,N_1268);
nand U2313 (N_2313,N_218,N_528);
xnor U2314 (N_2314,N_1389,N_1191);
and U2315 (N_2315,N_754,N_280);
nor U2316 (N_2316,N_778,N_698);
and U2317 (N_2317,N_1453,N_812);
nand U2318 (N_2318,N_104,N_1568);
nor U2319 (N_2319,N_310,N_731);
nand U2320 (N_2320,N_502,N_1616);
and U2321 (N_2321,N_1857,N_1327);
or U2322 (N_2322,N_1409,N_27);
nand U2323 (N_2323,N_1080,N_379);
or U2324 (N_2324,N_249,N_684);
nand U2325 (N_2325,N_1574,N_874);
nor U2326 (N_2326,N_1258,N_603);
nand U2327 (N_2327,N_1334,N_1673);
nand U2328 (N_2328,N_1125,N_1149);
nand U2329 (N_2329,N_1631,N_1302);
nand U2330 (N_2330,N_1951,N_1669);
nand U2331 (N_2331,N_1595,N_1682);
and U2332 (N_2332,N_954,N_1929);
and U2333 (N_2333,N_782,N_1707);
nand U2334 (N_2334,N_1860,N_1257);
or U2335 (N_2335,N_1676,N_1615);
nand U2336 (N_2336,N_50,N_1883);
and U2337 (N_2337,N_1396,N_1971);
and U2338 (N_2338,N_171,N_614);
nor U2339 (N_2339,N_685,N_1193);
or U2340 (N_2340,N_301,N_1074);
nand U2341 (N_2341,N_996,N_892);
nand U2342 (N_2342,N_1765,N_1117);
or U2343 (N_2343,N_1022,N_1);
or U2344 (N_2344,N_66,N_194);
nand U2345 (N_2345,N_465,N_1809);
xor U2346 (N_2346,N_1002,N_1375);
and U2347 (N_2347,N_1083,N_136);
and U2348 (N_2348,N_653,N_882);
or U2349 (N_2349,N_324,N_361);
nand U2350 (N_2350,N_1618,N_273);
and U2351 (N_2351,N_492,N_1009);
or U2352 (N_2352,N_1364,N_1341);
nand U2353 (N_2353,N_1036,N_1862);
xor U2354 (N_2354,N_15,N_497);
nand U2355 (N_2355,N_1639,N_1605);
and U2356 (N_2356,N_195,N_1917);
or U2357 (N_2357,N_1017,N_299);
nor U2358 (N_2358,N_1027,N_1532);
or U2359 (N_2359,N_1477,N_966);
nor U2360 (N_2360,N_1604,N_1602);
nand U2361 (N_2361,N_1158,N_1514);
nor U2362 (N_2362,N_167,N_1161);
xnor U2363 (N_2363,N_279,N_817);
or U2364 (N_2364,N_1267,N_370);
nor U2365 (N_2365,N_363,N_551);
nand U2366 (N_2366,N_844,N_1779);
and U2367 (N_2367,N_202,N_1246);
and U2368 (N_2368,N_1512,N_481);
nand U2369 (N_2369,N_586,N_1624);
and U2370 (N_2370,N_1990,N_245);
and U2371 (N_2371,N_1330,N_447);
nand U2372 (N_2372,N_1521,N_604);
nor U2373 (N_2373,N_1932,N_1542);
and U2374 (N_2374,N_1455,N_22);
nand U2375 (N_2375,N_548,N_1273);
nor U2376 (N_2376,N_1283,N_208);
nand U2377 (N_2377,N_1062,N_1309);
nor U2378 (N_2378,N_165,N_1388);
nor U2379 (N_2379,N_1724,N_1112);
or U2380 (N_2380,N_229,N_206);
and U2381 (N_2381,N_1393,N_3);
xnor U2382 (N_2382,N_725,N_323);
nor U2383 (N_2383,N_425,N_1935);
or U2384 (N_2384,N_1111,N_1429);
and U2385 (N_2385,N_611,N_1167);
and U2386 (N_2386,N_669,N_1363);
nor U2387 (N_2387,N_727,N_1254);
and U2388 (N_2388,N_1331,N_1046);
xnor U2389 (N_2389,N_744,N_1214);
and U2390 (N_2390,N_572,N_975);
and U2391 (N_2391,N_1280,N_322);
or U2392 (N_2392,N_786,N_1903);
nand U2393 (N_2393,N_1352,N_1977);
or U2394 (N_2394,N_1298,N_613);
and U2395 (N_2395,N_1960,N_177);
nor U2396 (N_2396,N_1175,N_1285);
nor U2397 (N_2397,N_1845,N_1256);
or U2398 (N_2398,N_1700,N_241);
nand U2399 (N_2399,N_1344,N_665);
or U2400 (N_2400,N_341,N_1222);
and U2401 (N_2401,N_138,N_1060);
or U2402 (N_2402,N_1230,N_1464);
nand U2403 (N_2403,N_451,N_332);
nor U2404 (N_2404,N_356,N_1381);
and U2405 (N_2405,N_1255,N_879);
and U2406 (N_2406,N_121,N_1742);
or U2407 (N_2407,N_1959,N_84);
or U2408 (N_2408,N_1168,N_455);
nand U2409 (N_2409,N_987,N_1939);
nor U2410 (N_2410,N_1882,N_1795);
xnor U2411 (N_2411,N_44,N_1217);
nor U2412 (N_2412,N_1995,N_117);
nor U2413 (N_2413,N_1431,N_739);
and U2414 (N_2414,N_540,N_618);
nand U2415 (N_2415,N_1648,N_147);
nor U2416 (N_2416,N_103,N_1701);
or U2417 (N_2417,N_146,N_1444);
and U2418 (N_2418,N_721,N_1359);
xor U2419 (N_2419,N_1249,N_1288);
nand U2420 (N_2420,N_516,N_1405);
nor U2421 (N_2421,N_737,N_991);
and U2422 (N_2422,N_1458,N_213);
xnor U2423 (N_2423,N_993,N_539);
or U2424 (N_2424,N_1677,N_1873);
xnor U2425 (N_2425,N_762,N_617);
or U2426 (N_2426,N_606,N_1638);
and U2427 (N_2427,N_800,N_681);
nor U2428 (N_2428,N_904,N_1840);
and U2429 (N_2429,N_1634,N_1242);
nand U2430 (N_2430,N_1688,N_1370);
xnor U2431 (N_2431,N_1520,N_1226);
or U2432 (N_2432,N_1383,N_102);
xor U2433 (N_2433,N_743,N_1142);
or U2434 (N_2434,N_1198,N_794);
or U2435 (N_2435,N_1501,N_1349);
nor U2436 (N_2436,N_21,N_1368);
nor U2437 (N_2437,N_1140,N_1710);
nor U2438 (N_2438,N_1178,N_1129);
or U2439 (N_2439,N_1019,N_1332);
or U2440 (N_2440,N_209,N_315);
and U2441 (N_2441,N_107,N_1637);
and U2442 (N_2442,N_496,N_1948);
or U2443 (N_2443,N_881,N_55);
or U2444 (N_2444,N_1419,N_1909);
nor U2445 (N_2445,N_870,N_704);
xnor U2446 (N_2446,N_758,N_1755);
nand U2447 (N_2447,N_527,N_491);
or U2448 (N_2448,N_112,N_1424);
or U2449 (N_2449,N_605,N_1620);
and U2450 (N_2450,N_1295,N_667);
and U2451 (N_2451,N_1030,N_347);
nand U2452 (N_2452,N_1667,N_1836);
or U2453 (N_2453,N_485,N_524);
nor U2454 (N_2454,N_584,N_482);
and U2455 (N_2455,N_493,N_1675);
nand U2456 (N_2456,N_395,N_1378);
nor U2457 (N_2457,N_216,N_916);
nor U2458 (N_2458,N_1018,N_274);
or U2459 (N_2459,N_1048,N_479);
nor U2460 (N_2460,N_1461,N_785);
or U2461 (N_2461,N_663,N_1575);
nor U2462 (N_2462,N_1607,N_1247);
and U2463 (N_2463,N_398,N_89);
xnor U2464 (N_2464,N_1227,N_1186);
nand U2465 (N_2465,N_1166,N_1705);
or U2466 (N_2466,N_751,N_937);
or U2467 (N_2467,N_672,N_30);
nand U2468 (N_2468,N_1962,N_1870);
or U2469 (N_2469,N_1852,N_841);
nand U2470 (N_2470,N_826,N_983);
nor U2471 (N_2471,N_219,N_748);
nor U2472 (N_2472,N_680,N_733);
and U2473 (N_2473,N_1244,N_1891);
and U2474 (N_2474,N_1738,N_776);
nand U2475 (N_2475,N_296,N_1735);
nand U2476 (N_2476,N_1793,N_239);
and U2477 (N_2477,N_1601,N_440);
and U2478 (N_2478,N_1182,N_695);
or U2479 (N_2479,N_1133,N_1970);
and U2480 (N_2480,N_675,N_1531);
nand U2481 (N_2481,N_843,N_772);
xnor U2482 (N_2482,N_938,N_1421);
nor U2483 (N_2483,N_867,N_595);
or U2484 (N_2484,N_964,N_557);
and U2485 (N_2485,N_1854,N_1055);
and U2486 (N_2486,N_510,N_1994);
and U2487 (N_2487,N_8,N_252);
nor U2488 (N_2488,N_1576,N_1137);
and U2489 (N_2489,N_1488,N_1794);
nor U2490 (N_2490,N_1164,N_1199);
or U2491 (N_2491,N_258,N_505);
xor U2492 (N_2492,N_1767,N_359);
and U2493 (N_2493,N_1702,N_1135);
and U2494 (N_2494,N_99,N_421);
or U2495 (N_2495,N_1672,N_525);
nand U2496 (N_2496,N_943,N_1827);
nand U2497 (N_2497,N_75,N_1808);
nor U2498 (N_2498,N_1613,N_1582);
nand U2499 (N_2499,N_1136,N_217);
and U2500 (N_2500,N_185,N_1899);
and U2501 (N_2501,N_79,N_150);
or U2502 (N_2502,N_948,N_997);
nand U2503 (N_2503,N_1486,N_590);
nor U2504 (N_2504,N_662,N_939);
xor U2505 (N_2505,N_1494,N_304);
or U2506 (N_2506,N_753,N_255);
and U2507 (N_2507,N_47,N_281);
nor U2508 (N_2508,N_1404,N_620);
and U2509 (N_2509,N_1154,N_686);
or U2510 (N_2510,N_445,N_236);
and U2511 (N_2511,N_470,N_1746);
or U2512 (N_2512,N_10,N_193);
xor U2513 (N_2513,N_1911,N_11);
nor U2514 (N_2514,N_1165,N_1093);
nand U2515 (N_2515,N_563,N_424);
and U2516 (N_2516,N_1587,N_1436);
nand U2517 (N_2517,N_1972,N_269);
nor U2518 (N_2518,N_905,N_1228);
and U2519 (N_2519,N_1989,N_1790);
nand U2520 (N_2520,N_581,N_1892);
nand U2521 (N_2521,N_31,N_796);
nand U2522 (N_2522,N_929,N_446);
and U2523 (N_2523,N_920,N_1919);
nor U2524 (N_2524,N_413,N_372);
and U2525 (N_2525,N_588,N_513);
or U2526 (N_2526,N_1014,N_25);
nor U2527 (N_2527,N_1976,N_1585);
nor U2528 (N_2528,N_1593,N_1291);
and U2529 (N_2529,N_1986,N_1180);
or U2530 (N_2530,N_597,N_1442);
or U2531 (N_2531,N_828,N_69);
or U2532 (N_2532,N_1861,N_635);
nor U2533 (N_2533,N_838,N_1425);
and U2534 (N_2534,N_898,N_226);
nor U2535 (N_2535,N_1833,N_989);
nor U2536 (N_2536,N_564,N_901);
nand U2537 (N_2537,N_520,N_729);
nor U2538 (N_2538,N_1068,N_382);
xor U2539 (N_2539,N_554,N_1863);
and U2540 (N_2540,N_1690,N_756);
nor U2541 (N_2541,N_593,N_183);
nor U2542 (N_2542,N_1402,N_1235);
and U2543 (N_2543,N_1039,N_414);
and U2544 (N_2544,N_1816,N_1454);
nand U2545 (N_2545,N_815,N_1536);
nor U2546 (N_2546,N_1713,N_1064);
nor U2547 (N_2547,N_1561,N_1982);
nor U2548 (N_2548,N_367,N_354);
nor U2549 (N_2549,N_876,N_1365);
xnor U2550 (N_2550,N_1558,N_692);
nor U2551 (N_2551,N_415,N_1610);
or U2552 (N_2552,N_773,N_1384);
and U2553 (N_2553,N_1452,N_1377);
nand U2554 (N_2554,N_1550,N_1603);
nor U2555 (N_2555,N_1880,N_314);
and U2556 (N_2556,N_298,N_1382);
nand U2557 (N_2557,N_1654,N_951);
nand U2558 (N_2558,N_1434,N_749);
or U2559 (N_2559,N_1510,N_235);
nor U2560 (N_2560,N_1612,N_128);
nand U2561 (N_2561,N_1966,N_890);
nand U2562 (N_2562,N_1838,N_1483);
nand U2563 (N_2563,N_1443,N_133);
and U2564 (N_2564,N_1769,N_1804);
nand U2565 (N_2565,N_1300,N_823);
or U2566 (N_2566,N_805,N_1522);
nand U2567 (N_2567,N_1786,N_833);
or U2568 (N_2568,N_713,N_710);
or U2569 (N_2569,N_515,N_961);
nor U2570 (N_2570,N_306,N_1063);
nand U2571 (N_2571,N_1659,N_140);
nor U2572 (N_2572,N_1524,N_1361);
nor U2573 (N_2573,N_1348,N_476);
or U2574 (N_2574,N_1475,N_1253);
nand U2575 (N_2575,N_362,N_1931);
or U2576 (N_2576,N_839,N_1876);
and U2577 (N_2577,N_1597,N_345);
nand U2578 (N_2578,N_769,N_1086);
nor U2579 (N_2579,N_1051,N_1451);
nand U2580 (N_2580,N_1347,N_526);
nor U2581 (N_2581,N_552,N_154);
nor U2582 (N_2582,N_1623,N_1697);
nor U2583 (N_2583,N_1196,N_175);
nor U2584 (N_2584,N_1636,N_1965);
and U2585 (N_2585,N_474,N_671);
and U2586 (N_2586,N_970,N_673);
or U2587 (N_2587,N_141,N_1414);
nand U2588 (N_2588,N_401,N_1239);
or U2589 (N_2589,N_659,N_1058);
nor U2590 (N_2590,N_1743,N_1848);
and U2591 (N_2591,N_1156,N_1271);
or U2592 (N_2592,N_851,N_957);
or U2593 (N_2593,N_317,N_862);
or U2594 (N_2594,N_1679,N_399);
nor U2595 (N_2595,N_53,N_735);
nand U2596 (N_2596,N_1694,N_460);
nand U2597 (N_2597,N_196,N_1544);
or U2598 (N_2598,N_1491,N_124);
or U2599 (N_2599,N_1949,N_62);
nand U2600 (N_2600,N_646,N_1759);
nor U2601 (N_2601,N_1803,N_602);
xor U2602 (N_2602,N_1884,N_535);
xnor U2603 (N_2603,N_690,N_1314);
or U2604 (N_2604,N_1555,N_371);
or U2605 (N_2605,N_1301,N_498);
nand U2606 (N_2606,N_1791,N_1340);
or U2607 (N_2607,N_1470,N_1220);
xnor U2608 (N_2608,N_734,N_1131);
and U2609 (N_2609,N_473,N_1933);
or U2610 (N_2610,N_20,N_509);
and U2611 (N_2611,N_1506,N_407);
xnor U2612 (N_2612,N_1010,N_1858);
nor U2613 (N_2613,N_392,N_1785);
and U2614 (N_2614,N_1683,N_689);
nor U2615 (N_2615,N_81,N_406);
nand U2616 (N_2616,N_316,N_968);
nand U2617 (N_2617,N_1066,N_499);
or U2618 (N_2618,N_1583,N_1503);
nor U2619 (N_2619,N_1049,N_678);
and U2620 (N_2620,N_583,N_1084);
nand U2621 (N_2621,N_254,N_253);
or U2622 (N_2622,N_893,N_1940);
nand U2623 (N_2623,N_917,N_1056);
or U2624 (N_2624,N_628,N_854);
xor U2625 (N_2625,N_1665,N_452);
and U2626 (N_2626,N_1311,N_831);
nor U2627 (N_2627,N_770,N_1801);
or U2628 (N_2628,N_125,N_1098);
nor U2629 (N_2629,N_1218,N_1934);
and U2630 (N_2630,N_1750,N_1813);
nand U2631 (N_2631,N_946,N_1930);
or U2632 (N_2632,N_203,N_35);
or U2633 (N_2633,N_1025,N_1723);
or U2634 (N_2634,N_958,N_98);
and U2635 (N_2635,N_1144,N_642);
nor U2636 (N_2636,N_1354,N_1005);
or U2637 (N_2637,N_1889,N_41);
and U2638 (N_2638,N_1973,N_151);
and U2639 (N_2639,N_490,N_224);
and U2640 (N_2640,N_576,N_1394);
nor U2641 (N_2641,N_1069,N_1869);
and U2642 (N_2642,N_1416,N_1763);
or U2643 (N_2643,N_1969,N_1719);
nor U2644 (N_2644,N_1034,N_1082);
nand U2645 (N_2645,N_986,N_1398);
xor U2646 (N_2646,N_360,N_872);
or U2647 (N_2647,N_1171,N_1213);
nand U2648 (N_2648,N_1617,N_1016);
and U2649 (N_2649,N_633,N_783);
nor U2650 (N_2650,N_875,N_1529);
nor U2651 (N_2651,N_290,N_1924);
and U2652 (N_2652,N_93,N_1240);
and U2653 (N_2653,N_1687,N_1729);
nand U2654 (N_2654,N_132,N_697);
or U2655 (N_2655,N_1918,N_707);
nand U2656 (N_2656,N_77,N_1928);
nor U2657 (N_2657,N_1353,N_1557);
nor U2658 (N_2658,N_1545,N_457);
and U2659 (N_2659,N_715,N_54);
nor U2660 (N_2660,N_1181,N_1162);
nand U2661 (N_2661,N_1445,N_1207);
nand U2662 (N_2662,N_766,N_369);
and U2663 (N_2663,N_1500,N_1481);
xor U2664 (N_2664,N_1073,N_311);
nand U2665 (N_2665,N_1812,N_1418);
or U2666 (N_2666,N_495,N_985);
and U2667 (N_2667,N_1864,N_575);
or U2668 (N_2668,N_346,N_1837);
nor U2669 (N_2669,N_16,N_1310);
nand U2670 (N_2670,N_444,N_461);
nor U2671 (N_2671,N_1277,N_164);
nor U2672 (N_2672,N_1726,N_911);
nand U2673 (N_2673,N_1287,N_169);
or U2674 (N_2674,N_1413,N_188);
nor U2675 (N_2675,N_1981,N_1927);
nand U2676 (N_2676,N_365,N_312);
or U2677 (N_2677,N_187,N_962);
and U2678 (N_2678,N_926,N_276);
nor U2679 (N_2679,N_172,N_1478);
nor U2680 (N_2680,N_106,N_1774);
and U2681 (N_2681,N_1564,N_1173);
nand U2682 (N_2682,N_1885,N_364);
nor U2683 (N_2683,N_501,N_68);
and U2684 (N_2684,N_984,N_1169);
nand U2685 (N_2685,N_1463,N_859);
and U2686 (N_2686,N_1118,N_1547);
and U2687 (N_2687,N_761,N_56);
nor U2688 (N_2688,N_471,N_1789);
and U2689 (N_2689,N_1233,N_1968);
nor U2690 (N_2690,N_1588,N_1745);
nor U2691 (N_2691,N_357,N_950);
nor U2692 (N_2692,N_1124,N_900);
nand U2693 (N_2693,N_1147,N_711);
nor U2694 (N_2694,N_1229,N_1001);
or U2695 (N_2695,N_227,N_741);
nor U2696 (N_2696,N_307,N_846);
nand U2697 (N_2697,N_1197,N_386);
nor U2698 (N_2698,N_918,N_1479);
nor U2699 (N_2699,N_1299,N_1872);
nand U2700 (N_2700,N_1415,N_396);
nor U2701 (N_2701,N_1839,N_1160);
or U2702 (N_2702,N_1263,N_560);
xnor U2703 (N_2703,N_1183,N_438);
or U2704 (N_2704,N_591,N_788);
nor U2705 (N_2705,N_1033,N_1031);
nand U2706 (N_2706,N_1947,N_1819);
and U2707 (N_2707,N_1185,N_1526);
and U2708 (N_2708,N_1139,N_1740);
nor U2709 (N_2709,N_71,N_1223);
nand U2710 (N_2710,N_661,N_546);
nand U2711 (N_2711,N_439,N_7);
xnor U2712 (N_2712,N_1708,N_36);
nor U2713 (N_2713,N_1766,N_1900);
or U2714 (N_2714,N_113,N_631);
nor U2715 (N_2715,N_40,N_855);
nor U2716 (N_2716,N_1071,N_718);
nand U2717 (N_2717,N_1307,N_771);
nand U2718 (N_2718,N_1412,N_1308);
nand U2719 (N_2719,N_1091,N_1992);
nor U2720 (N_2720,N_1539,N_668);
nand U2721 (N_2721,N_1141,N_1221);
nor U2722 (N_2722,N_1266,N_1799);
nand U2723 (N_2723,N_627,N_1490);
xnor U2724 (N_2724,N_1493,N_883);
or U2725 (N_2725,N_1628,N_1579);
or U2726 (N_2726,N_1052,N_283);
and U2727 (N_2727,N_1897,N_1422);
xor U2728 (N_2728,N_640,N_1570);
and U2729 (N_2729,N_300,N_325);
nand U2730 (N_2730,N_318,N_1997);
nor U2731 (N_2731,N_1121,N_51);
nor U2732 (N_2732,N_1006,N_1342);
nand U2733 (N_2733,N_1741,N_1760);
nand U2734 (N_2734,N_1265,N_264);
and U2735 (N_2735,N_1920,N_924);
and U2736 (N_2736,N_1709,N_1756);
nand U2737 (N_2737,N_1047,N_1518);
nand U2738 (N_2738,N_230,N_231);
or U2739 (N_2739,N_207,N_910);
and U2740 (N_2740,N_500,N_1890);
nand U2741 (N_2741,N_0,N_1343);
and U2742 (N_2742,N_275,N_573);
nand U2743 (N_2743,N_956,N_1441);
nor U2744 (N_2744,N_969,N_1633);
nand U2745 (N_2745,N_517,N_988);
nand U2746 (N_2746,N_1898,N_119);
nand U2747 (N_2747,N_1296,N_799);
and U2748 (N_2748,N_798,N_945);
and U2749 (N_2749,N_936,N_61);
or U2750 (N_2750,N_18,N_978);
nand U2751 (N_2751,N_1517,N_1336);
and U2752 (N_2752,N_580,N_1020);
nor U2753 (N_2753,N_1658,N_1157);
xnor U2754 (N_2754,N_293,N_940);
nand U2755 (N_2755,N_466,N_702);
and U2756 (N_2756,N_1787,N_1896);
xor U2757 (N_2757,N_863,N_848);
nand U2758 (N_2758,N_420,N_1621);
and U2759 (N_2759,N_28,N_19);
nand U2760 (N_2760,N_1875,N_1644);
xor U2761 (N_2761,N_337,N_1472);
or U2762 (N_2762,N_1356,N_1850);
nand U2763 (N_2763,N_806,N_100);
nand U2764 (N_2764,N_1187,N_1145);
nor U2765 (N_2765,N_763,N_636);
nor U2766 (N_2766,N_1655,N_443);
nand U2767 (N_2767,N_91,N_1484);
or U2768 (N_2768,N_1386,N_1264);
and U2769 (N_2769,N_441,N_1874);
nor U2770 (N_2770,N_714,N_210);
or U2771 (N_2771,N_263,N_1714);
nor U2772 (N_2772,N_779,N_601);
nand U2773 (N_2773,N_789,N_2);
nand U2774 (N_2774,N_712,N_4);
nor U2775 (N_2775,N_259,N_181);
and U2776 (N_2776,N_1188,N_303);
and U2777 (N_2777,N_1373,N_14);
and U2778 (N_2778,N_1905,N_1420);
nor U2779 (N_2779,N_1236,N_1523);
nor U2780 (N_2780,N_536,N_222);
and U2781 (N_2781,N_1528,N_533);
and U2782 (N_2782,N_1842,N_1459);
xnor U2783 (N_2783,N_1423,N_822);
nand U2784 (N_2784,N_1067,N_191);
nor U2785 (N_2785,N_1390,N_1853);
nand U2786 (N_2786,N_408,N_600);
nand U2787 (N_2787,N_1119,N_1106);
and U2788 (N_2788,N_243,N_1011);
or U2789 (N_2789,N_541,N_261);
or U2790 (N_2790,N_411,N_118);
and U2791 (N_2791,N_96,N_1820);
nor U2792 (N_2792,N_1023,N_288);
and U2793 (N_2793,N_860,N_433);
nand U2794 (N_2794,N_29,N_1608);
or U2795 (N_2795,N_97,N_547);
or U2796 (N_2796,N_1170,N_980);
and U2797 (N_2797,N_57,N_34);
nor U2798 (N_2798,N_1250,N_578);
and U2799 (N_2799,N_1802,N_1695);
or U2800 (N_2800,N_1408,N_393);
and U2801 (N_2801,N_608,N_1562);
or U2802 (N_2802,N_907,N_368);
nor U2803 (N_2803,N_1721,N_1814);
or U2804 (N_2804,N_374,N_716);
xnor U2805 (N_2805,N_1825,N_475);
and U2806 (N_2806,N_1433,N_906);
nand U2807 (N_2807,N_797,N_404);
nor U2808 (N_2808,N_126,N_1844);
nor U2809 (N_2809,N_162,N_1159);
and U2810 (N_2810,N_1826,N_1904);
or U2811 (N_2811,N_1998,N_795);
and U2812 (N_2812,N_1985,N_277);
nor U2813 (N_2813,N_1591,N_110);
xnor U2814 (N_2814,N_555,N_1571);
or U2815 (N_2815,N_1321,N_215);
and U2816 (N_2816,N_1540,N_840);
or U2817 (N_2817,N_1174,N_1392);
and U2818 (N_2818,N_933,N_1711);
or U2819 (N_2819,N_1916,N_1865);
and U2820 (N_2820,N_1984,N_78);
xor U2821 (N_2821,N_1466,N_1988);
nand U2822 (N_2822,N_1980,N_423);
and U2823 (N_2823,N_1163,N_1829);
nand U2824 (N_2824,N_158,N_131);
nand U2825 (N_2825,N_819,N_750);
nand U2826 (N_2826,N_1462,N_137);
nor U2827 (N_2827,N_1078,N_1674);
and U2828 (N_2828,N_1888,N_908);
nor U2829 (N_2829,N_1797,N_836);
nand U2830 (N_2830,N_1810,N_1021);
and U2831 (N_2831,N_64,N_699);
nor U2832 (N_2832,N_442,N_1238);
nor U2833 (N_2833,N_941,N_1527);
nand U2834 (N_2834,N_1333,N_682);
and U2835 (N_2835,N_932,N_694);
or U2836 (N_2836,N_1335,N_849);
nand U2837 (N_2837,N_1867,N_1739);
nand U2838 (N_2838,N_1241,N_1177);
and U2839 (N_2839,N_1274,N_1487);
and U2840 (N_2840,N_184,N_1201);
and U2841 (N_2841,N_530,N_921);
and U2842 (N_2842,N_1657,N_742);
and U2843 (N_2843,N_1088,N_272);
nand U2844 (N_2844,N_1385,N_378);
and U2845 (N_2845,N_871,N_1855);
nand U2846 (N_2846,N_639,N_1776);
nor U2847 (N_2847,N_1622,N_250);
nor U2848 (N_2848,N_1152,N_674);
and U2849 (N_2849,N_111,N_1380);
and U2850 (N_2850,N_144,N_1195);
nand U2851 (N_2851,N_1367,N_1293);
and U2852 (N_2852,N_1369,N_1457);
nand U2853 (N_2853,N_1943,N_1684);
nor U2854 (N_2854,N_260,N_1435);
and U2855 (N_2855,N_852,N_1736);
nor U2856 (N_2856,N_856,N_1663);
nand U2857 (N_2857,N_518,N_1495);
or U2858 (N_2858,N_1095,N_1279);
nand U2859 (N_2859,N_1440,N_1757);
xnor U2860 (N_2860,N_955,N_74);
or U2861 (N_2861,N_610,N_1012);
or U2862 (N_2862,N_1798,N_449);
and U2863 (N_2863,N_1072,N_1589);
nor U2864 (N_2864,N_1830,N_1113);
nand U2865 (N_2865,N_994,N_880);
nor U2866 (N_2866,N_1374,N_780);
nor U2867 (N_2867,N_1953,N_1224);
or U2868 (N_2868,N_170,N_1102);
nand U2869 (N_2869,N_331,N_426);
or U2870 (N_2870,N_221,N_1211);
nor U2871 (N_2871,N_960,N_376);
nor U2872 (N_2872,N_654,N_90);
and U2873 (N_2873,N_292,N_1456);
xnor U2874 (N_2874,N_148,N_637);
nor U2875 (N_2875,N_1772,N_387);
and U2876 (N_2876,N_1945,N_1116);
or U2877 (N_2877,N_1190,N_394);
and U2878 (N_2878,N_1586,N_1259);
xnor U2879 (N_2879,N_873,N_1678);
nor U2880 (N_2880,N_1003,N_1115);
nand U2881 (N_2881,N_607,N_1846);
and U2882 (N_2882,N_811,N_1818);
and U2883 (N_2883,N_705,N_810);
nand U2884 (N_2884,N_65,N_582);
nand U2885 (N_2885,N_914,N_1879);
xnor U2886 (N_2886,N_330,N_1698);
or U2887 (N_2887,N_514,N_1397);
nor U2888 (N_2888,N_1114,N_1626);
or U2889 (N_2889,N_1625,N_1303);
or U2890 (N_2890,N_232,N_173);
xnor U2891 (N_2891,N_416,N_1411);
and U2892 (N_2892,N_708,N_1635);
nand U2893 (N_2893,N_397,N_1783);
and U2894 (N_2894,N_1132,N_1543);
or U2895 (N_2895,N_1704,N_1761);
or U2896 (N_2896,N_1097,N_1357);
or U2897 (N_2897,N_268,N_1926);
nor U2898 (N_2898,N_85,N_1614);
nand U2899 (N_2899,N_1059,N_1316);
nor U2900 (N_2900,N_1476,N_1015);
nor U2901 (N_2901,N_1598,N_1513);
nor U2902 (N_2902,N_1209,N_1996);
or U2903 (N_2903,N_436,N_865);
or U2904 (N_2904,N_1815,N_1643);
nand U2905 (N_2905,N_73,N_802);
nand U2906 (N_2906,N_1319,N_180);
and U2907 (N_2907,N_622,N_1261);
nand U2908 (N_2908,N_1426,N_1525);
or U2909 (N_2909,N_1351,N_1427);
nor U2910 (N_2910,N_827,N_1323);
nand U2911 (N_2911,N_329,N_1450);
nand U2912 (N_2912,N_464,N_1294);
nor U2913 (N_2913,N_567,N_348);
and U2914 (N_2914,N_594,N_1796);
and U2915 (N_2915,N_979,N_76);
nand U2916 (N_2916,N_1245,N_1649);
or U2917 (N_2917,N_596,N_1128);
and U2918 (N_2918,N_626,N_814);
or U2919 (N_2919,N_486,N_1893);
and U2920 (N_2920,N_845,N_366);
or U2921 (N_2921,N_746,N_643);
nor U2922 (N_2922,N_1781,N_1584);
and U2923 (N_2923,N_842,N_1748);
nand U2924 (N_2924,N_587,N_971);
nor U2925 (N_2925,N_349,N_1627);
nor U2926 (N_2926,N_861,N_176);
nand U2927 (N_2927,N_286,N_130);
nand U2928 (N_2928,N_894,N_313);
and U2929 (N_2929,N_1219,N_634);
or U2930 (N_2930,N_1646,N_391);
nand U2931 (N_2931,N_1192,N_13);
nor U2932 (N_2932,N_1306,N_1632);
or U2933 (N_2933,N_1155,N_1032);
and U2934 (N_2934,N_251,N_1784);
or U2935 (N_2935,N_1952,N_550);
nor U2936 (N_2936,N_1686,N_1754);
nand U2937 (N_2937,N_1252,N_1600);
or U2938 (N_2938,N_1401,N_1553);
and U2939 (N_2939,N_534,N_1044);
or U2940 (N_2940,N_488,N_238);
and U2941 (N_2941,N_1859,N_529);
nor U2942 (N_2942,N_278,N_1516);
and U2943 (N_2943,N_723,N_1773);
and U2944 (N_2944,N_1770,N_83);
nand U2945 (N_2945,N_952,N_24);
nand U2946 (N_2946,N_738,N_1138);
or U2947 (N_2947,N_1717,N_569);
xnor U2948 (N_2948,N_598,N_651);
nand U2949 (N_2949,N_1727,N_850);
or U2950 (N_2950,N_1505,N_1448);
nand U2951 (N_2951,N_105,N_49);
nand U2952 (N_2952,N_1035,N_623);
and U2953 (N_2953,N_1081,N_1087);
nand U2954 (N_2954,N_1120,N_1851);
xnor U2955 (N_2955,N_43,N_1123);
and U2956 (N_2956,N_556,N_947);
nor U2957 (N_2957,N_212,N_1534);
or U2958 (N_2958,N_1502,N_52);
nor U2959 (N_2959,N_156,N_820);
xor U2960 (N_2960,N_585,N_326);
and U2961 (N_2961,N_899,N_722);
nand U2962 (N_2962,N_1877,N_225);
and U2963 (N_2963,N_915,N_1103);
xor U2964 (N_2964,N_736,N_657);
or U2965 (N_2965,N_558,N_1722);
or U2966 (N_2966,N_1913,N_658);
nor U2967 (N_2967,N_1007,N_1153);
nor U2968 (N_2968,N_1515,N_1730);
and U2969 (N_2969,N_930,N_1946);
or U2970 (N_2970,N_676,N_912);
xor U2971 (N_2971,N_992,N_1337);
nand U2972 (N_2972,N_853,N_1552);
nand U2973 (N_2973,N_522,N_157);
nand U2974 (N_2974,N_1329,N_878);
nand U2975 (N_2975,N_1936,N_1065);
nor U2976 (N_2976,N_134,N_428);
nand U2977 (N_2977,N_233,N_1070);
nor U2978 (N_2978,N_487,N_390);
or U2979 (N_2979,N_135,N_199);
nand U2980 (N_2980,N_532,N_380);
or U2981 (N_2981,N_619,N_1127);
xnor U2982 (N_2982,N_531,N_87);
or U2983 (N_2983,N_542,N_1577);
or U2984 (N_2984,N_1057,N_12);
nand U2985 (N_2985,N_847,N_1322);
nand U2986 (N_2986,N_885,N_1172);
nand U2987 (N_2987,N_1092,N_1275);
xor U2988 (N_2988,N_650,N_974);
nor U2989 (N_2989,N_807,N_652);
and U2990 (N_2990,N_1498,N_409);
nand U2991 (N_2991,N_1094,N_857);
nand U2992 (N_2992,N_791,N_467);
and U2993 (N_2993,N_437,N_877);
and U2994 (N_2994,N_696,N_1482);
and U2995 (N_2995,N_418,N_612);
or U2996 (N_2996,N_688,N_282);
and U2997 (N_2997,N_1573,N_142);
nor U2998 (N_2998,N_384,N_787);
nand U2999 (N_2999,N_923,N_1428);
or U3000 (N_3000,N_433,N_879);
and U3001 (N_3001,N_1303,N_1699);
nand U3002 (N_3002,N_362,N_51);
or U3003 (N_3003,N_1580,N_1212);
nand U3004 (N_3004,N_1847,N_288);
and U3005 (N_3005,N_229,N_50);
nor U3006 (N_3006,N_1847,N_153);
and U3007 (N_3007,N_1846,N_828);
and U3008 (N_3008,N_544,N_1472);
and U3009 (N_3009,N_784,N_379);
or U3010 (N_3010,N_88,N_1676);
nand U3011 (N_3011,N_735,N_1497);
or U3012 (N_3012,N_107,N_1875);
nand U3013 (N_3013,N_1998,N_867);
nor U3014 (N_3014,N_1789,N_91);
nand U3015 (N_3015,N_303,N_156);
and U3016 (N_3016,N_864,N_1532);
nor U3017 (N_3017,N_146,N_679);
nor U3018 (N_3018,N_767,N_108);
and U3019 (N_3019,N_599,N_1477);
nor U3020 (N_3020,N_401,N_870);
and U3021 (N_3021,N_782,N_1039);
xnor U3022 (N_3022,N_681,N_1140);
or U3023 (N_3023,N_1386,N_939);
or U3024 (N_3024,N_522,N_369);
nand U3025 (N_3025,N_712,N_1159);
or U3026 (N_3026,N_1073,N_1277);
nand U3027 (N_3027,N_955,N_840);
xnor U3028 (N_3028,N_1504,N_1810);
nand U3029 (N_3029,N_1260,N_1573);
or U3030 (N_3030,N_177,N_980);
and U3031 (N_3031,N_1933,N_156);
nand U3032 (N_3032,N_1266,N_1700);
and U3033 (N_3033,N_812,N_1101);
or U3034 (N_3034,N_1759,N_451);
and U3035 (N_3035,N_1389,N_972);
nand U3036 (N_3036,N_919,N_1671);
and U3037 (N_3037,N_259,N_1309);
or U3038 (N_3038,N_1077,N_455);
nand U3039 (N_3039,N_675,N_1059);
or U3040 (N_3040,N_1469,N_1529);
or U3041 (N_3041,N_833,N_39);
and U3042 (N_3042,N_1467,N_276);
nand U3043 (N_3043,N_1243,N_619);
and U3044 (N_3044,N_1592,N_568);
nand U3045 (N_3045,N_425,N_1652);
and U3046 (N_3046,N_902,N_1985);
nand U3047 (N_3047,N_745,N_1296);
and U3048 (N_3048,N_933,N_1449);
and U3049 (N_3049,N_970,N_992);
or U3050 (N_3050,N_1035,N_278);
nand U3051 (N_3051,N_855,N_924);
nand U3052 (N_3052,N_1695,N_1186);
nand U3053 (N_3053,N_99,N_1076);
xor U3054 (N_3054,N_1598,N_1410);
xnor U3055 (N_3055,N_1355,N_763);
or U3056 (N_3056,N_1257,N_1170);
nor U3057 (N_3057,N_354,N_1633);
or U3058 (N_3058,N_1568,N_533);
and U3059 (N_3059,N_711,N_511);
nand U3060 (N_3060,N_1120,N_414);
and U3061 (N_3061,N_1647,N_389);
and U3062 (N_3062,N_420,N_1733);
or U3063 (N_3063,N_1193,N_1779);
nand U3064 (N_3064,N_329,N_1692);
or U3065 (N_3065,N_1920,N_297);
nor U3066 (N_3066,N_1135,N_1962);
and U3067 (N_3067,N_588,N_1237);
nor U3068 (N_3068,N_1159,N_80);
and U3069 (N_3069,N_70,N_1413);
nand U3070 (N_3070,N_7,N_646);
or U3071 (N_3071,N_1818,N_1558);
nor U3072 (N_3072,N_441,N_791);
nand U3073 (N_3073,N_1157,N_231);
nand U3074 (N_3074,N_923,N_1636);
and U3075 (N_3075,N_1557,N_1276);
nand U3076 (N_3076,N_803,N_462);
nand U3077 (N_3077,N_1736,N_1249);
and U3078 (N_3078,N_1563,N_1738);
or U3079 (N_3079,N_913,N_1957);
and U3080 (N_3080,N_1949,N_170);
nand U3081 (N_3081,N_1861,N_1229);
or U3082 (N_3082,N_649,N_9);
nor U3083 (N_3083,N_1380,N_1127);
nor U3084 (N_3084,N_1253,N_617);
xnor U3085 (N_3085,N_520,N_533);
and U3086 (N_3086,N_593,N_1857);
and U3087 (N_3087,N_1886,N_636);
nor U3088 (N_3088,N_51,N_295);
xor U3089 (N_3089,N_500,N_22);
and U3090 (N_3090,N_1670,N_770);
nand U3091 (N_3091,N_828,N_928);
and U3092 (N_3092,N_512,N_288);
nor U3093 (N_3093,N_1557,N_103);
xor U3094 (N_3094,N_893,N_519);
and U3095 (N_3095,N_1039,N_990);
or U3096 (N_3096,N_324,N_43);
and U3097 (N_3097,N_518,N_583);
nand U3098 (N_3098,N_1571,N_1547);
and U3099 (N_3099,N_1635,N_1388);
and U3100 (N_3100,N_1037,N_855);
and U3101 (N_3101,N_252,N_1805);
nand U3102 (N_3102,N_472,N_263);
or U3103 (N_3103,N_69,N_1773);
and U3104 (N_3104,N_293,N_1764);
and U3105 (N_3105,N_879,N_1609);
or U3106 (N_3106,N_1306,N_43);
or U3107 (N_3107,N_1203,N_1797);
or U3108 (N_3108,N_1175,N_769);
or U3109 (N_3109,N_524,N_967);
and U3110 (N_3110,N_1385,N_211);
nand U3111 (N_3111,N_1596,N_337);
and U3112 (N_3112,N_1636,N_552);
nor U3113 (N_3113,N_707,N_173);
and U3114 (N_3114,N_1848,N_741);
and U3115 (N_3115,N_517,N_443);
and U3116 (N_3116,N_1441,N_1347);
xnor U3117 (N_3117,N_989,N_619);
nor U3118 (N_3118,N_43,N_1384);
nor U3119 (N_3119,N_1227,N_521);
and U3120 (N_3120,N_1833,N_695);
nand U3121 (N_3121,N_1119,N_198);
or U3122 (N_3122,N_816,N_1881);
nor U3123 (N_3123,N_204,N_227);
or U3124 (N_3124,N_1343,N_1065);
and U3125 (N_3125,N_1264,N_556);
or U3126 (N_3126,N_1160,N_1531);
nand U3127 (N_3127,N_1536,N_631);
nand U3128 (N_3128,N_1071,N_868);
nor U3129 (N_3129,N_270,N_1739);
nand U3130 (N_3130,N_1740,N_1731);
nand U3131 (N_3131,N_713,N_1648);
nand U3132 (N_3132,N_1742,N_1667);
xor U3133 (N_3133,N_1379,N_33);
nor U3134 (N_3134,N_1883,N_1781);
or U3135 (N_3135,N_1169,N_738);
nand U3136 (N_3136,N_28,N_262);
or U3137 (N_3137,N_259,N_1020);
or U3138 (N_3138,N_1132,N_1286);
nor U3139 (N_3139,N_232,N_709);
nor U3140 (N_3140,N_1130,N_1058);
nand U3141 (N_3141,N_1906,N_1023);
nand U3142 (N_3142,N_1017,N_13);
or U3143 (N_3143,N_1744,N_1942);
or U3144 (N_3144,N_750,N_122);
and U3145 (N_3145,N_437,N_1508);
xor U3146 (N_3146,N_392,N_545);
and U3147 (N_3147,N_872,N_1495);
and U3148 (N_3148,N_1141,N_904);
or U3149 (N_3149,N_1101,N_906);
nand U3150 (N_3150,N_1478,N_504);
and U3151 (N_3151,N_551,N_387);
or U3152 (N_3152,N_1031,N_1431);
nand U3153 (N_3153,N_237,N_1487);
xor U3154 (N_3154,N_1632,N_813);
or U3155 (N_3155,N_799,N_1673);
nor U3156 (N_3156,N_1635,N_156);
nand U3157 (N_3157,N_37,N_253);
or U3158 (N_3158,N_206,N_1520);
or U3159 (N_3159,N_881,N_392);
xnor U3160 (N_3160,N_516,N_620);
and U3161 (N_3161,N_1585,N_1197);
nand U3162 (N_3162,N_1475,N_211);
nor U3163 (N_3163,N_1548,N_1334);
nor U3164 (N_3164,N_1471,N_1790);
xnor U3165 (N_3165,N_1445,N_1231);
nand U3166 (N_3166,N_672,N_61);
or U3167 (N_3167,N_1831,N_341);
or U3168 (N_3168,N_701,N_884);
and U3169 (N_3169,N_55,N_1381);
nand U3170 (N_3170,N_1619,N_1096);
nand U3171 (N_3171,N_1928,N_1371);
nor U3172 (N_3172,N_1608,N_1321);
xor U3173 (N_3173,N_112,N_1129);
nand U3174 (N_3174,N_907,N_1536);
or U3175 (N_3175,N_1895,N_1694);
xor U3176 (N_3176,N_1936,N_1360);
nor U3177 (N_3177,N_799,N_247);
nand U3178 (N_3178,N_319,N_110);
xnor U3179 (N_3179,N_352,N_1078);
nor U3180 (N_3180,N_331,N_506);
nand U3181 (N_3181,N_1354,N_1379);
nand U3182 (N_3182,N_1807,N_92);
nand U3183 (N_3183,N_1950,N_792);
or U3184 (N_3184,N_491,N_25);
nand U3185 (N_3185,N_245,N_1178);
nand U3186 (N_3186,N_342,N_584);
or U3187 (N_3187,N_584,N_1016);
xnor U3188 (N_3188,N_415,N_1444);
or U3189 (N_3189,N_822,N_1236);
and U3190 (N_3190,N_585,N_1551);
xor U3191 (N_3191,N_959,N_1380);
nor U3192 (N_3192,N_505,N_817);
nand U3193 (N_3193,N_1825,N_981);
xor U3194 (N_3194,N_1238,N_1688);
and U3195 (N_3195,N_843,N_977);
or U3196 (N_3196,N_874,N_1845);
or U3197 (N_3197,N_915,N_1908);
and U3198 (N_3198,N_1032,N_609);
xnor U3199 (N_3199,N_1257,N_360);
or U3200 (N_3200,N_258,N_1174);
or U3201 (N_3201,N_460,N_11);
xor U3202 (N_3202,N_835,N_949);
and U3203 (N_3203,N_1586,N_1050);
or U3204 (N_3204,N_109,N_660);
xor U3205 (N_3205,N_475,N_166);
or U3206 (N_3206,N_956,N_1299);
xor U3207 (N_3207,N_1168,N_1138);
nor U3208 (N_3208,N_1650,N_808);
xnor U3209 (N_3209,N_39,N_1889);
nor U3210 (N_3210,N_1300,N_1735);
and U3211 (N_3211,N_477,N_1850);
nand U3212 (N_3212,N_1290,N_1749);
nor U3213 (N_3213,N_910,N_31);
and U3214 (N_3214,N_477,N_1070);
nor U3215 (N_3215,N_1510,N_930);
or U3216 (N_3216,N_874,N_287);
nor U3217 (N_3217,N_1008,N_954);
xnor U3218 (N_3218,N_1313,N_1012);
nor U3219 (N_3219,N_322,N_1358);
and U3220 (N_3220,N_1425,N_596);
or U3221 (N_3221,N_331,N_782);
nand U3222 (N_3222,N_475,N_755);
nor U3223 (N_3223,N_1671,N_876);
and U3224 (N_3224,N_1459,N_1422);
or U3225 (N_3225,N_1915,N_1140);
and U3226 (N_3226,N_309,N_960);
xnor U3227 (N_3227,N_1195,N_1987);
nand U3228 (N_3228,N_1215,N_1970);
and U3229 (N_3229,N_134,N_1214);
xor U3230 (N_3230,N_1010,N_1647);
and U3231 (N_3231,N_97,N_338);
nand U3232 (N_3232,N_1722,N_1017);
and U3233 (N_3233,N_210,N_1603);
nand U3234 (N_3234,N_1557,N_1872);
nor U3235 (N_3235,N_777,N_80);
nand U3236 (N_3236,N_809,N_795);
nor U3237 (N_3237,N_1736,N_445);
nor U3238 (N_3238,N_1641,N_330);
and U3239 (N_3239,N_1805,N_647);
and U3240 (N_3240,N_1295,N_687);
or U3241 (N_3241,N_711,N_414);
nand U3242 (N_3242,N_1753,N_1428);
and U3243 (N_3243,N_556,N_1836);
nand U3244 (N_3244,N_104,N_70);
or U3245 (N_3245,N_563,N_835);
and U3246 (N_3246,N_1795,N_251);
nand U3247 (N_3247,N_1319,N_775);
nor U3248 (N_3248,N_424,N_1177);
and U3249 (N_3249,N_750,N_74);
nand U3250 (N_3250,N_1873,N_675);
nand U3251 (N_3251,N_1989,N_1918);
or U3252 (N_3252,N_1639,N_1915);
and U3253 (N_3253,N_539,N_1606);
or U3254 (N_3254,N_614,N_1117);
and U3255 (N_3255,N_1238,N_67);
or U3256 (N_3256,N_226,N_1663);
nor U3257 (N_3257,N_855,N_1947);
or U3258 (N_3258,N_1027,N_720);
nand U3259 (N_3259,N_212,N_1163);
and U3260 (N_3260,N_1765,N_1142);
nand U3261 (N_3261,N_1083,N_1952);
nor U3262 (N_3262,N_148,N_900);
nor U3263 (N_3263,N_905,N_1995);
or U3264 (N_3264,N_298,N_822);
nor U3265 (N_3265,N_986,N_865);
nand U3266 (N_3266,N_974,N_850);
nor U3267 (N_3267,N_2,N_1642);
xnor U3268 (N_3268,N_1386,N_371);
and U3269 (N_3269,N_1430,N_1965);
nand U3270 (N_3270,N_482,N_1086);
or U3271 (N_3271,N_365,N_1122);
and U3272 (N_3272,N_1576,N_1738);
nand U3273 (N_3273,N_1576,N_1113);
nor U3274 (N_3274,N_1896,N_1728);
and U3275 (N_3275,N_829,N_1587);
and U3276 (N_3276,N_1383,N_346);
nor U3277 (N_3277,N_1996,N_222);
or U3278 (N_3278,N_802,N_1788);
nand U3279 (N_3279,N_1842,N_1446);
or U3280 (N_3280,N_1760,N_1873);
or U3281 (N_3281,N_1139,N_100);
and U3282 (N_3282,N_1301,N_590);
or U3283 (N_3283,N_179,N_68);
nand U3284 (N_3284,N_1370,N_1063);
and U3285 (N_3285,N_1675,N_918);
and U3286 (N_3286,N_444,N_473);
and U3287 (N_3287,N_1831,N_1982);
nor U3288 (N_3288,N_1148,N_916);
or U3289 (N_3289,N_755,N_1610);
and U3290 (N_3290,N_1792,N_198);
or U3291 (N_3291,N_1255,N_991);
nor U3292 (N_3292,N_1683,N_325);
or U3293 (N_3293,N_1927,N_514);
nand U3294 (N_3294,N_1939,N_1896);
or U3295 (N_3295,N_788,N_968);
xor U3296 (N_3296,N_1097,N_1749);
or U3297 (N_3297,N_991,N_275);
xor U3298 (N_3298,N_1290,N_38);
nand U3299 (N_3299,N_717,N_76);
or U3300 (N_3300,N_1308,N_1616);
and U3301 (N_3301,N_385,N_753);
nand U3302 (N_3302,N_50,N_923);
xnor U3303 (N_3303,N_449,N_684);
or U3304 (N_3304,N_1475,N_1414);
or U3305 (N_3305,N_1349,N_1391);
xor U3306 (N_3306,N_1841,N_1074);
nand U3307 (N_3307,N_394,N_1833);
nor U3308 (N_3308,N_636,N_219);
nor U3309 (N_3309,N_885,N_1939);
and U3310 (N_3310,N_1537,N_1315);
nand U3311 (N_3311,N_1212,N_705);
or U3312 (N_3312,N_892,N_356);
or U3313 (N_3313,N_255,N_952);
nand U3314 (N_3314,N_959,N_90);
xnor U3315 (N_3315,N_1662,N_1303);
nor U3316 (N_3316,N_481,N_1236);
xor U3317 (N_3317,N_1001,N_56);
and U3318 (N_3318,N_1284,N_1015);
nand U3319 (N_3319,N_294,N_929);
nand U3320 (N_3320,N_1236,N_984);
nor U3321 (N_3321,N_90,N_1428);
nand U3322 (N_3322,N_1714,N_810);
nand U3323 (N_3323,N_1257,N_1786);
nand U3324 (N_3324,N_1802,N_678);
and U3325 (N_3325,N_1138,N_425);
or U3326 (N_3326,N_638,N_1455);
and U3327 (N_3327,N_436,N_1222);
nor U3328 (N_3328,N_1577,N_902);
nand U3329 (N_3329,N_1837,N_1155);
nand U3330 (N_3330,N_1212,N_96);
nand U3331 (N_3331,N_1343,N_1247);
and U3332 (N_3332,N_1579,N_1);
or U3333 (N_3333,N_1801,N_1426);
nor U3334 (N_3334,N_977,N_908);
xnor U3335 (N_3335,N_969,N_268);
nand U3336 (N_3336,N_1738,N_1048);
nor U3337 (N_3337,N_1019,N_1470);
or U3338 (N_3338,N_735,N_182);
nand U3339 (N_3339,N_56,N_344);
xnor U3340 (N_3340,N_323,N_1651);
nand U3341 (N_3341,N_252,N_148);
and U3342 (N_3342,N_121,N_607);
nor U3343 (N_3343,N_393,N_260);
nor U3344 (N_3344,N_338,N_33);
nand U3345 (N_3345,N_1297,N_561);
nor U3346 (N_3346,N_1024,N_1537);
nand U3347 (N_3347,N_123,N_534);
and U3348 (N_3348,N_164,N_1381);
and U3349 (N_3349,N_316,N_262);
nor U3350 (N_3350,N_230,N_1147);
nand U3351 (N_3351,N_917,N_1952);
nand U3352 (N_3352,N_821,N_1316);
nor U3353 (N_3353,N_1864,N_636);
and U3354 (N_3354,N_956,N_1772);
nor U3355 (N_3355,N_1971,N_133);
and U3356 (N_3356,N_363,N_1882);
nor U3357 (N_3357,N_1438,N_584);
and U3358 (N_3358,N_1764,N_1680);
or U3359 (N_3359,N_581,N_963);
nand U3360 (N_3360,N_4,N_1621);
xnor U3361 (N_3361,N_1823,N_1619);
and U3362 (N_3362,N_220,N_196);
or U3363 (N_3363,N_562,N_1741);
xor U3364 (N_3364,N_257,N_1896);
xnor U3365 (N_3365,N_1375,N_1958);
and U3366 (N_3366,N_241,N_192);
and U3367 (N_3367,N_745,N_1986);
nand U3368 (N_3368,N_1635,N_881);
nand U3369 (N_3369,N_1538,N_558);
and U3370 (N_3370,N_1671,N_221);
nor U3371 (N_3371,N_246,N_450);
nand U3372 (N_3372,N_1190,N_647);
nand U3373 (N_3373,N_1004,N_1916);
nand U3374 (N_3374,N_908,N_70);
nor U3375 (N_3375,N_864,N_342);
nor U3376 (N_3376,N_1592,N_102);
or U3377 (N_3377,N_1135,N_1577);
nand U3378 (N_3378,N_1648,N_1014);
nand U3379 (N_3379,N_431,N_387);
xor U3380 (N_3380,N_1531,N_72);
and U3381 (N_3381,N_407,N_1212);
and U3382 (N_3382,N_869,N_1089);
or U3383 (N_3383,N_812,N_988);
nor U3384 (N_3384,N_1487,N_563);
xor U3385 (N_3385,N_960,N_660);
nand U3386 (N_3386,N_1315,N_17);
and U3387 (N_3387,N_607,N_1859);
and U3388 (N_3388,N_981,N_164);
nand U3389 (N_3389,N_149,N_368);
nor U3390 (N_3390,N_889,N_696);
nand U3391 (N_3391,N_694,N_1215);
and U3392 (N_3392,N_1436,N_1826);
nor U3393 (N_3393,N_1399,N_1866);
and U3394 (N_3394,N_698,N_1800);
nand U3395 (N_3395,N_1775,N_709);
nand U3396 (N_3396,N_1423,N_1687);
nor U3397 (N_3397,N_1055,N_295);
nand U3398 (N_3398,N_1914,N_721);
nand U3399 (N_3399,N_162,N_1627);
or U3400 (N_3400,N_475,N_692);
and U3401 (N_3401,N_1522,N_677);
or U3402 (N_3402,N_919,N_297);
or U3403 (N_3403,N_371,N_1855);
or U3404 (N_3404,N_1715,N_199);
or U3405 (N_3405,N_642,N_1299);
or U3406 (N_3406,N_1403,N_20);
and U3407 (N_3407,N_517,N_153);
xnor U3408 (N_3408,N_1434,N_280);
nor U3409 (N_3409,N_240,N_1714);
nor U3410 (N_3410,N_1022,N_426);
and U3411 (N_3411,N_1747,N_465);
nand U3412 (N_3412,N_604,N_864);
or U3413 (N_3413,N_1862,N_1395);
and U3414 (N_3414,N_883,N_1686);
nand U3415 (N_3415,N_447,N_1280);
nand U3416 (N_3416,N_1783,N_1100);
or U3417 (N_3417,N_71,N_785);
nand U3418 (N_3418,N_684,N_1311);
nor U3419 (N_3419,N_1683,N_440);
or U3420 (N_3420,N_1568,N_661);
nor U3421 (N_3421,N_1675,N_193);
or U3422 (N_3422,N_818,N_1564);
and U3423 (N_3423,N_1195,N_259);
nand U3424 (N_3424,N_1489,N_1870);
and U3425 (N_3425,N_198,N_1804);
and U3426 (N_3426,N_190,N_789);
nand U3427 (N_3427,N_154,N_523);
nor U3428 (N_3428,N_595,N_1616);
or U3429 (N_3429,N_94,N_1852);
nor U3430 (N_3430,N_1881,N_204);
nand U3431 (N_3431,N_1072,N_114);
and U3432 (N_3432,N_230,N_1469);
nand U3433 (N_3433,N_1372,N_1375);
nand U3434 (N_3434,N_1796,N_792);
xor U3435 (N_3435,N_450,N_687);
and U3436 (N_3436,N_1660,N_290);
nor U3437 (N_3437,N_817,N_220);
nand U3438 (N_3438,N_215,N_349);
nand U3439 (N_3439,N_385,N_46);
or U3440 (N_3440,N_1761,N_1036);
nor U3441 (N_3441,N_1913,N_1581);
nor U3442 (N_3442,N_731,N_990);
nor U3443 (N_3443,N_977,N_1966);
xor U3444 (N_3444,N_766,N_881);
nor U3445 (N_3445,N_1854,N_1550);
nand U3446 (N_3446,N_1980,N_820);
or U3447 (N_3447,N_1937,N_498);
and U3448 (N_3448,N_1445,N_1449);
and U3449 (N_3449,N_324,N_1679);
xor U3450 (N_3450,N_940,N_180);
nand U3451 (N_3451,N_1702,N_816);
xnor U3452 (N_3452,N_159,N_1455);
and U3453 (N_3453,N_1909,N_857);
nand U3454 (N_3454,N_405,N_223);
nor U3455 (N_3455,N_250,N_542);
and U3456 (N_3456,N_1396,N_1896);
and U3457 (N_3457,N_725,N_954);
nor U3458 (N_3458,N_1592,N_1478);
nor U3459 (N_3459,N_1743,N_792);
nor U3460 (N_3460,N_1427,N_640);
nand U3461 (N_3461,N_208,N_91);
and U3462 (N_3462,N_1293,N_173);
or U3463 (N_3463,N_1952,N_103);
nand U3464 (N_3464,N_326,N_225);
nand U3465 (N_3465,N_1682,N_419);
xnor U3466 (N_3466,N_1502,N_1944);
nand U3467 (N_3467,N_1379,N_1381);
nor U3468 (N_3468,N_880,N_1585);
xnor U3469 (N_3469,N_714,N_987);
nand U3470 (N_3470,N_733,N_1314);
nand U3471 (N_3471,N_1439,N_187);
and U3472 (N_3472,N_1882,N_12);
and U3473 (N_3473,N_690,N_751);
and U3474 (N_3474,N_134,N_828);
or U3475 (N_3475,N_1774,N_420);
nor U3476 (N_3476,N_668,N_516);
nand U3477 (N_3477,N_1323,N_170);
and U3478 (N_3478,N_1261,N_2);
and U3479 (N_3479,N_371,N_769);
and U3480 (N_3480,N_1395,N_1827);
or U3481 (N_3481,N_623,N_1736);
nand U3482 (N_3482,N_487,N_1204);
nand U3483 (N_3483,N_811,N_1075);
nor U3484 (N_3484,N_1297,N_1123);
and U3485 (N_3485,N_288,N_1918);
xor U3486 (N_3486,N_152,N_273);
nor U3487 (N_3487,N_1768,N_41);
xnor U3488 (N_3488,N_729,N_1944);
nand U3489 (N_3489,N_1758,N_1749);
nand U3490 (N_3490,N_1784,N_19);
nor U3491 (N_3491,N_154,N_301);
and U3492 (N_3492,N_522,N_462);
xor U3493 (N_3493,N_1208,N_1539);
nor U3494 (N_3494,N_448,N_530);
xor U3495 (N_3495,N_449,N_1011);
nor U3496 (N_3496,N_1754,N_558);
nor U3497 (N_3497,N_1590,N_212);
nand U3498 (N_3498,N_69,N_1842);
or U3499 (N_3499,N_955,N_264);
and U3500 (N_3500,N_1744,N_1260);
or U3501 (N_3501,N_1911,N_354);
nor U3502 (N_3502,N_1964,N_539);
nor U3503 (N_3503,N_305,N_278);
nor U3504 (N_3504,N_1204,N_1796);
nor U3505 (N_3505,N_1371,N_1630);
nand U3506 (N_3506,N_1397,N_1399);
nor U3507 (N_3507,N_1545,N_80);
or U3508 (N_3508,N_452,N_788);
nor U3509 (N_3509,N_1420,N_648);
and U3510 (N_3510,N_602,N_787);
or U3511 (N_3511,N_563,N_739);
nor U3512 (N_3512,N_797,N_1157);
nand U3513 (N_3513,N_1468,N_818);
xor U3514 (N_3514,N_433,N_145);
nand U3515 (N_3515,N_879,N_867);
or U3516 (N_3516,N_97,N_1652);
or U3517 (N_3517,N_1104,N_1651);
and U3518 (N_3518,N_978,N_56);
nor U3519 (N_3519,N_1699,N_1735);
and U3520 (N_3520,N_45,N_206);
or U3521 (N_3521,N_1566,N_1626);
or U3522 (N_3522,N_884,N_572);
nor U3523 (N_3523,N_803,N_1990);
nor U3524 (N_3524,N_773,N_1457);
nand U3525 (N_3525,N_230,N_237);
nand U3526 (N_3526,N_1175,N_1647);
and U3527 (N_3527,N_859,N_856);
nand U3528 (N_3528,N_135,N_1042);
nand U3529 (N_3529,N_1153,N_1815);
or U3530 (N_3530,N_1954,N_1466);
nor U3531 (N_3531,N_1833,N_1390);
and U3532 (N_3532,N_317,N_112);
nand U3533 (N_3533,N_1239,N_1786);
nand U3534 (N_3534,N_1701,N_559);
nor U3535 (N_3535,N_1161,N_1699);
xor U3536 (N_3536,N_1318,N_548);
xor U3537 (N_3537,N_1144,N_323);
nor U3538 (N_3538,N_84,N_604);
nand U3539 (N_3539,N_503,N_1935);
nand U3540 (N_3540,N_1100,N_1725);
nand U3541 (N_3541,N_1807,N_1551);
nand U3542 (N_3542,N_636,N_1134);
or U3543 (N_3543,N_500,N_596);
nand U3544 (N_3544,N_479,N_1545);
or U3545 (N_3545,N_16,N_89);
nand U3546 (N_3546,N_1086,N_845);
nand U3547 (N_3547,N_587,N_107);
and U3548 (N_3548,N_953,N_1372);
and U3549 (N_3549,N_719,N_1068);
or U3550 (N_3550,N_1636,N_237);
nor U3551 (N_3551,N_1945,N_1634);
and U3552 (N_3552,N_342,N_632);
and U3553 (N_3553,N_407,N_1428);
nand U3554 (N_3554,N_1692,N_1267);
or U3555 (N_3555,N_786,N_551);
nor U3556 (N_3556,N_496,N_1650);
nor U3557 (N_3557,N_138,N_1100);
xnor U3558 (N_3558,N_80,N_600);
nor U3559 (N_3559,N_514,N_1649);
nand U3560 (N_3560,N_106,N_1494);
nor U3561 (N_3561,N_698,N_1301);
nand U3562 (N_3562,N_336,N_1174);
or U3563 (N_3563,N_318,N_949);
and U3564 (N_3564,N_1148,N_1992);
and U3565 (N_3565,N_5,N_1448);
or U3566 (N_3566,N_1072,N_1365);
and U3567 (N_3567,N_1385,N_838);
nor U3568 (N_3568,N_261,N_326);
and U3569 (N_3569,N_1600,N_1908);
or U3570 (N_3570,N_343,N_229);
nor U3571 (N_3571,N_53,N_1380);
and U3572 (N_3572,N_1691,N_142);
nand U3573 (N_3573,N_810,N_1940);
nor U3574 (N_3574,N_1538,N_589);
nor U3575 (N_3575,N_1301,N_98);
and U3576 (N_3576,N_1965,N_617);
and U3577 (N_3577,N_467,N_1462);
or U3578 (N_3578,N_1336,N_1588);
nor U3579 (N_3579,N_13,N_624);
and U3580 (N_3580,N_1317,N_1120);
nand U3581 (N_3581,N_1433,N_1471);
or U3582 (N_3582,N_1870,N_166);
nor U3583 (N_3583,N_436,N_1938);
or U3584 (N_3584,N_1675,N_1862);
or U3585 (N_3585,N_78,N_256);
or U3586 (N_3586,N_569,N_975);
nor U3587 (N_3587,N_751,N_1462);
nor U3588 (N_3588,N_574,N_1740);
nand U3589 (N_3589,N_299,N_286);
and U3590 (N_3590,N_1335,N_1895);
or U3591 (N_3591,N_233,N_482);
xor U3592 (N_3592,N_1994,N_471);
nand U3593 (N_3593,N_1288,N_1320);
nor U3594 (N_3594,N_339,N_1023);
nand U3595 (N_3595,N_1486,N_1062);
nand U3596 (N_3596,N_97,N_1111);
or U3597 (N_3597,N_523,N_768);
and U3598 (N_3598,N_1957,N_926);
nand U3599 (N_3599,N_1263,N_1448);
xor U3600 (N_3600,N_1390,N_321);
nor U3601 (N_3601,N_1290,N_325);
nor U3602 (N_3602,N_1235,N_1733);
nor U3603 (N_3603,N_816,N_587);
nand U3604 (N_3604,N_1916,N_217);
xor U3605 (N_3605,N_1397,N_846);
and U3606 (N_3606,N_491,N_444);
or U3607 (N_3607,N_1454,N_838);
nor U3608 (N_3608,N_1905,N_553);
nor U3609 (N_3609,N_1176,N_36);
nand U3610 (N_3610,N_927,N_398);
and U3611 (N_3611,N_1949,N_1297);
nor U3612 (N_3612,N_1888,N_1724);
nor U3613 (N_3613,N_203,N_1840);
nor U3614 (N_3614,N_10,N_246);
or U3615 (N_3615,N_553,N_1569);
or U3616 (N_3616,N_1440,N_651);
or U3617 (N_3617,N_419,N_1329);
nand U3618 (N_3618,N_1586,N_1865);
and U3619 (N_3619,N_46,N_15);
nand U3620 (N_3620,N_40,N_912);
and U3621 (N_3621,N_1707,N_1703);
or U3622 (N_3622,N_1678,N_151);
nand U3623 (N_3623,N_676,N_240);
and U3624 (N_3624,N_1242,N_1396);
xnor U3625 (N_3625,N_1733,N_1767);
xnor U3626 (N_3626,N_601,N_130);
or U3627 (N_3627,N_44,N_1813);
nand U3628 (N_3628,N_72,N_271);
nor U3629 (N_3629,N_1174,N_208);
or U3630 (N_3630,N_411,N_1039);
nor U3631 (N_3631,N_1847,N_1524);
or U3632 (N_3632,N_1455,N_199);
and U3633 (N_3633,N_1285,N_694);
and U3634 (N_3634,N_1838,N_1655);
or U3635 (N_3635,N_1331,N_1696);
nand U3636 (N_3636,N_1742,N_413);
and U3637 (N_3637,N_1710,N_844);
nor U3638 (N_3638,N_745,N_1667);
or U3639 (N_3639,N_1095,N_839);
nand U3640 (N_3640,N_642,N_823);
nand U3641 (N_3641,N_1250,N_445);
and U3642 (N_3642,N_1484,N_1578);
nand U3643 (N_3643,N_1576,N_892);
or U3644 (N_3644,N_1113,N_276);
xor U3645 (N_3645,N_772,N_549);
and U3646 (N_3646,N_503,N_1604);
and U3647 (N_3647,N_1042,N_1950);
nor U3648 (N_3648,N_1770,N_729);
or U3649 (N_3649,N_1374,N_1485);
or U3650 (N_3650,N_1480,N_661);
and U3651 (N_3651,N_116,N_1661);
or U3652 (N_3652,N_298,N_574);
xnor U3653 (N_3653,N_370,N_1460);
or U3654 (N_3654,N_1158,N_1937);
nor U3655 (N_3655,N_1078,N_13);
nor U3656 (N_3656,N_1811,N_296);
nor U3657 (N_3657,N_1406,N_1695);
nor U3658 (N_3658,N_630,N_1481);
nor U3659 (N_3659,N_830,N_1927);
and U3660 (N_3660,N_1812,N_1090);
nand U3661 (N_3661,N_1867,N_1216);
or U3662 (N_3662,N_615,N_1192);
nand U3663 (N_3663,N_1755,N_444);
or U3664 (N_3664,N_1319,N_1831);
or U3665 (N_3665,N_776,N_353);
nand U3666 (N_3666,N_1988,N_921);
and U3667 (N_3667,N_131,N_1143);
nand U3668 (N_3668,N_674,N_576);
xor U3669 (N_3669,N_1957,N_1512);
and U3670 (N_3670,N_1967,N_1721);
nor U3671 (N_3671,N_512,N_270);
nand U3672 (N_3672,N_1245,N_1689);
and U3673 (N_3673,N_1685,N_1664);
and U3674 (N_3674,N_197,N_374);
xnor U3675 (N_3675,N_731,N_1312);
xnor U3676 (N_3676,N_785,N_962);
xnor U3677 (N_3677,N_407,N_1385);
nor U3678 (N_3678,N_1757,N_825);
nand U3679 (N_3679,N_1447,N_703);
or U3680 (N_3680,N_458,N_1263);
xor U3681 (N_3681,N_707,N_1810);
nand U3682 (N_3682,N_28,N_1982);
nand U3683 (N_3683,N_1277,N_726);
or U3684 (N_3684,N_511,N_973);
nor U3685 (N_3685,N_1414,N_712);
nand U3686 (N_3686,N_1727,N_1723);
nand U3687 (N_3687,N_229,N_1627);
nor U3688 (N_3688,N_1332,N_978);
and U3689 (N_3689,N_20,N_423);
and U3690 (N_3690,N_445,N_291);
nor U3691 (N_3691,N_1348,N_259);
nor U3692 (N_3692,N_744,N_1669);
nor U3693 (N_3693,N_673,N_428);
nor U3694 (N_3694,N_19,N_564);
xnor U3695 (N_3695,N_788,N_1634);
nor U3696 (N_3696,N_1795,N_539);
xnor U3697 (N_3697,N_352,N_1698);
nor U3698 (N_3698,N_1323,N_266);
nor U3699 (N_3699,N_995,N_1523);
nor U3700 (N_3700,N_149,N_955);
nor U3701 (N_3701,N_940,N_1541);
or U3702 (N_3702,N_815,N_1986);
and U3703 (N_3703,N_230,N_667);
or U3704 (N_3704,N_1703,N_1209);
nand U3705 (N_3705,N_28,N_223);
nor U3706 (N_3706,N_713,N_1676);
and U3707 (N_3707,N_1639,N_1011);
and U3708 (N_3708,N_1462,N_161);
and U3709 (N_3709,N_227,N_1021);
nor U3710 (N_3710,N_1361,N_768);
nand U3711 (N_3711,N_1618,N_1369);
nor U3712 (N_3712,N_84,N_747);
and U3713 (N_3713,N_1246,N_1610);
nor U3714 (N_3714,N_1361,N_1490);
xor U3715 (N_3715,N_99,N_943);
nor U3716 (N_3716,N_60,N_1259);
nor U3717 (N_3717,N_1713,N_604);
and U3718 (N_3718,N_1824,N_75);
nand U3719 (N_3719,N_797,N_1115);
nand U3720 (N_3720,N_1395,N_1075);
or U3721 (N_3721,N_521,N_1813);
xnor U3722 (N_3722,N_701,N_238);
or U3723 (N_3723,N_364,N_754);
or U3724 (N_3724,N_711,N_959);
xnor U3725 (N_3725,N_1982,N_116);
nand U3726 (N_3726,N_1212,N_975);
and U3727 (N_3727,N_1637,N_1752);
xor U3728 (N_3728,N_430,N_610);
or U3729 (N_3729,N_1401,N_1942);
nand U3730 (N_3730,N_1307,N_1640);
nor U3731 (N_3731,N_532,N_418);
and U3732 (N_3732,N_157,N_1605);
nand U3733 (N_3733,N_676,N_1260);
nand U3734 (N_3734,N_1536,N_1910);
and U3735 (N_3735,N_630,N_428);
and U3736 (N_3736,N_595,N_1981);
xnor U3737 (N_3737,N_324,N_561);
and U3738 (N_3738,N_1537,N_848);
or U3739 (N_3739,N_1423,N_928);
and U3740 (N_3740,N_963,N_1522);
xnor U3741 (N_3741,N_1343,N_1481);
nor U3742 (N_3742,N_829,N_1711);
or U3743 (N_3743,N_1697,N_797);
and U3744 (N_3744,N_1149,N_1794);
nand U3745 (N_3745,N_1450,N_51);
or U3746 (N_3746,N_204,N_1361);
or U3747 (N_3747,N_1137,N_1043);
nand U3748 (N_3748,N_28,N_798);
or U3749 (N_3749,N_725,N_1843);
nand U3750 (N_3750,N_1742,N_1695);
nand U3751 (N_3751,N_1222,N_889);
xor U3752 (N_3752,N_85,N_1327);
or U3753 (N_3753,N_1890,N_441);
or U3754 (N_3754,N_1463,N_524);
or U3755 (N_3755,N_485,N_1438);
nand U3756 (N_3756,N_1439,N_1188);
xor U3757 (N_3757,N_432,N_1987);
xor U3758 (N_3758,N_143,N_395);
xnor U3759 (N_3759,N_319,N_1763);
xnor U3760 (N_3760,N_1587,N_641);
nor U3761 (N_3761,N_1998,N_20);
or U3762 (N_3762,N_481,N_1453);
nor U3763 (N_3763,N_575,N_1536);
nor U3764 (N_3764,N_638,N_1335);
or U3765 (N_3765,N_947,N_1448);
nor U3766 (N_3766,N_879,N_1721);
nor U3767 (N_3767,N_335,N_455);
nand U3768 (N_3768,N_1787,N_51);
or U3769 (N_3769,N_655,N_1752);
xor U3770 (N_3770,N_440,N_1120);
and U3771 (N_3771,N_878,N_1723);
and U3772 (N_3772,N_279,N_998);
or U3773 (N_3773,N_964,N_930);
and U3774 (N_3774,N_1662,N_1742);
or U3775 (N_3775,N_80,N_520);
nor U3776 (N_3776,N_6,N_591);
and U3777 (N_3777,N_1209,N_1701);
or U3778 (N_3778,N_724,N_1910);
or U3779 (N_3779,N_887,N_119);
nor U3780 (N_3780,N_1424,N_1694);
nand U3781 (N_3781,N_898,N_1394);
and U3782 (N_3782,N_1260,N_1544);
or U3783 (N_3783,N_1729,N_1860);
nand U3784 (N_3784,N_316,N_1395);
nand U3785 (N_3785,N_1985,N_1979);
nand U3786 (N_3786,N_1936,N_1228);
nand U3787 (N_3787,N_791,N_580);
nor U3788 (N_3788,N_605,N_1911);
nor U3789 (N_3789,N_248,N_1882);
or U3790 (N_3790,N_673,N_371);
and U3791 (N_3791,N_1384,N_1642);
nor U3792 (N_3792,N_1233,N_1012);
xnor U3793 (N_3793,N_1823,N_685);
and U3794 (N_3794,N_490,N_657);
or U3795 (N_3795,N_1822,N_612);
and U3796 (N_3796,N_1524,N_296);
nand U3797 (N_3797,N_1781,N_1509);
nor U3798 (N_3798,N_139,N_1847);
and U3799 (N_3799,N_878,N_1624);
nand U3800 (N_3800,N_892,N_1936);
nor U3801 (N_3801,N_289,N_1356);
nand U3802 (N_3802,N_46,N_458);
and U3803 (N_3803,N_1469,N_1200);
xnor U3804 (N_3804,N_1923,N_977);
or U3805 (N_3805,N_284,N_199);
nand U3806 (N_3806,N_1280,N_1114);
or U3807 (N_3807,N_1856,N_467);
or U3808 (N_3808,N_1491,N_890);
or U3809 (N_3809,N_1079,N_198);
or U3810 (N_3810,N_328,N_1971);
nand U3811 (N_3811,N_42,N_1787);
and U3812 (N_3812,N_1211,N_1983);
nand U3813 (N_3813,N_1213,N_603);
nand U3814 (N_3814,N_103,N_416);
or U3815 (N_3815,N_1466,N_479);
nand U3816 (N_3816,N_1559,N_1348);
and U3817 (N_3817,N_955,N_635);
nand U3818 (N_3818,N_1966,N_1315);
nand U3819 (N_3819,N_663,N_65);
nand U3820 (N_3820,N_1681,N_1890);
nor U3821 (N_3821,N_1160,N_801);
or U3822 (N_3822,N_890,N_866);
xnor U3823 (N_3823,N_1944,N_1053);
xnor U3824 (N_3824,N_1008,N_1640);
nand U3825 (N_3825,N_764,N_1989);
and U3826 (N_3826,N_683,N_1071);
nand U3827 (N_3827,N_176,N_1613);
nand U3828 (N_3828,N_1252,N_228);
and U3829 (N_3829,N_1963,N_804);
nand U3830 (N_3830,N_1976,N_1440);
or U3831 (N_3831,N_380,N_854);
and U3832 (N_3832,N_1888,N_1134);
xor U3833 (N_3833,N_66,N_726);
or U3834 (N_3834,N_1506,N_869);
or U3835 (N_3835,N_291,N_1708);
or U3836 (N_3836,N_444,N_541);
or U3837 (N_3837,N_699,N_576);
nor U3838 (N_3838,N_98,N_1687);
nand U3839 (N_3839,N_1822,N_1040);
or U3840 (N_3840,N_997,N_594);
or U3841 (N_3841,N_219,N_120);
nand U3842 (N_3842,N_1146,N_492);
nand U3843 (N_3843,N_617,N_1243);
and U3844 (N_3844,N_582,N_1820);
nand U3845 (N_3845,N_1961,N_1194);
nand U3846 (N_3846,N_1313,N_1143);
nor U3847 (N_3847,N_306,N_42);
nor U3848 (N_3848,N_902,N_880);
and U3849 (N_3849,N_757,N_1224);
and U3850 (N_3850,N_276,N_187);
or U3851 (N_3851,N_205,N_1018);
and U3852 (N_3852,N_349,N_278);
nor U3853 (N_3853,N_1154,N_1725);
nand U3854 (N_3854,N_781,N_1589);
nand U3855 (N_3855,N_1017,N_293);
and U3856 (N_3856,N_1648,N_1213);
and U3857 (N_3857,N_1964,N_1499);
and U3858 (N_3858,N_1935,N_683);
and U3859 (N_3859,N_488,N_1759);
or U3860 (N_3860,N_913,N_1174);
and U3861 (N_3861,N_1571,N_268);
or U3862 (N_3862,N_340,N_392);
nor U3863 (N_3863,N_1361,N_1468);
or U3864 (N_3864,N_389,N_1637);
and U3865 (N_3865,N_1495,N_76);
or U3866 (N_3866,N_1710,N_1352);
nor U3867 (N_3867,N_242,N_455);
nand U3868 (N_3868,N_950,N_1626);
nand U3869 (N_3869,N_1285,N_783);
xnor U3870 (N_3870,N_1866,N_1314);
nand U3871 (N_3871,N_1015,N_326);
xnor U3872 (N_3872,N_32,N_1838);
and U3873 (N_3873,N_696,N_546);
nor U3874 (N_3874,N_209,N_1086);
nor U3875 (N_3875,N_26,N_1499);
nor U3876 (N_3876,N_619,N_898);
or U3877 (N_3877,N_1641,N_1911);
nor U3878 (N_3878,N_1528,N_1500);
and U3879 (N_3879,N_1667,N_1428);
nand U3880 (N_3880,N_1790,N_1910);
nand U3881 (N_3881,N_1602,N_517);
xnor U3882 (N_3882,N_529,N_279);
and U3883 (N_3883,N_1395,N_276);
or U3884 (N_3884,N_527,N_969);
and U3885 (N_3885,N_1725,N_119);
or U3886 (N_3886,N_1408,N_1986);
and U3887 (N_3887,N_1279,N_1645);
and U3888 (N_3888,N_385,N_865);
nand U3889 (N_3889,N_1387,N_428);
or U3890 (N_3890,N_1201,N_1421);
nor U3891 (N_3891,N_775,N_916);
and U3892 (N_3892,N_148,N_1825);
and U3893 (N_3893,N_490,N_1365);
nand U3894 (N_3894,N_629,N_57);
nor U3895 (N_3895,N_604,N_1548);
or U3896 (N_3896,N_487,N_1197);
nor U3897 (N_3897,N_873,N_751);
nor U3898 (N_3898,N_770,N_1977);
xnor U3899 (N_3899,N_1791,N_1507);
and U3900 (N_3900,N_1053,N_616);
xnor U3901 (N_3901,N_1239,N_606);
nand U3902 (N_3902,N_904,N_816);
and U3903 (N_3903,N_1386,N_542);
nand U3904 (N_3904,N_1978,N_925);
nor U3905 (N_3905,N_1221,N_982);
nor U3906 (N_3906,N_37,N_310);
or U3907 (N_3907,N_1939,N_1932);
or U3908 (N_3908,N_897,N_1130);
or U3909 (N_3909,N_224,N_882);
nand U3910 (N_3910,N_649,N_1904);
nor U3911 (N_3911,N_669,N_1235);
or U3912 (N_3912,N_1805,N_1701);
xor U3913 (N_3913,N_787,N_200);
and U3914 (N_3914,N_239,N_893);
xor U3915 (N_3915,N_1732,N_449);
nand U3916 (N_3916,N_1139,N_659);
nor U3917 (N_3917,N_1661,N_67);
nand U3918 (N_3918,N_660,N_1519);
nand U3919 (N_3919,N_885,N_989);
nor U3920 (N_3920,N_840,N_949);
nor U3921 (N_3921,N_922,N_731);
and U3922 (N_3922,N_1862,N_263);
nand U3923 (N_3923,N_563,N_1071);
nor U3924 (N_3924,N_1838,N_120);
nand U3925 (N_3925,N_363,N_1679);
nand U3926 (N_3926,N_1687,N_598);
or U3927 (N_3927,N_1181,N_1975);
nand U3928 (N_3928,N_1362,N_1064);
or U3929 (N_3929,N_928,N_759);
or U3930 (N_3930,N_780,N_1575);
nor U3931 (N_3931,N_1126,N_1039);
xnor U3932 (N_3932,N_1797,N_285);
and U3933 (N_3933,N_1888,N_501);
nand U3934 (N_3934,N_1368,N_672);
and U3935 (N_3935,N_1702,N_1118);
nand U3936 (N_3936,N_1404,N_1735);
or U3937 (N_3937,N_1862,N_940);
nor U3938 (N_3938,N_1391,N_985);
nor U3939 (N_3939,N_1112,N_1381);
nor U3940 (N_3940,N_1596,N_68);
nand U3941 (N_3941,N_1057,N_745);
nor U3942 (N_3942,N_4,N_1104);
or U3943 (N_3943,N_599,N_1601);
or U3944 (N_3944,N_1172,N_1474);
and U3945 (N_3945,N_1727,N_758);
nor U3946 (N_3946,N_1689,N_446);
nand U3947 (N_3947,N_965,N_1660);
or U3948 (N_3948,N_1554,N_616);
or U3949 (N_3949,N_662,N_1861);
nor U3950 (N_3950,N_330,N_220);
nand U3951 (N_3951,N_1034,N_837);
xor U3952 (N_3952,N_145,N_1580);
and U3953 (N_3953,N_1251,N_1664);
or U3954 (N_3954,N_1712,N_527);
nor U3955 (N_3955,N_1769,N_1306);
xor U3956 (N_3956,N_194,N_1890);
nand U3957 (N_3957,N_1378,N_1778);
xor U3958 (N_3958,N_1323,N_1051);
nand U3959 (N_3959,N_1453,N_1667);
and U3960 (N_3960,N_1459,N_393);
nand U3961 (N_3961,N_1179,N_1787);
or U3962 (N_3962,N_1194,N_722);
xnor U3963 (N_3963,N_1729,N_589);
xor U3964 (N_3964,N_652,N_524);
nand U3965 (N_3965,N_91,N_1482);
and U3966 (N_3966,N_90,N_276);
nor U3967 (N_3967,N_950,N_1854);
nand U3968 (N_3968,N_1532,N_489);
nand U3969 (N_3969,N_923,N_1956);
nor U3970 (N_3970,N_31,N_22);
or U3971 (N_3971,N_1873,N_1484);
and U3972 (N_3972,N_1381,N_1819);
and U3973 (N_3973,N_1011,N_995);
and U3974 (N_3974,N_87,N_1767);
and U3975 (N_3975,N_885,N_1429);
or U3976 (N_3976,N_1287,N_1811);
nand U3977 (N_3977,N_1712,N_1728);
or U3978 (N_3978,N_1749,N_277);
or U3979 (N_3979,N_138,N_1311);
nor U3980 (N_3980,N_1725,N_20);
and U3981 (N_3981,N_902,N_731);
nand U3982 (N_3982,N_356,N_109);
and U3983 (N_3983,N_314,N_1688);
xnor U3984 (N_3984,N_1959,N_1184);
and U3985 (N_3985,N_1933,N_1026);
nand U3986 (N_3986,N_882,N_718);
nand U3987 (N_3987,N_650,N_1469);
nor U3988 (N_3988,N_56,N_1106);
or U3989 (N_3989,N_1910,N_1163);
nor U3990 (N_3990,N_567,N_1173);
and U3991 (N_3991,N_1227,N_1265);
nor U3992 (N_3992,N_420,N_1807);
nor U3993 (N_3993,N_387,N_1923);
nor U3994 (N_3994,N_1852,N_595);
nand U3995 (N_3995,N_856,N_1101);
nand U3996 (N_3996,N_1576,N_1265);
or U3997 (N_3997,N_331,N_567);
or U3998 (N_3998,N_1468,N_1084);
and U3999 (N_3999,N_705,N_542);
and U4000 (N_4000,N_3730,N_2451);
nand U4001 (N_4001,N_3319,N_3809);
nand U4002 (N_4002,N_3143,N_2088);
or U4003 (N_4003,N_3772,N_3445);
and U4004 (N_4004,N_3263,N_3598);
nand U4005 (N_4005,N_3286,N_2548);
or U4006 (N_4006,N_2675,N_3641);
or U4007 (N_4007,N_2654,N_2078);
and U4008 (N_4008,N_3409,N_3656);
or U4009 (N_4009,N_3226,N_3469);
xnor U4010 (N_4010,N_2534,N_2850);
or U4011 (N_4011,N_2285,N_3278);
and U4012 (N_4012,N_3280,N_2708);
and U4013 (N_4013,N_2522,N_2752);
nand U4014 (N_4014,N_3979,N_3534);
and U4015 (N_4015,N_3491,N_3786);
xor U4016 (N_4016,N_2871,N_2460);
nor U4017 (N_4017,N_2709,N_3163);
or U4018 (N_4018,N_3905,N_3369);
nor U4019 (N_4019,N_3634,N_2583);
nand U4020 (N_4020,N_2086,N_2587);
or U4021 (N_4021,N_3745,N_3834);
nand U4022 (N_4022,N_3652,N_2818);
or U4023 (N_4023,N_3742,N_2938);
xor U4024 (N_4024,N_2765,N_3814);
nand U4025 (N_4025,N_2089,N_2431);
nand U4026 (N_4026,N_2356,N_3069);
and U4027 (N_4027,N_3014,N_3249);
or U4028 (N_4028,N_2268,N_2276);
and U4029 (N_4029,N_2710,N_3887);
and U4030 (N_4030,N_2994,N_2266);
nand U4031 (N_4031,N_3487,N_2560);
nor U4032 (N_4032,N_2726,N_2581);
nand U4033 (N_4033,N_2182,N_3894);
and U4034 (N_4034,N_2065,N_2662);
xnor U4035 (N_4035,N_3852,N_3315);
xor U4036 (N_4036,N_3031,N_3171);
and U4037 (N_4037,N_3843,N_3559);
and U4038 (N_4038,N_2097,N_3986);
nor U4039 (N_4039,N_3485,N_3855);
xor U4040 (N_4040,N_2509,N_3222);
nor U4041 (N_4041,N_2884,N_2371);
or U4042 (N_4042,N_2493,N_2364);
nor U4043 (N_4043,N_2847,N_2208);
nand U4044 (N_4044,N_2112,N_3784);
nor U4045 (N_4045,N_2976,N_2777);
and U4046 (N_4046,N_3414,N_2179);
or U4047 (N_4047,N_3845,N_3924);
nor U4048 (N_4048,N_2437,N_3696);
xnor U4049 (N_4049,N_2278,N_3618);
nor U4050 (N_4050,N_2164,N_3137);
and U4051 (N_4051,N_3350,N_3234);
and U4052 (N_4052,N_2462,N_2190);
or U4053 (N_4053,N_3704,N_3012);
nand U4054 (N_4054,N_3593,N_3099);
nand U4055 (N_4055,N_3705,N_3737);
nor U4056 (N_4056,N_3061,N_2108);
and U4057 (N_4057,N_3533,N_2554);
nor U4058 (N_4058,N_3376,N_3407);
nor U4059 (N_4059,N_2148,N_2215);
nand U4060 (N_4060,N_3346,N_3476);
nor U4061 (N_4061,N_3183,N_2690);
nor U4062 (N_4062,N_3964,N_3170);
nand U4063 (N_4063,N_2730,N_2337);
nor U4064 (N_4064,N_2012,N_3627);
xor U4065 (N_4065,N_3290,N_3220);
nand U4066 (N_4066,N_3150,N_3561);
xnor U4067 (N_4067,N_2128,N_3770);
xnor U4068 (N_4068,N_2742,N_2098);
or U4069 (N_4069,N_2645,N_2239);
and U4070 (N_4070,N_2605,N_3404);
xor U4071 (N_4071,N_2606,N_2345);
xnor U4072 (N_4072,N_3172,N_2805);
or U4073 (N_4073,N_3415,N_2433);
xnor U4074 (N_4074,N_2386,N_3366);
or U4075 (N_4075,N_2342,N_3000);
or U4076 (N_4076,N_2688,N_2323);
or U4077 (N_4077,N_2535,N_3570);
xnor U4078 (N_4078,N_2466,N_3273);
nand U4079 (N_4079,N_2205,N_3568);
nand U4080 (N_4080,N_3553,N_3307);
nand U4081 (N_4081,N_2010,N_2228);
nor U4082 (N_4082,N_3186,N_2832);
or U4083 (N_4083,N_2221,N_3755);
or U4084 (N_4084,N_3999,N_3078);
and U4085 (N_4085,N_2240,N_3914);
nor U4086 (N_4086,N_3578,N_3311);
nor U4087 (N_4087,N_2874,N_2840);
xor U4088 (N_4088,N_2019,N_3687);
and U4089 (N_4089,N_3646,N_2716);
or U4090 (N_4090,N_2826,N_2049);
and U4091 (N_4091,N_3925,N_2232);
or U4092 (N_4092,N_2326,N_2900);
or U4093 (N_4093,N_3953,N_3526);
nand U4094 (N_4094,N_2870,N_2816);
or U4095 (N_4095,N_2868,N_3289);
nor U4096 (N_4096,N_2246,N_3817);
nor U4097 (N_4097,N_3134,N_3276);
nand U4098 (N_4098,N_2695,N_3136);
and U4099 (N_4099,N_3856,N_2418);
and U4100 (N_4100,N_3810,N_2973);
xor U4101 (N_4101,N_3154,N_3668);
or U4102 (N_4102,N_2969,N_2919);
and U4103 (N_4103,N_3890,N_3522);
nor U4104 (N_4104,N_2291,N_3215);
and U4105 (N_4105,N_3565,N_3991);
or U4106 (N_4106,N_2700,N_2369);
nand U4107 (N_4107,N_2236,N_3962);
nor U4108 (N_4108,N_2833,N_2580);
nand U4109 (N_4109,N_3586,N_3402);
and U4110 (N_4110,N_2505,N_3191);
nand U4111 (N_4111,N_2125,N_2421);
nor U4112 (N_4112,N_2114,N_2811);
xnor U4113 (N_4113,N_2158,N_2821);
nor U4114 (N_4114,N_2885,N_2302);
or U4115 (N_4115,N_2389,N_3833);
or U4116 (N_4116,N_3574,N_2118);
nor U4117 (N_4117,N_2149,N_2017);
or U4118 (N_4118,N_3700,N_3601);
or U4119 (N_4119,N_3391,N_3442);
and U4120 (N_4120,N_3670,N_2497);
xnor U4121 (N_4121,N_2212,N_3217);
nor U4122 (N_4122,N_2152,N_2674);
nor U4123 (N_4123,N_3169,N_3033);
xor U4124 (N_4124,N_3081,N_3398);
and U4125 (N_4125,N_2819,N_2344);
nand U4126 (N_4126,N_3500,N_3537);
xnor U4127 (N_4127,N_2567,N_3957);
and U4128 (N_4128,N_2928,N_3348);
and U4129 (N_4129,N_2584,N_2477);
nand U4130 (N_4130,N_3096,N_2372);
nand U4131 (N_4131,N_3995,N_3201);
nand U4132 (N_4132,N_3686,N_3288);
and U4133 (N_4133,N_2672,N_3281);
nor U4134 (N_4134,N_3187,N_2090);
nand U4135 (N_4135,N_2753,N_3206);
nor U4136 (N_4136,N_3416,N_2296);
and U4137 (N_4137,N_2109,N_2363);
and U4138 (N_4138,N_3958,N_2478);
and U4139 (N_4139,N_2210,N_2775);
or U4140 (N_4140,N_3065,N_3503);
nand U4141 (N_4141,N_3071,N_3860);
nand U4142 (N_4142,N_2979,N_2604);
nor U4143 (N_4143,N_2166,N_2005);
xnor U4144 (N_4144,N_2541,N_2340);
or U4145 (N_4145,N_2234,N_3961);
and U4146 (N_4146,N_2436,N_3474);
or U4147 (N_4147,N_2521,N_2048);
and U4148 (N_4148,N_2848,N_3357);
or U4149 (N_4149,N_3279,N_2779);
nand U4150 (N_4150,N_2139,N_3417);
nand U4151 (N_4151,N_3003,N_2577);
and U4152 (N_4152,N_2898,N_2315);
xnor U4153 (N_4153,N_2008,N_2865);
nor U4154 (N_4154,N_2685,N_3254);
or U4155 (N_4155,N_2939,N_3877);
or U4156 (N_4156,N_3922,N_3753);
nor U4157 (N_4157,N_2855,N_2982);
or U4158 (N_4158,N_3535,N_2625);
nand U4159 (N_4159,N_3053,N_2718);
nor U4160 (N_4160,N_3177,N_2738);
nor U4161 (N_4161,N_3260,N_2707);
nor U4162 (N_4162,N_3316,N_3947);
nor U4163 (N_4163,N_3047,N_3883);
nand U4164 (N_4164,N_2837,N_3335);
or U4165 (N_4165,N_3589,N_3342);
or U4166 (N_4166,N_2656,N_3218);
nand U4167 (N_4167,N_2484,N_3420);
nor U4168 (N_4168,N_3899,N_3117);
and U4169 (N_4169,N_3788,N_2963);
nand U4170 (N_4170,N_2637,N_3250);
and U4171 (N_4171,N_3607,N_3910);
and U4172 (N_4172,N_2474,N_2209);
nand U4173 (N_4173,N_3956,N_3926);
and U4174 (N_4174,N_3089,N_3977);
or U4175 (N_4175,N_3198,N_3681);
nor U4176 (N_4176,N_2585,N_3354);
nand U4177 (N_4177,N_3966,N_3666);
nand U4178 (N_4178,N_3327,N_2183);
and U4179 (N_4179,N_2031,N_2788);
nor U4180 (N_4180,N_3841,N_3643);
nand U4181 (N_4181,N_2683,N_2551);
or U4182 (N_4182,N_2076,N_2988);
and U4183 (N_4183,N_3517,N_2122);
nand U4184 (N_4184,N_2443,N_2132);
nand U4185 (N_4185,N_2274,N_3543);
or U4186 (N_4186,N_3981,N_2957);
and U4187 (N_4187,N_2385,N_2888);
nor U4188 (N_4188,N_3195,N_3903);
nand U4189 (N_4189,N_3378,N_2754);
or U4190 (N_4190,N_3028,N_3359);
or U4191 (N_4191,N_3963,N_2129);
and U4192 (N_4192,N_3938,N_2487);
xor U4193 (N_4193,N_2666,N_2664);
and U4194 (N_4194,N_3111,N_2721);
and U4195 (N_4195,N_2226,N_3868);
or U4196 (N_4196,N_2354,N_2223);
xor U4197 (N_4197,N_2184,N_2697);
and U4198 (N_4198,N_3572,N_3757);
xor U4199 (N_4199,N_3236,N_2679);
or U4200 (N_4200,N_2127,N_3155);
or U4201 (N_4201,N_3913,N_3902);
nand U4202 (N_4202,N_3243,N_2773);
and U4203 (N_4203,N_2877,N_2021);
nand U4204 (N_4204,N_3489,N_3318);
xor U4205 (N_4205,N_2636,N_2768);
nor U4206 (N_4206,N_2055,N_3984);
or U4207 (N_4207,N_3383,N_3095);
or U4208 (N_4208,N_2760,N_3723);
and U4209 (N_4209,N_2862,N_2929);
and U4210 (N_4210,N_3308,N_3261);
or U4211 (N_4211,N_3408,N_3653);
nand U4212 (N_4212,N_3613,N_3472);
xnor U4213 (N_4213,N_3557,N_2204);
nand U4214 (N_4214,N_3508,N_2859);
and U4215 (N_4215,N_2176,N_2244);
nor U4216 (N_4216,N_2440,N_3412);
nor U4217 (N_4217,N_2990,N_3405);
nand U4218 (N_4218,N_2741,N_2943);
nand U4219 (N_4219,N_2542,N_2197);
nand U4220 (N_4220,N_3693,N_2039);
nor U4221 (N_4221,N_2022,N_2357);
and U4222 (N_4222,N_2838,N_2147);
or U4223 (N_4223,N_3101,N_2468);
and U4224 (N_4224,N_2347,N_2573);
nand U4225 (N_4225,N_3066,N_3840);
xor U4226 (N_4226,N_3050,N_2196);
xor U4227 (N_4227,N_3264,N_3235);
and U4228 (N_4228,N_2332,N_2875);
xnor U4229 (N_4229,N_3796,N_2959);
xnor U4230 (N_4230,N_2564,N_3556);
nand U4231 (N_4231,N_3462,N_3889);
xnor U4232 (N_4232,N_3725,N_3949);
or U4233 (N_4233,N_3683,N_3942);
or U4234 (N_4234,N_3648,N_2457);
xor U4235 (N_4235,N_3313,N_2558);
and U4236 (N_4236,N_2131,N_3118);
xnor U4237 (N_4237,N_2829,N_3265);
and U4238 (N_4238,N_2661,N_2787);
and U4239 (N_4239,N_2782,N_2277);
xor U4240 (N_4240,N_3591,N_3758);
xnor U4241 (N_4241,N_3312,N_2627);
and U4242 (N_4242,N_3042,N_2382);
nor U4243 (N_4243,N_2539,N_3709);
and U4244 (N_4244,N_3621,N_3021);
nor U4245 (N_4245,N_2294,N_2745);
nor U4246 (N_4246,N_3100,N_3457);
nor U4247 (N_4247,N_3923,N_2060);
nor U4248 (N_4248,N_2219,N_3002);
or U4249 (N_4249,N_2639,N_3630);
nor U4250 (N_4250,N_2248,N_2105);
and U4251 (N_4251,N_3030,N_2593);
nand U4252 (N_4252,N_3478,N_2781);
and U4253 (N_4253,N_2714,N_3427);
nor U4254 (N_4254,N_3600,N_2849);
nor U4255 (N_4255,N_3285,N_3739);
nand U4256 (N_4256,N_2992,N_3777);
nand U4257 (N_4257,N_3389,N_3639);
nor U4258 (N_4258,N_3023,N_2189);
and U4259 (N_4259,N_2794,N_2202);
or U4260 (N_4260,N_2673,N_3616);
nor U4261 (N_4261,N_2002,N_2691);
and U4262 (N_4262,N_3452,N_3716);
and U4263 (N_4263,N_3955,N_2698);
and U4264 (N_4264,N_2694,N_2866);
and U4265 (N_4265,N_3365,N_2603);
or U4266 (N_4266,N_2793,N_3514);
nor U4267 (N_4267,N_2009,N_3707);
nand U4268 (N_4268,N_2596,N_2759);
and U4269 (N_4269,N_3988,N_3467);
nor U4270 (N_4270,N_3767,N_3256);
nand U4271 (N_4271,N_3878,N_2056);
nand U4272 (N_4272,N_2744,N_2425);
nor U4273 (N_4273,N_2815,N_2452);
nor U4274 (N_4274,N_3818,N_2376);
xor U4275 (N_4275,N_3084,N_3300);
nor U4276 (N_4276,N_2544,N_2409);
xor U4277 (N_4277,N_2318,N_3004);
or U4278 (N_4278,N_3037,N_3481);
and U4279 (N_4279,N_3624,N_3258);
and U4280 (N_4280,N_2878,N_3917);
nor U4281 (N_4281,N_3293,N_2496);
nor U4282 (N_4282,N_2860,N_2731);
xor U4283 (N_4283,N_2613,N_2073);
nand U4284 (N_4284,N_3048,N_2093);
nor U4285 (N_4285,N_3347,N_3864);
nor U4286 (N_4286,N_3129,N_3204);
and U4287 (N_4287,N_2918,N_2934);
and U4288 (N_4288,N_3328,N_3985);
and U4289 (N_4289,N_2358,N_3178);
nand U4290 (N_4290,N_3588,N_3733);
nor U4291 (N_4291,N_2915,N_2499);
nor U4292 (N_4292,N_2589,N_3382);
and U4293 (N_4293,N_3199,N_2966);
nor U4294 (N_4294,N_3944,N_2640);
or U4295 (N_4295,N_3580,N_2444);
and U4296 (N_4296,N_3623,N_2750);
nand U4297 (N_4297,N_2485,N_3240);
xor U4298 (N_4298,N_3654,N_2776);
or U4299 (N_4299,N_3713,N_3872);
or U4300 (N_4300,N_3918,N_2789);
nor U4301 (N_4301,N_3244,N_3203);
xnor U4302 (N_4302,N_3519,N_2586);
nand U4303 (N_4303,N_3384,N_2936);
xnor U4304 (N_4304,N_2599,N_3025);
or U4305 (N_4305,N_2876,N_3035);
nor U4306 (N_4306,N_2308,N_3524);
nand U4307 (N_4307,N_2813,N_3443);
or U4308 (N_4308,N_3682,N_2727);
nand U4309 (N_4309,N_3688,N_2797);
nand U4310 (N_4310,N_3976,N_3388);
or U4311 (N_4311,N_3850,N_2163);
and U4312 (N_4312,N_2441,N_2703);
or U4313 (N_4313,N_3060,N_3403);
and U4314 (N_4314,N_2104,N_2540);
or U4315 (N_4315,N_2846,N_3946);
and U4316 (N_4316,N_2671,N_3464);
nand U4317 (N_4317,N_2379,N_3536);
nor U4318 (N_4318,N_3827,N_3680);
xor U4319 (N_4319,N_2766,N_3912);
or U4320 (N_4320,N_3743,N_2311);
or U4321 (N_4321,N_2882,N_2167);
and U4322 (N_4322,N_2912,N_3213);
or U4323 (N_4323,N_2217,N_3451);
nor U4324 (N_4324,N_3920,N_3396);
nor U4325 (N_4325,N_2297,N_3941);
or U4326 (N_4326,N_2159,N_3715);
nor U4327 (N_4327,N_3631,N_2545);
nor U4328 (N_4328,N_2728,N_2375);
and U4329 (N_4329,N_3530,N_2141);
or U4330 (N_4330,N_2486,N_2033);
nand U4331 (N_4331,N_2456,N_2284);
nand U4332 (N_4332,N_2942,N_2635);
nor U4333 (N_4333,N_3741,N_3675);
nand U4334 (N_4334,N_3016,N_2602);
nor U4335 (N_4335,N_2961,N_3728);
nor U4336 (N_4336,N_2761,N_2153);
nor U4337 (N_4337,N_2538,N_2503);
nand U4338 (N_4338,N_3992,N_2051);
nor U4339 (N_4339,N_3651,N_3246);
nor U4340 (N_4340,N_2434,N_2758);
nor U4341 (N_4341,N_2746,N_3554);
nand U4342 (N_4342,N_2867,N_3107);
nand U4343 (N_4343,N_2299,N_3305);
or U4344 (N_4344,N_3124,N_3615);
and U4345 (N_4345,N_3657,N_3783);
or U4346 (N_4346,N_2422,N_3635);
and U4347 (N_4347,N_2450,N_2306);
nor U4348 (N_4348,N_3584,N_3710);
or U4349 (N_4349,N_2615,N_2138);
or U4350 (N_4350,N_3038,N_2956);
or U4351 (N_4351,N_2520,N_3766);
nor U4352 (N_4352,N_2040,N_2999);
nand U4353 (N_4353,N_2381,N_2997);
xor U4354 (N_4354,N_2619,N_2643);
or U4355 (N_4355,N_3711,N_2186);
nand U4356 (N_4356,N_2445,N_3229);
nand U4357 (N_4357,N_3330,N_3399);
nand U4358 (N_4358,N_2388,N_3599);
or U4359 (N_4359,N_2135,N_3055);
nand U4360 (N_4360,N_3987,N_3665);
nand U4361 (N_4361,N_2262,N_3774);
nand U4362 (N_4362,N_3475,N_2926);
nor U4363 (N_4363,N_2067,N_2400);
or U4364 (N_4364,N_2028,N_3794);
and U4365 (N_4365,N_3950,N_3067);
or U4366 (N_4366,N_2955,N_3802);
or U4367 (N_4367,N_3994,N_2792);
nor U4368 (N_4368,N_2336,N_2095);
nor U4369 (N_4369,N_3232,N_3671);
or U4370 (N_4370,N_3406,N_2494);
and U4371 (N_4371,N_2143,N_3622);
nor U4372 (N_4372,N_2526,N_3769);
xnor U4373 (N_4373,N_2480,N_2804);
or U4374 (N_4374,N_2279,N_2629);
and U4375 (N_4375,N_2686,N_2074);
nand U4376 (N_4376,N_3862,N_3142);
or U4377 (N_4377,N_2230,N_3433);
and U4378 (N_4378,N_2140,N_2803);
or U4379 (N_4379,N_2638,N_3068);
or U4380 (N_4380,N_3619,N_2465);
xor U4381 (N_4381,N_2180,N_3642);
nor U4382 (N_4382,N_3585,N_3441);
or U4383 (N_4383,N_3094,N_3768);
and U4384 (N_4384,N_3965,N_3190);
nor U4385 (N_4385,N_2907,N_3857);
nor U4386 (N_4386,N_3807,N_3393);
or U4387 (N_4387,N_2631,N_2996);
or U4388 (N_4388,N_3041,N_2647);
xnor U4389 (N_4389,N_2853,N_3131);
and U4390 (N_4390,N_3270,N_2975);
or U4391 (N_4391,N_3908,N_2628);
nor U4392 (N_4392,N_2339,N_3039);
and U4393 (N_4393,N_3617,N_3760);
and U4394 (N_4394,N_2237,N_2762);
nand U4395 (N_4395,N_3801,N_3331);
nor U4396 (N_4396,N_3001,N_3560);
nor U4397 (N_4397,N_3013,N_3844);
and U4398 (N_4398,N_3080,N_2071);
nor U4399 (N_4399,N_3130,N_3812);
nor U4400 (N_4400,N_2784,N_3242);
nor U4401 (N_4401,N_3156,N_3302);
xnor U4402 (N_4402,N_2275,N_3811);
nor U4403 (N_4403,N_2570,N_3245);
or U4404 (N_4404,N_2978,N_2331);
nand U4405 (N_4405,N_3400,N_3509);
and U4406 (N_4406,N_3044,N_3090);
nor U4407 (N_4407,N_2003,N_2851);
and U4408 (N_4408,N_2007,N_2533);
xor U4409 (N_4409,N_3248,N_3377);
nor U4410 (N_4410,N_3729,N_3531);
nand U4411 (N_4411,N_3563,N_2319);
nand U4412 (N_4412,N_2927,N_3749);
nand U4413 (N_4413,N_3967,N_3892);
nor U4414 (N_4414,N_3835,N_3940);
and U4415 (N_4415,N_2968,N_3506);
or U4416 (N_4416,N_2949,N_2903);
xor U4417 (N_4417,N_2508,N_3180);
xnor U4418 (N_4418,N_2858,N_3983);
nor U4419 (N_4419,N_2207,N_2250);
nor U4420 (N_4420,N_3461,N_3609);
and U4421 (N_4421,N_2998,N_3571);
nand U4422 (N_4422,N_2026,N_3724);
or U4423 (N_4423,N_2165,N_3861);
nor U4424 (N_4424,N_3933,N_3230);
or U4425 (N_4425,N_3006,N_3971);
nor U4426 (N_4426,N_2507,N_2655);
or U4427 (N_4427,N_2490,N_3465);
nor U4428 (N_4428,N_2660,N_2359);
nand U4429 (N_4429,N_3297,N_3603);
nor U4430 (N_4430,N_3064,N_3109);
nand U4431 (N_4431,N_3336,N_3120);
or U4432 (N_4432,N_2195,N_2301);
nor U4433 (N_4433,N_3320,N_3027);
nand U4434 (N_4434,N_2038,N_2527);
or U4435 (N_4435,N_3368,N_3110);
and U4436 (N_4436,N_2702,N_2313);
nand U4437 (N_4437,N_3424,N_3735);
nand U4438 (N_4438,N_3092,N_2027);
or U4439 (N_4439,N_3998,N_2608);
or U4440 (N_4440,N_2470,N_2047);
and U4441 (N_4441,N_3401,N_3052);
and U4442 (N_4442,N_2783,N_2489);
or U4443 (N_4443,N_3604,N_2562);
or U4444 (N_4444,N_3825,N_3885);
nand U4445 (N_4445,N_3018,N_3165);
or U4446 (N_4446,N_3162,N_2940);
or U4447 (N_4447,N_3024,N_3516);
nand U4448 (N_4448,N_3765,N_3435);
or U4449 (N_4449,N_3262,N_3849);
nor U4450 (N_4450,N_3838,N_2293);
nor U4451 (N_4451,N_3492,N_2036);
and U4452 (N_4452,N_3972,N_3829);
nor U4453 (N_4453,N_3712,N_3214);
and U4454 (N_4454,N_2133,N_3164);
or U4455 (N_4455,N_3748,N_3296);
xnor U4456 (N_4456,N_3911,N_3138);
or U4457 (N_4457,N_3070,N_2150);
or U4458 (N_4458,N_2516,N_2397);
or U4459 (N_4459,N_2571,N_2680);
nand U4460 (N_4460,N_3460,N_3869);
or U4461 (N_4461,N_2050,N_3939);
nor U4462 (N_4462,N_2100,N_3421);
nand U4463 (N_4463,N_2475,N_3793);
or U4464 (N_4464,N_2964,N_3114);
nor U4465 (N_4465,N_2993,N_2252);
or U4466 (N_4466,N_2018,N_3895);
and U4467 (N_4467,N_2384,N_2199);
nor U4468 (N_4468,N_2235,N_3751);
or U4469 (N_4469,N_3523,N_3605);
nand U4470 (N_4470,N_2667,N_2528);
and U4471 (N_4471,N_3773,N_2600);
and U4472 (N_4472,N_2622,N_2177);
or U4473 (N_4473,N_3390,N_2426);
nand U4474 (N_4474,N_3626,N_3790);
and U4475 (N_4475,N_3370,N_2304);
nand U4476 (N_4476,N_3372,N_3754);
nand U4477 (N_4477,N_2170,N_2251);
nand U4478 (N_4478,N_3238,N_2825);
or U4479 (N_4479,N_2904,N_2430);
xor U4480 (N_4480,N_3132,N_3529);
nor U4481 (N_4481,N_2561,N_2264);
nor U4482 (N_4482,N_2392,N_3805);
nor U4483 (N_4483,N_3160,N_2734);
or U4484 (N_4484,N_3397,N_2053);
nor U4485 (N_4485,N_2864,N_3542);
nor U4486 (N_4486,N_2061,N_3550);
and U4487 (N_4487,N_3847,N_3640);
nor U4488 (N_4488,N_3510,N_2749);
nor U4489 (N_4489,N_2514,N_2863);
nand U4490 (N_4490,N_3009,N_2383);
nand U4491 (N_4491,N_3952,N_3361);
nor U4492 (N_4492,N_2947,N_2258);
and U4493 (N_4493,N_2501,N_2529);
nand U4494 (N_4494,N_3448,N_3928);
nor U4495 (N_4495,N_2481,N_3326);
nor U4496 (N_4496,N_2933,N_2764);
or U4497 (N_4497,N_2249,N_2404);
or U4498 (N_4498,N_2420,N_3973);
nand U4499 (N_4499,N_2856,N_3022);
and U4500 (N_4500,N_3655,N_3431);
nand U4501 (N_4501,N_2387,N_3821);
nand U4502 (N_4502,N_3853,N_3698);
nor U4503 (N_4503,N_3252,N_3919);
or U4504 (N_4504,N_2188,N_2395);
and U4505 (N_4505,N_2041,N_2836);
nor U4506 (N_4506,N_3674,N_2448);
and U4507 (N_4507,N_2830,N_2471);
nor U4508 (N_4508,N_3188,N_3468);
nand U4509 (N_4509,N_3780,N_3123);
and U4510 (N_4510,N_2663,N_3969);
xnor U4511 (N_4511,N_2909,N_3867);
xnor U4512 (N_4512,N_2068,N_2231);
or U4513 (N_4513,N_2890,N_2715);
nor U4514 (N_4514,N_2717,N_3893);
xor U4515 (N_4515,N_3210,N_3819);
and U4516 (N_4516,N_2417,N_2706);
nand U4517 (N_4517,N_2442,N_3555);
and U4518 (N_4518,N_2644,N_3564);
or U4519 (N_4519,N_2206,N_2362);
or U4520 (N_4520,N_3043,N_3239);
nor U4521 (N_4521,N_2980,N_2399);
or U4522 (N_4522,N_2873,N_3929);
nand U4523 (N_4523,N_2439,N_2595);
or U4524 (N_4524,N_3882,N_3225);
and U4525 (N_4525,N_3881,N_3192);
and U4526 (N_4526,N_3158,N_3521);
or U4527 (N_4527,N_3051,N_2312);
or U4528 (N_4528,N_2157,N_3722);
and U4529 (N_4529,N_2083,N_3358);
nor U4530 (N_4530,N_3590,N_3690);
or U4531 (N_4531,N_2737,N_2069);
nor U4532 (N_4532,N_2582,N_3951);
and U4533 (N_4533,N_2592,N_3450);
or U4534 (N_4534,N_3413,N_3996);
nand U4535 (N_4535,N_3104,N_3551);
and U4536 (N_4536,N_3685,N_2500);
nand U4537 (N_4537,N_3493,N_2006);
nor U4538 (N_4538,N_2124,N_2446);
nand U4539 (N_4539,N_2974,N_3495);
and U4540 (N_4540,N_2908,N_2123);
and U4541 (N_4541,N_3205,N_3746);
xor U4542 (N_4542,N_2659,N_2316);
or U4543 (N_4543,N_2879,N_3703);
and U4544 (N_4544,N_2214,N_3144);
nor U4545 (N_4545,N_2348,N_2739);
nand U4546 (N_4546,N_2515,N_3959);
nor U4547 (N_4547,N_2736,N_2724);
and U4548 (N_4548,N_2923,N_3738);
or U4549 (N_4549,N_3632,N_2591);
xnor U4550 (N_4550,N_2944,N_2822);
or U4551 (N_4551,N_3636,N_3673);
and U4552 (N_4552,N_2780,N_2227);
and U4553 (N_4553,N_3692,N_2705);
and U4554 (N_4554,N_2925,N_3058);
nand U4555 (N_4555,N_3119,N_2029);
or U4556 (N_4556,N_3614,N_2220);
nor U4557 (N_4557,N_2578,N_2416);
or U4558 (N_4558,N_3828,N_2886);
and U4559 (N_4559,N_3334,N_2984);
xnor U4560 (N_4560,N_2537,N_3638);
nor U4561 (N_4561,N_3989,N_3216);
nor U4562 (N_4562,N_2755,N_3539);
xor U4563 (N_4563,N_3778,N_3019);
nand U4564 (N_4564,N_2075,N_2064);
or U4565 (N_4565,N_3720,N_2620);
nand U4566 (N_4566,N_2000,N_3787);
and U4567 (N_4567,N_2081,N_3504);
and U4568 (N_4568,N_3432,N_2785);
nor U4569 (N_4569,N_2314,N_3582);
nand U4570 (N_4570,N_3221,N_3436);
or U4571 (N_4571,N_2621,N_3494);
and U4572 (N_4572,N_2004,N_2913);
nor U4573 (N_4573,N_2626,N_3083);
and U4574 (N_4574,N_3410,N_3549);
or U4575 (N_4575,N_2265,N_3317);
or U4576 (N_4576,N_3934,N_2820);
and U4577 (N_4577,N_2786,N_3367);
and U4578 (N_4578,N_2633,N_3993);
and U4579 (N_4579,N_2511,N_2914);
or U4580 (N_4580,N_2701,N_2532);
xnor U4581 (N_4581,N_2035,N_3102);
nor U4582 (N_4582,N_2365,N_3792);
and U4583 (N_4583,N_2971,N_3146);
or U4584 (N_4584,N_2648,N_2895);
nor U4585 (N_4585,N_2099,N_3063);
and U4586 (N_4586,N_2906,N_3870);
or U4587 (N_4587,N_3562,N_2046);
xor U4588 (N_4588,N_2831,N_3566);
or U4589 (N_4589,N_2651,N_3798);
or U4590 (N_4590,N_3085,N_3121);
nor U4591 (N_4591,N_3149,N_2676);
nand U4592 (N_4592,N_3185,N_3437);
and U4593 (N_4593,N_3046,N_2255);
xor U4594 (N_4594,N_3233,N_2463);
xnor U4595 (N_4595,N_3482,N_3439);
and U4596 (N_4596,N_2267,N_3816);
nor U4597 (N_4597,N_2343,N_2632);
and U4598 (N_4598,N_3804,N_3502);
nand U4599 (N_4599,N_3597,N_3228);
nor U4600 (N_4600,N_3789,N_3785);
and U4601 (N_4601,N_3647,N_2597);
and U4602 (N_4602,N_2617,N_2044);
nor U4603 (N_4603,N_3438,N_2225);
and U4604 (N_4604,N_3884,N_3837);
and U4605 (N_4605,N_3718,N_2115);
nor U4606 (N_4606,N_3936,N_3251);
nor U4607 (N_4607,N_2950,N_2052);
and U4608 (N_4608,N_2402,N_2747);
and U4609 (N_4609,N_3343,N_2174);
nor U4610 (N_4610,N_2238,N_2070);
nor U4611 (N_4611,N_2953,N_2960);
xor U4612 (N_4612,N_2325,N_2598);
and U4613 (N_4613,N_2366,N_3392);
or U4614 (N_4614,N_2795,N_3795);
nor U4615 (N_4615,N_2333,N_3105);
nor U4616 (N_4616,N_3677,N_3909);
nand U4617 (N_4617,N_2324,N_3077);
nor U4618 (N_4618,N_3363,N_2023);
nor U4619 (N_4619,N_2320,N_2809);
nor U4620 (N_4620,N_3449,N_3322);
and U4621 (N_4621,N_3611,N_3112);
and U4622 (N_4622,N_2552,N_3488);
or U4623 (N_4623,N_3208,N_2175);
or U4624 (N_4624,N_2142,N_2790);
or U4625 (N_4625,N_2305,N_3362);
nor U4626 (N_4626,N_3813,N_2130);
and U4627 (N_4627,N_2941,N_2889);
nor U4628 (N_4628,N_2733,N_2117);
or U4629 (N_4629,N_3227,N_3587);
and U4630 (N_4630,N_2770,N_3483);
xnor U4631 (N_4631,N_3511,N_2271);
or U4632 (N_4632,N_3701,N_2510);
nor U4633 (N_4633,N_3931,N_3595);
nand U4634 (N_4634,N_3166,N_2612);
nor U4635 (N_4635,N_2827,N_2396);
and U4636 (N_4636,N_2213,N_3193);
xor U4637 (N_4637,N_3823,N_3797);
nand U4638 (N_4638,N_3567,N_2835);
nor U4639 (N_4639,N_3072,N_3133);
xnor U4640 (N_4640,N_2492,N_2245);
nor U4641 (N_4641,N_2289,N_2247);
and U4642 (N_4642,N_3501,N_3292);
nor U4643 (N_4643,N_2473,N_2986);
and U4644 (N_4644,N_2203,N_2300);
or U4645 (N_4645,N_3697,N_3419);
or U4646 (N_4646,N_3341,N_3323);
nand U4647 (N_4647,N_2341,N_3576);
nor U4648 (N_4648,N_2924,N_2920);
xor U4649 (N_4649,N_3541,N_2161);
and U4650 (N_4650,N_2801,N_3310);
or U4651 (N_4651,N_3059,N_3338);
or U4652 (N_4652,N_2774,N_3997);
nand U4653 (N_4653,N_2464,N_2910);
and U4654 (N_4654,N_3694,N_2899);
and U4655 (N_4655,N_3202,N_2634);
or U4656 (N_4656,N_2557,N_2374);
nor U4657 (N_4657,N_3148,N_3219);
or U4658 (N_4658,N_3815,N_2461);
nor U4659 (N_4659,N_3458,N_2932);
xor U4660 (N_4660,N_2317,N_3126);
and U4661 (N_4661,N_3459,N_2699);
and U4662 (N_4662,N_3086,N_2410);
or U4663 (N_4663,N_2224,N_3394);
or U4664 (N_4664,N_3426,N_3904);
and U4665 (N_4665,N_2429,N_2732);
and U4666 (N_4666,N_2287,N_3345);
nor U4667 (N_4667,N_3649,N_2653);
or U4668 (N_4668,N_3268,N_2346);
or U4669 (N_4669,N_2751,N_3321);
or U4670 (N_4670,N_2151,N_2677);
xor U4671 (N_4671,N_3168,N_3153);
or U4672 (N_4672,N_3669,N_3224);
xnor U4673 (N_4673,N_3056,N_2704);
nor U4674 (N_4674,N_2987,N_2034);
or U4675 (N_4675,N_2281,N_2390);
nand U4676 (N_4676,N_2513,N_2665);
xnor U4677 (N_4677,N_2901,N_2309);
nor U4678 (N_4678,N_2310,N_3282);
nor U4679 (N_4679,N_2504,N_2576);
xor U4680 (N_4680,N_2995,N_2771);
and U4681 (N_4681,N_2911,N_3515);
nor U4682 (N_4682,N_2772,N_2373);
or U4683 (N_4683,N_3116,N_3267);
or U4684 (N_4684,N_3625,N_2432);
and U4685 (N_4685,N_2458,N_2769);
or U4686 (N_4686,N_2260,N_3891);
and U4687 (N_4687,N_2330,N_2016);
nor U4688 (N_4688,N_2218,N_3339);
and U4689 (N_4689,N_3147,N_3179);
nor U4690 (N_4690,N_3633,N_2917);
nand U4691 (N_4691,N_2546,N_3662);
nand U4692 (N_4692,N_2173,N_3381);
nand U4693 (N_4693,N_2024,N_2869);
and U4694 (N_4694,N_2192,N_3507);
nor U4695 (N_4695,N_2512,N_3866);
xnor U4696 (N_4696,N_2351,N_2292);
xor U4697 (N_4697,N_3152,N_3411);
nor U4698 (N_4698,N_2307,N_3091);
or U4699 (N_4699,N_3763,N_3842);
or U4700 (N_4700,N_2327,N_2828);
nor U4701 (N_4701,N_3937,N_3552);
xnor U4702 (N_4702,N_3295,N_3271);
or U4703 (N_4703,N_2172,N_3900);
or U4704 (N_4704,N_3098,N_2216);
and U4705 (N_4705,N_2958,N_3272);
and U4706 (N_4706,N_3699,N_2970);
and U4707 (N_4707,N_3752,N_2438);
or U4708 (N_4708,N_2322,N_3212);
xor U4709 (N_4709,N_3518,N_3645);
nand U4710 (N_4710,N_3846,N_2014);
and U4711 (N_4711,N_2242,N_3540);
and U4712 (N_4712,N_3283,N_3596);
and U4713 (N_4713,N_3499,N_3975);
nor U4714 (N_4714,N_2110,N_2162);
nor U4715 (N_4715,N_2280,N_2403);
nor U4716 (N_4716,N_2082,N_3008);
nor U4717 (N_4717,N_3606,N_2459);
or U4718 (N_4718,N_3097,N_2178);
xnor U4719 (N_4719,N_3269,N_2549);
xnor U4720 (N_4720,N_3371,N_3594);
or U4721 (N_4721,N_3294,N_3906);
and U4722 (N_4722,N_2854,N_3005);
or U4723 (N_4723,N_3299,N_3527);
nand U4724 (N_4724,N_2967,N_3253);
nor U4725 (N_4725,N_2349,N_3017);
xnor U4726 (N_4726,N_3211,N_3106);
xor U4727 (N_4727,N_2411,N_3423);
and U4728 (N_4728,N_3970,N_2807);
nor U4729 (N_4729,N_2491,N_3759);
nor U4730 (N_4730,N_2763,N_2286);
nand U4731 (N_4731,N_2556,N_2063);
nor U4732 (N_4732,N_2334,N_3678);
nor U4733 (N_4733,N_2712,N_3447);
or U4734 (N_4734,N_2469,N_3174);
nand U4735 (N_4735,N_3980,N_3546);
nand U4736 (N_4736,N_2618,N_3836);
and U4737 (N_4737,N_3418,N_3380);
nand U4738 (N_4738,N_2880,N_2616);
xnor U4739 (N_4739,N_2412,N_2530);
nand U4740 (N_4740,N_2256,N_2455);
or U4741 (N_4741,N_3125,N_2200);
nand U4742 (N_4742,N_2106,N_3429);
xor U4743 (N_4743,N_3954,N_3548);
or U4744 (N_4744,N_2930,N_3874);
nor U4745 (N_4745,N_3583,N_3352);
nand U4746 (N_4746,N_3806,N_3822);
nor U4747 (N_4747,N_2559,N_2335);
and U4748 (N_4748,N_2650,N_3127);
nand U4749 (N_4749,N_3344,N_2193);
or U4750 (N_4750,N_2611,N_3650);
xnor U4751 (N_4751,N_3573,N_2590);
nor U4752 (N_4752,N_2453,N_3455);
nand U4753 (N_4753,N_2896,N_3161);
nand U4754 (N_4754,N_3775,N_2181);
nor U4755 (N_4755,N_2488,N_2985);
xor U4756 (N_4756,N_2566,N_2091);
nor U4757 (N_4757,N_3247,N_2134);
and U4758 (N_4758,N_3329,N_3880);
and U4759 (N_4759,N_2609,N_2338);
nor U4760 (N_4760,N_3054,N_2791);
and U4761 (N_4761,N_3181,N_3497);
nand U4762 (N_4762,N_2107,N_2624);
nand U4763 (N_4763,N_3628,N_2054);
xor U4764 (N_4764,N_2020,N_2945);
or U4765 (N_4765,N_3440,N_3486);
nand U4766 (N_4766,N_3848,N_2435);
nor U4767 (N_4767,N_2575,N_2424);
and U4768 (N_4768,N_2922,N_3139);
nor U4769 (N_4769,N_3360,N_3151);
and U4770 (N_4770,N_3714,N_3706);
xor U4771 (N_4771,N_2298,N_3761);
and U4772 (N_4772,N_3799,N_2015);
nand U4773 (N_4773,N_3921,N_2057);
nand U4774 (N_4774,N_3672,N_3620);
xor U4775 (N_4775,N_3886,N_3176);
and U4776 (N_4776,N_3088,N_2419);
and U4777 (N_4777,N_2729,N_2991);
xnor U4778 (N_4778,N_2670,N_2693);
nand U4779 (N_4779,N_3932,N_2187);
nand U4780 (N_4780,N_2948,N_3479);
nor U4781 (N_4781,N_3333,N_2144);
and U4782 (N_4782,N_3782,N_2935);
xnor U4783 (N_4783,N_2059,N_2668);
or U4784 (N_4784,N_2146,N_2723);
and U4785 (N_4785,N_2011,N_2579);
nor U4786 (N_4786,N_2657,N_3140);
nand U4787 (N_4787,N_2547,N_2946);
or U4788 (N_4788,N_3477,N_2519);
nor U4789 (N_4789,N_2120,N_3658);
and U4790 (N_4790,N_3664,N_2812);
nor U4791 (N_4791,N_3879,N_2902);
nor U4792 (N_4792,N_2843,N_3351);
nand U4793 (N_4793,N_3901,N_3898);
xor U4794 (N_4794,N_3087,N_3851);
or U4795 (N_4795,N_2937,N_3740);
and U4796 (N_4796,N_2852,N_2735);
and U4797 (N_4797,N_2360,N_3076);
or U4798 (N_4798,N_2642,N_3237);
or U4799 (N_4799,N_3691,N_2623);
xor U4800 (N_4800,N_3309,N_3679);
nand U4801 (N_4801,N_2198,N_3943);
nand U4802 (N_4802,N_3820,N_2121);
and U4803 (N_4803,N_3513,N_2682);
nand U4804 (N_4804,N_2368,N_2415);
or U4805 (N_4805,N_3349,N_3525);
or U4806 (N_4806,N_2553,N_2495);
and U4807 (N_4807,N_3075,N_3717);
or U4808 (N_4808,N_3274,N_3387);
nand U4809 (N_4809,N_3314,N_2767);
and U4810 (N_4810,N_3434,N_3708);
nor U4811 (N_4811,N_2169,N_3762);
or U4812 (N_4812,N_2883,N_2072);
nor U4813 (N_4813,N_3734,N_2565);
or U4814 (N_4814,N_3667,N_2241);
nor U4815 (N_4815,N_3456,N_3978);
and U4816 (N_4816,N_3803,N_2887);
xnor U4817 (N_4817,N_3764,N_2394);
nor U4818 (N_4818,N_2817,N_3824);
or U4819 (N_4819,N_3637,N_3876);
xor U4820 (N_4820,N_3196,N_3082);
or U4821 (N_4821,N_3353,N_2834);
or U4822 (N_4822,N_3865,N_3209);
nand U4823 (N_4823,N_3663,N_3490);
nor U4824 (N_4824,N_3610,N_2380);
xor U4825 (N_4825,N_3689,N_3306);
nand U4826 (N_4826,N_2001,N_2401);
or U4827 (N_4827,N_3608,N_2861);
or U4828 (N_4828,N_2101,N_3744);
nor U4829 (N_4829,N_3103,N_3781);
and U4830 (N_4830,N_3197,N_2743);
nand U4831 (N_4831,N_2080,N_2523);
and U4832 (N_4832,N_2711,N_3207);
nand U4833 (N_4833,N_3026,N_3915);
nand U4834 (N_4834,N_2778,N_2610);
and U4835 (N_4835,N_2614,N_2194);
xnor U4836 (N_4836,N_3395,N_3430);
or U4837 (N_4837,N_3875,N_2798);
nand U4838 (N_4838,N_3520,N_3473);
and U4839 (N_4839,N_2066,N_2423);
or U4840 (N_4840,N_2408,N_3145);
and U4841 (N_4841,N_3927,N_2531);
nand U4842 (N_4842,N_2757,N_2329);
nor U4843 (N_4843,N_2037,N_2506);
or U4844 (N_4844,N_2449,N_2413);
or U4845 (N_4845,N_2824,N_3800);
or U4846 (N_4846,N_3945,N_2428);
or U4847 (N_4847,N_2649,N_2079);
xnor U4848 (N_4848,N_2156,N_2269);
or U4849 (N_4849,N_2962,N_3684);
nand U4850 (N_4850,N_2295,N_2096);
nor U4851 (N_4851,N_3115,N_3471);
nor U4852 (N_4852,N_2447,N_3324);
nor U4853 (N_4853,N_3277,N_2273);
nor U4854 (N_4854,N_2137,N_3808);
nor U4855 (N_4855,N_3045,N_3141);
or U4856 (N_4856,N_2370,N_2058);
xor U4857 (N_4857,N_2965,N_3428);
nor U4858 (N_4858,N_2257,N_2740);
and U4859 (N_4859,N_2894,N_2550);
and U4860 (N_4860,N_3661,N_2989);
or U4861 (N_4861,N_3466,N_2568);
or U4862 (N_4862,N_2377,N_3062);
or U4863 (N_4863,N_2756,N_3558);
nor U4864 (N_4864,N_2126,N_2032);
nand U4865 (N_4865,N_2454,N_2136);
nand U4866 (N_4866,N_2517,N_2525);
nand U4867 (N_4867,N_2952,N_2983);
and U4868 (N_4868,N_3301,N_3826);
xnor U4869 (N_4869,N_2087,N_3727);
and U4870 (N_4870,N_2406,N_3756);
or U4871 (N_4871,N_2841,N_2652);
and U4872 (N_4872,N_3659,N_2222);
nand U4873 (N_4873,N_2823,N_2800);
and U4874 (N_4874,N_3771,N_3577);
and U4875 (N_4875,N_2574,N_3385);
and U4876 (N_4876,N_3498,N_2282);
nand U4877 (N_4877,N_3266,N_2881);
nand U4878 (N_4878,N_2498,N_2243);
nor U4879 (N_4879,N_3015,N_2808);
nor U4880 (N_4880,N_3871,N_3079);
or U4881 (N_4881,N_3721,N_3287);
and U4882 (N_4882,N_3159,N_3332);
nor U4883 (N_4883,N_3453,N_2290);
xor U4884 (N_4884,N_3968,N_3231);
nand U4885 (N_4885,N_2563,N_2720);
nor U4886 (N_4886,N_3830,N_2272);
xor U4887 (N_4887,N_3896,N_2405);
nand U4888 (N_4888,N_3602,N_2092);
and U4889 (N_4889,N_2102,N_2355);
or U4890 (N_4890,N_3241,N_2113);
nand U4891 (N_4891,N_3776,N_2283);
nand U4892 (N_4892,N_3750,N_2893);
or U4893 (N_4893,N_3897,N_3298);
and U4894 (N_4894,N_2892,N_3444);
or U4895 (N_4895,N_2094,N_2972);
xor U4896 (N_4896,N_3982,N_2263);
or U4897 (N_4897,N_3355,N_3512);
nand U4898 (N_4898,N_3007,N_2077);
nand U4899 (N_4899,N_3859,N_3074);
xnor U4900 (N_4900,N_2483,N_3974);
nand U4901 (N_4901,N_2669,N_2191);
xor U4902 (N_4902,N_2482,N_3545);
nor U4903 (N_4903,N_3373,N_3538);
nand U4904 (N_4904,N_3747,N_2350);
or U4905 (N_4905,N_2681,N_2154);
or U4906 (N_4906,N_3644,N_2607);
nand U4907 (N_4907,N_3854,N_2641);
xor U4908 (N_4908,N_3791,N_2725);
and U4909 (N_4909,N_2270,N_2211);
nor U4910 (N_4910,N_2119,N_2502);
nand U4911 (N_4911,N_2378,N_3629);
xor U4912 (N_4912,N_3732,N_3907);
nand U4913 (N_4913,N_3592,N_2555);
or U4914 (N_4914,N_3020,N_3034);
nor U4915 (N_4915,N_3036,N_2806);
or U4916 (N_4916,N_2977,N_3726);
or U4917 (N_4917,N_2518,N_2692);
nor U4918 (N_4918,N_3175,N_3073);
nor U4919 (N_4919,N_2981,N_2810);
or U4920 (N_4920,N_3284,N_2572);
or U4921 (N_4921,N_2630,N_2427);
or U4922 (N_4922,N_2025,N_3291);
and U4923 (N_4923,N_2013,N_2536);
nor U4924 (N_4924,N_3935,N_2588);
nand U4925 (N_4925,N_2844,N_2391);
or U4926 (N_4926,N_2472,N_3364);
or U4927 (N_4927,N_2084,N_3189);
or U4928 (N_4928,N_2030,N_2288);
nor U4929 (N_4929,N_2479,N_2367);
nor U4930 (N_4930,N_2414,N_2062);
nor U4931 (N_4931,N_3948,N_3304);
xnor U4932 (N_4932,N_3676,N_2398);
and U4933 (N_4933,N_3930,N_2891);
or U4934 (N_4934,N_3544,N_2658);
or U4935 (N_4935,N_3470,N_2722);
and U4936 (N_4936,N_2259,N_3569);
xor U4937 (N_4937,N_3839,N_2328);
or U4938 (N_4938,N_3135,N_2796);
nor U4939 (N_4939,N_3888,N_3375);
or U4940 (N_4940,N_2201,N_3011);
nor U4941 (N_4941,N_2155,N_2689);
nor U4942 (N_4942,N_3032,N_3340);
xnor U4943 (N_4943,N_3863,N_2361);
and U4944 (N_4944,N_3374,N_3719);
and U4945 (N_4945,N_3579,N_3736);
and U4946 (N_4946,N_3113,N_2719);
and U4947 (N_4947,N_3612,N_2678);
and U4948 (N_4948,N_2233,N_2569);
and U4949 (N_4949,N_2045,N_2905);
or U4950 (N_4950,N_2160,N_3200);
nand U4951 (N_4951,N_3463,N_2467);
and U4952 (N_4952,N_3108,N_2353);
xor U4953 (N_4953,N_2594,N_2687);
nor U4954 (N_4954,N_2931,N_2407);
nand U4955 (N_4955,N_2897,N_3532);
nor U4956 (N_4956,N_3547,N_2042);
and U4957 (N_4957,N_2111,N_2696);
xor U4958 (N_4958,N_3660,N_3049);
and U4959 (N_4959,N_2857,N_3255);
or U4960 (N_4960,N_3990,N_3182);
and U4961 (N_4961,N_2043,N_3446);
nor U4962 (N_4962,N_2839,N_2748);
nor U4963 (N_4963,N_2543,N_3873);
xnor U4964 (N_4964,N_3379,N_2254);
xor U4965 (N_4965,N_3484,N_3779);
nand U4966 (N_4966,N_3223,N_2352);
nand U4967 (N_4967,N_3093,N_3858);
xor U4968 (N_4968,N_3505,N_2646);
nand U4969 (N_4969,N_3029,N_2684);
or U4970 (N_4970,N_3496,N_3832);
nand U4971 (N_4971,N_2916,N_2802);
or U4972 (N_4972,N_3731,N_3257);
nand U4973 (N_4973,N_2321,N_2476);
and U4974 (N_4974,N_3184,N_3194);
nand U4975 (N_4975,N_3057,N_3528);
and U4976 (N_4976,N_3480,N_3157);
and U4977 (N_4977,N_3337,N_3275);
nand U4978 (N_4978,N_2171,N_2168);
nor U4979 (N_4979,N_2103,N_2872);
and U4980 (N_4980,N_3122,N_3454);
or U4981 (N_4981,N_2303,N_2814);
xor U4982 (N_4982,N_2393,N_2229);
or U4983 (N_4983,N_2951,N_3581);
and U4984 (N_4984,N_3040,N_3128);
nor U4985 (N_4985,N_2713,N_2253);
or U4986 (N_4986,N_2845,N_3167);
or U4987 (N_4987,N_2921,N_2842);
xnor U4988 (N_4988,N_3386,N_2145);
or U4989 (N_4989,N_2954,N_3702);
nor U4990 (N_4990,N_3010,N_3575);
nand U4991 (N_4991,N_2601,N_3259);
and U4992 (N_4992,N_2116,N_3960);
and U4993 (N_4993,N_3325,N_2261);
nand U4994 (N_4994,N_3173,N_3422);
or U4995 (N_4995,N_3356,N_3695);
and U4996 (N_4996,N_2524,N_3425);
nor U4997 (N_4997,N_2799,N_3916);
nor U4998 (N_4998,N_3303,N_3831);
and U4999 (N_4999,N_2085,N_2185);
nor U5000 (N_5000,N_3778,N_2485);
nor U5001 (N_5001,N_2528,N_2857);
and U5002 (N_5002,N_2356,N_2843);
or U5003 (N_5003,N_2115,N_2208);
nand U5004 (N_5004,N_3391,N_3153);
and U5005 (N_5005,N_3945,N_3057);
and U5006 (N_5006,N_2859,N_2005);
and U5007 (N_5007,N_3571,N_3289);
nand U5008 (N_5008,N_2738,N_3128);
nand U5009 (N_5009,N_3816,N_3059);
or U5010 (N_5010,N_3824,N_3810);
and U5011 (N_5011,N_3668,N_2584);
nand U5012 (N_5012,N_2598,N_2015);
nor U5013 (N_5013,N_3671,N_2812);
and U5014 (N_5014,N_3370,N_2625);
xor U5015 (N_5015,N_2555,N_2702);
nor U5016 (N_5016,N_3772,N_2918);
nand U5017 (N_5017,N_2281,N_3985);
nor U5018 (N_5018,N_2705,N_2409);
and U5019 (N_5019,N_3446,N_2266);
nand U5020 (N_5020,N_3785,N_2125);
xnor U5021 (N_5021,N_2775,N_3545);
and U5022 (N_5022,N_2444,N_3204);
nand U5023 (N_5023,N_3092,N_3186);
or U5024 (N_5024,N_2800,N_3889);
nand U5025 (N_5025,N_2670,N_2884);
nor U5026 (N_5026,N_2496,N_3560);
and U5027 (N_5027,N_3623,N_2150);
or U5028 (N_5028,N_2531,N_2314);
xor U5029 (N_5029,N_2032,N_2246);
nor U5030 (N_5030,N_3104,N_2735);
and U5031 (N_5031,N_2271,N_3320);
or U5032 (N_5032,N_3594,N_3614);
or U5033 (N_5033,N_3377,N_2899);
nand U5034 (N_5034,N_3397,N_3984);
nand U5035 (N_5035,N_3980,N_3577);
and U5036 (N_5036,N_3926,N_3647);
or U5037 (N_5037,N_2196,N_2236);
or U5038 (N_5038,N_3445,N_3194);
nand U5039 (N_5039,N_3101,N_2033);
and U5040 (N_5040,N_3432,N_2390);
or U5041 (N_5041,N_3398,N_3276);
xnor U5042 (N_5042,N_3083,N_3017);
xnor U5043 (N_5043,N_3612,N_2026);
xnor U5044 (N_5044,N_2937,N_2272);
nor U5045 (N_5045,N_3344,N_2642);
nand U5046 (N_5046,N_3203,N_2947);
nor U5047 (N_5047,N_3071,N_2590);
and U5048 (N_5048,N_2814,N_3582);
and U5049 (N_5049,N_3280,N_3006);
or U5050 (N_5050,N_3074,N_2303);
nand U5051 (N_5051,N_2343,N_2942);
and U5052 (N_5052,N_2071,N_2994);
nor U5053 (N_5053,N_3048,N_3956);
nand U5054 (N_5054,N_3927,N_3903);
and U5055 (N_5055,N_2610,N_3471);
and U5056 (N_5056,N_2538,N_2243);
or U5057 (N_5057,N_2284,N_3513);
and U5058 (N_5058,N_3721,N_2494);
nor U5059 (N_5059,N_2846,N_3818);
nor U5060 (N_5060,N_2697,N_2889);
nor U5061 (N_5061,N_2087,N_3325);
nand U5062 (N_5062,N_2846,N_2339);
nand U5063 (N_5063,N_3757,N_3236);
nor U5064 (N_5064,N_3652,N_3473);
and U5065 (N_5065,N_3838,N_3933);
and U5066 (N_5066,N_3778,N_3103);
or U5067 (N_5067,N_2797,N_3857);
xor U5068 (N_5068,N_2312,N_2390);
and U5069 (N_5069,N_2315,N_3690);
and U5070 (N_5070,N_3867,N_2564);
xnor U5071 (N_5071,N_3118,N_3554);
or U5072 (N_5072,N_2873,N_3988);
nor U5073 (N_5073,N_2590,N_2324);
nor U5074 (N_5074,N_3851,N_2063);
or U5075 (N_5075,N_2278,N_3093);
and U5076 (N_5076,N_2556,N_2491);
or U5077 (N_5077,N_3284,N_3061);
xor U5078 (N_5078,N_3869,N_2034);
or U5079 (N_5079,N_3851,N_3520);
nand U5080 (N_5080,N_3463,N_2745);
or U5081 (N_5081,N_3206,N_3763);
and U5082 (N_5082,N_2001,N_2621);
and U5083 (N_5083,N_2666,N_2674);
nor U5084 (N_5084,N_3702,N_2671);
or U5085 (N_5085,N_3815,N_3530);
nand U5086 (N_5086,N_2687,N_3400);
nor U5087 (N_5087,N_2810,N_3737);
nor U5088 (N_5088,N_2363,N_3732);
and U5089 (N_5089,N_2002,N_2616);
nand U5090 (N_5090,N_3775,N_2273);
and U5091 (N_5091,N_3349,N_2412);
nand U5092 (N_5092,N_3360,N_3865);
nand U5093 (N_5093,N_2354,N_2991);
or U5094 (N_5094,N_2193,N_3642);
or U5095 (N_5095,N_3036,N_2701);
nand U5096 (N_5096,N_2079,N_3203);
and U5097 (N_5097,N_2092,N_2058);
nand U5098 (N_5098,N_2359,N_2283);
nor U5099 (N_5099,N_2991,N_3249);
xnor U5100 (N_5100,N_3843,N_3668);
or U5101 (N_5101,N_2983,N_3295);
nand U5102 (N_5102,N_3766,N_2467);
nor U5103 (N_5103,N_2796,N_2679);
and U5104 (N_5104,N_2487,N_2118);
or U5105 (N_5105,N_2349,N_2880);
xnor U5106 (N_5106,N_2564,N_2432);
or U5107 (N_5107,N_2139,N_2977);
or U5108 (N_5108,N_3388,N_3865);
and U5109 (N_5109,N_3909,N_3987);
xor U5110 (N_5110,N_3668,N_2273);
xor U5111 (N_5111,N_2032,N_2254);
or U5112 (N_5112,N_2106,N_3899);
nor U5113 (N_5113,N_3185,N_2148);
nor U5114 (N_5114,N_2640,N_3257);
nand U5115 (N_5115,N_2935,N_3534);
or U5116 (N_5116,N_3761,N_3376);
nor U5117 (N_5117,N_2583,N_3826);
nor U5118 (N_5118,N_3245,N_3745);
and U5119 (N_5119,N_3380,N_2977);
nand U5120 (N_5120,N_2213,N_2444);
nand U5121 (N_5121,N_2486,N_2980);
and U5122 (N_5122,N_2743,N_2646);
and U5123 (N_5123,N_2226,N_2807);
nand U5124 (N_5124,N_2973,N_3520);
nor U5125 (N_5125,N_3103,N_2726);
nand U5126 (N_5126,N_3678,N_3289);
nand U5127 (N_5127,N_2856,N_3952);
xor U5128 (N_5128,N_2444,N_2528);
nor U5129 (N_5129,N_3195,N_3587);
or U5130 (N_5130,N_3450,N_3511);
or U5131 (N_5131,N_3906,N_2352);
nand U5132 (N_5132,N_3632,N_2980);
and U5133 (N_5133,N_3111,N_2843);
and U5134 (N_5134,N_2215,N_3822);
or U5135 (N_5135,N_3741,N_2462);
nand U5136 (N_5136,N_2756,N_3330);
nand U5137 (N_5137,N_2763,N_2939);
or U5138 (N_5138,N_2303,N_3744);
or U5139 (N_5139,N_2234,N_3058);
and U5140 (N_5140,N_2312,N_3973);
nand U5141 (N_5141,N_2589,N_2029);
nor U5142 (N_5142,N_3674,N_2684);
xor U5143 (N_5143,N_2193,N_2212);
nor U5144 (N_5144,N_3485,N_2616);
and U5145 (N_5145,N_2926,N_3950);
nor U5146 (N_5146,N_3948,N_3984);
nor U5147 (N_5147,N_2069,N_3313);
and U5148 (N_5148,N_2577,N_2115);
or U5149 (N_5149,N_3276,N_2140);
nor U5150 (N_5150,N_3792,N_2707);
and U5151 (N_5151,N_3957,N_3487);
nor U5152 (N_5152,N_2780,N_3858);
xor U5153 (N_5153,N_2432,N_3507);
nor U5154 (N_5154,N_3667,N_2786);
nand U5155 (N_5155,N_3912,N_3085);
or U5156 (N_5156,N_3636,N_3716);
and U5157 (N_5157,N_3909,N_3442);
and U5158 (N_5158,N_3864,N_3131);
xor U5159 (N_5159,N_2077,N_2481);
or U5160 (N_5160,N_2387,N_2034);
or U5161 (N_5161,N_2414,N_3812);
nor U5162 (N_5162,N_2216,N_3443);
and U5163 (N_5163,N_3170,N_3742);
and U5164 (N_5164,N_2633,N_3451);
or U5165 (N_5165,N_3515,N_3136);
xor U5166 (N_5166,N_3886,N_3101);
nor U5167 (N_5167,N_3195,N_3161);
nor U5168 (N_5168,N_3846,N_3672);
or U5169 (N_5169,N_3762,N_2451);
or U5170 (N_5170,N_3737,N_2199);
nor U5171 (N_5171,N_2793,N_3340);
nor U5172 (N_5172,N_3662,N_3990);
nand U5173 (N_5173,N_2418,N_2071);
nor U5174 (N_5174,N_2166,N_3206);
nor U5175 (N_5175,N_3606,N_2225);
nor U5176 (N_5176,N_3640,N_3743);
nor U5177 (N_5177,N_3617,N_3749);
and U5178 (N_5178,N_2502,N_3907);
xor U5179 (N_5179,N_2906,N_3105);
and U5180 (N_5180,N_3442,N_3518);
nand U5181 (N_5181,N_3849,N_3497);
or U5182 (N_5182,N_2816,N_2786);
xnor U5183 (N_5183,N_3554,N_3388);
nor U5184 (N_5184,N_2177,N_3572);
and U5185 (N_5185,N_3481,N_3097);
nand U5186 (N_5186,N_3902,N_3278);
or U5187 (N_5187,N_3100,N_2398);
nand U5188 (N_5188,N_3678,N_3669);
or U5189 (N_5189,N_2665,N_3636);
or U5190 (N_5190,N_3152,N_2829);
and U5191 (N_5191,N_2416,N_3287);
nand U5192 (N_5192,N_3989,N_2899);
and U5193 (N_5193,N_2902,N_2929);
nand U5194 (N_5194,N_2118,N_3225);
nor U5195 (N_5195,N_3321,N_3257);
or U5196 (N_5196,N_2460,N_3682);
and U5197 (N_5197,N_2316,N_3109);
and U5198 (N_5198,N_2130,N_2967);
or U5199 (N_5199,N_3387,N_3658);
nand U5200 (N_5200,N_2524,N_2364);
xnor U5201 (N_5201,N_2223,N_2977);
or U5202 (N_5202,N_2948,N_3708);
nand U5203 (N_5203,N_3350,N_2648);
and U5204 (N_5204,N_3833,N_3777);
or U5205 (N_5205,N_3189,N_2846);
nand U5206 (N_5206,N_2795,N_3067);
nand U5207 (N_5207,N_2333,N_3157);
and U5208 (N_5208,N_3065,N_3772);
nand U5209 (N_5209,N_3681,N_2876);
and U5210 (N_5210,N_2850,N_2062);
and U5211 (N_5211,N_3247,N_3931);
nor U5212 (N_5212,N_2633,N_2500);
nand U5213 (N_5213,N_3680,N_2329);
or U5214 (N_5214,N_3344,N_2453);
nor U5215 (N_5215,N_2930,N_3056);
nor U5216 (N_5216,N_2388,N_3379);
nor U5217 (N_5217,N_2489,N_3839);
nor U5218 (N_5218,N_2377,N_3510);
and U5219 (N_5219,N_2297,N_2553);
and U5220 (N_5220,N_3574,N_3225);
or U5221 (N_5221,N_2248,N_2078);
nand U5222 (N_5222,N_3040,N_2364);
nand U5223 (N_5223,N_2151,N_3093);
and U5224 (N_5224,N_2137,N_3422);
nor U5225 (N_5225,N_3705,N_3432);
nor U5226 (N_5226,N_2878,N_3789);
nand U5227 (N_5227,N_2384,N_2815);
and U5228 (N_5228,N_2933,N_2826);
nor U5229 (N_5229,N_2761,N_2019);
nor U5230 (N_5230,N_3392,N_2307);
xnor U5231 (N_5231,N_2199,N_3320);
nand U5232 (N_5232,N_2939,N_3953);
nand U5233 (N_5233,N_3380,N_3632);
or U5234 (N_5234,N_2197,N_3366);
and U5235 (N_5235,N_3365,N_3994);
nand U5236 (N_5236,N_2327,N_2818);
and U5237 (N_5237,N_3413,N_2365);
or U5238 (N_5238,N_2830,N_2851);
or U5239 (N_5239,N_2925,N_2596);
nor U5240 (N_5240,N_2098,N_2084);
nand U5241 (N_5241,N_2755,N_3856);
nand U5242 (N_5242,N_3816,N_2715);
nand U5243 (N_5243,N_2167,N_3621);
or U5244 (N_5244,N_2156,N_3191);
and U5245 (N_5245,N_3821,N_2446);
or U5246 (N_5246,N_2707,N_3444);
nor U5247 (N_5247,N_3971,N_2935);
xor U5248 (N_5248,N_3765,N_3688);
and U5249 (N_5249,N_3355,N_3853);
or U5250 (N_5250,N_2581,N_2323);
and U5251 (N_5251,N_3267,N_3122);
nand U5252 (N_5252,N_3432,N_3481);
xor U5253 (N_5253,N_2588,N_3450);
nand U5254 (N_5254,N_2341,N_2656);
nand U5255 (N_5255,N_3286,N_3825);
nand U5256 (N_5256,N_2527,N_3643);
or U5257 (N_5257,N_3335,N_3441);
nor U5258 (N_5258,N_2226,N_2314);
nor U5259 (N_5259,N_3872,N_2040);
nor U5260 (N_5260,N_2671,N_3223);
xnor U5261 (N_5261,N_2926,N_2457);
nand U5262 (N_5262,N_3972,N_2637);
or U5263 (N_5263,N_2697,N_2220);
and U5264 (N_5264,N_3437,N_2608);
or U5265 (N_5265,N_3390,N_3663);
nand U5266 (N_5266,N_3996,N_3428);
and U5267 (N_5267,N_3983,N_3220);
nor U5268 (N_5268,N_2344,N_3274);
and U5269 (N_5269,N_2443,N_3494);
and U5270 (N_5270,N_3819,N_2144);
nor U5271 (N_5271,N_3870,N_2332);
nand U5272 (N_5272,N_2258,N_2659);
and U5273 (N_5273,N_2593,N_3715);
nor U5274 (N_5274,N_2432,N_2666);
nand U5275 (N_5275,N_2898,N_3734);
and U5276 (N_5276,N_3757,N_3117);
or U5277 (N_5277,N_2308,N_2751);
and U5278 (N_5278,N_3842,N_3771);
xnor U5279 (N_5279,N_2266,N_3004);
nand U5280 (N_5280,N_3590,N_3101);
and U5281 (N_5281,N_2416,N_2805);
nand U5282 (N_5282,N_2358,N_3580);
or U5283 (N_5283,N_3901,N_3789);
or U5284 (N_5284,N_2933,N_2848);
nor U5285 (N_5285,N_2451,N_3420);
and U5286 (N_5286,N_2605,N_3700);
or U5287 (N_5287,N_3042,N_2534);
nand U5288 (N_5288,N_2318,N_3319);
or U5289 (N_5289,N_2763,N_3862);
nor U5290 (N_5290,N_3362,N_2445);
nor U5291 (N_5291,N_3769,N_3784);
or U5292 (N_5292,N_2791,N_3592);
or U5293 (N_5293,N_3865,N_2666);
or U5294 (N_5294,N_3816,N_3340);
xor U5295 (N_5295,N_3079,N_3779);
or U5296 (N_5296,N_3885,N_2835);
xor U5297 (N_5297,N_2066,N_2808);
nand U5298 (N_5298,N_3854,N_3684);
or U5299 (N_5299,N_3587,N_3353);
xor U5300 (N_5300,N_3225,N_2921);
nand U5301 (N_5301,N_3574,N_2860);
nor U5302 (N_5302,N_2641,N_2004);
xnor U5303 (N_5303,N_2470,N_2688);
and U5304 (N_5304,N_3828,N_3117);
and U5305 (N_5305,N_3038,N_2404);
and U5306 (N_5306,N_2529,N_3622);
xor U5307 (N_5307,N_3886,N_2523);
or U5308 (N_5308,N_2929,N_2038);
and U5309 (N_5309,N_3872,N_3321);
or U5310 (N_5310,N_2617,N_3380);
xor U5311 (N_5311,N_3947,N_2605);
or U5312 (N_5312,N_3664,N_2305);
nand U5313 (N_5313,N_3786,N_3629);
nor U5314 (N_5314,N_3000,N_3024);
nor U5315 (N_5315,N_3096,N_2537);
nor U5316 (N_5316,N_2254,N_3450);
nor U5317 (N_5317,N_3650,N_2034);
nand U5318 (N_5318,N_2620,N_3733);
nor U5319 (N_5319,N_3577,N_3635);
nor U5320 (N_5320,N_3662,N_3297);
and U5321 (N_5321,N_2052,N_2929);
and U5322 (N_5322,N_2467,N_3608);
xor U5323 (N_5323,N_2060,N_2133);
nor U5324 (N_5324,N_2020,N_3896);
nor U5325 (N_5325,N_3831,N_3432);
and U5326 (N_5326,N_2758,N_3982);
and U5327 (N_5327,N_3338,N_3603);
or U5328 (N_5328,N_3318,N_3716);
or U5329 (N_5329,N_3022,N_2666);
and U5330 (N_5330,N_3975,N_3527);
nor U5331 (N_5331,N_3620,N_3581);
nand U5332 (N_5332,N_3756,N_3656);
and U5333 (N_5333,N_2503,N_3442);
nor U5334 (N_5334,N_3523,N_3117);
nor U5335 (N_5335,N_3011,N_2787);
nor U5336 (N_5336,N_2255,N_3414);
and U5337 (N_5337,N_2502,N_2752);
nand U5338 (N_5338,N_3453,N_3081);
and U5339 (N_5339,N_3003,N_3481);
xor U5340 (N_5340,N_2744,N_2837);
or U5341 (N_5341,N_2126,N_2901);
nand U5342 (N_5342,N_3509,N_3631);
nor U5343 (N_5343,N_3808,N_3474);
or U5344 (N_5344,N_2391,N_2501);
nor U5345 (N_5345,N_2290,N_2971);
and U5346 (N_5346,N_2556,N_3191);
or U5347 (N_5347,N_2884,N_3230);
xnor U5348 (N_5348,N_3515,N_3994);
nor U5349 (N_5349,N_3044,N_3878);
nand U5350 (N_5350,N_3620,N_2016);
nand U5351 (N_5351,N_3039,N_2482);
nand U5352 (N_5352,N_3009,N_3906);
nor U5353 (N_5353,N_3348,N_3709);
xor U5354 (N_5354,N_2993,N_2013);
nor U5355 (N_5355,N_3193,N_2306);
or U5356 (N_5356,N_3098,N_2764);
nor U5357 (N_5357,N_2533,N_2140);
nand U5358 (N_5358,N_2117,N_3878);
and U5359 (N_5359,N_3215,N_3324);
and U5360 (N_5360,N_3225,N_2401);
nand U5361 (N_5361,N_3570,N_2954);
and U5362 (N_5362,N_3647,N_2554);
nand U5363 (N_5363,N_3133,N_2561);
nor U5364 (N_5364,N_2110,N_2463);
nor U5365 (N_5365,N_3260,N_2775);
nor U5366 (N_5366,N_3813,N_2546);
and U5367 (N_5367,N_2116,N_2265);
nand U5368 (N_5368,N_3000,N_2539);
nand U5369 (N_5369,N_2532,N_2674);
nand U5370 (N_5370,N_3762,N_3028);
nor U5371 (N_5371,N_2109,N_3851);
nand U5372 (N_5372,N_2984,N_2028);
and U5373 (N_5373,N_2458,N_3527);
and U5374 (N_5374,N_3513,N_3908);
nor U5375 (N_5375,N_3980,N_3927);
and U5376 (N_5376,N_3575,N_3871);
or U5377 (N_5377,N_3688,N_2505);
and U5378 (N_5378,N_2750,N_2736);
nor U5379 (N_5379,N_2168,N_2790);
nor U5380 (N_5380,N_3599,N_2844);
nand U5381 (N_5381,N_3442,N_3381);
xnor U5382 (N_5382,N_3018,N_2813);
xor U5383 (N_5383,N_2538,N_2170);
nand U5384 (N_5384,N_3627,N_2089);
or U5385 (N_5385,N_2746,N_2757);
and U5386 (N_5386,N_3707,N_2532);
nand U5387 (N_5387,N_3521,N_3374);
nor U5388 (N_5388,N_2386,N_3214);
nand U5389 (N_5389,N_3259,N_3730);
and U5390 (N_5390,N_3712,N_3965);
or U5391 (N_5391,N_2501,N_2742);
nor U5392 (N_5392,N_2062,N_3240);
or U5393 (N_5393,N_2276,N_3679);
nand U5394 (N_5394,N_2869,N_3431);
nor U5395 (N_5395,N_3874,N_2154);
and U5396 (N_5396,N_2043,N_2656);
and U5397 (N_5397,N_2506,N_2468);
nor U5398 (N_5398,N_2297,N_3999);
and U5399 (N_5399,N_2003,N_2942);
nand U5400 (N_5400,N_3478,N_3244);
nand U5401 (N_5401,N_2817,N_3238);
or U5402 (N_5402,N_2393,N_3431);
nor U5403 (N_5403,N_2929,N_3400);
and U5404 (N_5404,N_3968,N_3014);
and U5405 (N_5405,N_2039,N_2370);
xor U5406 (N_5406,N_2866,N_2984);
nand U5407 (N_5407,N_2322,N_3226);
nand U5408 (N_5408,N_2723,N_2895);
nand U5409 (N_5409,N_3119,N_2406);
nor U5410 (N_5410,N_2569,N_2287);
nand U5411 (N_5411,N_3716,N_2390);
nand U5412 (N_5412,N_3587,N_2052);
or U5413 (N_5413,N_2345,N_3570);
and U5414 (N_5414,N_2674,N_2255);
or U5415 (N_5415,N_3310,N_3511);
or U5416 (N_5416,N_2711,N_2551);
nor U5417 (N_5417,N_2148,N_2983);
or U5418 (N_5418,N_2285,N_3975);
or U5419 (N_5419,N_3910,N_2973);
nor U5420 (N_5420,N_3769,N_2731);
nor U5421 (N_5421,N_2031,N_3162);
or U5422 (N_5422,N_3824,N_3658);
nand U5423 (N_5423,N_2134,N_2909);
nand U5424 (N_5424,N_3953,N_2290);
nor U5425 (N_5425,N_2842,N_3928);
nor U5426 (N_5426,N_3659,N_3880);
or U5427 (N_5427,N_3054,N_2861);
and U5428 (N_5428,N_3672,N_2659);
and U5429 (N_5429,N_2080,N_3583);
or U5430 (N_5430,N_2291,N_3011);
nor U5431 (N_5431,N_2749,N_2046);
nor U5432 (N_5432,N_3768,N_2991);
or U5433 (N_5433,N_3407,N_2882);
and U5434 (N_5434,N_2912,N_2817);
nand U5435 (N_5435,N_2990,N_3857);
nand U5436 (N_5436,N_3966,N_3381);
xnor U5437 (N_5437,N_2674,N_3301);
nand U5438 (N_5438,N_2761,N_2396);
xnor U5439 (N_5439,N_3053,N_2399);
or U5440 (N_5440,N_2613,N_3695);
and U5441 (N_5441,N_2421,N_2316);
or U5442 (N_5442,N_3565,N_3611);
nor U5443 (N_5443,N_3495,N_2817);
and U5444 (N_5444,N_3774,N_2657);
and U5445 (N_5445,N_2919,N_2925);
xor U5446 (N_5446,N_2654,N_2429);
nand U5447 (N_5447,N_3065,N_2931);
and U5448 (N_5448,N_2636,N_3701);
nand U5449 (N_5449,N_3411,N_2327);
xnor U5450 (N_5450,N_2573,N_3201);
and U5451 (N_5451,N_2934,N_2245);
nand U5452 (N_5452,N_2107,N_3514);
nor U5453 (N_5453,N_2706,N_2791);
and U5454 (N_5454,N_3836,N_2418);
nand U5455 (N_5455,N_2787,N_3694);
nor U5456 (N_5456,N_3975,N_3841);
nand U5457 (N_5457,N_2815,N_2762);
and U5458 (N_5458,N_2004,N_3637);
and U5459 (N_5459,N_3951,N_2635);
or U5460 (N_5460,N_3864,N_2822);
or U5461 (N_5461,N_2505,N_3156);
nand U5462 (N_5462,N_3848,N_2234);
and U5463 (N_5463,N_3958,N_2592);
or U5464 (N_5464,N_2526,N_2180);
nand U5465 (N_5465,N_2572,N_3328);
nand U5466 (N_5466,N_3362,N_3062);
nand U5467 (N_5467,N_2075,N_3880);
or U5468 (N_5468,N_3433,N_3574);
and U5469 (N_5469,N_3330,N_3707);
or U5470 (N_5470,N_3290,N_2460);
nor U5471 (N_5471,N_2886,N_3742);
and U5472 (N_5472,N_2442,N_3657);
and U5473 (N_5473,N_2158,N_3935);
nor U5474 (N_5474,N_2503,N_3799);
nor U5475 (N_5475,N_3097,N_2232);
nor U5476 (N_5476,N_3021,N_3446);
xor U5477 (N_5477,N_2722,N_3669);
nand U5478 (N_5478,N_3735,N_3906);
xnor U5479 (N_5479,N_3886,N_2155);
nor U5480 (N_5480,N_3466,N_3814);
nand U5481 (N_5481,N_2419,N_2556);
nand U5482 (N_5482,N_3546,N_2821);
nand U5483 (N_5483,N_3893,N_3121);
xnor U5484 (N_5484,N_2752,N_3813);
xor U5485 (N_5485,N_3932,N_3077);
nand U5486 (N_5486,N_2458,N_2806);
nand U5487 (N_5487,N_2667,N_2184);
nand U5488 (N_5488,N_2500,N_2595);
and U5489 (N_5489,N_3625,N_3855);
and U5490 (N_5490,N_2868,N_3843);
nand U5491 (N_5491,N_2628,N_2508);
xnor U5492 (N_5492,N_2433,N_3988);
or U5493 (N_5493,N_2826,N_3503);
nand U5494 (N_5494,N_2975,N_3154);
nor U5495 (N_5495,N_2485,N_3570);
or U5496 (N_5496,N_3865,N_2263);
nand U5497 (N_5497,N_2572,N_3886);
xor U5498 (N_5498,N_2462,N_2502);
nand U5499 (N_5499,N_3097,N_2408);
nand U5500 (N_5500,N_2103,N_2265);
nand U5501 (N_5501,N_3770,N_2695);
and U5502 (N_5502,N_2338,N_3497);
and U5503 (N_5503,N_2662,N_2964);
xor U5504 (N_5504,N_3402,N_3119);
and U5505 (N_5505,N_2819,N_3214);
nor U5506 (N_5506,N_3056,N_3769);
and U5507 (N_5507,N_3114,N_2904);
nor U5508 (N_5508,N_2657,N_3845);
nor U5509 (N_5509,N_2113,N_2166);
or U5510 (N_5510,N_3447,N_3092);
or U5511 (N_5511,N_2742,N_3381);
nor U5512 (N_5512,N_3301,N_2629);
or U5513 (N_5513,N_3859,N_2391);
xor U5514 (N_5514,N_3810,N_2630);
nand U5515 (N_5515,N_3927,N_2761);
or U5516 (N_5516,N_3528,N_2728);
nand U5517 (N_5517,N_3770,N_2783);
or U5518 (N_5518,N_3232,N_2454);
or U5519 (N_5519,N_3503,N_3773);
nand U5520 (N_5520,N_2543,N_2782);
and U5521 (N_5521,N_2990,N_3320);
nor U5522 (N_5522,N_2093,N_3830);
or U5523 (N_5523,N_2460,N_3488);
xnor U5524 (N_5524,N_3865,N_3206);
nor U5525 (N_5525,N_2646,N_3146);
nand U5526 (N_5526,N_2170,N_3421);
nand U5527 (N_5527,N_3943,N_2790);
nand U5528 (N_5528,N_3805,N_2676);
and U5529 (N_5529,N_2238,N_3541);
nand U5530 (N_5530,N_2169,N_3815);
or U5531 (N_5531,N_3898,N_3137);
xor U5532 (N_5532,N_2729,N_2111);
and U5533 (N_5533,N_3945,N_3887);
nor U5534 (N_5534,N_3084,N_2871);
and U5535 (N_5535,N_2824,N_3581);
and U5536 (N_5536,N_3063,N_3132);
nor U5537 (N_5537,N_3010,N_2958);
nor U5538 (N_5538,N_3913,N_2734);
or U5539 (N_5539,N_2625,N_3948);
nand U5540 (N_5540,N_2125,N_3598);
nand U5541 (N_5541,N_2026,N_3681);
nor U5542 (N_5542,N_3171,N_2217);
nor U5543 (N_5543,N_2178,N_3204);
or U5544 (N_5544,N_3953,N_3512);
xor U5545 (N_5545,N_2062,N_3559);
nand U5546 (N_5546,N_2248,N_2442);
and U5547 (N_5547,N_3866,N_3613);
nand U5548 (N_5548,N_2824,N_2741);
nor U5549 (N_5549,N_2151,N_2543);
or U5550 (N_5550,N_2186,N_3785);
nand U5551 (N_5551,N_2356,N_2661);
or U5552 (N_5552,N_3246,N_2491);
nor U5553 (N_5553,N_2991,N_2793);
or U5554 (N_5554,N_2714,N_2848);
xnor U5555 (N_5555,N_2615,N_3170);
and U5556 (N_5556,N_3618,N_2124);
nand U5557 (N_5557,N_2763,N_3690);
nand U5558 (N_5558,N_3508,N_3579);
and U5559 (N_5559,N_2639,N_2916);
nor U5560 (N_5560,N_2665,N_2807);
or U5561 (N_5561,N_2966,N_3619);
nand U5562 (N_5562,N_2024,N_3477);
nor U5563 (N_5563,N_3030,N_3156);
and U5564 (N_5564,N_2574,N_2751);
nand U5565 (N_5565,N_3592,N_2874);
or U5566 (N_5566,N_3121,N_2897);
and U5567 (N_5567,N_3030,N_3663);
nand U5568 (N_5568,N_2711,N_2952);
nor U5569 (N_5569,N_2674,N_2555);
nor U5570 (N_5570,N_2441,N_2922);
and U5571 (N_5571,N_2385,N_2554);
and U5572 (N_5572,N_3198,N_3811);
nand U5573 (N_5573,N_3376,N_3901);
nand U5574 (N_5574,N_3795,N_3349);
and U5575 (N_5575,N_3399,N_3670);
nor U5576 (N_5576,N_2310,N_2438);
or U5577 (N_5577,N_3099,N_3115);
nand U5578 (N_5578,N_2400,N_3359);
or U5579 (N_5579,N_2559,N_2394);
or U5580 (N_5580,N_3865,N_2657);
xnor U5581 (N_5581,N_3152,N_2585);
nor U5582 (N_5582,N_3901,N_2960);
nor U5583 (N_5583,N_3471,N_3014);
and U5584 (N_5584,N_3148,N_3397);
nand U5585 (N_5585,N_2453,N_3528);
xnor U5586 (N_5586,N_3429,N_3289);
nand U5587 (N_5587,N_3644,N_2708);
and U5588 (N_5588,N_3138,N_3516);
nand U5589 (N_5589,N_2981,N_3828);
nor U5590 (N_5590,N_3628,N_3251);
or U5591 (N_5591,N_3731,N_3857);
and U5592 (N_5592,N_2498,N_2902);
or U5593 (N_5593,N_3863,N_3385);
nand U5594 (N_5594,N_3146,N_2492);
or U5595 (N_5595,N_3579,N_3659);
or U5596 (N_5596,N_3824,N_2836);
or U5597 (N_5597,N_2713,N_2462);
nor U5598 (N_5598,N_3158,N_2293);
or U5599 (N_5599,N_3976,N_3550);
nor U5600 (N_5600,N_3087,N_2444);
nand U5601 (N_5601,N_2553,N_3414);
and U5602 (N_5602,N_2782,N_3376);
or U5603 (N_5603,N_2981,N_2767);
xor U5604 (N_5604,N_3928,N_2720);
and U5605 (N_5605,N_2105,N_2821);
nand U5606 (N_5606,N_3051,N_2413);
and U5607 (N_5607,N_3200,N_2880);
nand U5608 (N_5608,N_2636,N_2858);
nor U5609 (N_5609,N_2965,N_3156);
nor U5610 (N_5610,N_2114,N_2645);
or U5611 (N_5611,N_2094,N_3964);
nor U5612 (N_5612,N_3912,N_3023);
and U5613 (N_5613,N_3375,N_2482);
or U5614 (N_5614,N_3552,N_2915);
and U5615 (N_5615,N_2356,N_3572);
and U5616 (N_5616,N_2870,N_3121);
and U5617 (N_5617,N_3193,N_2291);
nor U5618 (N_5618,N_3295,N_2549);
xnor U5619 (N_5619,N_3243,N_2542);
xnor U5620 (N_5620,N_2345,N_2143);
or U5621 (N_5621,N_2345,N_3683);
or U5622 (N_5622,N_3533,N_3018);
and U5623 (N_5623,N_3465,N_2106);
nor U5624 (N_5624,N_3353,N_3854);
nor U5625 (N_5625,N_3358,N_3263);
xor U5626 (N_5626,N_2876,N_2817);
and U5627 (N_5627,N_3649,N_3715);
nand U5628 (N_5628,N_3356,N_3751);
nor U5629 (N_5629,N_3087,N_3288);
nand U5630 (N_5630,N_3941,N_3304);
and U5631 (N_5631,N_2251,N_3264);
and U5632 (N_5632,N_2615,N_2768);
and U5633 (N_5633,N_3480,N_2185);
or U5634 (N_5634,N_2166,N_2450);
nand U5635 (N_5635,N_3553,N_2102);
and U5636 (N_5636,N_2624,N_2001);
and U5637 (N_5637,N_2524,N_3617);
nand U5638 (N_5638,N_2424,N_3323);
and U5639 (N_5639,N_3359,N_2975);
nor U5640 (N_5640,N_2608,N_2797);
nor U5641 (N_5641,N_2701,N_3988);
or U5642 (N_5642,N_2967,N_2828);
and U5643 (N_5643,N_2687,N_2384);
and U5644 (N_5644,N_3483,N_2332);
nor U5645 (N_5645,N_2584,N_3518);
nor U5646 (N_5646,N_2260,N_3613);
nand U5647 (N_5647,N_2489,N_3115);
and U5648 (N_5648,N_3325,N_3995);
xor U5649 (N_5649,N_2773,N_3202);
nor U5650 (N_5650,N_2420,N_3152);
nand U5651 (N_5651,N_2704,N_2508);
nor U5652 (N_5652,N_3464,N_2422);
or U5653 (N_5653,N_3366,N_2053);
nor U5654 (N_5654,N_2182,N_2526);
nor U5655 (N_5655,N_2772,N_3946);
xnor U5656 (N_5656,N_2539,N_3461);
or U5657 (N_5657,N_3127,N_2993);
and U5658 (N_5658,N_2151,N_3025);
xnor U5659 (N_5659,N_3046,N_2091);
nand U5660 (N_5660,N_2893,N_3161);
nand U5661 (N_5661,N_3275,N_3960);
and U5662 (N_5662,N_2175,N_2653);
and U5663 (N_5663,N_2741,N_3764);
xor U5664 (N_5664,N_2131,N_3378);
xnor U5665 (N_5665,N_3810,N_2063);
and U5666 (N_5666,N_2523,N_2214);
xor U5667 (N_5667,N_2296,N_2250);
nand U5668 (N_5668,N_2495,N_3254);
or U5669 (N_5669,N_3222,N_2272);
or U5670 (N_5670,N_3371,N_2393);
nand U5671 (N_5671,N_3712,N_3500);
or U5672 (N_5672,N_2074,N_2855);
nand U5673 (N_5673,N_3872,N_3681);
nor U5674 (N_5674,N_3937,N_2310);
nand U5675 (N_5675,N_3012,N_3110);
nand U5676 (N_5676,N_3055,N_3330);
or U5677 (N_5677,N_2406,N_3769);
or U5678 (N_5678,N_2933,N_2331);
nor U5679 (N_5679,N_3582,N_3609);
nor U5680 (N_5680,N_3632,N_3220);
or U5681 (N_5681,N_3705,N_2566);
nand U5682 (N_5682,N_3724,N_3732);
and U5683 (N_5683,N_2902,N_3877);
and U5684 (N_5684,N_2144,N_3968);
xnor U5685 (N_5685,N_3091,N_2215);
nor U5686 (N_5686,N_3869,N_3999);
nor U5687 (N_5687,N_3471,N_3107);
and U5688 (N_5688,N_3734,N_3606);
nand U5689 (N_5689,N_3525,N_2318);
or U5690 (N_5690,N_3008,N_3736);
and U5691 (N_5691,N_2843,N_3800);
nor U5692 (N_5692,N_2384,N_2484);
nand U5693 (N_5693,N_3856,N_2412);
or U5694 (N_5694,N_2152,N_3666);
nor U5695 (N_5695,N_3854,N_3127);
nand U5696 (N_5696,N_3038,N_3830);
nor U5697 (N_5697,N_3963,N_3859);
and U5698 (N_5698,N_2486,N_2477);
or U5699 (N_5699,N_3931,N_2484);
nor U5700 (N_5700,N_2439,N_2954);
nand U5701 (N_5701,N_2463,N_2513);
nand U5702 (N_5702,N_2434,N_2371);
nor U5703 (N_5703,N_3247,N_2795);
or U5704 (N_5704,N_2035,N_2777);
and U5705 (N_5705,N_2604,N_3654);
nor U5706 (N_5706,N_2516,N_3192);
nand U5707 (N_5707,N_3699,N_3755);
nand U5708 (N_5708,N_3328,N_3550);
xnor U5709 (N_5709,N_2534,N_3080);
and U5710 (N_5710,N_3572,N_3975);
or U5711 (N_5711,N_3362,N_2416);
or U5712 (N_5712,N_2654,N_2914);
nor U5713 (N_5713,N_2601,N_2180);
and U5714 (N_5714,N_3763,N_3100);
and U5715 (N_5715,N_3676,N_2090);
and U5716 (N_5716,N_3314,N_2952);
nand U5717 (N_5717,N_2440,N_2279);
or U5718 (N_5718,N_2563,N_3379);
xnor U5719 (N_5719,N_3593,N_3062);
and U5720 (N_5720,N_2904,N_3927);
nor U5721 (N_5721,N_3245,N_2670);
or U5722 (N_5722,N_2362,N_3376);
xnor U5723 (N_5723,N_2096,N_2270);
nor U5724 (N_5724,N_2163,N_2386);
and U5725 (N_5725,N_2895,N_3602);
and U5726 (N_5726,N_2137,N_2276);
nor U5727 (N_5727,N_2851,N_3284);
or U5728 (N_5728,N_2583,N_2991);
or U5729 (N_5729,N_2439,N_3929);
nand U5730 (N_5730,N_2269,N_2987);
and U5731 (N_5731,N_2044,N_3270);
or U5732 (N_5732,N_3376,N_2639);
or U5733 (N_5733,N_2444,N_2520);
and U5734 (N_5734,N_3985,N_3647);
and U5735 (N_5735,N_3178,N_2184);
and U5736 (N_5736,N_3833,N_3876);
nand U5737 (N_5737,N_3554,N_3150);
xor U5738 (N_5738,N_2911,N_3303);
nor U5739 (N_5739,N_3141,N_2722);
nand U5740 (N_5740,N_2423,N_3121);
or U5741 (N_5741,N_3309,N_2039);
and U5742 (N_5742,N_3225,N_2570);
nor U5743 (N_5743,N_3012,N_2051);
nand U5744 (N_5744,N_2858,N_3084);
nand U5745 (N_5745,N_2959,N_3535);
nor U5746 (N_5746,N_3223,N_2493);
nand U5747 (N_5747,N_3561,N_2585);
or U5748 (N_5748,N_2365,N_3233);
xnor U5749 (N_5749,N_2599,N_3464);
or U5750 (N_5750,N_2846,N_2099);
or U5751 (N_5751,N_2487,N_2603);
and U5752 (N_5752,N_3526,N_3482);
and U5753 (N_5753,N_2739,N_3450);
or U5754 (N_5754,N_3264,N_2884);
nor U5755 (N_5755,N_3412,N_3070);
nand U5756 (N_5756,N_2406,N_2019);
nand U5757 (N_5757,N_2471,N_3887);
and U5758 (N_5758,N_3842,N_2348);
nand U5759 (N_5759,N_2606,N_3440);
nor U5760 (N_5760,N_2392,N_2233);
and U5761 (N_5761,N_3386,N_2894);
and U5762 (N_5762,N_2120,N_3159);
nor U5763 (N_5763,N_2147,N_2573);
nand U5764 (N_5764,N_2102,N_2752);
or U5765 (N_5765,N_2336,N_3584);
and U5766 (N_5766,N_2890,N_2894);
nor U5767 (N_5767,N_3624,N_2942);
nor U5768 (N_5768,N_3932,N_3873);
nand U5769 (N_5769,N_3066,N_2717);
nor U5770 (N_5770,N_3328,N_2428);
nor U5771 (N_5771,N_2006,N_3826);
nor U5772 (N_5772,N_2466,N_3495);
nor U5773 (N_5773,N_2655,N_3420);
nor U5774 (N_5774,N_3526,N_2580);
nor U5775 (N_5775,N_2915,N_2560);
or U5776 (N_5776,N_2664,N_3905);
nand U5777 (N_5777,N_3691,N_2998);
nand U5778 (N_5778,N_2170,N_3056);
and U5779 (N_5779,N_2887,N_2436);
or U5780 (N_5780,N_2555,N_2268);
nand U5781 (N_5781,N_2658,N_2154);
or U5782 (N_5782,N_2434,N_2105);
nand U5783 (N_5783,N_2500,N_3631);
nand U5784 (N_5784,N_2502,N_3682);
and U5785 (N_5785,N_3025,N_2778);
nand U5786 (N_5786,N_2623,N_2413);
or U5787 (N_5787,N_3919,N_2702);
nand U5788 (N_5788,N_3128,N_2980);
nand U5789 (N_5789,N_2045,N_3020);
and U5790 (N_5790,N_3787,N_2935);
nor U5791 (N_5791,N_2163,N_3178);
or U5792 (N_5792,N_2750,N_2394);
or U5793 (N_5793,N_3135,N_3648);
nor U5794 (N_5794,N_2182,N_2203);
nor U5795 (N_5795,N_2797,N_3044);
nor U5796 (N_5796,N_3359,N_3637);
xnor U5797 (N_5797,N_3370,N_3674);
or U5798 (N_5798,N_3582,N_3973);
nor U5799 (N_5799,N_3062,N_2685);
or U5800 (N_5800,N_3876,N_2347);
or U5801 (N_5801,N_2519,N_3849);
and U5802 (N_5802,N_2110,N_3858);
or U5803 (N_5803,N_3394,N_2508);
nand U5804 (N_5804,N_2285,N_2263);
nand U5805 (N_5805,N_2216,N_2580);
and U5806 (N_5806,N_2945,N_3191);
xor U5807 (N_5807,N_3036,N_2551);
and U5808 (N_5808,N_3506,N_2138);
xnor U5809 (N_5809,N_2324,N_2849);
nand U5810 (N_5810,N_2955,N_2094);
xnor U5811 (N_5811,N_3871,N_2479);
nand U5812 (N_5812,N_3931,N_3883);
nor U5813 (N_5813,N_2790,N_2858);
xnor U5814 (N_5814,N_2588,N_3004);
nand U5815 (N_5815,N_3536,N_3721);
nor U5816 (N_5816,N_3599,N_2264);
and U5817 (N_5817,N_2918,N_3762);
or U5818 (N_5818,N_3065,N_3440);
nand U5819 (N_5819,N_3473,N_3030);
or U5820 (N_5820,N_3619,N_2152);
nor U5821 (N_5821,N_3181,N_3759);
and U5822 (N_5822,N_2897,N_3049);
and U5823 (N_5823,N_2986,N_2931);
nand U5824 (N_5824,N_2789,N_3129);
and U5825 (N_5825,N_2059,N_2907);
xor U5826 (N_5826,N_2122,N_3384);
nand U5827 (N_5827,N_3634,N_3138);
nand U5828 (N_5828,N_3472,N_3565);
or U5829 (N_5829,N_3337,N_2123);
and U5830 (N_5830,N_3311,N_2863);
nor U5831 (N_5831,N_2440,N_2652);
nor U5832 (N_5832,N_2660,N_2608);
xnor U5833 (N_5833,N_2031,N_2282);
nor U5834 (N_5834,N_2525,N_2344);
nor U5835 (N_5835,N_3266,N_2847);
xor U5836 (N_5836,N_3953,N_2021);
or U5837 (N_5837,N_3105,N_2596);
nand U5838 (N_5838,N_2971,N_2500);
xor U5839 (N_5839,N_3692,N_3222);
nor U5840 (N_5840,N_2489,N_3855);
nand U5841 (N_5841,N_2857,N_3072);
or U5842 (N_5842,N_2835,N_3176);
nor U5843 (N_5843,N_3798,N_2098);
nor U5844 (N_5844,N_2324,N_3778);
nor U5845 (N_5845,N_2600,N_2794);
and U5846 (N_5846,N_2698,N_3315);
and U5847 (N_5847,N_2442,N_2761);
or U5848 (N_5848,N_2645,N_2891);
nand U5849 (N_5849,N_2203,N_2005);
or U5850 (N_5850,N_2183,N_3009);
nand U5851 (N_5851,N_2413,N_2409);
or U5852 (N_5852,N_3918,N_3132);
or U5853 (N_5853,N_3950,N_2435);
or U5854 (N_5854,N_3510,N_3238);
nand U5855 (N_5855,N_3214,N_2917);
nor U5856 (N_5856,N_2334,N_3864);
and U5857 (N_5857,N_2946,N_2496);
nand U5858 (N_5858,N_2774,N_3534);
or U5859 (N_5859,N_3595,N_2089);
or U5860 (N_5860,N_3679,N_3397);
and U5861 (N_5861,N_2292,N_3169);
nor U5862 (N_5862,N_2866,N_3362);
or U5863 (N_5863,N_3200,N_3573);
xor U5864 (N_5864,N_3594,N_3324);
nor U5865 (N_5865,N_2067,N_2647);
nor U5866 (N_5866,N_3260,N_3015);
and U5867 (N_5867,N_2066,N_2367);
or U5868 (N_5868,N_3430,N_3883);
and U5869 (N_5869,N_3170,N_3140);
nor U5870 (N_5870,N_3751,N_3696);
nor U5871 (N_5871,N_3167,N_3773);
nor U5872 (N_5872,N_3246,N_3158);
nor U5873 (N_5873,N_2581,N_3755);
and U5874 (N_5874,N_3219,N_3828);
nor U5875 (N_5875,N_3894,N_3508);
nand U5876 (N_5876,N_3251,N_3051);
and U5877 (N_5877,N_3627,N_3972);
and U5878 (N_5878,N_3948,N_2434);
and U5879 (N_5879,N_3960,N_3561);
xnor U5880 (N_5880,N_2286,N_2694);
nand U5881 (N_5881,N_3601,N_2974);
nor U5882 (N_5882,N_3701,N_2635);
nor U5883 (N_5883,N_2273,N_2463);
nand U5884 (N_5884,N_2960,N_3160);
nand U5885 (N_5885,N_3311,N_2624);
nand U5886 (N_5886,N_2403,N_2072);
and U5887 (N_5887,N_3109,N_3728);
nor U5888 (N_5888,N_3925,N_3141);
nor U5889 (N_5889,N_2544,N_3005);
nor U5890 (N_5890,N_2617,N_2686);
xnor U5891 (N_5891,N_3533,N_3724);
nor U5892 (N_5892,N_3498,N_2969);
and U5893 (N_5893,N_2215,N_2805);
and U5894 (N_5894,N_2716,N_2067);
xnor U5895 (N_5895,N_2514,N_2123);
or U5896 (N_5896,N_3594,N_3949);
nor U5897 (N_5897,N_2806,N_2162);
nor U5898 (N_5898,N_3649,N_2818);
or U5899 (N_5899,N_3471,N_2545);
nor U5900 (N_5900,N_3226,N_2855);
or U5901 (N_5901,N_2157,N_2518);
nor U5902 (N_5902,N_3833,N_3741);
nor U5903 (N_5903,N_3775,N_2323);
nor U5904 (N_5904,N_2552,N_2801);
or U5905 (N_5905,N_3046,N_3957);
or U5906 (N_5906,N_2181,N_3667);
and U5907 (N_5907,N_2625,N_2235);
or U5908 (N_5908,N_2182,N_3299);
or U5909 (N_5909,N_3389,N_3139);
nor U5910 (N_5910,N_3819,N_3349);
nor U5911 (N_5911,N_3131,N_2822);
nor U5912 (N_5912,N_3693,N_3536);
nand U5913 (N_5913,N_3798,N_2693);
or U5914 (N_5914,N_3289,N_2318);
and U5915 (N_5915,N_3402,N_3830);
and U5916 (N_5916,N_2779,N_2120);
or U5917 (N_5917,N_2674,N_3035);
nor U5918 (N_5918,N_2349,N_2971);
nor U5919 (N_5919,N_2639,N_2668);
nand U5920 (N_5920,N_2467,N_3281);
nand U5921 (N_5921,N_3880,N_3351);
and U5922 (N_5922,N_3421,N_2479);
nor U5923 (N_5923,N_3327,N_3648);
or U5924 (N_5924,N_2200,N_3462);
or U5925 (N_5925,N_3081,N_2805);
nand U5926 (N_5926,N_3324,N_2630);
or U5927 (N_5927,N_2837,N_2687);
nand U5928 (N_5928,N_2803,N_2106);
nor U5929 (N_5929,N_3616,N_2065);
nand U5930 (N_5930,N_3192,N_2876);
and U5931 (N_5931,N_2967,N_2054);
nor U5932 (N_5932,N_3676,N_3872);
xor U5933 (N_5933,N_3801,N_3928);
nand U5934 (N_5934,N_3859,N_2345);
nor U5935 (N_5935,N_3293,N_2631);
or U5936 (N_5936,N_3080,N_3826);
nor U5937 (N_5937,N_2315,N_2399);
nor U5938 (N_5938,N_2297,N_2904);
xnor U5939 (N_5939,N_3451,N_2177);
or U5940 (N_5940,N_2898,N_3071);
xnor U5941 (N_5941,N_3235,N_3846);
nand U5942 (N_5942,N_3603,N_3689);
nor U5943 (N_5943,N_2031,N_3731);
and U5944 (N_5944,N_2227,N_3539);
nand U5945 (N_5945,N_2572,N_3634);
and U5946 (N_5946,N_2049,N_2297);
or U5947 (N_5947,N_2207,N_3397);
nor U5948 (N_5948,N_2940,N_2648);
xnor U5949 (N_5949,N_2357,N_2096);
or U5950 (N_5950,N_2983,N_3913);
and U5951 (N_5951,N_3674,N_3279);
and U5952 (N_5952,N_3625,N_2596);
nor U5953 (N_5953,N_2429,N_3666);
nand U5954 (N_5954,N_3303,N_2908);
nand U5955 (N_5955,N_2027,N_2747);
nor U5956 (N_5956,N_3392,N_2719);
nand U5957 (N_5957,N_2385,N_3576);
nor U5958 (N_5958,N_2411,N_3607);
or U5959 (N_5959,N_2955,N_2138);
or U5960 (N_5960,N_2512,N_2977);
and U5961 (N_5961,N_3785,N_2031);
xor U5962 (N_5962,N_2656,N_2413);
nor U5963 (N_5963,N_3201,N_2072);
or U5964 (N_5964,N_3732,N_3226);
xor U5965 (N_5965,N_2360,N_2833);
nand U5966 (N_5966,N_3597,N_2211);
and U5967 (N_5967,N_2790,N_2987);
nand U5968 (N_5968,N_3007,N_2229);
or U5969 (N_5969,N_3318,N_3913);
or U5970 (N_5970,N_2314,N_2612);
and U5971 (N_5971,N_2120,N_3946);
nor U5972 (N_5972,N_2608,N_3322);
nor U5973 (N_5973,N_2568,N_2754);
xnor U5974 (N_5974,N_3497,N_3543);
nor U5975 (N_5975,N_3201,N_2499);
and U5976 (N_5976,N_3833,N_2903);
or U5977 (N_5977,N_2661,N_2000);
nand U5978 (N_5978,N_3852,N_2650);
nand U5979 (N_5979,N_3945,N_2238);
or U5980 (N_5980,N_2607,N_2754);
or U5981 (N_5981,N_3206,N_3055);
nand U5982 (N_5982,N_2565,N_3498);
nand U5983 (N_5983,N_3171,N_2479);
nor U5984 (N_5984,N_3434,N_3331);
nor U5985 (N_5985,N_3651,N_2024);
and U5986 (N_5986,N_3550,N_3003);
nor U5987 (N_5987,N_3631,N_3860);
xor U5988 (N_5988,N_2250,N_2463);
or U5989 (N_5989,N_3763,N_3617);
and U5990 (N_5990,N_3110,N_2213);
xor U5991 (N_5991,N_3396,N_2196);
and U5992 (N_5992,N_3587,N_2180);
and U5993 (N_5993,N_2251,N_3283);
xnor U5994 (N_5994,N_3908,N_2008);
or U5995 (N_5995,N_2560,N_3414);
nor U5996 (N_5996,N_2145,N_3544);
nor U5997 (N_5997,N_3454,N_2944);
and U5998 (N_5998,N_2849,N_2314);
nand U5999 (N_5999,N_2741,N_3498);
nor U6000 (N_6000,N_5646,N_5816);
and U6001 (N_6001,N_4498,N_5267);
or U6002 (N_6002,N_4957,N_4768);
nor U6003 (N_6003,N_4635,N_5985);
nand U6004 (N_6004,N_4572,N_5615);
or U6005 (N_6005,N_4160,N_4342);
nand U6006 (N_6006,N_5043,N_5122);
nand U6007 (N_6007,N_4774,N_4711);
and U6008 (N_6008,N_4413,N_5663);
nand U6009 (N_6009,N_4912,N_5876);
and U6010 (N_6010,N_5849,N_4049);
xor U6011 (N_6011,N_5319,N_5717);
nor U6012 (N_6012,N_5589,N_5020);
or U6013 (N_6013,N_4826,N_4325);
nand U6014 (N_6014,N_5834,N_4421);
or U6015 (N_6015,N_4204,N_4011);
or U6016 (N_6016,N_5377,N_5993);
and U6017 (N_6017,N_4257,N_5396);
xor U6018 (N_6018,N_5782,N_4535);
nor U6019 (N_6019,N_4215,N_5069);
nand U6020 (N_6020,N_4344,N_4240);
nand U6021 (N_6021,N_5071,N_4149);
nor U6022 (N_6022,N_5364,N_4391);
and U6023 (N_6023,N_5225,N_4403);
nand U6024 (N_6024,N_5897,N_5180);
nand U6025 (N_6025,N_5019,N_4546);
and U6026 (N_6026,N_4782,N_5945);
nand U6027 (N_6027,N_5832,N_4500);
nor U6028 (N_6028,N_5450,N_4292);
nor U6029 (N_6029,N_5779,N_4184);
and U6030 (N_6030,N_5695,N_4566);
nor U6031 (N_6031,N_4241,N_4616);
or U6032 (N_6032,N_5156,N_5508);
and U6033 (N_6033,N_4688,N_4940);
or U6034 (N_6034,N_4856,N_5644);
and U6035 (N_6035,N_5096,N_4908);
nand U6036 (N_6036,N_4933,N_5979);
or U6037 (N_6037,N_4227,N_5766);
nor U6038 (N_6038,N_5523,N_5463);
and U6039 (N_6039,N_4474,N_4612);
nand U6040 (N_6040,N_5098,N_4066);
nand U6041 (N_6041,N_4407,N_5776);
nand U6042 (N_6042,N_4857,N_4626);
nand U6043 (N_6043,N_4520,N_5496);
or U6044 (N_6044,N_5602,N_5103);
nand U6045 (N_6045,N_5517,N_5906);
xnor U6046 (N_6046,N_5253,N_4107);
nand U6047 (N_6047,N_5397,N_5207);
and U6048 (N_6048,N_4914,N_4586);
nor U6049 (N_6049,N_4036,N_5183);
or U6050 (N_6050,N_4271,N_5754);
nor U6051 (N_6051,N_5748,N_4420);
or U6052 (N_6052,N_5539,N_4796);
xor U6053 (N_6053,N_5248,N_5210);
nand U6054 (N_6054,N_5339,N_5120);
or U6055 (N_6055,N_4147,N_5469);
xnor U6056 (N_6056,N_4248,N_5407);
xor U6057 (N_6057,N_5161,N_5965);
or U6058 (N_6058,N_5164,N_5522);
nor U6059 (N_6059,N_4671,N_5574);
nand U6060 (N_6060,N_4358,N_5940);
or U6061 (N_6061,N_5318,N_4552);
xnor U6062 (N_6062,N_4141,N_5640);
and U6063 (N_6063,N_4966,N_5234);
nor U6064 (N_6064,N_4697,N_4724);
nand U6065 (N_6065,N_5725,N_5813);
and U6066 (N_6066,N_5184,N_4916);
or U6067 (N_6067,N_5817,N_5006);
or U6068 (N_6068,N_5636,N_5295);
or U6069 (N_6069,N_4847,N_5492);
nor U6070 (N_6070,N_4035,N_4621);
nor U6071 (N_6071,N_4641,N_4991);
nor U6072 (N_6072,N_4319,N_5730);
or U6073 (N_6073,N_4866,N_5034);
nand U6074 (N_6074,N_5514,N_4867);
and U6075 (N_6075,N_5625,N_4939);
nand U6076 (N_6076,N_4935,N_5360);
nand U6077 (N_6077,N_5053,N_4414);
nand U6078 (N_6078,N_4009,N_5200);
nor U6079 (N_6079,N_4506,N_4938);
or U6080 (N_6080,N_5938,N_4728);
xor U6081 (N_6081,N_4052,N_5510);
xnor U6082 (N_6082,N_5969,N_5280);
or U6083 (N_6083,N_4547,N_5762);
nor U6084 (N_6084,N_4484,N_4622);
and U6085 (N_6085,N_5935,N_4575);
or U6086 (N_6086,N_5362,N_5356);
nand U6087 (N_6087,N_4835,N_4401);
nor U6088 (N_6088,N_5307,N_4695);
xnor U6089 (N_6089,N_4639,N_5209);
and U6090 (N_6090,N_4814,N_5128);
nand U6091 (N_6091,N_4915,N_4368);
or U6092 (N_6092,N_5224,N_4214);
or U6093 (N_6093,N_5269,N_5076);
nor U6094 (N_6094,N_4383,N_4279);
and U6095 (N_6095,N_4651,N_5214);
and U6096 (N_6096,N_4744,N_4999);
nand U6097 (N_6097,N_5949,N_5216);
or U6098 (N_6098,N_4684,N_5616);
or U6099 (N_6099,N_5278,N_4462);
or U6100 (N_6100,N_4128,N_5500);
nor U6101 (N_6101,N_5349,N_4712);
nor U6102 (N_6102,N_5221,N_4137);
and U6103 (N_6103,N_4369,N_4628);
xor U6104 (N_6104,N_4540,N_4820);
nand U6105 (N_6105,N_5205,N_4627);
nor U6106 (N_6106,N_5871,N_5786);
nor U6107 (N_6107,N_5062,N_4256);
nor U6108 (N_6108,N_5327,N_5434);
or U6109 (N_6109,N_4564,N_4919);
nand U6110 (N_6110,N_5996,N_4062);
and U6111 (N_6111,N_5881,N_4336);
nand U6112 (N_6112,N_4219,N_5037);
xor U6113 (N_6113,N_4188,N_4771);
nor U6114 (N_6114,N_4941,N_4217);
or U6115 (N_6115,N_5070,N_5721);
nand U6116 (N_6116,N_5808,N_4258);
xor U6117 (N_6117,N_4901,N_4040);
or U6118 (N_6118,N_5647,N_5376);
nand U6119 (N_6119,N_4466,N_5995);
xor U6120 (N_6120,N_5271,N_5094);
or U6121 (N_6121,N_5005,N_4903);
or U6122 (N_6122,N_4296,N_4558);
xnor U6123 (N_6123,N_4291,N_4801);
nor U6124 (N_6124,N_5846,N_4508);
or U6125 (N_6125,N_5987,N_5722);
or U6126 (N_6126,N_4163,N_5954);
xnor U6127 (N_6127,N_4422,N_5951);
xor U6128 (N_6128,N_4216,N_4758);
xnor U6129 (N_6129,N_5038,N_4173);
xnor U6130 (N_6130,N_5102,N_5873);
nand U6131 (N_6131,N_4494,N_4755);
nor U6132 (N_6132,N_5335,N_5825);
or U6133 (N_6133,N_4287,N_5710);
xor U6134 (N_6134,N_4829,N_5892);
nand U6135 (N_6135,N_4849,N_5798);
nand U6136 (N_6136,N_5943,N_4263);
nand U6137 (N_6137,N_5361,N_4518);
and U6138 (N_6138,N_5761,N_5989);
nor U6139 (N_6139,N_4254,N_4813);
and U6140 (N_6140,N_5139,N_4614);
nand U6141 (N_6141,N_4117,N_4417);
or U6142 (N_6142,N_4511,N_5471);
or U6143 (N_6143,N_5066,N_4155);
and U6144 (N_6144,N_4306,N_4838);
nor U6145 (N_6145,N_5691,N_5457);
or U6146 (N_6146,N_4010,N_4153);
or U6147 (N_6147,N_4003,N_4436);
nor U6148 (N_6148,N_4580,N_5676);
or U6149 (N_6149,N_5187,N_5934);
nor U6150 (N_6150,N_5971,N_5412);
and U6151 (N_6151,N_5836,N_5991);
and U6152 (N_6152,N_5733,N_4893);
nor U6153 (N_6153,N_4174,N_5803);
and U6154 (N_6154,N_4557,N_5903);
nor U6155 (N_6155,N_4289,N_5932);
nand U6156 (N_6156,N_5445,N_5521);
xnor U6157 (N_6157,N_4677,N_4095);
nand U6158 (N_6158,N_5581,N_4778);
nand U6159 (N_6159,N_4666,N_5812);
and U6160 (N_6160,N_5531,N_5305);
xnor U6161 (N_6161,N_4740,N_5894);
nand U6162 (N_6162,N_5824,N_5952);
and U6163 (N_6163,N_5865,N_5707);
nand U6164 (N_6164,N_5970,N_5345);
or U6165 (N_6165,N_4603,N_5957);
or U6166 (N_6166,N_4058,N_5661);
xnor U6167 (N_6167,N_4555,N_4370);
nor U6168 (N_6168,N_4673,N_4875);
or U6169 (N_6169,N_5171,N_4583);
nor U6170 (N_6170,N_4016,N_5668);
nor U6171 (N_6171,N_5000,N_5092);
or U6172 (N_6172,N_5742,N_4180);
nand U6173 (N_6173,N_5618,N_4119);
nand U6174 (N_6174,N_5322,N_4069);
or U6175 (N_6175,N_4763,N_4834);
nand U6176 (N_6176,N_5314,N_5313);
or U6177 (N_6177,N_4101,N_4199);
nand U6178 (N_6178,N_4109,N_4410);
nand U6179 (N_6179,N_5308,N_4455);
nand U6180 (N_6180,N_5487,N_4309);
and U6181 (N_6181,N_5501,N_4642);
nand U6182 (N_6182,N_4266,N_4568);
or U6183 (N_6183,N_5788,N_4683);
nand U6184 (N_6184,N_4994,N_5587);
nand U6185 (N_6185,N_4221,N_4238);
nor U6186 (N_6186,N_5276,N_4176);
nand U6187 (N_6187,N_5185,N_5545);
nor U6188 (N_6188,N_4441,N_5226);
and U6189 (N_6189,N_5494,N_4571);
nand U6190 (N_6190,N_5720,N_5870);
nand U6191 (N_6191,N_5368,N_5114);
nand U6192 (N_6192,N_5666,N_5775);
nor U6193 (N_6193,N_5763,N_5099);
nor U6194 (N_6194,N_4738,N_4657);
or U6195 (N_6195,N_5435,N_4504);
or U6196 (N_6196,N_4213,N_4439);
nand U6197 (N_6197,N_4476,N_4708);
and U6198 (N_6198,N_5270,N_5538);
or U6199 (N_6199,N_5268,N_5734);
nor U6200 (N_6200,N_5402,N_4819);
and U6201 (N_6201,N_5452,N_4633);
nor U6202 (N_6202,N_4911,N_4091);
nor U6203 (N_6203,N_4977,N_4440);
and U6204 (N_6204,N_5854,N_4780);
nor U6205 (N_6205,N_4831,N_5049);
and U6206 (N_6206,N_4950,N_4717);
and U6207 (N_6207,N_5771,N_5374);
and U6208 (N_6208,N_5190,N_4843);
nor U6209 (N_6209,N_4607,N_5712);
nand U6210 (N_6210,N_5163,N_4136);
nand U6211 (N_6211,N_4273,N_5424);
xor U6212 (N_6212,N_5263,N_5518);
or U6213 (N_6213,N_4793,N_5512);
and U6214 (N_6214,N_4051,N_4714);
xor U6215 (N_6215,N_5036,N_4262);
or U6216 (N_6216,N_4970,N_5048);
nor U6217 (N_6217,N_5760,N_4519);
or U6218 (N_6218,N_5641,N_4467);
or U6219 (N_6219,N_5626,N_4874);
xor U6220 (N_6220,N_4952,N_5016);
nor U6221 (N_6221,N_4929,N_5199);
xor U6222 (N_6222,N_4301,N_5474);
nor U6223 (N_6223,N_5600,N_4753);
or U6224 (N_6224,N_4672,N_4170);
and U6225 (N_6225,N_5783,N_5887);
or U6226 (N_6226,N_5547,N_4037);
or U6227 (N_6227,N_4553,N_4667);
or U6228 (N_6228,N_5548,N_5148);
or U6229 (N_6229,N_4524,N_5843);
and U6230 (N_6230,N_5012,N_4779);
nor U6231 (N_6231,N_5426,N_5673);
nor U6232 (N_6232,N_4503,N_4249);
or U6233 (N_6233,N_4533,N_5429);
xnor U6234 (N_6234,N_4121,N_5388);
or U6235 (N_6235,N_4559,N_5853);
nand U6236 (N_6236,N_4944,N_5298);
or U6237 (N_6237,N_4828,N_4756);
nor U6238 (N_6238,N_4250,N_4807);
or U6239 (N_6239,N_5680,N_5557);
nor U6240 (N_6240,N_5525,N_5166);
nor U6241 (N_6241,N_4270,N_5389);
or U6242 (N_6242,N_4139,N_4229);
nor U6243 (N_6243,N_5242,N_4550);
nand U6244 (N_6244,N_4638,N_5095);
xor U6245 (N_6245,N_5024,N_4146);
xor U6246 (N_6246,N_5653,N_5632);
nor U6247 (N_6247,N_4936,N_5528);
and U6248 (N_6248,N_5919,N_4345);
and U6249 (N_6249,N_5874,N_5579);
and U6250 (N_6250,N_5231,N_4761);
nor U6251 (N_6251,N_4472,N_4767);
nand U6252 (N_6252,N_4839,N_4375);
and U6253 (N_6253,N_5976,N_4745);
nor U6254 (N_6254,N_4127,N_4031);
and U6255 (N_6255,N_4716,N_5802);
nand U6256 (N_6256,N_5009,N_4563);
or U6257 (N_6257,N_4093,N_5709);
xor U6258 (N_6258,N_5146,N_4205);
and U6259 (N_6259,N_5244,N_5915);
and U6260 (N_6260,N_4433,N_5840);
or U6261 (N_6261,N_4600,N_5460);
nand U6262 (N_6262,N_5273,N_5756);
or U6263 (N_6263,N_4418,N_4934);
xnor U6264 (N_6264,N_4220,N_5913);
and U6265 (N_6265,N_4398,N_4971);
nor U6266 (N_6266,N_4192,N_4181);
nand U6267 (N_6267,N_4430,N_5567);
or U6268 (N_6268,N_5385,N_5461);
nor U6269 (N_6269,N_5340,N_5240);
xnor U6270 (N_6270,N_5638,N_4754);
or U6271 (N_6271,N_4788,N_5559);
and U6272 (N_6272,N_5112,N_4024);
or U6273 (N_6273,N_4083,N_4060);
or U6274 (N_6274,N_5784,N_4231);
nand U6275 (N_6275,N_5852,N_4085);
and U6276 (N_6276,N_5065,N_4191);
nand U6277 (N_6277,N_5084,N_4570);
and U6278 (N_6278,N_4589,N_4623);
nor U6279 (N_6279,N_5681,N_4860);
or U6280 (N_6280,N_4056,N_5654);
or U6281 (N_6281,N_4619,N_5835);
or U6282 (N_6282,N_4833,N_5930);
nand U6283 (N_6283,N_5162,N_4159);
xnor U6284 (N_6284,N_4759,N_4898);
xnor U6285 (N_6285,N_4327,N_4526);
nor U6286 (N_6286,N_5830,N_5558);
nor U6287 (N_6287,N_5077,N_4615);
or U6288 (N_6288,N_4885,N_5131);
and U6289 (N_6289,N_4513,N_5260);
or U6290 (N_6290,N_5685,N_4481);
and U6291 (N_6291,N_4497,N_5612);
xor U6292 (N_6292,N_5002,N_4475);
and U6293 (N_6293,N_5885,N_5079);
nor U6294 (N_6294,N_4090,N_4340);
nor U6295 (N_6295,N_5841,N_5201);
xnor U6296 (N_6296,N_4380,N_5966);
or U6297 (N_6297,N_4084,N_5540);
xnor U6298 (N_6298,N_4193,N_5369);
or U6299 (N_6299,N_4203,N_4543);
xor U6300 (N_6300,N_4110,N_5399);
nand U6301 (N_6301,N_5904,N_4073);
nand U6302 (N_6302,N_4223,N_5342);
nand U6303 (N_6303,N_4371,N_5081);
and U6304 (N_6304,N_5806,N_4076);
nor U6305 (N_6305,N_5609,N_4208);
nor U6306 (N_6306,N_5110,N_4643);
nor U6307 (N_6307,N_5354,N_5197);
or U6308 (N_6308,N_5891,N_4341);
nor U6309 (N_6309,N_5366,N_4794);
and U6310 (N_6310,N_5866,N_5477);
and U6311 (N_6311,N_4842,N_4979);
nand U6312 (N_6312,N_4865,N_5439);
nor U6313 (N_6313,N_5029,N_5575);
nor U6314 (N_6314,N_5441,N_4313);
or U6315 (N_6315,N_5889,N_4048);
nor U6316 (N_6316,N_5879,N_4267);
nand U6317 (N_6317,N_4783,N_5422);
or U6318 (N_6318,N_5400,N_5455);
and U6319 (N_6319,N_5410,N_4545);
nor U6320 (N_6320,N_4588,N_5370);
or U6321 (N_6321,N_5583,N_4918);
nand U6322 (N_6322,N_4715,N_5924);
or U6323 (N_6323,N_5054,N_5864);
nor U6324 (N_6324,N_4157,N_5246);
or U6325 (N_6325,N_4485,N_4293);
nor U6326 (N_6326,N_4000,N_5704);
or U6327 (N_6327,N_5759,N_5427);
and U6328 (N_6328,N_5978,N_5923);
nand U6329 (N_6329,N_5614,N_5634);
or U6330 (N_6330,N_5927,N_4499);
or U6331 (N_6331,N_4057,N_5886);
nor U6332 (N_6332,N_4517,N_4253);
and U6333 (N_6333,N_5279,N_4338);
and U6334 (N_6334,N_5697,N_5014);
nand U6335 (N_6335,N_4297,N_4791);
or U6336 (N_6336,N_5981,N_4649);
and U6337 (N_6337,N_5315,N_5551);
xor U6338 (N_6338,N_5810,N_4265);
nand U6339 (N_6339,N_5117,N_4453);
nor U6340 (N_6340,N_4171,N_4429);
and U6341 (N_6341,N_4438,N_4165);
or U6342 (N_6342,N_4007,N_5888);
nand U6343 (N_6343,N_5105,N_4769);
nand U6344 (N_6344,N_5045,N_5287);
xnor U6345 (N_6345,N_4144,N_5630);
and U6346 (N_6346,N_4512,N_4790);
nand U6347 (N_6347,N_4804,N_5091);
or U6348 (N_6348,N_5617,N_5723);
or U6349 (N_6349,N_5419,N_4131);
nand U6350 (N_6350,N_4665,N_5905);
nor U6351 (N_6351,N_5532,N_5300);
nand U6352 (N_6352,N_4749,N_4937);
nor U6353 (N_6353,N_5140,N_4393);
nand U6354 (N_6354,N_4594,N_5144);
xnor U6355 (N_6355,N_4675,N_4284);
nor U6356 (N_6356,N_5700,N_5994);
nand U6357 (N_6357,N_4881,N_5807);
and U6358 (N_6358,N_5296,N_5107);
and U6359 (N_6359,N_4283,N_4674);
or U6360 (N_6360,N_5908,N_4739);
or U6361 (N_6361,N_4063,N_4987);
or U6362 (N_6362,N_4005,N_4887);
or U6363 (N_6363,N_5819,N_5650);
and U6364 (N_6364,N_5423,N_5421);
and U6365 (N_6365,N_5777,N_5683);
and U6366 (N_6366,N_4925,N_5556);
xor U6367 (N_6367,N_5344,N_4798);
xor U6368 (N_6368,N_5046,N_5309);
xor U6369 (N_6369,N_4045,N_5693);
and U6370 (N_6370,N_5250,N_5605);
nor U6371 (N_6371,N_4362,N_5708);
nand U6372 (N_6372,N_5592,N_4955);
nor U6373 (N_6373,N_5359,N_4502);
or U6374 (N_6374,N_4921,N_5925);
xnor U6375 (N_6375,N_4676,N_5235);
xnor U6376 (N_6376,N_4900,N_4479);
or U6377 (N_6377,N_4687,N_5506);
and U6378 (N_6378,N_5249,N_5677);
nand U6379 (N_6379,N_5288,N_5468);
and U6380 (N_6380,N_5052,N_5115);
nor U6381 (N_6381,N_5774,N_5057);
or U6382 (N_6382,N_4315,N_4509);
nand U6383 (N_6383,N_5619,N_5293);
xor U6384 (N_6384,N_4581,N_4452);
nor U6385 (N_6385,N_4274,N_4510);
nand U6386 (N_6386,N_4120,N_4932);
nand U6387 (N_6387,N_4967,N_4894);
nand U6388 (N_6388,N_5990,N_4008);
xnor U6389 (N_6389,N_4844,N_5526);
and U6390 (N_6390,N_5651,N_4766);
nand U6391 (N_6391,N_4544,N_4473);
xnor U6392 (N_6392,N_4548,N_5203);
or U6393 (N_6393,N_4681,N_4596);
and U6394 (N_6394,N_5003,N_4593);
nor U6395 (N_6395,N_5138,N_5236);
or U6396 (N_6396,N_4608,N_4388);
and U6397 (N_6397,N_5484,N_5660);
and U6398 (N_6398,N_4597,N_4152);
and U6399 (N_6399,N_5382,N_5025);
and U6400 (N_6400,N_4978,N_4381);
xnor U6401 (N_6401,N_4815,N_5855);
and U6402 (N_6402,N_4549,N_5233);
or U6403 (N_6403,N_5750,N_4721);
and U6404 (N_6404,N_5620,N_4537);
and U6405 (N_6405,N_4686,N_5237);
nand U6406 (N_6406,N_4140,N_5974);
nor U6407 (N_6407,N_5648,N_5039);
nor U6408 (N_6408,N_4311,N_4222);
and U6409 (N_6409,N_4318,N_4990);
nor U6410 (N_6410,N_4108,N_4074);
nand U6411 (N_6411,N_5372,N_5223);
and U6412 (N_6412,N_4142,N_5998);
and U6413 (N_6413,N_5737,N_4400);
nor U6414 (N_6414,N_4660,N_5432);
and U6415 (N_6415,N_4760,N_5827);
or U6416 (N_6416,N_4624,N_5061);
nor U6417 (N_6417,N_5780,N_4825);
or U6418 (N_6418,N_4189,N_5656);
or U6419 (N_6419,N_4878,N_5311);
and U6420 (N_6420,N_5153,N_4737);
or U6421 (N_6421,N_5466,N_5675);
nand U6422 (N_6422,N_4604,N_5912);
xnor U6423 (N_6423,N_5631,N_5502);
and U6424 (N_6424,N_4995,N_4840);
and U6425 (N_6425,N_5160,N_4425);
nor U6426 (N_6426,N_5628,N_4059);
or U6427 (N_6427,N_5021,N_4662);
nand U6428 (N_6428,N_4832,N_4072);
nor U6429 (N_6429,N_4488,N_5391);
and U6430 (N_6430,N_4985,N_5983);
or U6431 (N_6431,N_5174,N_4379);
nand U6432 (N_6432,N_5804,N_5482);
nand U6433 (N_6433,N_4496,N_4285);
and U6434 (N_6434,N_5056,N_5732);
or U6435 (N_6435,N_5509,N_5627);
and U6436 (N_6436,N_4126,N_5047);
nor U6437 (N_6437,N_4068,N_4312);
nand U6438 (N_6438,N_4435,N_4680);
and U6439 (N_6439,N_4786,N_5503);
nand U6440 (N_6440,N_5607,N_5895);
or U6441 (N_6441,N_5202,N_5304);
and U6442 (N_6442,N_4194,N_5652);
nand U6443 (N_6443,N_5393,N_5394);
nor U6444 (N_6444,N_4411,N_5584);
or U6445 (N_6445,N_5050,N_5831);
or U6446 (N_6446,N_5448,N_5169);
xor U6447 (N_6447,N_4487,N_4079);
nand U6448 (N_6448,N_5303,N_5358);
nor U6449 (N_6449,N_4732,N_4992);
or U6450 (N_6450,N_4478,N_5821);
or U6451 (N_6451,N_4752,N_4884);
xor U6452 (N_6452,N_4864,N_4777);
nand U6453 (N_6453,N_5338,N_5568);
nor U6454 (N_6454,N_4648,N_5022);
nor U6455 (N_6455,N_5942,N_5937);
nor U6456 (N_6456,N_4006,N_5189);
nand U6457 (N_6457,N_5962,N_5111);
nand U6458 (N_6458,N_4924,N_4501);
nand U6459 (N_6459,N_4308,N_5520);
nor U6460 (N_6460,N_4288,N_5769);
nand U6461 (N_6461,N_4295,N_4799);
and U6462 (N_6462,N_4605,N_4225);
nand U6463 (N_6463,N_5753,N_5515);
nand U6464 (N_6464,N_4196,N_5436);
or U6465 (N_6465,N_5247,N_4902);
xnor U6466 (N_6466,N_4945,N_4047);
and U6467 (N_6467,N_5489,N_4098);
or U6468 (N_6468,N_4354,N_5026);
or U6469 (N_6469,N_5067,N_5724);
nor U6470 (N_6470,N_4742,N_4450);
nand U6471 (N_6471,N_4404,N_4792);
nand U6472 (N_6472,N_4891,N_5013);
xor U6473 (N_6473,N_5384,N_5772);
nor U6474 (N_6474,N_5588,N_5752);
nor U6475 (N_6475,N_5473,N_5542);
nor U6476 (N_6476,N_5191,N_4187);
and U6477 (N_6477,N_4879,N_5544);
and U6478 (N_6478,N_4348,N_5524);
and U6479 (N_6479,N_5297,N_5175);
xnor U6480 (N_6480,N_5837,N_5578);
nor U6481 (N_6481,N_4100,N_5467);
nor U6482 (N_6482,N_4456,N_4961);
and U6483 (N_6483,N_4409,N_4726);
xor U6484 (N_6484,N_4800,N_4963);
or U6485 (N_6485,N_4175,N_5472);
or U6486 (N_6486,N_4416,N_4569);
xnor U6487 (N_6487,N_5089,N_4853);
and U6488 (N_6488,N_4361,N_4346);
or U6489 (N_6489,N_4423,N_4233);
or U6490 (N_6490,N_5916,N_4197);
nand U6491 (N_6491,N_4625,N_4521);
or U6492 (N_6492,N_4565,N_5306);
nor U6493 (N_6493,N_5491,N_4706);
xor U6494 (N_6494,N_5289,N_5714);
and U6495 (N_6495,N_5667,N_5058);
xor U6496 (N_6496,N_5814,N_5192);
nand U6497 (N_6497,N_5001,N_4670);
nand U6498 (N_6498,N_4631,N_5483);
nand U6499 (N_6499,N_5688,N_4718);
nor U6500 (N_6500,N_4969,N_4177);
or U6501 (N_6501,N_5324,N_5475);
and U6502 (N_6502,N_4574,N_4378);
nor U6503 (N_6503,N_5820,N_5686);
nand U6504 (N_6504,N_5655,N_4154);
and U6505 (N_6505,N_5861,N_5736);
and U6506 (N_6506,N_4071,N_4179);
xnor U6507 (N_6507,N_4195,N_4953);
or U6508 (N_6508,N_5499,N_5317);
or U6509 (N_6509,N_5251,N_5698);
xnor U6510 (N_6510,N_5797,N_5860);
xor U6511 (N_6511,N_5035,N_5571);
nand U6512 (N_6512,N_5256,N_5074);
nor U6513 (N_6513,N_4664,N_5425);
nand U6514 (N_6514,N_5862,N_4705);
nand U6515 (N_6515,N_4269,N_4931);
xnor U6516 (N_6516,N_5433,N_5590);
and U6517 (N_6517,N_4164,N_5124);
or U6518 (N_6518,N_4920,N_4172);
xnor U6519 (N_6519,N_4682,N_5657);
xnor U6520 (N_6520,N_5629,N_4629);
or U6521 (N_6521,N_4002,N_5893);
nand U6522 (N_6522,N_5684,N_4850);
and U6523 (N_6523,N_5516,N_5126);
and U6524 (N_6524,N_4463,N_5416);
nor U6525 (N_6525,N_4039,N_5261);
nand U6526 (N_6526,N_5781,N_4542);
nand U6527 (N_6527,N_5222,N_4691);
nand U6528 (N_6528,N_4202,N_4445);
nand U6529 (N_6529,N_4294,N_5476);
xnor U6530 (N_6530,N_5392,N_4235);
nor U6531 (N_6531,N_5386,N_4480);
nand U6532 (N_6532,N_4408,N_5706);
xor U6533 (N_6533,N_4352,N_5123);
and U6534 (N_6534,N_4789,N_5087);
nor U6535 (N_6535,N_4845,N_5449);
nor U6536 (N_6536,N_5580,N_5595);
nand U6537 (N_6537,N_5404,N_4679);
nand U6538 (N_6538,N_5444,N_5529);
and U6539 (N_6539,N_4367,N_4514);
nand U6540 (N_6540,N_5611,N_5086);
nor U6541 (N_6541,N_4030,N_5842);
and U6542 (N_6542,N_5051,N_4471);
nand U6543 (N_6543,N_4947,N_4236);
nor U6544 (N_6544,N_5859,N_4041);
nor U6545 (N_6545,N_5662,N_5428);
nand U6546 (N_6546,N_4951,N_4946);
or U6547 (N_6547,N_4734,N_5999);
or U6548 (N_6548,N_5920,N_4329);
or U6549 (N_6549,N_4114,N_4088);
nor U6550 (N_6550,N_4129,N_4310);
nand U6551 (N_6551,N_4888,N_5555);
and U6552 (N_6552,N_5778,N_4525);
nor U6553 (N_6553,N_5690,N_5911);
nand U6554 (N_6554,N_5848,N_4700);
and U6555 (N_6555,N_4178,N_4803);
or U6556 (N_6556,N_5847,N_4102);
nor U6557 (N_6557,N_5554,N_4356);
and U6558 (N_6558,N_5984,N_4252);
xnor U6559 (N_6559,N_4025,N_4337);
nor U6560 (N_6560,N_4873,N_4145);
xor U6561 (N_6561,N_5168,N_5552);
or U6562 (N_6562,N_4019,N_4067);
xnor U6563 (N_6563,N_5534,N_5975);
or U6564 (N_6564,N_4655,N_5505);
nor U6565 (N_6565,N_4246,N_5687);
xor U6566 (N_6566,N_5758,N_5299);
and U6567 (N_6567,N_5645,N_5451);
nand U6568 (N_6568,N_4810,N_4928);
or U6569 (N_6569,N_5822,N_5563);
nand U6570 (N_6570,N_5910,N_4713);
and U6571 (N_6571,N_5909,N_5497);
and U6572 (N_6572,N_5258,N_4134);
and U6573 (N_6573,N_5597,N_5219);
nand U6574 (N_6574,N_4895,N_5206);
nand U6575 (N_6575,N_4446,N_4906);
or U6576 (N_6576,N_4748,N_4989);
nor U6577 (N_6577,N_4851,N_5877);
or U6578 (N_6578,N_4904,N_5958);
nor U6579 (N_6579,N_5254,N_5703);
and U6580 (N_6580,N_5674,N_5792);
or U6581 (N_6581,N_4364,N_5643);
nand U6582 (N_6582,N_4261,N_5245);
nor U6583 (N_6583,N_4426,N_5430);
nor U6584 (N_6584,N_4143,N_4694);
nand U6585 (N_6585,N_4988,N_4078);
nor U6586 (N_6586,N_4601,N_5694);
nand U6587 (N_6587,N_4852,N_5790);
nor U6588 (N_6588,N_4573,N_5390);
or U6589 (N_6589,N_4659,N_5561);
and U6590 (N_6590,N_4018,N_4405);
xnor U6591 (N_6591,N_5576,N_5329);
xnor U6592 (N_6592,N_5333,N_5310);
and U6593 (N_6593,N_4802,N_4636);
nand U6594 (N_6594,N_5495,N_4650);
nand U6595 (N_6595,N_4943,N_5353);
nand U6596 (N_6596,N_5157,N_4489);
nor U6597 (N_6597,N_4861,N_5409);
nor U6598 (N_6598,N_4775,N_4247);
nor U6599 (N_6599,N_5642,N_5716);
xor U6600 (N_6600,N_4054,N_5281);
or U6601 (N_6601,N_5980,N_4723);
nor U6602 (N_6602,N_5977,N_4166);
and U6603 (N_6603,N_5383,N_5182);
nand U6604 (N_6604,N_4731,N_5063);
nor U6605 (N_6605,N_4206,N_4394);
and U6606 (N_6606,N_4399,N_5401);
xnor U6607 (N_6607,N_4910,N_4239);
nor U6608 (N_6608,N_5031,N_4897);
or U6609 (N_6609,N_4243,N_5826);
nor U6610 (N_6610,N_5536,N_4360);
nor U6611 (N_6611,N_5331,N_5015);
nand U6612 (N_6612,N_5040,N_5665);
nor U6613 (N_6613,N_5417,N_5513);
and U6614 (N_6614,N_5178,N_4099);
and U6615 (N_6615,N_5711,N_5418);
or U6616 (N_6616,N_5367,N_5947);
and U6617 (N_6617,N_5573,N_5751);
nor U6618 (N_6618,N_5490,N_4260);
nand U6619 (N_6619,N_4709,N_4907);
nor U6620 (N_6620,N_5901,N_4554);
and U6621 (N_6621,N_4776,N_4158);
nor U6622 (N_6622,N_4899,N_4703);
nor U6623 (N_6623,N_4493,N_5212);
nand U6624 (N_6624,N_5743,N_4505);
and U6625 (N_6625,N_5137,N_4454);
nor U6626 (N_6626,N_5498,N_4983);
xor U6627 (N_6627,N_4032,N_5088);
and U6628 (N_6628,N_4050,N_4530);
nor U6629 (N_6629,N_4896,N_5928);
nand U6630 (N_6630,N_4784,N_4268);
and U6631 (N_6631,N_4161,N_5032);
nor U6632 (N_6632,N_5917,N_4824);
nor U6633 (N_6633,N_4890,N_5464);
nor U6634 (N_6634,N_4654,N_4743);
or U6635 (N_6635,N_4491,N_4124);
or U6636 (N_6636,N_4442,N_4848);
and U6637 (N_6637,N_4585,N_4722);
or U6638 (N_6638,N_4150,N_4282);
nand U6639 (N_6639,N_5507,N_4384);
and U6640 (N_6640,N_5408,N_5381);
and U6641 (N_6641,N_4620,N_4698);
and U6642 (N_6642,N_4397,N_4300);
and U6643 (N_6643,N_5085,N_4640);
nor U6644 (N_6644,N_5764,N_5872);
nor U6645 (N_6645,N_5713,N_5145);
or U6646 (N_6646,N_5593,N_5351);
or U6647 (N_6647,N_5196,N_4877);
xnor U6648 (N_6648,N_4821,N_4773);
and U6649 (N_6649,N_4104,N_5346);
or U6650 (N_6650,N_4561,N_5108);
or U6651 (N_6651,N_4602,N_5170);
or U6652 (N_6652,N_4795,N_5447);
nand U6653 (N_6653,N_4658,N_5194);
xor U6654 (N_6654,N_4741,N_5078);
nor U6655 (N_6655,N_4112,N_4880);
and U6656 (N_6656,N_5833,N_5493);
xor U6657 (N_6657,N_4719,N_4096);
nand U6658 (N_6658,N_4613,N_5465);
nand U6659 (N_6659,N_5727,N_5283);
xor U6660 (N_6660,N_5577,N_5613);
xnor U6661 (N_6661,N_5330,N_4065);
or U6662 (N_6662,N_5794,N_4972);
nand U6663 (N_6663,N_5229,N_4551);
nor U6664 (N_6664,N_4770,N_5936);
and U6665 (N_6665,N_5929,N_4363);
xor U6666 (N_6666,N_4190,N_5129);
nand U6667 (N_6667,N_4747,N_4014);
nand U6668 (N_6668,N_4707,N_5565);
nor U6669 (N_6669,N_5735,N_4735);
or U6670 (N_6670,N_4765,N_5106);
or U6671 (N_6671,N_4245,N_5692);
and U6672 (N_6672,N_4528,N_4685);
or U6673 (N_6673,N_4012,N_4486);
xor U6674 (N_6674,N_4029,N_5914);
and U6675 (N_6675,N_5011,N_5731);
and U6676 (N_6676,N_5337,N_5302);
nor U6677 (N_6677,N_5082,N_5740);
or U6678 (N_6678,N_5130,N_4326);
and U6679 (N_6679,N_4837,N_4424);
or U6680 (N_6680,N_5420,N_5060);
or U6681 (N_6681,N_4314,N_5119);
nand U6682 (N_6682,N_4942,N_4316);
nor U6683 (N_6683,N_5252,N_5462);
xnor U6684 (N_6684,N_5121,N_4228);
nand U6685 (N_6685,N_4531,N_4459);
nor U6686 (N_6686,N_5218,N_4975);
nand U6687 (N_6687,N_5239,N_5159);
nand U6688 (N_6688,N_4307,N_5530);
and U6689 (N_6689,N_4647,N_4330);
nand U6690 (N_6690,N_4339,N_5649);
or U6691 (N_6691,N_4251,N_4606);
or U6692 (N_6692,N_5080,N_5438);
nand U6693 (N_6693,N_4492,N_4055);
or U6694 (N_6694,N_5230,N_5789);
nor U6695 (N_6695,N_4693,N_4332);
and U6696 (N_6696,N_5265,N_4038);
or U6697 (N_6697,N_5793,N_4587);
nor U6698 (N_6698,N_4043,N_4451);
xor U6699 (N_6699,N_5635,N_5073);
or U6700 (N_6700,N_4357,N_5023);
nor U6701 (N_6701,N_4061,N_4148);
or U6702 (N_6702,N_5437,N_5167);
and U6703 (N_6703,N_4652,N_4033);
and U6704 (N_6704,N_4412,N_4376);
nor U6705 (N_6705,N_5154,N_4868);
or U6706 (N_6706,N_5757,N_5352);
nor U6707 (N_6707,N_5044,N_5101);
or U6708 (N_6708,N_5755,N_5997);
nor U6709 (N_6709,N_5334,N_5274);
nor U6710 (N_6710,N_4111,N_5136);
nand U6711 (N_6711,N_5378,N_5869);
and U6712 (N_6712,N_5165,N_4637);
nand U6713 (N_6713,N_5549,N_5639);
xnor U6714 (N_6714,N_4389,N_4347);
nand U6715 (N_6715,N_4702,N_4169);
or U6716 (N_6716,N_4022,N_4334);
nand U6717 (N_6717,N_5132,N_5323);
and U6718 (N_6718,N_4954,N_4733);
and U6719 (N_6719,N_5257,N_4917);
xor U6720 (N_6720,N_5173,N_5227);
or U6721 (N_6721,N_5150,N_5569);
nor U6722 (N_6722,N_5442,N_5858);
or U6723 (N_6723,N_4428,N_5320);
nor U6724 (N_6724,N_5550,N_5326);
nand U6725 (N_6725,N_4390,N_4764);
and U6726 (N_6726,N_4396,N_5992);
xor U6727 (N_6727,N_5172,N_4053);
or U6728 (N_6728,N_5341,N_4958);
and U6729 (N_6729,N_4004,N_4105);
nor U6730 (N_6730,N_5125,N_5332);
nor U6731 (N_6731,N_5823,N_5259);
xnor U6732 (N_6732,N_4751,N_5606);
or U6733 (N_6733,N_4483,N_4725);
and U6734 (N_6734,N_4785,N_5973);
and U6735 (N_6735,N_4962,N_5090);
nand U6736 (N_6736,N_4230,N_4464);
or U6737 (N_6737,N_5585,N_5142);
or U6738 (N_6738,N_4729,N_4350);
nor U6739 (N_6739,N_5541,N_5950);
nand U6740 (N_6740,N_5478,N_5017);
and U6741 (N_6741,N_5072,N_4806);
or U6742 (N_6742,N_4212,N_4690);
nand U6743 (N_6743,N_5738,N_4949);
and U6744 (N_6744,N_5470,N_5604);
nand U6745 (N_6745,N_5800,N_5805);
or U6746 (N_6746,N_5010,N_4080);
or U6747 (N_6747,N_5678,N_5116);
nor U6748 (N_6748,N_4374,N_5582);
nor U6749 (N_6749,N_4232,N_5479);
nor U6750 (N_6750,N_5347,N_5850);
nand U6751 (N_6751,N_5208,N_4064);
and U6752 (N_6752,N_5705,N_4611);
and U6753 (N_6753,N_5375,N_5213);
xnor U6754 (N_6754,N_5097,N_5719);
nand U6755 (N_6755,N_4634,N_5387);
nand U6756 (N_6756,N_4757,N_4663);
nor U6757 (N_6757,N_5623,N_4089);
or U6758 (N_6758,N_4882,N_4817);
nand U6759 (N_6759,N_4964,N_4182);
and U6760 (N_6760,N_4772,N_5603);
or U6761 (N_6761,N_5773,N_5204);
and U6762 (N_6762,N_5294,N_4468);
xnor U6763 (N_6763,N_4689,N_4883);
and U6764 (N_6764,N_5485,N_5042);
nand U6765 (N_6765,N_5193,N_5033);
and U6766 (N_6766,N_4415,N_5637);
nor U6767 (N_6767,N_4841,N_4720);
nand U6768 (N_6768,N_5749,N_4913);
xnor U6769 (N_6769,N_5669,N_4211);
and U6770 (N_6770,N_4372,N_5828);
nand U6771 (N_6771,N_5964,N_5728);
nand U6772 (N_6772,N_4669,N_5215);
nor U6773 (N_6773,N_5312,N_5343);
nand U6774 (N_6774,N_4448,N_4226);
or U6775 (N_6775,N_4113,N_5291);
nand U6776 (N_6776,N_4982,N_4432);
xor U6777 (N_6777,N_4183,N_4632);
nor U6778 (N_6778,N_5679,N_4017);
nor U6779 (N_6779,N_5321,N_4385);
nand U6780 (N_6780,N_5379,N_4661);
nand U6781 (N_6781,N_5907,N_5586);
nand U6782 (N_6782,N_4816,N_4168);
nor U6783 (N_6783,N_4973,N_5931);
xor U6784 (N_6784,N_5179,N_5008);
nor U6785 (N_6785,N_4081,N_4290);
nand U6786 (N_6786,N_5564,N_4320);
and U6787 (N_6787,N_4889,N_4980);
nand U6788 (N_6788,N_4086,N_5591);
nor U6789 (N_6789,N_4387,N_4259);
or U6790 (N_6790,N_4272,N_4116);
or U6791 (N_6791,N_4997,N_4075);
and U6792 (N_6792,N_4026,N_5158);
nor U6793 (N_6793,N_4447,N_5527);
and U6794 (N_6794,N_5972,N_4013);
nor U6795 (N_6795,N_4118,N_4762);
nand U6796 (N_6796,N_4529,N_5878);
or U6797 (N_6797,N_4321,N_4138);
and U6798 (N_6798,N_5243,N_5147);
nor U6799 (N_6799,N_5718,N_5621);
nand U6800 (N_6800,N_4123,N_4351);
or U6801 (N_6801,N_4469,N_4132);
nand U6802 (N_6802,N_4846,N_4264);
nor U6803 (N_6803,N_4343,N_4948);
or U6804 (N_6804,N_4591,N_4609);
nand U6805 (N_6805,N_5282,N_5955);
nor U6806 (N_6806,N_4303,N_5325);
xnor U6807 (N_6807,N_4082,N_5880);
or U6808 (N_6808,N_4386,N_5610);
and U6809 (N_6809,N_5398,N_4818);
xor U6810 (N_6810,N_4750,N_5380);
nand U6811 (N_6811,N_5414,N_5007);
or U6812 (N_6812,N_5818,N_5488);
and U6813 (N_6813,N_5799,N_5519);
or U6814 (N_6814,N_4534,N_4809);
or U6815 (N_6815,N_4645,N_5238);
or U6816 (N_6816,N_5004,N_5104);
nor U6817 (N_6817,N_4998,N_5277);
or U6818 (N_6818,N_5041,N_4863);
and U6819 (N_6819,N_5152,N_5672);
nand U6820 (N_6820,N_4023,N_5922);
nand U6821 (N_6821,N_5533,N_4477);
or U6822 (N_6822,N_5944,N_5959);
xnor U6823 (N_6823,N_4242,N_5228);
or U6824 (N_6824,N_4610,N_4996);
and U6825 (N_6825,N_5553,N_5633);
or U6826 (N_6826,N_4470,N_5275);
nor U6827 (N_6827,N_4365,N_4133);
nor U6828 (N_6828,N_4905,N_5982);
and U6829 (N_6829,N_4324,N_4044);
and U6830 (N_6830,N_5961,N_4224);
nor U6831 (N_6831,N_5440,N_4704);
or U6832 (N_6832,N_5664,N_4302);
or U6833 (N_6833,N_5220,N_5953);
nand U6834 (N_6834,N_4618,N_4730);
or U6835 (N_6835,N_4927,N_5411);
nand U6836 (N_6836,N_5795,N_4317);
nand U6837 (N_6837,N_5151,N_4515);
and U6838 (N_6838,N_5292,N_4823);
and U6839 (N_6839,N_5403,N_5857);
nor U6840 (N_6840,N_4349,N_5701);
xnor U6841 (N_6841,N_5255,N_5921);
or U6842 (N_6842,N_5856,N_4200);
nand U6843 (N_6843,N_4331,N_4830);
nor U6844 (N_6844,N_4419,N_5658);
xnor U6845 (N_6845,N_4323,N_5815);
nor U6846 (N_6846,N_4644,N_5504);
or U6847 (N_6847,N_5018,N_5350);
and U6848 (N_6848,N_4366,N_5064);
nand U6849 (N_6849,N_4458,N_4275);
nand U6850 (N_6850,N_5241,N_4465);
nand U6851 (N_6851,N_5670,N_4495);
xor U6852 (N_6852,N_5918,N_5093);
or U6853 (N_6853,N_4736,N_4382);
or U6854 (N_6854,N_4130,N_5143);
nand U6855 (N_6855,N_5844,N_4077);
or U6856 (N_6856,N_5453,N_5195);
or U6857 (N_6857,N_5286,N_4567);
nand U6858 (N_6858,N_5745,N_4592);
nand U6859 (N_6859,N_5768,N_4746);
nand U6860 (N_6860,N_5181,N_5659);
nand U6861 (N_6861,N_4373,N_5284);
nor U6862 (N_6862,N_5682,N_5599);
nand U6863 (N_6863,N_5118,N_4922);
nor U6864 (N_6864,N_4578,N_4276);
and U6865 (N_6865,N_5413,N_4965);
or U6866 (N_6866,N_5598,N_4443);
and U6867 (N_6867,N_4167,N_4431);
or U6868 (N_6868,N_5355,N_4854);
nor U6869 (N_6869,N_5801,N_5217);
nor U6870 (N_6870,N_4959,N_4115);
nand U6871 (N_6871,N_4460,N_5373);
nor U6872 (N_6872,N_4993,N_5415);
or U6873 (N_6873,N_5395,N_4811);
nor U6874 (N_6874,N_4333,N_4255);
and U6875 (N_6875,N_4027,N_4960);
nand U6876 (N_6876,N_5608,N_5809);
and U6877 (N_6877,N_5141,N_5272);
or U6878 (N_6878,N_5967,N_5570);
nand U6879 (N_6879,N_5594,N_4872);
and U6880 (N_6880,N_5765,N_5135);
or U6881 (N_6881,N_5898,N_4377);
nor U6882 (N_6882,N_5845,N_5348);
or U6883 (N_6883,N_5232,N_4015);
and U6884 (N_6884,N_5405,N_5030);
or U6885 (N_6885,N_5336,N_5875);
and U6886 (N_6886,N_4070,N_4710);
nand U6887 (N_6887,N_5458,N_4201);
nand U6888 (N_6888,N_5454,N_4185);
xnor U6889 (N_6889,N_5211,N_5883);
nor U6890 (N_6890,N_4926,N_5537);
nor U6891 (N_6891,N_4678,N_5113);
nor U6892 (N_6892,N_5948,N_4359);
nor U6893 (N_6893,N_4237,N_4461);
nand U6894 (N_6894,N_5899,N_4210);
and U6895 (N_6895,N_4156,N_5702);
nand U6896 (N_6896,N_5868,N_4482);
or U6897 (N_6897,N_5262,N_5266);
and U6898 (N_6898,N_5785,N_5566);
or U6899 (N_6899,N_4103,N_5890);
or U6900 (N_6900,N_4162,N_4984);
or U6901 (N_6901,N_4001,N_5739);
or U6902 (N_6902,N_4305,N_4522);
nand U6903 (N_6903,N_4449,N_4577);
and U6904 (N_6904,N_5988,N_4097);
nor U6905 (N_6905,N_5480,N_4646);
xnor U6906 (N_6906,N_4322,N_5560);
or U6907 (N_6907,N_4781,N_5767);
nor U6908 (N_6908,N_4582,N_4151);
xnor U6909 (N_6909,N_4532,N_4209);
and U6910 (N_6910,N_4021,N_5431);
and U6911 (N_6911,N_4930,N_5572);
nand U6912 (N_6912,N_4886,N_5186);
nor U6913 (N_6913,N_4976,N_5176);
nand U6914 (N_6914,N_4536,N_5075);
nand U6915 (N_6915,N_5726,N_4584);
nor U6916 (N_6916,N_4402,N_4696);
nand U6917 (N_6917,N_4892,N_4871);
or U6918 (N_6918,N_5406,N_5083);
nor U6919 (N_6919,N_4207,N_4968);
and U6920 (N_6920,N_4278,N_4277);
nand U6921 (N_6921,N_4595,N_5622);
or U6922 (N_6922,N_5443,N_5941);
nor U6923 (N_6923,N_4986,N_5127);
and U6924 (N_6924,N_4701,N_5456);
xnor U6925 (N_6925,N_4656,N_4862);
and U6926 (N_6926,N_4858,N_4280);
nand U6927 (N_6927,N_5696,N_4556);
nand U6928 (N_6928,N_5900,N_5357);
nand U6929 (N_6929,N_5902,N_4981);
or U6930 (N_6930,N_4797,N_4808);
and U6931 (N_6931,N_5481,N_4876);
nand U6932 (N_6932,N_4590,N_4392);
nor U6933 (N_6933,N_4335,N_5134);
or U6934 (N_6934,N_5177,N_4087);
nor U6935 (N_6935,N_4444,N_5596);
nor U6936 (N_6936,N_5963,N_4560);
and U6937 (N_6937,N_4576,N_5459);
or U6938 (N_6938,N_5059,N_5624);
nand U6939 (N_6939,N_5896,N_5787);
nor U6940 (N_6940,N_4106,N_5511);
or U6941 (N_6941,N_5671,N_4198);
or U6942 (N_6942,N_4244,N_5796);
nor U6943 (N_6943,N_4974,N_5028);
nand U6944 (N_6944,N_5363,N_4599);
and U6945 (N_6945,N_5791,N_5838);
nand U6946 (N_6946,N_5960,N_5371);
nor U6947 (N_6947,N_5546,N_5986);
or U6948 (N_6948,N_4395,N_4034);
nor U6949 (N_6949,N_4028,N_4617);
xnor U6950 (N_6950,N_5068,N_5264);
and U6951 (N_6951,N_4457,N_4046);
nor U6952 (N_6952,N_4956,N_5689);
nand U6953 (N_6953,N_4427,N_4869);
and U6954 (N_6954,N_4218,N_5946);
xnor U6955 (N_6955,N_4042,N_4538);
and U6956 (N_6956,N_4304,N_5365);
and U6957 (N_6957,N_5188,N_5133);
or U6958 (N_6958,N_5811,N_4527);
or U6959 (N_6959,N_5155,N_5316);
nand U6960 (N_6960,N_5699,N_5149);
nor U6961 (N_6961,N_5729,N_4516);
and U6962 (N_6962,N_5601,N_5535);
or U6963 (N_6963,N_4328,N_5100);
or U6964 (N_6964,N_5882,N_4855);
or U6965 (N_6965,N_4507,N_5285);
or U6966 (N_6966,N_4186,N_5328);
nor U6967 (N_6967,N_5744,N_4125);
and U6968 (N_6968,N_5198,N_5956);
nand U6969 (N_6969,N_5884,N_4805);
nand U6970 (N_6970,N_5747,N_4298);
or U6971 (N_6971,N_4699,N_4598);
xnor U6972 (N_6972,N_5109,N_5926);
or U6973 (N_6973,N_5770,N_4822);
xor U6974 (N_6974,N_4827,N_4523);
and U6975 (N_6975,N_4653,N_4299);
or U6976 (N_6976,N_4562,N_4923);
nand U6977 (N_6977,N_4406,N_5851);
nor U6978 (N_6978,N_5746,N_4490);
nor U6979 (N_6979,N_5839,N_4135);
and U6980 (N_6980,N_5486,N_5562);
or U6981 (N_6981,N_4787,N_4668);
nand U6982 (N_6982,N_5543,N_4630);
nand U6983 (N_6983,N_5446,N_4286);
nor U6984 (N_6984,N_4092,N_4859);
and U6985 (N_6985,N_5301,N_5867);
xor U6986 (N_6986,N_4909,N_4353);
nand U6987 (N_6987,N_4434,N_5027);
and U6988 (N_6988,N_4094,N_5055);
nand U6989 (N_6989,N_5863,N_4870);
nand U6990 (N_6990,N_4020,N_4539);
nand U6991 (N_6991,N_5933,N_4437);
nor U6992 (N_6992,N_4727,N_5968);
nor U6993 (N_6993,N_5715,N_4234);
or U6994 (N_6994,N_4836,N_4541);
nor U6995 (N_6995,N_4355,N_5939);
nor U6996 (N_6996,N_4812,N_5290);
nor U6997 (N_6997,N_4122,N_5741);
and U6998 (N_6998,N_4281,N_4579);
and U6999 (N_6999,N_5829,N_4692);
or U7000 (N_7000,N_4648,N_5360);
or U7001 (N_7001,N_4058,N_4257);
nor U7002 (N_7002,N_5530,N_4292);
or U7003 (N_7003,N_4891,N_4164);
and U7004 (N_7004,N_5141,N_5999);
nand U7005 (N_7005,N_4060,N_4096);
nor U7006 (N_7006,N_5110,N_4199);
or U7007 (N_7007,N_5434,N_4290);
nand U7008 (N_7008,N_4736,N_5747);
nand U7009 (N_7009,N_4981,N_5819);
nor U7010 (N_7010,N_5887,N_5815);
nand U7011 (N_7011,N_5342,N_5765);
and U7012 (N_7012,N_5487,N_5858);
nor U7013 (N_7013,N_5114,N_4921);
or U7014 (N_7014,N_5582,N_4375);
or U7015 (N_7015,N_5750,N_5571);
or U7016 (N_7016,N_5162,N_5556);
and U7017 (N_7017,N_5472,N_5321);
xor U7018 (N_7018,N_5536,N_5896);
xnor U7019 (N_7019,N_5733,N_5672);
nand U7020 (N_7020,N_4766,N_4362);
or U7021 (N_7021,N_4240,N_4173);
and U7022 (N_7022,N_5260,N_4046);
nor U7023 (N_7023,N_5511,N_5128);
and U7024 (N_7024,N_4839,N_5931);
nand U7025 (N_7025,N_5522,N_4497);
nor U7026 (N_7026,N_4212,N_5086);
or U7027 (N_7027,N_5659,N_4952);
xnor U7028 (N_7028,N_5035,N_4647);
and U7029 (N_7029,N_4872,N_5340);
nand U7030 (N_7030,N_4290,N_5560);
and U7031 (N_7031,N_5017,N_5043);
nand U7032 (N_7032,N_5817,N_5327);
nor U7033 (N_7033,N_4035,N_4765);
nand U7034 (N_7034,N_4177,N_4210);
nand U7035 (N_7035,N_5062,N_5005);
xor U7036 (N_7036,N_5513,N_4686);
or U7037 (N_7037,N_5131,N_4172);
nor U7038 (N_7038,N_5111,N_4751);
nand U7039 (N_7039,N_5246,N_5440);
or U7040 (N_7040,N_5752,N_5320);
or U7041 (N_7041,N_4042,N_5616);
and U7042 (N_7042,N_5656,N_5790);
nand U7043 (N_7043,N_5025,N_5299);
nor U7044 (N_7044,N_5931,N_5525);
and U7045 (N_7045,N_4198,N_4296);
nor U7046 (N_7046,N_4635,N_4990);
xor U7047 (N_7047,N_4926,N_4864);
or U7048 (N_7048,N_5874,N_5607);
nand U7049 (N_7049,N_4214,N_5280);
and U7050 (N_7050,N_4131,N_4781);
nor U7051 (N_7051,N_4757,N_4382);
nand U7052 (N_7052,N_4395,N_5062);
nor U7053 (N_7053,N_4585,N_4125);
and U7054 (N_7054,N_4055,N_5319);
or U7055 (N_7055,N_5225,N_5906);
or U7056 (N_7056,N_5819,N_4319);
nand U7057 (N_7057,N_5832,N_4948);
xnor U7058 (N_7058,N_4974,N_5569);
nand U7059 (N_7059,N_4068,N_4037);
xnor U7060 (N_7060,N_4339,N_5495);
nand U7061 (N_7061,N_5750,N_4121);
nand U7062 (N_7062,N_4690,N_5459);
nor U7063 (N_7063,N_4535,N_4386);
nand U7064 (N_7064,N_4434,N_4666);
and U7065 (N_7065,N_5476,N_4516);
and U7066 (N_7066,N_4172,N_5303);
nor U7067 (N_7067,N_4635,N_4237);
nand U7068 (N_7068,N_5373,N_5250);
nand U7069 (N_7069,N_5851,N_4101);
nand U7070 (N_7070,N_4823,N_4425);
and U7071 (N_7071,N_4307,N_5359);
or U7072 (N_7072,N_5485,N_4908);
nand U7073 (N_7073,N_5891,N_4457);
and U7074 (N_7074,N_5201,N_5236);
or U7075 (N_7075,N_5393,N_5423);
xor U7076 (N_7076,N_4328,N_4849);
xnor U7077 (N_7077,N_4351,N_4634);
or U7078 (N_7078,N_5328,N_5184);
and U7079 (N_7079,N_4206,N_5651);
or U7080 (N_7080,N_4402,N_5329);
and U7081 (N_7081,N_4378,N_4224);
nor U7082 (N_7082,N_4863,N_4939);
or U7083 (N_7083,N_4282,N_4788);
nand U7084 (N_7084,N_5208,N_4005);
or U7085 (N_7085,N_4524,N_4433);
and U7086 (N_7086,N_5079,N_4400);
or U7087 (N_7087,N_5186,N_5955);
and U7088 (N_7088,N_5714,N_4126);
and U7089 (N_7089,N_5840,N_4293);
and U7090 (N_7090,N_5472,N_5294);
and U7091 (N_7091,N_5126,N_5718);
or U7092 (N_7092,N_4690,N_4456);
or U7093 (N_7093,N_5061,N_4243);
and U7094 (N_7094,N_4043,N_4199);
and U7095 (N_7095,N_4945,N_4629);
and U7096 (N_7096,N_5483,N_5230);
nand U7097 (N_7097,N_5651,N_4141);
xnor U7098 (N_7098,N_5366,N_5744);
or U7099 (N_7099,N_4471,N_4735);
nor U7100 (N_7100,N_5004,N_4862);
and U7101 (N_7101,N_4669,N_5845);
xor U7102 (N_7102,N_5141,N_5012);
nor U7103 (N_7103,N_4711,N_4653);
or U7104 (N_7104,N_4548,N_5463);
or U7105 (N_7105,N_5227,N_4283);
nand U7106 (N_7106,N_4405,N_4489);
nand U7107 (N_7107,N_4815,N_5179);
or U7108 (N_7108,N_4364,N_5525);
xor U7109 (N_7109,N_4583,N_4011);
nand U7110 (N_7110,N_5403,N_4283);
and U7111 (N_7111,N_4929,N_4387);
nor U7112 (N_7112,N_5200,N_4341);
nand U7113 (N_7113,N_4565,N_4095);
nand U7114 (N_7114,N_4650,N_5626);
and U7115 (N_7115,N_5541,N_4486);
nand U7116 (N_7116,N_4917,N_5621);
and U7117 (N_7117,N_5797,N_5615);
nand U7118 (N_7118,N_5969,N_5725);
xnor U7119 (N_7119,N_5016,N_4977);
nor U7120 (N_7120,N_5669,N_5511);
and U7121 (N_7121,N_4682,N_5614);
or U7122 (N_7122,N_5145,N_5013);
nand U7123 (N_7123,N_5516,N_4801);
or U7124 (N_7124,N_5101,N_4669);
nand U7125 (N_7125,N_4389,N_4144);
xor U7126 (N_7126,N_5834,N_5258);
nor U7127 (N_7127,N_4855,N_4621);
and U7128 (N_7128,N_5658,N_5805);
nand U7129 (N_7129,N_5799,N_4784);
nand U7130 (N_7130,N_4374,N_5779);
nand U7131 (N_7131,N_5049,N_5220);
nor U7132 (N_7132,N_5145,N_5359);
nor U7133 (N_7133,N_4196,N_5128);
nor U7134 (N_7134,N_5239,N_5739);
xor U7135 (N_7135,N_5222,N_4425);
nand U7136 (N_7136,N_5298,N_4140);
or U7137 (N_7137,N_4103,N_5086);
nor U7138 (N_7138,N_4965,N_5415);
xnor U7139 (N_7139,N_4223,N_4874);
nor U7140 (N_7140,N_4453,N_4774);
nand U7141 (N_7141,N_4921,N_5668);
nand U7142 (N_7142,N_5960,N_5805);
or U7143 (N_7143,N_5491,N_5932);
nor U7144 (N_7144,N_5089,N_4074);
nor U7145 (N_7145,N_4849,N_5965);
and U7146 (N_7146,N_4661,N_4048);
or U7147 (N_7147,N_5116,N_5227);
and U7148 (N_7148,N_4209,N_4013);
nand U7149 (N_7149,N_4717,N_5793);
nand U7150 (N_7150,N_4928,N_5192);
or U7151 (N_7151,N_5892,N_4950);
or U7152 (N_7152,N_5965,N_5868);
nor U7153 (N_7153,N_4485,N_5866);
xnor U7154 (N_7154,N_5989,N_4676);
or U7155 (N_7155,N_5812,N_4661);
nor U7156 (N_7156,N_5046,N_4407);
or U7157 (N_7157,N_4959,N_4308);
and U7158 (N_7158,N_5560,N_4310);
xor U7159 (N_7159,N_4674,N_5589);
nor U7160 (N_7160,N_5973,N_4364);
and U7161 (N_7161,N_5232,N_4274);
nand U7162 (N_7162,N_4423,N_5501);
and U7163 (N_7163,N_4627,N_5048);
nand U7164 (N_7164,N_5736,N_5599);
nor U7165 (N_7165,N_5424,N_4927);
xor U7166 (N_7166,N_5145,N_4938);
and U7167 (N_7167,N_4056,N_5542);
nor U7168 (N_7168,N_4694,N_5946);
or U7169 (N_7169,N_4869,N_5561);
or U7170 (N_7170,N_4217,N_4591);
and U7171 (N_7171,N_5487,N_4082);
and U7172 (N_7172,N_4551,N_5046);
nor U7173 (N_7173,N_5307,N_5012);
and U7174 (N_7174,N_4040,N_5764);
or U7175 (N_7175,N_4885,N_4987);
and U7176 (N_7176,N_4118,N_5427);
xor U7177 (N_7177,N_5903,N_5361);
and U7178 (N_7178,N_5908,N_4906);
and U7179 (N_7179,N_4948,N_4137);
nand U7180 (N_7180,N_4159,N_4748);
or U7181 (N_7181,N_4778,N_4658);
xnor U7182 (N_7182,N_4506,N_5119);
nand U7183 (N_7183,N_4523,N_4124);
and U7184 (N_7184,N_4301,N_4450);
and U7185 (N_7185,N_5715,N_4633);
nand U7186 (N_7186,N_5361,N_4945);
and U7187 (N_7187,N_5942,N_5172);
or U7188 (N_7188,N_5080,N_5778);
xor U7189 (N_7189,N_4401,N_4888);
nor U7190 (N_7190,N_5450,N_4342);
or U7191 (N_7191,N_5762,N_4061);
and U7192 (N_7192,N_5432,N_5045);
nand U7193 (N_7193,N_5385,N_4772);
or U7194 (N_7194,N_5950,N_5895);
nand U7195 (N_7195,N_4530,N_4882);
or U7196 (N_7196,N_5154,N_4982);
xnor U7197 (N_7197,N_5388,N_5447);
nor U7198 (N_7198,N_5423,N_4740);
and U7199 (N_7199,N_5798,N_5400);
or U7200 (N_7200,N_5386,N_4096);
or U7201 (N_7201,N_5532,N_5633);
and U7202 (N_7202,N_4619,N_4979);
nand U7203 (N_7203,N_4107,N_4240);
or U7204 (N_7204,N_5077,N_5090);
nor U7205 (N_7205,N_4238,N_4499);
nor U7206 (N_7206,N_5486,N_5069);
nor U7207 (N_7207,N_4984,N_4104);
or U7208 (N_7208,N_4545,N_5022);
nand U7209 (N_7209,N_5157,N_4714);
nor U7210 (N_7210,N_5606,N_4701);
or U7211 (N_7211,N_4125,N_4034);
xnor U7212 (N_7212,N_5678,N_4651);
nand U7213 (N_7213,N_5122,N_4989);
or U7214 (N_7214,N_5864,N_5220);
nor U7215 (N_7215,N_4470,N_4769);
or U7216 (N_7216,N_4096,N_4243);
and U7217 (N_7217,N_5466,N_5191);
nor U7218 (N_7218,N_5574,N_4274);
nand U7219 (N_7219,N_5253,N_4917);
and U7220 (N_7220,N_4329,N_4793);
xor U7221 (N_7221,N_5336,N_4911);
or U7222 (N_7222,N_5938,N_5998);
nor U7223 (N_7223,N_4188,N_5370);
nor U7224 (N_7224,N_4059,N_5479);
or U7225 (N_7225,N_5219,N_4247);
nand U7226 (N_7226,N_5325,N_5645);
nor U7227 (N_7227,N_4277,N_5310);
nor U7228 (N_7228,N_4825,N_5748);
or U7229 (N_7229,N_4080,N_5720);
and U7230 (N_7230,N_5482,N_4675);
and U7231 (N_7231,N_4472,N_4236);
xor U7232 (N_7232,N_5965,N_5283);
and U7233 (N_7233,N_5558,N_4192);
and U7234 (N_7234,N_4041,N_5832);
nand U7235 (N_7235,N_5908,N_5499);
nor U7236 (N_7236,N_5027,N_5784);
xor U7237 (N_7237,N_5156,N_4443);
and U7238 (N_7238,N_4431,N_5013);
nor U7239 (N_7239,N_4781,N_5034);
nand U7240 (N_7240,N_4319,N_5828);
nand U7241 (N_7241,N_4271,N_4770);
or U7242 (N_7242,N_4028,N_4591);
nor U7243 (N_7243,N_4943,N_5393);
nand U7244 (N_7244,N_4607,N_4749);
or U7245 (N_7245,N_5206,N_5865);
xor U7246 (N_7246,N_4581,N_5083);
nor U7247 (N_7247,N_5377,N_4075);
nor U7248 (N_7248,N_5358,N_4479);
or U7249 (N_7249,N_5357,N_5904);
xnor U7250 (N_7250,N_4597,N_5089);
nor U7251 (N_7251,N_4203,N_4878);
nand U7252 (N_7252,N_5424,N_5990);
nand U7253 (N_7253,N_5977,N_5280);
nand U7254 (N_7254,N_5820,N_5363);
nand U7255 (N_7255,N_4506,N_5835);
nand U7256 (N_7256,N_4937,N_4181);
nor U7257 (N_7257,N_5903,N_5933);
nand U7258 (N_7258,N_5102,N_5590);
nor U7259 (N_7259,N_5011,N_5631);
or U7260 (N_7260,N_5109,N_4571);
nor U7261 (N_7261,N_4449,N_4890);
xnor U7262 (N_7262,N_5828,N_4913);
nor U7263 (N_7263,N_5711,N_4153);
or U7264 (N_7264,N_4936,N_4060);
or U7265 (N_7265,N_4769,N_5717);
nand U7266 (N_7266,N_4952,N_4956);
or U7267 (N_7267,N_4192,N_5572);
nand U7268 (N_7268,N_5314,N_5961);
nand U7269 (N_7269,N_4232,N_4301);
xor U7270 (N_7270,N_5468,N_4779);
or U7271 (N_7271,N_5996,N_5299);
or U7272 (N_7272,N_4595,N_4247);
or U7273 (N_7273,N_4920,N_4893);
nand U7274 (N_7274,N_4592,N_5620);
or U7275 (N_7275,N_5671,N_5313);
nand U7276 (N_7276,N_4622,N_5749);
and U7277 (N_7277,N_4497,N_4663);
nand U7278 (N_7278,N_5428,N_4106);
xor U7279 (N_7279,N_4318,N_4908);
nand U7280 (N_7280,N_4485,N_4833);
and U7281 (N_7281,N_4204,N_4251);
or U7282 (N_7282,N_4765,N_5402);
or U7283 (N_7283,N_5441,N_5357);
or U7284 (N_7284,N_5996,N_4375);
or U7285 (N_7285,N_5342,N_4266);
nor U7286 (N_7286,N_5971,N_4432);
nand U7287 (N_7287,N_4828,N_5288);
nor U7288 (N_7288,N_4411,N_4280);
and U7289 (N_7289,N_5229,N_5015);
and U7290 (N_7290,N_5743,N_5597);
xor U7291 (N_7291,N_4317,N_5914);
nor U7292 (N_7292,N_4542,N_5266);
or U7293 (N_7293,N_5818,N_5343);
nor U7294 (N_7294,N_5878,N_5251);
nand U7295 (N_7295,N_5623,N_4436);
and U7296 (N_7296,N_5258,N_4690);
or U7297 (N_7297,N_5973,N_4707);
nor U7298 (N_7298,N_4803,N_4174);
nand U7299 (N_7299,N_5285,N_5282);
or U7300 (N_7300,N_4639,N_5399);
nand U7301 (N_7301,N_4799,N_4759);
nand U7302 (N_7302,N_5938,N_5907);
or U7303 (N_7303,N_5702,N_4624);
nor U7304 (N_7304,N_5577,N_5473);
or U7305 (N_7305,N_4404,N_4491);
xor U7306 (N_7306,N_4942,N_4234);
and U7307 (N_7307,N_5125,N_5221);
or U7308 (N_7308,N_5635,N_4461);
nand U7309 (N_7309,N_4751,N_4535);
and U7310 (N_7310,N_5085,N_4907);
or U7311 (N_7311,N_4291,N_5369);
nand U7312 (N_7312,N_4611,N_4967);
or U7313 (N_7313,N_4867,N_4448);
nand U7314 (N_7314,N_5677,N_5332);
nor U7315 (N_7315,N_5423,N_5651);
or U7316 (N_7316,N_4351,N_4329);
nand U7317 (N_7317,N_4979,N_5398);
and U7318 (N_7318,N_4098,N_5128);
nor U7319 (N_7319,N_5477,N_5871);
nor U7320 (N_7320,N_4925,N_4231);
nand U7321 (N_7321,N_5480,N_4543);
or U7322 (N_7322,N_4538,N_5484);
or U7323 (N_7323,N_4497,N_4025);
nand U7324 (N_7324,N_5532,N_4426);
xor U7325 (N_7325,N_4915,N_4503);
nand U7326 (N_7326,N_5007,N_4857);
nand U7327 (N_7327,N_5266,N_5209);
and U7328 (N_7328,N_5597,N_4830);
or U7329 (N_7329,N_5745,N_5545);
nor U7330 (N_7330,N_4028,N_4250);
xor U7331 (N_7331,N_5552,N_5825);
nand U7332 (N_7332,N_4621,N_4050);
xor U7333 (N_7333,N_4160,N_5539);
or U7334 (N_7334,N_5292,N_4158);
or U7335 (N_7335,N_5277,N_4434);
nand U7336 (N_7336,N_4263,N_5853);
nor U7337 (N_7337,N_5450,N_5184);
or U7338 (N_7338,N_4047,N_5451);
nor U7339 (N_7339,N_4478,N_4945);
xnor U7340 (N_7340,N_4137,N_4464);
nor U7341 (N_7341,N_4087,N_5822);
nor U7342 (N_7342,N_4562,N_4591);
and U7343 (N_7343,N_5670,N_4138);
or U7344 (N_7344,N_5154,N_5729);
nor U7345 (N_7345,N_5590,N_4654);
nor U7346 (N_7346,N_4893,N_5291);
nor U7347 (N_7347,N_4440,N_5840);
and U7348 (N_7348,N_4050,N_4597);
nand U7349 (N_7349,N_5374,N_4753);
nor U7350 (N_7350,N_4177,N_5990);
and U7351 (N_7351,N_4402,N_5097);
or U7352 (N_7352,N_4299,N_4759);
or U7353 (N_7353,N_4397,N_4591);
and U7354 (N_7354,N_4644,N_5281);
nor U7355 (N_7355,N_4811,N_5539);
and U7356 (N_7356,N_5117,N_4053);
nand U7357 (N_7357,N_4128,N_4372);
nor U7358 (N_7358,N_5076,N_5712);
or U7359 (N_7359,N_5492,N_4571);
nand U7360 (N_7360,N_5371,N_4685);
nor U7361 (N_7361,N_4370,N_4502);
nand U7362 (N_7362,N_4502,N_4466);
nand U7363 (N_7363,N_4476,N_4584);
nor U7364 (N_7364,N_5667,N_5624);
or U7365 (N_7365,N_5691,N_4277);
or U7366 (N_7366,N_5780,N_5244);
and U7367 (N_7367,N_4856,N_5759);
xnor U7368 (N_7368,N_5173,N_5995);
or U7369 (N_7369,N_5718,N_4882);
nor U7370 (N_7370,N_5497,N_5969);
or U7371 (N_7371,N_4160,N_5070);
and U7372 (N_7372,N_5500,N_5656);
nand U7373 (N_7373,N_4000,N_4607);
nor U7374 (N_7374,N_5331,N_5958);
and U7375 (N_7375,N_5581,N_4314);
nand U7376 (N_7376,N_5793,N_4916);
and U7377 (N_7377,N_5934,N_5379);
xnor U7378 (N_7378,N_5829,N_4435);
nand U7379 (N_7379,N_4541,N_4781);
nand U7380 (N_7380,N_5813,N_4927);
nor U7381 (N_7381,N_5056,N_5737);
and U7382 (N_7382,N_5343,N_4858);
nand U7383 (N_7383,N_5384,N_4790);
nor U7384 (N_7384,N_4201,N_4874);
nand U7385 (N_7385,N_4269,N_5848);
and U7386 (N_7386,N_5205,N_5902);
nor U7387 (N_7387,N_4538,N_4509);
or U7388 (N_7388,N_4594,N_5285);
nand U7389 (N_7389,N_4891,N_5083);
and U7390 (N_7390,N_4691,N_5377);
or U7391 (N_7391,N_4918,N_4555);
nor U7392 (N_7392,N_4128,N_5688);
xnor U7393 (N_7393,N_5855,N_4987);
xnor U7394 (N_7394,N_5420,N_4502);
or U7395 (N_7395,N_4760,N_5780);
nand U7396 (N_7396,N_5393,N_5549);
nor U7397 (N_7397,N_5150,N_5824);
nor U7398 (N_7398,N_5617,N_5855);
nor U7399 (N_7399,N_4192,N_4514);
or U7400 (N_7400,N_4174,N_4136);
and U7401 (N_7401,N_4378,N_5436);
nor U7402 (N_7402,N_5798,N_4760);
and U7403 (N_7403,N_5500,N_5937);
or U7404 (N_7404,N_5223,N_4285);
and U7405 (N_7405,N_4955,N_4081);
and U7406 (N_7406,N_4329,N_4188);
nor U7407 (N_7407,N_5127,N_5075);
nand U7408 (N_7408,N_5301,N_4299);
nand U7409 (N_7409,N_5052,N_4396);
or U7410 (N_7410,N_5216,N_4039);
or U7411 (N_7411,N_5963,N_4450);
nand U7412 (N_7412,N_5334,N_4198);
or U7413 (N_7413,N_5299,N_4594);
nand U7414 (N_7414,N_4686,N_4248);
nand U7415 (N_7415,N_5026,N_5272);
xnor U7416 (N_7416,N_5625,N_4785);
and U7417 (N_7417,N_4491,N_5974);
nand U7418 (N_7418,N_5843,N_4017);
and U7419 (N_7419,N_4558,N_5528);
or U7420 (N_7420,N_5147,N_5895);
or U7421 (N_7421,N_4886,N_5714);
xnor U7422 (N_7422,N_5353,N_4823);
nor U7423 (N_7423,N_4582,N_4382);
nor U7424 (N_7424,N_4473,N_5183);
or U7425 (N_7425,N_4957,N_4325);
nor U7426 (N_7426,N_5203,N_4542);
xnor U7427 (N_7427,N_5783,N_5818);
or U7428 (N_7428,N_4538,N_5873);
nor U7429 (N_7429,N_5468,N_5923);
xnor U7430 (N_7430,N_5223,N_5800);
or U7431 (N_7431,N_4436,N_5569);
nor U7432 (N_7432,N_5773,N_5043);
and U7433 (N_7433,N_4513,N_5692);
nand U7434 (N_7434,N_4623,N_5967);
nand U7435 (N_7435,N_4197,N_5650);
and U7436 (N_7436,N_5499,N_5646);
nand U7437 (N_7437,N_4517,N_5742);
nor U7438 (N_7438,N_5420,N_4662);
xor U7439 (N_7439,N_5414,N_5839);
and U7440 (N_7440,N_5873,N_4967);
and U7441 (N_7441,N_4291,N_5509);
and U7442 (N_7442,N_4835,N_5429);
and U7443 (N_7443,N_4262,N_4903);
nand U7444 (N_7444,N_5170,N_5542);
nor U7445 (N_7445,N_5983,N_4247);
or U7446 (N_7446,N_5413,N_5850);
and U7447 (N_7447,N_4024,N_5639);
nand U7448 (N_7448,N_5376,N_4856);
or U7449 (N_7449,N_4243,N_4489);
nand U7450 (N_7450,N_4623,N_5104);
or U7451 (N_7451,N_5484,N_5873);
or U7452 (N_7452,N_4314,N_5701);
nand U7453 (N_7453,N_5938,N_4022);
nand U7454 (N_7454,N_5916,N_4253);
xnor U7455 (N_7455,N_4065,N_5905);
or U7456 (N_7456,N_4556,N_4008);
and U7457 (N_7457,N_4680,N_5540);
xnor U7458 (N_7458,N_5689,N_4834);
nor U7459 (N_7459,N_4855,N_4305);
nand U7460 (N_7460,N_4747,N_4242);
xnor U7461 (N_7461,N_5021,N_4845);
nand U7462 (N_7462,N_5777,N_4516);
xnor U7463 (N_7463,N_4610,N_5441);
and U7464 (N_7464,N_4252,N_4897);
or U7465 (N_7465,N_4695,N_5942);
and U7466 (N_7466,N_5710,N_4329);
xnor U7467 (N_7467,N_4183,N_4598);
or U7468 (N_7468,N_5535,N_4567);
xnor U7469 (N_7469,N_4323,N_4793);
xnor U7470 (N_7470,N_4372,N_4094);
xnor U7471 (N_7471,N_4779,N_5043);
nand U7472 (N_7472,N_4394,N_5205);
nor U7473 (N_7473,N_4499,N_4764);
or U7474 (N_7474,N_5069,N_5404);
nor U7475 (N_7475,N_5649,N_5659);
and U7476 (N_7476,N_4549,N_4884);
nor U7477 (N_7477,N_5030,N_4474);
nand U7478 (N_7478,N_4196,N_4752);
or U7479 (N_7479,N_5954,N_4417);
or U7480 (N_7480,N_4589,N_4081);
or U7481 (N_7481,N_4186,N_4144);
nor U7482 (N_7482,N_5507,N_4561);
or U7483 (N_7483,N_5443,N_4448);
nand U7484 (N_7484,N_5452,N_5884);
nand U7485 (N_7485,N_5357,N_4717);
nand U7486 (N_7486,N_5299,N_5997);
nand U7487 (N_7487,N_4351,N_4218);
or U7488 (N_7488,N_5435,N_5614);
nand U7489 (N_7489,N_4918,N_5109);
nand U7490 (N_7490,N_5382,N_5284);
xor U7491 (N_7491,N_5593,N_5283);
and U7492 (N_7492,N_4700,N_5585);
and U7493 (N_7493,N_4095,N_5622);
nor U7494 (N_7494,N_4808,N_5175);
or U7495 (N_7495,N_4518,N_4273);
or U7496 (N_7496,N_4833,N_5162);
nor U7497 (N_7497,N_5731,N_5412);
and U7498 (N_7498,N_4751,N_5021);
and U7499 (N_7499,N_5671,N_5467);
or U7500 (N_7500,N_4215,N_4089);
xnor U7501 (N_7501,N_4608,N_5285);
and U7502 (N_7502,N_5769,N_5532);
nand U7503 (N_7503,N_5262,N_5863);
nor U7504 (N_7504,N_5828,N_4442);
nand U7505 (N_7505,N_4902,N_5209);
nor U7506 (N_7506,N_4682,N_5411);
xnor U7507 (N_7507,N_4518,N_4384);
nor U7508 (N_7508,N_4823,N_5145);
nor U7509 (N_7509,N_4829,N_4416);
xnor U7510 (N_7510,N_5934,N_5941);
xnor U7511 (N_7511,N_4715,N_5943);
nor U7512 (N_7512,N_4189,N_4844);
nand U7513 (N_7513,N_5583,N_4417);
and U7514 (N_7514,N_4360,N_5773);
xnor U7515 (N_7515,N_4209,N_4032);
nor U7516 (N_7516,N_5044,N_4799);
nor U7517 (N_7517,N_4939,N_4172);
and U7518 (N_7518,N_5114,N_5019);
nand U7519 (N_7519,N_5625,N_4987);
or U7520 (N_7520,N_5790,N_4945);
or U7521 (N_7521,N_4327,N_4660);
and U7522 (N_7522,N_4613,N_5325);
nor U7523 (N_7523,N_4706,N_5961);
and U7524 (N_7524,N_4824,N_5639);
nor U7525 (N_7525,N_4624,N_4689);
nor U7526 (N_7526,N_4471,N_4912);
nand U7527 (N_7527,N_5009,N_4991);
and U7528 (N_7528,N_4319,N_4960);
nand U7529 (N_7529,N_5892,N_5639);
or U7530 (N_7530,N_4736,N_5315);
or U7531 (N_7531,N_4616,N_5662);
and U7532 (N_7532,N_5371,N_4642);
nor U7533 (N_7533,N_5850,N_5394);
nand U7534 (N_7534,N_4703,N_5857);
or U7535 (N_7535,N_4471,N_4176);
and U7536 (N_7536,N_4265,N_4465);
and U7537 (N_7537,N_4900,N_5536);
and U7538 (N_7538,N_4502,N_4374);
and U7539 (N_7539,N_5175,N_4472);
or U7540 (N_7540,N_5738,N_4959);
nor U7541 (N_7541,N_4997,N_5706);
nand U7542 (N_7542,N_4453,N_4091);
nor U7543 (N_7543,N_5415,N_5075);
and U7544 (N_7544,N_4688,N_4619);
nand U7545 (N_7545,N_5180,N_5417);
nand U7546 (N_7546,N_5987,N_5707);
or U7547 (N_7547,N_5518,N_5754);
nor U7548 (N_7548,N_4839,N_4592);
nand U7549 (N_7549,N_4184,N_5893);
or U7550 (N_7550,N_5622,N_5983);
nor U7551 (N_7551,N_5347,N_5903);
nor U7552 (N_7552,N_4305,N_4934);
and U7553 (N_7553,N_4235,N_5261);
nor U7554 (N_7554,N_4224,N_5672);
nand U7555 (N_7555,N_5951,N_4728);
nor U7556 (N_7556,N_5280,N_5036);
nand U7557 (N_7557,N_4138,N_5161);
nor U7558 (N_7558,N_5708,N_4513);
and U7559 (N_7559,N_5144,N_5291);
nor U7560 (N_7560,N_4241,N_5012);
nor U7561 (N_7561,N_4951,N_4292);
nor U7562 (N_7562,N_4665,N_4940);
or U7563 (N_7563,N_5843,N_4813);
and U7564 (N_7564,N_4572,N_5547);
or U7565 (N_7565,N_5906,N_4710);
nand U7566 (N_7566,N_5901,N_5698);
nand U7567 (N_7567,N_5295,N_5577);
or U7568 (N_7568,N_5073,N_4509);
nand U7569 (N_7569,N_4821,N_5637);
or U7570 (N_7570,N_4332,N_4908);
nor U7571 (N_7571,N_5331,N_4496);
or U7572 (N_7572,N_4685,N_5970);
and U7573 (N_7573,N_4207,N_4085);
nor U7574 (N_7574,N_5342,N_5201);
nor U7575 (N_7575,N_4212,N_4120);
or U7576 (N_7576,N_5316,N_4577);
nand U7577 (N_7577,N_5059,N_4716);
nor U7578 (N_7578,N_4978,N_5492);
xnor U7579 (N_7579,N_5349,N_5631);
nand U7580 (N_7580,N_4272,N_5226);
and U7581 (N_7581,N_4985,N_4729);
nor U7582 (N_7582,N_4719,N_4567);
nor U7583 (N_7583,N_5812,N_4426);
or U7584 (N_7584,N_4244,N_4840);
and U7585 (N_7585,N_5757,N_4149);
nand U7586 (N_7586,N_5383,N_5362);
and U7587 (N_7587,N_4989,N_4848);
and U7588 (N_7588,N_5187,N_5606);
and U7589 (N_7589,N_5116,N_4459);
or U7590 (N_7590,N_4340,N_5752);
and U7591 (N_7591,N_4002,N_5232);
nor U7592 (N_7592,N_5553,N_4935);
xnor U7593 (N_7593,N_4570,N_5329);
or U7594 (N_7594,N_5321,N_5940);
xnor U7595 (N_7595,N_4841,N_5055);
nand U7596 (N_7596,N_5232,N_5176);
nor U7597 (N_7597,N_4497,N_5621);
or U7598 (N_7598,N_5187,N_5858);
or U7599 (N_7599,N_5004,N_4237);
and U7600 (N_7600,N_4106,N_5441);
or U7601 (N_7601,N_4540,N_5477);
or U7602 (N_7602,N_5261,N_4746);
nor U7603 (N_7603,N_4977,N_5008);
xnor U7604 (N_7604,N_4086,N_4962);
or U7605 (N_7605,N_5569,N_5540);
or U7606 (N_7606,N_5458,N_4326);
or U7607 (N_7607,N_4215,N_5860);
xor U7608 (N_7608,N_5249,N_4993);
xor U7609 (N_7609,N_4039,N_4091);
nor U7610 (N_7610,N_5124,N_4521);
nor U7611 (N_7611,N_4616,N_4648);
and U7612 (N_7612,N_4175,N_4725);
and U7613 (N_7613,N_4750,N_5873);
nand U7614 (N_7614,N_5026,N_4502);
xnor U7615 (N_7615,N_5893,N_4600);
nor U7616 (N_7616,N_4375,N_4431);
and U7617 (N_7617,N_4210,N_4390);
nor U7618 (N_7618,N_5945,N_5648);
or U7619 (N_7619,N_4307,N_4167);
or U7620 (N_7620,N_5165,N_4297);
nand U7621 (N_7621,N_4870,N_5860);
nor U7622 (N_7622,N_5763,N_4835);
nand U7623 (N_7623,N_4903,N_5619);
or U7624 (N_7624,N_4400,N_4905);
nor U7625 (N_7625,N_4481,N_5006);
and U7626 (N_7626,N_4375,N_4001);
or U7627 (N_7627,N_4693,N_5715);
or U7628 (N_7628,N_5897,N_4703);
nor U7629 (N_7629,N_4725,N_5287);
nor U7630 (N_7630,N_4526,N_4219);
and U7631 (N_7631,N_5783,N_5709);
and U7632 (N_7632,N_4713,N_4121);
and U7633 (N_7633,N_4610,N_4787);
xnor U7634 (N_7634,N_4409,N_5407);
and U7635 (N_7635,N_4214,N_5191);
and U7636 (N_7636,N_5011,N_5790);
nor U7637 (N_7637,N_4434,N_5444);
nor U7638 (N_7638,N_5057,N_5134);
nor U7639 (N_7639,N_4772,N_4866);
nor U7640 (N_7640,N_4346,N_5155);
nor U7641 (N_7641,N_5208,N_4561);
and U7642 (N_7642,N_4859,N_4299);
or U7643 (N_7643,N_5016,N_5407);
xor U7644 (N_7644,N_5421,N_5826);
or U7645 (N_7645,N_4197,N_5561);
or U7646 (N_7646,N_5873,N_4216);
nand U7647 (N_7647,N_5527,N_4990);
or U7648 (N_7648,N_4569,N_4825);
or U7649 (N_7649,N_4167,N_5713);
nand U7650 (N_7650,N_5938,N_4687);
nor U7651 (N_7651,N_5045,N_5840);
nor U7652 (N_7652,N_5252,N_5622);
nor U7653 (N_7653,N_5591,N_5373);
and U7654 (N_7654,N_4236,N_5279);
nand U7655 (N_7655,N_5585,N_4133);
and U7656 (N_7656,N_5957,N_4355);
or U7657 (N_7657,N_5763,N_5533);
and U7658 (N_7658,N_5853,N_5624);
and U7659 (N_7659,N_5570,N_5701);
or U7660 (N_7660,N_5905,N_4775);
or U7661 (N_7661,N_4536,N_5238);
and U7662 (N_7662,N_4096,N_4622);
nor U7663 (N_7663,N_4438,N_4453);
or U7664 (N_7664,N_4218,N_4437);
xor U7665 (N_7665,N_4730,N_5752);
xor U7666 (N_7666,N_5301,N_5891);
xor U7667 (N_7667,N_4705,N_4838);
nand U7668 (N_7668,N_5954,N_4234);
xor U7669 (N_7669,N_4233,N_5447);
and U7670 (N_7670,N_5026,N_5256);
and U7671 (N_7671,N_5618,N_5968);
nand U7672 (N_7672,N_4196,N_5071);
nor U7673 (N_7673,N_4254,N_5159);
and U7674 (N_7674,N_4314,N_4925);
xor U7675 (N_7675,N_5346,N_4742);
nor U7676 (N_7676,N_4690,N_4704);
nand U7677 (N_7677,N_4875,N_5963);
nand U7678 (N_7678,N_5792,N_4254);
nor U7679 (N_7679,N_5676,N_5073);
and U7680 (N_7680,N_4240,N_5723);
or U7681 (N_7681,N_5944,N_5008);
and U7682 (N_7682,N_5339,N_4465);
nor U7683 (N_7683,N_5911,N_5108);
or U7684 (N_7684,N_5703,N_5727);
and U7685 (N_7685,N_5805,N_5430);
nor U7686 (N_7686,N_5077,N_4882);
and U7687 (N_7687,N_5519,N_5024);
and U7688 (N_7688,N_4333,N_5796);
or U7689 (N_7689,N_4998,N_4711);
and U7690 (N_7690,N_4763,N_5156);
and U7691 (N_7691,N_5253,N_4848);
nor U7692 (N_7692,N_4447,N_5266);
nand U7693 (N_7693,N_4499,N_4924);
or U7694 (N_7694,N_4798,N_4353);
and U7695 (N_7695,N_4500,N_5991);
or U7696 (N_7696,N_4194,N_4950);
or U7697 (N_7697,N_4207,N_5494);
or U7698 (N_7698,N_4158,N_4813);
and U7699 (N_7699,N_4478,N_5716);
nor U7700 (N_7700,N_4778,N_4508);
or U7701 (N_7701,N_4642,N_5343);
nor U7702 (N_7702,N_4591,N_4540);
and U7703 (N_7703,N_4662,N_5396);
xor U7704 (N_7704,N_4560,N_4848);
or U7705 (N_7705,N_5341,N_4755);
or U7706 (N_7706,N_5133,N_4706);
xnor U7707 (N_7707,N_4218,N_4212);
and U7708 (N_7708,N_4122,N_5661);
nor U7709 (N_7709,N_4453,N_5555);
nand U7710 (N_7710,N_5162,N_4822);
nand U7711 (N_7711,N_4233,N_5319);
or U7712 (N_7712,N_5108,N_4408);
nor U7713 (N_7713,N_4843,N_4915);
xnor U7714 (N_7714,N_4000,N_4523);
and U7715 (N_7715,N_4140,N_5186);
nand U7716 (N_7716,N_4270,N_5811);
nor U7717 (N_7717,N_5625,N_4962);
or U7718 (N_7718,N_5372,N_5715);
nand U7719 (N_7719,N_4679,N_5737);
or U7720 (N_7720,N_5783,N_4956);
or U7721 (N_7721,N_4424,N_4378);
or U7722 (N_7722,N_5962,N_5451);
nor U7723 (N_7723,N_4531,N_5257);
and U7724 (N_7724,N_4911,N_4311);
nor U7725 (N_7725,N_4650,N_5851);
xor U7726 (N_7726,N_4205,N_4788);
or U7727 (N_7727,N_5053,N_4103);
nand U7728 (N_7728,N_4031,N_4514);
nand U7729 (N_7729,N_5174,N_5687);
xnor U7730 (N_7730,N_4970,N_4305);
and U7731 (N_7731,N_5172,N_5643);
nand U7732 (N_7732,N_5912,N_5836);
or U7733 (N_7733,N_5139,N_5969);
or U7734 (N_7734,N_5423,N_5442);
and U7735 (N_7735,N_5904,N_4721);
and U7736 (N_7736,N_5119,N_4560);
nand U7737 (N_7737,N_4948,N_4698);
nand U7738 (N_7738,N_4954,N_5913);
and U7739 (N_7739,N_4672,N_5527);
and U7740 (N_7740,N_5712,N_5885);
or U7741 (N_7741,N_5950,N_5726);
or U7742 (N_7742,N_4725,N_4438);
or U7743 (N_7743,N_4077,N_4887);
nand U7744 (N_7744,N_5472,N_5267);
or U7745 (N_7745,N_5927,N_4145);
xor U7746 (N_7746,N_5525,N_5313);
or U7747 (N_7747,N_4769,N_4811);
or U7748 (N_7748,N_4511,N_4345);
nor U7749 (N_7749,N_4839,N_5260);
nand U7750 (N_7750,N_4199,N_4423);
and U7751 (N_7751,N_5067,N_4686);
or U7752 (N_7752,N_5506,N_5197);
or U7753 (N_7753,N_5134,N_4689);
or U7754 (N_7754,N_5405,N_4908);
xor U7755 (N_7755,N_4173,N_5341);
nand U7756 (N_7756,N_5472,N_5803);
and U7757 (N_7757,N_4864,N_4934);
and U7758 (N_7758,N_5917,N_5364);
or U7759 (N_7759,N_4175,N_5079);
nand U7760 (N_7760,N_5177,N_5397);
nand U7761 (N_7761,N_4940,N_5668);
nor U7762 (N_7762,N_4637,N_4162);
nand U7763 (N_7763,N_5406,N_5865);
nand U7764 (N_7764,N_4877,N_4364);
nor U7765 (N_7765,N_4466,N_4375);
nand U7766 (N_7766,N_4286,N_4702);
and U7767 (N_7767,N_4211,N_5697);
or U7768 (N_7768,N_4219,N_4442);
nor U7769 (N_7769,N_5141,N_4364);
nor U7770 (N_7770,N_4788,N_4621);
nand U7771 (N_7771,N_4369,N_4782);
nor U7772 (N_7772,N_4459,N_5554);
and U7773 (N_7773,N_5664,N_5472);
and U7774 (N_7774,N_4847,N_4409);
and U7775 (N_7775,N_5086,N_4440);
and U7776 (N_7776,N_4098,N_5261);
and U7777 (N_7777,N_5160,N_4764);
or U7778 (N_7778,N_5932,N_4404);
nand U7779 (N_7779,N_4993,N_4338);
nor U7780 (N_7780,N_4599,N_5797);
or U7781 (N_7781,N_5153,N_5933);
nand U7782 (N_7782,N_5789,N_5985);
nor U7783 (N_7783,N_5494,N_4138);
and U7784 (N_7784,N_4277,N_4009);
nor U7785 (N_7785,N_5540,N_5394);
and U7786 (N_7786,N_4259,N_5398);
nand U7787 (N_7787,N_5124,N_4322);
or U7788 (N_7788,N_5961,N_5930);
nand U7789 (N_7789,N_4055,N_5181);
or U7790 (N_7790,N_4486,N_5674);
and U7791 (N_7791,N_5877,N_5247);
and U7792 (N_7792,N_4103,N_5459);
and U7793 (N_7793,N_5972,N_5123);
and U7794 (N_7794,N_4450,N_4778);
or U7795 (N_7795,N_4534,N_4308);
nand U7796 (N_7796,N_4454,N_5092);
nor U7797 (N_7797,N_4066,N_4261);
xor U7798 (N_7798,N_5333,N_5422);
xor U7799 (N_7799,N_5168,N_5953);
nand U7800 (N_7800,N_4824,N_5467);
or U7801 (N_7801,N_4716,N_4592);
and U7802 (N_7802,N_4745,N_5054);
nand U7803 (N_7803,N_4344,N_4050);
and U7804 (N_7804,N_5669,N_5487);
nor U7805 (N_7805,N_4801,N_5945);
nor U7806 (N_7806,N_4784,N_5053);
and U7807 (N_7807,N_4248,N_5084);
and U7808 (N_7808,N_5042,N_4296);
or U7809 (N_7809,N_4997,N_4938);
nor U7810 (N_7810,N_4799,N_4463);
or U7811 (N_7811,N_5951,N_4631);
and U7812 (N_7812,N_4055,N_5541);
nand U7813 (N_7813,N_4244,N_5372);
or U7814 (N_7814,N_4438,N_5142);
or U7815 (N_7815,N_5832,N_5954);
nand U7816 (N_7816,N_5508,N_4778);
nor U7817 (N_7817,N_5415,N_5558);
nor U7818 (N_7818,N_5402,N_5203);
nand U7819 (N_7819,N_4072,N_5044);
nand U7820 (N_7820,N_5652,N_5442);
nor U7821 (N_7821,N_5449,N_5975);
and U7822 (N_7822,N_5945,N_5793);
or U7823 (N_7823,N_5377,N_5757);
and U7824 (N_7824,N_4004,N_4159);
or U7825 (N_7825,N_5637,N_5537);
or U7826 (N_7826,N_5001,N_4135);
or U7827 (N_7827,N_4029,N_5417);
and U7828 (N_7828,N_5829,N_5712);
or U7829 (N_7829,N_4787,N_4085);
and U7830 (N_7830,N_5314,N_4290);
nor U7831 (N_7831,N_4084,N_4114);
nor U7832 (N_7832,N_4719,N_5162);
nor U7833 (N_7833,N_4864,N_5796);
nand U7834 (N_7834,N_5921,N_4424);
or U7835 (N_7835,N_5331,N_5425);
nor U7836 (N_7836,N_5119,N_5099);
nor U7837 (N_7837,N_5226,N_4437);
and U7838 (N_7838,N_4497,N_4001);
or U7839 (N_7839,N_5023,N_4756);
nor U7840 (N_7840,N_5193,N_4734);
or U7841 (N_7841,N_5339,N_4781);
nand U7842 (N_7842,N_4726,N_4829);
and U7843 (N_7843,N_4732,N_5516);
and U7844 (N_7844,N_4802,N_4037);
nor U7845 (N_7845,N_4087,N_5903);
nand U7846 (N_7846,N_4448,N_5008);
nand U7847 (N_7847,N_4619,N_5352);
and U7848 (N_7848,N_5096,N_4204);
and U7849 (N_7849,N_5863,N_4630);
nand U7850 (N_7850,N_4950,N_5598);
nand U7851 (N_7851,N_4511,N_5698);
nand U7852 (N_7852,N_5776,N_4990);
nor U7853 (N_7853,N_4068,N_4547);
nand U7854 (N_7854,N_5327,N_5940);
or U7855 (N_7855,N_5381,N_4787);
xnor U7856 (N_7856,N_4225,N_5779);
xor U7857 (N_7857,N_5881,N_4100);
xor U7858 (N_7858,N_5108,N_4214);
nand U7859 (N_7859,N_4159,N_4821);
and U7860 (N_7860,N_4553,N_5188);
nand U7861 (N_7861,N_4149,N_4534);
and U7862 (N_7862,N_4124,N_5728);
nor U7863 (N_7863,N_4364,N_5338);
nand U7864 (N_7864,N_4327,N_5336);
and U7865 (N_7865,N_4800,N_5100);
and U7866 (N_7866,N_5689,N_4776);
or U7867 (N_7867,N_4156,N_5362);
nor U7868 (N_7868,N_5180,N_4093);
nand U7869 (N_7869,N_5335,N_5814);
and U7870 (N_7870,N_5506,N_4233);
nor U7871 (N_7871,N_5798,N_5393);
xnor U7872 (N_7872,N_4692,N_4512);
nor U7873 (N_7873,N_5500,N_5040);
nor U7874 (N_7874,N_4980,N_4289);
xnor U7875 (N_7875,N_4915,N_5593);
nand U7876 (N_7876,N_5834,N_4926);
nor U7877 (N_7877,N_4319,N_4635);
nor U7878 (N_7878,N_4793,N_4313);
and U7879 (N_7879,N_5921,N_4413);
nand U7880 (N_7880,N_5845,N_5678);
and U7881 (N_7881,N_4225,N_5027);
nand U7882 (N_7882,N_5960,N_5607);
nand U7883 (N_7883,N_5738,N_5430);
or U7884 (N_7884,N_5166,N_4674);
and U7885 (N_7885,N_5520,N_5814);
nand U7886 (N_7886,N_4991,N_4003);
and U7887 (N_7887,N_5072,N_5440);
or U7888 (N_7888,N_4298,N_5491);
xor U7889 (N_7889,N_4559,N_5904);
xnor U7890 (N_7890,N_4666,N_5195);
or U7891 (N_7891,N_5262,N_4897);
nand U7892 (N_7892,N_5731,N_5516);
or U7893 (N_7893,N_4117,N_5886);
nand U7894 (N_7894,N_5141,N_5549);
or U7895 (N_7895,N_4928,N_4115);
or U7896 (N_7896,N_4313,N_5740);
or U7897 (N_7897,N_5263,N_5282);
or U7898 (N_7898,N_4051,N_5019);
nor U7899 (N_7899,N_5001,N_4576);
nor U7900 (N_7900,N_5996,N_4315);
nor U7901 (N_7901,N_4114,N_5262);
and U7902 (N_7902,N_5477,N_4765);
nand U7903 (N_7903,N_5512,N_4537);
nand U7904 (N_7904,N_4847,N_4181);
xor U7905 (N_7905,N_4280,N_5950);
nand U7906 (N_7906,N_5714,N_4490);
nor U7907 (N_7907,N_5932,N_4233);
xor U7908 (N_7908,N_5035,N_5733);
nand U7909 (N_7909,N_5640,N_4684);
xor U7910 (N_7910,N_4189,N_4108);
or U7911 (N_7911,N_4134,N_4200);
or U7912 (N_7912,N_5078,N_4230);
and U7913 (N_7913,N_4929,N_5035);
or U7914 (N_7914,N_4147,N_5030);
or U7915 (N_7915,N_5263,N_4121);
nand U7916 (N_7916,N_4463,N_4296);
nand U7917 (N_7917,N_4411,N_5283);
or U7918 (N_7918,N_4963,N_5549);
and U7919 (N_7919,N_5299,N_5243);
xnor U7920 (N_7920,N_5360,N_5007);
nor U7921 (N_7921,N_4025,N_5276);
or U7922 (N_7922,N_4852,N_4478);
nand U7923 (N_7923,N_4468,N_5662);
nor U7924 (N_7924,N_5022,N_4641);
nand U7925 (N_7925,N_5171,N_4237);
nand U7926 (N_7926,N_5967,N_4770);
and U7927 (N_7927,N_4840,N_4689);
nor U7928 (N_7928,N_5344,N_4384);
nand U7929 (N_7929,N_5446,N_4556);
nor U7930 (N_7930,N_4215,N_4845);
and U7931 (N_7931,N_4921,N_5868);
nor U7932 (N_7932,N_5072,N_4602);
nand U7933 (N_7933,N_4886,N_4717);
and U7934 (N_7934,N_4957,N_4963);
or U7935 (N_7935,N_4000,N_4859);
nor U7936 (N_7936,N_5946,N_5245);
or U7937 (N_7937,N_4409,N_5252);
or U7938 (N_7938,N_4615,N_4058);
or U7939 (N_7939,N_4848,N_5435);
and U7940 (N_7940,N_4977,N_5294);
nor U7941 (N_7941,N_5620,N_5457);
and U7942 (N_7942,N_4561,N_4133);
nor U7943 (N_7943,N_4005,N_4513);
nor U7944 (N_7944,N_5769,N_4884);
nor U7945 (N_7945,N_4964,N_5516);
nor U7946 (N_7946,N_4270,N_4137);
nor U7947 (N_7947,N_4202,N_4512);
nand U7948 (N_7948,N_5051,N_4273);
nor U7949 (N_7949,N_5669,N_4745);
xor U7950 (N_7950,N_4351,N_5036);
and U7951 (N_7951,N_5138,N_4017);
and U7952 (N_7952,N_4999,N_5964);
xnor U7953 (N_7953,N_5678,N_5749);
nor U7954 (N_7954,N_4256,N_4181);
nor U7955 (N_7955,N_4682,N_5065);
and U7956 (N_7956,N_5847,N_5623);
nor U7957 (N_7957,N_5837,N_4878);
or U7958 (N_7958,N_5518,N_5930);
or U7959 (N_7959,N_5137,N_5939);
and U7960 (N_7960,N_4107,N_4291);
nand U7961 (N_7961,N_5448,N_4885);
nor U7962 (N_7962,N_5255,N_5425);
nor U7963 (N_7963,N_4315,N_4185);
nor U7964 (N_7964,N_5979,N_4353);
nand U7965 (N_7965,N_4649,N_5840);
and U7966 (N_7966,N_5464,N_5781);
nand U7967 (N_7967,N_4652,N_4577);
xor U7968 (N_7968,N_5948,N_4663);
xor U7969 (N_7969,N_4583,N_4461);
nand U7970 (N_7970,N_5026,N_4169);
and U7971 (N_7971,N_5147,N_5771);
nor U7972 (N_7972,N_4507,N_5014);
xnor U7973 (N_7973,N_5849,N_4589);
nor U7974 (N_7974,N_4424,N_5568);
or U7975 (N_7975,N_5336,N_4006);
nor U7976 (N_7976,N_4898,N_5597);
xnor U7977 (N_7977,N_4987,N_4808);
and U7978 (N_7978,N_4221,N_5278);
and U7979 (N_7979,N_4251,N_4950);
nand U7980 (N_7980,N_5165,N_5077);
nor U7981 (N_7981,N_4679,N_4637);
and U7982 (N_7982,N_4738,N_4741);
and U7983 (N_7983,N_5945,N_5272);
nor U7984 (N_7984,N_5805,N_5792);
xor U7985 (N_7985,N_4594,N_4395);
and U7986 (N_7986,N_4022,N_5372);
and U7987 (N_7987,N_4848,N_5667);
or U7988 (N_7988,N_5739,N_5893);
nor U7989 (N_7989,N_5802,N_5284);
xnor U7990 (N_7990,N_5084,N_4753);
xor U7991 (N_7991,N_5443,N_4856);
nand U7992 (N_7992,N_5583,N_5249);
nor U7993 (N_7993,N_5555,N_4561);
or U7994 (N_7994,N_5774,N_5023);
nand U7995 (N_7995,N_5013,N_4249);
or U7996 (N_7996,N_4961,N_5679);
nor U7997 (N_7997,N_5737,N_4442);
nor U7998 (N_7998,N_5249,N_4102);
nor U7999 (N_7999,N_5896,N_4858);
and U8000 (N_8000,N_7068,N_6705);
nand U8001 (N_8001,N_7354,N_6586);
or U8002 (N_8002,N_7665,N_7848);
xnor U8003 (N_8003,N_6754,N_7855);
and U8004 (N_8004,N_7999,N_6522);
nand U8005 (N_8005,N_6882,N_7554);
and U8006 (N_8006,N_7419,N_6283);
and U8007 (N_8007,N_7424,N_6902);
nor U8008 (N_8008,N_6735,N_7019);
or U8009 (N_8009,N_6357,N_6079);
and U8010 (N_8010,N_6759,N_7044);
nand U8011 (N_8011,N_6342,N_6807);
nor U8012 (N_8012,N_6447,N_6276);
and U8013 (N_8013,N_7328,N_7616);
nor U8014 (N_8014,N_7923,N_7570);
nand U8015 (N_8015,N_6271,N_7789);
nor U8016 (N_8016,N_7064,N_7740);
xnor U8017 (N_8017,N_6279,N_7255);
or U8018 (N_8018,N_6779,N_7655);
or U8019 (N_8019,N_7608,N_6697);
nand U8020 (N_8020,N_6286,N_6461);
or U8021 (N_8021,N_7116,N_7784);
and U8022 (N_8022,N_6445,N_6041);
and U8023 (N_8023,N_7747,N_7672);
nor U8024 (N_8024,N_6804,N_6739);
and U8025 (N_8025,N_6275,N_7690);
xor U8026 (N_8026,N_7117,N_7439);
nand U8027 (N_8027,N_6856,N_6070);
xnor U8028 (N_8028,N_6703,N_7851);
and U8029 (N_8029,N_7399,N_7154);
and U8030 (N_8030,N_6732,N_7543);
nand U8031 (N_8031,N_7049,N_7664);
nor U8032 (N_8032,N_6415,N_6574);
nor U8033 (N_8033,N_6058,N_6277);
nand U8034 (N_8034,N_7507,N_6990);
nand U8035 (N_8035,N_7521,N_6570);
or U8036 (N_8036,N_7514,N_6490);
nor U8037 (N_8037,N_7421,N_6301);
nor U8038 (N_8038,N_7551,N_6323);
or U8039 (N_8039,N_7682,N_7921);
xnor U8040 (N_8040,N_7649,N_6519);
or U8041 (N_8041,N_7435,N_7752);
nand U8042 (N_8042,N_7646,N_7338);
nand U8043 (N_8043,N_6374,N_6842);
nand U8044 (N_8044,N_7363,N_7914);
and U8045 (N_8045,N_6532,N_6368);
or U8046 (N_8046,N_6840,N_7947);
and U8047 (N_8047,N_6404,N_7060);
and U8048 (N_8048,N_7323,N_7216);
or U8049 (N_8049,N_6941,N_6050);
xnor U8050 (N_8050,N_7810,N_6222);
nor U8051 (N_8051,N_6309,N_7557);
and U8052 (N_8052,N_7189,N_6505);
or U8053 (N_8053,N_7974,N_6425);
or U8054 (N_8054,N_7477,N_6051);
or U8055 (N_8055,N_6185,N_7148);
or U8056 (N_8056,N_7577,N_6053);
or U8057 (N_8057,N_6548,N_7245);
nor U8058 (N_8058,N_6282,N_7607);
nand U8059 (N_8059,N_7744,N_7517);
and U8060 (N_8060,N_7076,N_7907);
and U8061 (N_8061,N_7468,N_7768);
nor U8062 (N_8062,N_6326,N_7067);
nor U8063 (N_8063,N_7390,N_6546);
nand U8064 (N_8064,N_7005,N_6927);
nor U8065 (N_8065,N_6635,N_7047);
and U8066 (N_8066,N_7456,N_7425);
or U8067 (N_8067,N_7569,N_6375);
xor U8068 (N_8068,N_7769,N_6553);
and U8069 (N_8069,N_6600,N_7542);
nand U8070 (N_8070,N_7042,N_6813);
nor U8071 (N_8071,N_7678,N_7059);
or U8072 (N_8072,N_7611,N_6355);
or U8073 (N_8073,N_7164,N_6959);
xnor U8074 (N_8074,N_6075,N_7174);
and U8075 (N_8075,N_7736,N_7038);
or U8076 (N_8076,N_7699,N_7970);
nand U8077 (N_8077,N_7626,N_6479);
nor U8078 (N_8078,N_7509,N_7530);
and U8079 (N_8079,N_6741,N_6880);
nor U8080 (N_8080,N_7781,N_6698);
xor U8081 (N_8081,N_6560,N_7073);
nor U8082 (N_8082,N_7058,N_6469);
and U8083 (N_8083,N_6204,N_7968);
nand U8084 (N_8084,N_7162,N_6430);
nor U8085 (N_8085,N_7847,N_7290);
xor U8086 (N_8086,N_7670,N_6764);
or U8087 (N_8087,N_6762,N_6266);
nor U8088 (N_8088,N_7535,N_6508);
and U8089 (N_8089,N_7348,N_7911);
nand U8090 (N_8090,N_6158,N_7949);
and U8091 (N_8091,N_7955,N_7109);
or U8092 (N_8092,N_7802,N_7136);
or U8093 (N_8093,N_7175,N_7420);
xnor U8094 (N_8094,N_7447,N_6742);
xnor U8095 (N_8095,N_7428,N_7002);
or U8096 (N_8096,N_7078,N_6859);
and U8097 (N_8097,N_7644,N_6858);
and U8098 (N_8098,N_6230,N_7853);
nand U8099 (N_8099,N_6255,N_6778);
nand U8100 (N_8100,N_7755,N_6676);
nor U8101 (N_8101,N_7520,N_6181);
nand U8102 (N_8102,N_6552,N_7622);
nor U8103 (N_8103,N_7943,N_7777);
or U8104 (N_8104,N_7906,N_6881);
and U8105 (N_8105,N_6799,N_6908);
nor U8106 (N_8106,N_6573,N_7620);
or U8107 (N_8107,N_6884,N_6534);
and U8108 (N_8108,N_6809,N_7075);
nor U8109 (N_8109,N_6422,N_7088);
or U8110 (N_8110,N_6892,N_7180);
and U8111 (N_8111,N_7582,N_7774);
or U8112 (N_8112,N_6849,N_7751);
and U8113 (N_8113,N_7749,N_6584);
nor U8114 (N_8114,N_6599,N_6728);
or U8115 (N_8115,N_6943,N_7438);
or U8116 (N_8116,N_6776,N_7119);
nor U8117 (N_8117,N_6782,N_7578);
or U8118 (N_8118,N_7722,N_7294);
nand U8119 (N_8119,N_7273,N_7506);
xnor U8120 (N_8120,N_7219,N_7659);
or U8121 (N_8121,N_7131,N_6484);
nor U8122 (N_8122,N_6044,N_7138);
or U8123 (N_8123,N_7324,N_6605);
or U8124 (N_8124,N_6382,N_6246);
nand U8125 (N_8125,N_7391,N_7246);
nand U8126 (N_8126,N_6393,N_6085);
nand U8127 (N_8127,N_6037,N_6475);
and U8128 (N_8128,N_7220,N_7364);
and U8129 (N_8129,N_7203,N_7483);
and U8130 (N_8130,N_6839,N_7779);
nand U8131 (N_8131,N_7944,N_6977);
nand U8132 (N_8132,N_7077,N_7601);
nand U8133 (N_8133,N_6694,N_6032);
nand U8134 (N_8134,N_6285,N_6022);
xor U8135 (N_8135,N_6642,N_7964);
xnor U8136 (N_8136,N_6765,N_7927);
nand U8137 (N_8137,N_6607,N_7700);
nand U8138 (N_8138,N_6968,N_6156);
nand U8139 (N_8139,N_6601,N_6596);
xor U8140 (N_8140,N_6787,N_6583);
and U8141 (N_8141,N_7627,N_7368);
nor U8142 (N_8142,N_6094,N_7282);
nand U8143 (N_8143,N_7107,N_7981);
nor U8144 (N_8144,N_6589,N_7337);
or U8145 (N_8145,N_6630,N_6062);
and U8146 (N_8146,N_6870,N_6254);
or U8147 (N_8147,N_6716,N_7050);
nand U8148 (N_8148,N_6138,N_7919);
or U8149 (N_8149,N_7226,N_7941);
nor U8150 (N_8150,N_7718,N_6929);
nor U8151 (N_8151,N_6886,N_6503);
and U8152 (N_8152,N_7710,N_7493);
nand U8153 (N_8153,N_7153,N_7602);
nor U8154 (N_8154,N_7895,N_7634);
nor U8155 (N_8155,N_7029,N_6769);
nor U8156 (N_8156,N_6482,N_6480);
nor U8157 (N_8157,N_6499,N_6031);
nand U8158 (N_8158,N_7070,N_7978);
nand U8159 (N_8159,N_7928,N_6757);
nand U8160 (N_8160,N_6900,N_6825);
and U8161 (N_8161,N_7788,N_6916);
or U8162 (N_8162,N_6242,N_6449);
nand U8163 (N_8163,N_7773,N_7619);
nor U8164 (N_8164,N_6906,N_7563);
and U8165 (N_8165,N_6557,N_7152);
nor U8166 (N_8166,N_7207,N_7558);
nand U8167 (N_8167,N_7485,N_7685);
xor U8168 (N_8168,N_7086,N_7865);
nand U8169 (N_8169,N_6565,N_6695);
nand U8170 (N_8170,N_7315,N_7388);
nor U8171 (N_8171,N_6862,N_6452);
xnor U8172 (N_8172,N_7977,N_6917);
nand U8173 (N_8173,N_7043,N_7850);
or U8174 (N_8174,N_6590,N_7573);
nor U8175 (N_8175,N_6192,N_6626);
and U8176 (N_8176,N_7320,N_6260);
nor U8177 (N_8177,N_6946,N_7813);
or U8178 (N_8178,N_7552,N_6820);
and U8179 (N_8179,N_6481,N_6183);
nand U8180 (N_8180,N_6994,N_7271);
and U8181 (N_8181,N_6262,N_6344);
nand U8182 (N_8182,N_6702,N_6654);
nand U8183 (N_8183,N_7702,N_7357);
nor U8184 (N_8184,N_6010,N_7215);
nand U8185 (N_8185,N_7824,N_7142);
or U8186 (N_8186,N_6928,N_7403);
and U8187 (N_8187,N_7071,N_7385);
nor U8188 (N_8188,N_6609,N_6304);
and U8189 (N_8189,N_6024,N_6837);
or U8190 (N_8190,N_6738,N_7725);
or U8191 (N_8191,N_6296,N_6274);
and U8192 (N_8192,N_6592,N_7098);
xor U8193 (N_8193,N_6571,N_7798);
nand U8194 (N_8194,N_6633,N_6579);
nor U8195 (N_8195,N_7146,N_7816);
and U8196 (N_8196,N_6030,N_6352);
nor U8197 (N_8197,N_7475,N_6118);
nand U8198 (N_8198,N_6664,N_7597);
and U8199 (N_8199,N_7213,N_7492);
or U8200 (N_8200,N_6240,N_7952);
nor U8201 (N_8201,N_6369,N_7298);
nor U8202 (N_8202,N_7466,N_6073);
or U8203 (N_8203,N_6303,N_6652);
or U8204 (N_8204,N_7676,N_7680);
xnor U8205 (N_8205,N_7440,N_6487);
and U8206 (N_8206,N_6088,N_6507);
and U8207 (N_8207,N_6159,N_7459);
and U8208 (N_8208,N_7839,N_6077);
nor U8209 (N_8209,N_7464,N_7965);
and U8210 (N_8210,N_6965,N_6127);
nor U8211 (N_8211,N_6625,N_6029);
nand U8212 (N_8212,N_6023,N_7224);
nor U8213 (N_8213,N_7471,N_6896);
or U8214 (N_8214,N_6777,N_7147);
nand U8215 (N_8215,N_6651,N_6700);
or U8216 (N_8216,N_7904,N_6667);
and U8217 (N_8217,N_6647,N_7339);
nand U8218 (N_8218,N_6234,N_6253);
and U8219 (N_8219,N_6431,N_7361);
nand U8220 (N_8220,N_6749,N_6950);
and U8221 (N_8221,N_6349,N_6132);
or U8222 (N_8222,N_6019,N_7954);
or U8223 (N_8223,N_7272,N_7190);
nand U8224 (N_8224,N_6177,N_7818);
or U8225 (N_8225,N_6043,N_6243);
and U8226 (N_8226,N_6722,N_6049);
nor U8227 (N_8227,N_7922,N_6336);
xnor U8228 (N_8228,N_6383,N_7129);
nand U8229 (N_8229,N_7606,N_6551);
nand U8230 (N_8230,N_7931,N_6082);
or U8231 (N_8231,N_6021,N_6414);
nand U8232 (N_8232,N_6207,N_7861);
nand U8233 (N_8233,N_6934,N_7355);
nor U8234 (N_8234,N_7864,N_6151);
and U8235 (N_8235,N_7775,N_7946);
nand U8236 (N_8236,N_7441,N_7706);
and U8237 (N_8237,N_7961,N_6434);
nor U8238 (N_8238,N_6119,N_6143);
and U8239 (N_8239,N_7956,N_7504);
nor U8240 (N_8240,N_7694,N_6232);
or U8241 (N_8241,N_7892,N_7434);
xor U8242 (N_8242,N_6035,N_7958);
or U8243 (N_8243,N_6147,N_6515);
or U8244 (N_8244,N_6233,N_6623);
nor U8245 (N_8245,N_7080,N_6135);
or U8246 (N_8246,N_6624,N_6575);
or U8247 (N_8247,N_6729,N_7176);
or U8248 (N_8248,N_6270,N_6753);
nor U8249 (N_8249,N_6726,N_6918);
nor U8250 (N_8250,N_7111,N_6521);
nand U8251 (N_8251,N_6180,N_6381);
nor U8252 (N_8252,N_7327,N_7829);
and U8253 (N_8253,N_6331,N_6402);
or U8254 (N_8254,N_7442,N_6141);
nor U8255 (N_8255,N_6957,N_6198);
and U8256 (N_8256,N_6028,N_6974);
or U8257 (N_8257,N_6403,N_7647);
and U8258 (N_8258,N_7258,N_7598);
nor U8259 (N_8259,N_6872,N_7969);
nand U8260 (N_8260,N_6855,N_6910);
nor U8261 (N_8261,N_6125,N_7782);
nor U8262 (N_8262,N_6171,N_6712);
nor U8263 (N_8263,N_7871,N_6330);
xor U8264 (N_8264,N_7836,N_6953);
and U8265 (N_8265,N_7913,N_6106);
and U8266 (N_8266,N_7915,N_7643);
or U8267 (N_8267,N_7858,N_7177);
or U8268 (N_8268,N_6506,N_6766);
nand U8269 (N_8269,N_6743,N_7890);
or U8270 (N_8270,N_6737,N_6142);
and U8271 (N_8271,N_7395,N_6133);
nand U8272 (N_8272,N_6561,N_7663);
nand U8273 (N_8273,N_6289,N_7805);
and U8274 (N_8274,N_6078,N_7562);
nor U8275 (N_8275,N_6099,N_6148);
xor U8276 (N_8276,N_6670,N_6401);
nand U8277 (N_8277,N_7051,N_6907);
or U8278 (N_8278,N_7812,N_7971);
nand U8279 (N_8279,N_7486,N_6938);
xnor U8280 (N_8280,N_6163,N_6409);
nand U8281 (N_8281,N_6332,N_7287);
nand U8282 (N_8282,N_6400,N_7402);
or U8283 (N_8283,N_7645,N_6227);
nand U8284 (N_8284,N_7942,N_7863);
nor U8285 (N_8285,N_7584,N_6497);
nor U8286 (N_8286,N_7288,N_6850);
nor U8287 (N_8287,N_6912,N_6416);
or U8288 (N_8288,N_7345,N_7527);
nor U8289 (N_8289,N_7959,N_6576);
or U8290 (N_8290,N_6988,N_6975);
or U8291 (N_8291,N_6939,N_6366);
nand U8292 (N_8292,N_7589,N_7500);
nor U8293 (N_8293,N_6989,N_7040);
or U8294 (N_8294,N_7331,N_7344);
and U8295 (N_8295,N_6443,N_7349);
or U8296 (N_8296,N_6983,N_6115);
xnor U8297 (N_8297,N_6426,N_7405);
xnor U8298 (N_8298,N_6081,N_6423);
xnor U8299 (N_8299,N_6241,N_7408);
xnor U8300 (N_8300,N_6113,N_6788);
nor U8301 (N_8301,N_6815,N_7266);
nand U8302 (N_8302,N_7430,N_7329);
or U8303 (N_8303,N_6627,N_7992);
and U8304 (N_8304,N_6610,N_7732);
nand U8305 (N_8305,N_6209,N_6316);
and U8306 (N_8306,N_6772,N_7409);
nand U8307 (N_8307,N_6027,N_6001);
or U8308 (N_8308,N_7565,N_6930);
nand U8309 (N_8309,N_7362,N_6657);
nor U8310 (N_8310,N_7173,N_7593);
or U8311 (N_8311,N_7764,N_7874);
nand U8312 (N_8312,N_6608,N_6933);
and U8313 (N_8313,N_7238,N_7132);
nand U8314 (N_8314,N_6785,N_6827);
nand U8315 (N_8315,N_7975,N_7166);
nand U8316 (N_8316,N_7066,N_6725);
nand U8317 (N_8317,N_7794,N_7729);
nor U8318 (N_8318,N_7591,N_7041);
nand U8319 (N_8319,N_6202,N_6218);
or U8320 (N_8320,N_6587,N_6360);
and U8321 (N_8321,N_7698,N_6039);
or U8322 (N_8322,N_6767,N_6550);
or U8323 (N_8323,N_6682,N_6919);
or U8324 (N_8324,N_6294,N_6952);
xor U8325 (N_8325,N_7008,N_7118);
nand U8326 (N_8326,N_7575,N_6869);
nor U8327 (N_8327,N_7026,N_7145);
or U8328 (N_8328,N_7083,N_6922);
nand U8329 (N_8329,N_6976,N_7695);
nor U8330 (N_8330,N_7023,N_6543);
and U8331 (N_8331,N_6822,N_6714);
nand U8332 (N_8332,N_6281,N_6086);
and U8333 (N_8333,N_6853,N_6835);
nand U8334 (N_8334,N_7371,N_6894);
and U8335 (N_8335,N_7666,N_7667);
or U8336 (N_8336,N_6325,N_6478);
and U8337 (N_8337,N_6602,N_7418);
nor U8338 (N_8338,N_7717,N_7604);
and U8339 (N_8339,N_6925,N_6346);
and U8340 (N_8340,N_7738,N_7185);
nand U8341 (N_8341,N_6231,N_6102);
nor U8342 (N_8342,N_6693,N_7127);
and U8343 (N_8343,N_6083,N_7072);
or U8344 (N_8344,N_7708,N_6982);
or U8345 (N_8345,N_7003,N_7084);
nand U8346 (N_8346,N_7771,N_6666);
nor U8347 (N_8347,N_6069,N_6172);
xnor U8348 (N_8348,N_6878,N_6280);
nor U8349 (N_8349,N_7821,N_6092);
nor U8350 (N_8350,N_6969,N_6438);
or U8351 (N_8351,N_6628,N_6226);
nor U8352 (N_8352,N_6805,N_7024);
and U8353 (N_8353,N_7383,N_6887);
or U8354 (N_8354,N_7100,N_7511);
and U8355 (N_8355,N_6556,N_6129);
nor U8356 (N_8356,N_6686,N_7731);
and U8357 (N_8357,N_7297,N_7758);
and U8358 (N_8358,N_6370,N_7004);
and U8359 (N_8359,N_6828,N_7625);
and U8360 (N_8360,N_6225,N_6421);
or U8361 (N_8361,N_6056,N_7141);
and U8362 (N_8362,N_7536,N_6327);
or U8363 (N_8363,N_7962,N_6318);
nor U8364 (N_8364,N_6845,N_7237);
or U8365 (N_8365,N_7128,N_6756);
nor U8366 (N_8366,N_7687,N_7808);
xnor U8367 (N_8367,N_7735,N_7766);
and U8368 (N_8368,N_7534,N_7244);
xnor U8369 (N_8369,N_7233,N_6310);
nand U8370 (N_8370,N_6606,N_6992);
nand U8371 (N_8371,N_7691,N_7508);
nand U8372 (N_8372,N_7686,N_6942);
and U8373 (N_8373,N_6826,N_6410);
nor U8374 (N_8374,N_6528,N_7783);
or U8375 (N_8375,N_6167,N_6801);
and U8376 (N_8376,N_7759,N_6387);
nand U8377 (N_8377,N_7654,N_6354);
nand U8378 (N_8378,N_6932,N_6026);
and U8379 (N_8379,N_6643,N_7123);
nand U8380 (N_8380,N_7846,N_7559);
nand U8381 (N_8381,N_7924,N_6364);
or U8382 (N_8382,N_6103,N_7567);
nor U8383 (N_8383,N_6130,N_7202);
nand U8384 (N_8384,N_6834,N_6964);
or U8385 (N_8385,N_7704,N_6060);
nand U8386 (N_8386,N_6717,N_7115);
or U8387 (N_8387,N_7586,N_7025);
or U8388 (N_8388,N_6655,N_7436);
nor U8389 (N_8389,N_7413,N_7842);
xnor U8390 (N_8390,N_7837,N_6269);
nor U8391 (N_8391,N_6792,N_7746);
or U8392 (N_8392,N_6245,N_7679);
nor U8393 (N_8393,N_7204,N_6730);
nand U8394 (N_8394,N_7976,N_6559);
or U8395 (N_8395,N_7711,N_7417);
and U8396 (N_8396,N_6645,N_6340);
and U8397 (N_8397,N_7656,N_7229);
or U8398 (N_8398,N_6710,N_6263);
or U8399 (N_8399,N_6265,N_7636);
and U8400 (N_8400,N_6537,N_7762);
and U8401 (N_8401,N_7639,N_6208);
or U8402 (N_8402,N_7905,N_7519);
nand U8403 (N_8403,N_7491,N_6614);
nand U8404 (N_8404,N_7940,N_7222);
and U8405 (N_8405,N_7033,N_7300);
nand U8406 (N_8406,N_6157,N_6252);
or U8407 (N_8407,N_7510,N_7612);
or U8408 (N_8408,N_7487,N_6955);
nand U8409 (N_8409,N_6711,N_7986);
nand U8410 (N_8410,N_6101,N_6146);
nand U8411 (N_8411,N_7457,N_7130);
and U8412 (N_8412,N_6397,N_7133);
or U8413 (N_8413,N_7529,N_6257);
xnor U8414 (N_8414,N_7963,N_7372);
or U8415 (N_8415,N_6124,N_6526);
nor U8416 (N_8416,N_7550,N_6229);
nor U8417 (N_8417,N_6238,N_6413);
nor U8418 (N_8418,N_6420,N_7489);
or U8419 (N_8419,N_7617,N_7171);
xnor U8420 (N_8420,N_6109,N_7214);
and U8421 (N_8421,N_6205,N_7296);
and U8422 (N_8422,N_6436,N_7734);
and U8423 (N_8423,N_6709,N_6690);
xnor U8424 (N_8424,N_6384,N_6012);
nor U8425 (N_8425,N_6978,N_7209);
or U8426 (N_8426,N_7411,N_6396);
nand U8427 (N_8427,N_6439,N_7544);
nor U8428 (N_8428,N_6812,N_7165);
and U8429 (N_8429,N_6120,N_7887);
or U8430 (N_8430,N_7325,N_6678);
or U8431 (N_8431,N_6161,N_6187);
and U8432 (N_8432,N_7112,N_6220);
xnor U8433 (N_8433,N_7866,N_6372);
nor U8434 (N_8434,N_6493,N_7787);
nor U8435 (N_8435,N_7156,N_6456);
nor U8436 (N_8436,N_7289,N_6390);
or U8437 (N_8437,N_6668,N_7581);
and U8438 (N_8438,N_7106,N_6871);
nor U8439 (N_8439,N_6418,N_7313);
nand U8440 (N_8440,N_7767,N_7256);
nor U8441 (N_8441,N_6531,N_7467);
or U8442 (N_8442,N_7882,N_6446);
and U8443 (N_8443,N_7689,N_6006);
nor U8444 (N_8444,N_7994,N_6485);
or U8445 (N_8445,N_7228,N_7283);
or U8446 (N_8446,N_6793,N_6460);
and U8447 (N_8447,N_6221,N_6100);
and U8448 (N_8448,N_6833,N_7366);
xnor U8449 (N_8449,N_7832,N_7201);
and U8450 (N_8450,N_6914,N_7688);
nor U8451 (N_8451,N_7648,N_7316);
or U8452 (N_8452,N_6014,N_6137);
or U8453 (N_8453,N_7157,N_6860);
nand U8454 (N_8454,N_6477,N_6339);
nor U8455 (N_8455,N_7967,N_6541);
nand U8456 (N_8456,N_6305,N_7585);
and U8457 (N_8457,N_7079,N_7013);
nor U8458 (N_8458,N_7742,N_6816);
nand U8459 (N_8459,N_7675,N_6940);
or U8460 (N_8460,N_7849,N_7212);
nor U8461 (N_8461,N_7515,N_7929);
and U8462 (N_8462,N_7225,N_6800);
nand U8463 (N_8463,N_6677,N_6427);
and U8464 (N_8464,N_7367,N_6875);
xnor U8465 (N_8465,N_7948,N_7739);
or U8466 (N_8466,N_7628,N_7302);
and U8467 (N_8467,N_6435,N_6511);
nand U8468 (N_8468,N_7458,N_7538);
and U8469 (N_8469,N_6948,N_7712);
nor U8470 (N_8470,N_6966,N_6911);
nand U8471 (N_8471,N_7473,N_7737);
nor U8472 (N_8472,N_7274,N_7932);
or U8473 (N_8473,N_6162,N_7400);
or U8474 (N_8474,N_6903,N_6071);
and U8475 (N_8475,N_7281,N_6634);
or U8476 (N_8476,N_6065,N_7728);
and U8477 (N_8477,N_7785,N_7194);
and U8478 (N_8478,N_7444,N_7935);
xor U8479 (N_8479,N_6517,N_7295);
or U8480 (N_8480,N_7304,N_6046);
or U8481 (N_8481,N_6640,N_6611);
nand U8482 (N_8482,N_6453,N_7184);
nand U8483 (N_8483,N_6491,N_6052);
and U8484 (N_8484,N_6200,N_7482);
nor U8485 (N_8485,N_6954,N_6831);
xnor U8486 (N_8486,N_7898,N_7262);
xnor U8487 (N_8487,N_7183,N_6578);
nor U8488 (N_8488,N_6555,N_6740);
nor U8489 (N_8489,N_7134,N_7105);
or U8490 (N_8490,N_7450,N_7433);
and U8491 (N_8491,N_7208,N_6090);
xnor U8492 (N_8492,N_6199,N_7481);
nor U8493 (N_8493,N_7285,N_6501);
and U8494 (N_8494,N_7321,N_7776);
and U8495 (N_8495,N_6613,N_7571);
nand U8496 (N_8496,N_6140,N_7590);
or U8497 (N_8497,N_7632,N_6818);
and U8498 (N_8498,N_6495,N_6701);
and U8499 (N_8499,N_7650,N_7218);
and U8500 (N_8500,N_6399,N_7422);
nor U8501 (N_8501,N_6692,N_7843);
and U8502 (N_8502,N_7120,N_7104);
nand U8503 (N_8503,N_7760,N_7580);
nand U8504 (N_8504,N_6343,N_7406);
xnor U8505 (N_8505,N_6637,N_7753);
and U8506 (N_8506,N_7721,N_6388);
nand U8507 (N_8507,N_6371,N_7546);
or U8508 (N_8508,N_7502,N_7056);
and U8509 (N_8509,N_7251,N_6466);
or U8510 (N_8510,N_7236,N_6736);
xor U8511 (N_8511,N_7451,N_6945);
or U8512 (N_8512,N_6847,N_6707);
and U8513 (N_8513,N_6708,N_7280);
nor U8514 (N_8514,N_6385,N_6362);
or U8515 (N_8515,N_6504,N_7341);
xnor U8516 (N_8516,N_7340,N_7268);
nor U8517 (N_8517,N_6093,N_7693);
nand U8518 (N_8518,N_7637,N_7522);
nand U8519 (N_8519,N_6883,N_6525);
nand U8520 (N_8520,N_6193,N_7322);
nand U8521 (N_8521,N_7960,N_6873);
nand U8522 (N_8522,N_6554,N_6683);
and U8523 (N_8523,N_6971,N_7081);
nand U8524 (N_8524,N_7930,N_7099);
nor U8525 (N_8525,N_6061,N_6348);
nand U8526 (N_8526,N_7150,N_7793);
and U8527 (N_8527,N_7292,N_7819);
xor U8528 (N_8528,N_7181,N_6256);
nor U8529 (N_8529,N_7973,N_7653);
xnor U8530 (N_8530,N_7479,N_7566);
nor U8531 (N_8531,N_6530,N_6114);
nor U8532 (N_8532,N_6891,N_7091);
nand U8533 (N_8533,N_7378,N_6278);
xnor U8534 (N_8534,N_6259,N_6173);
nor U8535 (N_8535,N_7715,N_6632);
and U8536 (N_8536,N_7957,N_7726);
and U8537 (N_8537,N_7301,N_7560);
xnor U8538 (N_8538,N_6545,N_7488);
nor U8539 (N_8539,N_6136,N_6685);
nor U8540 (N_8540,N_7393,N_6080);
nor U8541 (N_8541,N_6798,N_6287);
nand U8542 (N_8542,N_6538,N_6733);
or U8543 (N_8543,N_7124,N_6470);
or U8544 (N_8544,N_7356,N_7614);
or U8545 (N_8545,N_7253,N_7140);
and U8546 (N_8546,N_7799,N_6638);
and U8547 (N_8547,N_7191,N_6539);
and U8548 (N_8548,N_6247,N_7917);
or U8549 (N_8549,N_7373,N_7270);
and U8550 (N_8550,N_6000,N_7265);
or U8551 (N_8551,N_7613,N_7114);
or U8552 (N_8552,N_7987,N_7903);
nor U8553 (N_8553,N_7461,N_6616);
nand U8554 (N_8554,N_7412,N_7350);
or U8555 (N_8555,N_7031,N_7852);
or U8556 (N_8556,N_7187,N_7092);
nor U8557 (N_8557,N_6644,N_6549);
and U8558 (N_8558,N_7293,N_7610);
nor U8559 (N_8559,N_6817,N_7370);
or U8560 (N_8560,N_6593,N_6688);
or U8561 (N_8561,N_7918,N_7668);
or U8562 (N_8562,N_6824,N_6025);
nand U8563 (N_8563,N_7242,N_6353);
and U8564 (N_8564,N_6631,N_6915);
nor U8565 (N_8565,N_6441,N_6373);
or U8566 (N_8566,N_6194,N_7404);
nand U8567 (N_8567,N_7048,N_6203);
xor U8568 (N_8568,N_7069,N_7885);
or U8569 (N_8569,N_6841,N_6621);
nor U8570 (N_8570,N_7772,N_7889);
nor U8571 (N_8571,N_7462,N_6582);
xnor U8572 (N_8572,N_6944,N_6433);
and U8573 (N_8573,N_6770,N_7791);
or U8574 (N_8574,N_6706,N_6214);
xor U8575 (N_8575,N_7902,N_6899);
and U8576 (N_8576,N_6797,N_7730);
nand U8577 (N_8577,N_7159,N_6224);
and U8578 (N_8578,N_6750,N_6182);
xor U8579 (N_8579,N_6540,N_6155);
or U8580 (N_8580,N_6991,N_6931);
nor U8581 (N_8581,N_7168,N_6498);
xor U8582 (N_8582,N_6312,N_7988);
nand U8583 (N_8583,N_7838,N_7375);
and U8584 (N_8584,N_6721,N_7696);
xnor U8585 (N_8585,N_6936,N_7476);
and U8586 (N_8586,N_7065,N_6923);
xnor U8587 (N_8587,N_6154,N_6486);
nor U8588 (N_8588,N_7426,N_7804);
or U8589 (N_8589,N_6217,N_6510);
nand U8590 (N_8590,N_7995,N_7684);
nand U8591 (N_8591,N_6144,N_6981);
and U8592 (N_8592,N_7155,N_7540);
xor U8593 (N_8593,N_6472,N_6746);
nor U8594 (N_8594,N_7910,N_7856);
or U8595 (N_8595,N_7920,N_7278);
or U8596 (N_8596,N_7936,N_6998);
and U8597 (N_8597,N_7063,N_7897);
nor U8598 (N_8598,N_7303,N_7006);
nor U8599 (N_8599,N_7835,N_6299);
or U8600 (N_8600,N_6329,N_7870);
and U8601 (N_8601,N_7651,N_7594);
nand U8602 (N_8602,N_7524,N_6066);
nand U8603 (N_8603,N_7991,N_7750);
nand U8604 (N_8604,N_6169,N_6720);
or U8605 (N_8605,N_6679,N_7110);
nor U8606 (N_8606,N_6680,N_6895);
nor U8607 (N_8607,N_6523,N_6865);
nor U8608 (N_8608,N_7326,N_7872);
or U8609 (N_8609,N_7352,N_6320);
nand U8610 (N_8610,N_6909,N_6297);
nor U8611 (N_8611,N_7093,N_7498);
xor U8612 (N_8612,N_6186,N_6488);
nor U8613 (N_8613,N_6361,N_7423);
and U8614 (N_8614,N_7478,N_7908);
xnor U8615 (N_8615,N_7223,N_7703);
nor U8616 (N_8616,N_6500,N_6057);
nand U8617 (N_8617,N_7778,N_7446);
and U8618 (N_8618,N_6832,N_7095);
and U8619 (N_8619,N_7392,N_7719);
or U8620 (N_8620,N_7556,N_6442);
or U8621 (N_8621,N_6411,N_7900);
and U8622 (N_8622,N_6313,N_6111);
or U8623 (N_8623,N_7279,N_6689);
nor U8624 (N_8624,N_6424,N_7925);
xnor U8625 (N_8625,N_7087,N_7227);
nor U8626 (N_8626,N_6580,N_7248);
nor U8627 (N_8627,N_6496,N_6806);
nor U8628 (N_8628,N_7609,N_6874);
nand U8629 (N_8629,N_6761,N_6572);
or U8630 (N_8630,N_6890,N_7912);
nor U8631 (N_8631,N_7454,N_7443);
and U8632 (N_8632,N_7583,N_6713);
and U8633 (N_8633,N_6660,N_6267);
and U8634 (N_8634,N_6684,N_7661);
nor U8635 (N_8635,N_7335,N_6175);
and U8636 (N_8636,N_6547,N_6150);
nor U8637 (N_8637,N_6512,N_7674);
nor U8638 (N_8638,N_6513,N_6317);
and U8639 (N_8639,N_6669,N_7307);
and U8640 (N_8640,N_7011,N_6112);
nand U8641 (N_8641,N_6567,N_7259);
nor U8642 (N_8642,N_7792,N_7193);
and U8643 (N_8643,N_6176,N_6731);
and U8644 (N_8644,N_6494,N_7990);
and U8645 (N_8645,N_6054,N_7333);
nor U8646 (N_8646,N_6836,N_6781);
and U8647 (N_8647,N_7501,N_6002);
and U8648 (N_8648,N_6064,N_7896);
nor U8649 (N_8649,N_7353,N_7603);
and U8650 (N_8650,N_6864,N_7770);
nand U8651 (N_8651,N_6951,N_6516);
xor U8652 (N_8652,N_6123,N_7455);
or U8653 (N_8653,N_6116,N_6350);
and U8654 (N_8654,N_6724,N_7939);
and U8655 (N_8655,N_6658,N_6937);
and U8656 (N_8656,N_7254,N_6314);
and U8657 (N_8657,N_7629,N_6018);
nor U8658 (N_8658,N_7801,N_6536);
nor U8659 (N_8659,N_6535,N_7757);
or U8660 (N_8660,N_7523,N_6365);
and U8661 (N_8661,N_7875,N_7239);
nand U8662 (N_8662,N_6876,N_6104);
and U8663 (N_8663,N_6188,N_6476);
and U8664 (N_8664,N_6577,N_6558);
nand U8665 (N_8665,N_6398,N_6780);
nor U8666 (N_8666,N_7669,N_7284);
or U8667 (N_8667,N_7564,N_6302);
nand U8668 (N_8668,N_7343,N_6802);
xnor U8669 (N_8669,N_6518,N_6542);
nor U8670 (N_8670,N_7480,N_7640);
or U8671 (N_8671,N_6451,N_6734);
nor U8672 (N_8672,N_6011,N_7036);
nor U8673 (N_8673,N_6636,N_7525);
and U8674 (N_8674,N_7319,N_7163);
and U8675 (N_8675,N_6956,N_7305);
or U8676 (N_8676,N_6126,N_7151);
nor U8677 (N_8677,N_7231,N_6394);
or U8678 (N_8678,N_6347,N_6960);
nand U8679 (N_8679,N_7260,N_6821);
nor U8680 (N_8680,N_6465,N_6790);
nand U8681 (N_8681,N_6190,N_7549);
nor U8682 (N_8682,N_6315,N_7122);
or U8683 (N_8683,N_6846,N_6897);
or U8684 (N_8684,N_6629,N_6893);
xor U8685 (N_8685,N_6432,N_7803);
and U8686 (N_8686,N_7526,N_6581);
nand U8687 (N_8687,N_6152,N_7600);
and U8688 (N_8688,N_6967,N_6857);
nor U8689 (N_8689,N_7539,N_6995);
and U8690 (N_8690,N_7877,N_7714);
nand U8691 (N_8691,N_7149,N_7630);
or U8692 (N_8692,N_7017,N_6904);
nor U8693 (N_8693,N_7448,N_6212);
nand U8694 (N_8694,N_6337,N_7061);
nand U8695 (N_8695,N_6696,N_6108);
xnor U8696 (N_8696,N_6017,N_7317);
nand U8697 (N_8697,N_7724,N_7179);
nor U8698 (N_8698,N_6921,N_6128);
or U8699 (N_8699,N_7334,N_6984);
and U8700 (N_8700,N_7822,N_7192);
nor U8701 (N_8701,N_6020,N_6844);
nor U8702 (N_8702,N_7276,N_7533);
or U8703 (N_8703,N_6087,N_6258);
xor U8704 (N_8704,N_6195,N_7720);
nand U8705 (N_8705,N_7496,N_6341);
or U8706 (N_8706,N_6356,N_7449);
and U8707 (N_8707,N_7094,N_6996);
nand U8708 (N_8708,N_7414,N_6250);
or U8709 (N_8709,N_6311,N_6174);
nand U8710 (N_8710,N_7101,N_7800);
xor U8711 (N_8711,N_6290,N_6795);
nand U8712 (N_8712,N_7828,N_6048);
nand U8713 (N_8713,N_6335,N_6999);
nand U8714 (N_8714,N_7673,N_7547);
or U8715 (N_8715,N_6013,N_6949);
or U8716 (N_8716,N_6751,N_7916);
xor U8717 (N_8717,N_6392,N_7823);
nand U8718 (N_8718,N_7234,N_6117);
and U8719 (N_8719,N_6533,N_6160);
and U8720 (N_8720,N_6924,N_7621);
nand U8721 (N_8721,N_6544,N_6704);
nand U8722 (N_8722,N_6009,N_7984);
or U8723 (N_8723,N_7881,N_6619);
and U8724 (N_8724,N_6196,N_7587);
or U8725 (N_8725,N_7859,N_7169);
or U8726 (N_8726,N_6620,N_6514);
nand U8727 (N_8727,N_6098,N_6288);
and U8728 (N_8728,N_7840,N_6848);
and U8729 (N_8729,N_7359,N_7474);
or U8730 (N_8730,N_6008,N_6178);
xnor U8731 (N_8731,N_6763,N_6040);
and U8732 (N_8732,N_7470,N_6829);
nand U8733 (N_8733,N_7756,N_7841);
nor U8734 (N_8734,N_7754,N_6378);
or U8735 (N_8735,N_6307,N_7347);
xnor U8736 (N_8736,N_7588,N_7427);
or U8737 (N_8737,N_7763,N_7379);
xor U8738 (N_8738,N_7827,N_7360);
or U8739 (N_8739,N_6055,N_6197);
or U8740 (N_8740,N_6851,N_6097);
nand U8741 (N_8741,N_6376,N_6211);
and U8742 (N_8742,N_7701,N_7980);
and U8743 (N_8743,N_7697,N_7553);
nand U8744 (N_8744,N_7358,N_6121);
or U8745 (N_8745,N_6189,N_6223);
nor U8746 (N_8746,N_6898,N_6963);
and U8747 (N_8747,N_6467,N_7018);
and U8748 (N_8748,N_6920,N_7662);
and U8749 (N_8749,N_6406,N_7318);
xnor U8750 (N_8750,N_7880,N_7232);
nor U8751 (N_8751,N_7716,N_7376);
and U8752 (N_8752,N_6168,N_6251);
nor U8753 (N_8753,N_6264,N_6889);
nor U8754 (N_8754,N_7709,N_7979);
nor U8755 (N_8755,N_7249,N_6673);
nor U8756 (N_8756,N_7250,N_7826);
nor U8757 (N_8757,N_7786,N_7888);
or U8758 (N_8758,N_7692,N_6237);
nand U8759 (N_8759,N_6206,N_7465);
nand U8760 (N_8760,N_6913,N_7096);
xnor U8761 (N_8761,N_7951,N_7257);
nor U8762 (N_8762,N_6681,N_7014);
nand U8763 (N_8763,N_6810,N_7909);
xor U8764 (N_8764,N_6389,N_7113);
or U8765 (N_8765,N_6653,N_7825);
and U8766 (N_8766,N_7139,N_7615);
and U8767 (N_8767,N_7592,N_6997);
or U8768 (N_8768,N_7452,N_6166);
and U8769 (N_8769,N_7045,N_7057);
xor U8770 (N_8770,N_6970,N_7997);
and U8771 (N_8771,N_6888,N_6489);
and U8772 (N_8772,N_7605,N_6184);
nand U8773 (N_8773,N_7332,N_6675);
or U8774 (N_8774,N_7365,N_6292);
nand U8775 (N_8775,N_7989,N_7886);
nor U8776 (N_8776,N_6661,N_7020);
xnor U8777 (N_8777,N_6284,N_7741);
or U8778 (N_8778,N_7167,N_7186);
and U8779 (N_8779,N_6437,N_7197);
or U8780 (N_8780,N_6867,N_6791);
and U8781 (N_8781,N_6755,N_6164);
or U8782 (N_8782,N_6509,N_7937);
and U8783 (N_8783,N_6215,N_7707);
nand U8784 (N_8784,N_7555,N_7765);
or U8785 (N_8785,N_6747,N_7369);
and U8786 (N_8786,N_7398,N_6134);
or U8787 (N_8787,N_6110,N_7878);
nor U8788 (N_8788,N_6719,N_7537);
or U8789 (N_8789,N_7623,N_6618);
nor U8790 (N_8790,N_7867,N_7311);
nand U8791 (N_8791,N_6321,N_7336);
nand U8792 (N_8792,N_6228,N_6905);
or U8793 (N_8793,N_6004,N_6170);
and U8794 (N_8794,N_7531,N_6760);
nand U8795 (N_8795,N_7382,N_6213);
nand U8796 (N_8796,N_6045,N_7873);
or U8797 (N_8797,N_6034,N_6646);
or U8798 (N_8798,N_7490,N_7235);
and U8799 (N_8799,N_7090,N_7381);
xor U8800 (N_8800,N_7007,N_7125);
nor U8801 (N_8801,N_6016,N_7576);
nor U8802 (N_8802,N_7683,N_7891);
and U8803 (N_8803,N_7857,N_6089);
xnor U8804 (N_8804,N_7346,N_6789);
and U8805 (N_8805,N_6568,N_7743);
nand U8806 (N_8806,N_6852,N_6239);
nor U8807 (N_8807,N_7195,N_7416);
nor U8808 (N_8808,N_6448,N_6985);
nand U8809 (N_8809,N_6139,N_7389);
or U8810 (N_8810,N_7545,N_7934);
and U8811 (N_8811,N_6492,N_7660);
nand U8812 (N_8812,N_6715,N_6773);
or U8813 (N_8813,N_6210,N_7291);
nand U8814 (N_8814,N_7121,N_7269);
nor U8815 (N_8815,N_7972,N_7437);
or U8816 (N_8816,N_7053,N_7460);
and U8817 (N_8817,N_6604,N_7267);
xor U8818 (N_8818,N_7484,N_7671);
nand U8819 (N_8819,N_6811,N_7055);
or U8820 (N_8820,N_6564,N_7351);
or U8821 (N_8821,N_6084,N_7631);
and U8822 (N_8822,N_7512,N_6322);
xnor U8823 (N_8823,N_6808,N_6622);
or U8824 (N_8824,N_7377,N_7796);
or U8825 (N_8825,N_6830,N_6775);
xnor U8826 (N_8826,N_7599,N_7009);
or U8827 (N_8827,N_7495,N_7314);
or U8828 (N_8828,N_6380,N_6784);
or U8829 (N_8829,N_6074,N_7286);
nor U8830 (N_8830,N_7384,N_7513);
xnor U8831 (N_8831,N_7021,N_6219);
and U8832 (N_8832,N_7854,N_6603);
or U8833 (N_8833,N_7844,N_6474);
nor U8834 (N_8834,N_7830,N_7950);
and U8835 (N_8835,N_7503,N_6351);
and U8836 (N_8836,N_6980,N_7182);
nor U8837 (N_8837,N_6615,N_6165);
and U8838 (N_8838,N_7401,N_6333);
or U8839 (N_8839,N_6444,N_7681);
nand U8840 (N_8840,N_7494,N_7170);
nand U8841 (N_8841,N_7178,N_6015);
and U8842 (N_8842,N_6718,N_6727);
and U8843 (N_8843,N_6529,N_6823);
or U8844 (N_8844,N_6562,N_6261);
and U8845 (N_8845,N_6563,N_7221);
and U8846 (N_8846,N_6300,N_6483);
and U8847 (N_8847,N_6377,N_7983);
and U8848 (N_8848,N_6674,N_7472);
nor U8849 (N_8849,N_6462,N_7993);
nor U8850 (N_8850,N_7733,N_6745);
or U8851 (N_8851,N_6650,N_7809);
nor U8852 (N_8852,N_7879,N_7938);
nor U8853 (N_8853,N_7985,N_7374);
or U8854 (N_8854,N_6149,N_7312);
nor U8855 (N_8855,N_6617,N_6405);
nor U8856 (N_8856,N_7407,N_7135);
or U8857 (N_8857,N_7723,N_7309);
or U8858 (N_8858,N_7306,N_7883);
xor U8859 (N_8859,N_6926,N_7966);
or U8860 (N_8860,N_6868,N_6866);
nand U8861 (N_8861,N_6987,N_6649);
xor U8862 (N_8862,N_6334,N_7211);
nand U8863 (N_8863,N_6972,N_7926);
and U8864 (N_8864,N_7431,N_6659);
or U8865 (N_8865,N_7532,N_7396);
or U8866 (N_8866,N_6291,N_7518);
nand U8867 (N_8867,N_7196,N_7205);
nor U8868 (N_8868,N_6819,N_7015);
nand U8869 (N_8869,N_7933,N_6463);
or U8870 (N_8870,N_6248,N_7869);
or U8871 (N_8871,N_6244,N_6961);
nor U8872 (N_8872,N_7032,N_6063);
and U8873 (N_8873,N_7275,N_7497);
nor U8874 (N_8874,N_7677,N_6973);
and U8875 (N_8875,N_7658,N_6429);
xnor U8876 (N_8876,N_6319,N_6007);
nand U8877 (N_8877,N_7945,N_7000);
nand U8878 (N_8878,N_7261,N_7039);
or U8879 (N_8879,N_6386,N_6662);
nor U8880 (N_8880,N_7642,N_7453);
or U8881 (N_8881,N_7263,N_6455);
nand U8882 (N_8882,N_6962,N_6408);
and U8883 (N_8883,N_7012,N_6363);
or U8884 (N_8884,N_7052,N_6458);
nor U8885 (N_8885,N_7572,N_7103);
nor U8886 (N_8886,N_7568,N_6520);
nor U8887 (N_8887,N_7505,N_7815);
and U8888 (N_8888,N_6993,N_6235);
and U8889 (N_8889,N_7862,N_7342);
nand U8890 (N_8890,N_6648,N_7126);
and U8891 (N_8891,N_7820,N_7618);
nor U8892 (N_8892,N_6379,N_6843);
xnor U8893 (N_8893,N_7469,N_7243);
and U8894 (N_8894,N_7579,N_7528);
and U8895 (N_8895,N_7834,N_6216);
nor U8896 (N_8896,N_6105,N_7814);
nor U8897 (N_8897,N_7996,N_7745);
or U8898 (N_8898,N_7574,N_7028);
nand U8899 (N_8899,N_7240,N_7241);
or U8900 (N_8900,N_7097,N_7144);
nor U8901 (N_8901,N_7633,N_6639);
nand U8902 (N_8902,N_7210,N_7198);
nand U8903 (N_8903,N_6338,N_6131);
nor U8904 (N_8904,N_6038,N_7035);
nand U8905 (N_8905,N_7387,N_6524);
and U8906 (N_8906,N_6440,N_7397);
or U8907 (N_8907,N_6814,N_6748);
nand U8908 (N_8908,N_7595,N_7108);
nor U8909 (N_8909,N_6468,N_6665);
nor U8910 (N_8910,N_7199,N_6308);
and U8911 (N_8911,N_6691,N_6663);
or U8912 (N_8912,N_6854,N_7230);
or U8913 (N_8913,N_6358,N_6298);
or U8914 (N_8914,N_7089,N_7868);
or U8915 (N_8915,N_7022,N_6771);
or U8916 (N_8916,N_7780,N_6145);
or U8917 (N_8917,N_6272,N_7380);
xor U8918 (N_8918,N_7217,N_7102);
nand U8919 (N_8919,N_7884,N_6588);
or U8920 (N_8920,N_6598,N_6095);
xor U8921 (N_8921,N_7160,N_6047);
xnor U8922 (N_8922,N_7806,N_7463);
nor U8923 (N_8923,N_6885,N_7206);
and U8924 (N_8924,N_7713,N_6059);
and U8925 (N_8925,N_7761,N_6459);
and U8926 (N_8926,N_7085,N_7062);
nand U8927 (N_8927,N_6324,N_7860);
nand U8928 (N_8928,N_7705,N_7016);
nand U8929 (N_8929,N_6671,N_6947);
nand U8930 (N_8930,N_6612,N_6419);
nor U8931 (N_8931,N_6122,N_7748);
nand U8932 (N_8932,N_7415,N_7264);
or U8933 (N_8933,N_6863,N_6179);
xnor U8934 (N_8934,N_6768,N_7445);
or U8935 (N_8935,N_7657,N_6412);
or U8936 (N_8936,N_7516,N_7833);
and U8937 (N_8937,N_7635,N_6794);
nand U8938 (N_8938,N_6838,N_6774);
xor U8939 (N_8939,N_7299,N_7624);
or U8940 (N_8940,N_6457,N_6407);
or U8941 (N_8941,N_6107,N_6901);
xnor U8942 (N_8942,N_6861,N_6033);
or U8943 (N_8943,N_7172,N_6752);
nand U8944 (N_8944,N_7727,N_6036);
xor U8945 (N_8945,N_6641,N_6796);
and U8946 (N_8946,N_7432,N_6687);
nor U8947 (N_8947,N_7797,N_6473);
and U8948 (N_8948,N_6656,N_6153);
or U8949 (N_8949,N_6003,N_6464);
or U8950 (N_8950,N_6958,N_6471);
xnor U8951 (N_8951,N_7790,N_6454);
nand U8952 (N_8952,N_7034,N_7074);
nor U8953 (N_8953,N_6201,N_6345);
xnor U8954 (N_8954,N_6594,N_7308);
xor U8955 (N_8955,N_6367,N_7831);
and U8956 (N_8956,N_6359,N_7310);
nor U8957 (N_8957,N_7158,N_6042);
xnor U8958 (N_8958,N_6803,N_7330);
or U8959 (N_8959,N_6597,N_7410);
nand U8960 (N_8960,N_6273,N_7054);
nand U8961 (N_8961,N_7817,N_7638);
nand U8962 (N_8962,N_7596,N_6450);
and U8963 (N_8963,N_6076,N_6758);
nand U8964 (N_8964,N_7188,N_6672);
nand U8965 (N_8965,N_7807,N_7143);
nor U8966 (N_8966,N_6879,N_6566);
nand U8967 (N_8967,N_7953,N_6986);
xor U8968 (N_8968,N_6249,N_6502);
nand U8969 (N_8969,N_6979,N_6786);
nor U8970 (N_8970,N_7998,N_6306);
nand U8971 (N_8971,N_6723,N_7027);
or U8972 (N_8972,N_7046,N_7561);
nand U8973 (N_8973,N_7252,N_7247);
and U8974 (N_8974,N_7161,N_6783);
nand U8975 (N_8975,N_7030,N_6744);
nand U8976 (N_8976,N_7082,N_7876);
nor U8977 (N_8977,N_6527,N_7001);
and U8978 (N_8978,N_6068,N_6067);
nor U8979 (N_8979,N_7429,N_7641);
or U8980 (N_8980,N_7894,N_6395);
and U8981 (N_8981,N_6935,N_7394);
nor U8982 (N_8982,N_6293,N_7010);
and U8983 (N_8983,N_7137,N_7277);
and U8984 (N_8984,N_6005,N_6569);
nor U8985 (N_8985,N_6428,N_7845);
and U8986 (N_8986,N_6699,N_7541);
nand U8987 (N_8987,N_7901,N_7386);
and U8988 (N_8988,N_6191,N_7499);
nand U8989 (N_8989,N_6096,N_7811);
nand U8990 (N_8990,N_7037,N_6877);
or U8991 (N_8991,N_7795,N_6072);
nand U8992 (N_8992,N_6295,N_6585);
nand U8993 (N_8993,N_7899,N_6328);
and U8994 (N_8994,N_6236,N_7548);
nor U8995 (N_8995,N_6417,N_6268);
xor U8996 (N_8996,N_7200,N_6591);
nor U8997 (N_8997,N_6091,N_7652);
nor U8998 (N_8998,N_7982,N_7893);
or U8999 (N_8999,N_6595,N_6391);
or U9000 (N_9000,N_7540,N_7052);
xnor U9001 (N_9001,N_7749,N_7646);
nand U9002 (N_9002,N_7431,N_6546);
and U9003 (N_9003,N_7608,N_7374);
nor U9004 (N_9004,N_6774,N_6672);
nor U9005 (N_9005,N_6059,N_7490);
and U9006 (N_9006,N_7656,N_6595);
nand U9007 (N_9007,N_6747,N_6971);
or U9008 (N_9008,N_6138,N_6518);
nor U9009 (N_9009,N_7180,N_7930);
nand U9010 (N_9010,N_6320,N_7805);
nand U9011 (N_9011,N_6703,N_6397);
nand U9012 (N_9012,N_6868,N_7283);
or U9013 (N_9013,N_7288,N_6913);
or U9014 (N_9014,N_7539,N_6519);
and U9015 (N_9015,N_7738,N_6328);
nand U9016 (N_9016,N_6890,N_6192);
and U9017 (N_9017,N_6635,N_6466);
or U9018 (N_9018,N_6767,N_7408);
xnor U9019 (N_9019,N_7585,N_6343);
nand U9020 (N_9020,N_6029,N_7143);
nor U9021 (N_9021,N_7770,N_7020);
and U9022 (N_9022,N_7286,N_7139);
nand U9023 (N_9023,N_6632,N_7020);
nand U9024 (N_9024,N_7738,N_6612);
nor U9025 (N_9025,N_7855,N_6906);
nor U9026 (N_9026,N_7610,N_6851);
nand U9027 (N_9027,N_7980,N_6259);
and U9028 (N_9028,N_7542,N_7323);
or U9029 (N_9029,N_6891,N_7992);
and U9030 (N_9030,N_6421,N_7629);
or U9031 (N_9031,N_6812,N_7314);
and U9032 (N_9032,N_6188,N_6359);
nand U9033 (N_9033,N_7383,N_6419);
nand U9034 (N_9034,N_7190,N_6045);
or U9035 (N_9035,N_6613,N_6657);
nand U9036 (N_9036,N_6657,N_7827);
nand U9037 (N_9037,N_6510,N_7319);
and U9038 (N_9038,N_6900,N_7117);
and U9039 (N_9039,N_7040,N_6087);
xor U9040 (N_9040,N_6627,N_7498);
and U9041 (N_9041,N_7315,N_7546);
and U9042 (N_9042,N_7078,N_7208);
and U9043 (N_9043,N_7564,N_7909);
nand U9044 (N_9044,N_6718,N_7854);
and U9045 (N_9045,N_6071,N_6070);
or U9046 (N_9046,N_6896,N_6863);
nand U9047 (N_9047,N_6716,N_7607);
nand U9048 (N_9048,N_6685,N_6230);
nor U9049 (N_9049,N_7274,N_7641);
and U9050 (N_9050,N_7422,N_7247);
or U9051 (N_9051,N_7074,N_7456);
and U9052 (N_9052,N_7181,N_7926);
nor U9053 (N_9053,N_6070,N_6074);
and U9054 (N_9054,N_7017,N_6228);
nand U9055 (N_9055,N_7291,N_6749);
nor U9056 (N_9056,N_6330,N_6286);
or U9057 (N_9057,N_6100,N_7722);
and U9058 (N_9058,N_6124,N_6504);
and U9059 (N_9059,N_7155,N_6575);
and U9060 (N_9060,N_7572,N_6952);
or U9061 (N_9061,N_6217,N_6688);
nand U9062 (N_9062,N_6487,N_7378);
nand U9063 (N_9063,N_6654,N_6601);
nand U9064 (N_9064,N_6219,N_6776);
and U9065 (N_9065,N_6374,N_7696);
and U9066 (N_9066,N_6258,N_6391);
nand U9067 (N_9067,N_7372,N_7732);
or U9068 (N_9068,N_7938,N_7800);
nand U9069 (N_9069,N_6650,N_6946);
or U9070 (N_9070,N_6521,N_6593);
nor U9071 (N_9071,N_7190,N_6241);
nand U9072 (N_9072,N_6084,N_7580);
and U9073 (N_9073,N_7989,N_6542);
nand U9074 (N_9074,N_7804,N_7733);
nand U9075 (N_9075,N_6481,N_7860);
nand U9076 (N_9076,N_7089,N_7719);
nand U9077 (N_9077,N_6156,N_6270);
nor U9078 (N_9078,N_7992,N_7954);
nor U9079 (N_9079,N_6703,N_7057);
nor U9080 (N_9080,N_7820,N_7047);
or U9081 (N_9081,N_7064,N_7581);
and U9082 (N_9082,N_7350,N_6328);
and U9083 (N_9083,N_7880,N_7124);
nor U9084 (N_9084,N_7363,N_7027);
nor U9085 (N_9085,N_7874,N_7179);
or U9086 (N_9086,N_7407,N_6642);
nand U9087 (N_9087,N_6427,N_6909);
nor U9088 (N_9088,N_7848,N_6845);
or U9089 (N_9089,N_7097,N_7462);
and U9090 (N_9090,N_6959,N_7182);
nand U9091 (N_9091,N_7102,N_7745);
xor U9092 (N_9092,N_6328,N_7449);
and U9093 (N_9093,N_7980,N_7550);
nand U9094 (N_9094,N_6102,N_6456);
and U9095 (N_9095,N_7355,N_6232);
xor U9096 (N_9096,N_7063,N_6155);
and U9097 (N_9097,N_7050,N_6467);
or U9098 (N_9098,N_7824,N_6769);
or U9099 (N_9099,N_6317,N_7137);
and U9100 (N_9100,N_7017,N_7421);
nor U9101 (N_9101,N_7063,N_7614);
and U9102 (N_9102,N_7156,N_6315);
and U9103 (N_9103,N_6348,N_6460);
nand U9104 (N_9104,N_7658,N_7610);
or U9105 (N_9105,N_7057,N_7379);
or U9106 (N_9106,N_6010,N_6962);
nor U9107 (N_9107,N_7351,N_6018);
nand U9108 (N_9108,N_6700,N_7949);
and U9109 (N_9109,N_6392,N_6371);
nand U9110 (N_9110,N_6437,N_6293);
or U9111 (N_9111,N_6056,N_6952);
or U9112 (N_9112,N_6990,N_7821);
and U9113 (N_9113,N_7131,N_7010);
or U9114 (N_9114,N_7192,N_7203);
nand U9115 (N_9115,N_7464,N_6534);
xor U9116 (N_9116,N_7017,N_6268);
nor U9117 (N_9117,N_6941,N_7930);
nor U9118 (N_9118,N_6098,N_7745);
nand U9119 (N_9119,N_7321,N_7118);
nand U9120 (N_9120,N_6888,N_6562);
or U9121 (N_9121,N_7979,N_6985);
nand U9122 (N_9122,N_7549,N_7850);
and U9123 (N_9123,N_7251,N_7669);
nand U9124 (N_9124,N_7366,N_7364);
nand U9125 (N_9125,N_7745,N_6605);
and U9126 (N_9126,N_7626,N_7174);
nand U9127 (N_9127,N_6302,N_7717);
nand U9128 (N_9128,N_6375,N_6058);
and U9129 (N_9129,N_7761,N_6657);
nand U9130 (N_9130,N_7459,N_7179);
or U9131 (N_9131,N_6018,N_6082);
nor U9132 (N_9132,N_6333,N_6308);
or U9133 (N_9133,N_6766,N_7927);
nor U9134 (N_9134,N_7707,N_6650);
and U9135 (N_9135,N_6802,N_7173);
nand U9136 (N_9136,N_7414,N_7688);
nor U9137 (N_9137,N_6543,N_6152);
xor U9138 (N_9138,N_7765,N_7961);
nand U9139 (N_9139,N_7809,N_6151);
nor U9140 (N_9140,N_7061,N_7163);
nand U9141 (N_9141,N_7117,N_7985);
nand U9142 (N_9142,N_7224,N_7199);
or U9143 (N_9143,N_6750,N_7589);
nor U9144 (N_9144,N_7610,N_7915);
or U9145 (N_9145,N_7184,N_7975);
nor U9146 (N_9146,N_7022,N_7885);
and U9147 (N_9147,N_7423,N_6794);
nor U9148 (N_9148,N_7730,N_7997);
and U9149 (N_9149,N_6358,N_7641);
nand U9150 (N_9150,N_6546,N_6861);
and U9151 (N_9151,N_6961,N_6578);
and U9152 (N_9152,N_7340,N_7573);
or U9153 (N_9153,N_6428,N_7326);
xor U9154 (N_9154,N_7730,N_7882);
nor U9155 (N_9155,N_6210,N_7461);
and U9156 (N_9156,N_6414,N_6667);
nor U9157 (N_9157,N_7001,N_7746);
or U9158 (N_9158,N_7054,N_6203);
and U9159 (N_9159,N_6304,N_7689);
xnor U9160 (N_9160,N_6980,N_7186);
or U9161 (N_9161,N_6823,N_6836);
xor U9162 (N_9162,N_6818,N_6019);
or U9163 (N_9163,N_7823,N_7702);
xor U9164 (N_9164,N_7724,N_7313);
xor U9165 (N_9165,N_7089,N_7070);
nand U9166 (N_9166,N_6781,N_6556);
and U9167 (N_9167,N_7944,N_6663);
and U9168 (N_9168,N_7490,N_7698);
nor U9169 (N_9169,N_6880,N_6660);
and U9170 (N_9170,N_7180,N_7457);
and U9171 (N_9171,N_7217,N_6316);
nor U9172 (N_9172,N_6409,N_6528);
nand U9173 (N_9173,N_7986,N_6999);
nor U9174 (N_9174,N_6149,N_7440);
nand U9175 (N_9175,N_6198,N_6435);
nand U9176 (N_9176,N_7374,N_7582);
nand U9177 (N_9177,N_6140,N_7227);
nor U9178 (N_9178,N_6483,N_7411);
or U9179 (N_9179,N_6645,N_7675);
nand U9180 (N_9180,N_7929,N_7825);
nor U9181 (N_9181,N_6508,N_7492);
nor U9182 (N_9182,N_6352,N_6767);
nand U9183 (N_9183,N_7925,N_6350);
xnor U9184 (N_9184,N_6697,N_6479);
nand U9185 (N_9185,N_6757,N_7698);
nand U9186 (N_9186,N_6817,N_7912);
nand U9187 (N_9187,N_7297,N_6174);
nand U9188 (N_9188,N_6135,N_6940);
nand U9189 (N_9189,N_7446,N_7484);
nand U9190 (N_9190,N_6970,N_7880);
or U9191 (N_9191,N_6190,N_7162);
nand U9192 (N_9192,N_6887,N_7482);
or U9193 (N_9193,N_7321,N_6956);
and U9194 (N_9194,N_6504,N_7385);
xnor U9195 (N_9195,N_6264,N_6136);
nor U9196 (N_9196,N_6867,N_7187);
and U9197 (N_9197,N_7613,N_7609);
nor U9198 (N_9198,N_6354,N_7785);
xor U9199 (N_9199,N_6157,N_7941);
and U9200 (N_9200,N_6928,N_7447);
nor U9201 (N_9201,N_7446,N_6075);
or U9202 (N_9202,N_7741,N_7775);
and U9203 (N_9203,N_7327,N_7133);
nand U9204 (N_9204,N_6496,N_6306);
nor U9205 (N_9205,N_7427,N_6985);
nand U9206 (N_9206,N_7666,N_6516);
or U9207 (N_9207,N_6889,N_6689);
nor U9208 (N_9208,N_7888,N_6354);
and U9209 (N_9209,N_6186,N_7749);
and U9210 (N_9210,N_6707,N_6405);
or U9211 (N_9211,N_7666,N_6628);
or U9212 (N_9212,N_6445,N_6378);
nand U9213 (N_9213,N_7984,N_6013);
nor U9214 (N_9214,N_6098,N_7283);
nand U9215 (N_9215,N_7760,N_7238);
nand U9216 (N_9216,N_6156,N_7195);
xor U9217 (N_9217,N_6787,N_6614);
nand U9218 (N_9218,N_6836,N_6204);
or U9219 (N_9219,N_6770,N_7521);
or U9220 (N_9220,N_6228,N_7461);
or U9221 (N_9221,N_6010,N_6372);
nor U9222 (N_9222,N_7140,N_6535);
nor U9223 (N_9223,N_7772,N_6751);
xor U9224 (N_9224,N_6272,N_7045);
nand U9225 (N_9225,N_7612,N_6729);
nand U9226 (N_9226,N_6096,N_6414);
or U9227 (N_9227,N_7432,N_6711);
and U9228 (N_9228,N_6635,N_6843);
or U9229 (N_9229,N_7908,N_7438);
nor U9230 (N_9230,N_6830,N_6726);
nand U9231 (N_9231,N_7597,N_6730);
nor U9232 (N_9232,N_6974,N_7296);
nor U9233 (N_9233,N_6575,N_7866);
or U9234 (N_9234,N_7839,N_6817);
nand U9235 (N_9235,N_7244,N_6427);
or U9236 (N_9236,N_6180,N_6232);
nor U9237 (N_9237,N_7575,N_7443);
nor U9238 (N_9238,N_7186,N_7164);
nand U9239 (N_9239,N_7587,N_7525);
nand U9240 (N_9240,N_7415,N_6984);
xor U9241 (N_9241,N_7887,N_6549);
and U9242 (N_9242,N_6843,N_6024);
nand U9243 (N_9243,N_6667,N_7997);
xor U9244 (N_9244,N_6471,N_7466);
or U9245 (N_9245,N_6643,N_6502);
nor U9246 (N_9246,N_7365,N_7997);
or U9247 (N_9247,N_7985,N_6441);
nor U9248 (N_9248,N_6670,N_7242);
or U9249 (N_9249,N_6641,N_7820);
nor U9250 (N_9250,N_7470,N_7244);
or U9251 (N_9251,N_7783,N_6716);
xor U9252 (N_9252,N_7992,N_6335);
nor U9253 (N_9253,N_7934,N_7925);
and U9254 (N_9254,N_6984,N_7368);
and U9255 (N_9255,N_7571,N_6303);
and U9256 (N_9256,N_6418,N_7126);
and U9257 (N_9257,N_6040,N_6588);
nor U9258 (N_9258,N_6712,N_7941);
nor U9259 (N_9259,N_6307,N_6047);
nand U9260 (N_9260,N_7053,N_6340);
and U9261 (N_9261,N_7730,N_7437);
or U9262 (N_9262,N_7033,N_7118);
xor U9263 (N_9263,N_7537,N_7434);
nand U9264 (N_9264,N_7693,N_7194);
and U9265 (N_9265,N_6174,N_7735);
and U9266 (N_9266,N_7794,N_6349);
or U9267 (N_9267,N_6068,N_7373);
xor U9268 (N_9268,N_6394,N_7004);
nand U9269 (N_9269,N_6607,N_7450);
xor U9270 (N_9270,N_7158,N_6184);
nor U9271 (N_9271,N_6392,N_6877);
or U9272 (N_9272,N_6778,N_7137);
or U9273 (N_9273,N_7137,N_6938);
or U9274 (N_9274,N_7102,N_6054);
xor U9275 (N_9275,N_6813,N_6157);
and U9276 (N_9276,N_7850,N_7426);
xnor U9277 (N_9277,N_6357,N_7536);
or U9278 (N_9278,N_7082,N_6735);
xor U9279 (N_9279,N_6501,N_6739);
xor U9280 (N_9280,N_6807,N_6114);
and U9281 (N_9281,N_7611,N_6026);
and U9282 (N_9282,N_7272,N_6654);
xnor U9283 (N_9283,N_7301,N_7378);
or U9284 (N_9284,N_7581,N_6050);
or U9285 (N_9285,N_7506,N_6727);
nand U9286 (N_9286,N_6929,N_6529);
or U9287 (N_9287,N_6775,N_6628);
and U9288 (N_9288,N_6951,N_6429);
or U9289 (N_9289,N_7638,N_6707);
nand U9290 (N_9290,N_6859,N_6525);
nor U9291 (N_9291,N_6111,N_6796);
or U9292 (N_9292,N_7109,N_6075);
or U9293 (N_9293,N_7968,N_6888);
nand U9294 (N_9294,N_7404,N_7837);
or U9295 (N_9295,N_7784,N_7890);
and U9296 (N_9296,N_7375,N_6517);
nor U9297 (N_9297,N_6724,N_6156);
or U9298 (N_9298,N_6881,N_7251);
and U9299 (N_9299,N_7430,N_7835);
and U9300 (N_9300,N_7842,N_7503);
nor U9301 (N_9301,N_7874,N_7033);
or U9302 (N_9302,N_6093,N_7097);
and U9303 (N_9303,N_7264,N_7861);
nor U9304 (N_9304,N_7211,N_6921);
nor U9305 (N_9305,N_7698,N_6241);
nor U9306 (N_9306,N_7959,N_6246);
or U9307 (N_9307,N_7577,N_7270);
xor U9308 (N_9308,N_7841,N_6880);
or U9309 (N_9309,N_7213,N_7135);
nand U9310 (N_9310,N_6282,N_7164);
nor U9311 (N_9311,N_6956,N_7977);
and U9312 (N_9312,N_6071,N_7449);
nor U9313 (N_9313,N_7460,N_6924);
and U9314 (N_9314,N_6921,N_7537);
and U9315 (N_9315,N_7462,N_7311);
nor U9316 (N_9316,N_6208,N_7880);
nor U9317 (N_9317,N_7630,N_7217);
and U9318 (N_9318,N_7576,N_7303);
xnor U9319 (N_9319,N_7455,N_6133);
xnor U9320 (N_9320,N_7721,N_7257);
and U9321 (N_9321,N_6546,N_7846);
xnor U9322 (N_9322,N_6036,N_6102);
nor U9323 (N_9323,N_6426,N_7355);
and U9324 (N_9324,N_6057,N_7471);
nand U9325 (N_9325,N_6097,N_6107);
or U9326 (N_9326,N_6033,N_6694);
and U9327 (N_9327,N_7193,N_6604);
nand U9328 (N_9328,N_6527,N_6406);
or U9329 (N_9329,N_7400,N_7276);
and U9330 (N_9330,N_7552,N_6580);
xnor U9331 (N_9331,N_6739,N_6082);
nor U9332 (N_9332,N_6308,N_6823);
xor U9333 (N_9333,N_7823,N_6692);
and U9334 (N_9334,N_6325,N_7299);
and U9335 (N_9335,N_6320,N_7997);
and U9336 (N_9336,N_6314,N_7634);
or U9337 (N_9337,N_6676,N_7562);
nor U9338 (N_9338,N_6359,N_6513);
nand U9339 (N_9339,N_6495,N_7623);
nor U9340 (N_9340,N_6812,N_7054);
or U9341 (N_9341,N_6201,N_7898);
nor U9342 (N_9342,N_7324,N_7964);
or U9343 (N_9343,N_7393,N_6984);
nor U9344 (N_9344,N_7021,N_7790);
or U9345 (N_9345,N_6394,N_6381);
nor U9346 (N_9346,N_6110,N_6710);
nand U9347 (N_9347,N_7024,N_6523);
nor U9348 (N_9348,N_7602,N_7576);
and U9349 (N_9349,N_6717,N_6521);
and U9350 (N_9350,N_6425,N_7424);
and U9351 (N_9351,N_6230,N_7038);
and U9352 (N_9352,N_6688,N_7984);
nor U9353 (N_9353,N_7581,N_7526);
xor U9354 (N_9354,N_6241,N_6820);
xor U9355 (N_9355,N_6556,N_7640);
xor U9356 (N_9356,N_6700,N_6029);
nor U9357 (N_9357,N_7981,N_7513);
and U9358 (N_9358,N_7144,N_6053);
nor U9359 (N_9359,N_6027,N_7396);
or U9360 (N_9360,N_7717,N_6817);
nand U9361 (N_9361,N_6042,N_6040);
xor U9362 (N_9362,N_7617,N_7376);
nand U9363 (N_9363,N_6998,N_7497);
nor U9364 (N_9364,N_6874,N_7447);
and U9365 (N_9365,N_6311,N_6555);
and U9366 (N_9366,N_6291,N_7685);
or U9367 (N_9367,N_6767,N_6603);
nand U9368 (N_9368,N_6964,N_7895);
and U9369 (N_9369,N_6976,N_6227);
nand U9370 (N_9370,N_6093,N_6490);
nand U9371 (N_9371,N_6731,N_6021);
nor U9372 (N_9372,N_7139,N_6373);
nor U9373 (N_9373,N_7185,N_6226);
or U9374 (N_9374,N_6482,N_7595);
nor U9375 (N_9375,N_6975,N_6265);
and U9376 (N_9376,N_6274,N_6170);
nor U9377 (N_9377,N_6096,N_6233);
or U9378 (N_9378,N_6819,N_7220);
and U9379 (N_9379,N_6038,N_7257);
nor U9380 (N_9380,N_6038,N_6165);
and U9381 (N_9381,N_6563,N_7384);
or U9382 (N_9382,N_7510,N_7251);
and U9383 (N_9383,N_7533,N_6489);
nor U9384 (N_9384,N_6146,N_7870);
nor U9385 (N_9385,N_7469,N_6060);
nand U9386 (N_9386,N_6947,N_7659);
nor U9387 (N_9387,N_7943,N_7882);
nor U9388 (N_9388,N_6136,N_7699);
and U9389 (N_9389,N_7241,N_6799);
xnor U9390 (N_9390,N_7754,N_6358);
nor U9391 (N_9391,N_6677,N_6717);
and U9392 (N_9392,N_7762,N_7293);
nor U9393 (N_9393,N_7237,N_6759);
or U9394 (N_9394,N_6411,N_6608);
or U9395 (N_9395,N_7274,N_6021);
or U9396 (N_9396,N_7883,N_6979);
and U9397 (N_9397,N_7583,N_7042);
nor U9398 (N_9398,N_7110,N_6903);
or U9399 (N_9399,N_6716,N_7515);
and U9400 (N_9400,N_7979,N_7508);
or U9401 (N_9401,N_7098,N_6274);
nand U9402 (N_9402,N_6343,N_7951);
and U9403 (N_9403,N_6386,N_6027);
and U9404 (N_9404,N_7253,N_7717);
nand U9405 (N_9405,N_6960,N_6867);
or U9406 (N_9406,N_7778,N_7089);
and U9407 (N_9407,N_6816,N_6793);
or U9408 (N_9408,N_7475,N_7271);
or U9409 (N_9409,N_7407,N_7286);
nor U9410 (N_9410,N_7031,N_7747);
or U9411 (N_9411,N_7544,N_7367);
nor U9412 (N_9412,N_6061,N_6682);
nor U9413 (N_9413,N_6517,N_7895);
nor U9414 (N_9414,N_7384,N_6464);
or U9415 (N_9415,N_6522,N_6901);
and U9416 (N_9416,N_7400,N_7110);
nor U9417 (N_9417,N_7136,N_6277);
or U9418 (N_9418,N_7798,N_7244);
nand U9419 (N_9419,N_7346,N_7395);
or U9420 (N_9420,N_6715,N_7832);
nand U9421 (N_9421,N_6578,N_6866);
or U9422 (N_9422,N_7780,N_6537);
nand U9423 (N_9423,N_7367,N_6067);
and U9424 (N_9424,N_6781,N_7171);
and U9425 (N_9425,N_7737,N_7169);
nor U9426 (N_9426,N_6534,N_7640);
and U9427 (N_9427,N_7020,N_6764);
nor U9428 (N_9428,N_7609,N_6121);
or U9429 (N_9429,N_6049,N_7797);
nand U9430 (N_9430,N_6829,N_7663);
nand U9431 (N_9431,N_7343,N_6074);
nand U9432 (N_9432,N_7711,N_6564);
and U9433 (N_9433,N_7197,N_7352);
nor U9434 (N_9434,N_7175,N_6322);
or U9435 (N_9435,N_7784,N_7725);
nor U9436 (N_9436,N_7193,N_6453);
nor U9437 (N_9437,N_7798,N_6940);
nand U9438 (N_9438,N_7018,N_6046);
and U9439 (N_9439,N_6184,N_6586);
nor U9440 (N_9440,N_6130,N_6010);
or U9441 (N_9441,N_6111,N_6104);
or U9442 (N_9442,N_7665,N_6659);
nor U9443 (N_9443,N_7099,N_7787);
or U9444 (N_9444,N_6966,N_6215);
nor U9445 (N_9445,N_7660,N_6478);
and U9446 (N_9446,N_7061,N_7399);
nand U9447 (N_9447,N_7925,N_7573);
nand U9448 (N_9448,N_6469,N_6034);
or U9449 (N_9449,N_7867,N_6064);
nand U9450 (N_9450,N_7463,N_6817);
and U9451 (N_9451,N_6507,N_7529);
nor U9452 (N_9452,N_7190,N_6094);
and U9453 (N_9453,N_6245,N_6006);
and U9454 (N_9454,N_7062,N_7859);
nand U9455 (N_9455,N_6414,N_6971);
and U9456 (N_9456,N_6689,N_7111);
nor U9457 (N_9457,N_7049,N_7298);
or U9458 (N_9458,N_6662,N_6693);
and U9459 (N_9459,N_7856,N_6109);
and U9460 (N_9460,N_6078,N_6040);
xnor U9461 (N_9461,N_6004,N_7997);
and U9462 (N_9462,N_7910,N_7141);
or U9463 (N_9463,N_7536,N_7793);
or U9464 (N_9464,N_7215,N_6505);
xnor U9465 (N_9465,N_6201,N_7777);
nand U9466 (N_9466,N_7779,N_7443);
nand U9467 (N_9467,N_7501,N_7992);
nor U9468 (N_9468,N_7412,N_6850);
nand U9469 (N_9469,N_6247,N_7095);
and U9470 (N_9470,N_7726,N_6723);
or U9471 (N_9471,N_7022,N_6031);
nor U9472 (N_9472,N_7054,N_7249);
nor U9473 (N_9473,N_6189,N_7180);
and U9474 (N_9474,N_7082,N_6483);
and U9475 (N_9475,N_6482,N_6766);
nand U9476 (N_9476,N_6573,N_6260);
or U9477 (N_9477,N_7686,N_7759);
and U9478 (N_9478,N_6258,N_7172);
and U9479 (N_9479,N_6836,N_6979);
nand U9480 (N_9480,N_6603,N_6244);
nor U9481 (N_9481,N_6169,N_7730);
or U9482 (N_9482,N_7460,N_7392);
or U9483 (N_9483,N_7875,N_7574);
nand U9484 (N_9484,N_6797,N_7008);
nor U9485 (N_9485,N_6466,N_7147);
nor U9486 (N_9486,N_6709,N_7685);
xnor U9487 (N_9487,N_7922,N_6047);
and U9488 (N_9488,N_6265,N_6897);
and U9489 (N_9489,N_7155,N_7557);
nand U9490 (N_9490,N_7680,N_7347);
or U9491 (N_9491,N_6055,N_6024);
nand U9492 (N_9492,N_7176,N_7287);
or U9493 (N_9493,N_7026,N_6603);
and U9494 (N_9494,N_7259,N_7908);
and U9495 (N_9495,N_7370,N_6882);
and U9496 (N_9496,N_7550,N_6947);
or U9497 (N_9497,N_6753,N_7830);
nor U9498 (N_9498,N_6549,N_7720);
nand U9499 (N_9499,N_7813,N_6025);
or U9500 (N_9500,N_6471,N_7819);
and U9501 (N_9501,N_7921,N_6260);
or U9502 (N_9502,N_6924,N_7922);
nor U9503 (N_9503,N_6951,N_6771);
xnor U9504 (N_9504,N_6684,N_7749);
nand U9505 (N_9505,N_6865,N_6014);
or U9506 (N_9506,N_7630,N_6311);
nand U9507 (N_9507,N_6513,N_7436);
nand U9508 (N_9508,N_6471,N_6785);
nor U9509 (N_9509,N_6288,N_6554);
and U9510 (N_9510,N_6733,N_7361);
nand U9511 (N_9511,N_6206,N_7103);
and U9512 (N_9512,N_7307,N_6975);
or U9513 (N_9513,N_7324,N_6533);
and U9514 (N_9514,N_7043,N_7071);
or U9515 (N_9515,N_6324,N_7397);
and U9516 (N_9516,N_7225,N_7967);
nor U9517 (N_9517,N_6980,N_6858);
nor U9518 (N_9518,N_7945,N_6106);
or U9519 (N_9519,N_7745,N_7362);
and U9520 (N_9520,N_6089,N_6026);
or U9521 (N_9521,N_6189,N_7526);
nor U9522 (N_9522,N_7595,N_7067);
and U9523 (N_9523,N_6938,N_7454);
and U9524 (N_9524,N_6274,N_6035);
or U9525 (N_9525,N_7800,N_6145);
xnor U9526 (N_9526,N_7682,N_6857);
nand U9527 (N_9527,N_6920,N_7211);
nor U9528 (N_9528,N_7429,N_7280);
nand U9529 (N_9529,N_7038,N_7240);
and U9530 (N_9530,N_6174,N_6139);
or U9531 (N_9531,N_7251,N_7726);
and U9532 (N_9532,N_6460,N_7971);
nand U9533 (N_9533,N_7102,N_6412);
nor U9534 (N_9534,N_7435,N_7007);
and U9535 (N_9535,N_6378,N_7010);
nor U9536 (N_9536,N_6176,N_7662);
nor U9537 (N_9537,N_7158,N_7908);
xnor U9538 (N_9538,N_7787,N_7449);
nand U9539 (N_9539,N_6284,N_7197);
nor U9540 (N_9540,N_6661,N_6662);
nand U9541 (N_9541,N_6576,N_6271);
and U9542 (N_9542,N_7458,N_6608);
or U9543 (N_9543,N_7041,N_6352);
nor U9544 (N_9544,N_7759,N_7693);
nand U9545 (N_9545,N_7637,N_6547);
xnor U9546 (N_9546,N_6692,N_6595);
or U9547 (N_9547,N_7167,N_6523);
or U9548 (N_9548,N_6692,N_7733);
nand U9549 (N_9549,N_6870,N_7631);
or U9550 (N_9550,N_7200,N_7256);
and U9551 (N_9551,N_6366,N_7993);
or U9552 (N_9552,N_6002,N_6330);
nor U9553 (N_9553,N_7228,N_7998);
nand U9554 (N_9554,N_6761,N_6239);
xnor U9555 (N_9555,N_6926,N_7312);
nand U9556 (N_9556,N_7731,N_6438);
nor U9557 (N_9557,N_6032,N_6664);
xnor U9558 (N_9558,N_7649,N_7605);
and U9559 (N_9559,N_7965,N_6683);
or U9560 (N_9560,N_7719,N_7198);
and U9561 (N_9561,N_7578,N_6398);
nor U9562 (N_9562,N_6326,N_7273);
or U9563 (N_9563,N_7448,N_7689);
nand U9564 (N_9564,N_7634,N_7576);
or U9565 (N_9565,N_7535,N_6894);
and U9566 (N_9566,N_7054,N_7034);
or U9567 (N_9567,N_7708,N_7396);
or U9568 (N_9568,N_6752,N_7144);
nand U9569 (N_9569,N_6566,N_6121);
nor U9570 (N_9570,N_7682,N_6393);
and U9571 (N_9571,N_6216,N_6635);
nor U9572 (N_9572,N_7481,N_7245);
nand U9573 (N_9573,N_6867,N_6680);
nand U9574 (N_9574,N_6165,N_7624);
xor U9575 (N_9575,N_6467,N_7430);
nor U9576 (N_9576,N_7423,N_6506);
or U9577 (N_9577,N_6459,N_7090);
nand U9578 (N_9578,N_6473,N_7262);
nand U9579 (N_9579,N_7471,N_7192);
nor U9580 (N_9580,N_6741,N_7729);
nand U9581 (N_9581,N_7542,N_6369);
nor U9582 (N_9582,N_6797,N_7211);
nor U9583 (N_9583,N_7542,N_7685);
and U9584 (N_9584,N_7374,N_6501);
nor U9585 (N_9585,N_6705,N_6819);
nor U9586 (N_9586,N_7220,N_7583);
and U9587 (N_9587,N_7295,N_7395);
xnor U9588 (N_9588,N_7715,N_7328);
or U9589 (N_9589,N_6135,N_6592);
nand U9590 (N_9590,N_7756,N_7814);
xor U9591 (N_9591,N_6876,N_7297);
or U9592 (N_9592,N_7757,N_7007);
or U9593 (N_9593,N_7590,N_6260);
and U9594 (N_9594,N_7596,N_7000);
nand U9595 (N_9595,N_6514,N_6190);
and U9596 (N_9596,N_6311,N_7986);
nand U9597 (N_9597,N_6424,N_7180);
nor U9598 (N_9598,N_7205,N_6711);
nand U9599 (N_9599,N_6743,N_7021);
xor U9600 (N_9600,N_6875,N_6352);
and U9601 (N_9601,N_6389,N_6395);
nand U9602 (N_9602,N_7543,N_6109);
and U9603 (N_9603,N_7885,N_7569);
nor U9604 (N_9604,N_7108,N_7813);
or U9605 (N_9605,N_7276,N_6723);
and U9606 (N_9606,N_7452,N_6620);
and U9607 (N_9607,N_7352,N_6192);
nor U9608 (N_9608,N_6676,N_6756);
nor U9609 (N_9609,N_7596,N_6240);
or U9610 (N_9610,N_6548,N_7338);
and U9611 (N_9611,N_7519,N_6359);
nor U9612 (N_9612,N_7081,N_6304);
nand U9613 (N_9613,N_6553,N_7845);
and U9614 (N_9614,N_7619,N_6082);
or U9615 (N_9615,N_7967,N_6485);
or U9616 (N_9616,N_7492,N_6083);
or U9617 (N_9617,N_7916,N_7537);
and U9618 (N_9618,N_7675,N_6826);
or U9619 (N_9619,N_7513,N_7476);
nand U9620 (N_9620,N_7666,N_7950);
nor U9621 (N_9621,N_7199,N_6463);
xor U9622 (N_9622,N_6721,N_6741);
nor U9623 (N_9623,N_6677,N_6088);
nor U9624 (N_9624,N_6797,N_7001);
and U9625 (N_9625,N_7322,N_7593);
nand U9626 (N_9626,N_7446,N_6358);
nand U9627 (N_9627,N_7077,N_6794);
or U9628 (N_9628,N_7168,N_6444);
or U9629 (N_9629,N_7996,N_6625);
nand U9630 (N_9630,N_7780,N_7030);
or U9631 (N_9631,N_6615,N_6213);
and U9632 (N_9632,N_7199,N_6167);
nand U9633 (N_9633,N_6977,N_6278);
and U9634 (N_9634,N_7063,N_7703);
and U9635 (N_9635,N_7379,N_7979);
or U9636 (N_9636,N_7979,N_7352);
and U9637 (N_9637,N_7589,N_6250);
nand U9638 (N_9638,N_6400,N_7591);
nand U9639 (N_9639,N_7109,N_6423);
or U9640 (N_9640,N_7075,N_7928);
nor U9641 (N_9641,N_7697,N_7760);
nand U9642 (N_9642,N_7536,N_7546);
nor U9643 (N_9643,N_6870,N_7708);
or U9644 (N_9644,N_7608,N_7568);
nor U9645 (N_9645,N_6152,N_6814);
or U9646 (N_9646,N_7788,N_7953);
and U9647 (N_9647,N_7017,N_6284);
nand U9648 (N_9648,N_6679,N_6029);
or U9649 (N_9649,N_7710,N_6918);
nor U9650 (N_9650,N_7471,N_6710);
or U9651 (N_9651,N_7923,N_7563);
nor U9652 (N_9652,N_7086,N_7355);
and U9653 (N_9653,N_7745,N_7561);
and U9654 (N_9654,N_6851,N_7779);
and U9655 (N_9655,N_7797,N_6891);
xnor U9656 (N_9656,N_6195,N_6269);
and U9657 (N_9657,N_7272,N_6602);
or U9658 (N_9658,N_7882,N_6792);
nor U9659 (N_9659,N_6041,N_6689);
and U9660 (N_9660,N_7235,N_7393);
nor U9661 (N_9661,N_6908,N_6663);
or U9662 (N_9662,N_6203,N_7080);
nor U9663 (N_9663,N_7911,N_7280);
nand U9664 (N_9664,N_6129,N_7245);
or U9665 (N_9665,N_7652,N_7242);
xnor U9666 (N_9666,N_7210,N_6679);
xnor U9667 (N_9667,N_7951,N_7110);
nor U9668 (N_9668,N_6173,N_7659);
nor U9669 (N_9669,N_7573,N_7806);
nor U9670 (N_9670,N_7870,N_7655);
nor U9671 (N_9671,N_6171,N_7631);
nor U9672 (N_9672,N_7464,N_6622);
or U9673 (N_9673,N_7430,N_6487);
and U9674 (N_9674,N_6218,N_6919);
nand U9675 (N_9675,N_7687,N_7294);
or U9676 (N_9676,N_7582,N_6037);
or U9677 (N_9677,N_7707,N_6468);
xnor U9678 (N_9678,N_6412,N_6650);
xor U9679 (N_9679,N_7174,N_6507);
nor U9680 (N_9680,N_7170,N_7538);
or U9681 (N_9681,N_6439,N_7459);
xnor U9682 (N_9682,N_7214,N_7021);
nand U9683 (N_9683,N_6139,N_6747);
nand U9684 (N_9684,N_6398,N_7133);
nand U9685 (N_9685,N_6601,N_7359);
xor U9686 (N_9686,N_7550,N_7589);
nand U9687 (N_9687,N_7792,N_6237);
or U9688 (N_9688,N_7775,N_7844);
or U9689 (N_9689,N_7530,N_6459);
nor U9690 (N_9690,N_6688,N_7906);
and U9691 (N_9691,N_6457,N_6945);
nor U9692 (N_9692,N_6128,N_7290);
nor U9693 (N_9693,N_6932,N_6236);
and U9694 (N_9694,N_7237,N_6636);
nor U9695 (N_9695,N_6545,N_7119);
and U9696 (N_9696,N_6908,N_7589);
nand U9697 (N_9697,N_6303,N_6675);
and U9698 (N_9698,N_7198,N_6939);
or U9699 (N_9699,N_6275,N_7153);
xor U9700 (N_9700,N_7844,N_6358);
and U9701 (N_9701,N_6079,N_7274);
nand U9702 (N_9702,N_6106,N_7658);
and U9703 (N_9703,N_6443,N_6955);
nor U9704 (N_9704,N_7680,N_7348);
and U9705 (N_9705,N_6755,N_6394);
nor U9706 (N_9706,N_6895,N_7971);
nor U9707 (N_9707,N_6175,N_6279);
or U9708 (N_9708,N_6569,N_7947);
nand U9709 (N_9709,N_6599,N_7026);
or U9710 (N_9710,N_7151,N_7771);
nor U9711 (N_9711,N_6250,N_7749);
or U9712 (N_9712,N_7153,N_7288);
nand U9713 (N_9713,N_7217,N_7291);
nand U9714 (N_9714,N_6370,N_7035);
and U9715 (N_9715,N_6947,N_6958);
nor U9716 (N_9716,N_7211,N_6942);
nand U9717 (N_9717,N_6183,N_7763);
or U9718 (N_9718,N_6336,N_7705);
or U9719 (N_9719,N_6794,N_7732);
or U9720 (N_9720,N_7367,N_7017);
or U9721 (N_9721,N_6775,N_7275);
nor U9722 (N_9722,N_6671,N_6448);
and U9723 (N_9723,N_7204,N_6491);
nand U9724 (N_9724,N_7761,N_7145);
nor U9725 (N_9725,N_7024,N_7587);
nand U9726 (N_9726,N_7651,N_7636);
nor U9727 (N_9727,N_7747,N_6894);
nor U9728 (N_9728,N_7970,N_7639);
nand U9729 (N_9729,N_7751,N_7575);
and U9730 (N_9730,N_7738,N_6978);
nor U9731 (N_9731,N_7109,N_6178);
nor U9732 (N_9732,N_7062,N_7586);
xor U9733 (N_9733,N_6934,N_7944);
and U9734 (N_9734,N_7769,N_7336);
nor U9735 (N_9735,N_7146,N_6262);
or U9736 (N_9736,N_7841,N_7092);
xor U9737 (N_9737,N_7286,N_7390);
nor U9738 (N_9738,N_6771,N_7470);
nor U9739 (N_9739,N_6504,N_7876);
or U9740 (N_9740,N_7675,N_6312);
nand U9741 (N_9741,N_7063,N_6687);
nand U9742 (N_9742,N_7139,N_7680);
and U9743 (N_9743,N_7351,N_6323);
and U9744 (N_9744,N_7211,N_7054);
and U9745 (N_9745,N_6833,N_6135);
or U9746 (N_9746,N_6364,N_6146);
and U9747 (N_9747,N_7645,N_6436);
nand U9748 (N_9748,N_7551,N_6446);
nand U9749 (N_9749,N_6751,N_6344);
and U9750 (N_9750,N_7170,N_6306);
or U9751 (N_9751,N_6721,N_6310);
nor U9752 (N_9752,N_7460,N_7293);
nand U9753 (N_9753,N_6308,N_6168);
nor U9754 (N_9754,N_7638,N_7379);
or U9755 (N_9755,N_7710,N_7056);
or U9756 (N_9756,N_6729,N_7677);
nor U9757 (N_9757,N_6582,N_7578);
nor U9758 (N_9758,N_7058,N_6066);
and U9759 (N_9759,N_6676,N_6126);
nand U9760 (N_9760,N_7050,N_7855);
nand U9761 (N_9761,N_7136,N_6227);
nor U9762 (N_9762,N_7363,N_7876);
xor U9763 (N_9763,N_7515,N_7374);
nand U9764 (N_9764,N_7245,N_7364);
nor U9765 (N_9765,N_6823,N_7329);
or U9766 (N_9766,N_6441,N_7159);
xnor U9767 (N_9767,N_7472,N_6537);
and U9768 (N_9768,N_6482,N_6823);
and U9769 (N_9769,N_6704,N_7620);
nand U9770 (N_9770,N_7373,N_7414);
or U9771 (N_9771,N_7145,N_6929);
and U9772 (N_9772,N_6464,N_6501);
and U9773 (N_9773,N_6655,N_7999);
and U9774 (N_9774,N_6305,N_6850);
nand U9775 (N_9775,N_7416,N_7240);
or U9776 (N_9776,N_7473,N_6367);
or U9777 (N_9777,N_6836,N_7235);
or U9778 (N_9778,N_6457,N_6037);
nand U9779 (N_9779,N_6800,N_7562);
or U9780 (N_9780,N_6978,N_7922);
or U9781 (N_9781,N_6189,N_7405);
xor U9782 (N_9782,N_6563,N_7875);
nor U9783 (N_9783,N_7444,N_6963);
xor U9784 (N_9784,N_7705,N_6564);
and U9785 (N_9785,N_6657,N_7869);
nand U9786 (N_9786,N_7484,N_6833);
xor U9787 (N_9787,N_7714,N_6143);
and U9788 (N_9788,N_7367,N_7460);
or U9789 (N_9789,N_6742,N_6103);
nor U9790 (N_9790,N_7826,N_7351);
nor U9791 (N_9791,N_6697,N_7868);
and U9792 (N_9792,N_7618,N_6835);
or U9793 (N_9793,N_6220,N_7432);
or U9794 (N_9794,N_6159,N_7776);
nor U9795 (N_9795,N_6387,N_6496);
or U9796 (N_9796,N_6079,N_6827);
and U9797 (N_9797,N_6376,N_6103);
or U9798 (N_9798,N_7312,N_7275);
nand U9799 (N_9799,N_6191,N_7330);
nor U9800 (N_9800,N_6877,N_7240);
nand U9801 (N_9801,N_6788,N_7188);
nor U9802 (N_9802,N_7079,N_6236);
and U9803 (N_9803,N_6187,N_7734);
or U9804 (N_9804,N_6678,N_6198);
and U9805 (N_9805,N_7367,N_6615);
or U9806 (N_9806,N_7147,N_6225);
or U9807 (N_9807,N_7055,N_6402);
nand U9808 (N_9808,N_6182,N_6062);
nor U9809 (N_9809,N_6549,N_6666);
nand U9810 (N_9810,N_7448,N_7186);
nand U9811 (N_9811,N_6495,N_6328);
nand U9812 (N_9812,N_6753,N_6554);
and U9813 (N_9813,N_7161,N_6431);
nor U9814 (N_9814,N_6088,N_6769);
and U9815 (N_9815,N_6585,N_6291);
nand U9816 (N_9816,N_7812,N_7005);
and U9817 (N_9817,N_7424,N_6854);
and U9818 (N_9818,N_7119,N_6052);
xnor U9819 (N_9819,N_7561,N_6473);
nand U9820 (N_9820,N_6475,N_7702);
nand U9821 (N_9821,N_7295,N_7792);
or U9822 (N_9822,N_7642,N_6466);
nand U9823 (N_9823,N_7549,N_6828);
nand U9824 (N_9824,N_7355,N_7722);
and U9825 (N_9825,N_7371,N_7685);
nand U9826 (N_9826,N_7762,N_7577);
or U9827 (N_9827,N_7020,N_7011);
xnor U9828 (N_9828,N_6536,N_6787);
nand U9829 (N_9829,N_7792,N_7427);
and U9830 (N_9830,N_6987,N_7166);
nand U9831 (N_9831,N_7262,N_7565);
and U9832 (N_9832,N_6395,N_6308);
nor U9833 (N_9833,N_7925,N_6022);
nand U9834 (N_9834,N_7349,N_7793);
nor U9835 (N_9835,N_7620,N_7501);
nor U9836 (N_9836,N_7099,N_6505);
and U9837 (N_9837,N_6968,N_6242);
nor U9838 (N_9838,N_6548,N_6583);
nor U9839 (N_9839,N_6102,N_7082);
xnor U9840 (N_9840,N_7571,N_7278);
nor U9841 (N_9841,N_7090,N_7269);
or U9842 (N_9842,N_6695,N_7357);
and U9843 (N_9843,N_6548,N_6194);
or U9844 (N_9844,N_7067,N_7809);
and U9845 (N_9845,N_7475,N_6972);
and U9846 (N_9846,N_6118,N_7496);
or U9847 (N_9847,N_6361,N_7065);
nand U9848 (N_9848,N_6843,N_6143);
or U9849 (N_9849,N_7428,N_7202);
and U9850 (N_9850,N_7355,N_6349);
or U9851 (N_9851,N_7836,N_6311);
and U9852 (N_9852,N_7724,N_7904);
nand U9853 (N_9853,N_6385,N_7880);
nor U9854 (N_9854,N_6077,N_7770);
nor U9855 (N_9855,N_7470,N_7133);
nand U9856 (N_9856,N_7669,N_6736);
and U9857 (N_9857,N_6355,N_6295);
and U9858 (N_9858,N_6801,N_7215);
or U9859 (N_9859,N_7015,N_7690);
nor U9860 (N_9860,N_7276,N_6876);
nand U9861 (N_9861,N_6572,N_7041);
or U9862 (N_9862,N_7553,N_7435);
nand U9863 (N_9863,N_6857,N_7730);
nand U9864 (N_9864,N_6951,N_6367);
nand U9865 (N_9865,N_7441,N_7230);
or U9866 (N_9866,N_7512,N_7986);
nand U9867 (N_9867,N_6171,N_6904);
nor U9868 (N_9868,N_6182,N_7397);
nor U9869 (N_9869,N_6301,N_6928);
nor U9870 (N_9870,N_7590,N_7704);
nand U9871 (N_9871,N_7425,N_7723);
nor U9872 (N_9872,N_6099,N_6963);
nand U9873 (N_9873,N_7888,N_6345);
nand U9874 (N_9874,N_6729,N_7252);
nand U9875 (N_9875,N_7029,N_6644);
nor U9876 (N_9876,N_7551,N_7841);
nor U9877 (N_9877,N_6248,N_7032);
xnor U9878 (N_9878,N_6765,N_7059);
nor U9879 (N_9879,N_7209,N_6130);
nand U9880 (N_9880,N_6987,N_7691);
nand U9881 (N_9881,N_7921,N_7445);
nand U9882 (N_9882,N_6340,N_7878);
nor U9883 (N_9883,N_7941,N_7663);
or U9884 (N_9884,N_7529,N_7659);
xnor U9885 (N_9885,N_7112,N_7949);
or U9886 (N_9886,N_7999,N_7011);
nor U9887 (N_9887,N_6926,N_7113);
and U9888 (N_9888,N_7064,N_6244);
or U9889 (N_9889,N_6988,N_6049);
or U9890 (N_9890,N_6449,N_7448);
and U9891 (N_9891,N_7631,N_6983);
or U9892 (N_9892,N_6963,N_6672);
or U9893 (N_9893,N_6235,N_6185);
nand U9894 (N_9894,N_6089,N_6967);
or U9895 (N_9895,N_7435,N_7269);
or U9896 (N_9896,N_7982,N_7227);
or U9897 (N_9897,N_6668,N_6130);
nor U9898 (N_9898,N_7257,N_6998);
nor U9899 (N_9899,N_6830,N_6555);
xnor U9900 (N_9900,N_6991,N_7268);
nor U9901 (N_9901,N_7059,N_7365);
nand U9902 (N_9902,N_7857,N_6300);
or U9903 (N_9903,N_6760,N_6758);
nor U9904 (N_9904,N_7626,N_7725);
and U9905 (N_9905,N_6841,N_6126);
or U9906 (N_9906,N_7819,N_6954);
nand U9907 (N_9907,N_7830,N_6628);
xnor U9908 (N_9908,N_7573,N_7881);
nand U9909 (N_9909,N_6574,N_7265);
nor U9910 (N_9910,N_7262,N_6487);
nor U9911 (N_9911,N_6687,N_7090);
or U9912 (N_9912,N_7895,N_7582);
nor U9913 (N_9913,N_7013,N_7087);
nor U9914 (N_9914,N_6945,N_6396);
nor U9915 (N_9915,N_7060,N_6887);
nand U9916 (N_9916,N_7858,N_6802);
nand U9917 (N_9917,N_7531,N_6329);
nand U9918 (N_9918,N_7956,N_7318);
and U9919 (N_9919,N_7907,N_6263);
and U9920 (N_9920,N_6648,N_7437);
and U9921 (N_9921,N_7348,N_6631);
nand U9922 (N_9922,N_6464,N_7661);
or U9923 (N_9923,N_7757,N_7718);
and U9924 (N_9924,N_6517,N_7185);
and U9925 (N_9925,N_7464,N_7564);
and U9926 (N_9926,N_6763,N_7008);
nand U9927 (N_9927,N_6402,N_6152);
xnor U9928 (N_9928,N_7539,N_7467);
or U9929 (N_9929,N_6231,N_7327);
nand U9930 (N_9930,N_7622,N_6686);
xnor U9931 (N_9931,N_7286,N_6921);
and U9932 (N_9932,N_6219,N_6813);
and U9933 (N_9933,N_6733,N_6622);
nand U9934 (N_9934,N_7190,N_7336);
nand U9935 (N_9935,N_6496,N_6317);
nand U9936 (N_9936,N_6540,N_6911);
nor U9937 (N_9937,N_6839,N_6171);
nor U9938 (N_9938,N_7878,N_6328);
nor U9939 (N_9939,N_6867,N_6932);
nand U9940 (N_9940,N_7035,N_7030);
or U9941 (N_9941,N_7760,N_6179);
and U9942 (N_9942,N_7383,N_7320);
nor U9943 (N_9943,N_6177,N_7230);
and U9944 (N_9944,N_6414,N_7468);
or U9945 (N_9945,N_6960,N_7271);
nor U9946 (N_9946,N_7747,N_6648);
and U9947 (N_9947,N_6029,N_7615);
and U9948 (N_9948,N_6420,N_7607);
xor U9949 (N_9949,N_7365,N_7828);
nor U9950 (N_9950,N_6422,N_7571);
xor U9951 (N_9951,N_7594,N_6120);
xnor U9952 (N_9952,N_7469,N_7347);
nand U9953 (N_9953,N_7666,N_6879);
or U9954 (N_9954,N_6224,N_7502);
or U9955 (N_9955,N_7183,N_7979);
and U9956 (N_9956,N_7212,N_7766);
and U9957 (N_9957,N_6039,N_6398);
nor U9958 (N_9958,N_7120,N_7191);
and U9959 (N_9959,N_7424,N_7964);
or U9960 (N_9960,N_7507,N_6767);
or U9961 (N_9961,N_7875,N_7140);
and U9962 (N_9962,N_6698,N_7561);
nor U9963 (N_9963,N_6338,N_6638);
nand U9964 (N_9964,N_7855,N_6262);
nand U9965 (N_9965,N_7791,N_7213);
xnor U9966 (N_9966,N_7087,N_7683);
or U9967 (N_9967,N_7303,N_6315);
nand U9968 (N_9968,N_7528,N_6157);
nor U9969 (N_9969,N_6567,N_7692);
and U9970 (N_9970,N_7131,N_6201);
xor U9971 (N_9971,N_7705,N_7240);
nand U9972 (N_9972,N_7277,N_7552);
and U9973 (N_9973,N_7602,N_6007);
nor U9974 (N_9974,N_7880,N_6051);
and U9975 (N_9975,N_6998,N_6828);
xor U9976 (N_9976,N_6467,N_6263);
xnor U9977 (N_9977,N_7906,N_7724);
and U9978 (N_9978,N_7638,N_7316);
and U9979 (N_9979,N_6689,N_7362);
nor U9980 (N_9980,N_7494,N_7181);
nand U9981 (N_9981,N_7340,N_6416);
nor U9982 (N_9982,N_7978,N_7545);
nor U9983 (N_9983,N_6771,N_6189);
or U9984 (N_9984,N_7404,N_7970);
xnor U9985 (N_9985,N_6501,N_7120);
nor U9986 (N_9986,N_6591,N_7676);
nand U9987 (N_9987,N_6876,N_6111);
or U9988 (N_9988,N_6290,N_6834);
and U9989 (N_9989,N_6887,N_6905);
and U9990 (N_9990,N_6868,N_6870);
nand U9991 (N_9991,N_6528,N_7531);
or U9992 (N_9992,N_7625,N_7847);
or U9993 (N_9993,N_6824,N_7976);
nand U9994 (N_9994,N_6376,N_7701);
nor U9995 (N_9995,N_7308,N_6573);
and U9996 (N_9996,N_7046,N_7234);
or U9997 (N_9997,N_7024,N_7931);
xor U9998 (N_9998,N_6746,N_6333);
nor U9999 (N_9999,N_6778,N_6926);
or U10000 (N_10000,N_8568,N_8847);
and U10001 (N_10001,N_8199,N_8581);
or U10002 (N_10002,N_9628,N_9732);
and U10003 (N_10003,N_8660,N_9170);
and U10004 (N_10004,N_8153,N_9115);
or U10005 (N_10005,N_9895,N_9190);
xnor U10006 (N_10006,N_8948,N_8493);
and U10007 (N_10007,N_9045,N_9702);
nor U10008 (N_10008,N_9405,N_9990);
or U10009 (N_10009,N_9695,N_9878);
and U10010 (N_10010,N_9159,N_8713);
nor U10011 (N_10011,N_8030,N_8941);
nand U10012 (N_10012,N_9266,N_9243);
or U10013 (N_10013,N_8132,N_8538);
and U10014 (N_10014,N_9198,N_8155);
nor U10015 (N_10015,N_8088,N_8247);
nand U10016 (N_10016,N_9263,N_8221);
or U10017 (N_10017,N_8683,N_8490);
xor U10018 (N_10018,N_8913,N_8016);
and U10019 (N_10019,N_9284,N_8354);
and U10020 (N_10020,N_8494,N_8257);
and U10021 (N_10021,N_9697,N_9731);
and U10022 (N_10022,N_8682,N_9656);
or U10023 (N_10023,N_8436,N_8933);
or U10024 (N_10024,N_9829,N_9722);
or U10025 (N_10025,N_9467,N_8842);
and U10026 (N_10026,N_8350,N_8495);
nand U10027 (N_10027,N_8499,N_8266);
xnor U10028 (N_10028,N_9674,N_9298);
and U10029 (N_10029,N_9452,N_9007);
xnor U10030 (N_10030,N_8073,N_9772);
nand U10031 (N_10031,N_8277,N_8053);
nand U10032 (N_10032,N_8236,N_8512);
or U10033 (N_10033,N_8105,N_8458);
nor U10034 (N_10034,N_8498,N_8692);
and U10035 (N_10035,N_9804,N_8622);
nor U10036 (N_10036,N_9141,N_8849);
nand U10037 (N_10037,N_8846,N_9589);
and U10038 (N_10038,N_9939,N_9093);
nor U10039 (N_10039,N_8628,N_8218);
nor U10040 (N_10040,N_9853,N_9867);
and U10041 (N_10041,N_8644,N_9565);
or U10042 (N_10042,N_9180,N_8778);
and U10043 (N_10043,N_8852,N_9124);
and U10044 (N_10044,N_8742,N_8533);
and U10045 (N_10045,N_9634,N_9175);
and U10046 (N_10046,N_9071,N_8601);
and U10047 (N_10047,N_8427,N_8780);
nor U10048 (N_10048,N_9142,N_9983);
or U10049 (N_10049,N_9610,N_9578);
or U10050 (N_10050,N_8051,N_9363);
nor U10051 (N_10051,N_9670,N_9640);
and U10052 (N_10052,N_9612,N_8511);
and U10053 (N_10053,N_9929,N_8025);
xor U10054 (N_10054,N_9129,N_9967);
and U10055 (N_10055,N_8796,N_9718);
nand U10056 (N_10056,N_8641,N_8484);
and U10057 (N_10057,N_8187,N_8943);
and U10058 (N_10058,N_8888,N_8031);
and U10059 (N_10059,N_8974,N_8283);
or U10060 (N_10060,N_9104,N_9861);
xor U10061 (N_10061,N_9092,N_9993);
xnor U10062 (N_10062,N_9328,N_9451);
nand U10063 (N_10063,N_9537,N_9655);
nor U10064 (N_10064,N_9755,N_8930);
or U10065 (N_10065,N_9027,N_8067);
nor U10066 (N_10066,N_8824,N_9608);
nor U10067 (N_10067,N_9036,N_9133);
and U10068 (N_10068,N_8977,N_9176);
or U10069 (N_10069,N_9669,N_9905);
nand U10070 (N_10070,N_8034,N_9766);
nand U10071 (N_10071,N_9040,N_8906);
xnor U10072 (N_10072,N_9552,N_9013);
nand U10073 (N_10073,N_9316,N_8927);
nand U10074 (N_10074,N_9339,N_9843);
or U10075 (N_10075,N_8563,N_8021);
or U10076 (N_10076,N_9283,N_9020);
nor U10077 (N_10077,N_8275,N_8989);
nor U10078 (N_10078,N_8522,N_8612);
nand U10079 (N_10079,N_8551,N_9618);
nand U10080 (N_10080,N_8246,N_8839);
nor U10081 (N_10081,N_8673,N_9764);
or U10082 (N_10082,N_9106,N_9423);
or U10083 (N_10083,N_8315,N_8599);
nand U10084 (N_10084,N_9816,N_9495);
xor U10085 (N_10085,N_9560,N_9987);
and U10086 (N_10086,N_9728,N_9430);
nand U10087 (N_10087,N_9836,N_9218);
nor U10088 (N_10088,N_8773,N_9822);
or U10089 (N_10089,N_8988,N_8443);
nand U10090 (N_10090,N_9418,N_8777);
and U10091 (N_10091,N_9450,N_9672);
or U10092 (N_10092,N_8461,N_8997);
nand U10093 (N_10093,N_9401,N_9951);
and U10094 (N_10094,N_9579,N_9077);
nand U10095 (N_10095,N_9315,N_9973);
and U10096 (N_10096,N_8099,N_9681);
or U10097 (N_10097,N_8864,N_9114);
and U10098 (N_10098,N_8899,N_9015);
and U10099 (N_10099,N_8419,N_8667);
nor U10100 (N_10100,N_8543,N_9546);
and U10101 (N_10101,N_9594,N_8194);
nand U10102 (N_10102,N_8395,N_9111);
nor U10103 (N_10103,N_9089,N_8929);
and U10104 (N_10104,N_9548,N_9684);
nand U10105 (N_10105,N_9394,N_8691);
nor U10106 (N_10106,N_8619,N_8144);
xnor U10107 (N_10107,N_9699,N_8302);
nand U10108 (N_10108,N_8148,N_9748);
nor U10109 (N_10109,N_9392,N_8002);
xnor U10110 (N_10110,N_8135,N_8120);
and U10111 (N_10111,N_9140,N_8784);
and U10112 (N_10112,N_9868,N_8642);
or U10113 (N_10113,N_8862,N_9158);
or U10114 (N_10114,N_8103,N_8009);
nor U10115 (N_10115,N_9319,N_9821);
nor U10116 (N_10116,N_9883,N_8771);
nand U10117 (N_10117,N_9269,N_9700);
and U10118 (N_10118,N_8217,N_8195);
nor U10119 (N_10119,N_9194,N_8500);
nor U10120 (N_10120,N_9119,N_9519);
nand U10121 (N_10121,N_8071,N_8985);
nand U10122 (N_10122,N_8014,N_8529);
and U10123 (N_10123,N_8727,N_8333);
nand U10124 (N_10124,N_9241,N_8424);
xor U10125 (N_10125,N_9500,N_9245);
nand U10126 (N_10126,N_8238,N_8441);
nand U10127 (N_10127,N_8129,N_8542);
and U10128 (N_10128,N_9481,N_8739);
nand U10129 (N_10129,N_9889,N_9955);
and U10130 (N_10130,N_8373,N_9833);
nor U10131 (N_10131,N_8478,N_8222);
xor U10132 (N_10132,N_9979,N_9149);
nor U10133 (N_10133,N_9614,N_9652);
nand U10134 (N_10134,N_8553,N_9910);
or U10135 (N_10135,N_8624,N_9370);
or U10136 (N_10136,N_8305,N_8074);
or U10137 (N_10137,N_8621,N_9575);
or U10138 (N_10138,N_9862,N_8766);
nor U10139 (N_10139,N_8335,N_9447);
xor U10140 (N_10140,N_9323,N_8104);
xor U10141 (N_10141,N_8794,N_9953);
nor U10142 (N_10142,N_9908,N_8184);
nor U10143 (N_10143,N_8801,N_9812);
nor U10144 (N_10144,N_8806,N_9424);
nor U10145 (N_10145,N_9116,N_8385);
xor U10146 (N_10146,N_9580,N_8935);
nor U10147 (N_10147,N_8240,N_8598);
xor U10148 (N_10148,N_9120,N_8370);
and U10149 (N_10149,N_8361,N_8161);
nor U10150 (N_10150,N_8438,N_8274);
nor U10151 (N_10151,N_8003,N_9597);
and U10152 (N_10152,N_9417,N_9557);
nor U10153 (N_10153,N_8804,N_8168);
nor U10154 (N_10154,N_8202,N_8027);
or U10155 (N_10155,N_8420,N_8557);
nor U10156 (N_10156,N_9980,N_9576);
and U10157 (N_10157,N_8853,N_8750);
and U10158 (N_10158,N_9056,N_8109);
or U10159 (N_10159,N_8625,N_9280);
or U10160 (N_10160,N_8540,N_8059);
nand U10161 (N_10161,N_9113,N_9123);
and U10162 (N_10162,N_8911,N_9039);
nand U10163 (N_10163,N_9033,N_9872);
xor U10164 (N_10164,N_9130,N_8431);
nand U10165 (N_10165,N_8376,N_9353);
and U10166 (N_10166,N_8799,N_9617);
or U10167 (N_10167,N_9105,N_9765);
xnor U10168 (N_10168,N_9288,N_9625);
nor U10169 (N_10169,N_8907,N_8102);
or U10170 (N_10170,N_8303,N_8614);
nor U10171 (N_10171,N_9197,N_9223);
nand U10172 (N_10172,N_9247,N_9646);
and U10173 (N_10173,N_8939,N_9923);
nand U10174 (N_10174,N_9227,N_9879);
xor U10175 (N_10175,N_9305,N_9870);
or U10176 (N_10176,N_8355,N_8092);
or U10177 (N_10177,N_9312,N_8632);
or U10178 (N_10178,N_9512,N_8825);
or U10179 (N_10179,N_9402,N_9382);
nor U10180 (N_10180,N_8158,N_8487);
nand U10181 (N_10181,N_9442,N_9320);
or U10182 (N_10182,N_9167,N_8963);
or U10183 (N_10183,N_9746,N_9375);
nor U10184 (N_10184,N_8765,N_8139);
or U10185 (N_10185,N_8291,N_9068);
nand U10186 (N_10186,N_9915,N_8508);
or U10187 (N_10187,N_9239,N_9273);
nand U10188 (N_10188,N_9744,N_9445);
nand U10189 (N_10189,N_9381,N_8390);
nor U10190 (N_10190,N_8815,N_9547);
nand U10191 (N_10191,N_8085,N_8084);
nand U10192 (N_10192,N_9146,N_8552);
nand U10193 (N_10193,N_9310,N_8191);
or U10194 (N_10194,N_8164,N_9739);
and U10195 (N_10195,N_9584,N_9911);
or U10196 (N_10196,N_9668,N_9187);
or U10197 (N_10197,N_8669,N_8838);
or U10198 (N_10198,N_9260,N_9135);
and U10199 (N_10199,N_9012,N_8924);
xnor U10200 (N_10200,N_8213,N_9107);
xor U10201 (N_10201,N_8735,N_9464);
or U10202 (N_10202,N_9636,N_8342);
and U10203 (N_10203,N_9561,N_8101);
nor U10204 (N_10204,N_8124,N_9759);
and U10205 (N_10205,N_9409,N_8952);
and U10206 (N_10206,N_8887,N_8634);
nor U10207 (N_10207,N_9361,N_9293);
or U10208 (N_10208,N_9769,N_8122);
nor U10209 (N_10209,N_9005,N_8582);
or U10210 (N_10210,N_9265,N_9162);
xnor U10211 (N_10211,N_8017,N_8416);
nand U10212 (N_10212,N_8772,N_9181);
nor U10213 (N_10213,N_8362,N_9942);
or U10214 (N_10214,N_8203,N_9696);
nand U10215 (N_10215,N_9360,N_9721);
nor U10216 (N_10216,N_8392,N_8740);
and U10217 (N_10217,N_9019,N_8703);
or U10218 (N_10218,N_9134,N_9834);
or U10219 (N_10219,N_8128,N_9904);
nor U10220 (N_10220,N_8647,N_8080);
nor U10221 (N_10221,N_9386,N_9796);
nor U10222 (N_10222,N_8358,N_8928);
nand U10223 (N_10223,N_8770,N_9794);
or U10224 (N_10224,N_9301,N_8248);
or U10225 (N_10225,N_9059,N_8319);
nand U10226 (N_10226,N_9309,N_8915);
or U10227 (N_10227,N_9808,N_8343);
nor U10228 (N_10228,N_9102,N_8201);
nand U10229 (N_10229,N_8078,N_8475);
nand U10230 (N_10230,N_8593,N_8147);
nor U10231 (N_10231,N_8993,N_9685);
nand U10232 (N_10232,N_9719,N_9469);
and U10233 (N_10233,N_8212,N_8942);
and U10234 (N_10234,N_9734,N_9551);
nor U10235 (N_10235,N_8950,N_8759);
nand U10236 (N_10236,N_9132,N_9016);
and U10237 (N_10237,N_8239,N_9406);
nor U10238 (N_10238,N_9413,N_8616);
nand U10239 (N_10239,N_9959,N_9863);
nand U10240 (N_10240,N_8752,N_8353);
nor U10241 (N_10241,N_9508,N_8836);
and U10242 (N_10242,N_9860,N_8169);
and U10243 (N_10243,N_8962,N_8447);
and U10244 (N_10244,N_8477,N_8066);
nand U10245 (N_10245,N_8680,N_8702);
and U10246 (N_10246,N_8959,N_8653);
nand U10247 (N_10247,N_9048,N_8117);
nand U10248 (N_10248,N_8068,N_9126);
and U10249 (N_10249,N_9025,N_9400);
and U10250 (N_10250,N_8288,N_9434);
nand U10251 (N_10251,N_8798,N_9877);
or U10252 (N_10252,N_8297,N_8757);
nand U10253 (N_10253,N_8638,N_8197);
nand U10254 (N_10254,N_8398,N_8774);
and U10255 (N_10255,N_8276,N_8571);
nor U10256 (N_10256,N_9727,N_8242);
or U10257 (N_10257,N_9588,N_8412);
nand U10258 (N_10258,N_8701,N_8877);
nand U10259 (N_10259,N_8873,N_8425);
or U10260 (N_10260,N_8448,N_9920);
or U10261 (N_10261,N_9186,N_8955);
and U10262 (N_10262,N_8805,N_8459);
nand U10263 (N_10263,N_8586,N_8687);
nand U10264 (N_10264,N_8786,N_9497);
xor U10265 (N_10265,N_8630,N_8445);
xor U10266 (N_10266,N_9549,N_9072);
nor U10267 (N_10267,N_8045,N_8397);
or U10268 (N_10268,N_8039,N_8507);
xnor U10269 (N_10269,N_9277,N_8324);
and U10270 (N_10270,N_9460,N_8043);
nor U10271 (N_10271,N_9524,N_8520);
and U10272 (N_10272,N_9928,N_9898);
and U10273 (N_10273,N_8211,N_9483);
nor U10274 (N_10274,N_9026,N_8548);
nand U10275 (N_10275,N_8695,N_8063);
xor U10276 (N_10276,N_9014,N_8751);
nor U10277 (N_10277,N_8761,N_9869);
and U10278 (N_10278,N_8000,N_8994);
xnor U10279 (N_10279,N_9654,N_9244);
or U10280 (N_10280,N_8190,N_9645);
xnor U10281 (N_10281,N_8142,N_9419);
or U10282 (N_10282,N_8175,N_8999);
nand U10283 (N_10283,N_8954,N_9938);
nand U10284 (N_10284,N_8684,N_9485);
xor U10285 (N_10285,N_9886,N_8883);
nand U10286 (N_10286,N_9463,N_9738);
nand U10287 (N_10287,N_9693,N_8400);
nor U10288 (N_10288,N_9338,N_8393);
nor U10289 (N_10289,N_9712,N_8781);
and U10290 (N_10290,N_8467,N_9838);
and U10291 (N_10291,N_9178,N_9842);
or U10292 (N_10292,N_8259,N_9611);
or U10293 (N_10293,N_8131,N_9493);
xor U10294 (N_10294,N_9008,N_8947);
nand U10295 (N_10295,N_8094,N_8789);
xor U10296 (N_10296,N_8371,N_9080);
or U10297 (N_10297,N_9665,N_9028);
or U10298 (N_10298,N_8617,N_9342);
nor U10299 (N_10299,N_9678,N_8719);
nor U10300 (N_10300,N_9371,N_9995);
nor U10301 (N_10301,N_9488,N_9408);
and U10302 (N_10302,N_8473,N_8829);
and U10303 (N_10303,N_8706,N_9644);
nor U10304 (N_10304,N_8383,N_8566);
nand U10305 (N_10305,N_8280,N_8707);
nand U10306 (N_10306,N_9211,N_8645);
nand U10307 (N_10307,N_9062,N_8262);
nor U10308 (N_10308,N_9233,N_8850);
nor U10309 (N_10309,N_8626,N_8296);
xnor U10310 (N_10310,N_9365,N_8439);
nand U10311 (N_10311,N_8256,N_9737);
nor U10312 (N_10312,N_9224,N_9367);
or U10313 (N_10313,N_9925,N_9088);
nor U10314 (N_10314,N_9474,N_8969);
xnor U10315 (N_10315,N_9567,N_8417);
or U10316 (N_10316,N_8575,N_9171);
nor U10317 (N_10317,N_8813,N_9758);
and U10318 (N_10318,N_9096,N_8882);
or U10319 (N_10319,N_9825,N_8869);
xor U10320 (N_10320,N_8972,N_8418);
or U10321 (N_10321,N_9377,N_8173);
xnor U10322 (N_10322,N_9216,N_9926);
nand U10323 (N_10323,N_9606,N_9057);
or U10324 (N_10324,N_9703,N_9961);
and U10325 (N_10325,N_8042,N_8001);
nand U10326 (N_10326,N_9466,N_9276);
nor U10327 (N_10327,N_9087,N_8162);
nand U10328 (N_10328,N_8670,N_9304);
or U10329 (N_10329,N_9875,N_8513);
or U10330 (N_10330,N_9701,N_8921);
or U10331 (N_10331,N_9374,N_8650);
and U10332 (N_10332,N_8833,N_9345);
nand U10333 (N_10333,N_8384,N_9192);
nor U10334 (N_10334,N_8038,N_9456);
nor U10335 (N_10335,N_9694,N_8206);
and U10336 (N_10336,N_9540,N_9675);
xnor U10337 (N_10337,N_8545,N_9065);
nand U10338 (N_10338,N_9968,N_9038);
nand U10339 (N_10339,N_8064,N_8534);
or U10340 (N_10340,N_9687,N_9615);
nand U10341 (N_10341,N_9658,N_9137);
and U10342 (N_10342,N_8841,N_8937);
nand U10343 (N_10343,N_8802,N_9780);
and U10344 (N_10344,N_9553,N_9826);
nor U10345 (N_10345,N_8388,N_9775);
nand U10346 (N_10346,N_9099,N_8356);
and U10347 (N_10347,N_9237,N_8318);
nor U10348 (N_10348,N_8474,N_9590);
and U10349 (N_10349,N_8934,N_9225);
or U10350 (N_10350,N_9683,N_9498);
or U10351 (N_10351,N_9357,N_9972);
nand U10352 (N_10352,N_8951,N_8558);
or U10353 (N_10353,N_9607,N_8666);
nor U10354 (N_10354,N_9396,N_8811);
nor U10355 (N_10355,N_9936,N_8504);
nand U10356 (N_10356,N_9757,N_9422);
nor U10357 (N_10357,N_8651,N_9586);
and U10358 (N_10358,N_9730,N_8896);
or U10359 (N_10359,N_9482,N_9458);
and U10360 (N_10360,N_9841,N_9541);
nand U10361 (N_10361,N_8313,N_8900);
or U10362 (N_10362,N_8295,N_8329);
or U10363 (N_10363,N_9499,N_9391);
nand U10364 (N_10364,N_9801,N_9195);
or U10365 (N_10365,N_8229,N_8501);
or U10366 (N_10366,N_9046,N_8378);
nor U10367 (N_10367,N_9996,N_8006);
or U10368 (N_10368,N_8260,N_9024);
or U10369 (N_10369,N_9449,N_9632);
or U10370 (N_10370,N_8531,N_9828);
nand U10371 (N_10371,N_8049,N_9070);
and U10372 (N_10372,N_9663,N_8047);
xnor U10373 (N_10373,N_8547,N_9462);
or U10374 (N_10374,N_8956,N_8434);
or U10375 (N_10375,N_9041,N_8555);
and U10376 (N_10376,N_8269,N_9956);
nor U10377 (N_10377,N_8341,N_8118);
nor U10378 (N_10378,N_9577,N_8032);
and U10379 (N_10379,N_8851,N_8251);
xor U10380 (N_10380,N_9415,N_8483);
and U10381 (N_10381,N_9529,N_8033);
nor U10382 (N_10382,N_8154,N_8826);
nor U10383 (N_10383,N_9934,N_8608);
nor U10384 (N_10384,N_9522,N_9443);
nor U10385 (N_10385,N_8535,N_9032);
and U10386 (N_10386,N_8056,N_9994);
or U10387 (N_10387,N_8013,N_9121);
nor U10388 (N_10388,N_9521,N_9332);
and U10389 (N_10389,N_8724,N_8380);
or U10390 (N_10390,N_9667,N_9144);
or U10391 (N_10391,N_8116,N_9252);
nor U10392 (N_10392,N_8189,N_9108);
and U10393 (N_10393,N_9118,N_9799);
or U10394 (N_10394,N_9716,N_9962);
nor U10395 (N_10395,N_8061,N_8468);
nor U10396 (N_10396,N_9621,N_8481);
nand U10397 (N_10397,N_8141,N_9950);
and U10398 (N_10398,N_9604,N_8729);
nand U10399 (N_10399,N_9350,N_9865);
nand U10400 (N_10400,N_9333,N_8235);
xnor U10401 (N_10401,N_8840,N_9366);
nand U10402 (N_10402,N_9783,N_8479);
or U10403 (N_10403,N_9643,N_9969);
and U10404 (N_10404,N_9790,N_9037);
or U10405 (N_10405,N_9885,N_8885);
nor U10406 (N_10406,N_8115,N_9294);
nor U10407 (N_10407,N_9525,N_9322);
nor U10408 (N_10408,N_9380,N_9944);
nor U10409 (N_10409,N_8565,N_8491);
nand U10410 (N_10410,N_8620,N_8278);
or U10411 (N_10411,N_9595,N_9978);
nor U10412 (N_10412,N_9717,N_9930);
and U10413 (N_10413,N_8506,N_9421);
or U10414 (N_10414,N_8265,N_9635);
nand U10415 (N_10415,N_9185,N_8405);
nor U10416 (N_10416,N_9715,N_8872);
and U10417 (N_10417,N_9436,N_9177);
nand U10418 (N_10418,N_9184,N_8556);
nor U10419 (N_10419,N_9516,N_9605);
nand U10420 (N_10420,N_8605,N_8200);
nand U10421 (N_10421,N_9937,N_8486);
xor U10422 (N_10422,N_8709,N_8986);
nand U10423 (N_10423,N_9420,N_9486);
or U10424 (N_10424,N_9624,N_8185);
xor U10425 (N_10425,N_9676,N_9573);
nor U10426 (N_10426,N_9690,N_8909);
or U10427 (N_10427,N_9334,N_8748);
nand U10428 (N_10428,N_8055,N_9079);
nand U10429 (N_10429,N_8402,N_8987);
and U10430 (N_10430,N_8681,N_9164);
nor U10431 (N_10431,N_9490,N_9754);
and U10432 (N_10432,N_8738,N_9344);
and U10433 (N_10433,N_8346,N_9289);
xnor U10434 (N_10434,N_9563,N_8455);
and U10435 (N_10435,N_8889,N_8600);
and U10436 (N_10436,N_8391,N_8657);
or U10437 (N_10437,N_9086,N_9234);
or U10438 (N_10438,N_8127,N_8328);
and U10439 (N_10439,N_8640,N_8633);
xor U10440 (N_10440,N_9921,N_8020);
nand U10441 (N_10441,N_9156,N_9199);
nand U10442 (N_10442,N_8176,N_9791);
or U10443 (N_10443,N_9183,N_9591);
nor U10444 (N_10444,N_9971,N_8263);
nor U10445 (N_10445,N_8255,N_9531);
nor U10446 (N_10446,N_9642,N_9906);
and U10447 (N_10447,N_8415,N_8146);
xor U10448 (N_10448,N_8528,N_9880);
and U10449 (N_10449,N_9726,N_8241);
and U10450 (N_10450,N_8591,N_8914);
nand U10451 (N_10451,N_9907,N_9329);
xor U10452 (N_10452,N_9303,N_9711);
nor U10453 (N_10453,N_9602,N_9922);
nand U10454 (N_10454,N_9941,N_9564);
nor U10455 (N_10455,N_9803,N_8525);
xor U10456 (N_10456,N_9848,N_9168);
nand U10457 (N_10457,N_8159,N_9558);
xor U10458 (N_10458,N_8648,N_9847);
and U10459 (N_10459,N_8228,N_8866);
or U10460 (N_10460,N_9063,N_8602);
nand U10461 (N_10461,N_9255,N_8432);
or U10462 (N_10462,N_8270,N_9347);
nor U10463 (N_10463,N_9314,N_9050);
nor U10464 (N_10464,N_9795,N_9281);
or U10465 (N_10465,N_9657,N_9976);
nand U10466 (N_10466,N_8949,N_9637);
nor U10467 (N_10467,N_9250,N_8423);
nor U10468 (N_10468,N_8451,N_9661);
or U10469 (N_10469,N_9998,N_8902);
nand U10470 (N_10470,N_9182,N_8379);
nand U10471 (N_10471,N_8816,N_8442);
or U10472 (N_10472,N_9492,N_9837);
xor U10473 (N_10473,N_8476,N_9550);
nand U10474 (N_10474,N_8465,N_9208);
nand U10475 (N_10475,N_9047,N_8220);
nor U10476 (N_10476,N_8696,N_9901);
xor U10477 (N_10477,N_8879,N_9044);
nor U10478 (N_10478,N_9480,N_9932);
nor U10479 (N_10479,N_9776,N_9258);
nand U10480 (N_10480,N_8012,N_8497);
nor U10481 (N_10481,N_8521,N_9818);
or U10482 (N_10482,N_9686,N_9279);
xor U10483 (N_10483,N_9136,N_9627);
xor U10484 (N_10484,N_8023,N_8271);
xnor U10485 (N_10485,N_9832,N_9429);
and U10486 (N_10486,N_8298,N_9372);
and U10487 (N_10487,N_8093,N_9587);
nor U10488 (N_10488,N_9774,N_9631);
nand U10489 (N_10489,N_8062,N_9982);
nand U10490 (N_10490,N_8615,N_9484);
nand U10491 (N_10491,N_8450,N_9035);
and U10492 (N_10492,N_8452,N_9854);
or U10493 (N_10493,N_9975,N_8060);
nor U10494 (N_10494,N_9364,N_9957);
xnor U10495 (N_10495,N_8855,N_8904);
or U10496 (N_10496,N_9054,N_8897);
nor U10497 (N_10497,N_8688,N_9807);
nand U10498 (N_10498,N_8810,N_9336);
nand U10499 (N_10499,N_9507,N_8808);
nand U10500 (N_10500,N_9899,N_9346);
nor U10501 (N_10501,N_9708,N_8453);
and U10502 (N_10502,N_8375,N_8953);
or U10503 (N_10503,N_9914,N_8496);
xor U10504 (N_10504,N_9317,N_8741);
nor U10505 (N_10505,N_9489,N_9206);
and U10506 (N_10506,N_9752,N_9515);
and U10507 (N_10507,N_8800,N_8254);
nor U10508 (N_10508,N_9152,N_8569);
nand U10509 (N_10509,N_8606,N_8720);
nor U10510 (N_10510,N_9228,N_9725);
or U10511 (N_10511,N_9128,N_8690);
nor U10512 (N_10512,N_8316,N_9749);
or U10513 (N_10513,N_8292,N_9403);
and U10514 (N_10514,N_8198,N_8050);
and U10515 (N_10515,N_8880,N_9511);
or U10516 (N_10516,N_8932,N_9532);
xnor U10517 (N_10517,N_9984,N_8273);
nand U10518 (N_10518,N_9022,N_9388);
or U10519 (N_10519,N_8110,N_8193);
or U10520 (N_10520,N_8733,N_8961);
xor U10521 (N_10521,N_8040,N_8422);
and U10522 (N_10522,N_9473,N_9539);
nor U10523 (N_10523,N_9154,N_9491);
nand U10524 (N_10524,N_8519,N_9362);
nor U10525 (N_10525,N_8881,N_8243);
and U10526 (N_10526,N_8289,N_8325);
nand U10527 (N_10527,N_9100,N_9010);
nand U10528 (N_10528,N_8188,N_8998);
or U10529 (N_10529,N_9527,N_9659);
nor U10530 (N_10530,N_8435,N_9902);
and U10531 (N_10531,N_9313,N_8138);
nand U10532 (N_10532,N_9351,N_8208);
or U10533 (N_10533,N_8564,N_9148);
nor U10534 (N_10534,N_9592,N_8480);
nor U10535 (N_10535,N_8232,N_8026);
xor U10536 (N_10536,N_8230,N_9435);
nand U10537 (N_10537,N_8510,N_9859);
nand U10538 (N_10538,N_8732,N_8734);
and U10539 (N_10539,N_9166,N_9431);
nand U10540 (N_10540,N_8968,N_8404);
or U10541 (N_10541,N_8783,N_9083);
nor U10542 (N_10542,N_8814,N_8244);
and U10543 (N_10543,N_8196,N_9426);
and U10544 (N_10544,N_9751,N_9444);
nor U10545 (N_10545,N_8076,N_8449);
and U10546 (N_10546,N_8387,N_9866);
or U10547 (N_10547,N_9954,N_9254);
nand U10548 (N_10548,N_8665,N_9720);
or U10549 (N_10549,N_8351,N_9554);
nor U10550 (N_10550,N_9977,N_8433);
or U10551 (N_10551,N_9249,N_9713);
nand U10552 (N_10552,N_8886,N_8967);
nand U10553 (N_10553,N_9949,N_8100);
and U10554 (N_10554,N_9236,N_9292);
and U10555 (N_10555,N_8758,N_9204);
xor U10556 (N_10556,N_9763,N_9471);
nand U10557 (N_10557,N_8186,N_8819);
and U10558 (N_10558,N_8743,N_9958);
nand U10559 (N_10559,N_9295,N_9891);
nand U10560 (N_10560,N_9425,N_9067);
and U10561 (N_10561,N_9997,N_9510);
nand U10562 (N_10562,N_8524,N_8386);
or U10563 (N_10563,N_8082,N_9324);
or U10564 (N_10564,N_8736,N_9398);
or U10565 (N_10565,N_9066,N_8544);
nor U10566 (N_10566,N_8527,N_9542);
nor U10567 (N_10567,N_9756,N_9191);
nor U10568 (N_10568,N_8382,N_9896);
nand U10569 (N_10569,N_9049,N_8674);
nand U10570 (N_10570,N_8536,N_9031);
nor U10571 (N_10571,N_9061,N_9074);
nand U10572 (N_10572,N_8157,N_8635);
nand U10573 (N_10573,N_9287,N_8469);
nand U10574 (N_10574,N_8293,N_9461);
nor U10575 (N_10575,N_9813,N_8643);
and U10576 (N_10576,N_8523,N_8069);
nand U10577 (N_10577,N_8174,N_8845);
nand U10578 (N_10578,N_9536,N_9155);
and U10579 (N_10579,N_9321,N_8337);
and U10580 (N_10580,N_8209,N_8210);
or U10581 (N_10581,N_8170,N_8561);
xnor U10582 (N_10582,N_9784,N_9457);
or U10583 (N_10583,N_8264,N_9098);
nor U10584 (N_10584,N_9169,N_8588);
nand U10585 (N_10585,N_8089,N_8891);
or U10586 (N_10586,N_9581,N_8090);
and U10587 (N_10587,N_8179,N_8369);
xor U10588 (N_10588,N_8817,N_9845);
and U10589 (N_10589,N_8347,N_9110);
and U10590 (N_10590,N_8321,N_8981);
or U10591 (N_10591,N_9356,N_8134);
xnor U10592 (N_10592,N_8106,N_9530);
nor U10593 (N_10593,N_9017,N_8396);
or U10594 (N_10594,N_8587,N_8868);
nand U10595 (N_10595,N_8177,N_8145);
nand U10596 (N_10596,N_9138,N_8119);
nand U10597 (N_10597,N_8916,N_8675);
and U10598 (N_10598,N_8097,N_8308);
nor U10599 (N_10599,N_8151,N_9242);
or U10600 (N_10600,N_8699,N_9131);
nor U10601 (N_10601,N_9707,N_8596);
nand U10602 (N_10602,N_9143,N_9871);
nand U10603 (N_10603,N_8573,N_8166);
and U10604 (N_10604,N_8492,N_8005);
and U10605 (N_10605,N_9545,N_9543);
xor U10606 (N_10606,N_9477,N_9714);
xor U10607 (N_10607,N_9097,N_8214);
and U10608 (N_10608,N_8854,N_8820);
or U10609 (N_10609,N_8803,N_9733);
nand U10610 (N_10610,N_8137,N_8966);
nand U10611 (N_10611,N_9109,N_9526);
nor U10612 (N_10612,N_9055,N_9337);
or U10613 (N_10613,N_8821,N_9259);
and U10614 (N_10614,N_8414,N_9003);
or U10615 (N_10615,N_8182,N_8652);
nand U10616 (N_10616,N_8046,N_8957);
xnor U10617 (N_10617,N_8183,N_9161);
or U10618 (N_10618,N_9147,N_9566);
nand U10619 (N_10619,N_8662,N_9018);
and U10620 (N_10620,N_9876,N_8590);
or U10621 (N_10621,N_8931,N_8923);
xor U10622 (N_10622,N_8580,N_9626);
xnor U10623 (N_10623,N_8488,N_9556);
nand U10624 (N_10624,N_8505,N_8268);
nor U10625 (N_10625,N_8697,N_8574);
nor U10626 (N_10626,N_8357,N_8744);
nor U10627 (N_10627,N_8300,N_9201);
and U10628 (N_10628,N_8982,N_8912);
nand U10629 (N_10629,N_9085,N_9705);
xnor U10630 (N_10630,N_8411,N_8992);
nor U10631 (N_10631,N_8304,N_9459);
and U10632 (N_10632,N_8509,N_9963);
or U10633 (N_10633,N_9704,N_9448);
nor U10634 (N_10634,N_8482,N_8463);
xnor U10635 (N_10635,N_8782,N_9384);
nand U10636 (N_10636,N_8549,N_8167);
nand U10637 (N_10637,N_8250,N_8693);
and U10638 (N_10638,N_9060,N_9267);
or U10639 (N_10639,N_8515,N_9638);
nor U10640 (N_10640,N_9011,N_8181);
nor U10641 (N_10641,N_8654,N_8875);
nand U10642 (N_10642,N_8472,N_8792);
and U10643 (N_10643,N_8095,N_9679);
nor U10644 (N_10644,N_9992,N_8649);
and U10645 (N_10645,N_9603,N_8595);
nor U10646 (N_10646,N_8152,N_9850);
nor U10647 (N_10647,N_9051,N_9270);
nor U10648 (N_10648,N_8717,N_9327);
or U10649 (N_10649,N_9819,N_8136);
and U10650 (N_10650,N_8604,N_9916);
and U10651 (N_10651,N_8426,N_8537);
nand U10652 (N_10652,N_8081,N_9517);
or U10653 (N_10653,N_9620,N_9203);
xor U10654 (N_10654,N_8015,N_8114);
xor U10655 (N_10655,N_9884,N_8224);
nand U10656 (N_10656,N_8456,N_8083);
or U10657 (N_10657,N_9221,N_8637);
and U10658 (N_10658,N_9352,N_9985);
and U10659 (N_10659,N_9747,N_9882);
nand U10660 (N_10660,N_8381,N_8828);
nand U10661 (N_10661,N_9533,N_8871);
or U10662 (N_10662,N_8294,N_8978);
nor U10663 (N_10663,N_9622,N_9986);
nand U10664 (N_10664,N_9009,N_8611);
nor U10665 (N_10665,N_8079,N_9817);
nor U10666 (N_10666,N_8299,N_8018);
and U10667 (N_10667,N_9318,N_8700);
and U10668 (N_10668,N_8111,N_9890);
or U10669 (N_10669,N_9509,N_8848);
or U10670 (N_10670,N_9771,N_8306);
and U10671 (N_10671,N_8940,N_9948);
or U10672 (N_10672,N_8857,N_8859);
and U10673 (N_10673,N_9981,N_9619);
nand U10674 (N_10674,N_9407,N_9153);
nor U10675 (N_10675,N_9023,N_9504);
xor U10676 (N_10676,N_8489,N_9742);
or U10677 (N_10677,N_8330,N_8087);
nor U10678 (N_10678,N_8207,N_8360);
or U10679 (N_10679,N_9571,N_8205);
or U10680 (N_10680,N_8834,N_8925);
nand U10681 (N_10681,N_9379,N_8389);
xor U10682 (N_10682,N_8327,N_9874);
and U10683 (N_10683,N_9770,N_9789);
nor U10684 (N_10684,N_9090,N_9785);
nand U10685 (N_10685,N_9735,N_8310);
xor U10686 (N_10686,N_9501,N_8795);
xor U10687 (N_10687,N_8656,N_8309);
and U10688 (N_10688,N_9212,N_8394);
and U10689 (N_10689,N_8517,N_8618);
and U10690 (N_10690,N_9369,N_8570);
nor U10691 (N_10691,N_9680,N_8130);
and U10692 (N_10692,N_8756,N_8901);
nand U10693 (N_10693,N_8970,N_8920);
or U10694 (N_10694,N_8311,N_8374);
nor U10695 (N_10695,N_9815,N_8975);
or U10696 (N_10696,N_8530,N_8143);
xor U10697 (N_10697,N_8822,N_9290);
nor U10698 (N_10698,N_9222,N_9673);
and U10699 (N_10699,N_8661,N_9296);
or U10700 (N_10700,N_8514,N_9437);
nor U10701 (N_10701,N_8113,N_9651);
nand U10702 (N_10702,N_9373,N_9736);
nor U10703 (N_10703,N_8823,N_8831);
nor U10704 (N_10704,N_8058,N_9030);
nand U10705 (N_10705,N_9455,N_8589);
nor U10706 (N_10706,N_8503,N_9830);
and U10707 (N_10707,N_9506,N_8922);
or U10708 (N_10708,N_9900,N_8677);
or U10709 (N_10709,N_8065,N_9122);
or U10710 (N_10710,N_9940,N_8075);
nand U10711 (N_10711,N_8746,N_8457);
and U10712 (N_10712,N_9325,N_9034);
or U10713 (N_10713,N_9855,N_9432);
or U10714 (N_10714,N_9918,N_8585);
nand U10715 (N_10715,N_9781,N_9285);
nor U10716 (N_10716,N_9150,N_9741);
xor U10717 (N_10717,N_9302,N_9069);
xor U10718 (N_10718,N_9535,N_9893);
nand U10719 (N_10719,N_9649,N_8898);
nor U10720 (N_10720,N_9630,N_8964);
xor U10721 (N_10721,N_8171,N_8938);
nand U10722 (N_10722,N_8613,N_9805);
and U10723 (N_10723,N_8516,N_9613);
or U10724 (N_10724,N_8287,N_9230);
and U10725 (N_10725,N_9538,N_9387);
or U10726 (N_10726,N_9094,N_9857);
or U10727 (N_10727,N_8532,N_9188);
xnor U10728 (N_10728,N_9933,N_9840);
nor U10729 (N_10729,N_9570,N_9827);
or U10730 (N_10730,N_9991,N_9760);
and U10731 (N_10731,N_9650,N_8464);
xnor U10732 (N_10732,N_9753,N_8908);
or U10733 (N_10733,N_9677,N_9809);
and U10734 (N_10734,N_8809,N_9307);
nor U10735 (N_10735,N_8764,N_8261);
or U10736 (N_10736,N_8787,N_8579);
and U10737 (N_10737,N_8919,N_8052);
nor U10738 (N_10738,N_8332,N_8219);
or U10739 (N_10739,N_9073,N_8726);
xor U10740 (N_10740,N_9706,N_8679);
or U10741 (N_10741,N_8004,N_9585);
nand U10742 (N_10742,N_9446,N_9214);
nor U10743 (N_10743,N_9648,N_8267);
or U10744 (N_10744,N_8718,N_8408);
or U10745 (N_10745,N_9274,N_9692);
nand U10746 (N_10746,N_8471,N_8678);
nand U10747 (N_10747,N_8035,N_9202);
nor U10748 (N_10748,N_9209,N_8903);
nor U10749 (N_10749,N_9810,N_9219);
nand U10750 (N_10750,N_8072,N_9773);
nor U10751 (N_10751,N_9856,N_9278);
nor U10752 (N_10752,N_9792,N_8562);
nor U10753 (N_10753,N_8320,N_8708);
and U10754 (N_10754,N_8070,N_8466);
and U10755 (N_10755,N_8984,N_8437);
nand U10756 (N_10756,N_8769,N_8231);
nand U10757 (N_10757,N_9786,N_8686);
nand U10758 (N_10758,N_8285,N_9112);
nor U10759 (N_10759,N_9710,N_8584);
nor U10760 (N_10760,N_8234,N_8312);
xnor U10761 (N_10761,N_9205,N_9139);
nor U10762 (N_10762,N_8165,N_8827);
or U10763 (N_10763,N_9213,N_9623);
nand U10764 (N_10764,N_8403,N_9616);
or U10765 (N_10765,N_8890,N_9468);
nor U10766 (N_10766,N_9306,N_8960);
or U10767 (N_10767,N_9664,N_8936);
nor U10768 (N_10768,N_8745,N_8976);
nand U10769 (N_10769,N_9582,N_8314);
nand U10770 (N_10770,N_9814,N_9887);
or U10771 (N_10771,N_9001,N_9502);
or U10772 (N_10772,N_9518,N_9964);
nand U10773 (N_10773,N_8788,N_8286);
nor U10774 (N_10774,N_8730,N_8550);
and U10775 (N_10775,N_9946,N_9454);
nand U10776 (N_10776,N_9743,N_9262);
nor U10777 (N_10777,N_9698,N_9919);
or U10778 (N_10778,N_9688,N_9157);
and U10779 (N_10779,N_9000,N_9888);
nor U10780 (N_10780,N_8812,N_8858);
or U10781 (N_10781,N_9404,N_8108);
nor U10782 (N_10782,N_9641,N_8123);
xor U10783 (N_10783,N_8022,N_8658);
and U10784 (N_10784,N_8659,N_8133);
and U10785 (N_10785,N_9246,N_8973);
or U10786 (N_10786,N_9689,N_9475);
or U10787 (N_10787,N_8712,N_8150);
nand U10788 (N_10788,N_8603,N_8024);
or U10789 (N_10789,N_9913,N_9793);
or U10790 (N_10790,N_8037,N_8755);
xor U10791 (N_10791,N_8572,N_9839);
nor U10792 (N_10792,N_8577,N_9389);
nor U10793 (N_10793,N_8019,N_8180);
nand U10794 (N_10794,N_8791,N_9797);
nand U10795 (N_10795,N_9410,N_8249);
nand U10796 (N_10796,N_9505,N_9952);
nor U10797 (N_10797,N_8352,N_9151);
nand U10798 (N_10798,N_8227,N_9660);
and U10799 (N_10799,N_9528,N_8044);
xnor U10800 (N_10800,N_8779,N_9965);
nor U10801 (N_10801,N_8560,N_8098);
nand U10802 (N_10802,N_8583,N_9311);
nand U10803 (N_10803,N_9042,N_9849);
xor U10804 (N_10804,N_9076,N_9671);
or U10805 (N_10805,N_9091,N_9666);
and U10806 (N_10806,N_9395,N_8163);
nand U10807 (N_10807,N_9924,N_8639);
nor U10808 (N_10808,N_8077,N_9229);
nor U10809 (N_10809,N_9682,N_8884);
nor U10810 (N_10810,N_9745,N_9798);
and U10811 (N_10811,N_8754,N_9174);
nor U10812 (N_10812,N_9523,N_8991);
and U10813 (N_10813,N_8192,N_8711);
nor U10814 (N_10814,N_8366,N_8233);
nand U10815 (N_10815,N_8636,N_9767);
nand U10816 (N_10816,N_8223,N_8594);
and U10817 (N_10817,N_8763,N_8454);
and U10818 (N_10818,N_8793,N_9256);
nand U10819 (N_10819,N_9002,N_9927);
nand U10820 (N_10820,N_9341,N_8344);
nand U10821 (N_10821,N_9084,N_9021);
nor U10822 (N_10822,N_9358,N_9058);
or U10823 (N_10823,N_8971,N_9340);
nand U10824 (N_10824,N_8725,N_8860);
or U10825 (N_10825,N_9947,N_8609);
and U10826 (N_10826,N_8835,N_9349);
nand U10827 (N_10827,N_8172,N_9385);
nor U10828 (N_10828,N_9376,N_9297);
and U10829 (N_10829,N_9330,N_8364);
nor U10830 (N_10830,N_8983,N_9778);
nor U10831 (N_10831,N_8996,N_9892);
nor U10832 (N_10832,N_8767,N_9569);
nor U10833 (N_10833,N_9235,N_9647);
nor U10834 (N_10834,N_9846,N_9160);
or U10835 (N_10835,N_8440,N_9609);
and U10836 (N_10836,N_8762,N_9271);
or U10837 (N_10837,N_8226,N_8567);
and U10838 (N_10838,N_8057,N_9691);
nand U10839 (N_10839,N_9897,N_9207);
xor U10840 (N_10840,N_8301,N_8290);
and U10841 (N_10841,N_9572,N_9397);
or U10842 (N_10842,N_8258,N_9308);
or U10843 (N_10843,N_9248,N_9662);
and U10844 (N_10844,N_8958,N_9782);
nand U10845 (N_10845,N_9568,N_9125);
and U10846 (N_10846,N_9326,N_9251);
nor U10847 (N_10847,N_8502,N_9064);
nand U10848 (N_10848,N_8905,N_9354);
nand U10849 (N_10849,N_8631,N_9844);
and U10850 (N_10850,N_9852,N_9831);
nor U10851 (N_10851,N_9966,N_9476);
nand U10852 (N_10852,N_8140,N_9261);
and U10853 (N_10853,N_9127,N_8737);
and U10854 (N_10854,N_8546,N_9851);
or U10855 (N_10855,N_8365,N_8775);
nor U10856 (N_10856,N_8429,N_8216);
xnor U10857 (N_10857,N_8460,N_8338);
nand U10858 (N_10858,N_9974,N_8554);
and U10859 (N_10859,N_9513,N_9988);
xor U10860 (N_10860,N_9433,N_9231);
nand U10861 (N_10861,N_9881,N_9999);
and U10862 (N_10862,N_8331,N_8237);
or U10863 (N_10863,N_8407,N_9439);
nand U10864 (N_10864,N_9858,N_8979);
or U10865 (N_10865,N_9800,N_8377);
nor U10866 (N_10866,N_8944,N_8722);
nand U10867 (N_10867,N_9653,N_9864);
nand U10868 (N_10868,N_9163,N_9257);
nor U10869 (N_10869,N_8446,N_9078);
nand U10870 (N_10870,N_8870,N_8863);
and U10871 (N_10871,N_8990,N_8413);
xor U10872 (N_10872,N_8036,N_9393);
nand U10873 (N_10873,N_8253,N_9779);
nand U10874 (N_10874,N_9544,N_8749);
and U10875 (N_10875,N_8627,N_9823);
xor U10876 (N_10876,N_8878,N_8918);
xnor U10877 (N_10877,N_8367,N_9052);
xor U10878 (N_10878,N_8401,N_8676);
or U10879 (N_10879,N_8470,N_9082);
or U10880 (N_10880,N_8215,N_8610);
and U10881 (N_10881,N_9383,N_9299);
nor U10882 (N_10882,N_8867,N_9599);
or U10883 (N_10883,N_9935,N_8121);
nand U10884 (N_10884,N_9210,N_9494);
nand U10885 (N_10885,N_9179,N_9004);
nand U10886 (N_10886,N_9368,N_8856);
or U10887 (N_10887,N_9399,N_9411);
or U10888 (N_10888,N_9788,N_8348);
nor U10889 (N_10889,N_8797,N_8965);
or U10890 (N_10890,N_8245,N_8054);
nor U10891 (N_10891,N_8668,N_9378);
nor U10892 (N_10892,N_9600,N_9750);
nand U10893 (N_10893,N_8279,N_9275);
and U10894 (N_10894,N_8518,N_9633);
and U10895 (N_10895,N_8723,N_8368);
nand U10896 (N_10896,N_8716,N_8372);
nand U10897 (N_10897,N_9479,N_8349);
or U10898 (N_10898,N_9272,N_8980);
nor U10899 (N_10899,N_8156,N_9970);
and U10900 (N_10900,N_8663,N_8832);
or U10901 (N_10901,N_9075,N_9478);
and U10902 (N_10902,N_9598,N_9811);
or U10903 (N_10903,N_9802,N_8406);
nand U10904 (N_10904,N_9238,N_8041);
nand U10905 (N_10905,N_9200,N_8790);
xor U10906 (N_10906,N_8307,N_8917);
nor U10907 (N_10907,N_9331,N_8698);
or U10908 (N_10908,N_8843,N_8876);
or U10909 (N_10909,N_8444,N_9960);
and U10910 (N_10910,N_8028,N_9189);
nand U10911 (N_10911,N_8048,N_9335);
or U10912 (N_10912,N_8893,N_8007);
and U10913 (N_10913,N_8526,N_9232);
xor U10914 (N_10914,N_8672,N_8664);
and U10915 (N_10915,N_9253,N_9820);
nand U10916 (N_10916,N_8892,N_9215);
nor U10917 (N_10917,N_9709,N_9286);
nor U10918 (N_10918,N_9496,N_8776);
and U10919 (N_10919,N_9348,N_8607);
nor U10920 (N_10920,N_8428,N_9440);
or U10921 (N_10921,N_9503,N_9917);
or U10922 (N_10922,N_8107,N_8623);
nand U10923 (N_10923,N_9359,N_9268);
nor U10924 (N_10924,N_9583,N_9217);
nor U10925 (N_10925,N_8334,N_8317);
and U10926 (N_10926,N_9103,N_8731);
nand U10927 (N_10927,N_9723,N_9806);
nor U10928 (N_10928,N_9193,N_8091);
xnor U10929 (N_10929,N_9043,N_8844);
or U10930 (N_10930,N_8830,N_9006);
and U10931 (N_10931,N_9220,N_8714);
or U10932 (N_10932,N_9989,N_8768);
and U10933 (N_10933,N_9053,N_8125);
or U10934 (N_10934,N_8861,N_8462);
xnor U10935 (N_10935,N_8409,N_9903);
nor U10936 (N_10936,N_9264,N_8485);
and U10937 (N_10937,N_8807,N_9416);
xnor U10938 (N_10938,N_8284,N_8694);
nand U10939 (N_10939,N_9534,N_8029);
nand U10940 (N_10940,N_8837,N_8895);
xnor U10941 (N_10941,N_8874,N_9145);
and U10942 (N_10942,N_9520,N_8282);
and U10943 (N_10943,N_9427,N_8410);
nor U10944 (N_10944,N_8894,N_8399);
and U10945 (N_10945,N_9943,N_9824);
and U10946 (N_10946,N_8126,N_8336);
nand U10947 (N_10947,N_9601,N_9931);
nor U10948 (N_10948,N_9291,N_9453);
nand U10949 (N_10949,N_8340,N_8011);
or U10950 (N_10950,N_8945,N_9559);
and U10951 (N_10951,N_8760,N_8578);
nor U10952 (N_10952,N_8421,N_8322);
xnor U10953 (N_10953,N_8685,N_9412);
nor U10954 (N_10954,N_8655,N_9196);
and U10955 (N_10955,N_9095,N_8204);
or U10956 (N_10956,N_9300,N_9414);
and U10957 (N_10957,N_8728,N_9555);
nor U10958 (N_10958,N_8225,N_8363);
nand U10959 (N_10959,N_8541,N_8281);
or U10960 (N_10960,N_9945,N_8721);
or U10961 (N_10961,N_9173,N_9562);
or U10962 (N_10962,N_8710,N_8096);
nor U10963 (N_10963,N_8926,N_8592);
nand U10964 (N_10964,N_8178,N_8149);
and U10965 (N_10965,N_9724,N_8785);
and U10966 (N_10966,N_8646,N_8160);
nand U10967 (N_10967,N_9465,N_9172);
nor U10968 (N_10968,N_9282,N_8430);
and U10969 (N_10969,N_9873,N_9029);
nand U10970 (N_10970,N_9487,N_9639);
nand U10971 (N_10971,N_9343,N_9240);
nor U10972 (N_10972,N_8539,N_9574);
xor U10973 (N_10973,N_9593,N_8010);
xnor U10974 (N_10974,N_9761,N_8252);
and U10975 (N_10975,N_8865,N_9438);
nand U10976 (N_10976,N_9165,N_9909);
or U10977 (N_10977,N_9596,N_8272);
nand U10978 (N_10978,N_8086,N_9787);
nand U10979 (N_10979,N_8910,N_8671);
xnor U10980 (N_10980,N_9912,N_9355);
or U10981 (N_10981,N_8339,N_9390);
nor U10982 (N_10982,N_8705,N_8689);
and U10983 (N_10983,N_9428,N_8818);
and U10984 (N_10984,N_9835,N_9470);
nor U10985 (N_10985,N_8715,N_9472);
and U10986 (N_10986,N_9117,N_8946);
and U10987 (N_10987,N_8597,N_8323);
and U10988 (N_10988,N_8008,N_8559);
or U10989 (N_10989,N_8995,N_9226);
nand U10990 (N_10990,N_9441,N_9081);
or U10991 (N_10991,N_8359,N_9777);
or U10992 (N_10992,N_9514,N_9894);
and U10993 (N_10993,N_8345,N_9768);
xnor U10994 (N_10994,N_9762,N_8747);
or U10995 (N_10995,N_9101,N_8326);
and U10996 (N_10996,N_9629,N_9729);
and U10997 (N_10997,N_8704,N_8629);
and U10998 (N_10998,N_8112,N_8753);
xnor U10999 (N_10999,N_9740,N_8576);
or U11000 (N_11000,N_9492,N_8843);
nand U11001 (N_11001,N_8952,N_8328);
or U11002 (N_11002,N_9132,N_9696);
nor U11003 (N_11003,N_9148,N_8798);
and U11004 (N_11004,N_9977,N_8682);
nand U11005 (N_11005,N_9858,N_8208);
or U11006 (N_11006,N_8132,N_9585);
or U11007 (N_11007,N_9587,N_8518);
nand U11008 (N_11008,N_9497,N_8345);
nor U11009 (N_11009,N_8107,N_8366);
nor U11010 (N_11010,N_9009,N_8337);
nand U11011 (N_11011,N_9680,N_8078);
nand U11012 (N_11012,N_9775,N_8957);
or U11013 (N_11013,N_9022,N_8392);
xor U11014 (N_11014,N_8271,N_8097);
nand U11015 (N_11015,N_9808,N_8289);
nand U11016 (N_11016,N_8648,N_9006);
nor U11017 (N_11017,N_8564,N_9885);
or U11018 (N_11018,N_8461,N_8905);
nor U11019 (N_11019,N_8618,N_9452);
xor U11020 (N_11020,N_8665,N_9763);
nand U11021 (N_11021,N_8928,N_8348);
nor U11022 (N_11022,N_9748,N_8113);
or U11023 (N_11023,N_9263,N_9024);
nor U11024 (N_11024,N_8871,N_8841);
or U11025 (N_11025,N_8728,N_9097);
nor U11026 (N_11026,N_9666,N_8902);
nor U11027 (N_11027,N_9840,N_8548);
or U11028 (N_11028,N_8141,N_9452);
nand U11029 (N_11029,N_8472,N_9049);
xor U11030 (N_11030,N_8223,N_8325);
nor U11031 (N_11031,N_9683,N_8100);
nand U11032 (N_11032,N_9710,N_8214);
xor U11033 (N_11033,N_9771,N_9566);
and U11034 (N_11034,N_8568,N_9885);
nand U11035 (N_11035,N_8987,N_9347);
xor U11036 (N_11036,N_9542,N_8441);
nor U11037 (N_11037,N_8275,N_9288);
and U11038 (N_11038,N_8491,N_9316);
and U11039 (N_11039,N_8421,N_8150);
or U11040 (N_11040,N_8762,N_9347);
nand U11041 (N_11041,N_9265,N_9684);
nor U11042 (N_11042,N_9022,N_9813);
xnor U11043 (N_11043,N_8959,N_9024);
and U11044 (N_11044,N_9394,N_9743);
nand U11045 (N_11045,N_8916,N_9869);
nand U11046 (N_11046,N_9166,N_9422);
or U11047 (N_11047,N_9583,N_8707);
or U11048 (N_11048,N_9887,N_8103);
or U11049 (N_11049,N_9681,N_8387);
xor U11050 (N_11050,N_8573,N_9618);
or U11051 (N_11051,N_8044,N_9704);
or U11052 (N_11052,N_8676,N_9228);
nor U11053 (N_11053,N_9218,N_8552);
or U11054 (N_11054,N_9408,N_8092);
nor U11055 (N_11055,N_8736,N_9043);
nand U11056 (N_11056,N_8326,N_9627);
and U11057 (N_11057,N_8909,N_9040);
and U11058 (N_11058,N_8279,N_8758);
nor U11059 (N_11059,N_8386,N_9742);
nor U11060 (N_11060,N_8654,N_9896);
or U11061 (N_11061,N_9126,N_9760);
xor U11062 (N_11062,N_9306,N_9001);
nor U11063 (N_11063,N_9307,N_9487);
nand U11064 (N_11064,N_9210,N_8611);
and U11065 (N_11065,N_9810,N_9965);
nor U11066 (N_11066,N_9975,N_9468);
or U11067 (N_11067,N_8114,N_8387);
or U11068 (N_11068,N_8011,N_8937);
nor U11069 (N_11069,N_9272,N_8545);
nand U11070 (N_11070,N_9208,N_8850);
nand U11071 (N_11071,N_9152,N_8015);
nand U11072 (N_11072,N_9038,N_9888);
nor U11073 (N_11073,N_8540,N_8223);
nor U11074 (N_11074,N_9522,N_8885);
nand U11075 (N_11075,N_9334,N_9559);
and U11076 (N_11076,N_8636,N_8959);
or U11077 (N_11077,N_8749,N_8162);
or U11078 (N_11078,N_8106,N_9503);
nor U11079 (N_11079,N_8325,N_8400);
nor U11080 (N_11080,N_9749,N_8348);
nand U11081 (N_11081,N_9420,N_9711);
nor U11082 (N_11082,N_8888,N_9877);
nor U11083 (N_11083,N_9799,N_9628);
nor U11084 (N_11084,N_9275,N_9964);
or U11085 (N_11085,N_9277,N_9880);
xor U11086 (N_11086,N_9179,N_9194);
nor U11087 (N_11087,N_8856,N_9557);
and U11088 (N_11088,N_8748,N_8124);
nand U11089 (N_11089,N_9885,N_8830);
or U11090 (N_11090,N_8754,N_8638);
nand U11091 (N_11091,N_9980,N_9315);
nand U11092 (N_11092,N_8919,N_8089);
nor U11093 (N_11093,N_8984,N_9953);
nor U11094 (N_11094,N_8662,N_9656);
and U11095 (N_11095,N_9892,N_9025);
xor U11096 (N_11096,N_8485,N_8810);
or U11097 (N_11097,N_8112,N_9448);
nor U11098 (N_11098,N_9780,N_9275);
or U11099 (N_11099,N_9238,N_8170);
and U11100 (N_11100,N_8632,N_8915);
nor U11101 (N_11101,N_9589,N_9770);
nand U11102 (N_11102,N_8382,N_9237);
or U11103 (N_11103,N_8578,N_8192);
or U11104 (N_11104,N_9322,N_9554);
or U11105 (N_11105,N_9034,N_8051);
nand U11106 (N_11106,N_8819,N_9863);
xnor U11107 (N_11107,N_8794,N_9972);
and U11108 (N_11108,N_9954,N_8888);
nor U11109 (N_11109,N_8293,N_9023);
and U11110 (N_11110,N_8117,N_8491);
or U11111 (N_11111,N_9898,N_9392);
nand U11112 (N_11112,N_8645,N_9060);
nand U11113 (N_11113,N_8266,N_9090);
nor U11114 (N_11114,N_9711,N_9450);
xnor U11115 (N_11115,N_8628,N_8401);
or U11116 (N_11116,N_9538,N_9147);
nand U11117 (N_11117,N_9538,N_9227);
nand U11118 (N_11118,N_8184,N_9249);
nor U11119 (N_11119,N_8295,N_9470);
nand U11120 (N_11120,N_9395,N_8148);
and U11121 (N_11121,N_9883,N_8628);
and U11122 (N_11122,N_8829,N_9333);
and U11123 (N_11123,N_8954,N_9211);
and U11124 (N_11124,N_8315,N_8909);
and U11125 (N_11125,N_9715,N_9017);
nand U11126 (N_11126,N_9594,N_9714);
nor U11127 (N_11127,N_8456,N_8453);
or U11128 (N_11128,N_9828,N_8701);
and U11129 (N_11129,N_9012,N_9528);
and U11130 (N_11130,N_8143,N_8582);
and U11131 (N_11131,N_8875,N_9427);
nor U11132 (N_11132,N_8453,N_8408);
nand U11133 (N_11133,N_9204,N_9510);
xnor U11134 (N_11134,N_8191,N_9420);
nand U11135 (N_11135,N_8717,N_8419);
nor U11136 (N_11136,N_8523,N_9019);
nor U11137 (N_11137,N_9573,N_9838);
nand U11138 (N_11138,N_8780,N_8231);
and U11139 (N_11139,N_8424,N_8842);
and U11140 (N_11140,N_9850,N_8387);
xor U11141 (N_11141,N_9721,N_9775);
or U11142 (N_11142,N_8914,N_8169);
or U11143 (N_11143,N_9427,N_8901);
or U11144 (N_11144,N_9832,N_9246);
nor U11145 (N_11145,N_8490,N_8000);
nand U11146 (N_11146,N_9629,N_9922);
nand U11147 (N_11147,N_8733,N_9551);
nand U11148 (N_11148,N_8534,N_8956);
nor U11149 (N_11149,N_8995,N_9111);
or U11150 (N_11150,N_8240,N_9566);
and U11151 (N_11151,N_8162,N_9453);
nand U11152 (N_11152,N_8525,N_9997);
or U11153 (N_11153,N_9052,N_9066);
and U11154 (N_11154,N_8195,N_8547);
xnor U11155 (N_11155,N_8677,N_8936);
nand U11156 (N_11156,N_9997,N_8132);
nor U11157 (N_11157,N_9204,N_8641);
nand U11158 (N_11158,N_8162,N_9952);
nand U11159 (N_11159,N_9986,N_8753);
or U11160 (N_11160,N_9647,N_9163);
and U11161 (N_11161,N_9049,N_9299);
nor U11162 (N_11162,N_8263,N_8779);
nor U11163 (N_11163,N_8217,N_9961);
nand U11164 (N_11164,N_8097,N_8282);
and U11165 (N_11165,N_9733,N_9535);
xor U11166 (N_11166,N_9108,N_9034);
or U11167 (N_11167,N_8147,N_8016);
nand U11168 (N_11168,N_8260,N_8419);
nand U11169 (N_11169,N_8911,N_8997);
nor U11170 (N_11170,N_9078,N_8039);
xnor U11171 (N_11171,N_9350,N_9586);
or U11172 (N_11172,N_9204,N_8473);
or U11173 (N_11173,N_8494,N_9981);
nand U11174 (N_11174,N_8487,N_9008);
nand U11175 (N_11175,N_8060,N_9747);
and U11176 (N_11176,N_8923,N_9321);
or U11177 (N_11177,N_8116,N_9939);
xor U11178 (N_11178,N_9350,N_8904);
nand U11179 (N_11179,N_9098,N_8268);
nor U11180 (N_11180,N_8854,N_9337);
or U11181 (N_11181,N_8799,N_8687);
and U11182 (N_11182,N_8522,N_9694);
and U11183 (N_11183,N_8460,N_9727);
or U11184 (N_11184,N_8280,N_8514);
nand U11185 (N_11185,N_8022,N_9645);
nor U11186 (N_11186,N_8942,N_8185);
xor U11187 (N_11187,N_9536,N_9791);
nand U11188 (N_11188,N_9088,N_9356);
and U11189 (N_11189,N_9334,N_8928);
or U11190 (N_11190,N_8562,N_9049);
nand U11191 (N_11191,N_8614,N_8475);
nor U11192 (N_11192,N_8413,N_8096);
or U11193 (N_11193,N_9153,N_9866);
xnor U11194 (N_11194,N_9660,N_9886);
nor U11195 (N_11195,N_8558,N_9275);
nand U11196 (N_11196,N_9160,N_8654);
xor U11197 (N_11197,N_9658,N_8454);
and U11198 (N_11198,N_9530,N_9969);
nor U11199 (N_11199,N_8604,N_9271);
xnor U11200 (N_11200,N_9203,N_9493);
nand U11201 (N_11201,N_9389,N_9146);
or U11202 (N_11202,N_8676,N_9600);
nor U11203 (N_11203,N_8676,N_9660);
and U11204 (N_11204,N_8427,N_8592);
or U11205 (N_11205,N_9023,N_8390);
nand U11206 (N_11206,N_9903,N_9199);
or U11207 (N_11207,N_8658,N_8344);
nor U11208 (N_11208,N_8401,N_8638);
or U11209 (N_11209,N_9084,N_8863);
xnor U11210 (N_11210,N_9426,N_9659);
xnor U11211 (N_11211,N_9103,N_8554);
nor U11212 (N_11212,N_9070,N_9544);
nor U11213 (N_11213,N_8091,N_9921);
and U11214 (N_11214,N_8028,N_8384);
and U11215 (N_11215,N_8236,N_9986);
nor U11216 (N_11216,N_9912,N_9047);
and U11217 (N_11217,N_8541,N_9260);
nand U11218 (N_11218,N_8023,N_9464);
or U11219 (N_11219,N_9694,N_9970);
nand U11220 (N_11220,N_9287,N_8281);
nand U11221 (N_11221,N_9107,N_9425);
nand U11222 (N_11222,N_9920,N_8589);
nor U11223 (N_11223,N_9604,N_9633);
nand U11224 (N_11224,N_8455,N_8544);
nand U11225 (N_11225,N_8409,N_8935);
or U11226 (N_11226,N_8541,N_9791);
or U11227 (N_11227,N_8801,N_8323);
nand U11228 (N_11228,N_8416,N_8853);
or U11229 (N_11229,N_9712,N_9777);
and U11230 (N_11230,N_8749,N_9454);
nand U11231 (N_11231,N_8536,N_9788);
nor U11232 (N_11232,N_8965,N_9308);
nor U11233 (N_11233,N_9372,N_9124);
or U11234 (N_11234,N_9083,N_8765);
and U11235 (N_11235,N_9124,N_8802);
or U11236 (N_11236,N_9504,N_8310);
and U11237 (N_11237,N_8865,N_9694);
and U11238 (N_11238,N_9733,N_9695);
nor U11239 (N_11239,N_9753,N_8316);
nand U11240 (N_11240,N_9949,N_9131);
xor U11241 (N_11241,N_8495,N_9830);
nand U11242 (N_11242,N_8262,N_8957);
or U11243 (N_11243,N_8970,N_9560);
nand U11244 (N_11244,N_8169,N_9771);
or U11245 (N_11245,N_8464,N_9049);
or U11246 (N_11246,N_8305,N_8763);
or U11247 (N_11247,N_9638,N_8691);
and U11248 (N_11248,N_9617,N_8135);
or U11249 (N_11249,N_8503,N_8463);
and U11250 (N_11250,N_9840,N_8132);
and U11251 (N_11251,N_8179,N_8697);
or U11252 (N_11252,N_9505,N_9341);
nor U11253 (N_11253,N_8950,N_9935);
and U11254 (N_11254,N_8300,N_9025);
and U11255 (N_11255,N_8833,N_9803);
and U11256 (N_11256,N_9173,N_9223);
or U11257 (N_11257,N_9603,N_8990);
or U11258 (N_11258,N_9348,N_9045);
nor U11259 (N_11259,N_9150,N_9339);
nand U11260 (N_11260,N_9258,N_8306);
or U11261 (N_11261,N_8477,N_9009);
nand U11262 (N_11262,N_8974,N_8212);
and U11263 (N_11263,N_9605,N_9980);
nor U11264 (N_11264,N_8517,N_8583);
nor U11265 (N_11265,N_9266,N_8070);
nand U11266 (N_11266,N_9544,N_9960);
or U11267 (N_11267,N_8377,N_8468);
nand U11268 (N_11268,N_8316,N_9306);
xor U11269 (N_11269,N_8304,N_8220);
or U11270 (N_11270,N_8744,N_9913);
and U11271 (N_11271,N_9124,N_8564);
nand U11272 (N_11272,N_8837,N_9674);
or U11273 (N_11273,N_9826,N_8309);
and U11274 (N_11274,N_8942,N_8433);
and U11275 (N_11275,N_8965,N_8679);
and U11276 (N_11276,N_9850,N_8474);
nand U11277 (N_11277,N_9052,N_8370);
and U11278 (N_11278,N_8639,N_9484);
xnor U11279 (N_11279,N_8884,N_8314);
and U11280 (N_11280,N_9613,N_9248);
or U11281 (N_11281,N_9314,N_9005);
or U11282 (N_11282,N_8209,N_8011);
nand U11283 (N_11283,N_8539,N_9736);
nor U11284 (N_11284,N_9735,N_8297);
nand U11285 (N_11285,N_9669,N_8860);
nor U11286 (N_11286,N_8851,N_8440);
xor U11287 (N_11287,N_8947,N_9042);
nor U11288 (N_11288,N_9143,N_9819);
and U11289 (N_11289,N_8059,N_9845);
nand U11290 (N_11290,N_9097,N_9072);
or U11291 (N_11291,N_9574,N_8026);
xnor U11292 (N_11292,N_8345,N_8311);
nand U11293 (N_11293,N_9378,N_8659);
xor U11294 (N_11294,N_9282,N_8923);
or U11295 (N_11295,N_9085,N_8519);
nor U11296 (N_11296,N_8110,N_8789);
or U11297 (N_11297,N_9469,N_8577);
and U11298 (N_11298,N_8058,N_8811);
nor U11299 (N_11299,N_9338,N_9993);
nand U11300 (N_11300,N_8648,N_8205);
nand U11301 (N_11301,N_8772,N_8776);
or U11302 (N_11302,N_8786,N_8871);
or U11303 (N_11303,N_8576,N_9515);
and U11304 (N_11304,N_8960,N_8946);
xor U11305 (N_11305,N_8729,N_9361);
and U11306 (N_11306,N_8179,N_8691);
xnor U11307 (N_11307,N_9168,N_8521);
nand U11308 (N_11308,N_8304,N_8674);
and U11309 (N_11309,N_9442,N_8887);
nor U11310 (N_11310,N_8265,N_9705);
or U11311 (N_11311,N_9824,N_8179);
and U11312 (N_11312,N_8712,N_8027);
or U11313 (N_11313,N_9138,N_9184);
xnor U11314 (N_11314,N_9922,N_8516);
nor U11315 (N_11315,N_9491,N_9170);
xnor U11316 (N_11316,N_9607,N_8257);
or U11317 (N_11317,N_9139,N_8029);
nor U11318 (N_11318,N_9657,N_9136);
or U11319 (N_11319,N_8947,N_9463);
nor U11320 (N_11320,N_8498,N_9342);
or U11321 (N_11321,N_8207,N_9811);
nor U11322 (N_11322,N_9115,N_9141);
nor U11323 (N_11323,N_9586,N_8759);
nand U11324 (N_11324,N_8261,N_8156);
or U11325 (N_11325,N_9765,N_8995);
nand U11326 (N_11326,N_9935,N_9213);
and U11327 (N_11327,N_9275,N_8678);
nor U11328 (N_11328,N_9514,N_8102);
and U11329 (N_11329,N_9377,N_8586);
nor U11330 (N_11330,N_9349,N_8734);
or U11331 (N_11331,N_8865,N_8955);
xor U11332 (N_11332,N_9543,N_8537);
and U11333 (N_11333,N_9011,N_8448);
or U11334 (N_11334,N_8763,N_8602);
or U11335 (N_11335,N_9521,N_8744);
nand U11336 (N_11336,N_9269,N_8724);
nand U11337 (N_11337,N_8679,N_8081);
nand U11338 (N_11338,N_8807,N_9211);
and U11339 (N_11339,N_8605,N_9861);
nand U11340 (N_11340,N_9767,N_8004);
nor U11341 (N_11341,N_8601,N_9544);
xnor U11342 (N_11342,N_9177,N_8329);
or U11343 (N_11343,N_9192,N_9233);
or U11344 (N_11344,N_9227,N_9281);
and U11345 (N_11345,N_8435,N_8059);
nand U11346 (N_11346,N_9323,N_8099);
and U11347 (N_11347,N_9465,N_9894);
or U11348 (N_11348,N_9084,N_8336);
or U11349 (N_11349,N_9427,N_8022);
or U11350 (N_11350,N_9471,N_9900);
and U11351 (N_11351,N_9596,N_8534);
xor U11352 (N_11352,N_8118,N_9217);
and U11353 (N_11353,N_8564,N_9315);
nor U11354 (N_11354,N_9024,N_9886);
and U11355 (N_11355,N_8862,N_8246);
nor U11356 (N_11356,N_9810,N_8883);
nand U11357 (N_11357,N_8736,N_9317);
or U11358 (N_11358,N_9556,N_9909);
nor U11359 (N_11359,N_8501,N_8934);
nand U11360 (N_11360,N_9495,N_8185);
nor U11361 (N_11361,N_8337,N_9026);
xor U11362 (N_11362,N_8714,N_9383);
nor U11363 (N_11363,N_8360,N_8007);
nand U11364 (N_11364,N_9062,N_8266);
nor U11365 (N_11365,N_8345,N_9083);
nor U11366 (N_11366,N_8378,N_8367);
or U11367 (N_11367,N_8916,N_9795);
or U11368 (N_11368,N_8153,N_8764);
nand U11369 (N_11369,N_9205,N_9813);
xor U11370 (N_11370,N_8644,N_8740);
and U11371 (N_11371,N_9907,N_8212);
nor U11372 (N_11372,N_8407,N_8478);
and U11373 (N_11373,N_8895,N_8115);
or U11374 (N_11374,N_8975,N_8447);
and U11375 (N_11375,N_8704,N_8598);
nor U11376 (N_11376,N_9244,N_9353);
nand U11377 (N_11377,N_9490,N_9315);
or U11378 (N_11378,N_9020,N_9791);
or U11379 (N_11379,N_8570,N_9923);
or U11380 (N_11380,N_9128,N_9801);
or U11381 (N_11381,N_8420,N_8025);
nor U11382 (N_11382,N_9030,N_9267);
nand U11383 (N_11383,N_8422,N_8322);
and U11384 (N_11384,N_9071,N_8185);
or U11385 (N_11385,N_8329,N_9043);
or U11386 (N_11386,N_8669,N_8822);
nor U11387 (N_11387,N_8481,N_9886);
or U11388 (N_11388,N_8181,N_8250);
and U11389 (N_11389,N_8754,N_9284);
nand U11390 (N_11390,N_9522,N_8624);
xor U11391 (N_11391,N_9407,N_9830);
nor U11392 (N_11392,N_9360,N_9296);
nor U11393 (N_11393,N_9006,N_8311);
or U11394 (N_11394,N_9896,N_8154);
and U11395 (N_11395,N_8490,N_8637);
nand U11396 (N_11396,N_8045,N_9764);
nor U11397 (N_11397,N_9071,N_9831);
nor U11398 (N_11398,N_8653,N_8074);
or U11399 (N_11399,N_8396,N_8064);
and U11400 (N_11400,N_9665,N_8296);
and U11401 (N_11401,N_8686,N_9506);
and U11402 (N_11402,N_8373,N_9139);
nand U11403 (N_11403,N_8814,N_9655);
and U11404 (N_11404,N_9530,N_8349);
nor U11405 (N_11405,N_8153,N_8358);
or U11406 (N_11406,N_9397,N_8407);
or U11407 (N_11407,N_8601,N_9546);
xnor U11408 (N_11408,N_8650,N_9886);
and U11409 (N_11409,N_8001,N_9153);
or U11410 (N_11410,N_9062,N_8572);
nor U11411 (N_11411,N_8546,N_8116);
and U11412 (N_11412,N_8088,N_9319);
and U11413 (N_11413,N_9686,N_9324);
nor U11414 (N_11414,N_9306,N_8121);
and U11415 (N_11415,N_9366,N_9915);
or U11416 (N_11416,N_9094,N_8754);
and U11417 (N_11417,N_9669,N_8506);
and U11418 (N_11418,N_8622,N_8567);
xor U11419 (N_11419,N_9330,N_8142);
nor U11420 (N_11420,N_9572,N_9757);
xor U11421 (N_11421,N_9990,N_9631);
or U11422 (N_11422,N_9541,N_8231);
and U11423 (N_11423,N_8776,N_9148);
and U11424 (N_11424,N_9463,N_9648);
xor U11425 (N_11425,N_9564,N_8886);
and U11426 (N_11426,N_8268,N_9863);
nand U11427 (N_11427,N_8522,N_8660);
nor U11428 (N_11428,N_9228,N_8976);
and U11429 (N_11429,N_8784,N_9784);
or U11430 (N_11430,N_8931,N_8810);
nand U11431 (N_11431,N_9447,N_8068);
or U11432 (N_11432,N_9788,N_9370);
and U11433 (N_11433,N_8676,N_8550);
nor U11434 (N_11434,N_9932,N_8889);
nand U11435 (N_11435,N_9624,N_9436);
nand U11436 (N_11436,N_9139,N_9898);
nand U11437 (N_11437,N_8913,N_8098);
nand U11438 (N_11438,N_9105,N_9561);
nor U11439 (N_11439,N_8635,N_8212);
xor U11440 (N_11440,N_8081,N_9247);
nor U11441 (N_11441,N_9977,N_9631);
and U11442 (N_11442,N_8487,N_8254);
and U11443 (N_11443,N_8801,N_9905);
nand U11444 (N_11444,N_8692,N_8345);
and U11445 (N_11445,N_9565,N_9407);
xnor U11446 (N_11446,N_8313,N_9101);
xor U11447 (N_11447,N_8181,N_9217);
xor U11448 (N_11448,N_8034,N_9269);
and U11449 (N_11449,N_8416,N_9074);
and U11450 (N_11450,N_9339,N_8994);
nand U11451 (N_11451,N_8882,N_9015);
and U11452 (N_11452,N_8712,N_8009);
nor U11453 (N_11453,N_9308,N_9679);
or U11454 (N_11454,N_8469,N_9627);
nor U11455 (N_11455,N_9604,N_8760);
nand U11456 (N_11456,N_9516,N_9960);
or U11457 (N_11457,N_8367,N_9473);
nor U11458 (N_11458,N_8092,N_9034);
xnor U11459 (N_11459,N_9385,N_8973);
and U11460 (N_11460,N_8648,N_8190);
nor U11461 (N_11461,N_9476,N_8026);
nand U11462 (N_11462,N_9197,N_8062);
and U11463 (N_11463,N_9105,N_9896);
nand U11464 (N_11464,N_9170,N_9980);
or U11465 (N_11465,N_9389,N_9249);
or U11466 (N_11466,N_9154,N_9963);
or U11467 (N_11467,N_8853,N_8886);
or U11468 (N_11468,N_9334,N_9634);
nor U11469 (N_11469,N_8254,N_9450);
nor U11470 (N_11470,N_9235,N_8619);
and U11471 (N_11471,N_9930,N_8433);
nand U11472 (N_11472,N_8257,N_8607);
and U11473 (N_11473,N_8423,N_8929);
nor U11474 (N_11474,N_9614,N_9910);
and U11475 (N_11475,N_9894,N_8840);
or U11476 (N_11476,N_8451,N_9685);
or U11477 (N_11477,N_8995,N_9541);
nand U11478 (N_11478,N_8564,N_9130);
xor U11479 (N_11479,N_8796,N_8252);
nor U11480 (N_11480,N_9694,N_9996);
or U11481 (N_11481,N_8945,N_8582);
or U11482 (N_11482,N_8626,N_8861);
or U11483 (N_11483,N_8458,N_8435);
nor U11484 (N_11484,N_9598,N_9841);
nand U11485 (N_11485,N_8549,N_8552);
nor U11486 (N_11486,N_8423,N_8477);
xnor U11487 (N_11487,N_9463,N_8806);
nand U11488 (N_11488,N_9628,N_8534);
nor U11489 (N_11489,N_8825,N_9635);
nand U11490 (N_11490,N_8036,N_9907);
nand U11491 (N_11491,N_9042,N_9121);
nand U11492 (N_11492,N_9821,N_9915);
nor U11493 (N_11493,N_8449,N_9833);
nand U11494 (N_11494,N_9707,N_9868);
and U11495 (N_11495,N_9235,N_9803);
nor U11496 (N_11496,N_9786,N_8833);
nand U11497 (N_11497,N_8158,N_8038);
or U11498 (N_11498,N_9317,N_8766);
and U11499 (N_11499,N_9783,N_9871);
or U11500 (N_11500,N_8502,N_9095);
nand U11501 (N_11501,N_8037,N_8760);
or U11502 (N_11502,N_9679,N_9161);
xor U11503 (N_11503,N_9005,N_9887);
and U11504 (N_11504,N_8345,N_8239);
and U11505 (N_11505,N_8782,N_9769);
and U11506 (N_11506,N_8667,N_8405);
and U11507 (N_11507,N_9154,N_9417);
or U11508 (N_11508,N_8921,N_8840);
xnor U11509 (N_11509,N_8504,N_8268);
nand U11510 (N_11510,N_8101,N_8319);
nand U11511 (N_11511,N_9064,N_9861);
xnor U11512 (N_11512,N_9987,N_9535);
nor U11513 (N_11513,N_8533,N_9109);
and U11514 (N_11514,N_8060,N_9579);
nor U11515 (N_11515,N_9995,N_9487);
nor U11516 (N_11516,N_9184,N_8493);
and U11517 (N_11517,N_8363,N_8126);
nor U11518 (N_11518,N_9034,N_8830);
xor U11519 (N_11519,N_8115,N_9012);
nor U11520 (N_11520,N_8433,N_9001);
and U11521 (N_11521,N_9712,N_9279);
nand U11522 (N_11522,N_8764,N_9078);
and U11523 (N_11523,N_9604,N_9622);
nand U11524 (N_11524,N_9994,N_8494);
nor U11525 (N_11525,N_8030,N_8642);
nand U11526 (N_11526,N_8459,N_8193);
and U11527 (N_11527,N_8750,N_8827);
nand U11528 (N_11528,N_8616,N_9563);
or U11529 (N_11529,N_9840,N_9185);
and U11530 (N_11530,N_9531,N_9353);
nor U11531 (N_11531,N_8460,N_8747);
and U11532 (N_11532,N_9607,N_8810);
or U11533 (N_11533,N_9859,N_8787);
and U11534 (N_11534,N_8648,N_9394);
nand U11535 (N_11535,N_8494,N_9396);
nand U11536 (N_11536,N_8677,N_9096);
xnor U11537 (N_11537,N_8728,N_8190);
or U11538 (N_11538,N_8892,N_8675);
or U11539 (N_11539,N_9524,N_9140);
nor U11540 (N_11540,N_9178,N_8165);
or U11541 (N_11541,N_9556,N_8331);
nor U11542 (N_11542,N_8034,N_8161);
and U11543 (N_11543,N_8856,N_8584);
nor U11544 (N_11544,N_9818,N_9704);
and U11545 (N_11545,N_9567,N_9537);
nand U11546 (N_11546,N_8257,N_8138);
nand U11547 (N_11547,N_9042,N_8175);
nor U11548 (N_11548,N_9888,N_8799);
and U11549 (N_11549,N_8031,N_8172);
nand U11550 (N_11550,N_9622,N_8068);
nand U11551 (N_11551,N_9422,N_9967);
and U11552 (N_11552,N_9286,N_9007);
nor U11553 (N_11553,N_9660,N_9641);
nand U11554 (N_11554,N_8578,N_9281);
or U11555 (N_11555,N_8545,N_9770);
or U11556 (N_11556,N_8834,N_8577);
and U11557 (N_11557,N_8687,N_8576);
or U11558 (N_11558,N_8309,N_9055);
nand U11559 (N_11559,N_9799,N_9052);
or U11560 (N_11560,N_9342,N_8395);
and U11561 (N_11561,N_8089,N_9610);
nand U11562 (N_11562,N_8804,N_9708);
xnor U11563 (N_11563,N_9691,N_8958);
and U11564 (N_11564,N_8223,N_9294);
and U11565 (N_11565,N_8194,N_8873);
and U11566 (N_11566,N_8579,N_9773);
and U11567 (N_11567,N_8516,N_9835);
nand U11568 (N_11568,N_8455,N_8745);
and U11569 (N_11569,N_9262,N_9672);
and U11570 (N_11570,N_9175,N_8189);
nand U11571 (N_11571,N_9621,N_9106);
nor U11572 (N_11572,N_8166,N_8437);
nor U11573 (N_11573,N_8793,N_8627);
and U11574 (N_11574,N_8162,N_9435);
nor U11575 (N_11575,N_8323,N_8642);
and U11576 (N_11576,N_8388,N_8799);
or U11577 (N_11577,N_9701,N_9813);
xor U11578 (N_11578,N_9422,N_9108);
or U11579 (N_11579,N_8292,N_9512);
nor U11580 (N_11580,N_8635,N_9207);
xnor U11581 (N_11581,N_9456,N_8146);
nand U11582 (N_11582,N_8336,N_8748);
and U11583 (N_11583,N_8155,N_8931);
and U11584 (N_11584,N_8061,N_8773);
or U11585 (N_11585,N_8990,N_9645);
nor U11586 (N_11586,N_8646,N_9903);
nor U11587 (N_11587,N_8640,N_8448);
nand U11588 (N_11588,N_8321,N_9403);
nor U11589 (N_11589,N_8531,N_8322);
and U11590 (N_11590,N_9633,N_9480);
nand U11591 (N_11591,N_9736,N_9666);
nand U11592 (N_11592,N_9812,N_9776);
xor U11593 (N_11593,N_8715,N_8497);
nor U11594 (N_11594,N_8565,N_9747);
xnor U11595 (N_11595,N_9874,N_8501);
nor U11596 (N_11596,N_9588,N_9646);
and U11597 (N_11597,N_9020,N_9751);
or U11598 (N_11598,N_8704,N_8151);
xor U11599 (N_11599,N_9627,N_8691);
or U11600 (N_11600,N_8595,N_8189);
nand U11601 (N_11601,N_9379,N_9193);
and U11602 (N_11602,N_9042,N_8818);
nor U11603 (N_11603,N_8934,N_8874);
xor U11604 (N_11604,N_9201,N_9199);
nand U11605 (N_11605,N_8015,N_8800);
nand U11606 (N_11606,N_8082,N_8564);
and U11607 (N_11607,N_8127,N_9598);
and U11608 (N_11608,N_9235,N_8170);
xnor U11609 (N_11609,N_9618,N_9919);
or U11610 (N_11610,N_8184,N_9943);
and U11611 (N_11611,N_9622,N_9569);
nor U11612 (N_11612,N_9573,N_8508);
or U11613 (N_11613,N_9391,N_8116);
or U11614 (N_11614,N_8132,N_8319);
nand U11615 (N_11615,N_8293,N_8702);
nand U11616 (N_11616,N_9833,N_9847);
nand U11617 (N_11617,N_8959,N_8413);
nand U11618 (N_11618,N_8479,N_8857);
nor U11619 (N_11619,N_9642,N_9308);
nor U11620 (N_11620,N_9301,N_9530);
xor U11621 (N_11621,N_9175,N_9144);
and U11622 (N_11622,N_9152,N_8316);
and U11623 (N_11623,N_9734,N_8449);
or U11624 (N_11624,N_8941,N_9991);
and U11625 (N_11625,N_8333,N_8014);
nand U11626 (N_11626,N_9985,N_9341);
or U11627 (N_11627,N_8043,N_9587);
or U11628 (N_11628,N_9322,N_9988);
or U11629 (N_11629,N_9706,N_8626);
or U11630 (N_11630,N_9780,N_8612);
or U11631 (N_11631,N_8103,N_8712);
xnor U11632 (N_11632,N_9757,N_9402);
nand U11633 (N_11633,N_8894,N_8209);
or U11634 (N_11634,N_9282,N_9731);
nand U11635 (N_11635,N_8492,N_9868);
and U11636 (N_11636,N_8416,N_8296);
nor U11637 (N_11637,N_9177,N_8731);
and U11638 (N_11638,N_9065,N_8084);
xnor U11639 (N_11639,N_8772,N_9220);
nor U11640 (N_11640,N_8981,N_8087);
xnor U11641 (N_11641,N_9818,N_9504);
or U11642 (N_11642,N_9845,N_8722);
or U11643 (N_11643,N_9113,N_9906);
nand U11644 (N_11644,N_9493,N_9006);
nand U11645 (N_11645,N_9025,N_9877);
or U11646 (N_11646,N_9420,N_8050);
or U11647 (N_11647,N_8076,N_8206);
or U11648 (N_11648,N_9600,N_8890);
and U11649 (N_11649,N_9327,N_8457);
nand U11650 (N_11650,N_9255,N_9036);
nand U11651 (N_11651,N_8213,N_9490);
nand U11652 (N_11652,N_9901,N_8955);
or U11653 (N_11653,N_9798,N_8802);
or U11654 (N_11654,N_8013,N_9339);
or U11655 (N_11655,N_9922,N_9927);
and U11656 (N_11656,N_9620,N_9250);
nor U11657 (N_11657,N_9324,N_8680);
and U11658 (N_11658,N_8139,N_9560);
nor U11659 (N_11659,N_9336,N_8246);
nor U11660 (N_11660,N_8959,N_9192);
or U11661 (N_11661,N_9206,N_8586);
and U11662 (N_11662,N_9019,N_8871);
or U11663 (N_11663,N_8675,N_8900);
nor U11664 (N_11664,N_8842,N_8136);
or U11665 (N_11665,N_9949,N_9165);
nor U11666 (N_11666,N_8090,N_9643);
nor U11667 (N_11667,N_9642,N_8736);
and U11668 (N_11668,N_9269,N_9076);
nor U11669 (N_11669,N_8938,N_8288);
and U11670 (N_11670,N_9774,N_8918);
or U11671 (N_11671,N_8387,N_8808);
or U11672 (N_11672,N_9598,N_9387);
nand U11673 (N_11673,N_9069,N_8681);
or U11674 (N_11674,N_9637,N_9728);
or U11675 (N_11675,N_8698,N_8323);
and U11676 (N_11676,N_9410,N_8127);
and U11677 (N_11677,N_9721,N_9428);
nand U11678 (N_11678,N_9978,N_8351);
nand U11679 (N_11679,N_9257,N_9990);
or U11680 (N_11680,N_9075,N_8692);
nor U11681 (N_11681,N_9445,N_9878);
nor U11682 (N_11682,N_8838,N_9152);
and U11683 (N_11683,N_9392,N_8078);
nand U11684 (N_11684,N_8070,N_9670);
and U11685 (N_11685,N_8008,N_9938);
and U11686 (N_11686,N_9412,N_9058);
nand U11687 (N_11687,N_9281,N_9339);
nor U11688 (N_11688,N_9202,N_8699);
nor U11689 (N_11689,N_8949,N_8026);
and U11690 (N_11690,N_8929,N_9100);
xnor U11691 (N_11691,N_9835,N_9901);
nor U11692 (N_11692,N_8249,N_8675);
nor U11693 (N_11693,N_9565,N_9176);
nor U11694 (N_11694,N_9627,N_8827);
or U11695 (N_11695,N_8039,N_9885);
nand U11696 (N_11696,N_8635,N_9530);
xnor U11697 (N_11697,N_8236,N_9927);
and U11698 (N_11698,N_8113,N_8022);
and U11699 (N_11699,N_9582,N_9631);
nor U11700 (N_11700,N_8166,N_8749);
nor U11701 (N_11701,N_9885,N_9818);
or U11702 (N_11702,N_9679,N_8427);
nand U11703 (N_11703,N_9789,N_9267);
nand U11704 (N_11704,N_9875,N_8573);
or U11705 (N_11705,N_8479,N_9410);
or U11706 (N_11706,N_8919,N_8317);
nor U11707 (N_11707,N_8225,N_8373);
xnor U11708 (N_11708,N_8646,N_8354);
or U11709 (N_11709,N_8267,N_9094);
xor U11710 (N_11710,N_8963,N_8889);
or U11711 (N_11711,N_9199,N_9487);
nor U11712 (N_11712,N_8656,N_8784);
or U11713 (N_11713,N_8200,N_8874);
and U11714 (N_11714,N_8625,N_8246);
nor U11715 (N_11715,N_8060,N_9984);
nand U11716 (N_11716,N_9438,N_8819);
nor U11717 (N_11717,N_9729,N_9932);
and U11718 (N_11718,N_9149,N_9404);
nand U11719 (N_11719,N_8931,N_8776);
nand U11720 (N_11720,N_8196,N_8918);
or U11721 (N_11721,N_8444,N_9315);
xnor U11722 (N_11722,N_8311,N_9373);
nand U11723 (N_11723,N_8417,N_9549);
nand U11724 (N_11724,N_8416,N_8124);
nand U11725 (N_11725,N_9674,N_8068);
or U11726 (N_11726,N_8073,N_9814);
or U11727 (N_11727,N_9866,N_9796);
nor U11728 (N_11728,N_9805,N_8010);
nor U11729 (N_11729,N_9312,N_9078);
and U11730 (N_11730,N_9266,N_8443);
xor U11731 (N_11731,N_9949,N_9920);
or U11732 (N_11732,N_8541,N_9016);
or U11733 (N_11733,N_8546,N_8324);
or U11734 (N_11734,N_9288,N_8178);
and U11735 (N_11735,N_8210,N_9124);
nand U11736 (N_11736,N_8162,N_8107);
or U11737 (N_11737,N_9220,N_8710);
or U11738 (N_11738,N_8056,N_9672);
nand U11739 (N_11739,N_9589,N_9142);
and U11740 (N_11740,N_9827,N_8091);
or U11741 (N_11741,N_9706,N_9781);
nand U11742 (N_11742,N_9419,N_9695);
nand U11743 (N_11743,N_8521,N_8844);
nand U11744 (N_11744,N_9658,N_9096);
or U11745 (N_11745,N_8928,N_8776);
nand U11746 (N_11746,N_9459,N_9708);
nand U11747 (N_11747,N_9754,N_8657);
xnor U11748 (N_11748,N_9786,N_8187);
xnor U11749 (N_11749,N_8146,N_9103);
nand U11750 (N_11750,N_9618,N_9729);
nand U11751 (N_11751,N_9702,N_9556);
and U11752 (N_11752,N_8603,N_9450);
nor U11753 (N_11753,N_9325,N_8797);
or U11754 (N_11754,N_8063,N_8156);
nand U11755 (N_11755,N_9301,N_9439);
and U11756 (N_11756,N_8037,N_9443);
nand U11757 (N_11757,N_9379,N_8555);
or U11758 (N_11758,N_9207,N_8136);
nand U11759 (N_11759,N_9023,N_9297);
nand U11760 (N_11760,N_8744,N_9460);
nor U11761 (N_11761,N_9720,N_9445);
or U11762 (N_11762,N_8045,N_8933);
nor U11763 (N_11763,N_8506,N_8090);
and U11764 (N_11764,N_9285,N_9768);
or U11765 (N_11765,N_8047,N_8530);
nand U11766 (N_11766,N_8024,N_9230);
nor U11767 (N_11767,N_9985,N_8612);
nor U11768 (N_11768,N_9609,N_9735);
or U11769 (N_11769,N_8670,N_8399);
nor U11770 (N_11770,N_9003,N_8409);
and U11771 (N_11771,N_8079,N_8434);
nor U11772 (N_11772,N_8159,N_9800);
nor U11773 (N_11773,N_8311,N_9583);
nand U11774 (N_11774,N_9111,N_8760);
or U11775 (N_11775,N_8834,N_9930);
nor U11776 (N_11776,N_8448,N_8162);
or U11777 (N_11777,N_8420,N_9210);
and U11778 (N_11778,N_8660,N_9673);
nand U11779 (N_11779,N_9721,N_8480);
nand U11780 (N_11780,N_9410,N_8163);
xnor U11781 (N_11781,N_8512,N_8077);
nand U11782 (N_11782,N_9973,N_9960);
and U11783 (N_11783,N_8368,N_8659);
or U11784 (N_11784,N_9536,N_9858);
xor U11785 (N_11785,N_9917,N_8558);
nand U11786 (N_11786,N_9179,N_9947);
nand U11787 (N_11787,N_9672,N_9123);
xnor U11788 (N_11788,N_8182,N_8895);
and U11789 (N_11789,N_8248,N_8397);
nand U11790 (N_11790,N_8069,N_8058);
and U11791 (N_11791,N_8190,N_9660);
or U11792 (N_11792,N_8534,N_8625);
nand U11793 (N_11793,N_9164,N_9706);
and U11794 (N_11794,N_8264,N_8611);
nand U11795 (N_11795,N_8945,N_9467);
nand U11796 (N_11796,N_9122,N_8020);
and U11797 (N_11797,N_8211,N_9509);
or U11798 (N_11798,N_8048,N_9643);
or U11799 (N_11799,N_9190,N_8232);
or U11800 (N_11800,N_8868,N_9617);
nor U11801 (N_11801,N_8951,N_9401);
nor U11802 (N_11802,N_9700,N_8451);
nor U11803 (N_11803,N_9420,N_8154);
nor U11804 (N_11804,N_9456,N_8062);
nand U11805 (N_11805,N_8712,N_8750);
nor U11806 (N_11806,N_9530,N_9465);
or U11807 (N_11807,N_8249,N_8548);
or U11808 (N_11808,N_8620,N_9139);
xor U11809 (N_11809,N_8577,N_9058);
and U11810 (N_11810,N_8852,N_8183);
and U11811 (N_11811,N_9012,N_8452);
nand U11812 (N_11812,N_8107,N_9020);
nor U11813 (N_11813,N_9023,N_8796);
nand U11814 (N_11814,N_9660,N_8975);
nand U11815 (N_11815,N_9395,N_8300);
nor U11816 (N_11816,N_9378,N_9224);
nand U11817 (N_11817,N_9789,N_9208);
nor U11818 (N_11818,N_8745,N_8452);
nor U11819 (N_11819,N_9154,N_8817);
and U11820 (N_11820,N_9361,N_8280);
and U11821 (N_11821,N_9678,N_9175);
nand U11822 (N_11822,N_8171,N_8791);
and U11823 (N_11823,N_8334,N_9940);
nand U11824 (N_11824,N_8710,N_8302);
or U11825 (N_11825,N_9824,N_9370);
or U11826 (N_11826,N_9498,N_8409);
xor U11827 (N_11827,N_9095,N_9595);
and U11828 (N_11828,N_8648,N_9451);
xor U11829 (N_11829,N_9634,N_8936);
or U11830 (N_11830,N_9445,N_8574);
and U11831 (N_11831,N_9397,N_9172);
or U11832 (N_11832,N_8676,N_8418);
or U11833 (N_11833,N_8325,N_8775);
or U11834 (N_11834,N_8173,N_8736);
and U11835 (N_11835,N_8931,N_8383);
nand U11836 (N_11836,N_9705,N_8291);
or U11837 (N_11837,N_9232,N_9638);
nor U11838 (N_11838,N_9941,N_8236);
xor U11839 (N_11839,N_8716,N_8829);
nor U11840 (N_11840,N_8229,N_9533);
and U11841 (N_11841,N_9214,N_8230);
nor U11842 (N_11842,N_9783,N_9599);
or U11843 (N_11843,N_8306,N_9701);
nor U11844 (N_11844,N_9318,N_8836);
nor U11845 (N_11845,N_8128,N_9648);
xnor U11846 (N_11846,N_8486,N_9423);
and U11847 (N_11847,N_9116,N_8199);
nor U11848 (N_11848,N_9774,N_9304);
or U11849 (N_11849,N_8216,N_9548);
or U11850 (N_11850,N_8202,N_9244);
nand U11851 (N_11851,N_8869,N_8052);
and U11852 (N_11852,N_9139,N_9416);
and U11853 (N_11853,N_9092,N_8672);
or U11854 (N_11854,N_9628,N_9896);
nand U11855 (N_11855,N_8091,N_8621);
nor U11856 (N_11856,N_9565,N_8569);
xnor U11857 (N_11857,N_8335,N_9970);
nand U11858 (N_11858,N_8500,N_9358);
and U11859 (N_11859,N_9944,N_9764);
and U11860 (N_11860,N_8163,N_8358);
nor U11861 (N_11861,N_9836,N_8051);
nand U11862 (N_11862,N_8582,N_9475);
nor U11863 (N_11863,N_9698,N_8451);
nor U11864 (N_11864,N_9389,N_8509);
nor U11865 (N_11865,N_8669,N_8154);
nor U11866 (N_11866,N_8202,N_8242);
or U11867 (N_11867,N_9856,N_8117);
or U11868 (N_11868,N_9359,N_9052);
and U11869 (N_11869,N_9842,N_9532);
or U11870 (N_11870,N_8099,N_9911);
nor U11871 (N_11871,N_8107,N_9741);
or U11872 (N_11872,N_8676,N_8954);
and U11873 (N_11873,N_8375,N_8435);
xor U11874 (N_11874,N_9968,N_9120);
nand U11875 (N_11875,N_9315,N_8917);
nand U11876 (N_11876,N_9183,N_9862);
nand U11877 (N_11877,N_8000,N_9234);
nand U11878 (N_11878,N_9363,N_8663);
or U11879 (N_11879,N_9348,N_9745);
or U11880 (N_11880,N_8352,N_8527);
xor U11881 (N_11881,N_8365,N_9444);
xnor U11882 (N_11882,N_9127,N_8932);
and U11883 (N_11883,N_8624,N_9989);
nor U11884 (N_11884,N_8214,N_9526);
nor U11885 (N_11885,N_8884,N_8484);
nor U11886 (N_11886,N_9637,N_9247);
nand U11887 (N_11887,N_8532,N_9298);
and U11888 (N_11888,N_9857,N_8795);
or U11889 (N_11889,N_9179,N_9214);
nor U11890 (N_11890,N_8081,N_8670);
xor U11891 (N_11891,N_9569,N_8902);
or U11892 (N_11892,N_8379,N_8385);
nor U11893 (N_11893,N_9186,N_8092);
or U11894 (N_11894,N_8815,N_8748);
nor U11895 (N_11895,N_8434,N_9484);
or U11896 (N_11896,N_9626,N_9179);
xnor U11897 (N_11897,N_8999,N_8193);
and U11898 (N_11898,N_9989,N_9120);
nand U11899 (N_11899,N_9343,N_8057);
nand U11900 (N_11900,N_9412,N_9398);
nor U11901 (N_11901,N_9749,N_8694);
nor U11902 (N_11902,N_8630,N_8969);
or U11903 (N_11903,N_9765,N_9949);
nor U11904 (N_11904,N_8768,N_8685);
xor U11905 (N_11905,N_9908,N_9767);
nor U11906 (N_11906,N_8202,N_9006);
or U11907 (N_11907,N_8987,N_8635);
or U11908 (N_11908,N_9395,N_9563);
and U11909 (N_11909,N_9155,N_8952);
nor U11910 (N_11910,N_9853,N_8979);
nand U11911 (N_11911,N_8942,N_9802);
or U11912 (N_11912,N_8328,N_9125);
nand U11913 (N_11913,N_9064,N_9114);
or U11914 (N_11914,N_9381,N_9305);
nor U11915 (N_11915,N_9016,N_8800);
nand U11916 (N_11916,N_8972,N_9834);
nor U11917 (N_11917,N_8908,N_8127);
nor U11918 (N_11918,N_9101,N_8790);
nand U11919 (N_11919,N_9203,N_9902);
xor U11920 (N_11920,N_9344,N_8342);
nand U11921 (N_11921,N_8148,N_9895);
and U11922 (N_11922,N_9908,N_9179);
nor U11923 (N_11923,N_8977,N_8356);
or U11924 (N_11924,N_9500,N_8256);
xor U11925 (N_11925,N_8795,N_9795);
or U11926 (N_11926,N_9548,N_8424);
and U11927 (N_11927,N_8653,N_8433);
and U11928 (N_11928,N_9629,N_8209);
or U11929 (N_11929,N_8595,N_9767);
or U11930 (N_11930,N_9671,N_8108);
and U11931 (N_11931,N_8502,N_8442);
or U11932 (N_11932,N_9194,N_9080);
nor U11933 (N_11933,N_8098,N_9781);
and U11934 (N_11934,N_9306,N_8931);
nand U11935 (N_11935,N_9608,N_8795);
nand U11936 (N_11936,N_8871,N_9133);
or U11937 (N_11937,N_8864,N_8347);
nand U11938 (N_11938,N_8782,N_8513);
and U11939 (N_11939,N_9456,N_8156);
nor U11940 (N_11940,N_9152,N_8404);
or U11941 (N_11941,N_9916,N_9260);
nand U11942 (N_11942,N_8137,N_8963);
xor U11943 (N_11943,N_9293,N_9752);
xnor U11944 (N_11944,N_9845,N_9777);
and U11945 (N_11945,N_9294,N_8677);
xnor U11946 (N_11946,N_8341,N_8340);
nand U11947 (N_11947,N_9065,N_8074);
nor U11948 (N_11948,N_9678,N_8211);
nand U11949 (N_11949,N_8850,N_8924);
or U11950 (N_11950,N_9257,N_9143);
and U11951 (N_11951,N_9088,N_9648);
and U11952 (N_11952,N_9970,N_8747);
nand U11953 (N_11953,N_9545,N_9771);
xor U11954 (N_11954,N_8709,N_9478);
nor U11955 (N_11955,N_9038,N_9177);
nor U11956 (N_11956,N_9131,N_9713);
and U11957 (N_11957,N_9686,N_9718);
and U11958 (N_11958,N_8249,N_9685);
nand U11959 (N_11959,N_8651,N_9380);
nand U11960 (N_11960,N_9475,N_9141);
nor U11961 (N_11961,N_8090,N_8631);
xnor U11962 (N_11962,N_8853,N_8131);
nand U11963 (N_11963,N_9308,N_9511);
nor U11964 (N_11964,N_8089,N_8290);
xnor U11965 (N_11965,N_8001,N_8959);
nand U11966 (N_11966,N_9576,N_8750);
nand U11967 (N_11967,N_9966,N_9938);
or U11968 (N_11968,N_8590,N_9623);
nand U11969 (N_11969,N_8134,N_8679);
xnor U11970 (N_11970,N_9704,N_9595);
nand U11971 (N_11971,N_9302,N_9191);
nand U11972 (N_11972,N_8728,N_8750);
or U11973 (N_11973,N_8846,N_9011);
and U11974 (N_11974,N_8922,N_9021);
nand U11975 (N_11975,N_8620,N_9274);
and U11976 (N_11976,N_8179,N_9799);
nor U11977 (N_11977,N_8127,N_8640);
xor U11978 (N_11978,N_8100,N_9485);
or U11979 (N_11979,N_9106,N_9247);
nand U11980 (N_11980,N_9430,N_9949);
and U11981 (N_11981,N_8708,N_9606);
nor U11982 (N_11982,N_8457,N_9620);
and U11983 (N_11983,N_9453,N_9431);
xnor U11984 (N_11984,N_8802,N_8470);
xor U11985 (N_11985,N_9107,N_9904);
nand U11986 (N_11986,N_9847,N_8894);
nand U11987 (N_11987,N_9479,N_9273);
nor U11988 (N_11988,N_8391,N_8125);
xor U11989 (N_11989,N_8504,N_9482);
or U11990 (N_11990,N_9852,N_9593);
and U11991 (N_11991,N_9113,N_9004);
and U11992 (N_11992,N_9514,N_8930);
nor U11993 (N_11993,N_9073,N_8036);
nand U11994 (N_11994,N_9977,N_9983);
and U11995 (N_11995,N_9409,N_9057);
nand U11996 (N_11996,N_9550,N_9429);
and U11997 (N_11997,N_8888,N_9935);
or U11998 (N_11998,N_8763,N_9440);
nor U11999 (N_11999,N_9728,N_8742);
nor U12000 (N_12000,N_11242,N_11093);
and U12001 (N_12001,N_11855,N_11091);
or U12002 (N_12002,N_10523,N_11929);
nor U12003 (N_12003,N_10299,N_10019);
and U12004 (N_12004,N_11560,N_11489);
and U12005 (N_12005,N_10797,N_10823);
nor U12006 (N_12006,N_10511,N_10982);
nor U12007 (N_12007,N_10754,N_10188);
nor U12008 (N_12008,N_10879,N_11388);
xnor U12009 (N_12009,N_10300,N_11657);
nand U12010 (N_12010,N_10281,N_10762);
or U12011 (N_12011,N_11050,N_11038);
and U12012 (N_12012,N_10681,N_10286);
nor U12013 (N_12013,N_11908,N_10657);
nand U12014 (N_12014,N_10857,N_11613);
nor U12015 (N_12015,N_11788,N_11090);
nor U12016 (N_12016,N_10131,N_10859);
or U12017 (N_12017,N_10105,N_11956);
and U12018 (N_12018,N_10396,N_11431);
nand U12019 (N_12019,N_11060,N_10705);
xnor U12020 (N_12020,N_11025,N_10507);
nand U12021 (N_12021,N_10533,N_11372);
and U12022 (N_12022,N_10854,N_11684);
nand U12023 (N_12023,N_10592,N_10519);
xnor U12024 (N_12024,N_10684,N_10383);
and U12025 (N_12025,N_10626,N_10976);
nand U12026 (N_12026,N_10205,N_11963);
nand U12027 (N_12027,N_11408,N_11650);
xor U12028 (N_12028,N_10127,N_11449);
and U12029 (N_12029,N_10962,N_11339);
nor U12030 (N_12030,N_11151,N_11678);
nor U12031 (N_12031,N_11858,N_10183);
or U12032 (N_12032,N_11222,N_11728);
or U12033 (N_12033,N_10166,N_10469);
and U12034 (N_12034,N_11216,N_10891);
and U12035 (N_12035,N_10339,N_11481);
nor U12036 (N_12036,N_10306,N_10997);
nor U12037 (N_12037,N_11261,N_11535);
nand U12038 (N_12038,N_10654,N_11764);
and U12039 (N_12039,N_10191,N_11685);
and U12040 (N_12040,N_11354,N_11695);
and U12041 (N_12041,N_11348,N_10913);
and U12042 (N_12042,N_10027,N_11290);
or U12043 (N_12043,N_11513,N_11530);
nor U12044 (N_12044,N_11207,N_10426);
and U12045 (N_12045,N_10789,N_10922);
xnor U12046 (N_12046,N_10742,N_11832);
nor U12047 (N_12047,N_11082,N_11037);
xor U12048 (N_12048,N_11720,N_11971);
nor U12049 (N_12049,N_11053,N_10959);
and U12050 (N_12050,N_11759,N_11309);
and U12051 (N_12051,N_10569,N_11812);
nor U12052 (N_12052,N_10169,N_11308);
or U12053 (N_12053,N_11555,N_10370);
nand U12054 (N_12054,N_11406,N_11105);
nand U12055 (N_12055,N_11174,N_10835);
nor U12056 (N_12056,N_10757,N_11891);
or U12057 (N_12057,N_11487,N_11241);
and U12058 (N_12058,N_11572,N_11273);
xor U12059 (N_12059,N_10867,N_10101);
or U12060 (N_12060,N_11807,N_10672);
and U12061 (N_12061,N_10969,N_11023);
and U12062 (N_12062,N_10362,N_11141);
or U12063 (N_12063,N_10572,N_11550);
or U12064 (N_12064,N_11444,N_10830);
nor U12065 (N_12065,N_11604,N_11722);
and U12066 (N_12066,N_11860,N_10594);
and U12067 (N_12067,N_11588,N_10722);
and U12068 (N_12068,N_11006,N_10452);
nand U12069 (N_12069,N_11517,N_11991);
nand U12070 (N_12070,N_11785,N_10844);
xnor U12071 (N_12071,N_10294,N_10893);
and U12072 (N_12072,N_11413,N_10801);
nor U12073 (N_12073,N_11815,N_10025);
and U12074 (N_12074,N_10925,N_11122);
or U12075 (N_12075,N_11526,N_11959);
xor U12076 (N_12076,N_11341,N_10028);
nor U12077 (N_12077,N_11321,N_10768);
nor U12078 (N_12078,N_11218,N_10400);
or U12079 (N_12079,N_11169,N_10713);
nand U12080 (N_12080,N_11559,N_10630);
or U12081 (N_12081,N_10418,N_10571);
nor U12082 (N_12082,N_10087,N_11160);
or U12083 (N_12083,N_10590,N_10676);
nand U12084 (N_12084,N_11393,N_11987);
or U12085 (N_12085,N_11689,N_11292);
or U12086 (N_12086,N_11574,N_10735);
nand U12087 (N_12087,N_10750,N_11410);
nand U12088 (N_12088,N_11751,N_10556);
nand U12089 (N_12089,N_10391,N_11755);
nor U12090 (N_12090,N_11894,N_10054);
or U12091 (N_12091,N_11276,N_11178);
and U12092 (N_12092,N_10256,N_10435);
xnor U12093 (N_12093,N_10740,N_11827);
nand U12094 (N_12094,N_11916,N_10161);
or U12095 (N_12095,N_10202,N_11289);
nand U12096 (N_12096,N_10326,N_10449);
or U12097 (N_12097,N_10692,N_11671);
and U12098 (N_12098,N_11066,N_11663);
or U12099 (N_12099,N_10580,N_11236);
nor U12100 (N_12100,N_10352,N_10539);
or U12101 (N_12101,N_11801,N_11020);
nor U12102 (N_12102,N_10165,N_11012);
and U12103 (N_12103,N_11655,N_10344);
nand U12104 (N_12104,N_10864,N_10024);
nand U12105 (N_12105,N_11592,N_10049);
and U12106 (N_12106,N_10160,N_10777);
nand U12107 (N_12107,N_10275,N_10090);
nand U12108 (N_12108,N_10896,N_11412);
or U12109 (N_12109,N_10701,N_11317);
and U12110 (N_12110,N_11761,N_11601);
and U12111 (N_12111,N_10341,N_10374);
nor U12112 (N_12112,N_11948,N_11673);
nor U12113 (N_12113,N_11705,N_10515);
or U12114 (N_12114,N_11669,N_11735);
nor U12115 (N_12115,N_11727,N_10494);
nand U12116 (N_12116,N_11039,N_10671);
nor U12117 (N_12117,N_11584,N_11459);
nand U12118 (N_12118,N_11681,N_10910);
and U12119 (N_12119,N_11538,N_10960);
nor U12120 (N_12120,N_10586,N_10059);
and U12121 (N_12121,N_10051,N_10516);
nor U12122 (N_12122,N_11000,N_11575);
or U12123 (N_12123,N_10380,N_11201);
nor U12124 (N_12124,N_11153,N_10780);
and U12125 (N_12125,N_10399,N_10081);
xor U12126 (N_12126,N_11239,N_11131);
nand U12127 (N_12127,N_10625,N_10290);
nor U12128 (N_12128,N_10955,N_11647);
nor U12129 (N_12129,N_10669,N_11456);
nor U12130 (N_12130,N_10357,N_10497);
nand U12131 (N_12131,N_10634,N_10477);
or U12132 (N_12132,N_11355,N_10840);
or U12133 (N_12133,N_10337,N_10884);
or U12134 (N_12134,N_11437,N_10509);
nand U12135 (N_12135,N_10858,N_11223);
nand U12136 (N_12136,N_10582,N_11344);
xor U12137 (N_12137,N_11934,N_11464);
nor U12138 (N_12138,N_10407,N_10645);
nor U12139 (N_12139,N_11774,N_11072);
nand U12140 (N_12140,N_11175,N_10283);
nand U12141 (N_12141,N_10708,N_10086);
and U12142 (N_12142,N_11073,N_10624);
nor U12143 (N_12143,N_10904,N_10597);
or U12144 (N_12144,N_10150,N_11804);
and U12145 (N_12145,N_10929,N_11757);
or U12146 (N_12146,N_10030,N_11220);
or U12147 (N_12147,N_10679,N_11704);
and U12148 (N_12148,N_10318,N_10570);
nor U12149 (N_12149,N_11590,N_11612);
nor U12150 (N_12150,N_11307,N_10207);
nand U12151 (N_12151,N_10464,N_11899);
nor U12152 (N_12152,N_11300,N_10685);
nor U12153 (N_12153,N_10619,N_10486);
or U12154 (N_12154,N_11578,N_10832);
or U12155 (N_12155,N_10727,N_11277);
and U12156 (N_12156,N_10147,N_11966);
or U12157 (N_12157,N_10401,N_11362);
or U12158 (N_12158,N_11946,N_10782);
or U12159 (N_12159,N_10691,N_11244);
nor U12160 (N_12160,N_11754,N_10993);
and U12161 (N_12161,N_10136,N_10312);
and U12162 (N_12162,N_10375,N_11753);
or U12163 (N_12163,N_11779,N_10920);
xnor U12164 (N_12164,N_10239,N_11686);
nand U12165 (N_12165,N_11556,N_10791);
nand U12166 (N_12166,N_10089,N_10529);
and U12167 (N_12167,N_11896,N_10552);
nand U12168 (N_12168,N_10074,N_11096);
xnor U12169 (N_12169,N_11405,N_11425);
or U12170 (N_12170,N_11763,N_10898);
nand U12171 (N_12171,N_10513,N_10839);
nand U12172 (N_12172,N_10874,N_11134);
nor U12173 (N_12173,N_11429,N_10121);
xor U12174 (N_12174,N_11507,N_10588);
nand U12175 (N_12175,N_10083,N_10919);
nand U12176 (N_12176,N_11192,N_11340);
and U12177 (N_12177,N_10536,N_10114);
or U12178 (N_12178,N_10940,N_10044);
nand U12179 (N_12179,N_11052,N_10720);
nand U12180 (N_12180,N_10482,N_10700);
nor U12181 (N_12181,N_10765,N_11435);
or U12182 (N_12182,N_10408,N_10084);
nor U12183 (N_12183,N_10289,N_10875);
nor U12184 (N_12184,N_10741,N_11977);
and U12185 (N_12185,N_10650,N_10862);
nor U12186 (N_12186,N_10103,N_10208);
nor U12187 (N_12187,N_11204,N_10724);
nor U12188 (N_12188,N_11111,N_11798);
and U12189 (N_12189,N_11646,N_10377);
nor U12190 (N_12190,N_10259,N_10038);
nor U12191 (N_12191,N_10316,N_11250);
and U12192 (N_12192,N_10825,N_11842);
nand U12193 (N_12193,N_10887,N_11208);
or U12194 (N_12194,N_10524,N_10699);
and U12195 (N_12195,N_10404,N_11497);
or U12196 (N_12196,N_11397,N_10512);
or U12197 (N_12197,N_11295,N_10332);
nand U12198 (N_12198,N_10423,N_11771);
nor U12199 (N_12199,N_10313,N_10773);
nor U12200 (N_12200,N_10790,N_10829);
or U12201 (N_12201,N_11426,N_11453);
nor U12202 (N_12202,N_10865,N_10296);
nand U12203 (N_12203,N_11627,N_10379);
or U12204 (N_12204,N_10023,N_10770);
nand U12205 (N_12205,N_11994,N_11071);
and U12206 (N_12206,N_10719,N_10595);
xor U12207 (N_12207,N_10340,N_10579);
xor U12208 (N_12208,N_10055,N_11510);
and U12209 (N_12209,N_10753,N_10371);
nor U12210 (N_12210,N_11196,N_10113);
or U12211 (N_12211,N_10944,N_10468);
xnor U12212 (N_12212,N_11455,N_11599);
xnor U12213 (N_12213,N_10124,N_11126);
nand U12214 (N_12214,N_10022,N_10903);
and U12215 (N_12215,N_10682,N_11524);
nand U12216 (N_12216,N_11694,N_10419);
nor U12217 (N_12217,N_11452,N_10029);
or U12218 (N_12218,N_10437,N_10847);
nand U12219 (N_12219,N_11143,N_10834);
nor U12220 (N_12220,N_10409,N_11715);
xor U12221 (N_12221,N_11644,N_10334);
and U12222 (N_12222,N_10298,N_10227);
or U12223 (N_12223,N_11521,N_11389);
nor U12224 (N_12224,N_10032,N_11569);
and U12225 (N_12225,N_11664,N_10432);
or U12226 (N_12226,N_11005,N_10080);
and U12227 (N_12227,N_11205,N_11494);
nand U12228 (N_12228,N_11373,N_10343);
nor U12229 (N_12229,N_10557,N_10703);
nor U12230 (N_12230,N_11427,N_11214);
nor U12231 (N_12231,N_10881,N_10013);
or U12232 (N_12232,N_10309,N_11514);
or U12233 (N_12233,N_11128,N_11619);
or U12234 (N_12234,N_11856,N_10336);
or U12235 (N_12235,N_11306,N_11029);
or U12236 (N_12236,N_11527,N_10238);
or U12237 (N_12237,N_10690,N_11632);
nand U12238 (N_12238,N_10510,N_11329);
or U12239 (N_12239,N_10333,N_10082);
nand U12240 (N_12240,N_11747,N_11607);
and U12241 (N_12241,N_11256,N_11132);
or U12242 (N_12242,N_11358,N_11305);
or U12243 (N_12243,N_11215,N_10430);
nor U12244 (N_12244,N_11106,N_10346);
nand U12245 (N_12245,N_11401,N_11395);
nand U12246 (N_12246,N_10350,N_11182);
or U12247 (N_12247,N_11819,N_10984);
xor U12248 (N_12248,N_11721,N_11528);
or U12249 (N_12249,N_10849,N_11904);
xor U12250 (N_12250,N_11921,N_11769);
nor U12251 (N_12251,N_11600,N_10545);
nor U12252 (N_12252,N_10304,N_10226);
nand U12253 (N_12253,N_10577,N_11017);
xor U12254 (N_12254,N_10048,N_11936);
or U12255 (N_12255,N_11149,N_11648);
and U12256 (N_12256,N_10267,N_10220);
nor U12257 (N_12257,N_11442,N_11279);
xnor U12258 (N_12258,N_11187,N_11964);
and U12259 (N_12259,N_11396,N_11782);
nand U12260 (N_12260,N_11716,N_10810);
and U12261 (N_12261,N_10912,N_10584);
xor U12262 (N_12262,N_11176,N_11859);
or U12263 (N_12263,N_11076,N_11784);
xor U12264 (N_12264,N_10675,N_11291);
and U12265 (N_12265,N_10195,N_10627);
nand U12266 (N_12266,N_11707,N_10821);
or U12267 (N_12267,N_10598,N_10585);
nor U12268 (N_12268,N_10623,N_11152);
nor U12269 (N_12269,N_11806,N_11974);
and U12270 (N_12270,N_11548,N_11184);
nor U12271 (N_12271,N_11033,N_11359);
or U12272 (N_12272,N_11258,N_11047);
nand U12273 (N_12273,N_11577,N_10359);
nand U12274 (N_12274,N_11928,N_10674);
nand U12275 (N_12275,N_10637,N_11675);
nand U12276 (N_12276,N_11432,N_11976);
xor U12277 (N_12277,N_10167,N_11310);
nand U12278 (N_12278,N_11474,N_10269);
nor U12279 (N_12279,N_10097,N_10020);
or U12280 (N_12280,N_11349,N_11316);
and U12281 (N_12281,N_10402,N_11700);
nand U12282 (N_12282,N_10123,N_11089);
or U12283 (N_12283,N_10353,N_10758);
and U12284 (N_12284,N_10365,N_11377);
or U12285 (N_12285,N_10521,N_10258);
nor U12286 (N_12286,N_11995,N_11366);
and U12287 (N_12287,N_11793,N_11156);
and U12288 (N_12288,N_10071,N_10604);
or U12289 (N_12289,N_11210,N_10983);
and U12290 (N_12290,N_10179,N_11014);
and U12291 (N_12291,N_10855,N_10144);
and U12292 (N_12292,N_11498,N_10924);
xnor U12293 (N_12293,N_10643,N_10268);
nand U12294 (N_12294,N_11299,N_10172);
nand U12295 (N_12295,N_11937,N_11888);
or U12296 (N_12296,N_10039,N_11044);
nand U12297 (N_12297,N_10870,N_10905);
nor U12298 (N_12298,N_10567,N_11056);
nor U12299 (N_12299,N_11814,N_10366);
and U12300 (N_12300,N_10171,N_11233);
and U12301 (N_12301,N_11630,N_10257);
nand U12302 (N_12302,N_11315,N_10991);
nor U12303 (N_12303,N_11835,N_10246);
and U12304 (N_12304,N_11084,N_10528);
or U12305 (N_12305,N_11123,N_10841);
nand U12306 (N_12306,N_11749,N_11197);
and U12307 (N_12307,N_10527,N_10743);
or U12308 (N_12308,N_10249,N_11752);
xnor U12309 (N_12309,N_11980,N_10118);
or U12310 (N_12310,N_11235,N_11267);
nor U12311 (N_12311,N_10578,N_11616);
xor U12312 (N_12312,N_11202,N_11119);
and U12313 (N_12313,N_10827,N_11424);
xnor U12314 (N_12314,N_10351,N_10961);
xnor U12315 (N_12315,N_11463,N_10210);
nand U12316 (N_12316,N_10058,N_11311);
nor U12317 (N_12317,N_10878,N_10649);
or U12318 (N_12318,N_11330,N_11108);
nor U12319 (N_12319,N_10759,N_10731);
and U12320 (N_12320,N_10695,N_11731);
nor U12321 (N_12321,N_11733,N_10236);
and U12322 (N_12322,N_10093,N_11159);
nand U12323 (N_12323,N_10831,N_10868);
nand U12324 (N_12324,N_11077,N_11150);
nor U12325 (N_12325,N_10125,N_10219);
or U12326 (N_12326,N_11003,N_11505);
and U12327 (N_12327,N_10617,N_10693);
nor U12328 (N_12328,N_10706,N_11826);
or U12329 (N_12329,N_10367,N_11623);
or U12330 (N_12330,N_10481,N_11110);
nand U12331 (N_12331,N_10499,N_10621);
and U12332 (N_12332,N_10242,N_10522);
and U12333 (N_12333,N_10288,N_10551);
or U12334 (N_12334,N_11737,N_10788);
nand U12335 (N_12335,N_10576,N_11611);
and U12336 (N_12336,N_11048,N_11462);
xor U12337 (N_12337,N_10369,N_11129);
nand U12338 (N_12338,N_10095,N_11515);
and U12339 (N_12339,N_11996,N_10804);
nand U12340 (N_12340,N_10185,N_11209);
and U12341 (N_12341,N_10263,N_11387);
and U12342 (N_12342,N_10558,N_11167);
nor U12343 (N_12343,N_11802,N_11661);
nor U12344 (N_12344,N_11847,N_10541);
or U12345 (N_12345,N_11817,N_10253);
or U12346 (N_12346,N_11732,N_10361);
or U12347 (N_12347,N_11007,N_10411);
nand U12348 (N_12348,N_10007,N_10687);
xnor U12349 (N_12349,N_10382,N_11165);
and U12350 (N_12350,N_11911,N_10614);
or U12351 (N_12351,N_10434,N_11058);
and U12352 (N_12352,N_11190,N_11602);
and U12353 (N_12353,N_10968,N_10808);
nor U12354 (N_12354,N_10096,N_11629);
or U12355 (N_12355,N_10311,N_11672);
nor U12356 (N_12356,N_11186,N_10378);
xor U12357 (N_12357,N_11844,N_10769);
nand U12358 (N_12358,N_10270,N_11490);
nand U12359 (N_12359,N_10518,N_11869);
and U12360 (N_12360,N_11975,N_10974);
nor U12361 (N_12361,N_11351,N_10548);
nand U12362 (N_12362,N_10661,N_10648);
or U12363 (N_12363,N_10110,N_11484);
nand U12364 (N_12364,N_11376,N_10153);
xor U12365 (N_12365,N_10342,N_11512);
and U12366 (N_12366,N_11617,N_10457);
and U12367 (N_12367,N_11703,N_11533);
nand U12368 (N_12368,N_10421,N_10941);
and U12369 (N_12369,N_10662,N_11579);
nor U12370 (N_12370,N_10152,N_11252);
and U12371 (N_12371,N_10806,N_11713);
nand U12372 (N_12372,N_11953,N_11508);
or U12373 (N_12373,N_10099,N_11845);
and U12374 (N_12374,N_10534,N_11944);
nor U12375 (N_12375,N_11460,N_10129);
and U12376 (N_12376,N_11016,N_11138);
and U12377 (N_12377,N_11065,N_10349);
nand U12378 (N_12378,N_10209,N_10372);
nand U12379 (N_12379,N_11320,N_11420);
and U12380 (N_12380,N_10601,N_10602);
nor U12381 (N_12381,N_11880,N_11714);
xor U12382 (N_12382,N_10668,N_11285);
nand U12383 (N_12383,N_11443,N_11046);
and U12384 (N_12384,N_11097,N_10031);
nor U12385 (N_12385,N_10502,N_11822);
or U12386 (N_12386,N_11766,N_10363);
nand U12387 (N_12387,N_11098,N_10995);
or U12388 (N_12388,N_10888,N_11898);
nand U12389 (N_12389,N_11799,N_11158);
or U12390 (N_12390,N_11568,N_11967);
nand U12391 (N_12391,N_10139,N_11796);
nor U12392 (N_12392,N_11853,N_10838);
and U12393 (N_12393,N_10321,N_11969);
and U12394 (N_12394,N_10673,N_11718);
and U12395 (N_12395,N_10658,N_11691);
or U12396 (N_12396,N_10193,N_10730);
or U12397 (N_12397,N_11841,N_11502);
xnor U12398 (N_12398,N_11773,N_11368);
or U12399 (N_12399,N_11837,N_10215);
or U12400 (N_12400,N_10424,N_11386);
and U12401 (N_12401,N_11392,N_11537);
xor U12402 (N_12402,N_11544,N_11297);
or U12403 (N_12403,N_11876,N_11177);
nor U12404 (N_12404,N_11318,N_10412);
or U12405 (N_12405,N_11608,N_11570);
or U12406 (N_12406,N_11166,N_10799);
and U12407 (N_12407,N_10729,N_11545);
or U12408 (N_12408,N_10948,N_11962);
and U12409 (N_12409,N_10140,N_11468);
xnor U12410 (N_12410,N_10917,N_11595);
and U12411 (N_12411,N_10926,N_11935);
and U12412 (N_12412,N_10135,N_10973);
and U12413 (N_12413,N_11461,N_11683);
or U12414 (N_12414,N_11411,N_11283);
or U12415 (N_12415,N_10532,N_11659);
nand U12416 (N_12416,N_11760,N_10989);
nor U12417 (N_12417,N_10772,N_11852);
and U12418 (N_12418,N_10264,N_10711);
xor U12419 (N_12419,N_11631,N_11229);
nor U12420 (N_12420,N_11345,N_10237);
and U12421 (N_12421,N_11818,N_11246);
or U12422 (N_12422,N_11055,N_11002);
xnor U12423 (N_12423,N_11088,N_11193);
xnor U12424 (N_12424,N_10608,N_10873);
and U12425 (N_12425,N_10324,N_10501);
nand U12426 (N_12426,N_10970,N_11848);
and U12427 (N_12427,N_11925,N_10653);
nand U12428 (N_12428,N_11428,N_11225);
xor U12429 (N_12429,N_11251,N_10683);
nand U12430 (N_12430,N_10384,N_11902);
and U12431 (N_12431,N_10760,N_10323);
and U12432 (N_12432,N_11857,N_11907);
or U12433 (N_12433,N_11085,N_10128);
or U12434 (N_12434,N_11866,N_11473);
nor U12435 (N_12435,N_10106,N_11451);
or U12436 (N_12436,N_10328,N_10639);
nor U12437 (N_12437,N_11228,N_11580);
nor U12438 (N_12438,N_11940,N_11624);
xnor U12439 (N_12439,N_11115,N_10999);
or U12440 (N_12440,N_11206,N_10416);
or U12441 (N_12441,N_10543,N_11999);
or U12442 (N_12442,N_11506,N_11677);
or U12443 (N_12443,N_11816,N_10491);
nand U12444 (N_12444,N_10307,N_10120);
nand U12445 (N_12445,N_11360,N_10260);
and U12446 (N_12446,N_11838,N_11370);
nor U12447 (N_12447,N_10189,N_10222);
nor U12448 (N_12448,N_11958,N_11711);
and U12449 (N_12449,N_10927,N_11864);
nor U12450 (N_12450,N_10479,N_10145);
or U12451 (N_12451,N_11712,N_10981);
and U12452 (N_12452,N_10109,N_10301);
nand U12453 (N_12453,N_11952,N_11850);
or U12454 (N_12454,N_11063,N_11271);
xor U12455 (N_12455,N_10748,N_10764);
nor U12456 (N_12456,N_10117,N_11062);
xnor U12457 (N_12457,N_10410,N_11022);
nand U12458 (N_12458,N_10141,N_11419);
nor U12459 (N_12459,N_10656,N_10302);
nor U12460 (N_12460,N_10072,N_11674);
nor U12461 (N_12461,N_10142,N_10148);
nor U12462 (N_12462,N_11043,N_11811);
nor U12463 (N_12463,N_10800,N_10663);
xnor U12464 (N_12464,N_10815,N_10725);
nor U12465 (N_12465,N_11547,N_10229);
nor U12466 (N_12466,N_10037,N_10204);
xor U12467 (N_12467,N_10021,N_10733);
nand U12468 (N_12468,N_11791,N_10364);
and U12469 (N_12469,N_10348,N_11069);
nor U12470 (N_12470,N_11399,N_10231);
and U12471 (N_12471,N_11924,N_10317);
nand U12472 (N_12472,N_10641,N_10394);
or U12473 (N_12473,N_10980,N_10698);
nor U12474 (N_12474,N_10073,N_10012);
or U12475 (N_12475,N_11148,N_10493);
and U12476 (N_12476,N_10894,N_11203);
or U12477 (N_12477,N_11238,N_10694);
xnor U12478 (N_12478,N_10882,N_11185);
xor U12479 (N_12479,N_10274,N_10498);
nand U12480 (N_12480,N_10633,N_10480);
nor U12481 (N_12481,N_11031,N_10549);
and U12482 (N_12482,N_11334,N_10575);
nor U12483 (N_12483,N_11906,N_11180);
xnor U12484 (N_12484,N_11790,N_11313);
or U12485 (N_12485,N_10064,N_11918);
or U12486 (N_12486,N_10992,N_11019);
nand U12487 (N_12487,N_10395,N_10453);
nand U12488 (N_12488,N_10990,N_10848);
nor U12489 (N_12489,N_10589,N_10736);
xor U12490 (N_12490,N_11171,N_11163);
or U12491 (N_12491,N_10420,N_10943);
nand U12492 (N_12492,N_10547,N_11622);
or U12493 (N_12493,N_11116,N_11482);
or U12494 (N_12494,N_10303,N_11384);
nand U12495 (N_12495,N_11080,N_11380);
or U12496 (N_12496,N_11941,N_10415);
nor U12497 (N_12497,N_10360,N_10355);
xnor U12498 (N_12498,N_11518,N_10285);
xnor U12499 (N_12499,N_11516,N_11625);
or U12500 (N_12500,N_11536,N_10609);
xnor U12501 (N_12501,N_10537,N_10387);
nor U12502 (N_12502,N_11100,N_11418);
nand U12503 (N_12503,N_11319,N_11083);
and U12504 (N_12504,N_10642,N_10986);
and U12505 (N_12505,N_11543,N_10755);
nor U12506 (N_12506,N_10062,N_11421);
nand U12507 (N_12507,N_11563,N_10473);
nand U12508 (N_12508,N_10240,N_10795);
or U12509 (N_12509,N_10282,N_10902);
and U12510 (N_12510,N_10738,N_11912);
nand U12511 (N_12511,N_11746,N_10385);
and U12512 (N_12512,N_10972,N_11724);
or U12513 (N_12513,N_10130,N_10756);
xnor U12514 (N_12514,N_11287,N_10890);
nand U12515 (N_12515,N_10386,N_10255);
and U12516 (N_12516,N_11219,N_10812);
and U12517 (N_12517,N_11667,N_11662);
nand U12518 (N_12518,N_10816,N_11154);
nor U12519 (N_12519,N_10824,N_11326);
and U12520 (N_12520,N_11092,N_10373);
and U12521 (N_12521,N_11051,N_10600);
nor U12522 (N_12522,N_10988,N_11087);
nand U12523 (N_12523,N_11541,N_11145);
and U12524 (N_12524,N_11028,N_10003);
nor U12525 (N_12525,N_11382,N_10016);
and U12526 (N_12526,N_10503,N_11628);
nor U12527 (N_12527,N_11394,N_10798);
and U12528 (N_12528,N_10817,N_10544);
nor U12529 (N_12529,N_11332,N_11554);
nor U12530 (N_12530,N_10718,N_11933);
nand U12531 (N_12531,N_10381,N_11834);
nand U12532 (N_12532,N_10554,N_11939);
or U12533 (N_12533,N_11364,N_10077);
or U12534 (N_12534,N_10964,N_10900);
and U12535 (N_12535,N_11270,N_11978);
or U12536 (N_12536,N_11404,N_11440);
or U12537 (N_12537,N_11454,N_10949);
nand U12538 (N_12538,N_10175,N_11409);
nor U12539 (N_12539,N_11086,N_10715);
nor U12540 (N_12540,N_11610,N_10248);
and U12541 (N_12541,N_10149,N_10194);
xnor U12542 (N_12542,N_11057,N_10428);
nor U12543 (N_12543,N_11068,N_10937);
nand U12544 (N_12544,N_10843,N_10112);
xnor U12545 (N_12545,N_10462,N_10895);
xor U12546 (N_12546,N_11476,N_10425);
xor U12547 (N_12547,N_10433,N_10471);
or U12548 (N_12548,N_11895,N_10247);
or U12549 (N_12549,N_11736,N_11905);
nor U12550 (N_12550,N_10047,N_10610);
and U12551 (N_12551,N_10809,N_11532);
and U12552 (N_12552,N_10635,N_11865);
nor U12553 (N_12553,N_11079,N_10198);
and U12554 (N_12554,N_11130,N_10901);
and U12555 (N_12555,N_11447,N_10506);
and U12556 (N_12556,N_11227,N_11155);
or U12557 (N_12557,N_11803,N_11640);
nor U12558 (N_12558,N_10892,N_10035);
and U12559 (N_12559,N_11993,N_11765);
nor U12560 (N_12560,N_10233,N_11240);
nand U12561 (N_12561,N_11945,N_11275);
and U12562 (N_12562,N_11884,N_11194);
nor U12563 (N_12563,N_11820,N_10292);
or U12564 (N_12564,N_11293,N_11810);
xor U12565 (N_12565,N_10459,N_10555);
nand U12566 (N_12566,N_11660,N_10390);
nand U12567 (N_12567,N_10241,N_11795);
or U12568 (N_12568,N_10587,N_11531);
nand U12569 (N_12569,N_10448,N_11217);
or U12570 (N_12570,N_11162,N_11036);
xnor U12571 (N_12571,N_10566,N_11257);
or U12572 (N_12572,N_10444,N_11676);
or U12573 (N_12573,N_10603,N_10043);
and U12574 (N_12574,N_11565,N_10538);
nor U12575 (N_12575,N_10465,N_11915);
and U12576 (N_12576,N_11571,N_10245);
or U12577 (N_12577,N_11558,N_10442);
or U12578 (N_12578,N_10751,N_11402);
xor U12579 (N_12579,N_11259,N_10975);
nand U12580 (N_12580,N_11018,N_11525);
nor U12581 (N_12581,N_10230,N_10611);
and U12582 (N_12582,N_11890,N_11961);
nor U12583 (N_12583,N_10775,N_10098);
or U12584 (N_12584,N_10476,N_11979);
xnor U12585 (N_12585,N_11423,N_11873);
xnor U12586 (N_12586,N_11789,N_10934);
xor U12587 (N_12587,N_11248,N_11998);
and U12588 (N_12588,N_10413,N_10792);
and U12589 (N_12589,N_10445,N_11247);
or U12590 (N_12590,N_11523,N_11709);
nand U12591 (N_12591,N_11726,N_10162);
or U12592 (N_12592,N_10060,N_10911);
and U12593 (N_12593,N_10484,N_11133);
nor U12594 (N_12594,N_10935,N_11539);
xor U12595 (N_12595,N_10945,N_10327);
and U12596 (N_12596,N_10787,N_11030);
xor U12597 (N_12597,N_11337,N_10042);
or U12598 (N_12598,N_10261,N_11074);
or U12599 (N_12599,N_11112,N_11263);
or U12600 (N_12600,N_11540,N_10947);
nor U12601 (N_12601,N_11226,N_10763);
nor U12602 (N_12602,N_10803,N_11943);
nor U12603 (N_12603,N_10151,N_11298);
or U12604 (N_12604,N_11723,N_10392);
nand U12605 (N_12605,N_10591,N_10217);
and U12606 (N_12606,N_11139,N_11549);
xor U12607 (N_12607,N_10581,N_10977);
nor U12608 (N_12608,N_11621,N_10192);
or U12609 (N_12609,N_11626,N_10406);
or U12610 (N_12610,N_10779,N_11797);
nor U12611 (N_12611,N_10956,N_11181);
nor U12612 (N_12612,N_10613,N_10243);
nor U12613 (N_12613,N_11519,N_11231);
nand U12614 (N_12614,N_11212,N_11363);
xor U12615 (N_12615,N_10950,N_11687);
nand U12616 (N_12616,N_11434,N_11323);
nor U12617 (N_12617,N_10017,N_10397);
nand U12618 (N_12618,N_10707,N_11288);
nor U12619 (N_12619,N_10046,N_10001);
xor U12620 (N_12620,N_10771,N_10811);
nand U12621 (N_12621,N_11741,N_11479);
and U12622 (N_12622,N_10265,N_10813);
nor U12623 (N_12623,N_10146,N_11829);
or U12624 (N_12624,N_10200,N_10646);
or U12625 (N_12625,N_11234,N_11189);
nor U12626 (N_12626,N_10774,N_11897);
nor U12627 (N_12627,N_11142,N_11059);
nand U12628 (N_12628,N_11777,N_11679);
nor U12629 (N_12629,N_11942,N_11243);
and U12630 (N_12630,N_11809,N_10137);
or U12631 (N_12631,N_11839,N_10115);
nor U12632 (N_12632,N_11828,N_10271);
or U12633 (N_12633,N_11775,N_11213);
and U12634 (N_12634,N_11170,N_11794);
or U12635 (N_12635,N_11919,N_11534);
or U12636 (N_12636,N_11436,N_11808);
or U12637 (N_12637,N_10008,N_10889);
or U12638 (N_12638,N_10796,N_10504);
nor U12639 (N_12639,N_11830,N_11583);
nand U12640 (N_12640,N_10869,N_10347);
and U12641 (N_12641,N_10918,N_10936);
xnor U12642 (N_12642,N_11407,N_11322);
xnor U12643 (N_12643,N_10186,N_11094);
or U12644 (N_12644,N_11179,N_10427);
nor U12645 (N_12645,N_11356,N_10886);
and U12646 (N_12646,N_11325,N_10856);
and U12647 (N_12647,N_11347,N_11950);
and U12648 (N_12648,N_10996,N_11649);
and U12649 (N_12649,N_10173,N_10000);
and U12650 (N_12650,N_11034,N_10710);
or U12651 (N_12651,N_10659,N_11103);
nand U12652 (N_12652,N_11265,N_10784);
or U12653 (N_12653,N_11889,N_10853);
and U12654 (N_12654,N_10436,N_10102);
and U12655 (N_12655,N_10957,N_11433);
or U12656 (N_12656,N_11562,N_11717);
and U12657 (N_12657,N_10712,N_10517);
or U12658 (N_12658,N_10052,N_11740);
nor U12659 (N_12659,N_11743,N_10004);
and U12660 (N_12660,N_11886,N_11118);
or U12661 (N_12661,N_10234,N_11938);
nor U12662 (N_12662,N_10607,N_11268);
nor U12663 (N_12663,N_10250,N_10747);
and U12664 (N_12664,N_11863,N_10987);
or U12665 (N_12665,N_11652,N_10485);
and U12666 (N_12666,N_10907,N_10266);
nand U12667 (N_12667,N_11872,N_11883);
or U12668 (N_12668,N_10915,N_11027);
or U12669 (N_12669,N_10201,N_11417);
nor U12670 (N_12670,N_11493,N_10164);
or U12671 (N_12671,N_11744,N_10100);
and U12672 (N_12672,N_11472,N_10388);
nand U12673 (N_12673,N_11614,N_10376);
xor U12674 (N_12674,N_10006,N_10315);
or U12675 (N_12675,N_11157,N_11104);
nor U12676 (N_12676,N_11414,N_10085);
nor U12677 (N_12677,N_11296,N_10820);
or U12678 (N_12678,N_10168,N_11557);
nor U12679 (N_12679,N_11328,N_11121);
nand U12680 (N_12680,N_11843,N_11109);
nor U12681 (N_12681,N_10156,N_11573);
nor U12682 (N_12682,N_11706,N_10057);
nor U12683 (N_12683,N_10923,N_11985);
nand U12684 (N_12684,N_11144,N_10026);
and U12685 (N_12685,N_10015,N_11781);
nor U12686 (N_12686,N_10599,N_11172);
and U12687 (N_12687,N_10079,N_11221);
or U12688 (N_12688,N_11361,N_10472);
and U12689 (N_12689,N_10794,N_11970);
nand U12690 (N_12690,N_10273,N_11913);
nor U12691 (N_12691,N_10852,N_10221);
nand U12692 (N_12692,N_10930,N_10647);
nor U12693 (N_12693,N_11107,N_10319);
or U12694 (N_12694,N_11787,N_10651);
or U12695 (N_12695,N_11988,N_10688);
and U12696 (N_12696,N_10574,N_11255);
nand U12697 (N_12697,N_10414,N_10967);
nand U12698 (N_12698,N_10846,N_10050);
and U12699 (N_12699,N_11824,N_11078);
and U12700 (N_12700,N_11719,N_10966);
xor U12701 (N_12701,N_10908,N_10190);
and U12702 (N_12702,N_11992,N_10478);
nand U12703 (N_12703,N_10492,N_11303);
nand U12704 (N_12704,N_11585,N_11237);
nor U12705 (N_12705,N_10914,N_10429);
nand U12706 (N_12706,N_10931,N_10837);
nor U12707 (N_12707,N_11920,N_10180);
xor U12708 (N_12708,N_11688,N_11725);
and U12709 (N_12709,N_10065,N_10631);
or U12710 (N_12710,N_10439,N_10063);
nand U12711 (N_12711,N_10573,N_10877);
and U12712 (N_12712,N_11164,N_10778);
and U12713 (N_12713,N_11441,N_11643);
or U12714 (N_12714,N_11471,N_11013);
nor U12715 (N_12715,N_11874,N_10487);
and U12716 (N_12716,N_11114,N_11639);
and U12717 (N_12717,N_11117,N_11365);
nor U12718 (N_12718,N_10203,N_10540);
xnor U12719 (N_12719,N_11520,N_10583);
nand U12720 (N_12720,N_10897,N_10330);
and U12721 (N_12721,N_10196,N_10978);
nor U12722 (N_12722,N_10354,N_10612);
nor U12723 (N_12723,N_10356,N_10746);
nor U12724 (N_12724,N_10716,N_11870);
and U12725 (N_12725,N_11338,N_11477);
nor U12726 (N_12726,N_10542,N_11651);
xnor U12727 (N_12727,N_11955,N_10018);
nand U12728 (N_12728,N_11102,N_10615);
nand U12729 (N_12729,N_10629,N_11885);
or U12730 (N_12730,N_10785,N_11466);
nand U12731 (N_12731,N_11501,N_11282);
and U12732 (N_12732,N_10670,N_11183);
or U12733 (N_12733,N_10279,N_11698);
nor U12734 (N_12734,N_10091,N_11280);
nor U12735 (N_12735,N_10696,N_10531);
and U12736 (N_12736,N_11892,N_11400);
nand U12737 (N_12737,N_11783,N_10040);
and U12738 (N_12738,N_10946,N_10916);
or U12739 (N_12739,N_10405,N_11770);
and U12740 (N_12740,N_10776,N_11591);
nor U12741 (N_12741,N_10461,N_10280);
nand U12742 (N_12742,N_11278,N_11041);
nor U12743 (N_12743,N_10644,N_10254);
or U12744 (N_12744,N_11606,N_11101);
or U12745 (N_12745,N_11982,N_11742);
nand U12746 (N_12746,N_11734,N_10187);
nand U12747 (N_12747,N_10971,N_11374);
or U12748 (N_12748,N_11483,N_11887);
nor U12749 (N_12749,N_11140,N_11881);
nor U12750 (N_12750,N_11274,N_11862);
or U12751 (N_12751,N_11371,N_11136);
and U12752 (N_12752,N_10805,N_11656);
nor U12753 (N_12753,N_10845,N_10677);
nand U12754 (N_12754,N_11702,N_10014);
nand U12755 (N_12755,N_11882,N_10002);
or U12756 (N_12756,N_11825,N_11909);
nor U12757 (N_12757,N_11846,N_11893);
xnor U12758 (N_12758,N_10717,N_11161);
and U12759 (N_12759,N_11990,N_11861);
or U12760 (N_12760,N_11780,N_10010);
xor U12761 (N_12761,N_11951,N_10998);
nand U12762 (N_12762,N_11930,N_10628);
or U12763 (N_12763,N_10075,N_10033);
and U12764 (N_12764,N_11272,N_10550);
nor U12765 (N_12765,N_10559,N_11762);
nand U12766 (N_12766,N_10958,N_10616);
nor U12767 (N_12767,N_10483,N_11439);
or U12768 (N_12768,N_11485,N_10885);
nand U12769 (N_12769,N_11075,N_11986);
xor U12770 (N_12770,N_11262,N_10389);
or U12771 (N_12771,N_10447,N_10514);
and U12772 (N_12772,N_10530,N_11957);
and U12773 (N_12773,N_10496,N_10728);
and U12774 (N_12774,N_11302,N_10451);
and U12775 (N_12775,N_10223,N_10826);
nor U12776 (N_12776,N_11369,N_11984);
xor U12777 (N_12777,N_11284,N_11923);
nand U12778 (N_12778,N_10163,N_10561);
nand U12779 (N_12779,N_10505,N_10814);
xnor U12780 (N_12780,N_10070,N_11597);
nor U12781 (N_12781,N_10861,N_10994);
nand U12782 (N_12782,N_10475,N_11581);
or U12783 (N_12783,N_10470,N_11586);
and U12784 (N_12784,N_11561,N_10134);
or U12785 (N_12785,N_10842,N_10067);
nand U12786 (N_12786,N_10822,N_11813);
xnor U12787 (N_12787,N_10358,N_11260);
and U12788 (N_12788,N_11851,N_11499);
xnor U12789 (N_12789,N_11776,N_11576);
or U12790 (N_12790,N_10618,N_11367);
and U12791 (N_12791,N_11750,N_10181);
nand U12792 (N_12792,N_11692,N_11032);
or U12793 (N_12793,N_10325,N_10985);
xor U12794 (N_12794,N_11015,N_10562);
nand U12795 (N_12795,N_10116,N_10655);
nand U12796 (N_12796,N_11343,N_11566);
and U12797 (N_12797,N_11448,N_11596);
and U12798 (N_12798,N_10564,N_11879);
nand U12799 (N_12799,N_10338,N_11665);
and U12800 (N_12800,N_10640,N_11965);
nand U12801 (N_12801,N_10721,N_11949);
nand U12802 (N_12802,N_10450,N_10170);
or U12803 (N_12803,N_10211,N_11324);
or U12804 (N_12804,N_11509,N_11756);
xnor U12805 (N_12805,N_11511,N_10159);
nor U12806 (N_12806,N_10560,N_10766);
nor U12807 (N_12807,N_11067,N_10745);
or U12808 (N_12808,N_10939,N_11469);
xor U12809 (N_12809,N_11342,N_11636);
or U12810 (N_12810,N_10866,N_11868);
nand U12811 (N_12811,N_11878,N_11049);
xor U12812 (N_12812,N_11931,N_10954);
and U12813 (N_12813,N_11927,N_10078);
nand U12814 (N_12814,N_10345,N_10749);
and U12815 (N_12815,N_11496,N_10568);
and U12816 (N_12816,N_11333,N_10965);
nand U12817 (N_12817,N_10818,N_10704);
or U12818 (N_12818,N_10709,N_10606);
and U12819 (N_12819,N_10440,N_10678);
nor U12820 (N_12820,N_10297,N_11188);
nand U12821 (N_12821,N_11710,N_10723);
and U12822 (N_12822,N_11230,N_11475);
nand U12823 (N_12823,N_11697,N_11582);
nand U12824 (N_12824,N_10122,N_11211);
nor U12825 (N_12825,N_10702,N_11805);
or U12826 (N_12826,N_10474,N_11010);
or U12827 (N_12827,N_11772,N_10938);
nor U12828 (N_12828,N_10737,N_10526);
xor U12829 (N_12829,N_10088,N_10214);
and U12830 (N_12830,N_10284,N_11137);
nor U12831 (N_12831,N_10443,N_10322);
nand U12832 (N_12832,N_10652,N_10138);
or U12833 (N_12833,N_11245,N_11422);
nand U12834 (N_12834,N_11232,N_11040);
and U12835 (N_12835,N_11035,N_10178);
or U12836 (N_12836,N_11312,N_10620);
and U12837 (N_12837,N_10689,N_11503);
nand U12838 (N_12838,N_11821,N_10441);
or U12839 (N_12839,N_11294,N_10157);
nor U12840 (N_12840,N_10488,N_11973);
nand U12841 (N_12841,N_11635,N_11064);
or U12842 (N_12842,N_10295,N_11304);
or U12843 (N_12843,N_10011,N_11598);
or U12844 (N_12844,N_11701,N_11350);
or U12845 (N_12845,N_11385,N_11900);
or U12846 (N_12846,N_10056,N_10596);
nor U12847 (N_12847,N_11670,N_11658);
or U12848 (N_12848,N_11492,N_11127);
and U12849 (N_12849,N_10906,N_10680);
or U12850 (N_12850,N_11989,N_11054);
and U12851 (N_12851,N_10212,N_11932);
nand U12852 (N_12852,N_11011,N_10520);
and U12853 (N_12853,N_11195,N_11001);
nor U12854 (N_12854,N_11615,N_10293);
and U12855 (N_12855,N_11070,N_11768);
nand U12856 (N_12856,N_10726,N_10793);
nor U12857 (N_12857,N_11378,N_10921);
and U12858 (N_12858,N_10495,N_11833);
xor U12859 (N_12859,N_10697,N_10872);
or U12860 (N_12860,N_10262,N_11042);
or U12861 (N_12861,N_10438,N_11542);
or U12862 (N_12862,N_10819,N_11739);
and U12863 (N_12863,N_10605,N_10744);
or U12864 (N_12864,N_10182,N_11609);
nor U12865 (N_12865,N_11390,N_10107);
nand U12866 (N_12866,N_11379,N_10422);
xnor U12867 (N_12867,N_10490,N_10206);
or U12868 (N_12868,N_10732,N_11529);
nor U12869 (N_12869,N_11254,N_10752);
and U12870 (N_12870,N_10225,N_10761);
nand U12871 (N_12871,N_10320,N_11004);
or U12872 (N_12872,N_11249,N_10224);
nand U12873 (N_12873,N_10807,N_10714);
or U12874 (N_12874,N_11603,N_10883);
or U12875 (N_12875,N_11696,N_10833);
and U12876 (N_12876,N_11346,N_10660);
nand U12877 (N_12877,N_10119,N_11849);
nand U12878 (N_12878,N_10009,N_10216);
and U12879 (N_12879,N_11173,N_10287);
and U12880 (N_12880,N_11269,N_11926);
or U12881 (N_12881,N_11191,N_11264);
nor U12882 (N_12882,N_11831,N_10563);
or U12883 (N_12883,N_10593,N_11901);
or U12884 (N_12884,N_11854,N_10158);
and U12885 (N_12885,N_11641,N_11301);
nand U12886 (N_12886,N_10403,N_11800);
xnor U12887 (N_12887,N_11375,N_10783);
xnor U12888 (N_12888,N_11564,N_11488);
and U12889 (N_12889,N_11653,N_10314);
nand U12890 (N_12890,N_10069,N_10734);
nor U12891 (N_12891,N_10005,N_10880);
nand U12892 (N_12892,N_11954,N_10041);
or U12893 (N_12893,N_10466,N_10143);
nor U12894 (N_12894,N_11767,N_11026);
or U12895 (N_12895,N_10331,N_11281);
and U12896 (N_12896,N_10933,N_11690);
nand U12897 (N_12897,N_10111,N_11922);
xnor U12898 (N_12898,N_11120,N_10310);
nand U12899 (N_12899,N_10068,N_10686);
and U12900 (N_12900,N_10053,N_11587);
nor U12901 (N_12901,N_11495,N_10154);
nor U12902 (N_12902,N_10932,N_10850);
xor U12903 (N_12903,N_11666,N_11008);
nor U12904 (N_12904,N_11336,N_10460);
xor U12905 (N_12905,N_11470,N_11383);
nor U12906 (N_12906,N_10508,N_11403);
nor U12907 (N_12907,N_10489,N_10963);
or U12908 (N_12908,N_10132,N_10277);
nor U12909 (N_12909,N_10045,N_10546);
nand U12910 (N_12910,N_10851,N_11708);
nor U12911 (N_12911,N_11633,N_11981);
nor U12912 (N_12912,N_10638,N_11682);
and U12913 (N_12913,N_11593,N_10928);
or U12914 (N_12914,N_10066,N_11553);
or U12915 (N_12915,N_11125,N_10431);
nor U12916 (N_12916,N_10454,N_11867);
and U12917 (N_12917,N_11786,N_10235);
nand U12918 (N_12918,N_10553,N_11357);
or U12919 (N_12919,N_11021,N_11398);
or U12920 (N_12920,N_10218,N_11353);
nand U12921 (N_12921,N_11823,N_11836);
or U12922 (N_12922,N_11224,N_10177);
nor U12923 (N_12923,N_11972,N_11445);
or U12924 (N_12924,N_10176,N_10456);
nor U12925 (N_12925,N_11352,N_11668);
nor U12926 (N_12926,N_11730,N_11061);
or U12927 (N_12927,N_10767,N_10276);
nor U12928 (N_12928,N_11467,N_11286);
or U12929 (N_12929,N_11504,N_10199);
and U12930 (N_12930,N_11748,N_11009);
nand U12931 (N_12931,N_10899,N_10665);
and U12932 (N_12932,N_11792,N_11654);
nor U12933 (N_12933,N_11095,N_10666);
or U12934 (N_12934,N_11415,N_11618);
xor U12935 (N_12935,N_10368,N_10184);
or U12936 (N_12936,N_11546,N_11605);
or U12937 (N_12937,N_10565,N_11567);
nor U12938 (N_12938,N_10979,N_10305);
nand U12939 (N_12939,N_10500,N_10458);
nor U12940 (N_12940,N_10876,N_10952);
nor U12941 (N_12941,N_11680,N_11910);
or U12942 (N_12942,N_10251,N_11266);
nand U12943 (N_12943,N_10133,N_11438);
and U12944 (N_12944,N_11199,N_10781);
nand U12945 (N_12945,N_11903,N_10174);
or U12946 (N_12946,N_11465,N_11968);
nor U12947 (N_12947,N_10467,N_11486);
and U12948 (N_12948,N_10108,N_10525);
and U12949 (N_12949,N_10061,N_10942);
nor U12950 (N_12950,N_11917,N_11314);
or U12951 (N_12951,N_11500,N_11738);
and U12952 (N_12952,N_10278,N_10871);
xor U12953 (N_12953,N_10094,N_11458);
and U12954 (N_12954,N_11099,N_10126);
or U12955 (N_12955,N_10076,N_11198);
nor U12956 (N_12956,N_10636,N_11491);
and U12957 (N_12957,N_10329,N_10836);
xor U12958 (N_12958,N_10802,N_11457);
nand U12959 (N_12959,N_11997,N_11146);
nor U12960 (N_12960,N_11168,N_11446);
or U12961 (N_12961,N_11875,N_10664);
nor U12962 (N_12962,N_11589,N_11478);
nor U12963 (N_12963,N_11758,N_11200);
or U12964 (N_12964,N_10244,N_10455);
nand U12965 (N_12965,N_10828,N_11552);
nand U12966 (N_12966,N_10034,N_10213);
and U12967 (N_12967,N_10036,N_10272);
or U12968 (N_12968,N_11024,N_11729);
or U12969 (N_12969,N_10335,N_11693);
and U12970 (N_12970,N_11253,N_11335);
nand U12971 (N_12971,N_11045,N_10953);
and U12972 (N_12972,N_11840,N_10155);
or U12973 (N_12973,N_11594,N_10446);
nor U12974 (N_12974,N_10197,N_11983);
nand U12975 (N_12975,N_10228,N_11391);
nor U12976 (N_12976,N_10393,N_10622);
nand U12977 (N_12977,N_10252,N_11620);
nand U12978 (N_12978,N_10951,N_11871);
nand U12979 (N_12979,N_11645,N_11877);
xnor U12980 (N_12980,N_11914,N_11634);
or U12981 (N_12981,N_11778,N_11637);
and U12982 (N_12982,N_10909,N_10308);
or U12983 (N_12983,N_10291,N_11381);
xnor U12984 (N_12984,N_11135,N_10667);
xnor U12985 (N_12985,N_11699,N_11081);
nor U12986 (N_12986,N_10739,N_10463);
or U12987 (N_12987,N_11522,N_11947);
xor U12988 (N_12988,N_11124,N_11450);
or U12989 (N_12989,N_11416,N_11327);
nor U12990 (N_12990,N_10535,N_11331);
and U12991 (N_12991,N_11551,N_10104);
nand U12992 (N_12992,N_10417,N_11430);
or U12993 (N_12993,N_11480,N_11113);
or U12994 (N_12994,N_11745,N_11147);
or U12995 (N_12995,N_11642,N_10232);
nor U12996 (N_12996,N_10632,N_10863);
nor U12997 (N_12997,N_10092,N_11638);
xnor U12998 (N_12998,N_11960,N_10786);
nand U12999 (N_12999,N_10860,N_10398);
and U13000 (N_13000,N_11034,N_10792);
xor U13001 (N_13001,N_10687,N_10003);
and U13002 (N_13002,N_10064,N_11753);
nand U13003 (N_13003,N_10515,N_11874);
or U13004 (N_13004,N_11092,N_11452);
nor U13005 (N_13005,N_10507,N_10728);
nand U13006 (N_13006,N_11071,N_11133);
xor U13007 (N_13007,N_10223,N_11408);
or U13008 (N_13008,N_10013,N_11929);
or U13009 (N_13009,N_10977,N_11643);
nor U13010 (N_13010,N_10904,N_11659);
nor U13011 (N_13011,N_11645,N_11501);
nand U13012 (N_13012,N_11165,N_11725);
nand U13013 (N_13013,N_11864,N_10004);
or U13014 (N_13014,N_10102,N_10517);
and U13015 (N_13015,N_11674,N_11838);
or U13016 (N_13016,N_11567,N_11645);
nor U13017 (N_13017,N_11688,N_10634);
nand U13018 (N_13018,N_10192,N_10063);
xnor U13019 (N_13019,N_11465,N_10972);
and U13020 (N_13020,N_11328,N_10904);
or U13021 (N_13021,N_10562,N_10300);
or U13022 (N_13022,N_10570,N_11073);
and U13023 (N_13023,N_10050,N_10545);
nand U13024 (N_13024,N_10506,N_10501);
xor U13025 (N_13025,N_11385,N_10235);
nand U13026 (N_13026,N_10266,N_10872);
nand U13027 (N_13027,N_10730,N_11693);
or U13028 (N_13028,N_11734,N_11679);
xor U13029 (N_13029,N_10620,N_10000);
and U13030 (N_13030,N_11146,N_10370);
nand U13031 (N_13031,N_11820,N_10037);
nand U13032 (N_13032,N_10234,N_10625);
and U13033 (N_13033,N_10965,N_10612);
nor U13034 (N_13034,N_11885,N_11728);
or U13035 (N_13035,N_10978,N_11117);
or U13036 (N_13036,N_10260,N_10521);
nand U13037 (N_13037,N_11820,N_10380);
xor U13038 (N_13038,N_11029,N_11994);
nand U13039 (N_13039,N_11951,N_11266);
nand U13040 (N_13040,N_10759,N_11921);
xnor U13041 (N_13041,N_11675,N_10336);
and U13042 (N_13042,N_11498,N_10968);
and U13043 (N_13043,N_11558,N_10902);
nor U13044 (N_13044,N_11110,N_10260);
nand U13045 (N_13045,N_10071,N_10853);
and U13046 (N_13046,N_10338,N_11855);
and U13047 (N_13047,N_10923,N_11629);
nor U13048 (N_13048,N_11789,N_11285);
xnor U13049 (N_13049,N_11792,N_10175);
nor U13050 (N_13050,N_11061,N_11975);
nand U13051 (N_13051,N_10741,N_11112);
xnor U13052 (N_13052,N_10039,N_10727);
or U13053 (N_13053,N_11084,N_10185);
or U13054 (N_13054,N_11249,N_10624);
nor U13055 (N_13055,N_10940,N_11087);
nand U13056 (N_13056,N_10303,N_10191);
nor U13057 (N_13057,N_11574,N_11185);
or U13058 (N_13058,N_10362,N_10038);
nor U13059 (N_13059,N_11326,N_10807);
nand U13060 (N_13060,N_11978,N_10929);
or U13061 (N_13061,N_10048,N_11944);
nor U13062 (N_13062,N_10698,N_10988);
nor U13063 (N_13063,N_11109,N_10750);
nor U13064 (N_13064,N_11714,N_10925);
xor U13065 (N_13065,N_10625,N_11898);
xnor U13066 (N_13066,N_11492,N_11461);
nand U13067 (N_13067,N_10323,N_11292);
nand U13068 (N_13068,N_10156,N_11534);
or U13069 (N_13069,N_10393,N_10133);
nand U13070 (N_13070,N_11387,N_11207);
nor U13071 (N_13071,N_11222,N_10014);
and U13072 (N_13072,N_11514,N_11529);
or U13073 (N_13073,N_10677,N_10113);
and U13074 (N_13074,N_11479,N_11401);
and U13075 (N_13075,N_10513,N_10055);
and U13076 (N_13076,N_10422,N_11357);
and U13077 (N_13077,N_10385,N_10467);
nor U13078 (N_13078,N_11278,N_10388);
and U13079 (N_13079,N_10060,N_10714);
nor U13080 (N_13080,N_11794,N_11452);
nand U13081 (N_13081,N_10947,N_11912);
and U13082 (N_13082,N_11657,N_10421);
nand U13083 (N_13083,N_10543,N_10284);
and U13084 (N_13084,N_11036,N_11964);
nand U13085 (N_13085,N_10699,N_11454);
or U13086 (N_13086,N_10222,N_11704);
nor U13087 (N_13087,N_11204,N_10071);
nor U13088 (N_13088,N_11203,N_11004);
xor U13089 (N_13089,N_11806,N_10723);
and U13090 (N_13090,N_10290,N_10359);
and U13091 (N_13091,N_11327,N_10422);
and U13092 (N_13092,N_10371,N_11619);
nor U13093 (N_13093,N_11859,N_11268);
nor U13094 (N_13094,N_10031,N_10409);
nor U13095 (N_13095,N_11525,N_10058);
nand U13096 (N_13096,N_11737,N_11103);
or U13097 (N_13097,N_10309,N_11774);
nand U13098 (N_13098,N_10579,N_10919);
nand U13099 (N_13099,N_11730,N_10310);
or U13100 (N_13100,N_10259,N_11543);
xnor U13101 (N_13101,N_11857,N_11480);
or U13102 (N_13102,N_11608,N_11186);
and U13103 (N_13103,N_10640,N_10831);
and U13104 (N_13104,N_11824,N_11205);
or U13105 (N_13105,N_11826,N_10593);
xor U13106 (N_13106,N_10251,N_10756);
nor U13107 (N_13107,N_10032,N_11821);
and U13108 (N_13108,N_11949,N_10596);
nand U13109 (N_13109,N_10134,N_11890);
nand U13110 (N_13110,N_11502,N_10622);
nor U13111 (N_13111,N_10208,N_11663);
nand U13112 (N_13112,N_11375,N_10596);
nand U13113 (N_13113,N_10277,N_11567);
nand U13114 (N_13114,N_11326,N_10189);
nand U13115 (N_13115,N_11492,N_11459);
and U13116 (N_13116,N_11226,N_10427);
or U13117 (N_13117,N_10726,N_11929);
nor U13118 (N_13118,N_11280,N_11705);
nor U13119 (N_13119,N_10005,N_10571);
or U13120 (N_13120,N_11194,N_10369);
or U13121 (N_13121,N_11108,N_11444);
xor U13122 (N_13122,N_11801,N_11281);
and U13123 (N_13123,N_11987,N_11566);
and U13124 (N_13124,N_10770,N_11960);
nand U13125 (N_13125,N_10727,N_10005);
or U13126 (N_13126,N_11112,N_10108);
nor U13127 (N_13127,N_11445,N_10795);
nor U13128 (N_13128,N_10474,N_11277);
or U13129 (N_13129,N_11719,N_11279);
and U13130 (N_13130,N_10834,N_11013);
nor U13131 (N_13131,N_11175,N_10870);
xor U13132 (N_13132,N_10137,N_11142);
xnor U13133 (N_13133,N_11230,N_11633);
and U13134 (N_13134,N_11379,N_10993);
xor U13135 (N_13135,N_11322,N_10705);
nand U13136 (N_13136,N_11876,N_11597);
and U13137 (N_13137,N_10834,N_11736);
nor U13138 (N_13138,N_11219,N_11177);
and U13139 (N_13139,N_10058,N_10186);
nand U13140 (N_13140,N_11998,N_11589);
xor U13141 (N_13141,N_11174,N_11375);
nor U13142 (N_13142,N_11654,N_11738);
and U13143 (N_13143,N_11963,N_10606);
nand U13144 (N_13144,N_11117,N_10718);
or U13145 (N_13145,N_10792,N_11560);
and U13146 (N_13146,N_10236,N_10705);
nand U13147 (N_13147,N_11829,N_10754);
nor U13148 (N_13148,N_11917,N_11137);
and U13149 (N_13149,N_10238,N_10477);
xor U13150 (N_13150,N_11563,N_11587);
nor U13151 (N_13151,N_10905,N_10243);
or U13152 (N_13152,N_11557,N_10345);
nor U13153 (N_13153,N_10568,N_10997);
nand U13154 (N_13154,N_10178,N_11442);
xnor U13155 (N_13155,N_10339,N_11676);
nand U13156 (N_13156,N_11073,N_10222);
or U13157 (N_13157,N_11931,N_10499);
nand U13158 (N_13158,N_11885,N_10251);
nor U13159 (N_13159,N_10874,N_11405);
or U13160 (N_13160,N_11847,N_10879);
and U13161 (N_13161,N_11085,N_10027);
and U13162 (N_13162,N_10204,N_10239);
nor U13163 (N_13163,N_10473,N_11953);
and U13164 (N_13164,N_11297,N_11362);
or U13165 (N_13165,N_11089,N_11173);
and U13166 (N_13166,N_11476,N_10602);
nand U13167 (N_13167,N_11423,N_11211);
xnor U13168 (N_13168,N_11894,N_11029);
nand U13169 (N_13169,N_11055,N_11830);
and U13170 (N_13170,N_10676,N_10506);
and U13171 (N_13171,N_11842,N_10492);
nor U13172 (N_13172,N_10108,N_11354);
nand U13173 (N_13173,N_10505,N_10192);
or U13174 (N_13174,N_10570,N_10564);
nand U13175 (N_13175,N_10263,N_11271);
and U13176 (N_13176,N_10839,N_11860);
nor U13177 (N_13177,N_11543,N_10781);
nand U13178 (N_13178,N_11612,N_10836);
nand U13179 (N_13179,N_11691,N_11845);
xnor U13180 (N_13180,N_11354,N_11866);
and U13181 (N_13181,N_11518,N_10650);
nand U13182 (N_13182,N_10975,N_11186);
and U13183 (N_13183,N_11345,N_10757);
xor U13184 (N_13184,N_11984,N_10580);
and U13185 (N_13185,N_10031,N_11071);
or U13186 (N_13186,N_10242,N_10593);
or U13187 (N_13187,N_11048,N_10607);
and U13188 (N_13188,N_11588,N_10206);
nand U13189 (N_13189,N_11042,N_10367);
and U13190 (N_13190,N_11156,N_10310);
and U13191 (N_13191,N_10539,N_11443);
or U13192 (N_13192,N_11827,N_10577);
and U13193 (N_13193,N_11133,N_10529);
xnor U13194 (N_13194,N_10155,N_11962);
nand U13195 (N_13195,N_11587,N_11276);
nand U13196 (N_13196,N_11858,N_10812);
and U13197 (N_13197,N_10271,N_11984);
xnor U13198 (N_13198,N_11535,N_11911);
nand U13199 (N_13199,N_10828,N_11144);
or U13200 (N_13200,N_10858,N_10137);
xnor U13201 (N_13201,N_10273,N_10535);
xnor U13202 (N_13202,N_11242,N_11681);
nand U13203 (N_13203,N_10392,N_11768);
nor U13204 (N_13204,N_10782,N_10148);
nand U13205 (N_13205,N_10520,N_10450);
or U13206 (N_13206,N_11877,N_10571);
nor U13207 (N_13207,N_10045,N_11044);
or U13208 (N_13208,N_11085,N_11831);
xor U13209 (N_13209,N_10297,N_10074);
or U13210 (N_13210,N_10877,N_10809);
or U13211 (N_13211,N_11917,N_11203);
or U13212 (N_13212,N_11271,N_11630);
nand U13213 (N_13213,N_10464,N_11012);
nor U13214 (N_13214,N_10081,N_11032);
or U13215 (N_13215,N_11249,N_10232);
and U13216 (N_13216,N_10221,N_10864);
nand U13217 (N_13217,N_10049,N_11829);
nor U13218 (N_13218,N_11719,N_10636);
or U13219 (N_13219,N_10627,N_10089);
and U13220 (N_13220,N_10649,N_11408);
or U13221 (N_13221,N_11296,N_11513);
nor U13222 (N_13222,N_10950,N_11369);
and U13223 (N_13223,N_10464,N_11405);
or U13224 (N_13224,N_11459,N_10706);
nand U13225 (N_13225,N_11639,N_11174);
nand U13226 (N_13226,N_11503,N_10912);
or U13227 (N_13227,N_10094,N_10360);
xor U13228 (N_13228,N_11325,N_11023);
and U13229 (N_13229,N_11466,N_11242);
and U13230 (N_13230,N_10275,N_11679);
nand U13231 (N_13231,N_11808,N_10010);
xnor U13232 (N_13232,N_10135,N_10983);
nand U13233 (N_13233,N_10128,N_10193);
xor U13234 (N_13234,N_10578,N_11226);
nand U13235 (N_13235,N_11253,N_11787);
nand U13236 (N_13236,N_10646,N_10893);
or U13237 (N_13237,N_11886,N_10119);
and U13238 (N_13238,N_10939,N_10625);
nand U13239 (N_13239,N_10710,N_10409);
nor U13240 (N_13240,N_11520,N_10354);
nor U13241 (N_13241,N_10323,N_11077);
nand U13242 (N_13242,N_11228,N_11575);
nand U13243 (N_13243,N_11853,N_11889);
and U13244 (N_13244,N_10447,N_11093);
and U13245 (N_13245,N_11567,N_11506);
nor U13246 (N_13246,N_10208,N_10180);
nor U13247 (N_13247,N_10107,N_11839);
nand U13248 (N_13248,N_10700,N_10178);
nor U13249 (N_13249,N_10406,N_11368);
nor U13250 (N_13250,N_10915,N_11011);
nand U13251 (N_13251,N_11729,N_11509);
nand U13252 (N_13252,N_11602,N_11763);
nand U13253 (N_13253,N_11658,N_11493);
or U13254 (N_13254,N_10044,N_11202);
nor U13255 (N_13255,N_11293,N_11915);
and U13256 (N_13256,N_11405,N_10584);
xor U13257 (N_13257,N_10436,N_11794);
and U13258 (N_13258,N_10771,N_10792);
nand U13259 (N_13259,N_10365,N_11710);
and U13260 (N_13260,N_11773,N_11393);
nand U13261 (N_13261,N_11020,N_10857);
or U13262 (N_13262,N_11731,N_11852);
nor U13263 (N_13263,N_10414,N_11934);
nor U13264 (N_13264,N_10123,N_10952);
nor U13265 (N_13265,N_10088,N_11179);
nand U13266 (N_13266,N_10733,N_10503);
or U13267 (N_13267,N_11593,N_11052);
or U13268 (N_13268,N_10568,N_11738);
nor U13269 (N_13269,N_11094,N_11761);
and U13270 (N_13270,N_10707,N_11082);
nand U13271 (N_13271,N_10244,N_10190);
nor U13272 (N_13272,N_11391,N_11346);
nand U13273 (N_13273,N_11865,N_10249);
or U13274 (N_13274,N_11759,N_11968);
and U13275 (N_13275,N_11537,N_10979);
nor U13276 (N_13276,N_10539,N_11629);
and U13277 (N_13277,N_10141,N_11980);
nor U13278 (N_13278,N_11180,N_10271);
nand U13279 (N_13279,N_11219,N_10510);
or U13280 (N_13280,N_10346,N_10318);
and U13281 (N_13281,N_11984,N_11068);
nand U13282 (N_13282,N_10240,N_10648);
nand U13283 (N_13283,N_11499,N_11153);
nor U13284 (N_13284,N_10442,N_11045);
xnor U13285 (N_13285,N_10344,N_10109);
or U13286 (N_13286,N_11497,N_10809);
and U13287 (N_13287,N_10226,N_10990);
or U13288 (N_13288,N_10647,N_11296);
nand U13289 (N_13289,N_10616,N_10545);
or U13290 (N_13290,N_10896,N_10743);
nand U13291 (N_13291,N_11775,N_11781);
and U13292 (N_13292,N_11641,N_11122);
or U13293 (N_13293,N_11498,N_10289);
xor U13294 (N_13294,N_11561,N_10210);
or U13295 (N_13295,N_11269,N_11696);
and U13296 (N_13296,N_11368,N_11076);
nand U13297 (N_13297,N_10736,N_11561);
nor U13298 (N_13298,N_11122,N_10090);
xor U13299 (N_13299,N_11790,N_10204);
and U13300 (N_13300,N_11537,N_11457);
nor U13301 (N_13301,N_11830,N_10084);
nand U13302 (N_13302,N_10383,N_11211);
or U13303 (N_13303,N_11915,N_11901);
xor U13304 (N_13304,N_10342,N_11902);
or U13305 (N_13305,N_11794,N_11222);
and U13306 (N_13306,N_10011,N_11087);
and U13307 (N_13307,N_10986,N_11541);
or U13308 (N_13308,N_11282,N_11067);
or U13309 (N_13309,N_11289,N_11024);
and U13310 (N_13310,N_10747,N_10372);
xnor U13311 (N_13311,N_11282,N_11735);
nand U13312 (N_13312,N_11775,N_10090);
nand U13313 (N_13313,N_11043,N_11315);
nor U13314 (N_13314,N_10460,N_11550);
or U13315 (N_13315,N_10416,N_11291);
and U13316 (N_13316,N_10577,N_11921);
xnor U13317 (N_13317,N_11177,N_10524);
or U13318 (N_13318,N_10475,N_10721);
or U13319 (N_13319,N_11479,N_11325);
nand U13320 (N_13320,N_10639,N_10629);
nand U13321 (N_13321,N_10312,N_11814);
nor U13322 (N_13322,N_11894,N_10697);
and U13323 (N_13323,N_10988,N_10442);
nor U13324 (N_13324,N_10983,N_10737);
nor U13325 (N_13325,N_11432,N_10609);
and U13326 (N_13326,N_11074,N_11566);
xor U13327 (N_13327,N_11140,N_11742);
xnor U13328 (N_13328,N_10356,N_11523);
nand U13329 (N_13329,N_11574,N_11781);
or U13330 (N_13330,N_10116,N_11823);
nor U13331 (N_13331,N_10320,N_11915);
or U13332 (N_13332,N_10660,N_11072);
nand U13333 (N_13333,N_11354,N_11231);
xor U13334 (N_13334,N_10558,N_11817);
nand U13335 (N_13335,N_11862,N_10745);
or U13336 (N_13336,N_11578,N_11870);
or U13337 (N_13337,N_11854,N_10757);
or U13338 (N_13338,N_10396,N_11419);
and U13339 (N_13339,N_11980,N_10788);
nand U13340 (N_13340,N_11403,N_10155);
xnor U13341 (N_13341,N_10405,N_10478);
and U13342 (N_13342,N_10391,N_11211);
nor U13343 (N_13343,N_10763,N_11157);
or U13344 (N_13344,N_11311,N_10564);
nor U13345 (N_13345,N_11759,N_11379);
nor U13346 (N_13346,N_11900,N_11949);
xor U13347 (N_13347,N_10413,N_11764);
xnor U13348 (N_13348,N_11770,N_11136);
nand U13349 (N_13349,N_11313,N_11624);
or U13350 (N_13350,N_11513,N_10475);
nor U13351 (N_13351,N_11606,N_11966);
or U13352 (N_13352,N_11068,N_10451);
and U13353 (N_13353,N_10193,N_10787);
and U13354 (N_13354,N_10872,N_10573);
nor U13355 (N_13355,N_11901,N_10735);
or U13356 (N_13356,N_10505,N_11764);
or U13357 (N_13357,N_10777,N_10062);
xnor U13358 (N_13358,N_11622,N_11976);
and U13359 (N_13359,N_11326,N_10407);
and U13360 (N_13360,N_11523,N_10910);
nor U13361 (N_13361,N_11168,N_11583);
nor U13362 (N_13362,N_10701,N_11482);
xor U13363 (N_13363,N_11698,N_10715);
nor U13364 (N_13364,N_11691,N_10684);
or U13365 (N_13365,N_11191,N_10961);
or U13366 (N_13366,N_11752,N_10169);
or U13367 (N_13367,N_10642,N_10932);
nand U13368 (N_13368,N_10057,N_10816);
nor U13369 (N_13369,N_10469,N_10271);
and U13370 (N_13370,N_10866,N_10729);
nand U13371 (N_13371,N_11294,N_11025);
nand U13372 (N_13372,N_10523,N_10583);
or U13373 (N_13373,N_10610,N_10433);
and U13374 (N_13374,N_10393,N_11795);
and U13375 (N_13375,N_10811,N_10101);
and U13376 (N_13376,N_10090,N_10303);
or U13377 (N_13377,N_10723,N_10045);
xor U13378 (N_13378,N_10870,N_11248);
nand U13379 (N_13379,N_10795,N_10738);
nand U13380 (N_13380,N_11851,N_11234);
nand U13381 (N_13381,N_10460,N_10161);
nand U13382 (N_13382,N_11937,N_10600);
nor U13383 (N_13383,N_10626,N_11959);
nor U13384 (N_13384,N_10099,N_11255);
nor U13385 (N_13385,N_11988,N_10529);
or U13386 (N_13386,N_11601,N_10552);
or U13387 (N_13387,N_10632,N_11171);
or U13388 (N_13388,N_11823,N_11367);
nor U13389 (N_13389,N_11335,N_10312);
nand U13390 (N_13390,N_10425,N_10982);
nor U13391 (N_13391,N_11399,N_11129);
nor U13392 (N_13392,N_11095,N_11751);
or U13393 (N_13393,N_10722,N_10859);
xnor U13394 (N_13394,N_11506,N_11544);
and U13395 (N_13395,N_10256,N_10815);
and U13396 (N_13396,N_11880,N_11978);
nand U13397 (N_13397,N_10281,N_10188);
nor U13398 (N_13398,N_11020,N_10472);
and U13399 (N_13399,N_11565,N_11197);
or U13400 (N_13400,N_11260,N_10304);
or U13401 (N_13401,N_10259,N_11213);
nor U13402 (N_13402,N_10663,N_10389);
and U13403 (N_13403,N_11690,N_11320);
or U13404 (N_13404,N_11317,N_11237);
nor U13405 (N_13405,N_11028,N_11884);
nor U13406 (N_13406,N_10872,N_11744);
nor U13407 (N_13407,N_11598,N_10121);
or U13408 (N_13408,N_10715,N_11727);
or U13409 (N_13409,N_10011,N_11138);
xnor U13410 (N_13410,N_11247,N_11836);
or U13411 (N_13411,N_11375,N_11571);
xor U13412 (N_13412,N_10052,N_11260);
nor U13413 (N_13413,N_11074,N_10635);
xnor U13414 (N_13414,N_10492,N_11526);
xor U13415 (N_13415,N_11932,N_10485);
nor U13416 (N_13416,N_11336,N_10479);
nor U13417 (N_13417,N_11779,N_11216);
nor U13418 (N_13418,N_10353,N_10254);
nor U13419 (N_13419,N_10076,N_11184);
and U13420 (N_13420,N_10785,N_10955);
and U13421 (N_13421,N_11513,N_11935);
nand U13422 (N_13422,N_10657,N_11540);
nand U13423 (N_13423,N_11166,N_11473);
or U13424 (N_13424,N_10168,N_10541);
and U13425 (N_13425,N_10989,N_10721);
nand U13426 (N_13426,N_10516,N_11066);
nor U13427 (N_13427,N_10349,N_10433);
nand U13428 (N_13428,N_10933,N_10021);
nand U13429 (N_13429,N_10588,N_10599);
nor U13430 (N_13430,N_11516,N_10910);
nor U13431 (N_13431,N_10309,N_11015);
xnor U13432 (N_13432,N_10630,N_11856);
nor U13433 (N_13433,N_10298,N_11678);
or U13434 (N_13434,N_10023,N_10738);
nand U13435 (N_13435,N_10309,N_10494);
nand U13436 (N_13436,N_11085,N_10615);
or U13437 (N_13437,N_11725,N_10821);
and U13438 (N_13438,N_11819,N_11162);
nor U13439 (N_13439,N_10307,N_10558);
nand U13440 (N_13440,N_11700,N_11542);
nand U13441 (N_13441,N_11847,N_11472);
or U13442 (N_13442,N_11110,N_10388);
or U13443 (N_13443,N_11947,N_10124);
nand U13444 (N_13444,N_10449,N_11640);
or U13445 (N_13445,N_10106,N_10924);
or U13446 (N_13446,N_11410,N_10543);
nand U13447 (N_13447,N_11012,N_10043);
and U13448 (N_13448,N_11220,N_10440);
and U13449 (N_13449,N_10591,N_11283);
or U13450 (N_13450,N_11750,N_11485);
or U13451 (N_13451,N_11515,N_11576);
or U13452 (N_13452,N_11531,N_11845);
or U13453 (N_13453,N_11838,N_11675);
nor U13454 (N_13454,N_11805,N_10190);
nor U13455 (N_13455,N_11090,N_10262);
and U13456 (N_13456,N_10779,N_11505);
nor U13457 (N_13457,N_11018,N_10697);
or U13458 (N_13458,N_11534,N_10477);
or U13459 (N_13459,N_10039,N_11848);
nand U13460 (N_13460,N_10027,N_10844);
nand U13461 (N_13461,N_11867,N_10495);
and U13462 (N_13462,N_10318,N_11539);
and U13463 (N_13463,N_11690,N_11675);
nor U13464 (N_13464,N_10473,N_11191);
and U13465 (N_13465,N_11392,N_11152);
nand U13466 (N_13466,N_11630,N_11358);
or U13467 (N_13467,N_10943,N_10864);
and U13468 (N_13468,N_10703,N_11357);
nand U13469 (N_13469,N_10157,N_11923);
and U13470 (N_13470,N_10240,N_11167);
nand U13471 (N_13471,N_11625,N_11495);
or U13472 (N_13472,N_11051,N_11557);
and U13473 (N_13473,N_11579,N_11059);
or U13474 (N_13474,N_11477,N_10215);
nand U13475 (N_13475,N_11061,N_11494);
nand U13476 (N_13476,N_10725,N_11435);
xor U13477 (N_13477,N_11207,N_10498);
nor U13478 (N_13478,N_11384,N_10321);
nand U13479 (N_13479,N_11084,N_10324);
nor U13480 (N_13480,N_11805,N_10117);
or U13481 (N_13481,N_11742,N_10715);
and U13482 (N_13482,N_11222,N_11750);
nor U13483 (N_13483,N_10452,N_10500);
nor U13484 (N_13484,N_10823,N_11331);
and U13485 (N_13485,N_10194,N_10338);
and U13486 (N_13486,N_11769,N_10355);
xor U13487 (N_13487,N_10154,N_10037);
and U13488 (N_13488,N_11772,N_11953);
nor U13489 (N_13489,N_11609,N_11086);
xnor U13490 (N_13490,N_11669,N_10477);
nand U13491 (N_13491,N_11670,N_10812);
nor U13492 (N_13492,N_10560,N_11446);
xor U13493 (N_13493,N_10039,N_10390);
nor U13494 (N_13494,N_11556,N_10576);
and U13495 (N_13495,N_11939,N_10121);
nor U13496 (N_13496,N_10803,N_11692);
or U13497 (N_13497,N_10548,N_10217);
xor U13498 (N_13498,N_11339,N_11512);
nand U13499 (N_13499,N_11697,N_10863);
nor U13500 (N_13500,N_11730,N_10242);
nand U13501 (N_13501,N_10839,N_10332);
and U13502 (N_13502,N_11815,N_11242);
nand U13503 (N_13503,N_10467,N_11459);
nand U13504 (N_13504,N_11074,N_11540);
nor U13505 (N_13505,N_10201,N_10689);
or U13506 (N_13506,N_11972,N_11584);
nand U13507 (N_13507,N_11573,N_11452);
and U13508 (N_13508,N_10672,N_11974);
and U13509 (N_13509,N_11763,N_10820);
nor U13510 (N_13510,N_10804,N_11935);
xnor U13511 (N_13511,N_11327,N_10668);
nor U13512 (N_13512,N_11197,N_10168);
and U13513 (N_13513,N_11684,N_10240);
nor U13514 (N_13514,N_10287,N_11416);
or U13515 (N_13515,N_10075,N_11619);
or U13516 (N_13516,N_11656,N_10283);
xor U13517 (N_13517,N_10547,N_10288);
or U13518 (N_13518,N_11682,N_11943);
nor U13519 (N_13519,N_11927,N_10694);
or U13520 (N_13520,N_11697,N_11021);
nor U13521 (N_13521,N_10655,N_10001);
nand U13522 (N_13522,N_10771,N_10742);
or U13523 (N_13523,N_10103,N_11244);
or U13524 (N_13524,N_11596,N_10245);
nor U13525 (N_13525,N_10278,N_10189);
nand U13526 (N_13526,N_11258,N_10978);
nand U13527 (N_13527,N_11716,N_11819);
and U13528 (N_13528,N_11973,N_11560);
nor U13529 (N_13529,N_11029,N_11690);
xnor U13530 (N_13530,N_10984,N_11094);
xor U13531 (N_13531,N_11569,N_11458);
and U13532 (N_13532,N_10798,N_10551);
or U13533 (N_13533,N_11987,N_11952);
nand U13534 (N_13534,N_10719,N_10958);
xnor U13535 (N_13535,N_11244,N_10030);
nand U13536 (N_13536,N_11339,N_11605);
and U13537 (N_13537,N_11589,N_11845);
nor U13538 (N_13538,N_10992,N_11812);
nor U13539 (N_13539,N_11269,N_10963);
nor U13540 (N_13540,N_11170,N_11883);
and U13541 (N_13541,N_10815,N_10325);
nor U13542 (N_13542,N_11892,N_11790);
nand U13543 (N_13543,N_10429,N_11392);
nor U13544 (N_13544,N_10800,N_10534);
and U13545 (N_13545,N_10736,N_11384);
or U13546 (N_13546,N_11135,N_11655);
xor U13547 (N_13547,N_11932,N_10822);
nor U13548 (N_13548,N_10538,N_10951);
and U13549 (N_13549,N_10441,N_10628);
and U13550 (N_13550,N_11831,N_10583);
or U13551 (N_13551,N_10651,N_10257);
and U13552 (N_13552,N_11326,N_10757);
and U13553 (N_13553,N_11608,N_10755);
xor U13554 (N_13554,N_11319,N_10970);
nor U13555 (N_13555,N_10427,N_11537);
nor U13556 (N_13556,N_10861,N_11349);
xor U13557 (N_13557,N_10358,N_10798);
nand U13558 (N_13558,N_10052,N_10868);
nand U13559 (N_13559,N_10737,N_10265);
and U13560 (N_13560,N_11555,N_11738);
or U13561 (N_13561,N_11052,N_10182);
or U13562 (N_13562,N_10265,N_11817);
and U13563 (N_13563,N_10561,N_11260);
nand U13564 (N_13564,N_10308,N_11910);
or U13565 (N_13565,N_10520,N_10801);
or U13566 (N_13566,N_11518,N_11988);
nand U13567 (N_13567,N_11273,N_10535);
nor U13568 (N_13568,N_10940,N_10011);
or U13569 (N_13569,N_11865,N_11164);
and U13570 (N_13570,N_11440,N_11141);
or U13571 (N_13571,N_11071,N_10986);
or U13572 (N_13572,N_10964,N_11864);
and U13573 (N_13573,N_10443,N_10841);
nor U13574 (N_13574,N_10452,N_11915);
and U13575 (N_13575,N_10689,N_11719);
and U13576 (N_13576,N_10479,N_11305);
and U13577 (N_13577,N_10284,N_11469);
xnor U13578 (N_13578,N_10855,N_10511);
and U13579 (N_13579,N_10519,N_10051);
or U13580 (N_13580,N_10049,N_10018);
xnor U13581 (N_13581,N_11073,N_11674);
xnor U13582 (N_13582,N_10296,N_10218);
or U13583 (N_13583,N_11235,N_10286);
nand U13584 (N_13584,N_11080,N_10082);
or U13585 (N_13585,N_10361,N_11971);
or U13586 (N_13586,N_11756,N_11444);
nand U13587 (N_13587,N_10183,N_11823);
nand U13588 (N_13588,N_11209,N_10645);
nand U13589 (N_13589,N_10321,N_10366);
or U13590 (N_13590,N_10937,N_10923);
nand U13591 (N_13591,N_10705,N_10615);
xor U13592 (N_13592,N_10804,N_10945);
nor U13593 (N_13593,N_11248,N_10878);
and U13594 (N_13594,N_11929,N_10411);
or U13595 (N_13595,N_11774,N_10655);
and U13596 (N_13596,N_11727,N_10052);
or U13597 (N_13597,N_10711,N_10695);
or U13598 (N_13598,N_11818,N_11062);
and U13599 (N_13599,N_11492,N_10299);
or U13600 (N_13600,N_11984,N_11741);
and U13601 (N_13601,N_11066,N_11466);
or U13602 (N_13602,N_11884,N_11036);
nor U13603 (N_13603,N_11071,N_10000);
nor U13604 (N_13604,N_11296,N_10957);
or U13605 (N_13605,N_10030,N_10343);
and U13606 (N_13606,N_11230,N_11046);
or U13607 (N_13607,N_10246,N_10055);
nand U13608 (N_13608,N_11012,N_10681);
nand U13609 (N_13609,N_11775,N_11736);
or U13610 (N_13610,N_11115,N_11781);
and U13611 (N_13611,N_11885,N_10199);
and U13612 (N_13612,N_11466,N_10985);
nor U13613 (N_13613,N_10278,N_10711);
nor U13614 (N_13614,N_10879,N_10806);
nor U13615 (N_13615,N_10967,N_11312);
or U13616 (N_13616,N_10343,N_10785);
or U13617 (N_13617,N_10182,N_10473);
xnor U13618 (N_13618,N_10640,N_11710);
nand U13619 (N_13619,N_11734,N_11005);
and U13620 (N_13620,N_10796,N_11418);
or U13621 (N_13621,N_10460,N_10072);
and U13622 (N_13622,N_10961,N_10334);
xor U13623 (N_13623,N_10164,N_10662);
nand U13624 (N_13624,N_11594,N_10059);
nand U13625 (N_13625,N_10335,N_10923);
nor U13626 (N_13626,N_10078,N_11018);
or U13627 (N_13627,N_10927,N_10969);
or U13628 (N_13628,N_11970,N_10396);
and U13629 (N_13629,N_11154,N_10690);
nand U13630 (N_13630,N_10783,N_11536);
and U13631 (N_13631,N_10471,N_10848);
nand U13632 (N_13632,N_11607,N_11179);
nor U13633 (N_13633,N_11565,N_10528);
xnor U13634 (N_13634,N_10635,N_10873);
or U13635 (N_13635,N_11592,N_11514);
or U13636 (N_13636,N_11973,N_11020);
nor U13637 (N_13637,N_11629,N_11512);
or U13638 (N_13638,N_11332,N_11614);
xor U13639 (N_13639,N_10582,N_10890);
and U13640 (N_13640,N_10584,N_11967);
nor U13641 (N_13641,N_11090,N_11383);
or U13642 (N_13642,N_10826,N_10396);
nand U13643 (N_13643,N_11885,N_11800);
xnor U13644 (N_13644,N_11728,N_10122);
and U13645 (N_13645,N_10394,N_11461);
nor U13646 (N_13646,N_10398,N_11324);
and U13647 (N_13647,N_11126,N_10079);
nand U13648 (N_13648,N_11779,N_10068);
or U13649 (N_13649,N_11427,N_10976);
nor U13650 (N_13650,N_11683,N_10836);
nand U13651 (N_13651,N_10073,N_11486);
or U13652 (N_13652,N_11381,N_11792);
and U13653 (N_13653,N_10337,N_11546);
and U13654 (N_13654,N_11735,N_10772);
and U13655 (N_13655,N_10732,N_10878);
and U13656 (N_13656,N_11933,N_10518);
nand U13657 (N_13657,N_10877,N_11607);
nand U13658 (N_13658,N_11746,N_10576);
nor U13659 (N_13659,N_10971,N_11148);
nor U13660 (N_13660,N_11807,N_10478);
xnor U13661 (N_13661,N_10288,N_11053);
nand U13662 (N_13662,N_10299,N_10822);
nor U13663 (N_13663,N_10469,N_11527);
xnor U13664 (N_13664,N_10350,N_11359);
and U13665 (N_13665,N_10163,N_10590);
or U13666 (N_13666,N_10679,N_10165);
and U13667 (N_13667,N_10711,N_11039);
and U13668 (N_13668,N_11816,N_11336);
nand U13669 (N_13669,N_11486,N_11248);
nand U13670 (N_13670,N_11097,N_10748);
nand U13671 (N_13671,N_11841,N_10619);
and U13672 (N_13672,N_10942,N_10703);
and U13673 (N_13673,N_10650,N_10049);
or U13674 (N_13674,N_10373,N_10589);
nand U13675 (N_13675,N_10931,N_11597);
and U13676 (N_13676,N_10768,N_10276);
nand U13677 (N_13677,N_10079,N_11831);
or U13678 (N_13678,N_11989,N_10848);
and U13679 (N_13679,N_10336,N_11628);
and U13680 (N_13680,N_10050,N_11603);
nand U13681 (N_13681,N_10430,N_10589);
or U13682 (N_13682,N_11359,N_10402);
xnor U13683 (N_13683,N_11528,N_11113);
or U13684 (N_13684,N_11072,N_10948);
nor U13685 (N_13685,N_11305,N_11516);
nor U13686 (N_13686,N_10708,N_10078);
nor U13687 (N_13687,N_10726,N_10626);
nor U13688 (N_13688,N_11384,N_11822);
or U13689 (N_13689,N_11370,N_11358);
and U13690 (N_13690,N_10278,N_11535);
nand U13691 (N_13691,N_11966,N_10851);
nor U13692 (N_13692,N_10621,N_10513);
or U13693 (N_13693,N_10101,N_11548);
and U13694 (N_13694,N_10652,N_11936);
nor U13695 (N_13695,N_11186,N_10102);
nand U13696 (N_13696,N_11748,N_11257);
and U13697 (N_13697,N_10954,N_10347);
nor U13698 (N_13698,N_11215,N_10347);
nand U13699 (N_13699,N_10266,N_11679);
and U13700 (N_13700,N_11031,N_10884);
xnor U13701 (N_13701,N_11121,N_10579);
nand U13702 (N_13702,N_11910,N_11110);
and U13703 (N_13703,N_11678,N_10649);
nor U13704 (N_13704,N_10037,N_11706);
or U13705 (N_13705,N_10970,N_10060);
nor U13706 (N_13706,N_10766,N_10657);
or U13707 (N_13707,N_11649,N_10751);
and U13708 (N_13708,N_10116,N_11231);
nor U13709 (N_13709,N_11206,N_10191);
and U13710 (N_13710,N_11618,N_11127);
nand U13711 (N_13711,N_11625,N_11626);
and U13712 (N_13712,N_11040,N_10979);
and U13713 (N_13713,N_10228,N_10300);
or U13714 (N_13714,N_10168,N_10114);
nand U13715 (N_13715,N_11797,N_11543);
nor U13716 (N_13716,N_11160,N_10884);
nand U13717 (N_13717,N_10369,N_10860);
xnor U13718 (N_13718,N_11388,N_10533);
and U13719 (N_13719,N_10593,N_11339);
and U13720 (N_13720,N_10235,N_10730);
xnor U13721 (N_13721,N_11391,N_11718);
or U13722 (N_13722,N_11695,N_11763);
nor U13723 (N_13723,N_11941,N_10852);
and U13724 (N_13724,N_11610,N_10393);
and U13725 (N_13725,N_10171,N_11078);
nor U13726 (N_13726,N_11986,N_11987);
and U13727 (N_13727,N_11905,N_10704);
and U13728 (N_13728,N_10342,N_11191);
nor U13729 (N_13729,N_10263,N_11186);
or U13730 (N_13730,N_11482,N_10554);
nand U13731 (N_13731,N_10820,N_11357);
or U13732 (N_13732,N_10140,N_11939);
and U13733 (N_13733,N_10250,N_10002);
nor U13734 (N_13734,N_11672,N_11254);
nor U13735 (N_13735,N_10351,N_11356);
xor U13736 (N_13736,N_11111,N_11752);
and U13737 (N_13737,N_11167,N_11135);
xor U13738 (N_13738,N_10006,N_10936);
nand U13739 (N_13739,N_10742,N_11371);
nor U13740 (N_13740,N_11021,N_10677);
xor U13741 (N_13741,N_10859,N_11390);
xor U13742 (N_13742,N_10068,N_10878);
or U13743 (N_13743,N_11089,N_11687);
and U13744 (N_13744,N_10200,N_11788);
nand U13745 (N_13745,N_10858,N_10982);
or U13746 (N_13746,N_11490,N_11596);
nor U13747 (N_13747,N_10677,N_11381);
nand U13748 (N_13748,N_10150,N_10792);
nand U13749 (N_13749,N_11034,N_10031);
nor U13750 (N_13750,N_10435,N_11608);
or U13751 (N_13751,N_10160,N_11845);
nand U13752 (N_13752,N_11370,N_11606);
nor U13753 (N_13753,N_11982,N_10118);
and U13754 (N_13754,N_11628,N_11366);
or U13755 (N_13755,N_11817,N_11217);
or U13756 (N_13756,N_10786,N_10248);
nor U13757 (N_13757,N_11814,N_10884);
nand U13758 (N_13758,N_10487,N_10082);
nor U13759 (N_13759,N_10392,N_10311);
nand U13760 (N_13760,N_11622,N_10097);
or U13761 (N_13761,N_11404,N_11074);
and U13762 (N_13762,N_11393,N_10546);
and U13763 (N_13763,N_11259,N_10390);
nor U13764 (N_13764,N_11729,N_11395);
and U13765 (N_13765,N_11509,N_10134);
and U13766 (N_13766,N_10426,N_11461);
or U13767 (N_13767,N_11466,N_11679);
nor U13768 (N_13768,N_11573,N_11748);
or U13769 (N_13769,N_10909,N_11377);
and U13770 (N_13770,N_11951,N_11601);
or U13771 (N_13771,N_11959,N_11098);
or U13772 (N_13772,N_10993,N_11611);
nand U13773 (N_13773,N_11884,N_10198);
nand U13774 (N_13774,N_10214,N_11413);
and U13775 (N_13775,N_10797,N_10725);
nor U13776 (N_13776,N_11531,N_10228);
nand U13777 (N_13777,N_11868,N_11068);
nand U13778 (N_13778,N_11866,N_11599);
nand U13779 (N_13779,N_11820,N_10309);
nand U13780 (N_13780,N_11963,N_10249);
or U13781 (N_13781,N_11233,N_11847);
nand U13782 (N_13782,N_10479,N_11570);
nor U13783 (N_13783,N_10846,N_11512);
xor U13784 (N_13784,N_10160,N_11879);
and U13785 (N_13785,N_10377,N_10184);
nor U13786 (N_13786,N_11365,N_11712);
nand U13787 (N_13787,N_11636,N_11977);
nor U13788 (N_13788,N_10346,N_11651);
nand U13789 (N_13789,N_11693,N_11089);
or U13790 (N_13790,N_10274,N_11042);
and U13791 (N_13791,N_10349,N_11233);
and U13792 (N_13792,N_10763,N_11437);
nand U13793 (N_13793,N_11320,N_10376);
or U13794 (N_13794,N_10174,N_10140);
and U13795 (N_13795,N_10506,N_10192);
nand U13796 (N_13796,N_11066,N_11072);
nor U13797 (N_13797,N_11227,N_10919);
or U13798 (N_13798,N_11836,N_11118);
and U13799 (N_13799,N_10906,N_11959);
and U13800 (N_13800,N_11951,N_11588);
nand U13801 (N_13801,N_10238,N_11246);
nand U13802 (N_13802,N_11340,N_10888);
nor U13803 (N_13803,N_11483,N_11093);
and U13804 (N_13804,N_10444,N_11579);
nor U13805 (N_13805,N_11198,N_10523);
xor U13806 (N_13806,N_10769,N_10072);
and U13807 (N_13807,N_11044,N_11621);
and U13808 (N_13808,N_11256,N_11045);
nor U13809 (N_13809,N_10015,N_10329);
xor U13810 (N_13810,N_10489,N_11643);
xnor U13811 (N_13811,N_10672,N_11884);
nand U13812 (N_13812,N_10018,N_10576);
or U13813 (N_13813,N_11250,N_11064);
or U13814 (N_13814,N_10416,N_11974);
and U13815 (N_13815,N_11918,N_11501);
nand U13816 (N_13816,N_10137,N_11744);
nand U13817 (N_13817,N_11367,N_10935);
xnor U13818 (N_13818,N_10500,N_10814);
nor U13819 (N_13819,N_11173,N_11464);
and U13820 (N_13820,N_10761,N_10686);
or U13821 (N_13821,N_11862,N_11646);
xor U13822 (N_13822,N_11732,N_10423);
xnor U13823 (N_13823,N_10364,N_10358);
nor U13824 (N_13824,N_10159,N_10748);
and U13825 (N_13825,N_10376,N_11929);
nor U13826 (N_13826,N_11541,N_10884);
nor U13827 (N_13827,N_11844,N_11474);
and U13828 (N_13828,N_11004,N_10999);
and U13829 (N_13829,N_10656,N_11194);
nor U13830 (N_13830,N_11853,N_11425);
or U13831 (N_13831,N_11948,N_11890);
nor U13832 (N_13832,N_10311,N_10565);
nand U13833 (N_13833,N_11285,N_10145);
or U13834 (N_13834,N_11111,N_10662);
xnor U13835 (N_13835,N_11523,N_11024);
and U13836 (N_13836,N_11626,N_11016);
nand U13837 (N_13837,N_10225,N_10940);
nor U13838 (N_13838,N_10989,N_10260);
xor U13839 (N_13839,N_10138,N_11765);
or U13840 (N_13840,N_11747,N_10120);
and U13841 (N_13841,N_10204,N_10882);
and U13842 (N_13842,N_10239,N_11247);
nor U13843 (N_13843,N_10698,N_11983);
and U13844 (N_13844,N_11335,N_10721);
nand U13845 (N_13845,N_10914,N_11695);
nor U13846 (N_13846,N_10386,N_10647);
or U13847 (N_13847,N_11440,N_11955);
or U13848 (N_13848,N_10465,N_10726);
and U13849 (N_13849,N_11902,N_10705);
xnor U13850 (N_13850,N_10460,N_10748);
nor U13851 (N_13851,N_11347,N_10846);
nor U13852 (N_13852,N_11514,N_10414);
or U13853 (N_13853,N_11615,N_10010);
or U13854 (N_13854,N_11561,N_11439);
nor U13855 (N_13855,N_11381,N_10388);
nand U13856 (N_13856,N_11764,N_11946);
xnor U13857 (N_13857,N_11362,N_10980);
xor U13858 (N_13858,N_10296,N_11535);
or U13859 (N_13859,N_10830,N_10956);
nor U13860 (N_13860,N_10683,N_11567);
xor U13861 (N_13861,N_11995,N_10549);
nor U13862 (N_13862,N_11508,N_10189);
nand U13863 (N_13863,N_11908,N_11030);
nand U13864 (N_13864,N_11275,N_11103);
nor U13865 (N_13865,N_10950,N_10398);
nor U13866 (N_13866,N_11111,N_10793);
nand U13867 (N_13867,N_11040,N_11732);
xnor U13868 (N_13868,N_11073,N_11247);
and U13869 (N_13869,N_11319,N_11712);
nor U13870 (N_13870,N_10085,N_10962);
or U13871 (N_13871,N_10869,N_10791);
and U13872 (N_13872,N_10940,N_10013);
and U13873 (N_13873,N_11662,N_11434);
nand U13874 (N_13874,N_11900,N_11383);
and U13875 (N_13875,N_10466,N_10287);
or U13876 (N_13876,N_10500,N_10373);
nor U13877 (N_13877,N_11909,N_11196);
nand U13878 (N_13878,N_11987,N_11270);
nand U13879 (N_13879,N_10825,N_10381);
or U13880 (N_13880,N_10929,N_11674);
nor U13881 (N_13881,N_11617,N_10272);
or U13882 (N_13882,N_10942,N_11301);
and U13883 (N_13883,N_11568,N_10806);
nand U13884 (N_13884,N_11540,N_10218);
and U13885 (N_13885,N_11928,N_11568);
nor U13886 (N_13886,N_11900,N_10413);
xnor U13887 (N_13887,N_10560,N_11914);
and U13888 (N_13888,N_11216,N_10198);
nor U13889 (N_13889,N_10929,N_10993);
nand U13890 (N_13890,N_10046,N_11308);
nor U13891 (N_13891,N_11563,N_11106);
nand U13892 (N_13892,N_11411,N_10293);
or U13893 (N_13893,N_11056,N_10514);
nor U13894 (N_13894,N_11427,N_11924);
or U13895 (N_13895,N_10962,N_10171);
nor U13896 (N_13896,N_10747,N_11661);
or U13897 (N_13897,N_11154,N_11629);
or U13898 (N_13898,N_10198,N_10880);
nand U13899 (N_13899,N_11693,N_11826);
nor U13900 (N_13900,N_10436,N_10540);
nor U13901 (N_13901,N_10834,N_11273);
or U13902 (N_13902,N_11033,N_10917);
nand U13903 (N_13903,N_10428,N_10107);
and U13904 (N_13904,N_10919,N_10871);
and U13905 (N_13905,N_10090,N_10163);
or U13906 (N_13906,N_10942,N_11920);
or U13907 (N_13907,N_10501,N_11073);
xnor U13908 (N_13908,N_11938,N_10181);
nor U13909 (N_13909,N_10496,N_11931);
or U13910 (N_13910,N_11718,N_11861);
or U13911 (N_13911,N_10732,N_10711);
or U13912 (N_13912,N_11829,N_11588);
nand U13913 (N_13913,N_11193,N_10084);
and U13914 (N_13914,N_10635,N_10749);
nand U13915 (N_13915,N_11744,N_10357);
or U13916 (N_13916,N_11500,N_11029);
or U13917 (N_13917,N_10470,N_10076);
nand U13918 (N_13918,N_10153,N_10535);
nand U13919 (N_13919,N_11230,N_10517);
nor U13920 (N_13920,N_10604,N_11307);
and U13921 (N_13921,N_11343,N_10709);
xnor U13922 (N_13922,N_10628,N_10993);
or U13923 (N_13923,N_11272,N_10300);
or U13924 (N_13924,N_11548,N_11854);
nor U13925 (N_13925,N_11443,N_10938);
nand U13926 (N_13926,N_10127,N_10834);
nand U13927 (N_13927,N_10340,N_11402);
nand U13928 (N_13928,N_10550,N_11942);
xor U13929 (N_13929,N_11182,N_10701);
nand U13930 (N_13930,N_11542,N_10415);
nor U13931 (N_13931,N_10279,N_10244);
or U13932 (N_13932,N_10060,N_11042);
or U13933 (N_13933,N_10443,N_11628);
nand U13934 (N_13934,N_10510,N_11672);
and U13935 (N_13935,N_11108,N_10630);
or U13936 (N_13936,N_11324,N_10604);
nor U13937 (N_13937,N_10251,N_11594);
and U13938 (N_13938,N_10678,N_10327);
or U13939 (N_13939,N_10404,N_11507);
nand U13940 (N_13940,N_10096,N_11985);
nor U13941 (N_13941,N_10254,N_11360);
or U13942 (N_13942,N_10117,N_10382);
or U13943 (N_13943,N_10575,N_10986);
nand U13944 (N_13944,N_11628,N_11253);
nand U13945 (N_13945,N_11872,N_11558);
or U13946 (N_13946,N_11359,N_11422);
nand U13947 (N_13947,N_10281,N_11416);
nand U13948 (N_13948,N_10972,N_11942);
and U13949 (N_13949,N_10647,N_10948);
xor U13950 (N_13950,N_10143,N_11271);
nor U13951 (N_13951,N_11834,N_10278);
nor U13952 (N_13952,N_10849,N_11197);
and U13953 (N_13953,N_10747,N_10736);
and U13954 (N_13954,N_11631,N_11901);
or U13955 (N_13955,N_11266,N_10802);
nand U13956 (N_13956,N_11765,N_10486);
nand U13957 (N_13957,N_10029,N_11602);
nand U13958 (N_13958,N_10165,N_11699);
nor U13959 (N_13959,N_10335,N_11180);
nor U13960 (N_13960,N_10722,N_10750);
nor U13961 (N_13961,N_10563,N_10387);
xor U13962 (N_13962,N_10834,N_10635);
nor U13963 (N_13963,N_11537,N_10499);
nand U13964 (N_13964,N_10032,N_10617);
nor U13965 (N_13965,N_11700,N_11379);
nor U13966 (N_13966,N_11521,N_10821);
nor U13967 (N_13967,N_10004,N_10544);
nand U13968 (N_13968,N_11054,N_10053);
nand U13969 (N_13969,N_11340,N_10239);
and U13970 (N_13970,N_10936,N_10433);
xor U13971 (N_13971,N_11743,N_11227);
nor U13972 (N_13972,N_11095,N_11692);
or U13973 (N_13973,N_10327,N_10593);
nand U13974 (N_13974,N_11272,N_10880);
nand U13975 (N_13975,N_10579,N_11587);
nand U13976 (N_13976,N_11323,N_11486);
nor U13977 (N_13977,N_11295,N_11117);
and U13978 (N_13978,N_11164,N_10064);
and U13979 (N_13979,N_10155,N_10347);
nor U13980 (N_13980,N_10525,N_11061);
nand U13981 (N_13981,N_10720,N_10155);
or U13982 (N_13982,N_10052,N_11005);
and U13983 (N_13983,N_11263,N_10935);
nand U13984 (N_13984,N_10165,N_10564);
xnor U13985 (N_13985,N_10048,N_10567);
and U13986 (N_13986,N_10464,N_10910);
or U13987 (N_13987,N_10516,N_11614);
and U13988 (N_13988,N_11679,N_10868);
and U13989 (N_13989,N_11791,N_10512);
or U13990 (N_13990,N_10430,N_10009);
or U13991 (N_13991,N_10662,N_11981);
or U13992 (N_13992,N_10716,N_11331);
and U13993 (N_13993,N_10566,N_10277);
xor U13994 (N_13994,N_10466,N_11263);
nand U13995 (N_13995,N_10900,N_10207);
and U13996 (N_13996,N_10576,N_10897);
or U13997 (N_13997,N_10902,N_10341);
nor U13998 (N_13998,N_10511,N_11242);
nand U13999 (N_13999,N_11632,N_10742);
and U14000 (N_14000,N_12391,N_13176);
or U14001 (N_14001,N_13410,N_13085);
and U14002 (N_14002,N_12564,N_13451);
or U14003 (N_14003,N_12197,N_12857);
nor U14004 (N_14004,N_12121,N_13734);
or U14005 (N_14005,N_13735,N_12575);
nor U14006 (N_14006,N_13530,N_13387);
or U14007 (N_14007,N_13098,N_13415);
and U14008 (N_14008,N_13532,N_12210);
xor U14009 (N_14009,N_13980,N_12088);
and U14010 (N_14010,N_12383,N_12682);
xor U14011 (N_14011,N_13761,N_12450);
nand U14012 (N_14012,N_13611,N_12980);
nand U14013 (N_14013,N_12590,N_12619);
xnor U14014 (N_14014,N_13405,N_13135);
nor U14015 (N_14015,N_12139,N_13153);
nand U14016 (N_14016,N_13615,N_13445);
nor U14017 (N_14017,N_13575,N_12530);
nor U14018 (N_14018,N_13065,N_12111);
nor U14019 (N_14019,N_12021,N_12230);
or U14020 (N_14020,N_12705,N_12563);
or U14021 (N_14021,N_12870,N_12819);
xnor U14022 (N_14022,N_12908,N_12712);
and U14023 (N_14023,N_12262,N_12739);
and U14024 (N_14024,N_13378,N_13221);
and U14025 (N_14025,N_13740,N_13330);
or U14026 (N_14026,N_13016,N_12919);
nor U14027 (N_14027,N_13897,N_12834);
nand U14028 (N_14028,N_12978,N_12370);
nand U14029 (N_14029,N_12580,N_12814);
nand U14030 (N_14030,N_12104,N_12767);
nand U14031 (N_14031,N_13909,N_12124);
and U14032 (N_14032,N_12985,N_12611);
xor U14033 (N_14033,N_12146,N_13170);
nand U14034 (N_14034,N_12656,N_12764);
and U14035 (N_14035,N_12147,N_13797);
and U14036 (N_14036,N_13296,N_13664);
nand U14037 (N_14037,N_12500,N_12892);
or U14038 (N_14038,N_12244,N_12482);
nand U14039 (N_14039,N_13419,N_12367);
nor U14040 (N_14040,N_13268,N_13137);
nand U14041 (N_14041,N_12013,N_13332);
nand U14042 (N_14042,N_12159,N_13516);
and U14043 (N_14043,N_12950,N_12792);
or U14044 (N_14044,N_12079,N_13235);
nor U14045 (N_14045,N_12898,N_13524);
nand U14046 (N_14046,N_13818,N_12969);
nor U14047 (N_14047,N_13705,N_13787);
or U14048 (N_14048,N_13109,N_13527);
and U14049 (N_14049,N_13113,N_12699);
and U14050 (N_14050,N_12650,N_12274);
and U14051 (N_14051,N_13878,N_12377);
or U14052 (N_14052,N_12382,N_12700);
or U14053 (N_14053,N_13219,N_12544);
and U14054 (N_14054,N_13630,N_13793);
or U14055 (N_14055,N_13783,N_13713);
nor U14056 (N_14056,N_12502,N_12306);
nand U14057 (N_14057,N_12279,N_13188);
xor U14058 (N_14058,N_12489,N_12932);
nand U14059 (N_14059,N_13782,N_12976);
nand U14060 (N_14060,N_13964,N_12490);
and U14061 (N_14061,N_13968,N_12223);
and U14062 (N_14062,N_13139,N_12505);
nand U14063 (N_14063,N_12901,N_13181);
and U14064 (N_14064,N_13939,N_13059);
and U14065 (N_14065,N_12518,N_13003);
nor U14066 (N_14066,N_13839,N_13376);
xor U14067 (N_14067,N_13313,N_13895);
nand U14068 (N_14068,N_12368,N_13609);
xor U14069 (N_14069,N_12143,N_13066);
xor U14070 (N_14070,N_12430,N_13600);
or U14071 (N_14071,N_13730,N_13351);
nand U14072 (N_14072,N_13894,N_13288);
xor U14073 (N_14073,N_13222,N_13256);
xnor U14074 (N_14074,N_13916,N_12278);
xor U14075 (N_14075,N_13820,N_13438);
nor U14076 (N_14076,N_12869,N_12059);
or U14077 (N_14077,N_12192,N_12707);
nor U14078 (N_14078,N_12228,N_12484);
nor U14079 (N_14079,N_13463,N_13460);
nor U14080 (N_14080,N_12053,N_12584);
and U14081 (N_14081,N_13294,N_12045);
and U14082 (N_14082,N_12636,N_12273);
and U14083 (N_14083,N_13739,N_13996);
nor U14084 (N_14084,N_13110,N_13197);
nand U14085 (N_14085,N_13473,N_13537);
xnor U14086 (N_14086,N_12922,N_13815);
and U14087 (N_14087,N_13727,N_13622);
or U14088 (N_14088,N_12878,N_12661);
nor U14089 (N_14089,N_12338,N_13706);
nand U14090 (N_14090,N_12441,N_12763);
and U14091 (N_14091,N_12945,N_12158);
or U14092 (N_14092,N_12649,N_12001);
nand U14093 (N_14093,N_12182,N_12145);
nand U14094 (N_14094,N_12125,N_12588);
or U14095 (N_14095,N_13765,N_13464);
nand U14096 (N_14096,N_12780,N_12481);
nand U14097 (N_14097,N_13425,N_12290);
nand U14098 (N_14098,N_13645,N_12188);
nand U14099 (N_14099,N_13114,N_12187);
and U14100 (N_14100,N_13206,N_12536);
nor U14101 (N_14101,N_12073,N_13928);
nand U14102 (N_14102,N_12690,N_13062);
nor U14103 (N_14103,N_13407,N_12810);
nand U14104 (N_14104,N_13886,N_13444);
nor U14105 (N_14105,N_13619,N_13041);
xnor U14106 (N_14106,N_12806,N_12291);
or U14107 (N_14107,N_12170,N_12305);
nor U14108 (N_14108,N_12300,N_12087);
xnor U14109 (N_14109,N_13970,N_12548);
nand U14110 (N_14110,N_13273,N_12746);
or U14111 (N_14111,N_12742,N_13014);
or U14112 (N_14112,N_13323,N_12222);
nor U14113 (N_14113,N_12349,N_13573);
or U14114 (N_14114,N_12421,N_13890);
nor U14115 (N_14115,N_13690,N_13339);
and U14116 (N_14116,N_12123,N_13564);
or U14117 (N_14117,N_13678,N_12164);
nand U14118 (N_14118,N_12628,N_12555);
nand U14119 (N_14119,N_12108,N_12981);
nand U14120 (N_14120,N_13314,N_12473);
nand U14121 (N_14121,N_12102,N_12875);
nand U14122 (N_14122,N_13060,N_13321);
nand U14123 (N_14123,N_13480,N_12836);
and U14124 (N_14124,N_12256,N_12779);
and U14125 (N_14125,N_12783,N_12352);
or U14126 (N_14126,N_13354,N_12497);
nand U14127 (N_14127,N_13311,N_13079);
or U14128 (N_14128,N_12406,N_12698);
and U14129 (N_14129,N_13251,N_13724);
nor U14130 (N_14130,N_12292,N_12024);
or U14131 (N_14131,N_12596,N_13819);
nor U14132 (N_14132,N_13493,N_13603);
or U14133 (N_14133,N_12852,N_12521);
xor U14134 (N_14134,N_12748,N_12949);
nor U14135 (N_14135,N_12299,N_13394);
and U14136 (N_14136,N_13649,N_12671);
nand U14137 (N_14137,N_12016,N_13566);
nor U14138 (N_14138,N_12612,N_13809);
nand U14139 (N_14139,N_13501,N_13398);
and U14140 (N_14140,N_13495,N_13048);
or U14141 (N_14141,N_13057,N_13164);
nand U14142 (N_14142,N_12689,N_12265);
or U14143 (N_14143,N_13174,N_12263);
or U14144 (N_14144,N_12941,N_12466);
and U14145 (N_14145,N_12409,N_12952);
or U14146 (N_14146,N_12847,N_13371);
and U14147 (N_14147,N_12327,N_12601);
or U14148 (N_14148,N_13402,N_12178);
nor U14149 (N_14149,N_12736,N_13917);
xor U14150 (N_14150,N_13190,N_13353);
or U14151 (N_14151,N_13610,N_12692);
or U14152 (N_14152,N_12082,N_13310);
and U14153 (N_14153,N_12965,N_12328);
or U14154 (N_14154,N_13904,N_13281);
or U14155 (N_14155,N_13274,N_13557);
and U14156 (N_14156,N_12851,N_13008);
nand U14157 (N_14157,N_12993,N_12660);
nand U14158 (N_14158,N_12303,N_12740);
or U14159 (N_14159,N_12030,N_12090);
nand U14160 (N_14160,N_13150,N_13364);
nor U14161 (N_14161,N_13467,N_12253);
xor U14162 (N_14162,N_13350,N_13806);
or U14163 (N_14163,N_13414,N_13335);
nor U14164 (N_14164,N_13101,N_12591);
and U14165 (N_14165,N_13726,N_13831);
or U14166 (N_14166,N_13020,N_12522);
nand U14167 (N_14167,N_13342,N_12051);
or U14168 (N_14168,N_13266,N_13978);
nor U14169 (N_14169,N_13331,N_12238);
or U14170 (N_14170,N_13112,N_12854);
or U14171 (N_14171,N_13363,N_12936);
and U14172 (N_14172,N_13952,N_12116);
nor U14173 (N_14173,N_12618,N_12958);
nand U14174 (N_14174,N_12859,N_12570);
nand U14175 (N_14175,N_13182,N_13036);
nor U14176 (N_14176,N_13319,N_13312);
or U14177 (N_14177,N_12982,N_12943);
nor U14178 (N_14178,N_13659,N_13064);
nor U14179 (N_14179,N_12236,N_12597);
nand U14180 (N_14180,N_12003,N_13618);
xnor U14181 (N_14181,N_13393,N_13748);
and U14182 (N_14182,N_12647,N_13992);
or U14183 (N_14183,N_12297,N_12755);
nor U14184 (N_14184,N_13116,N_13111);
and U14185 (N_14185,N_13729,N_13867);
or U14186 (N_14186,N_12662,N_13237);
and U14187 (N_14187,N_12100,N_13853);
nor U14188 (N_14188,N_13923,N_13503);
xnor U14189 (N_14189,N_13033,N_12678);
and U14190 (N_14190,N_13644,N_13198);
xnor U14191 (N_14191,N_13650,N_12224);
and U14192 (N_14192,N_12302,N_13544);
and U14193 (N_14193,N_12702,N_12239);
nand U14194 (N_14194,N_13329,N_13902);
or U14195 (N_14195,N_13490,N_12405);
nand U14196 (N_14196,N_13333,N_13680);
and U14197 (N_14197,N_12160,N_13800);
nand U14198 (N_14198,N_13590,N_12453);
nor U14199 (N_14199,N_13519,N_13648);
xor U14200 (N_14200,N_13594,N_12757);
or U14201 (N_14201,N_13234,N_13750);
or U14202 (N_14202,N_12358,N_13891);
or U14203 (N_14203,N_13443,N_12670);
or U14204 (N_14204,N_13756,N_12110);
and U14205 (N_14205,N_12944,N_12663);
xnor U14206 (N_14206,N_13143,N_13187);
or U14207 (N_14207,N_13122,N_12371);
or U14208 (N_14208,N_13391,N_12876);
nor U14209 (N_14209,N_13465,N_13699);
nand U14210 (N_14210,N_13986,N_13427);
nor U14211 (N_14211,N_13998,N_13293);
and U14212 (N_14212,N_12495,N_13720);
and U14213 (N_14213,N_13944,N_13432);
or U14214 (N_14214,N_12275,N_12773);
or U14215 (N_14215,N_12803,N_13587);
and U14216 (N_14216,N_13439,N_13869);
nor U14217 (N_14217,N_13366,N_13966);
and U14218 (N_14218,N_12259,N_12267);
nand U14219 (N_14219,N_12434,N_12479);
and U14220 (N_14220,N_12823,N_13924);
nand U14221 (N_14221,N_12799,N_13226);
or U14222 (N_14222,N_13933,N_13441);
nand U14223 (N_14223,N_12133,N_12269);
and U14224 (N_14224,N_13022,N_13728);
or U14225 (N_14225,N_13982,N_12821);
and U14226 (N_14226,N_12173,N_12233);
nand U14227 (N_14227,N_13192,N_13517);
and U14228 (N_14228,N_12510,N_13055);
nor U14229 (N_14229,N_12042,N_12753);
nor U14230 (N_14230,N_13259,N_12545);
and U14231 (N_14231,N_12499,N_13086);
or U14232 (N_14232,N_13795,N_13478);
or U14233 (N_14233,N_12568,N_12390);
or U14234 (N_14234,N_12861,N_12728);
nand U14235 (N_14235,N_13934,N_13299);
nand U14236 (N_14236,N_12048,N_13951);
nand U14237 (N_14237,N_13956,N_12156);
or U14238 (N_14238,N_12750,N_13858);
nand U14239 (N_14239,N_12401,N_13863);
xor U14240 (N_14240,N_13344,N_13225);
and U14241 (N_14241,N_13384,N_12389);
and U14242 (N_14242,N_13668,N_12150);
or U14243 (N_14243,N_12720,N_12828);
or U14244 (N_14244,N_12282,N_13042);
xnor U14245 (N_14245,N_13262,N_12056);
xor U14246 (N_14246,N_12218,N_12986);
or U14247 (N_14247,N_12883,N_13882);
or U14248 (N_14248,N_13211,N_13385);
or U14249 (N_14249,N_13263,N_13334);
nand U14250 (N_14250,N_13682,N_12062);
nor U14251 (N_14251,N_12415,N_13798);
nor U14252 (N_14252,N_12659,N_12622);
or U14253 (N_14253,N_13741,N_13861);
xnor U14254 (N_14254,N_13301,N_12397);
and U14255 (N_14255,N_12380,N_12846);
and U14256 (N_14256,N_13272,N_12900);
or U14257 (N_14257,N_12906,N_13687);
and U14258 (N_14258,N_12557,N_13477);
or U14259 (N_14259,N_13302,N_12805);
and U14260 (N_14260,N_12953,N_12395);
xor U14261 (N_14261,N_13083,N_12142);
nand U14262 (N_14262,N_13777,N_12446);
or U14263 (N_14263,N_13812,N_13635);
and U14264 (N_14264,N_12507,N_13808);
and U14265 (N_14265,N_12054,N_12573);
nand U14266 (N_14266,N_12762,N_13096);
nand U14267 (N_14267,N_13718,N_12138);
nor U14268 (N_14268,N_13614,N_12934);
or U14269 (N_14269,N_12019,N_13571);
or U14270 (N_14270,N_13077,N_13838);
nor U14271 (N_14271,N_13922,N_13579);
or U14272 (N_14272,N_12768,N_12185);
nor U14273 (N_14273,N_13128,N_12938);
nand U14274 (N_14274,N_13044,N_13759);
or U14275 (N_14275,N_13358,N_12988);
nand U14276 (N_14276,N_12798,N_13429);
xnor U14277 (N_14277,N_12057,N_12340);
or U14278 (N_14278,N_12560,N_12344);
or U14279 (N_14279,N_12322,N_13565);
or U14280 (N_14280,N_12576,N_12926);
and U14281 (N_14281,N_12411,N_13873);
or U14282 (N_14282,N_13762,N_13859);
nor U14283 (N_14283,N_12227,N_13217);
or U14284 (N_14284,N_13534,N_13141);
nand U14285 (N_14285,N_12250,N_12475);
nand U14286 (N_14286,N_12315,N_12726);
and U14287 (N_14287,N_12927,N_12963);
nand U14288 (N_14288,N_13269,N_12891);
or U14289 (N_14289,N_12716,N_12996);
or U14290 (N_14290,N_12688,N_12168);
nand U14291 (N_14291,N_13854,N_13608);
nor U14292 (N_14292,N_13860,N_13686);
nand U14293 (N_14293,N_12888,N_12913);
nand U14294 (N_14294,N_12141,N_13291);
and U14295 (N_14295,N_13675,N_13658);
or U14296 (N_14296,N_12119,N_12071);
and U14297 (N_14297,N_13071,N_12418);
and U14298 (N_14298,N_12211,N_12258);
or U14299 (N_14299,N_13169,N_13390);
nand U14300 (N_14300,N_12684,N_12089);
nor U14301 (N_14301,N_13108,N_12072);
nor U14302 (N_14302,N_13813,N_13521);
nor U14303 (N_14303,N_12915,N_12533);
or U14304 (N_14304,N_12640,N_12838);
nand U14305 (N_14305,N_12594,N_12766);
nand U14306 (N_14306,N_12171,N_13758);
nor U14307 (N_14307,N_12330,N_13504);
and U14308 (N_14308,N_13006,N_12445);
or U14309 (N_14309,N_12527,N_12665);
xor U14310 (N_14310,N_12179,N_13957);
nand U14311 (N_14311,N_12078,N_13577);
nor U14312 (N_14312,N_13560,N_13123);
and U14313 (N_14313,N_13037,N_13136);
or U14314 (N_14314,N_13975,N_12216);
nor U14315 (N_14315,N_12646,N_12586);
nand U14316 (N_14316,N_13243,N_12027);
nor U14317 (N_14317,N_12680,N_13732);
nor U14318 (N_14318,N_13877,N_12261);
or U14319 (N_14319,N_12975,N_13367);
nor U14320 (N_14320,N_13945,N_13612);
nor U14321 (N_14321,N_12751,N_12165);
nand U14322 (N_14322,N_12874,N_13155);
or U14323 (N_14323,N_13639,N_13487);
nand U14324 (N_14324,N_13160,N_13948);
and U14325 (N_14325,N_13595,N_12129);
xor U14326 (N_14326,N_12283,N_13663);
nor U14327 (N_14327,N_13715,N_13196);
nand U14328 (N_14328,N_12558,N_13545);
nand U14329 (N_14329,N_12225,N_13242);
nor U14330 (N_14330,N_12077,N_12924);
and U14331 (N_14331,N_12339,N_12569);
or U14332 (N_14332,N_12356,N_12971);
nand U14333 (N_14333,N_12691,N_12882);
nor U14334 (N_14334,N_12960,N_13885);
nand U14335 (N_14335,N_12643,N_13855);
and U14336 (N_14336,N_12206,N_12504);
and U14337 (N_14337,N_12333,N_13409);
or U14338 (N_14338,N_13010,N_13498);
nor U14339 (N_14339,N_12137,N_13736);
xor U14340 (N_14340,N_12458,N_13320);
nand U14341 (N_14341,N_12542,N_13670);
nand U14342 (N_14342,N_13814,N_13757);
xor U14343 (N_14343,N_13983,N_12935);
xnor U14344 (N_14344,N_12342,N_13584);
or U14345 (N_14345,N_13803,N_12581);
and U14346 (N_14346,N_13624,N_13442);
or U14347 (N_14347,N_13623,N_13872);
or U14348 (N_14348,N_12106,N_13078);
nor U14349 (N_14349,N_13397,N_12324);
nand U14350 (N_14350,N_12967,N_13195);
nand U14351 (N_14351,N_13834,N_13850);
or U14352 (N_14352,N_13823,N_12651);
and U14353 (N_14353,N_12193,N_13954);
and U14354 (N_14354,N_12134,N_13248);
or U14355 (N_14355,N_12839,N_12719);
nor U14356 (N_14356,N_12709,N_12589);
nand U14357 (N_14357,N_13275,N_12005);
or U14358 (N_14358,N_12268,N_13851);
xor U14359 (N_14359,N_12131,N_13911);
and U14360 (N_14360,N_13961,N_13840);
nand U14361 (N_14361,N_13989,N_13025);
and U14362 (N_14362,N_12972,N_12610);
or U14363 (N_14363,N_13238,N_13901);
and U14364 (N_14364,N_12345,N_13028);
and U14365 (N_14365,N_12229,N_12373);
and U14366 (N_14366,N_12508,N_13893);
and U14367 (N_14367,N_13172,N_12697);
xor U14368 (N_14368,N_13270,N_12863);
nor U14369 (N_14369,N_12737,N_13063);
nand U14370 (N_14370,N_13280,N_13383);
or U14371 (N_14371,N_13514,N_13540);
or U14372 (N_14372,N_13475,N_13203);
and U14373 (N_14373,N_12872,N_13697);
and U14374 (N_14374,N_13026,N_12459);
nand U14375 (N_14375,N_13349,N_13550);
xnor U14376 (N_14376,N_13969,N_12701);
and U14377 (N_14377,N_13636,N_12826);
nand U14378 (N_14378,N_13142,N_13486);
and U14379 (N_14379,N_12365,N_12744);
nor U14380 (N_14380,N_13186,N_12868);
nand U14381 (N_14381,N_13159,N_13596);
or U14382 (N_14382,N_13535,N_13133);
or U14383 (N_14383,N_13348,N_12885);
nand U14384 (N_14384,N_13709,N_13529);
and U14385 (N_14385,N_13087,N_12451);
nand U14386 (N_14386,N_12687,N_12644);
or U14387 (N_14387,N_13708,N_13552);
nor U14388 (N_14388,N_13254,N_13082);
and U14389 (N_14389,N_13888,N_12007);
nand U14390 (N_14390,N_13396,N_13202);
xor U14391 (N_14391,N_13693,N_13346);
nor U14392 (N_14392,N_12970,N_13990);
nor U14393 (N_14393,N_13215,N_12990);
xor U14394 (N_14394,N_13892,N_12956);
and U14395 (N_14395,N_13661,N_12896);
and U14396 (N_14396,N_13528,N_12918);
nand U14397 (N_14397,N_12422,N_13640);
xor U14398 (N_14398,N_13887,N_12832);
or U14399 (N_14399,N_13583,N_13775);
or U14400 (N_14400,N_13147,N_12673);
xnor U14401 (N_14401,N_13868,N_12582);
nand U14402 (N_14402,N_12562,N_13488);
and U14403 (N_14403,N_13337,N_13286);
nand U14404 (N_14404,N_12176,N_12068);
nand U14405 (N_14405,N_12621,N_13052);
nor U14406 (N_14406,N_13375,N_12317);
and U14407 (N_14407,N_12652,N_13841);
or U14408 (N_14408,N_12811,N_13536);
nor U14409 (N_14409,N_13880,N_13290);
or U14410 (N_14410,N_12703,N_13449);
nand U14411 (N_14411,N_12378,N_13771);
and U14412 (N_14412,N_12633,N_12234);
nor U14413 (N_14413,N_13903,N_13070);
or U14414 (N_14414,N_13184,N_13669);
nand U14415 (N_14415,N_12733,N_12392);
or U14416 (N_14416,N_12135,N_13688);
or U14417 (N_14417,N_12237,N_13011);
or U14418 (N_14418,N_13345,N_12055);
or U14419 (N_14419,N_12122,N_13258);
or U14420 (N_14420,N_13769,N_12483);
and U14421 (N_14421,N_13481,N_12022);
and U14422 (N_14422,N_13742,N_12132);
or U14423 (N_14423,N_13325,N_12921);
xor U14424 (N_14424,N_13279,N_12402);
nand U14425 (N_14425,N_12784,N_12221);
nand U14426 (N_14426,N_12093,N_12000);
and U14427 (N_14427,N_13817,N_13586);
and U14428 (N_14428,N_13714,N_12075);
nand U14429 (N_14429,N_12512,N_12860);
and U14430 (N_14430,N_12095,N_12052);
and U14431 (N_14431,N_12487,N_13666);
nand U14432 (N_14432,N_12815,N_13788);
or U14433 (N_14433,N_12532,N_12528);
nor U14434 (N_14434,N_12749,N_12770);
nor U14435 (N_14435,N_12220,N_12722);
xor U14436 (N_14436,N_13165,N_13090);
nand U14437 (N_14437,N_13205,N_13352);
xnor U14438 (N_14438,N_12332,N_13471);
nor U14439 (N_14439,N_12894,N_12476);
or U14440 (N_14440,N_12552,N_12020);
nor U14441 (N_14441,N_13204,N_12477);
and U14442 (N_14442,N_12759,N_12127);
nor U14443 (N_14443,N_12280,N_13326);
nor U14444 (N_14444,N_12272,N_12028);
and U14445 (N_14445,N_12669,N_12091);
nand U14446 (N_14446,N_12494,N_13479);
nand U14447 (N_14447,N_13921,N_13252);
nor U14448 (N_14448,N_12404,N_13355);
or U14449 (N_14449,N_12714,N_13826);
xnor U14450 (N_14450,N_13412,N_13031);
nor U14451 (N_14451,N_13870,N_12658);
and U14452 (N_14452,N_12008,N_12947);
nand U14453 (N_14453,N_12795,N_13068);
and U14454 (N_14454,N_13450,N_12668);
or U14455 (N_14455,N_12706,N_13620);
xor U14456 (N_14456,N_13553,N_12565);
or U14457 (N_14457,N_12103,N_13685);
nor U14458 (N_14458,N_12710,N_12181);
or U14459 (N_14459,N_13546,N_13074);
nand U14460 (N_14460,N_12999,N_13949);
or U14461 (N_14461,N_12252,N_12765);
and U14462 (N_14462,N_12353,N_13656);
nand U14463 (N_14463,N_13703,N_13462);
and U14464 (N_14464,N_13925,N_12964);
nor U14465 (N_14465,N_13510,N_12226);
nor U14466 (N_14466,N_12105,N_13027);
and U14467 (N_14467,N_13781,N_12567);
or U14468 (N_14468,N_12511,N_12928);
nor U14469 (N_14469,N_12524,N_12554);
xor U14470 (N_14470,N_13760,N_12336);
or U14471 (N_14471,N_12480,N_13030);
nor U14472 (N_14472,N_13124,N_12498);
nand U14473 (N_14473,N_12114,N_12249);
nand U14474 (N_14474,N_12592,N_12912);
xnor U14475 (N_14475,N_13844,N_12136);
and U14476 (N_14476,N_13569,N_13874);
nand U14477 (N_14477,N_13733,N_12468);
nor U14478 (N_14478,N_13131,N_13167);
xnor U14479 (N_14479,N_12412,N_13175);
and U14480 (N_14480,N_13846,N_12471);
nor U14481 (N_14481,N_12616,N_12191);
nand U14482 (N_14482,N_13454,N_13810);
or U14483 (N_14483,N_12295,N_13214);
or U14484 (N_14484,N_13896,N_13912);
nor U14485 (N_14485,N_12066,N_12350);
xnor U14486 (N_14486,N_13754,N_13621);
or U14487 (N_14487,N_12989,N_12357);
or U14488 (N_14488,N_12550,N_13357);
nor U14489 (N_14489,N_12432,N_12424);
nand U14490 (N_14490,N_13738,N_12410);
nor U14491 (N_14491,N_13513,N_12664);
nand U14492 (N_14492,N_12531,N_12676);
nor U14493 (N_14493,N_13499,N_13694);
and U14494 (N_14494,N_13606,N_12977);
nor U14495 (N_14495,N_12856,N_12169);
and U14496 (N_14496,N_12070,N_13317);
or U14497 (N_14497,N_12437,N_13837);
nor U14498 (N_14498,N_12693,N_13081);
nor U14499 (N_14499,N_13930,N_12516);
xnor U14500 (N_14500,N_13145,N_13300);
nor U14501 (N_14501,N_13199,N_12496);
xor U14502 (N_14502,N_12318,N_13240);
nand U14503 (N_14503,N_12625,N_13072);
and U14504 (N_14504,N_12172,N_12825);
and U14505 (N_14505,N_12630,N_12440);
or U14506 (N_14506,N_12820,N_13725);
nor U14507 (N_14507,N_12320,N_12376);
nor U14508 (N_14508,N_12148,N_12509);
nand U14509 (N_14509,N_12893,N_12004);
nor U14510 (N_14510,N_12895,N_13991);
and U14511 (N_14511,N_13431,N_13825);
and U14512 (N_14512,N_13395,N_13864);
and U14513 (N_14513,N_13768,N_13701);
nand U14514 (N_14514,N_12175,N_12384);
nand U14515 (N_14515,N_12667,N_12152);
nand U14516 (N_14516,N_12923,N_13960);
nand U14517 (N_14517,N_12775,N_12540);
or U14518 (N_14518,N_12890,N_12506);
or U14519 (N_14519,N_12571,N_12843);
or U14520 (N_14520,N_12448,N_13277);
nor U14521 (N_14521,N_13264,N_12974);
xor U14522 (N_14522,N_13436,N_12735);
and U14523 (N_14523,N_12065,N_13763);
nor U14524 (N_14524,N_12011,N_12312);
nand U14525 (N_14525,N_12623,N_12802);
nor U14526 (N_14526,N_13794,N_13018);
nand U14527 (N_14527,N_12771,N_13149);
nor U14528 (N_14528,N_13328,N_13657);
nor U14529 (N_14529,N_12002,N_12493);
nand U14530 (N_14530,N_13413,N_13336);
xor U14531 (N_14531,N_12617,N_13447);
and U14532 (N_14532,N_13613,N_13505);
or U14533 (N_14533,N_13570,N_13148);
nand U14534 (N_14534,N_13216,N_13001);
or U14535 (N_14535,N_13843,N_13588);
or U14536 (N_14536,N_12155,N_12653);
nand U14537 (N_14537,N_12217,N_13856);
and U14538 (N_14538,N_13056,N_12523);
and U14539 (N_14539,N_12323,N_12313);
nor U14540 (N_14540,N_12118,N_13946);
and U14541 (N_14541,N_13097,N_12727);
nor U14542 (N_14542,N_13700,N_13404);
nand U14543 (N_14543,N_13899,N_12015);
or U14544 (N_14544,N_13012,N_12049);
nand U14545 (N_14545,N_13824,N_13852);
nand U14546 (N_14546,N_12879,N_12423);
xor U14547 (N_14547,N_12973,N_12427);
xor U14548 (N_14548,N_12645,N_13241);
or U14549 (N_14549,N_13972,N_12032);
nand U14550 (N_14550,N_12606,N_12696);
or U14551 (N_14551,N_12388,N_13024);
or U14552 (N_14552,N_12801,N_12354);
nand U14553 (N_14553,N_12271,N_13589);
nor U14554 (N_14554,N_12807,N_12128);
nand U14555 (N_14555,N_13292,N_12264);
nand U14556 (N_14556,N_12648,N_13049);
or U14557 (N_14557,N_12425,N_13193);
nand U14558 (N_14558,N_13076,N_13549);
nand U14559 (N_14559,N_12429,N_13907);
nor U14560 (N_14560,N_13993,N_13261);
nand U14561 (N_14561,N_13561,N_12107);
and U14562 (N_14562,N_12608,N_13842);
or U14563 (N_14563,N_12513,N_13491);
nand U14564 (N_14564,N_12454,N_12064);
or U14565 (N_14565,N_13994,N_12627);
nand U14566 (N_14566,N_12130,N_12553);
nor U14567 (N_14567,N_13157,N_12240);
nor U14568 (N_14568,N_12364,N_12587);
nand U14569 (N_14569,N_12491,N_13338);
nor U14570 (N_14570,N_12101,N_13426);
nor U14571 (N_14571,N_12046,N_12478);
nand U14572 (N_14572,N_13433,N_13023);
nand U14573 (N_14573,N_12036,N_12578);
and U14574 (N_14574,N_12844,N_12871);
nor U14575 (N_14575,N_12385,N_12363);
or U14576 (N_14576,N_12822,N_12760);
nor U14577 (N_14577,N_13913,N_13179);
nand U14578 (N_14578,N_13971,N_12235);
nor U14579 (N_14579,N_12154,N_12756);
nand U14580 (N_14580,N_13051,N_12257);
nand U14581 (N_14581,N_12449,N_13053);
nor U14582 (N_14582,N_13218,N_13629);
nand U14583 (N_14583,N_13672,N_12743);
and U14584 (N_14584,N_13093,N_13021);
and U14585 (N_14585,N_13973,N_13132);
nand U14586 (N_14586,N_13780,N_13652);
nor U14587 (N_14587,N_13616,N_13212);
or U14588 (N_14588,N_12774,N_12026);
and U14589 (N_14589,N_13602,N_13017);
nor U14590 (N_14590,N_13766,N_13283);
nand U14591 (N_14591,N_12162,N_13045);
nor U14592 (N_14592,N_13472,N_13963);
and U14593 (N_14593,N_12417,N_13035);
nand U14594 (N_14594,N_13107,N_13876);
and U14595 (N_14595,N_13009,N_12247);
nor U14596 (N_14596,N_13926,N_13828);
or U14597 (N_14597,N_13497,N_13400);
nand U14598 (N_14598,N_13526,N_12215);
and U14599 (N_14599,N_13180,N_13653);
nand U14600 (N_14600,N_12629,N_13642);
or U14601 (N_14601,N_12600,N_12827);
and U14602 (N_14602,N_12745,N_13702);
and U14603 (N_14603,N_12747,N_13908);
and U14604 (N_14604,N_13434,N_13191);
and U14605 (N_14605,N_13435,N_13667);
nor U14606 (N_14606,N_12685,N_13919);
nor U14607 (N_14607,N_13731,N_13054);
xor U14608 (N_14608,N_12679,N_13168);
or U14609 (N_14609,N_13717,N_13255);
and U14610 (N_14610,N_13201,N_12902);
nor U14611 (N_14611,N_12808,N_13297);
or U14612 (N_14612,N_13470,N_13029);
or U14613 (N_14613,N_13126,N_13104);
and U14614 (N_14614,N_13744,N_13559);
or U14615 (N_14615,N_13785,N_13643);
nor U14616 (N_14616,N_12301,N_13977);
nor U14617 (N_14617,N_13307,N_12599);
nand U14618 (N_14618,N_12374,N_13633);
nor U14619 (N_14619,N_13095,N_12833);
nand U14620 (N_14620,N_13941,N_12288);
nand U14621 (N_14621,N_13257,N_12060);
and U14622 (N_14622,N_12800,N_12294);
and U14623 (N_14623,N_13089,N_12866);
nand U14624 (N_14624,N_12202,N_13173);
or U14625 (N_14625,N_12817,N_12341);
nor U14626 (N_14626,N_13340,N_13073);
nand U14627 (N_14627,N_12204,N_12347);
xnor U14628 (N_14628,N_12905,N_13134);
nand U14629 (N_14629,N_13723,N_12438);
nor U14630 (N_14630,N_12704,N_13746);
or U14631 (N_14631,N_12602,N_13628);
and U14632 (N_14632,N_12166,N_12213);
nand U14633 (N_14633,N_12270,N_12515);
and U14634 (N_14634,N_13483,N_12190);
or U14635 (N_14635,N_12266,N_12526);
xnor U14636 (N_14636,N_13118,N_13711);
or U14637 (N_14637,N_12012,N_13563);
and U14638 (N_14638,N_13267,N_13452);
or U14639 (N_14639,N_13737,N_12683);
nand U14640 (N_14640,N_13625,N_12556);
nor U14641 (N_14641,N_12120,N_13210);
nand U14642 (N_14642,N_12797,N_12157);
xor U14643 (N_14643,N_13722,N_13361);
nand U14644 (N_14644,N_12607,N_13430);
and U14645 (N_14645,N_12713,N_12631);
nand U14646 (N_14646,N_12598,N_13651);
nand U14647 (N_14647,N_12566,N_13562);
nor U14648 (N_14648,N_13372,N_13306);
or U14649 (N_14649,N_12334,N_12031);
or U14650 (N_14650,N_12675,N_12387);
nor U14651 (N_14651,N_12848,N_12862);
and U14652 (N_14652,N_12804,N_12998);
nor U14653 (N_14653,N_12831,N_13509);
or U14654 (N_14654,N_12010,N_13692);
nor U14655 (N_14655,N_12251,N_12194);
nor U14656 (N_14656,N_13790,N_13551);
or U14657 (N_14657,N_13120,N_12375);
or U14658 (N_14658,N_13581,N_13898);
nor U14659 (N_14659,N_12177,N_13677);
xor U14660 (N_14660,N_12897,N_12463);
nand U14661 (N_14661,N_13224,N_13284);
or U14662 (N_14662,N_13500,N_13940);
xor U14663 (N_14663,N_12654,N_12925);
or U14664 (N_14664,N_13360,N_13848);
xor U14665 (N_14665,N_12325,N_13631);
and U14666 (N_14666,N_13654,N_13929);
and U14667 (N_14667,N_12254,N_12398);
nand U14668 (N_14668,N_13271,N_12951);
xor U14669 (N_14669,N_13161,N_12413);
and U14670 (N_14670,N_13368,N_12074);
and U14671 (N_14671,N_13572,N_13260);
nand U14672 (N_14672,N_12887,N_13647);
and U14673 (N_14673,N_13716,N_12583);
nand U14674 (N_14674,N_13002,N_13604);
or U14675 (N_14675,N_13200,N_13665);
nand U14676 (N_14676,N_13543,N_12529);
nand U14677 (N_14677,N_13322,N_12837);
or U14678 (N_14678,N_13105,N_13721);
nor U14679 (N_14679,N_13512,N_13632);
and U14680 (N_14680,N_12461,N_12433);
nand U14681 (N_14681,N_13712,N_12431);
xnor U14682 (N_14682,N_13247,N_13947);
or U14683 (N_14683,N_12098,N_13476);
or U14684 (N_14684,N_13796,N_12281);
or U14685 (N_14685,N_12731,N_13459);
nand U14686 (N_14686,N_12455,N_13671);
and U14687 (N_14687,N_13004,N_13229);
nand U14688 (N_14688,N_12585,N_13764);
or U14689 (N_14689,N_12609,N_13466);
nor U14690 (N_14690,N_12346,N_12626);
nor U14691 (N_14691,N_13423,N_12501);
or U14692 (N_14692,N_13719,N_12991);
nor U14693 (N_14693,N_13422,N_12782);
or U14694 (N_14694,N_12407,N_12083);
nor U14695 (N_14695,N_12316,N_12962);
and U14696 (N_14696,N_13100,N_13508);
and U14697 (N_14697,N_13936,N_12298);
and U14698 (N_14698,N_13518,N_13377);
nand U14699 (N_14699,N_12721,N_13879);
xor U14700 (N_14700,N_13138,N_13538);
and U14701 (N_14701,N_12937,N_13457);
nor U14702 (N_14702,N_12777,N_13511);
xor U14703 (N_14703,N_13213,N_13684);
nand U14704 (N_14704,N_13568,N_13558);
nor U14705 (N_14705,N_13318,N_13359);
or U14706 (N_14706,N_13626,N_12144);
and U14707 (N_14707,N_12242,N_12920);
nor U14708 (N_14708,N_12884,N_12789);
nor U14709 (N_14709,N_13755,N_13601);
or U14710 (N_14710,N_12914,N_12035);
nand U14711 (N_14711,N_12723,N_13324);
nor U14712 (N_14712,N_13347,N_12140);
xnor U14713 (N_14713,N_13784,N_13592);
xor U14714 (N_14714,N_12724,N_12574);
nor U14715 (N_14715,N_12907,N_12525);
nor U14716 (N_14716,N_12439,N_12219);
or U14717 (N_14717,N_13774,N_12708);
nor U14718 (N_14718,N_13231,N_12018);
nor U14719 (N_14719,N_13094,N_13389);
or U14720 (N_14720,N_13485,N_12039);
or U14721 (N_14721,N_12386,N_13959);
and U14722 (N_14722,N_13484,N_13931);
nor U14723 (N_14723,N_13305,N_13773);
and U14724 (N_14724,N_12979,N_12624);
nand U14725 (N_14725,N_13156,N_13249);
or U14726 (N_14726,N_13401,N_12308);
and U14727 (N_14727,N_13151,N_13791);
and U14728 (N_14728,N_12741,N_12604);
or U14729 (N_14729,N_12841,N_12205);
or U14730 (N_14730,N_12541,N_13239);
or U14731 (N_14731,N_13469,N_12293);
and U14732 (N_14732,N_12355,N_12209);
and U14733 (N_14733,N_13069,N_13683);
nand U14734 (N_14734,N_12520,N_12734);
or U14735 (N_14735,N_13468,N_13177);
nor U14736 (N_14736,N_13938,N_13278);
and U14737 (N_14737,N_12718,N_12196);
or U14738 (N_14738,N_13745,N_13289);
and U14739 (N_14739,N_12277,N_13163);
and U14740 (N_14740,N_12877,N_13038);
or U14741 (N_14741,N_13356,N_13821);
nor U14742 (N_14742,N_13786,N_12420);
and U14743 (N_14743,N_12248,N_13811);
nor U14744 (N_14744,N_13343,N_12809);
or U14745 (N_14745,N_13679,N_12099);
or U14746 (N_14746,N_12853,N_12472);
xor U14747 (N_14747,N_12058,N_12994);
and U14748 (N_14748,N_13767,N_12287);
and U14749 (N_14749,N_12539,N_13743);
or U14750 (N_14750,N_13129,N_12637);
xnor U14751 (N_14751,N_13080,N_12725);
or U14752 (N_14752,N_13845,N_13084);
nand U14753 (N_14753,N_12968,N_13520);
nor U14754 (N_14754,N_12639,N_12337);
xor U14755 (N_14755,N_12889,N_13574);
xor U14756 (N_14756,N_13776,N_12199);
nand U14757 (N_14757,N_12403,N_13556);
xnor U14758 (N_14758,N_13935,N_12014);
and U14759 (N_14759,N_13075,N_12711);
nand U14760 (N_14760,N_13875,N_12537);
nand U14761 (N_14761,N_12006,N_13220);
xnor U14762 (N_14762,N_13166,N_13802);
or U14763 (N_14763,N_13920,N_13121);
and U14764 (N_14764,N_12372,N_12881);
or U14765 (N_14765,N_12824,N_12180);
and U14766 (N_14766,N_12519,N_12435);
and U14767 (N_14767,N_13492,N_13531);
nor U14768 (N_14768,N_13953,N_13091);
nand U14769 (N_14769,N_12864,N_12517);
or U14770 (N_14770,N_12931,N_12715);
or U14771 (N_14771,N_12911,N_12400);
or U14772 (N_14772,N_12758,N_12635);
nand U14773 (N_14773,N_13236,N_13304);
nor U14774 (N_14774,N_13871,N_12034);
nor U14775 (N_14775,N_13627,N_12729);
and U14776 (N_14776,N_12260,N_13507);
nor U14777 (N_14777,N_13778,N_13130);
nand U14778 (N_14778,N_12304,N_12457);
xor U14779 (N_14779,N_13233,N_12289);
xnor U14780 (N_14780,N_12310,N_13411);
or U14781 (N_14781,N_12916,N_12984);
nor U14782 (N_14782,N_12781,N_12444);
and U14783 (N_14783,N_13995,N_13303);
and U14784 (N_14784,N_13370,N_13676);
nor U14785 (N_14785,N_13827,N_12009);
nand U14786 (N_14786,N_13833,N_13883);
and U14787 (N_14787,N_12394,N_12790);
and U14788 (N_14788,N_13067,N_13223);
nor U14789 (N_14789,N_12813,N_13927);
nand U14790 (N_14790,N_12577,N_13597);
nand U14791 (N_14791,N_12997,N_12452);
xnor U14792 (N_14792,N_13607,N_12436);
and U14793 (N_14793,N_13502,N_12085);
nand U14794 (N_14794,N_13585,N_13981);
nand U14795 (N_14795,N_12769,N_13707);
and U14796 (N_14796,N_12044,N_13747);
nand U14797 (N_14797,N_12954,N_12214);
nand U14798 (N_14798,N_12615,N_12942);
and U14799 (N_14799,N_12816,N_12241);
and U14800 (N_14800,N_13976,N_12910);
or U14801 (N_14801,N_13362,N_12603);
and U14802 (N_14802,N_13932,N_12428);
nand U14803 (N_14803,N_13578,N_13158);
and U14804 (N_14804,N_13900,N_13458);
and U14805 (N_14805,N_12677,N_13380);
or U14806 (N_14806,N_13374,N_12092);
or U14807 (N_14807,N_13034,N_13655);
nand U14808 (N_14808,N_12787,N_12948);
and U14809 (N_14809,N_13691,N_12666);
xor U14810 (N_14810,N_13695,N_12686);
xnor U14811 (N_14811,N_13847,N_13244);
xnor U14812 (N_14812,N_13789,N_12930);
nand U14813 (N_14813,N_12785,N_13421);
nand U14814 (N_14814,N_12348,N_12465);
nand U14815 (N_14815,N_13474,N_13541);
or U14816 (N_14816,N_13660,N_13987);
xor U14817 (N_14817,N_13593,N_12243);
and U14818 (N_14818,N_13144,N_13127);
nand U14819 (N_14819,N_12084,N_13040);
nor U14820 (N_14820,N_12189,N_13634);
xor U14821 (N_14821,N_12835,N_12321);
and U14822 (N_14822,N_13539,N_13061);
nand U14823 (N_14823,N_13772,N_13849);
xnor U14824 (N_14824,N_13555,N_12067);
or U14825 (N_14825,N_12360,N_13792);
or U14826 (N_14826,N_13388,N_12025);
nor U14827 (N_14827,N_13032,N_13779);
and U14828 (N_14828,N_12485,N_13617);
and U14829 (N_14829,N_13245,N_13282);
or U14830 (N_14830,N_13246,N_12917);
nor U14831 (N_14831,N_13937,N_12983);
nor U14832 (N_14832,N_13751,N_12393);
and U14833 (N_14833,N_13440,N_12366);
xor U14834 (N_14834,N_12761,N_12778);
nand U14835 (N_14835,N_13250,N_12207);
and U14836 (N_14836,N_13576,N_13816);
xor U14837 (N_14837,N_12867,N_12419);
xnor U14838 (N_14838,N_12231,N_12579);
nor U14839 (N_14839,N_13437,N_13494);
or U14840 (N_14840,N_13591,N_13985);
or U14841 (N_14841,N_13453,N_13194);
nand U14842 (N_14842,N_12642,N_12153);
or U14843 (N_14843,N_12309,N_13547);
or U14844 (N_14844,N_13988,N_13496);
or U14845 (N_14845,N_13386,N_13914);
and U14846 (N_14846,N_12559,N_12245);
and U14847 (N_14847,N_13208,N_13232);
nand U14848 (N_14848,N_12830,N_13865);
and U14849 (N_14849,N_13943,N_13013);
and U14850 (N_14850,N_12638,N_13308);
or U14851 (N_14851,N_13461,N_12063);
nand U14852 (N_14852,N_12314,N_12776);
and U14853 (N_14853,N_13102,N_12311);
nand U14854 (N_14854,N_12396,N_12381);
and U14855 (N_14855,N_13881,N_12561);
nor U14856 (N_14856,N_12029,N_13424);
or U14857 (N_14857,N_12903,N_13807);
and U14858 (N_14858,N_12362,N_13580);
and U14859 (N_14859,N_13207,N_13341);
or U14860 (N_14860,N_13408,N_12186);
xnor U14861 (N_14861,N_13152,N_12995);
and U14862 (N_14862,N_12041,N_13832);
or U14863 (N_14863,N_12940,N_12593);
nor U14864 (N_14864,N_12880,N_12717);
xor U14865 (N_14865,N_13316,N_13522);
or U14866 (N_14866,N_12788,N_12939);
nand U14867 (N_14867,N_12456,N_13327);
nor U14868 (N_14868,N_12109,N_13482);
xor U14869 (N_14869,N_13178,N_13910);
nand U14870 (N_14870,N_13836,N_13448);
and U14871 (N_14871,N_13805,N_13523);
nand U14872 (N_14872,N_12069,N_12361);
nor U14873 (N_14873,N_13119,N_12772);
nand U14874 (N_14874,N_12047,N_13889);
and U14875 (N_14875,N_13905,N_13106);
xnor U14876 (N_14876,N_13489,N_13822);
nand U14877 (N_14877,N_12551,N_13230);
nor U14878 (N_14878,N_12359,N_12987);
nand U14879 (N_14879,N_12605,N_12329);
or U14880 (N_14880,N_12276,N_12246);
nand U14881 (N_14881,N_12929,N_13770);
or U14882 (N_14882,N_13696,N_12634);
and U14883 (N_14883,N_12149,N_13884);
and U14884 (N_14884,N_13418,N_12379);
xnor U14885 (N_14885,N_12076,N_13125);
or U14886 (N_14886,N_12208,N_13804);
nor U14887 (N_14887,N_13582,N_13605);
nor U14888 (N_14888,N_13997,N_12488);
nand U14889 (N_14889,N_12200,N_12184);
and U14890 (N_14890,N_12416,N_13047);
or U14891 (N_14891,N_13369,N_13227);
nor U14892 (N_14892,N_13950,N_13253);
nor U14893 (N_14893,N_13801,N_12904);
nand U14894 (N_14894,N_12117,N_12543);
nor U14895 (N_14895,N_12037,N_12096);
nor U14896 (N_14896,N_12183,N_12460);
nor U14897 (N_14897,N_13183,N_12201);
nor U14898 (N_14898,N_13710,N_12595);
or U14899 (N_14899,N_12657,N_12113);
nand U14900 (N_14900,N_12730,N_12842);
xnor U14901 (N_14901,N_13115,N_12335);
and U14902 (N_14902,N_13146,N_12080);
and U14903 (N_14903,N_12514,N_12319);
or U14904 (N_14904,N_13554,N_13315);
nand U14905 (N_14905,N_13456,N_12212);
and U14906 (N_14906,N_13689,N_12167);
nand U14907 (N_14907,N_13019,N_13455);
nand U14908 (N_14908,N_13752,N_12467);
nor U14909 (N_14909,N_12793,N_13965);
nand U14910 (N_14910,N_13140,N_13525);
and U14911 (N_14911,N_13381,N_12151);
nor U14912 (N_14912,N_12812,N_13830);
and U14913 (N_14913,N_13403,N_12620);
nand U14914 (N_14914,N_13674,N_13698);
and U14915 (N_14915,N_12946,N_13185);
or U14916 (N_14916,N_12865,N_12033);
nand U14917 (N_14917,N_12909,N_12794);
nand U14918 (N_14918,N_12672,N_13646);
nor U14919 (N_14919,N_12126,N_13958);
nand U14920 (N_14920,N_12538,N_13058);
nand U14921 (N_14921,N_13542,N_12161);
and U14922 (N_14922,N_13637,N_13753);
or U14923 (N_14923,N_12534,N_13189);
and U14924 (N_14924,N_12695,N_13599);
or U14925 (N_14925,N_12818,N_13088);
xnor U14926 (N_14926,N_12203,N_12017);
or U14927 (N_14927,N_12613,N_12462);
or U14928 (N_14928,N_12326,N_13287);
nand U14929 (N_14929,N_12786,N_13382);
nand U14930 (N_14930,N_12255,N_12955);
and U14931 (N_14931,N_13392,N_12023);
or U14932 (N_14932,N_12933,N_12040);
and U14933 (N_14933,N_12845,N_13984);
or U14934 (N_14934,N_12849,N_13567);
and U14935 (N_14935,N_12681,N_12081);
nor U14936 (N_14936,N_12535,N_12443);
nand U14937 (N_14937,N_12694,N_13309);
or U14938 (N_14938,N_12546,N_13673);
or U14939 (N_14939,N_12840,N_12195);
nor U14940 (N_14940,N_13638,N_13276);
and U14941 (N_14941,N_13265,N_12655);
and U14942 (N_14942,N_13662,N_12547);
xnor U14943 (N_14943,N_12873,N_13039);
and U14944 (N_14944,N_12572,N_13598);
xnor U14945 (N_14945,N_13428,N_12464);
xnor U14946 (N_14946,N_12732,N_12850);
and U14947 (N_14947,N_13918,N_12331);
nor U14948 (N_14948,N_13416,N_12752);
or U14949 (N_14949,N_12447,N_13548);
and U14950 (N_14950,N_12285,N_13857);
xor U14951 (N_14951,N_12408,N_12549);
nor U14952 (N_14952,N_12043,N_13942);
nand U14953 (N_14953,N_12296,N_13154);
nand U14954 (N_14954,N_13162,N_13515);
or U14955 (N_14955,N_12992,N_12174);
nor U14956 (N_14956,N_12086,N_12754);
xor U14957 (N_14957,N_13373,N_13799);
and U14958 (N_14958,N_13099,N_12858);
or U14959 (N_14959,N_12351,N_12232);
nand U14960 (N_14960,N_12163,N_12674);
nand U14961 (N_14961,N_13285,N_13406);
or U14962 (N_14962,N_13974,N_13209);
nand U14963 (N_14963,N_13365,N_13866);
nand U14964 (N_14964,N_12198,N_12632);
nor U14965 (N_14965,N_12503,N_12115);
or U14966 (N_14966,N_12426,N_12957);
and U14967 (N_14967,N_12414,N_12050);
and U14968 (N_14968,N_12855,N_12899);
nand U14969 (N_14969,N_12369,N_12094);
or U14970 (N_14970,N_12038,N_12469);
or U14971 (N_14971,N_13446,N_13962);
or U14972 (N_14972,N_13704,N_13906);
and U14973 (N_14973,N_13749,N_13043);
nor U14974 (N_14974,N_13979,N_12486);
xnor U14975 (N_14975,N_13000,N_13103);
nand U14976 (N_14976,N_13420,N_13298);
or U14977 (N_14977,N_13641,N_12286);
nand U14978 (N_14978,N_12284,N_13171);
nand U14979 (N_14979,N_13417,N_13955);
or U14980 (N_14980,N_13999,N_12343);
nand U14981 (N_14981,N_13379,N_13829);
or U14982 (N_14982,N_12614,N_12959);
nand U14983 (N_14983,N_13005,N_12791);
nand U14984 (N_14984,N_12442,N_13506);
nand U14985 (N_14985,N_13015,N_12112);
nor U14986 (N_14986,N_12829,N_12796);
nand U14987 (N_14987,N_12399,N_13915);
nor U14988 (N_14988,N_12738,N_13399);
or U14989 (N_14989,N_13046,N_12470);
and U14990 (N_14990,N_12961,N_13967);
or U14991 (N_14991,N_12061,N_13050);
nand U14992 (N_14992,N_13007,N_13295);
nor U14993 (N_14993,N_12492,N_13681);
nor U14994 (N_14994,N_13533,N_13862);
or U14995 (N_14995,N_13117,N_12886);
and U14996 (N_14996,N_12641,N_12307);
or U14997 (N_14997,N_13228,N_13835);
or U14998 (N_14998,N_12966,N_13092);
or U14999 (N_14999,N_12474,N_12097);
or U15000 (N_15000,N_13085,N_12024);
nor U15001 (N_15001,N_12357,N_13341);
nand U15002 (N_15002,N_12315,N_13277);
nand U15003 (N_15003,N_13444,N_12138);
and U15004 (N_15004,N_12044,N_13961);
or U15005 (N_15005,N_12323,N_13126);
xnor U15006 (N_15006,N_13891,N_13307);
or U15007 (N_15007,N_13030,N_13629);
nand U15008 (N_15008,N_13466,N_13707);
nand U15009 (N_15009,N_13594,N_13368);
xnor U15010 (N_15010,N_13428,N_12443);
nor U15011 (N_15011,N_13640,N_12192);
or U15012 (N_15012,N_12205,N_12315);
nand U15013 (N_15013,N_13091,N_13490);
nor U15014 (N_15014,N_12489,N_13544);
and U15015 (N_15015,N_13951,N_12524);
nand U15016 (N_15016,N_13298,N_12461);
or U15017 (N_15017,N_13530,N_13132);
or U15018 (N_15018,N_13353,N_12662);
nand U15019 (N_15019,N_13616,N_12728);
and U15020 (N_15020,N_12723,N_12134);
xor U15021 (N_15021,N_12002,N_13288);
nor U15022 (N_15022,N_13008,N_13665);
or U15023 (N_15023,N_12928,N_13876);
nor U15024 (N_15024,N_13595,N_13569);
nand U15025 (N_15025,N_12373,N_12231);
nand U15026 (N_15026,N_12011,N_13505);
or U15027 (N_15027,N_13827,N_12516);
or U15028 (N_15028,N_13576,N_12311);
and U15029 (N_15029,N_13447,N_12447);
nor U15030 (N_15030,N_13323,N_12449);
and U15031 (N_15031,N_13112,N_12082);
and U15032 (N_15032,N_13583,N_13746);
nor U15033 (N_15033,N_12202,N_12594);
and U15034 (N_15034,N_12917,N_13190);
or U15035 (N_15035,N_13607,N_12155);
nor U15036 (N_15036,N_12733,N_12260);
and U15037 (N_15037,N_12862,N_13021);
xnor U15038 (N_15038,N_13585,N_13197);
and U15039 (N_15039,N_12106,N_13733);
or U15040 (N_15040,N_13350,N_12752);
xnor U15041 (N_15041,N_13409,N_13017);
nand U15042 (N_15042,N_12297,N_13616);
and U15043 (N_15043,N_13520,N_13124);
or U15044 (N_15044,N_13907,N_13506);
nor U15045 (N_15045,N_13449,N_13393);
nand U15046 (N_15046,N_13926,N_13345);
or U15047 (N_15047,N_12076,N_13679);
nand U15048 (N_15048,N_13875,N_12135);
nand U15049 (N_15049,N_12882,N_12953);
nor U15050 (N_15050,N_13292,N_13588);
nor U15051 (N_15051,N_13281,N_12509);
nand U15052 (N_15052,N_13895,N_12313);
and U15053 (N_15053,N_13443,N_13525);
or U15054 (N_15054,N_12503,N_13610);
nor U15055 (N_15055,N_13049,N_13133);
nor U15056 (N_15056,N_12034,N_12546);
nor U15057 (N_15057,N_12160,N_12614);
xnor U15058 (N_15058,N_12887,N_12191);
nor U15059 (N_15059,N_12885,N_13017);
and U15060 (N_15060,N_12535,N_12189);
and U15061 (N_15061,N_13067,N_12746);
and U15062 (N_15062,N_12668,N_13793);
and U15063 (N_15063,N_13672,N_13352);
and U15064 (N_15064,N_12624,N_12208);
and U15065 (N_15065,N_13499,N_12752);
xnor U15066 (N_15066,N_13758,N_12326);
or U15067 (N_15067,N_13845,N_13836);
nor U15068 (N_15068,N_13098,N_13579);
nor U15069 (N_15069,N_13643,N_13073);
nand U15070 (N_15070,N_12503,N_12654);
and U15071 (N_15071,N_13245,N_13009);
and U15072 (N_15072,N_12114,N_12432);
and U15073 (N_15073,N_13770,N_12928);
nor U15074 (N_15074,N_13117,N_12468);
xnor U15075 (N_15075,N_13491,N_13381);
nand U15076 (N_15076,N_12766,N_13001);
and U15077 (N_15077,N_12022,N_12309);
or U15078 (N_15078,N_12944,N_13219);
and U15079 (N_15079,N_13384,N_12963);
and U15080 (N_15080,N_13094,N_13735);
nand U15081 (N_15081,N_12343,N_13308);
nor U15082 (N_15082,N_12361,N_12425);
and U15083 (N_15083,N_12650,N_12164);
and U15084 (N_15084,N_12812,N_12428);
and U15085 (N_15085,N_12994,N_13143);
and U15086 (N_15086,N_13435,N_13867);
nor U15087 (N_15087,N_12964,N_12286);
nor U15088 (N_15088,N_13002,N_13469);
or U15089 (N_15089,N_13373,N_12375);
and U15090 (N_15090,N_13185,N_12591);
xor U15091 (N_15091,N_12692,N_12444);
xor U15092 (N_15092,N_12239,N_13575);
nor U15093 (N_15093,N_12454,N_12058);
nand U15094 (N_15094,N_13859,N_12772);
nor U15095 (N_15095,N_13044,N_12201);
nor U15096 (N_15096,N_13844,N_13104);
nand U15097 (N_15097,N_13485,N_12721);
and U15098 (N_15098,N_12879,N_13222);
or U15099 (N_15099,N_13275,N_13957);
xnor U15100 (N_15100,N_13577,N_13563);
or U15101 (N_15101,N_12415,N_13724);
nor U15102 (N_15102,N_13914,N_12718);
and U15103 (N_15103,N_12909,N_12024);
or U15104 (N_15104,N_12117,N_12317);
nand U15105 (N_15105,N_12200,N_13313);
xor U15106 (N_15106,N_12983,N_13929);
nor U15107 (N_15107,N_13380,N_13348);
nand U15108 (N_15108,N_12494,N_13690);
nand U15109 (N_15109,N_13767,N_13732);
or U15110 (N_15110,N_13615,N_13468);
xor U15111 (N_15111,N_13005,N_12733);
nand U15112 (N_15112,N_13465,N_13991);
or U15113 (N_15113,N_12427,N_13764);
and U15114 (N_15114,N_13342,N_13327);
or U15115 (N_15115,N_12593,N_12292);
or U15116 (N_15116,N_13722,N_12654);
or U15117 (N_15117,N_13451,N_13596);
nor U15118 (N_15118,N_12115,N_13586);
nor U15119 (N_15119,N_13649,N_12273);
nor U15120 (N_15120,N_12238,N_13886);
and U15121 (N_15121,N_12297,N_12147);
nand U15122 (N_15122,N_13508,N_12868);
nor U15123 (N_15123,N_12839,N_13486);
and U15124 (N_15124,N_13416,N_13410);
nand U15125 (N_15125,N_12565,N_12746);
or U15126 (N_15126,N_12752,N_12793);
or U15127 (N_15127,N_13885,N_12651);
and U15128 (N_15128,N_13359,N_13463);
xor U15129 (N_15129,N_12760,N_13352);
nor U15130 (N_15130,N_13402,N_12638);
or U15131 (N_15131,N_12045,N_12864);
nand U15132 (N_15132,N_13064,N_13532);
and U15133 (N_15133,N_12489,N_12351);
nand U15134 (N_15134,N_13664,N_13694);
and U15135 (N_15135,N_12696,N_12772);
or U15136 (N_15136,N_13428,N_13242);
and U15137 (N_15137,N_13358,N_13845);
nor U15138 (N_15138,N_13207,N_13735);
and U15139 (N_15139,N_13174,N_13476);
xor U15140 (N_15140,N_13068,N_12853);
and U15141 (N_15141,N_13901,N_13714);
and U15142 (N_15142,N_13082,N_12692);
nor U15143 (N_15143,N_12791,N_13453);
xor U15144 (N_15144,N_12936,N_13883);
nor U15145 (N_15145,N_12866,N_12355);
and U15146 (N_15146,N_12850,N_12364);
nand U15147 (N_15147,N_13569,N_13629);
and U15148 (N_15148,N_13666,N_12877);
or U15149 (N_15149,N_12789,N_12199);
nor U15150 (N_15150,N_13321,N_13191);
nor U15151 (N_15151,N_13614,N_12124);
nor U15152 (N_15152,N_12540,N_13309);
nor U15153 (N_15153,N_13271,N_12206);
or U15154 (N_15154,N_13039,N_13706);
or U15155 (N_15155,N_12163,N_12320);
xor U15156 (N_15156,N_12167,N_13124);
xor U15157 (N_15157,N_12339,N_12321);
or U15158 (N_15158,N_12041,N_13772);
nor U15159 (N_15159,N_13511,N_12244);
xor U15160 (N_15160,N_12268,N_12829);
nor U15161 (N_15161,N_12888,N_13608);
xor U15162 (N_15162,N_12304,N_12657);
nor U15163 (N_15163,N_12647,N_13363);
nor U15164 (N_15164,N_13261,N_12170);
and U15165 (N_15165,N_12440,N_13825);
nand U15166 (N_15166,N_12312,N_12075);
nand U15167 (N_15167,N_12949,N_13995);
nor U15168 (N_15168,N_12989,N_13180);
nand U15169 (N_15169,N_13015,N_12341);
nand U15170 (N_15170,N_13451,N_13375);
nor U15171 (N_15171,N_13245,N_12280);
nor U15172 (N_15172,N_13603,N_12636);
xor U15173 (N_15173,N_12829,N_12982);
and U15174 (N_15174,N_13702,N_13488);
or U15175 (N_15175,N_13107,N_12028);
nand U15176 (N_15176,N_13313,N_13490);
nor U15177 (N_15177,N_12618,N_13121);
nand U15178 (N_15178,N_13673,N_13943);
nand U15179 (N_15179,N_12666,N_12234);
and U15180 (N_15180,N_12685,N_13049);
nor U15181 (N_15181,N_13505,N_12935);
or U15182 (N_15182,N_13788,N_12608);
nor U15183 (N_15183,N_13612,N_12086);
nand U15184 (N_15184,N_12340,N_13137);
nor U15185 (N_15185,N_12470,N_13004);
or U15186 (N_15186,N_13652,N_12119);
or U15187 (N_15187,N_12991,N_13847);
nor U15188 (N_15188,N_12784,N_13995);
nor U15189 (N_15189,N_13777,N_12790);
and U15190 (N_15190,N_13648,N_13186);
and U15191 (N_15191,N_13627,N_12088);
and U15192 (N_15192,N_12120,N_12834);
nor U15193 (N_15193,N_13468,N_13379);
nor U15194 (N_15194,N_13140,N_13125);
or U15195 (N_15195,N_13969,N_12048);
xor U15196 (N_15196,N_12796,N_13292);
nand U15197 (N_15197,N_12283,N_13490);
nor U15198 (N_15198,N_13860,N_13953);
nand U15199 (N_15199,N_12608,N_13387);
xor U15200 (N_15200,N_13464,N_13411);
or U15201 (N_15201,N_13505,N_13528);
nand U15202 (N_15202,N_13612,N_13011);
or U15203 (N_15203,N_12885,N_12130);
xor U15204 (N_15204,N_12896,N_13017);
nand U15205 (N_15205,N_12279,N_13550);
nand U15206 (N_15206,N_12080,N_12649);
nor U15207 (N_15207,N_13631,N_13351);
or U15208 (N_15208,N_13358,N_12381);
nand U15209 (N_15209,N_12014,N_13431);
or U15210 (N_15210,N_13830,N_12607);
nor U15211 (N_15211,N_13545,N_12705);
nor U15212 (N_15212,N_12196,N_13758);
and U15213 (N_15213,N_12032,N_12365);
and U15214 (N_15214,N_12072,N_13363);
nand U15215 (N_15215,N_12217,N_13897);
and U15216 (N_15216,N_13802,N_12042);
and U15217 (N_15217,N_12470,N_13208);
or U15218 (N_15218,N_13837,N_13261);
and U15219 (N_15219,N_12592,N_12086);
nand U15220 (N_15220,N_13379,N_13736);
and U15221 (N_15221,N_12313,N_12655);
xnor U15222 (N_15222,N_13144,N_13582);
or U15223 (N_15223,N_13736,N_12740);
nor U15224 (N_15224,N_13084,N_13810);
or U15225 (N_15225,N_13659,N_13412);
or U15226 (N_15226,N_13801,N_13495);
or U15227 (N_15227,N_13907,N_13981);
and U15228 (N_15228,N_13048,N_13438);
nor U15229 (N_15229,N_13868,N_12279);
nor U15230 (N_15230,N_13022,N_13005);
and U15231 (N_15231,N_13416,N_13993);
nor U15232 (N_15232,N_12348,N_12437);
nor U15233 (N_15233,N_13790,N_12637);
nor U15234 (N_15234,N_13284,N_13858);
nand U15235 (N_15235,N_13362,N_12604);
or U15236 (N_15236,N_12722,N_12688);
and U15237 (N_15237,N_13514,N_12906);
nor U15238 (N_15238,N_13854,N_12335);
nand U15239 (N_15239,N_12204,N_13774);
or U15240 (N_15240,N_13722,N_12364);
and U15241 (N_15241,N_13644,N_13638);
xor U15242 (N_15242,N_12411,N_12398);
nor U15243 (N_15243,N_13645,N_13172);
nor U15244 (N_15244,N_13021,N_12941);
nor U15245 (N_15245,N_13570,N_13604);
nor U15246 (N_15246,N_12066,N_13421);
nand U15247 (N_15247,N_12920,N_12551);
nor U15248 (N_15248,N_13168,N_13220);
nand U15249 (N_15249,N_13772,N_12691);
nor U15250 (N_15250,N_13111,N_13584);
nor U15251 (N_15251,N_12523,N_12542);
and U15252 (N_15252,N_13554,N_12468);
or U15253 (N_15253,N_13511,N_13128);
nand U15254 (N_15254,N_12114,N_13948);
nand U15255 (N_15255,N_12643,N_13431);
nand U15256 (N_15256,N_13819,N_12602);
and U15257 (N_15257,N_13397,N_12836);
nand U15258 (N_15258,N_12310,N_13025);
nor U15259 (N_15259,N_13151,N_13216);
nor U15260 (N_15260,N_12953,N_12344);
nand U15261 (N_15261,N_13215,N_12493);
nand U15262 (N_15262,N_12921,N_13957);
nor U15263 (N_15263,N_12439,N_12929);
nor U15264 (N_15264,N_13886,N_12182);
nor U15265 (N_15265,N_12758,N_13512);
xnor U15266 (N_15266,N_12296,N_13653);
nand U15267 (N_15267,N_12087,N_13555);
and U15268 (N_15268,N_12993,N_13790);
nor U15269 (N_15269,N_13401,N_12679);
nand U15270 (N_15270,N_12171,N_13131);
or U15271 (N_15271,N_12639,N_13210);
nand U15272 (N_15272,N_13854,N_13175);
nand U15273 (N_15273,N_13029,N_13376);
or U15274 (N_15274,N_12802,N_13172);
xnor U15275 (N_15275,N_13756,N_13449);
nand U15276 (N_15276,N_12333,N_13464);
nand U15277 (N_15277,N_12747,N_12905);
nor U15278 (N_15278,N_13915,N_12218);
nor U15279 (N_15279,N_13387,N_13373);
xnor U15280 (N_15280,N_12359,N_12037);
nand U15281 (N_15281,N_12994,N_13288);
xor U15282 (N_15282,N_13028,N_13157);
nand U15283 (N_15283,N_13570,N_12641);
nand U15284 (N_15284,N_13674,N_13908);
xor U15285 (N_15285,N_12704,N_13727);
nand U15286 (N_15286,N_12296,N_12010);
nand U15287 (N_15287,N_13257,N_12907);
and U15288 (N_15288,N_12835,N_12998);
or U15289 (N_15289,N_13431,N_13722);
nor U15290 (N_15290,N_12259,N_12975);
nor U15291 (N_15291,N_13406,N_12891);
and U15292 (N_15292,N_12291,N_12841);
or U15293 (N_15293,N_12076,N_12070);
or U15294 (N_15294,N_12847,N_13382);
or U15295 (N_15295,N_13137,N_13930);
nor U15296 (N_15296,N_13843,N_12681);
nand U15297 (N_15297,N_13673,N_13068);
or U15298 (N_15298,N_13670,N_13037);
nand U15299 (N_15299,N_12704,N_12844);
or U15300 (N_15300,N_13281,N_12389);
nand U15301 (N_15301,N_13967,N_12679);
nor U15302 (N_15302,N_12023,N_12265);
or U15303 (N_15303,N_12813,N_12645);
and U15304 (N_15304,N_12291,N_13013);
and U15305 (N_15305,N_12383,N_13058);
and U15306 (N_15306,N_12816,N_12274);
or U15307 (N_15307,N_13600,N_12807);
or U15308 (N_15308,N_13000,N_12451);
xnor U15309 (N_15309,N_12242,N_13024);
nand U15310 (N_15310,N_12353,N_12116);
xor U15311 (N_15311,N_13275,N_12868);
nand U15312 (N_15312,N_12697,N_12545);
nor U15313 (N_15313,N_12656,N_12108);
and U15314 (N_15314,N_12210,N_13230);
and U15315 (N_15315,N_13246,N_13457);
nand U15316 (N_15316,N_12926,N_12173);
nor U15317 (N_15317,N_13046,N_13667);
or U15318 (N_15318,N_12435,N_12140);
or U15319 (N_15319,N_13815,N_12660);
and U15320 (N_15320,N_13456,N_12432);
nand U15321 (N_15321,N_12874,N_12153);
xnor U15322 (N_15322,N_12046,N_12228);
or U15323 (N_15323,N_12696,N_13574);
nor U15324 (N_15324,N_12006,N_13514);
nor U15325 (N_15325,N_13019,N_13559);
or U15326 (N_15326,N_13002,N_13450);
nand U15327 (N_15327,N_13865,N_13555);
or U15328 (N_15328,N_13620,N_13383);
nand U15329 (N_15329,N_12796,N_13903);
nor U15330 (N_15330,N_13672,N_12273);
nor U15331 (N_15331,N_13253,N_13446);
and U15332 (N_15332,N_13324,N_12769);
or U15333 (N_15333,N_13593,N_13408);
or U15334 (N_15334,N_12903,N_13982);
and U15335 (N_15335,N_12404,N_13262);
xnor U15336 (N_15336,N_13780,N_13721);
or U15337 (N_15337,N_13592,N_12110);
xor U15338 (N_15338,N_12082,N_12389);
and U15339 (N_15339,N_12069,N_13448);
and U15340 (N_15340,N_12500,N_12986);
nand U15341 (N_15341,N_13055,N_13016);
or U15342 (N_15342,N_12045,N_12028);
nor U15343 (N_15343,N_13086,N_13233);
or U15344 (N_15344,N_12474,N_12099);
nand U15345 (N_15345,N_13298,N_12213);
nand U15346 (N_15346,N_13597,N_13228);
xnor U15347 (N_15347,N_12044,N_13837);
or U15348 (N_15348,N_12570,N_13617);
nand U15349 (N_15349,N_13455,N_12141);
and U15350 (N_15350,N_13072,N_13711);
nand U15351 (N_15351,N_12239,N_12518);
and U15352 (N_15352,N_12413,N_13938);
or U15353 (N_15353,N_13716,N_12001);
and U15354 (N_15354,N_12277,N_12153);
nor U15355 (N_15355,N_12067,N_13602);
nand U15356 (N_15356,N_12218,N_12626);
nand U15357 (N_15357,N_13965,N_12953);
and U15358 (N_15358,N_12105,N_12383);
xor U15359 (N_15359,N_12795,N_12485);
nor U15360 (N_15360,N_13929,N_12961);
or U15361 (N_15361,N_12536,N_12625);
or U15362 (N_15362,N_13112,N_12969);
nor U15363 (N_15363,N_12451,N_12958);
nor U15364 (N_15364,N_13878,N_12046);
xnor U15365 (N_15365,N_12895,N_13140);
nor U15366 (N_15366,N_12513,N_13878);
nand U15367 (N_15367,N_12472,N_12129);
nand U15368 (N_15368,N_12482,N_12440);
and U15369 (N_15369,N_12856,N_12954);
xor U15370 (N_15370,N_13968,N_13360);
nor U15371 (N_15371,N_12312,N_13648);
nor U15372 (N_15372,N_12683,N_12101);
nand U15373 (N_15373,N_12170,N_13118);
or U15374 (N_15374,N_12923,N_12474);
nand U15375 (N_15375,N_13484,N_13261);
xnor U15376 (N_15376,N_12019,N_13460);
nand U15377 (N_15377,N_12914,N_12837);
and U15378 (N_15378,N_13353,N_13482);
or U15379 (N_15379,N_12893,N_12443);
xnor U15380 (N_15380,N_13450,N_12551);
nand U15381 (N_15381,N_13705,N_13623);
xnor U15382 (N_15382,N_12536,N_13816);
and U15383 (N_15383,N_12969,N_13082);
and U15384 (N_15384,N_13068,N_13170);
and U15385 (N_15385,N_12000,N_13967);
or U15386 (N_15386,N_12631,N_12558);
nor U15387 (N_15387,N_12710,N_12718);
nor U15388 (N_15388,N_12446,N_13951);
xnor U15389 (N_15389,N_13234,N_13132);
or U15390 (N_15390,N_13196,N_13160);
nor U15391 (N_15391,N_13803,N_13290);
or U15392 (N_15392,N_13609,N_12458);
and U15393 (N_15393,N_13468,N_12164);
and U15394 (N_15394,N_12625,N_13967);
and U15395 (N_15395,N_13482,N_12566);
or U15396 (N_15396,N_12636,N_13128);
nor U15397 (N_15397,N_13056,N_13281);
nor U15398 (N_15398,N_13203,N_13620);
and U15399 (N_15399,N_13793,N_13245);
nand U15400 (N_15400,N_13582,N_13532);
nor U15401 (N_15401,N_13171,N_13882);
nand U15402 (N_15402,N_13954,N_12465);
xnor U15403 (N_15403,N_12409,N_13638);
xnor U15404 (N_15404,N_13531,N_13956);
and U15405 (N_15405,N_13181,N_13698);
nor U15406 (N_15406,N_12815,N_13009);
and U15407 (N_15407,N_13410,N_12501);
nand U15408 (N_15408,N_13543,N_13667);
nand U15409 (N_15409,N_13552,N_12550);
nor U15410 (N_15410,N_13582,N_13080);
nor U15411 (N_15411,N_13379,N_13289);
nor U15412 (N_15412,N_12252,N_13543);
and U15413 (N_15413,N_13934,N_13828);
and U15414 (N_15414,N_12846,N_13460);
or U15415 (N_15415,N_12079,N_13811);
or U15416 (N_15416,N_12935,N_13666);
xor U15417 (N_15417,N_13319,N_12196);
or U15418 (N_15418,N_13552,N_12609);
and U15419 (N_15419,N_12388,N_13330);
or U15420 (N_15420,N_12433,N_13924);
and U15421 (N_15421,N_13715,N_12451);
or U15422 (N_15422,N_13333,N_13643);
nor U15423 (N_15423,N_12144,N_13925);
nand U15424 (N_15424,N_13785,N_12399);
or U15425 (N_15425,N_13831,N_12579);
or U15426 (N_15426,N_13904,N_13707);
nor U15427 (N_15427,N_13990,N_12346);
and U15428 (N_15428,N_12849,N_12644);
or U15429 (N_15429,N_13912,N_13822);
or U15430 (N_15430,N_13913,N_12741);
or U15431 (N_15431,N_13324,N_12434);
nand U15432 (N_15432,N_12484,N_13152);
nand U15433 (N_15433,N_12847,N_13875);
or U15434 (N_15434,N_12481,N_12742);
xor U15435 (N_15435,N_13214,N_13640);
nor U15436 (N_15436,N_12453,N_13107);
or U15437 (N_15437,N_12376,N_12706);
or U15438 (N_15438,N_13309,N_13722);
nand U15439 (N_15439,N_13103,N_12422);
and U15440 (N_15440,N_12034,N_12296);
and U15441 (N_15441,N_13899,N_12504);
and U15442 (N_15442,N_13348,N_12901);
nor U15443 (N_15443,N_13335,N_12302);
nand U15444 (N_15444,N_12657,N_13089);
nand U15445 (N_15445,N_13208,N_13609);
nand U15446 (N_15446,N_12445,N_13181);
or U15447 (N_15447,N_12779,N_13423);
or U15448 (N_15448,N_12845,N_13079);
nand U15449 (N_15449,N_12080,N_13905);
xnor U15450 (N_15450,N_12265,N_13228);
and U15451 (N_15451,N_12434,N_13930);
and U15452 (N_15452,N_12019,N_13212);
and U15453 (N_15453,N_13711,N_12096);
nand U15454 (N_15454,N_12707,N_13939);
or U15455 (N_15455,N_12675,N_12245);
nor U15456 (N_15456,N_12530,N_13742);
nand U15457 (N_15457,N_12661,N_12339);
nand U15458 (N_15458,N_12462,N_13808);
nor U15459 (N_15459,N_12850,N_13059);
nor U15460 (N_15460,N_13425,N_12951);
and U15461 (N_15461,N_12522,N_12299);
xor U15462 (N_15462,N_12824,N_13616);
nor U15463 (N_15463,N_13498,N_12850);
nand U15464 (N_15464,N_12994,N_13182);
xnor U15465 (N_15465,N_13258,N_13086);
or U15466 (N_15466,N_13119,N_13105);
nor U15467 (N_15467,N_13134,N_12760);
and U15468 (N_15468,N_12677,N_12933);
xor U15469 (N_15469,N_12406,N_12792);
nand U15470 (N_15470,N_12525,N_13841);
nand U15471 (N_15471,N_12939,N_13074);
nand U15472 (N_15472,N_12425,N_12554);
nand U15473 (N_15473,N_12156,N_13466);
or U15474 (N_15474,N_13749,N_12473);
and U15475 (N_15475,N_13487,N_13442);
or U15476 (N_15476,N_13689,N_12615);
or U15477 (N_15477,N_13155,N_12587);
and U15478 (N_15478,N_13062,N_13504);
or U15479 (N_15479,N_13222,N_12047);
and U15480 (N_15480,N_12202,N_12413);
nor U15481 (N_15481,N_13176,N_13212);
nand U15482 (N_15482,N_13021,N_12997);
and U15483 (N_15483,N_12317,N_13168);
nor U15484 (N_15484,N_12354,N_13602);
and U15485 (N_15485,N_13989,N_13506);
nor U15486 (N_15486,N_12268,N_13893);
or U15487 (N_15487,N_12866,N_13456);
nor U15488 (N_15488,N_13334,N_13563);
or U15489 (N_15489,N_13476,N_13224);
or U15490 (N_15490,N_13229,N_13899);
and U15491 (N_15491,N_12063,N_13518);
nand U15492 (N_15492,N_12701,N_12212);
and U15493 (N_15493,N_12852,N_12908);
nor U15494 (N_15494,N_12255,N_13740);
xnor U15495 (N_15495,N_12401,N_12849);
nand U15496 (N_15496,N_13030,N_12732);
nor U15497 (N_15497,N_13514,N_13118);
nand U15498 (N_15498,N_13842,N_12315);
and U15499 (N_15499,N_12557,N_12046);
nor U15500 (N_15500,N_13684,N_13196);
or U15501 (N_15501,N_12023,N_12794);
and U15502 (N_15502,N_13055,N_13922);
nor U15503 (N_15503,N_13377,N_13115);
nand U15504 (N_15504,N_12152,N_13957);
and U15505 (N_15505,N_12701,N_13391);
and U15506 (N_15506,N_13462,N_13373);
nor U15507 (N_15507,N_13634,N_13247);
and U15508 (N_15508,N_13782,N_12456);
or U15509 (N_15509,N_13275,N_13728);
and U15510 (N_15510,N_12402,N_13444);
xor U15511 (N_15511,N_12432,N_13274);
or U15512 (N_15512,N_12924,N_12736);
and U15513 (N_15513,N_13891,N_13711);
xor U15514 (N_15514,N_12000,N_13925);
or U15515 (N_15515,N_12122,N_13865);
nand U15516 (N_15516,N_13797,N_13199);
nand U15517 (N_15517,N_12835,N_13182);
nor U15518 (N_15518,N_13816,N_12876);
nor U15519 (N_15519,N_13949,N_12652);
and U15520 (N_15520,N_13738,N_12535);
nand U15521 (N_15521,N_13157,N_12617);
and U15522 (N_15522,N_13869,N_13510);
or U15523 (N_15523,N_12100,N_12994);
nand U15524 (N_15524,N_13484,N_12706);
or U15525 (N_15525,N_12912,N_13178);
or U15526 (N_15526,N_12644,N_13675);
nor U15527 (N_15527,N_12945,N_13859);
nand U15528 (N_15528,N_12313,N_13883);
and U15529 (N_15529,N_12962,N_12088);
nor U15530 (N_15530,N_12954,N_13586);
nor U15531 (N_15531,N_13094,N_13653);
xnor U15532 (N_15532,N_12749,N_12240);
nand U15533 (N_15533,N_12536,N_12296);
xor U15534 (N_15534,N_13602,N_12528);
nor U15535 (N_15535,N_13455,N_12833);
nand U15536 (N_15536,N_13172,N_12605);
nand U15537 (N_15537,N_12696,N_12839);
nand U15538 (N_15538,N_12844,N_13324);
and U15539 (N_15539,N_12724,N_12062);
or U15540 (N_15540,N_13010,N_12806);
xnor U15541 (N_15541,N_13369,N_12053);
nand U15542 (N_15542,N_12745,N_12725);
or U15543 (N_15543,N_12741,N_12424);
nand U15544 (N_15544,N_13855,N_13969);
nor U15545 (N_15545,N_13852,N_13427);
xnor U15546 (N_15546,N_12503,N_13700);
nand U15547 (N_15547,N_13172,N_13379);
xnor U15548 (N_15548,N_13164,N_12346);
nand U15549 (N_15549,N_13562,N_12967);
nor U15550 (N_15550,N_13841,N_12631);
xor U15551 (N_15551,N_12902,N_13211);
nand U15552 (N_15552,N_13659,N_12284);
and U15553 (N_15553,N_13984,N_13105);
and U15554 (N_15554,N_12562,N_13397);
nor U15555 (N_15555,N_12197,N_13158);
nor U15556 (N_15556,N_12107,N_12230);
nand U15557 (N_15557,N_13358,N_12051);
and U15558 (N_15558,N_12850,N_13072);
nor U15559 (N_15559,N_13882,N_13340);
nor U15560 (N_15560,N_12943,N_12440);
nand U15561 (N_15561,N_12771,N_12496);
or U15562 (N_15562,N_13647,N_12886);
nor U15563 (N_15563,N_12471,N_13049);
or U15564 (N_15564,N_13757,N_13882);
nor U15565 (N_15565,N_12905,N_12899);
nand U15566 (N_15566,N_12660,N_12779);
nor U15567 (N_15567,N_13545,N_12584);
nor U15568 (N_15568,N_13705,N_12439);
and U15569 (N_15569,N_12213,N_13784);
nand U15570 (N_15570,N_12886,N_13008);
and U15571 (N_15571,N_13935,N_13907);
nand U15572 (N_15572,N_13014,N_12125);
nor U15573 (N_15573,N_13113,N_13825);
nor U15574 (N_15574,N_12912,N_13165);
and U15575 (N_15575,N_13182,N_12657);
or U15576 (N_15576,N_13015,N_13149);
nand U15577 (N_15577,N_12441,N_13992);
nor U15578 (N_15578,N_12975,N_13673);
and U15579 (N_15579,N_13227,N_12738);
nand U15580 (N_15580,N_12867,N_12819);
and U15581 (N_15581,N_13521,N_12063);
and U15582 (N_15582,N_12299,N_12553);
or U15583 (N_15583,N_13239,N_12939);
nand U15584 (N_15584,N_12622,N_13019);
nor U15585 (N_15585,N_13605,N_13192);
and U15586 (N_15586,N_12043,N_12473);
and U15587 (N_15587,N_12435,N_12887);
and U15588 (N_15588,N_12225,N_13809);
or U15589 (N_15589,N_12624,N_13014);
nand U15590 (N_15590,N_13352,N_12619);
and U15591 (N_15591,N_13471,N_12261);
nand U15592 (N_15592,N_12088,N_13315);
and U15593 (N_15593,N_12853,N_13527);
nor U15594 (N_15594,N_13456,N_12001);
and U15595 (N_15595,N_13490,N_13426);
nand U15596 (N_15596,N_13899,N_13464);
nor U15597 (N_15597,N_12497,N_12198);
nand U15598 (N_15598,N_12218,N_13818);
or U15599 (N_15599,N_12825,N_13832);
or U15600 (N_15600,N_12577,N_12055);
or U15601 (N_15601,N_12577,N_13318);
and U15602 (N_15602,N_13486,N_12306);
nand U15603 (N_15603,N_12026,N_13335);
nor U15604 (N_15604,N_12799,N_13530);
or U15605 (N_15605,N_13261,N_12903);
or U15606 (N_15606,N_13679,N_13984);
nor U15607 (N_15607,N_13407,N_13914);
nand U15608 (N_15608,N_13785,N_13151);
nand U15609 (N_15609,N_12496,N_13857);
nor U15610 (N_15610,N_13541,N_12763);
or U15611 (N_15611,N_12572,N_13739);
xnor U15612 (N_15612,N_13290,N_12479);
or U15613 (N_15613,N_13800,N_12013);
or U15614 (N_15614,N_13506,N_13064);
and U15615 (N_15615,N_12783,N_12547);
nor U15616 (N_15616,N_13818,N_12860);
and U15617 (N_15617,N_12140,N_12132);
and U15618 (N_15618,N_13798,N_13694);
nor U15619 (N_15619,N_12045,N_13936);
xor U15620 (N_15620,N_12692,N_13895);
and U15621 (N_15621,N_13947,N_13401);
nor U15622 (N_15622,N_12655,N_13012);
nor U15623 (N_15623,N_13067,N_12898);
nor U15624 (N_15624,N_12285,N_13892);
nor U15625 (N_15625,N_12659,N_12371);
nand U15626 (N_15626,N_13586,N_12097);
and U15627 (N_15627,N_12818,N_12244);
or U15628 (N_15628,N_13809,N_13993);
nor U15629 (N_15629,N_13272,N_12523);
nand U15630 (N_15630,N_12220,N_12386);
xnor U15631 (N_15631,N_13511,N_13075);
nand U15632 (N_15632,N_13596,N_12561);
and U15633 (N_15633,N_13490,N_13875);
and U15634 (N_15634,N_12484,N_13715);
xnor U15635 (N_15635,N_13722,N_13619);
nand U15636 (N_15636,N_13806,N_13858);
nand U15637 (N_15637,N_13934,N_13712);
xor U15638 (N_15638,N_12374,N_13601);
or U15639 (N_15639,N_12205,N_13113);
nand U15640 (N_15640,N_13358,N_12751);
nand U15641 (N_15641,N_12871,N_12986);
nor U15642 (N_15642,N_13102,N_13976);
nor U15643 (N_15643,N_12456,N_12861);
nor U15644 (N_15644,N_12184,N_13710);
or U15645 (N_15645,N_13113,N_12779);
or U15646 (N_15646,N_13487,N_12542);
nor U15647 (N_15647,N_12135,N_12878);
nand U15648 (N_15648,N_13776,N_12990);
or U15649 (N_15649,N_13401,N_12862);
and U15650 (N_15650,N_13919,N_12007);
or U15651 (N_15651,N_12477,N_12593);
nand U15652 (N_15652,N_13467,N_12484);
nand U15653 (N_15653,N_13461,N_12501);
or U15654 (N_15654,N_13800,N_13368);
or U15655 (N_15655,N_13957,N_13109);
and U15656 (N_15656,N_13668,N_12777);
and U15657 (N_15657,N_12978,N_12402);
nor U15658 (N_15658,N_12677,N_13990);
and U15659 (N_15659,N_13885,N_13993);
and U15660 (N_15660,N_12837,N_12823);
and U15661 (N_15661,N_12194,N_13500);
nand U15662 (N_15662,N_13538,N_12355);
nor U15663 (N_15663,N_13043,N_13860);
and U15664 (N_15664,N_13968,N_12001);
nand U15665 (N_15665,N_12469,N_13163);
nand U15666 (N_15666,N_13940,N_12257);
nor U15667 (N_15667,N_12588,N_12500);
nand U15668 (N_15668,N_12756,N_13341);
xnor U15669 (N_15669,N_13688,N_12426);
nor U15670 (N_15670,N_12497,N_12735);
nand U15671 (N_15671,N_12773,N_13356);
nor U15672 (N_15672,N_13890,N_13630);
xor U15673 (N_15673,N_13757,N_12918);
nor U15674 (N_15674,N_13833,N_13262);
xnor U15675 (N_15675,N_12551,N_12408);
and U15676 (N_15676,N_12874,N_12010);
nand U15677 (N_15677,N_13845,N_13510);
nor U15678 (N_15678,N_13171,N_12928);
and U15679 (N_15679,N_13225,N_12609);
and U15680 (N_15680,N_12528,N_12022);
or U15681 (N_15681,N_12686,N_12134);
or U15682 (N_15682,N_12404,N_12003);
nor U15683 (N_15683,N_13247,N_13322);
nor U15684 (N_15684,N_13872,N_13284);
nand U15685 (N_15685,N_13490,N_12962);
or U15686 (N_15686,N_12249,N_13515);
and U15687 (N_15687,N_13773,N_13964);
nand U15688 (N_15688,N_13379,N_13613);
xor U15689 (N_15689,N_12064,N_12638);
nor U15690 (N_15690,N_12600,N_13260);
or U15691 (N_15691,N_12766,N_13891);
and U15692 (N_15692,N_12813,N_12100);
xor U15693 (N_15693,N_12148,N_13033);
xnor U15694 (N_15694,N_12928,N_12965);
or U15695 (N_15695,N_13968,N_12391);
or U15696 (N_15696,N_12588,N_13074);
nand U15697 (N_15697,N_12474,N_13024);
nor U15698 (N_15698,N_13232,N_12643);
nand U15699 (N_15699,N_13972,N_12694);
and U15700 (N_15700,N_13089,N_12882);
nor U15701 (N_15701,N_12077,N_12599);
nor U15702 (N_15702,N_12715,N_12283);
and U15703 (N_15703,N_12907,N_13534);
nor U15704 (N_15704,N_13390,N_12928);
nand U15705 (N_15705,N_12914,N_12867);
or U15706 (N_15706,N_12501,N_13445);
nand U15707 (N_15707,N_13081,N_13391);
or U15708 (N_15708,N_12736,N_13032);
or U15709 (N_15709,N_13277,N_13777);
nand U15710 (N_15710,N_12076,N_12490);
and U15711 (N_15711,N_12918,N_13302);
nor U15712 (N_15712,N_12574,N_12825);
nand U15713 (N_15713,N_13374,N_12815);
nand U15714 (N_15714,N_13020,N_13016);
xnor U15715 (N_15715,N_12834,N_12873);
nor U15716 (N_15716,N_13342,N_12348);
and U15717 (N_15717,N_12599,N_12450);
nor U15718 (N_15718,N_12271,N_13532);
and U15719 (N_15719,N_12004,N_13733);
or U15720 (N_15720,N_12917,N_13808);
nand U15721 (N_15721,N_12719,N_13378);
nor U15722 (N_15722,N_12938,N_12478);
and U15723 (N_15723,N_12815,N_12681);
and U15724 (N_15724,N_12691,N_12360);
nor U15725 (N_15725,N_12868,N_12857);
or U15726 (N_15726,N_13382,N_13320);
xnor U15727 (N_15727,N_13768,N_12722);
and U15728 (N_15728,N_12913,N_13967);
and U15729 (N_15729,N_13564,N_12781);
and U15730 (N_15730,N_13113,N_12466);
nor U15731 (N_15731,N_13763,N_13921);
xor U15732 (N_15732,N_13410,N_12826);
and U15733 (N_15733,N_12125,N_13681);
xnor U15734 (N_15734,N_12653,N_13611);
nand U15735 (N_15735,N_12497,N_12628);
nor U15736 (N_15736,N_13716,N_13582);
and U15737 (N_15737,N_12072,N_13291);
or U15738 (N_15738,N_13101,N_12167);
nand U15739 (N_15739,N_13106,N_12559);
xnor U15740 (N_15740,N_12548,N_12881);
xor U15741 (N_15741,N_13315,N_12925);
xor U15742 (N_15742,N_13213,N_12039);
and U15743 (N_15743,N_13953,N_13402);
nor U15744 (N_15744,N_12412,N_13525);
nor U15745 (N_15745,N_12248,N_13412);
and U15746 (N_15746,N_13862,N_13114);
nor U15747 (N_15747,N_12197,N_13374);
nand U15748 (N_15748,N_12750,N_12441);
and U15749 (N_15749,N_12874,N_12435);
or U15750 (N_15750,N_13556,N_13397);
nor U15751 (N_15751,N_13143,N_13095);
xor U15752 (N_15752,N_12932,N_12101);
or U15753 (N_15753,N_12383,N_12948);
nor U15754 (N_15754,N_12659,N_13350);
xnor U15755 (N_15755,N_12346,N_13791);
or U15756 (N_15756,N_12840,N_12206);
nand U15757 (N_15757,N_13705,N_12559);
and U15758 (N_15758,N_12853,N_12592);
nand U15759 (N_15759,N_13099,N_12727);
nand U15760 (N_15760,N_13442,N_13307);
xnor U15761 (N_15761,N_12195,N_13995);
nand U15762 (N_15762,N_12626,N_13221);
or U15763 (N_15763,N_12580,N_12662);
or U15764 (N_15764,N_13702,N_12726);
nand U15765 (N_15765,N_13790,N_12398);
nand U15766 (N_15766,N_13064,N_13337);
and U15767 (N_15767,N_12326,N_12744);
xor U15768 (N_15768,N_13420,N_12662);
nor U15769 (N_15769,N_12787,N_13927);
nor U15770 (N_15770,N_13755,N_13588);
nand U15771 (N_15771,N_12152,N_12969);
and U15772 (N_15772,N_12607,N_12786);
nand U15773 (N_15773,N_13724,N_13994);
nor U15774 (N_15774,N_13811,N_12765);
or U15775 (N_15775,N_12893,N_13034);
and U15776 (N_15776,N_13989,N_12257);
and U15777 (N_15777,N_12588,N_12472);
or U15778 (N_15778,N_12057,N_13706);
xor U15779 (N_15779,N_12773,N_13375);
and U15780 (N_15780,N_12989,N_13218);
nand U15781 (N_15781,N_12066,N_13890);
nand U15782 (N_15782,N_13283,N_13308);
nor U15783 (N_15783,N_13742,N_13882);
nor U15784 (N_15784,N_13782,N_13923);
nor U15785 (N_15785,N_12406,N_13707);
and U15786 (N_15786,N_13316,N_13459);
or U15787 (N_15787,N_13979,N_13397);
or U15788 (N_15788,N_12170,N_13736);
and U15789 (N_15789,N_13212,N_13231);
or U15790 (N_15790,N_13298,N_12540);
nand U15791 (N_15791,N_13014,N_12636);
nand U15792 (N_15792,N_13826,N_12621);
nand U15793 (N_15793,N_13305,N_13317);
xnor U15794 (N_15794,N_12143,N_12093);
nor U15795 (N_15795,N_12667,N_13583);
xnor U15796 (N_15796,N_12004,N_13190);
nand U15797 (N_15797,N_13101,N_13779);
nand U15798 (N_15798,N_13843,N_12622);
or U15799 (N_15799,N_12395,N_13023);
nor U15800 (N_15800,N_13649,N_12498);
and U15801 (N_15801,N_12155,N_13847);
and U15802 (N_15802,N_12982,N_12925);
nor U15803 (N_15803,N_12530,N_13342);
nand U15804 (N_15804,N_12468,N_12817);
nor U15805 (N_15805,N_13250,N_13037);
and U15806 (N_15806,N_12265,N_13576);
and U15807 (N_15807,N_12094,N_12738);
nor U15808 (N_15808,N_12687,N_13729);
and U15809 (N_15809,N_12644,N_12570);
and U15810 (N_15810,N_13418,N_13141);
nand U15811 (N_15811,N_13114,N_13060);
or U15812 (N_15812,N_13461,N_13206);
and U15813 (N_15813,N_12722,N_12090);
or U15814 (N_15814,N_12152,N_13610);
and U15815 (N_15815,N_13320,N_12908);
and U15816 (N_15816,N_13627,N_13582);
nand U15817 (N_15817,N_13852,N_13280);
or U15818 (N_15818,N_12513,N_13887);
nand U15819 (N_15819,N_12869,N_13042);
nand U15820 (N_15820,N_13894,N_12377);
and U15821 (N_15821,N_13031,N_12015);
or U15822 (N_15822,N_13227,N_12199);
and U15823 (N_15823,N_12245,N_13131);
nor U15824 (N_15824,N_12683,N_13631);
nand U15825 (N_15825,N_12144,N_12448);
nor U15826 (N_15826,N_13783,N_12747);
or U15827 (N_15827,N_13647,N_13178);
nor U15828 (N_15828,N_13672,N_13337);
or U15829 (N_15829,N_13507,N_12883);
and U15830 (N_15830,N_13300,N_12779);
and U15831 (N_15831,N_13657,N_13077);
or U15832 (N_15832,N_13286,N_12741);
or U15833 (N_15833,N_12589,N_13394);
and U15834 (N_15834,N_13494,N_13199);
and U15835 (N_15835,N_13451,N_12574);
and U15836 (N_15836,N_13234,N_12900);
nor U15837 (N_15837,N_13725,N_13290);
and U15838 (N_15838,N_12659,N_13978);
xor U15839 (N_15839,N_13902,N_13791);
and U15840 (N_15840,N_13986,N_12556);
and U15841 (N_15841,N_12120,N_13385);
nand U15842 (N_15842,N_13184,N_12541);
nand U15843 (N_15843,N_13552,N_12169);
nand U15844 (N_15844,N_13692,N_13260);
and U15845 (N_15845,N_13497,N_12319);
nand U15846 (N_15846,N_12225,N_12471);
and U15847 (N_15847,N_12911,N_13862);
or U15848 (N_15848,N_12731,N_13583);
xnor U15849 (N_15849,N_12229,N_13574);
nand U15850 (N_15850,N_12262,N_12182);
nand U15851 (N_15851,N_12292,N_12705);
nor U15852 (N_15852,N_13832,N_13309);
nor U15853 (N_15853,N_12765,N_13515);
nor U15854 (N_15854,N_12204,N_12371);
and U15855 (N_15855,N_12128,N_13104);
nor U15856 (N_15856,N_12240,N_12044);
or U15857 (N_15857,N_12160,N_13263);
or U15858 (N_15858,N_12785,N_13832);
and U15859 (N_15859,N_12652,N_12904);
nor U15860 (N_15860,N_13147,N_12696);
or U15861 (N_15861,N_13675,N_13733);
nand U15862 (N_15862,N_13103,N_13637);
or U15863 (N_15863,N_12130,N_12406);
nand U15864 (N_15864,N_13895,N_13092);
or U15865 (N_15865,N_12629,N_12493);
nand U15866 (N_15866,N_13236,N_12179);
and U15867 (N_15867,N_13987,N_12905);
nor U15868 (N_15868,N_13689,N_12190);
or U15869 (N_15869,N_13235,N_13253);
and U15870 (N_15870,N_13649,N_12326);
nand U15871 (N_15871,N_12117,N_13768);
nor U15872 (N_15872,N_13498,N_13951);
xnor U15873 (N_15873,N_12483,N_12245);
xnor U15874 (N_15874,N_12403,N_13336);
nand U15875 (N_15875,N_13631,N_12339);
nor U15876 (N_15876,N_13897,N_13881);
and U15877 (N_15877,N_12873,N_13264);
or U15878 (N_15878,N_12597,N_12206);
and U15879 (N_15879,N_12059,N_12713);
or U15880 (N_15880,N_12480,N_13703);
xor U15881 (N_15881,N_13078,N_12390);
or U15882 (N_15882,N_12599,N_13079);
nand U15883 (N_15883,N_12213,N_12635);
and U15884 (N_15884,N_12490,N_13638);
or U15885 (N_15885,N_13402,N_12115);
nand U15886 (N_15886,N_12215,N_13066);
or U15887 (N_15887,N_13435,N_13967);
or U15888 (N_15888,N_12691,N_13650);
nor U15889 (N_15889,N_13124,N_13777);
nor U15890 (N_15890,N_12619,N_12267);
xnor U15891 (N_15891,N_12834,N_13787);
nand U15892 (N_15892,N_13361,N_13309);
nor U15893 (N_15893,N_12749,N_13358);
xor U15894 (N_15894,N_12971,N_12049);
nand U15895 (N_15895,N_12041,N_13595);
or U15896 (N_15896,N_12585,N_13812);
nand U15897 (N_15897,N_12799,N_12647);
xnor U15898 (N_15898,N_12285,N_12977);
xnor U15899 (N_15899,N_13288,N_13400);
xor U15900 (N_15900,N_13303,N_12510);
nor U15901 (N_15901,N_13558,N_13313);
xor U15902 (N_15902,N_13951,N_12232);
xor U15903 (N_15903,N_12124,N_13879);
nor U15904 (N_15904,N_12208,N_12764);
and U15905 (N_15905,N_12312,N_13865);
xor U15906 (N_15906,N_13311,N_12050);
and U15907 (N_15907,N_13893,N_12058);
or U15908 (N_15908,N_13801,N_13989);
or U15909 (N_15909,N_13774,N_13444);
nand U15910 (N_15910,N_12266,N_13148);
xor U15911 (N_15911,N_13546,N_13322);
and U15912 (N_15912,N_13566,N_13202);
and U15913 (N_15913,N_12479,N_13448);
nor U15914 (N_15914,N_13430,N_13616);
nor U15915 (N_15915,N_12130,N_12318);
and U15916 (N_15916,N_12305,N_12367);
nand U15917 (N_15917,N_13630,N_12320);
and U15918 (N_15918,N_13764,N_13465);
nand U15919 (N_15919,N_12094,N_12835);
nand U15920 (N_15920,N_13899,N_12953);
or U15921 (N_15921,N_12627,N_12135);
nand U15922 (N_15922,N_13664,N_12776);
and U15923 (N_15923,N_12855,N_12439);
nand U15924 (N_15924,N_12289,N_12630);
and U15925 (N_15925,N_13456,N_13351);
nand U15926 (N_15926,N_12227,N_12377);
xor U15927 (N_15927,N_12628,N_12924);
xor U15928 (N_15928,N_13698,N_13987);
nand U15929 (N_15929,N_13377,N_13522);
nand U15930 (N_15930,N_12717,N_12583);
and U15931 (N_15931,N_12580,N_13066);
xor U15932 (N_15932,N_12478,N_12392);
or U15933 (N_15933,N_13088,N_13203);
nand U15934 (N_15934,N_12416,N_13891);
nand U15935 (N_15935,N_12115,N_12082);
xor U15936 (N_15936,N_12838,N_13126);
and U15937 (N_15937,N_12996,N_12133);
or U15938 (N_15938,N_12966,N_13532);
nand U15939 (N_15939,N_12454,N_12372);
and U15940 (N_15940,N_12735,N_13268);
and U15941 (N_15941,N_12794,N_13320);
nand U15942 (N_15942,N_12282,N_12715);
nand U15943 (N_15943,N_12483,N_12833);
nor U15944 (N_15944,N_13068,N_12890);
nand U15945 (N_15945,N_12330,N_13765);
or U15946 (N_15946,N_12863,N_13693);
or U15947 (N_15947,N_13393,N_12137);
or U15948 (N_15948,N_13127,N_13848);
and U15949 (N_15949,N_13410,N_13819);
nor U15950 (N_15950,N_13912,N_12905);
nor U15951 (N_15951,N_13109,N_13784);
and U15952 (N_15952,N_13368,N_12558);
and U15953 (N_15953,N_13782,N_12511);
nor U15954 (N_15954,N_13371,N_12410);
or U15955 (N_15955,N_13899,N_13999);
nor U15956 (N_15956,N_13044,N_13574);
or U15957 (N_15957,N_12626,N_12157);
or U15958 (N_15958,N_12569,N_12417);
nor U15959 (N_15959,N_13050,N_13070);
nor U15960 (N_15960,N_12255,N_12085);
nand U15961 (N_15961,N_13136,N_12708);
or U15962 (N_15962,N_13899,N_12533);
and U15963 (N_15963,N_12404,N_12989);
nor U15964 (N_15964,N_13891,N_13038);
and U15965 (N_15965,N_13088,N_13706);
and U15966 (N_15966,N_13557,N_12444);
nor U15967 (N_15967,N_12564,N_12358);
xor U15968 (N_15968,N_12485,N_13835);
nor U15969 (N_15969,N_12151,N_12997);
and U15970 (N_15970,N_13780,N_13149);
nor U15971 (N_15971,N_12710,N_13970);
nor U15972 (N_15972,N_12838,N_12730);
nor U15973 (N_15973,N_12153,N_12162);
or U15974 (N_15974,N_13087,N_12935);
nand U15975 (N_15975,N_12874,N_13236);
nand U15976 (N_15976,N_12630,N_12687);
xnor U15977 (N_15977,N_12316,N_12463);
nor U15978 (N_15978,N_12804,N_12943);
nand U15979 (N_15979,N_13812,N_12292);
and U15980 (N_15980,N_13428,N_12393);
and U15981 (N_15981,N_13475,N_12135);
nor U15982 (N_15982,N_12781,N_12459);
or U15983 (N_15983,N_13974,N_13381);
and U15984 (N_15984,N_13188,N_12457);
nand U15985 (N_15985,N_13691,N_13392);
and U15986 (N_15986,N_13260,N_12721);
nand U15987 (N_15987,N_12009,N_13285);
and U15988 (N_15988,N_13666,N_12964);
or U15989 (N_15989,N_13547,N_13280);
nand U15990 (N_15990,N_12668,N_13537);
and U15991 (N_15991,N_12764,N_13146);
xor U15992 (N_15992,N_12188,N_12089);
or U15993 (N_15993,N_12372,N_13443);
nor U15994 (N_15994,N_13345,N_12563);
xnor U15995 (N_15995,N_13768,N_13082);
nor U15996 (N_15996,N_12656,N_12627);
nor U15997 (N_15997,N_12434,N_13808);
and U15998 (N_15998,N_12350,N_12393);
or U15999 (N_15999,N_12445,N_12073);
and U16000 (N_16000,N_14336,N_14856);
nand U16001 (N_16001,N_14561,N_15412);
nor U16002 (N_16002,N_14044,N_15806);
nand U16003 (N_16003,N_15071,N_15441);
nor U16004 (N_16004,N_15431,N_14032);
and U16005 (N_16005,N_15583,N_15502);
nand U16006 (N_16006,N_14004,N_15773);
and U16007 (N_16007,N_14490,N_14277);
nor U16008 (N_16008,N_14242,N_15152);
or U16009 (N_16009,N_14581,N_14025);
nand U16010 (N_16010,N_15627,N_15788);
nor U16011 (N_16011,N_14316,N_14462);
or U16012 (N_16012,N_14565,N_14435);
or U16013 (N_16013,N_14546,N_14501);
nor U16014 (N_16014,N_14439,N_15758);
or U16015 (N_16015,N_14793,N_15260);
nand U16016 (N_16016,N_14589,N_14408);
or U16017 (N_16017,N_15148,N_15452);
nor U16018 (N_16018,N_15633,N_15369);
nand U16019 (N_16019,N_15008,N_14094);
or U16020 (N_16020,N_15537,N_14688);
and U16021 (N_16021,N_14558,N_14517);
and U16022 (N_16022,N_14858,N_15529);
nor U16023 (N_16023,N_14058,N_15573);
nand U16024 (N_16024,N_14560,N_14878);
and U16025 (N_16025,N_14986,N_15415);
and U16026 (N_16026,N_14897,N_14876);
and U16027 (N_16027,N_15011,N_14474);
nor U16028 (N_16028,N_14243,N_15549);
or U16029 (N_16029,N_14397,N_15158);
nor U16030 (N_16030,N_14197,N_14742);
nor U16031 (N_16031,N_14750,N_14206);
nand U16032 (N_16032,N_14678,N_14342);
xor U16033 (N_16033,N_14670,N_15799);
and U16034 (N_16034,N_14607,N_15443);
nor U16035 (N_16035,N_15337,N_14028);
nand U16036 (N_16036,N_15893,N_14837);
or U16037 (N_16037,N_15681,N_14707);
xnor U16038 (N_16038,N_15669,N_15997);
nand U16039 (N_16039,N_15548,N_15182);
nor U16040 (N_16040,N_15798,N_15058);
or U16041 (N_16041,N_14403,N_14968);
nand U16042 (N_16042,N_14674,N_15559);
nor U16043 (N_16043,N_15654,N_14461);
and U16044 (N_16044,N_15905,N_15034);
or U16045 (N_16045,N_14606,N_15367);
nand U16046 (N_16046,N_14945,N_14161);
nor U16047 (N_16047,N_15046,N_14690);
nand U16048 (N_16048,N_15881,N_15590);
and U16049 (N_16049,N_15041,N_15777);
and U16050 (N_16050,N_15744,N_15283);
and U16051 (N_16051,N_15919,N_14761);
nor U16052 (N_16052,N_15749,N_14100);
nor U16053 (N_16053,N_14131,N_14812);
nand U16054 (N_16054,N_15585,N_15714);
xnor U16055 (N_16055,N_14913,N_15849);
or U16056 (N_16056,N_14465,N_14267);
nand U16057 (N_16057,N_15349,N_14709);
xnor U16058 (N_16058,N_14062,N_14413);
and U16059 (N_16059,N_14958,N_14220);
xor U16060 (N_16060,N_14425,N_15520);
and U16061 (N_16061,N_14360,N_15424);
xnor U16062 (N_16062,N_14308,N_14621);
nand U16063 (N_16063,N_15730,N_15747);
or U16064 (N_16064,N_14034,N_15699);
nand U16065 (N_16065,N_14522,N_14843);
nor U16066 (N_16066,N_14012,N_15380);
and U16067 (N_16067,N_15086,N_15159);
and U16068 (N_16068,N_14060,N_14999);
nand U16069 (N_16069,N_14226,N_15004);
and U16070 (N_16070,N_15293,N_14721);
or U16071 (N_16071,N_14971,N_15241);
and U16072 (N_16072,N_14427,N_14671);
and U16073 (N_16073,N_14792,N_15474);
or U16074 (N_16074,N_14973,N_15753);
nor U16075 (N_16075,N_14319,N_14450);
nand U16076 (N_16076,N_15936,N_15170);
or U16077 (N_16077,N_14230,N_15561);
or U16078 (N_16078,N_14163,N_14673);
and U16079 (N_16079,N_15056,N_15628);
nor U16080 (N_16080,N_15792,N_14079);
and U16081 (N_16081,N_15939,N_15718);
nand U16082 (N_16082,N_14748,N_14978);
nand U16083 (N_16083,N_14346,N_15707);
and U16084 (N_16084,N_14263,N_14251);
xnor U16085 (N_16085,N_14001,N_14315);
nand U16086 (N_16086,N_14572,N_14901);
nor U16087 (N_16087,N_15575,N_15751);
nor U16088 (N_16088,N_14874,N_14662);
nand U16089 (N_16089,N_14739,N_15832);
or U16090 (N_16090,N_14771,N_15683);
and U16091 (N_16091,N_14594,N_15602);
and U16092 (N_16092,N_14393,N_14337);
nand U16093 (N_16093,N_15787,N_15187);
xor U16094 (N_16094,N_14550,N_14066);
nor U16095 (N_16095,N_14563,N_14653);
nor U16096 (N_16096,N_15519,N_15780);
nor U16097 (N_16097,N_14406,N_14138);
or U16098 (N_16098,N_14357,N_14074);
nor U16099 (N_16099,N_14993,N_15358);
or U16100 (N_16100,N_14173,N_15295);
or U16101 (N_16101,N_14005,N_14189);
nor U16102 (N_16102,N_15605,N_14452);
and U16103 (N_16103,N_15425,N_14087);
xor U16104 (N_16104,N_14557,N_14362);
or U16105 (N_16105,N_15906,N_14312);
nor U16106 (N_16106,N_14836,N_14174);
nand U16107 (N_16107,N_15268,N_15272);
and U16108 (N_16108,N_15342,N_15965);
or U16109 (N_16109,N_15813,N_14193);
and U16110 (N_16110,N_14885,N_14859);
nand U16111 (N_16111,N_14642,N_15302);
or U16112 (N_16112,N_15735,N_14753);
or U16113 (N_16113,N_15517,N_14726);
nor U16114 (N_16114,N_15623,N_15454);
or U16115 (N_16115,N_14939,N_15870);
or U16116 (N_16116,N_14424,N_14283);
or U16117 (N_16117,N_14417,N_14054);
and U16118 (N_16118,N_15348,N_15174);
or U16119 (N_16119,N_15850,N_15661);
or U16120 (N_16120,N_14307,N_14834);
nor U16121 (N_16121,N_15782,N_14070);
nor U16122 (N_16122,N_15663,N_14137);
nor U16123 (N_16123,N_15866,N_14203);
or U16124 (N_16124,N_14727,N_15479);
nor U16125 (N_16125,N_14619,N_15088);
nor U16126 (N_16126,N_15442,N_15554);
xor U16127 (N_16127,N_14564,N_15809);
nand U16128 (N_16128,N_15713,N_15399);
nor U16129 (N_16129,N_15419,N_14962);
or U16130 (N_16130,N_14228,N_14281);
or U16131 (N_16131,N_15523,N_14373);
or U16132 (N_16132,N_14860,N_14593);
nand U16133 (N_16133,N_15667,N_15255);
nand U16134 (N_16134,N_14905,N_15157);
and U16135 (N_16135,N_15353,N_15609);
xnor U16136 (N_16136,N_14445,N_14447);
nand U16137 (N_16137,N_15971,N_15993);
nor U16138 (N_16138,N_15636,N_14575);
nor U16139 (N_16139,N_15259,N_15160);
xor U16140 (N_16140,N_14440,N_14227);
and U16141 (N_16141,N_14578,N_14795);
nand U16142 (N_16142,N_14341,N_14322);
xor U16143 (N_16143,N_15942,N_14358);
and U16144 (N_16144,N_14240,N_14912);
nor U16145 (N_16145,N_15469,N_14102);
and U16146 (N_16146,N_14253,N_15673);
nor U16147 (N_16147,N_14915,N_14588);
nor U16148 (N_16148,N_14365,N_14482);
or U16149 (N_16149,N_15384,N_15748);
nor U16150 (N_16150,N_15533,N_14190);
nor U16151 (N_16151,N_14259,N_14518);
xnor U16152 (N_16152,N_15334,N_15564);
nand U16153 (N_16153,N_15409,N_14198);
or U16154 (N_16154,N_15060,N_15113);
nand U16155 (N_16155,N_14504,N_15463);
or U16156 (N_16156,N_15134,N_15410);
or U16157 (N_16157,N_15389,N_15381);
nor U16158 (N_16158,N_14509,N_15625);
nand U16159 (N_16159,N_15242,N_15239);
or U16160 (N_16160,N_14029,N_15503);
or U16161 (N_16161,N_14676,N_14015);
nand U16162 (N_16162,N_14059,N_14486);
or U16163 (N_16163,N_14617,N_14496);
nor U16164 (N_16164,N_14171,N_15282);
and U16165 (N_16165,N_15542,N_14646);
and U16166 (N_16166,N_15974,N_15457);
and U16167 (N_16167,N_14115,N_14460);
nand U16168 (N_16168,N_15033,N_14489);
nor U16169 (N_16169,N_15488,N_14442);
and U16170 (N_16170,N_14983,N_14468);
and U16171 (N_16171,N_14271,N_14457);
xor U16172 (N_16172,N_15901,N_15446);
nor U16173 (N_16173,N_15770,N_15213);
and U16174 (N_16174,N_14738,N_14903);
and U16175 (N_16175,N_15948,N_14666);
and U16176 (N_16176,N_15240,N_15280);
nor U16177 (N_16177,N_14041,N_14906);
and U16178 (N_16178,N_15140,N_14743);
and U16179 (N_16179,N_15066,N_14667);
nand U16180 (N_16180,N_14080,N_14908);
and U16181 (N_16181,N_15721,N_14369);
nor U16182 (N_16182,N_15161,N_15087);
nor U16183 (N_16183,N_15217,N_15765);
nand U16184 (N_16184,N_14356,N_14233);
nor U16185 (N_16185,N_14311,N_15889);
nor U16186 (N_16186,N_15235,N_15385);
nand U16187 (N_16187,N_14825,N_15364);
nor U16188 (N_16188,N_15332,N_15729);
xor U16189 (N_16189,N_15914,N_14835);
and U16190 (N_16190,N_14953,N_15551);
nor U16191 (N_16191,N_15584,N_14869);
or U16192 (N_16192,N_15499,N_15432);
nor U16193 (N_16193,N_15902,N_14021);
xor U16194 (N_16194,N_15275,N_14791);
or U16195 (N_16195,N_15145,N_14849);
nor U16196 (N_16196,N_14261,N_14349);
xor U16197 (N_16197,N_15698,N_14776);
nand U16198 (N_16198,N_15245,N_14188);
or U16199 (N_16199,N_14716,N_14555);
or U16200 (N_16200,N_14257,N_14567);
and U16201 (N_16201,N_14615,N_15422);
and U16202 (N_16202,N_15444,N_15124);
and U16203 (N_16203,N_14980,N_14275);
or U16204 (N_16204,N_15007,N_14057);
and U16205 (N_16205,N_14286,N_14954);
nor U16206 (N_16206,N_14643,N_14347);
nor U16207 (N_16207,N_15279,N_15171);
and U16208 (N_16208,N_15691,N_14067);
or U16209 (N_16209,N_15390,N_14657);
and U16210 (N_16210,N_15818,N_15518);
xor U16211 (N_16211,N_14212,N_14782);
xnor U16212 (N_16212,N_15922,N_14630);
nand U16213 (N_16213,N_15843,N_14314);
and U16214 (N_16214,N_14331,N_14804);
nand U16215 (N_16215,N_15761,N_15677);
nand U16216 (N_16216,N_15556,N_14612);
nand U16217 (N_16217,N_15668,N_14252);
nand U16218 (N_16218,N_15992,N_15234);
or U16219 (N_16219,N_14078,N_15377);
and U16220 (N_16220,N_14754,N_15210);
nor U16221 (N_16221,N_14601,N_14478);
and U16222 (N_16222,N_14963,N_14184);
nor U16223 (N_16223,N_14807,N_14225);
and U16224 (N_16224,N_14103,N_15097);
nor U16225 (N_16225,N_15859,N_14819);
nand U16226 (N_16226,N_15986,N_15169);
nand U16227 (N_16227,N_15167,N_15897);
or U16228 (N_16228,N_14455,N_14881);
or U16229 (N_16229,N_15243,N_15652);
or U16230 (N_16230,N_14491,N_14135);
and U16231 (N_16231,N_14568,N_15231);
nor U16232 (N_16232,N_15076,N_15237);
and U16233 (N_16233,N_15393,N_14466);
or U16234 (N_16234,N_14351,N_15137);
nand U16235 (N_16235,N_14592,N_14152);
nor U16236 (N_16236,N_15980,N_15312);
and U16237 (N_16237,N_14877,N_15995);
nand U16238 (N_16238,N_15970,N_15614);
and U16239 (N_16239,N_14039,N_15065);
nand U16240 (N_16240,N_14177,N_14042);
nand U16241 (N_16241,N_15955,N_15769);
and U16242 (N_16242,N_14566,N_14632);
xnor U16243 (N_16243,N_15853,N_15362);
nor U16244 (N_16244,N_14096,N_14888);
nand U16245 (N_16245,N_14868,N_14472);
and U16246 (N_16246,N_15374,N_15990);
and U16247 (N_16247,N_15418,N_15984);
and U16248 (N_16248,N_15195,N_14543);
or U16249 (N_16249,N_15665,N_15851);
and U16250 (N_16250,N_14916,N_14763);
or U16251 (N_16251,N_14608,N_14961);
nor U16252 (N_16252,N_15299,N_14086);
nand U16253 (N_16253,N_15482,N_14158);
nor U16254 (N_16254,N_14562,N_15720);
nor U16255 (N_16255,N_14441,N_14810);
xnor U16256 (N_16256,N_15869,N_14757);
or U16257 (N_16257,N_14473,N_14165);
or U16258 (N_16258,N_15184,N_14960);
nand U16259 (N_16259,N_14285,N_15895);
and U16260 (N_16260,N_15156,N_14910);
nor U16261 (N_16261,N_15039,N_14605);
and U16262 (N_16262,N_15841,N_14048);
nor U16263 (N_16263,N_15733,N_14049);
nor U16264 (N_16264,N_15928,N_14924);
and U16265 (N_16265,N_15724,N_15998);
nor U16266 (N_16266,N_15305,N_14668);
nand U16267 (N_16267,N_14687,N_14118);
or U16268 (N_16268,N_14700,N_15596);
or U16269 (N_16269,N_14199,N_14778);
or U16270 (N_16270,N_15212,N_14772);
and U16271 (N_16271,N_14428,N_15028);
or U16272 (N_16272,N_14348,N_15608);
or U16273 (N_16273,N_15630,N_15968);
nor U16274 (N_16274,N_14416,N_15705);
and U16275 (N_16275,N_14631,N_14586);
nor U16276 (N_16276,N_15946,N_14647);
or U16277 (N_16277,N_15128,N_15094);
and U16278 (N_16278,N_14533,N_15979);
xnor U16279 (N_16279,N_14443,N_15983);
nor U16280 (N_16280,N_14796,N_14239);
nand U16281 (N_16281,N_15553,N_14531);
nand U16282 (N_16282,N_14523,N_15396);
nor U16283 (N_16283,N_14513,N_15168);
or U16284 (N_16284,N_15485,N_14683);
nand U16285 (N_16285,N_14585,N_15106);
nor U16286 (N_16286,N_14681,N_15301);
or U16287 (N_16287,N_14368,N_14061);
and U16288 (N_16288,N_14786,N_14372);
nor U16289 (N_16289,N_15460,N_14480);
xnor U16290 (N_16290,N_14651,N_15985);
nor U16291 (N_16291,N_15285,N_14987);
xnor U16292 (N_16292,N_14981,N_15453);
nor U16293 (N_16293,N_15373,N_14579);
and U16294 (N_16294,N_14056,N_14089);
xnor U16295 (N_16295,N_15513,N_15570);
or U16296 (N_16296,N_14528,N_15339);
nor U16297 (N_16297,N_15712,N_14011);
and U16298 (N_16298,N_14318,N_14300);
or U16299 (N_16299,N_15634,N_14390);
nand U16300 (N_16300,N_15219,N_15082);
and U16301 (N_16301,N_15030,N_15198);
or U16302 (N_16302,N_15571,N_14422);
nand U16303 (N_16303,N_14040,N_14355);
nand U16304 (N_16304,N_15021,N_15150);
nor U16305 (N_16305,N_15200,N_15956);
or U16306 (N_16306,N_14556,N_15202);
and U16307 (N_16307,N_15296,N_14733);
or U16308 (N_16308,N_15372,N_15582);
or U16309 (N_16309,N_14712,N_15805);
nand U16310 (N_16310,N_15797,N_15580);
or U16311 (N_16311,N_14182,N_15833);
nor U16312 (N_16312,N_15888,N_14409);
xor U16313 (N_16313,N_14569,N_15016);
xnor U16314 (N_16314,N_14031,N_14655);
nor U16315 (N_16315,N_15102,N_15643);
xor U16316 (N_16316,N_15105,N_14405);
nand U16317 (N_16317,N_14529,N_14296);
nand U16318 (N_16318,N_15686,N_15035);
and U16319 (N_16319,N_15904,N_15436);
nand U16320 (N_16320,N_14598,N_14280);
nand U16321 (N_16321,N_14400,N_14838);
nor U16322 (N_16322,N_15108,N_14321);
or U16323 (N_16323,N_15493,N_15692);
nand U16324 (N_16324,N_15639,N_15327);
or U16325 (N_16325,N_14515,N_15143);
nand U16326 (N_16326,N_15031,N_15051);
xor U16327 (N_16327,N_14803,N_14415);
nor U16328 (N_16328,N_14799,N_14429);
nand U16329 (N_16329,N_14583,N_15890);
nand U16330 (N_16330,N_15426,N_14185);
or U16331 (N_16331,N_14110,N_15680);
nand U16332 (N_16332,N_15000,N_14144);
or U16333 (N_16333,N_15131,N_14142);
or U16334 (N_16334,N_15900,N_15702);
or U16335 (N_16335,N_14366,N_14340);
or U16336 (N_16336,N_14934,N_14840);
nor U16337 (N_16337,N_14007,N_15879);
and U16338 (N_16338,N_15656,N_14832);
nand U16339 (N_16339,N_15975,N_15915);
nor U16340 (N_16340,N_14749,N_14597);
nand U16341 (N_16341,N_15541,N_15802);
or U16342 (N_16342,N_15629,N_14374);
or U16343 (N_16343,N_14045,N_15024);
xor U16344 (N_16344,N_15052,N_14737);
or U16345 (N_16345,N_15209,N_14927);
nor U16346 (N_16346,N_15837,N_15416);
nor U16347 (N_16347,N_15586,N_14133);
nor U16348 (N_16348,N_15294,N_15945);
nand U16349 (N_16349,N_14191,N_15032);
and U16350 (N_16350,N_14932,N_14701);
and U16351 (N_16351,N_15943,N_14882);
nor U16352 (N_16352,N_14614,N_14183);
or U16353 (N_16353,N_15784,N_15764);
and U16354 (N_16354,N_14291,N_14991);
nor U16355 (N_16355,N_15827,N_15616);
and U16356 (N_16356,N_15601,N_15355);
nor U16357 (N_16357,N_15246,N_15675);
nor U16358 (N_16358,N_15599,N_15635);
nand U16359 (N_16359,N_15215,N_15188);
and U16360 (N_16360,N_15467,N_14814);
and U16361 (N_16361,N_14787,N_14935);
or U16362 (N_16362,N_15522,N_15081);
or U16363 (N_16363,N_14656,N_15164);
nand U16364 (N_16364,N_15069,N_14327);
or U16365 (N_16365,N_15844,N_15684);
or U16366 (N_16366,N_14205,N_14909);
or U16367 (N_16367,N_14446,N_15040);
and U16368 (N_16368,N_14436,N_14241);
nor U16369 (N_16369,N_15957,N_15121);
nor U16370 (N_16370,N_14279,N_14010);
nand U16371 (N_16371,N_15978,N_15546);
and U16372 (N_16372,N_14266,N_14487);
nor U16373 (N_16373,N_14353,N_15054);
nand U16374 (N_16374,N_14830,N_15696);
or U16375 (N_16375,N_14704,N_14887);
or U16376 (N_16376,N_14343,N_15501);
or U16377 (N_16377,N_14833,N_14535);
and U16378 (N_16378,N_15738,N_14985);
and U16379 (N_16379,N_14250,N_15961);
and U16380 (N_16380,N_14037,N_14904);
nor U16381 (N_16381,N_14534,N_14820);
nor U16382 (N_16382,N_14644,N_14124);
or U16383 (N_16383,N_15951,N_14591);
and U16384 (N_16384,N_15923,N_14485);
nand U16385 (N_16385,N_15394,N_14943);
and U16386 (N_16386,N_14976,N_14997);
and U16387 (N_16387,N_15185,N_15595);
nor U16388 (N_16388,N_14264,N_14722);
or U16389 (N_16389,N_14549,N_14289);
nor U16390 (N_16390,N_15794,N_15593);
or U16391 (N_16391,N_15898,N_15743);
nand U16392 (N_16392,N_15531,N_14870);
and U16393 (N_16393,N_14313,N_14375);
and U16394 (N_16394,N_15703,N_15083);
and U16395 (N_16395,N_15080,N_14800);
nand U16396 (N_16396,N_15288,N_15003);
and U16397 (N_16397,N_14990,N_14845);
and U16398 (N_16398,N_14853,N_15600);
or U16399 (N_16399,N_14329,N_15015);
nor U16400 (N_16400,N_14894,N_15804);
and U16401 (N_16401,N_15592,N_14641);
and U16402 (N_16402,N_15310,N_14276);
or U16403 (N_16403,N_14411,N_15896);
and U16404 (N_16404,N_14317,N_15456);
nand U16405 (N_16405,N_14036,N_15057);
or U16406 (N_16406,N_14889,N_14119);
or U16407 (N_16407,N_15341,N_14287);
or U16408 (N_16408,N_14950,N_14270);
xnor U16409 (N_16409,N_14724,N_14846);
and U16410 (N_16410,N_15067,N_14895);
nand U16411 (N_16411,N_15524,N_14571);
nand U16412 (N_16412,N_14675,N_15934);
and U16413 (N_16413,N_15973,N_15176);
xor U16414 (N_16414,N_15711,N_14109);
nand U16415 (N_16415,N_15528,N_14172);
nand U16416 (N_16416,N_14023,N_14129);
nor U16417 (N_16417,N_14539,N_15093);
nor U16418 (N_16418,N_15370,N_15731);
nand U16419 (N_16419,N_15642,N_14937);
xnor U16420 (N_16420,N_15823,N_14069);
or U16421 (N_16421,N_15434,N_15878);
nand U16422 (N_16422,N_14731,N_14992);
or U16423 (N_16423,N_14995,N_14302);
nor U16424 (N_16424,N_15194,N_15112);
nor U16425 (N_16425,N_14774,N_15578);
nand U16426 (N_16426,N_14364,N_15835);
nor U16427 (N_16427,N_14214,N_14444);
xor U16428 (N_16428,N_15745,N_14946);
nor U16429 (N_16429,N_14952,N_14577);
nand U16430 (N_16430,N_14524,N_14180);
nand U16431 (N_16431,N_15173,N_15371);
or U16432 (N_16432,N_15262,N_15572);
xnor U16433 (N_16433,N_14951,N_15096);
or U16434 (N_16434,N_14116,N_15812);
nand U16435 (N_16435,N_15695,N_14175);
and U16436 (N_16436,N_14827,N_14097);
and U16437 (N_16437,N_15512,N_14505);
nand U16438 (N_16438,N_15865,N_14050);
nor U16439 (N_16439,N_14745,N_15196);
nor U16440 (N_16440,N_14328,N_15954);
or U16441 (N_16441,N_14552,N_15658);
or U16442 (N_16442,N_14117,N_14122);
or U16443 (N_16443,N_15828,N_15289);
xnor U16444 (N_16444,N_14256,N_14652);
nor U16445 (N_16445,N_14431,N_15292);
xor U16446 (N_16446,N_15976,N_14649);
nor U16447 (N_16447,N_14231,N_14719);
nor U16448 (N_16448,N_14284,N_14498);
and U16449 (N_16449,N_14363,N_14817);
xor U16450 (N_16450,N_14326,N_15644);
and U16451 (N_16451,N_15473,N_15500);
or U16452 (N_16452,N_15653,N_15248);
nor U16453 (N_16453,N_14600,N_15461);
nor U16454 (N_16454,N_14027,N_15911);
and U16455 (N_16455,N_15350,N_15206);
nor U16456 (N_16456,N_14736,N_15563);
nor U16457 (N_16457,N_15162,N_14956);
or U16458 (N_16458,N_15382,N_15871);
nand U16459 (N_16459,N_15181,N_15615);
nor U16460 (N_16460,N_15750,N_14638);
xnor U16461 (N_16461,N_14294,N_15138);
or U16462 (N_16462,N_14107,N_14650);
and U16463 (N_16463,N_15264,N_15830);
and U16464 (N_16464,N_15801,N_14017);
nand U16465 (N_16465,N_15119,N_14922);
or U16466 (N_16466,N_14038,N_15064);
or U16467 (N_16467,N_15892,N_15505);
nor U16468 (N_16468,N_15756,N_15178);
and U16469 (N_16469,N_15821,N_15613);
nand U16470 (N_16470,N_15950,N_14634);
nor U16471 (N_16471,N_14580,N_14223);
and U16472 (N_16472,N_14179,N_15886);
and U16473 (N_16473,N_14187,N_14695);
and U16474 (N_16474,N_14146,N_14636);
nand U16475 (N_16475,N_14325,N_14371);
nand U16476 (N_16476,N_14113,N_15079);
nand U16477 (N_16477,N_15981,N_14862);
or U16478 (N_16478,N_14758,N_15315);
nor U16479 (N_16479,N_14269,N_15638);
or U16480 (N_16480,N_15803,N_15917);
nand U16481 (N_16481,N_14728,N_14537);
xor U16482 (N_16482,N_14640,N_14711);
xor U16483 (N_16483,N_15438,N_14940);
or U16484 (N_16484,N_15376,N_14414);
xnor U16485 (N_16485,N_15462,N_15701);
or U16486 (N_16486,N_15877,N_14768);
nor U16487 (N_16487,N_14033,N_14141);
or U16488 (N_16488,N_15100,N_15214);
nand U16489 (N_16489,N_14752,N_14162);
nor U16490 (N_16490,N_14682,N_15190);
nand U16491 (N_16491,N_15130,N_15736);
nor U16492 (N_16492,N_14430,N_15723);
and U16493 (N_16493,N_14379,N_14570);
nand U16494 (N_16494,N_15648,N_14469);
and U16495 (N_16495,N_14419,N_15487);
or U16496 (N_16496,N_14923,N_15579);
nand U16497 (N_16497,N_14710,N_15300);
nor U16498 (N_16498,N_15754,N_15786);
nand U16499 (N_16499,N_14884,N_14516);
nand U16500 (N_16500,N_15063,N_15347);
and U16501 (N_16501,N_15423,N_15375);
or U16502 (N_16502,N_14030,N_15953);
or U16503 (N_16503,N_15155,N_15365);
xnor U16504 (N_16504,N_15962,N_15498);
nand U16505 (N_16505,N_14850,N_15256);
or U16506 (N_16506,N_14599,N_14551);
and U16507 (N_16507,N_15147,N_15047);
nand U16508 (N_16508,N_15958,N_14729);
or U16509 (N_16509,N_15103,N_15455);
and U16510 (N_16510,N_14548,N_14627);
nand U16511 (N_16511,N_15941,N_14775);
nand U16512 (N_16512,N_15427,N_15550);
nor U16513 (N_16513,N_15133,N_14128);
and U16514 (N_16514,N_14407,N_14169);
and U16515 (N_16515,N_15604,N_15552);
xor U16516 (N_16516,N_15224,N_14767);
nand U16517 (N_16517,N_14944,N_15254);
nor U16518 (N_16518,N_15343,N_14385);
and U16519 (N_16519,N_14892,N_14016);
or U16520 (N_16520,N_15038,N_15336);
nor U16521 (N_16521,N_14022,N_15739);
nor U16522 (N_16522,N_14273,N_15111);
and U16523 (N_16523,N_15316,N_15811);
or U16524 (N_16524,N_14633,N_15920);
and U16525 (N_16525,N_14477,N_15311);
nand U16526 (N_16526,N_15603,N_15783);
and U16527 (N_16527,N_14111,N_15776);
and U16528 (N_16528,N_14121,N_14635);
xnor U16529 (N_16529,N_15197,N_14809);
or U16530 (N_16530,N_15208,N_15061);
nor U16531 (N_16531,N_15331,N_14399);
xor U16532 (N_16532,N_14802,N_14301);
nor U16533 (N_16533,N_14201,N_14766);
xnor U16534 (N_16534,N_14933,N_14507);
and U16535 (N_16535,N_15304,N_15359);
or U16536 (N_16536,N_15340,N_15972);
or U16537 (N_16537,N_15645,N_14808);
nor U16538 (N_16538,N_14967,N_14765);
nand U16539 (N_16539,N_15746,N_14154);
nand U16540 (N_16540,N_15921,N_15391);
xor U16541 (N_16541,N_15117,N_14931);
or U16542 (N_16542,N_15048,N_14381);
and U16543 (N_16543,N_14759,N_15250);
and U16544 (N_16544,N_14898,N_15937);
or U16545 (N_16545,N_15072,N_15075);
nor U16546 (N_16546,N_15022,N_14900);
or U16547 (N_16547,N_15598,N_15508);
or U16548 (N_16548,N_15144,N_15688);
nor U16549 (N_16549,N_15029,N_14783);
nor U16550 (N_16550,N_15309,N_15126);
xnor U16551 (N_16551,N_14150,N_14204);
xnor U16552 (N_16552,N_14178,N_15507);
nor U16553 (N_16553,N_15284,N_15481);
nand U16554 (N_16554,N_14333,N_15538);
nor U16555 (N_16555,N_14218,N_15949);
nand U16556 (N_16556,N_14616,N_14713);
or U16557 (N_16557,N_15314,N_14009);
and U16558 (N_16558,N_14964,N_14497);
nor U16559 (N_16559,N_14780,N_14723);
nor U16560 (N_16560,N_15509,N_15516);
and U16561 (N_16561,N_14104,N_15617);
and U16562 (N_16562,N_14458,N_15940);
nor U16563 (N_16563,N_15495,N_14930);
or U16564 (N_16564,N_15233,N_15876);
nor U16565 (N_16565,N_14789,N_14519);
nor U16566 (N_16566,N_14665,N_15741);
xnor U16567 (N_16567,N_15660,N_15351);
nor U16568 (N_16568,N_15591,N_15848);
nand U16569 (N_16569,N_15388,N_14434);
nor U16570 (N_16570,N_15435,N_15023);
and U16571 (N_16571,N_15321,N_15840);
and U16572 (N_16572,N_15361,N_15858);
and U16573 (N_16573,N_14977,N_14698);
nor U16574 (N_16574,N_15662,N_15291);
and U16575 (N_16575,N_14391,N_14829);
nand U16576 (N_16576,N_14278,N_14207);
and U16577 (N_16577,N_14604,N_14229);
or U16578 (N_16578,N_14857,N_15092);
nand U16579 (N_16579,N_15287,N_14918);
nand U16580 (N_16580,N_14064,N_14000);
nand U16581 (N_16581,N_15611,N_15228);
nor U16582 (N_16582,N_15139,N_15055);
and U16583 (N_16583,N_14730,N_15191);
and U16584 (N_16584,N_14396,N_14216);
nor U16585 (N_16585,N_15597,N_15346);
or U16586 (N_16586,N_14512,N_14663);
or U16587 (N_16587,N_15118,N_15569);
nand U16588 (N_16588,N_14970,N_14831);
nand U16589 (N_16589,N_14156,N_14969);
and U16590 (N_16590,N_15856,N_14493);
or U16591 (N_16591,N_14153,N_14899);
nor U16592 (N_16592,N_14367,N_15253);
xor U16593 (N_16593,N_15966,N_14035);
or U16594 (N_16594,N_14088,N_14818);
or U16595 (N_16595,N_15449,N_15471);
or U16596 (N_16596,N_15925,N_14658);
xor U16597 (N_16597,N_15084,N_14288);
nand U16598 (N_16598,N_14813,N_14324);
xor U16599 (N_16599,N_14260,N_14404);
nand U16600 (N_16600,N_14875,N_15014);
or U16601 (N_16601,N_15760,N_15478);
nor U16602 (N_16602,N_14692,N_14526);
nor U16603 (N_16603,N_15318,N_15298);
and U16604 (N_16604,N_15791,N_15447);
nor U16605 (N_16605,N_14083,N_15496);
nor U16606 (N_16606,N_15091,N_15335);
or U16607 (N_16607,N_15223,N_15179);
and U16608 (N_16608,N_15562,N_14538);
nor U16609 (N_16609,N_14603,N_14382);
and U16610 (N_16610,N_14982,N_14618);
and U16611 (N_16611,N_14844,N_15618);
nor U16612 (N_16612,N_15952,N_14412);
nor U16613 (N_16613,N_14148,N_14388);
nand U16614 (N_16614,N_14865,N_14684);
or U16615 (N_16615,N_15996,N_15269);
nand U16616 (N_16616,N_14705,N_15098);
nand U16617 (N_16617,N_15480,N_15737);
nand U16618 (N_16618,N_15115,N_14941);
nor U16619 (N_16619,N_15429,N_15543);
or U16620 (N_16620,N_14541,N_15544);
or U16621 (N_16621,N_15672,N_15059);
nand U16622 (N_16622,N_15323,N_15308);
nand U16623 (N_16623,N_15817,N_15402);
nand U16624 (N_16624,N_15319,N_14265);
and U16625 (N_16625,N_14101,N_15816);
nor U16626 (N_16626,N_14483,N_15854);
or U16627 (N_16627,N_15400,N_14290);
nand U16628 (N_16628,N_15440,N_15666);
nand U16629 (N_16629,N_14664,N_14864);
or U16630 (N_16630,N_15655,N_15967);
xnor U16631 (N_16631,N_15464,N_15710);
nand U16632 (N_16632,N_14925,N_14330);
and U16633 (N_16633,N_15560,N_15037);
nor U16634 (N_16634,N_15430,N_14902);
nor U16635 (N_16635,N_14454,N_14624);
nand U16636 (N_16636,N_14420,N_14208);
nand U16637 (N_16637,N_15244,N_14975);
nand U16638 (N_16638,N_14988,N_14718);
xor U16639 (N_16639,N_15330,N_14166);
xor U16640 (N_16640,N_15766,N_14691);
or U16641 (N_16641,N_15433,N_14866);
or U16642 (N_16642,N_14136,N_14254);
nand U16643 (N_16643,N_14741,N_15099);
and U16644 (N_16644,N_15175,N_15492);
nand U16645 (N_16645,N_14019,N_15822);
and U16646 (N_16646,N_14350,N_15774);
xor U16647 (N_16647,N_15068,N_15755);
nand U16648 (N_16648,N_14295,N_15328);
or U16649 (N_16649,N_15982,N_15271);
xor U16650 (N_16650,N_14911,N_14195);
nand U16651 (N_16651,N_15078,N_14090);
nor U16652 (N_16652,N_14693,N_14781);
and U16653 (N_16653,N_14433,N_15650);
or U16654 (N_16654,N_15413,N_14609);
and U16655 (N_16655,N_15685,N_14760);
and U16656 (N_16656,N_14735,N_14755);
or U16657 (N_16657,N_15565,N_15910);
nor U16658 (N_16658,N_14536,N_14159);
nand U16659 (N_16659,N_14510,N_14145);
nor U16660 (N_16660,N_15682,N_15326);
nor U16661 (N_16661,N_15875,N_14547);
or U16662 (N_16662,N_14068,N_14449);
or U16663 (N_16663,N_14972,N_15778);
nand U16664 (N_16664,N_15709,N_15193);
nand U16665 (N_16665,N_15727,N_14816);
xnor U16666 (N_16666,N_15401,N_14451);
nor U16667 (N_16667,N_14576,N_14209);
and U16668 (N_16668,N_14706,N_14297);
and U16669 (N_16669,N_14130,N_14361);
and U16670 (N_16670,N_15222,N_14886);
or U16671 (N_16671,N_15366,N_14339);
or U16672 (N_16672,N_14914,N_15763);
nand U16673 (N_16673,N_14625,N_15988);
or U16674 (N_16674,N_15860,N_15872);
and U16675 (N_16675,N_15290,N_15042);
or U16676 (N_16676,N_15510,N_14715);
and U16677 (N_16677,N_15504,N_14105);
or U16678 (N_16678,N_15540,N_14320);
and U16679 (N_16679,N_14785,N_14387);
nor U16680 (N_16680,N_15236,N_15815);
or U16681 (N_16681,N_15693,N_15506);
and U16682 (N_16682,N_14221,N_15964);
and U16683 (N_16683,N_15428,N_15511);
nand U16684 (N_16684,N_15205,N_14861);
nand U16685 (N_16685,N_14626,N_15344);
and U16686 (N_16686,N_15793,N_15490);
nor U16687 (N_16687,N_14779,N_15368);
or U16688 (N_16688,N_14584,N_14126);
nor U16689 (N_16689,N_15525,N_15722);
nand U16690 (N_16690,N_15790,N_14732);
xor U16691 (N_16691,N_15862,N_14127);
nor U16692 (N_16692,N_15360,N_15932);
nand U16693 (N_16693,N_15908,N_15220);
nand U16694 (N_16694,N_14893,N_14092);
nor U16695 (N_16695,N_15530,N_15417);
nor U16696 (N_16696,N_14344,N_15676);
or U16697 (N_16697,N_14573,N_15470);
nor U16698 (N_16698,N_14680,N_14725);
xnor U16699 (N_16699,N_14305,N_15297);
nand U16700 (N_16700,N_15826,N_15883);
nor U16701 (N_16701,N_14359,N_14648);
or U16702 (N_16702,N_15322,N_15249);
and U16703 (N_16703,N_14699,N_14484);
xnor U16704 (N_16704,N_15532,N_14703);
and U16705 (N_16705,N_15820,N_14395);
nor U16706 (N_16706,N_14542,N_15847);
or U16707 (N_16707,N_15880,N_15670);
nand U16708 (N_16708,N_14076,N_14770);
or U16709 (N_16709,N_15286,N_14151);
xor U16710 (N_16710,N_14114,N_15218);
nand U16711 (N_16711,N_14024,N_14611);
xnor U16712 (N_16712,N_15270,N_14677);
or U16713 (N_16713,N_15810,N_15136);
and U16714 (N_16714,N_15477,N_14764);
or U16715 (N_16715,N_14996,N_15539);
nor U16716 (N_16716,N_14494,N_14181);
nand U16717 (N_16717,N_15742,N_14421);
or U16718 (N_16718,N_14052,N_14574);
nand U16719 (N_16719,N_15363,N_14863);
xnor U16720 (N_16720,N_15407,N_14530);
and U16721 (N_16721,N_15439,N_14160);
or U16722 (N_16722,N_14075,N_15594);
nor U16723 (N_16723,N_15010,N_15789);
or U16724 (N_16724,N_14920,N_15013);
nand U16725 (N_16725,N_14046,N_15252);
nand U16726 (N_16726,N_15527,N_15947);
nand U16727 (N_16727,N_14237,N_15725);
and U16728 (N_16728,N_14467,N_15345);
or U16729 (N_16729,N_14352,N_14426);
xor U16730 (N_16730,N_15587,N_15306);
nand U16731 (N_16731,N_15406,N_14746);
nor U16732 (N_16732,N_14232,N_15887);
and U16733 (N_16733,N_14306,N_14410);
nand U16734 (N_16734,N_15819,N_14756);
nand U16735 (N_16735,N_14282,N_14492);
nor U16736 (N_16736,N_14043,N_15626);
and U16737 (N_16737,N_15163,N_14448);
xor U16738 (N_16738,N_15225,N_15716);
and U16739 (N_16739,N_14432,N_14013);
xor U16740 (N_16740,N_14938,N_15172);
nor U16741 (N_16741,N_15386,N_15017);
or U16742 (N_16742,N_15090,N_15383);
or U16743 (N_16743,N_14471,N_14470);
and U16744 (N_16744,N_15036,N_15012);
nor U16745 (N_16745,N_14170,N_15451);
nor U16746 (N_16746,N_15005,N_15588);
and U16747 (N_16747,N_14377,N_15907);
and U16748 (N_16748,N_14694,N_14401);
nand U16749 (N_16749,N_14559,N_15153);
or U16750 (N_16750,N_15472,N_15273);
and U16751 (N_16751,N_14222,N_14773);
xor U16752 (N_16752,N_15397,N_14246);
nor U16753 (N_16753,N_14392,N_15929);
xor U16754 (N_16754,N_14847,N_14595);
or U16755 (N_16755,N_14801,N_14871);
xnor U16756 (N_16756,N_15873,N_14824);
nand U16757 (N_16757,N_15278,N_15944);
xor U16758 (N_16758,N_15867,N_14553);
or U16759 (N_16759,N_15785,N_15674);
or U16760 (N_16760,N_15891,N_14055);
or U16761 (N_16761,N_15281,N_14140);
and U16762 (N_16762,N_14098,N_14093);
nor U16763 (N_16763,N_14176,N_14091);
nand U16764 (N_16764,N_15664,N_14686);
nand U16765 (N_16765,N_15640,N_14697);
nor U16766 (N_16766,N_15885,N_15211);
xnor U16767 (N_16767,N_15489,N_14966);
and U16768 (N_16768,N_14544,N_15963);
nand U16769 (N_16769,N_14777,N_14402);
nor U16770 (N_16770,N_14823,N_14873);
and U16771 (N_16771,N_14891,N_15899);
or U16772 (N_16772,N_15095,N_15232);
or U16773 (N_16773,N_15317,N_14073);
nor U16774 (N_16774,N_14855,N_14955);
or U16775 (N_16775,N_14003,N_15107);
nand U16776 (N_16776,N_15192,N_15186);
nor U16777 (N_16777,N_15123,N_14155);
or U16778 (N_16778,N_14047,N_14811);
nand U16779 (N_16779,N_14132,N_15576);
or U16780 (N_16780,N_15557,N_15484);
and U16781 (N_16781,N_14112,N_14672);
nor U16782 (N_16782,N_15762,N_14797);
or U16783 (N_16783,N_14095,N_15129);
nor U16784 (N_16784,N_14645,N_14268);
nand U16785 (N_16785,N_14437,N_15894);
nand U16786 (N_16786,N_15637,N_14303);
nor U16787 (N_16787,N_14247,N_15475);
nor U16788 (N_16788,N_14628,N_14734);
and U16789 (N_16789,N_15230,N_15558);
and U16790 (N_16790,N_15912,N_14841);
nand U16791 (N_16791,N_15694,N_15049);
nor U16792 (N_16792,N_15001,N_14907);
nand U16793 (N_16793,N_14540,N_15357);
nand U16794 (N_16794,N_14453,N_15325);
and U16795 (N_16795,N_15933,N_15574);
nor U16796 (N_16796,N_15547,N_15732);
or U16797 (N_16797,N_14398,N_14545);
and U16798 (N_16798,N_15476,N_14848);
nand U16799 (N_16799,N_14679,N_15437);
and U16800 (N_16800,N_14508,N_15987);
nand U16801 (N_16801,N_15324,N_15606);
or U16802 (N_16802,N_14917,N_15109);
and U16803 (N_16803,N_15258,N_15831);
nor U16804 (N_16804,N_14926,N_14063);
and U16805 (N_16805,N_14500,N_15977);
and U16806 (N_16806,N_14805,N_15855);
nand U16807 (N_16807,N_14610,N_15641);
and U16808 (N_16808,N_15135,N_14249);
or U16809 (N_16809,N_15116,N_15276);
and U16810 (N_16810,N_14383,N_14929);
nor U16811 (N_16811,N_14720,N_15913);
nand U16812 (N_16812,N_15534,N_15465);
nand U16813 (N_16813,N_14394,N_14272);
nand U16814 (N_16814,N_14298,N_15483);
nor U16815 (N_16815,N_15146,N_15352);
nand U16816 (N_16816,N_14085,N_14702);
xnor U16817 (N_16817,N_15846,N_15568);
nor U16818 (N_16818,N_15839,N_15420);
and U16819 (N_16819,N_14502,N_14139);
nand U16820 (N_16820,N_14511,N_14389);
nand U16821 (N_16821,N_15612,N_15545);
and U16822 (N_16822,N_14806,N_15151);
nand U16823 (N_16823,N_14890,N_14077);
and U16824 (N_16824,N_14051,N_15740);
nor U16825 (N_16825,N_14143,N_15659);
nand U16826 (N_16826,N_14613,N_15610);
and U16827 (N_16827,N_15227,N_15927);
and U16828 (N_16828,N_15166,N_15303);
nor U16829 (N_16829,N_15277,N_15070);
or U16830 (N_16830,N_15808,N_14949);
nor U16831 (N_16831,N_15221,N_14659);
nor U16832 (N_16832,N_15189,N_15903);
nand U16833 (N_16833,N_15404,N_15313);
and U16834 (N_16834,N_15807,N_15581);
nand U16835 (N_16835,N_14590,N_15719);
or U16836 (N_16836,N_15589,N_14108);
or U16837 (N_16837,N_14790,N_15631);
and U16838 (N_16838,N_14488,N_15752);
nand U16839 (N_16839,N_14826,N_14217);
and U16840 (N_16840,N_14255,N_14192);
nand U16841 (N_16841,N_15577,N_15829);
xnor U16842 (N_16842,N_15649,N_14423);
and U16843 (N_16843,N_14639,N_15715);
nand U16844 (N_16844,N_15959,N_15909);
nand U16845 (N_16845,N_14018,N_14994);
nor U16846 (N_16846,N_15050,N_15053);
and U16847 (N_16847,N_15497,N_15387);
xnor U16848 (N_16848,N_15651,N_15657);
nand U16849 (N_16849,N_14919,N_15020);
and U16850 (N_16850,N_15999,N_15607);
or U16851 (N_16851,N_14506,N_14587);
xor U16852 (N_16852,N_15991,N_15916);
or U16853 (N_16853,N_14238,N_14200);
and U16854 (N_16854,N_14084,N_14008);
and U16855 (N_16855,N_14965,N_14525);
nor U16856 (N_16856,N_14872,N_14202);
or U16857 (N_16857,N_15204,N_15796);
nand U16858 (N_16858,N_14134,N_15632);
nor U16859 (N_16859,N_14002,N_15207);
nor U16860 (N_16860,N_15403,N_14338);
and U16861 (N_16861,N_15142,N_15960);
or U16862 (N_16862,N_14106,N_15926);
nor U16863 (N_16863,N_15814,N_14463);
or U16864 (N_16864,N_14464,N_14164);
xor U16865 (N_16865,N_14310,N_15445);
and U16866 (N_16866,N_15073,N_15333);
or U16867 (N_16867,N_15043,N_15226);
or U16868 (N_16868,N_14880,N_15825);
nand U16869 (N_16869,N_15154,N_15378);
or U16870 (N_16870,N_15536,N_15918);
and U16871 (N_16871,N_14532,N_14293);
or U16872 (N_16872,N_15180,N_15775);
nand U16873 (N_16873,N_14637,N_14157);
nand U16874 (N_16874,N_15085,N_15411);
or U16875 (N_16875,N_14224,N_15535);
nand U16876 (N_16876,N_15019,N_14685);
and U16877 (N_16877,N_15274,N_14386);
and U16878 (N_16878,N_15263,N_15408);
nand U16879 (N_16879,N_15622,N_14815);
nor U16880 (N_16880,N_14167,N_15356);
and U16881 (N_16881,N_14622,N_14006);
nor U16882 (N_16882,N_14274,N_14370);
or U16883 (N_16883,N_14186,N_15177);
nand U16884 (N_16884,N_15026,N_14883);
or U16885 (N_16885,N_15852,N_15120);
nor U16886 (N_16886,N_14762,N_15405);
nor U16887 (N_16887,N_15354,N_15767);
nand U16888 (N_16888,N_15863,N_14149);
or U16889 (N_16889,N_15938,N_14081);
and U16890 (N_16890,N_14828,N_14481);
xor U16891 (N_16891,N_15257,N_15687);
or U16892 (N_16892,N_15450,N_15935);
or U16893 (N_16893,N_14196,N_15141);
and U16894 (N_16894,N_14099,N_15619);
nand U16895 (N_16895,N_15884,N_14499);
and U16896 (N_16896,N_14747,N_14521);
or U16897 (N_16897,N_14354,N_15734);
nand U16898 (N_16898,N_15101,N_14947);
or U16899 (N_16899,N_14495,N_14065);
nand U16900 (N_16900,N_14194,N_14384);
nand U16901 (N_16901,N_14602,N_15044);
or U16902 (N_16902,N_14794,N_15772);
or U16903 (N_16903,N_15768,N_14989);
nand U16904 (N_16904,N_14788,N_15165);
nand U16905 (N_16905,N_14744,N_14669);
nor U16906 (N_16906,N_15216,N_14629);
nand U16907 (N_16907,N_15679,N_14654);
or U16908 (N_16908,N_14071,N_15700);
or U16909 (N_16909,N_14696,N_14120);
and U16910 (N_16910,N_14304,N_15781);
nor U16911 (N_16911,N_14438,N_14258);
xnor U16912 (N_16912,N_14380,N_15329);
and U16913 (N_16913,N_15646,N_14851);
or U16914 (N_16914,N_14376,N_15989);
nor U16915 (N_16915,N_15027,N_14211);
and U16916 (N_16916,N_15110,N_14514);
and U16917 (N_16917,N_14842,N_14854);
and U16918 (N_16918,N_15834,N_15521);
nor U16919 (N_16919,N_15006,N_14053);
nand U16920 (N_16920,N_14740,N_14234);
nor U16921 (N_16921,N_15199,N_15842);
or U16922 (N_16922,N_15708,N_15421);
or U16923 (N_16923,N_14520,N_15468);
nor U16924 (N_16924,N_15759,N_15690);
nand U16925 (N_16925,N_14751,N_15994);
or U16926 (N_16926,N_15229,N_15874);
or U16927 (N_16927,N_15491,N_15486);
nand U16928 (N_16928,N_15267,N_15074);
or U16929 (N_16929,N_15127,N_15671);
nor U16930 (N_16930,N_14852,N_14020);
or U16931 (N_16931,N_15089,N_15689);
nor U16932 (N_16932,N_15838,N_14026);
xor U16933 (N_16933,N_15122,N_14957);
nand U16934 (N_16934,N_15247,N_14948);
or U16935 (N_16935,N_15458,N_15002);
or U16936 (N_16936,N_14168,N_15836);
or U16937 (N_16937,N_15266,N_15931);
nor U16938 (N_16938,N_15466,N_15620);
or U16939 (N_16939,N_15555,N_14503);
and U16940 (N_16940,N_15624,N_15678);
nand U16941 (N_16941,N_14822,N_14921);
or U16942 (N_16942,N_14717,N_14959);
nand U16943 (N_16943,N_14125,N_15728);
nand U16944 (N_16944,N_14459,N_14244);
nor U16945 (N_16945,N_14147,N_14620);
or U16946 (N_16946,N_15930,N_15704);
or U16947 (N_16947,N_15104,N_14215);
and U16948 (N_16948,N_15924,N_15448);
nand U16949 (N_16949,N_14210,N_14798);
nand U16950 (N_16950,N_15882,N_15238);
xor U16951 (N_16951,N_15697,N_15132);
and U16952 (N_16952,N_14345,N_14839);
or U16953 (N_16953,N_15261,N_15861);
nand U16954 (N_16954,N_14292,N_15621);
and U16955 (N_16955,N_14476,N_14236);
nand U16956 (N_16956,N_15149,N_15515);
and U16957 (N_16957,N_14213,N_15757);
or U16958 (N_16958,N_15062,N_14582);
nor U16959 (N_16959,N_14689,N_15824);
nor U16960 (N_16960,N_14879,N_14378);
nor U16961 (N_16961,N_15717,N_15395);
or U16962 (N_16962,N_15414,N_15779);
nand U16963 (N_16963,N_15045,N_14979);
and U16964 (N_16964,N_15647,N_14245);
or U16965 (N_16965,N_14896,N_15526);
nand U16966 (N_16966,N_14309,N_14262);
and U16967 (N_16967,N_14479,N_15201);
nand U16968 (N_16968,N_15706,N_14072);
or U16969 (N_16969,N_15307,N_14596);
nor U16970 (N_16970,N_14418,N_15125);
nand U16971 (N_16971,N_15864,N_14936);
nor U16972 (N_16972,N_14235,N_15379);
nand U16973 (N_16973,N_14248,N_14998);
nand U16974 (N_16974,N_15459,N_15251);
or U16975 (N_16975,N_15857,N_14984);
xnor U16976 (N_16976,N_14867,N_14299);
or U16977 (N_16977,N_15114,N_14942);
or U16978 (N_16978,N_14714,N_14334);
and U16979 (N_16979,N_15203,N_15338);
nor U16980 (N_16980,N_15320,N_14475);
nor U16981 (N_16981,N_14928,N_14123);
or U16982 (N_16982,N_15800,N_14219);
and U16983 (N_16983,N_14335,N_14323);
nand U16984 (N_16984,N_14456,N_14784);
nand U16985 (N_16985,N_15771,N_14974);
nor U16986 (N_16986,N_15025,N_15969);
and U16987 (N_16987,N_14821,N_14623);
and U16988 (N_16988,N_15077,N_15392);
nor U16989 (N_16989,N_14554,N_15183);
and U16990 (N_16990,N_15845,N_14014);
nor U16991 (N_16991,N_14527,N_15018);
xor U16992 (N_16992,N_15265,N_15868);
nand U16993 (N_16993,N_14660,N_15494);
and U16994 (N_16994,N_15566,N_15009);
nand U16995 (N_16995,N_14082,N_15567);
and U16996 (N_16996,N_15514,N_14332);
xnor U16997 (N_16997,N_14661,N_15726);
and U16998 (N_16998,N_15398,N_14769);
and U16999 (N_16999,N_15795,N_14708);
or U17000 (N_17000,N_15601,N_14969);
nor U17001 (N_17001,N_15998,N_14919);
xor U17002 (N_17002,N_14312,N_14112);
or U17003 (N_17003,N_15323,N_15466);
xnor U17004 (N_17004,N_15021,N_15327);
xnor U17005 (N_17005,N_14286,N_15620);
nand U17006 (N_17006,N_14092,N_14022);
or U17007 (N_17007,N_15581,N_15286);
xnor U17008 (N_17008,N_14273,N_15923);
nand U17009 (N_17009,N_14798,N_15550);
or U17010 (N_17010,N_14628,N_14065);
nor U17011 (N_17011,N_14718,N_14257);
xor U17012 (N_17012,N_15670,N_14813);
or U17013 (N_17013,N_15330,N_14185);
or U17014 (N_17014,N_14002,N_15903);
nand U17015 (N_17015,N_15209,N_15000);
nor U17016 (N_17016,N_15495,N_15632);
or U17017 (N_17017,N_15203,N_14471);
or U17018 (N_17018,N_15292,N_14724);
or U17019 (N_17019,N_14962,N_14999);
xnor U17020 (N_17020,N_15707,N_14872);
nor U17021 (N_17021,N_14542,N_15042);
or U17022 (N_17022,N_14550,N_15717);
nor U17023 (N_17023,N_14359,N_15603);
nand U17024 (N_17024,N_14777,N_14919);
xnor U17025 (N_17025,N_15557,N_15513);
or U17026 (N_17026,N_14394,N_15067);
and U17027 (N_17027,N_14661,N_15691);
xor U17028 (N_17028,N_14142,N_14957);
or U17029 (N_17029,N_14317,N_14004);
nand U17030 (N_17030,N_15822,N_15782);
xnor U17031 (N_17031,N_15495,N_15652);
and U17032 (N_17032,N_15261,N_14343);
nor U17033 (N_17033,N_15314,N_15152);
nor U17034 (N_17034,N_15046,N_15465);
xnor U17035 (N_17035,N_15145,N_15450);
and U17036 (N_17036,N_14696,N_14412);
or U17037 (N_17037,N_15974,N_14360);
or U17038 (N_17038,N_14740,N_15809);
nor U17039 (N_17039,N_14691,N_15373);
xnor U17040 (N_17040,N_14379,N_14577);
or U17041 (N_17041,N_15167,N_14172);
nand U17042 (N_17042,N_15964,N_14465);
and U17043 (N_17043,N_14197,N_14274);
nand U17044 (N_17044,N_15778,N_15538);
and U17045 (N_17045,N_15446,N_15161);
nor U17046 (N_17046,N_14584,N_15213);
nor U17047 (N_17047,N_15012,N_14038);
or U17048 (N_17048,N_15716,N_15123);
or U17049 (N_17049,N_14915,N_14384);
and U17050 (N_17050,N_15463,N_15467);
and U17051 (N_17051,N_14961,N_15757);
nand U17052 (N_17052,N_15374,N_14152);
xnor U17053 (N_17053,N_15787,N_15325);
nor U17054 (N_17054,N_15035,N_15116);
nor U17055 (N_17055,N_14572,N_14336);
and U17056 (N_17056,N_15597,N_14117);
or U17057 (N_17057,N_15362,N_14155);
and U17058 (N_17058,N_15603,N_15028);
or U17059 (N_17059,N_15939,N_14779);
or U17060 (N_17060,N_14757,N_14743);
and U17061 (N_17061,N_14730,N_14625);
and U17062 (N_17062,N_15541,N_15827);
nor U17063 (N_17063,N_15417,N_14603);
nor U17064 (N_17064,N_15935,N_15049);
or U17065 (N_17065,N_15159,N_14834);
nand U17066 (N_17066,N_14917,N_15305);
and U17067 (N_17067,N_15191,N_14804);
nor U17068 (N_17068,N_15428,N_14946);
nor U17069 (N_17069,N_14960,N_15942);
nor U17070 (N_17070,N_14113,N_14239);
or U17071 (N_17071,N_14748,N_15292);
or U17072 (N_17072,N_15004,N_15979);
nor U17073 (N_17073,N_14170,N_14549);
nor U17074 (N_17074,N_15923,N_15438);
nand U17075 (N_17075,N_15124,N_14162);
xor U17076 (N_17076,N_15049,N_15044);
nand U17077 (N_17077,N_15809,N_15876);
or U17078 (N_17078,N_15402,N_14816);
nand U17079 (N_17079,N_15380,N_15552);
and U17080 (N_17080,N_15861,N_15369);
nor U17081 (N_17081,N_15947,N_15060);
nor U17082 (N_17082,N_14213,N_14968);
nor U17083 (N_17083,N_14641,N_15133);
nand U17084 (N_17084,N_15829,N_15090);
nand U17085 (N_17085,N_15118,N_14743);
or U17086 (N_17086,N_15968,N_14681);
nand U17087 (N_17087,N_15033,N_15694);
xor U17088 (N_17088,N_15796,N_15703);
nand U17089 (N_17089,N_15581,N_15893);
or U17090 (N_17090,N_14542,N_15383);
or U17091 (N_17091,N_15128,N_15322);
xnor U17092 (N_17092,N_15260,N_15928);
and U17093 (N_17093,N_14910,N_15374);
nand U17094 (N_17094,N_14964,N_15422);
or U17095 (N_17095,N_14315,N_15492);
nor U17096 (N_17096,N_15678,N_15919);
nand U17097 (N_17097,N_14952,N_15134);
and U17098 (N_17098,N_14068,N_14586);
or U17099 (N_17099,N_14549,N_15711);
xor U17100 (N_17100,N_15340,N_14210);
nand U17101 (N_17101,N_14257,N_15647);
nand U17102 (N_17102,N_15696,N_14872);
nand U17103 (N_17103,N_14616,N_14008);
and U17104 (N_17104,N_14564,N_14385);
nand U17105 (N_17105,N_15353,N_15265);
nor U17106 (N_17106,N_14658,N_14458);
nor U17107 (N_17107,N_14708,N_14605);
or U17108 (N_17108,N_14318,N_15167);
nor U17109 (N_17109,N_15453,N_14648);
nor U17110 (N_17110,N_14124,N_15918);
nor U17111 (N_17111,N_15817,N_14330);
xnor U17112 (N_17112,N_15663,N_14537);
xnor U17113 (N_17113,N_15615,N_14901);
nor U17114 (N_17114,N_14734,N_15077);
or U17115 (N_17115,N_15615,N_15154);
nand U17116 (N_17116,N_14830,N_14570);
or U17117 (N_17117,N_14166,N_14173);
nand U17118 (N_17118,N_14012,N_15944);
nand U17119 (N_17119,N_14956,N_14059);
nand U17120 (N_17120,N_15867,N_14788);
nor U17121 (N_17121,N_14750,N_15066);
xnor U17122 (N_17122,N_15229,N_14609);
and U17123 (N_17123,N_14418,N_14996);
nand U17124 (N_17124,N_15111,N_15803);
or U17125 (N_17125,N_14805,N_15383);
or U17126 (N_17126,N_15768,N_14030);
nor U17127 (N_17127,N_14078,N_15230);
and U17128 (N_17128,N_15194,N_14779);
or U17129 (N_17129,N_14207,N_14437);
nand U17130 (N_17130,N_14682,N_15485);
and U17131 (N_17131,N_14005,N_14880);
nand U17132 (N_17132,N_15060,N_14293);
xnor U17133 (N_17133,N_15431,N_15401);
nor U17134 (N_17134,N_15330,N_15947);
and U17135 (N_17135,N_15190,N_14273);
nor U17136 (N_17136,N_15360,N_14949);
nand U17137 (N_17137,N_15322,N_15261);
nand U17138 (N_17138,N_14271,N_15724);
nor U17139 (N_17139,N_14177,N_14345);
nor U17140 (N_17140,N_15851,N_15459);
nand U17141 (N_17141,N_14086,N_15637);
nand U17142 (N_17142,N_15130,N_15719);
nand U17143 (N_17143,N_15073,N_14257);
nor U17144 (N_17144,N_15033,N_14017);
nand U17145 (N_17145,N_14293,N_15844);
or U17146 (N_17146,N_14369,N_15434);
and U17147 (N_17147,N_15960,N_15513);
nor U17148 (N_17148,N_14416,N_15556);
nand U17149 (N_17149,N_15869,N_15087);
nor U17150 (N_17150,N_14862,N_15874);
and U17151 (N_17151,N_15262,N_14471);
or U17152 (N_17152,N_14768,N_15582);
or U17153 (N_17153,N_14499,N_14167);
or U17154 (N_17154,N_14392,N_14203);
nor U17155 (N_17155,N_15362,N_15147);
and U17156 (N_17156,N_15433,N_15670);
xnor U17157 (N_17157,N_14242,N_15746);
xnor U17158 (N_17158,N_14119,N_15086);
and U17159 (N_17159,N_14652,N_14410);
or U17160 (N_17160,N_15687,N_14803);
nand U17161 (N_17161,N_14864,N_15591);
xnor U17162 (N_17162,N_14996,N_15644);
xor U17163 (N_17163,N_15856,N_15531);
and U17164 (N_17164,N_15882,N_15088);
or U17165 (N_17165,N_14252,N_15556);
or U17166 (N_17166,N_15040,N_15046);
or U17167 (N_17167,N_14646,N_15074);
nand U17168 (N_17168,N_14657,N_14839);
and U17169 (N_17169,N_15907,N_14164);
nor U17170 (N_17170,N_14215,N_14053);
or U17171 (N_17171,N_14158,N_15868);
or U17172 (N_17172,N_15753,N_14245);
nor U17173 (N_17173,N_14629,N_15662);
and U17174 (N_17174,N_14659,N_14354);
or U17175 (N_17175,N_15808,N_14721);
or U17176 (N_17176,N_15357,N_14061);
and U17177 (N_17177,N_15666,N_15119);
or U17178 (N_17178,N_15013,N_14923);
nand U17179 (N_17179,N_15675,N_15610);
and U17180 (N_17180,N_14415,N_14346);
nand U17181 (N_17181,N_14068,N_14063);
and U17182 (N_17182,N_14113,N_15699);
and U17183 (N_17183,N_14366,N_14952);
and U17184 (N_17184,N_15322,N_14680);
and U17185 (N_17185,N_15327,N_15111);
xnor U17186 (N_17186,N_14059,N_15440);
nor U17187 (N_17187,N_15386,N_14941);
or U17188 (N_17188,N_15472,N_14426);
nor U17189 (N_17189,N_14408,N_14622);
nand U17190 (N_17190,N_15282,N_15829);
and U17191 (N_17191,N_15305,N_14242);
and U17192 (N_17192,N_15792,N_15997);
and U17193 (N_17193,N_15221,N_14500);
nor U17194 (N_17194,N_15279,N_14144);
and U17195 (N_17195,N_14385,N_15567);
nand U17196 (N_17196,N_15028,N_15419);
nor U17197 (N_17197,N_15249,N_15026);
nor U17198 (N_17198,N_15976,N_15072);
or U17199 (N_17199,N_14489,N_14123);
and U17200 (N_17200,N_15904,N_14857);
or U17201 (N_17201,N_15637,N_14621);
nor U17202 (N_17202,N_15814,N_14891);
nand U17203 (N_17203,N_15134,N_14614);
nor U17204 (N_17204,N_14973,N_15069);
and U17205 (N_17205,N_15222,N_14132);
and U17206 (N_17206,N_15478,N_14197);
and U17207 (N_17207,N_14776,N_14507);
and U17208 (N_17208,N_14725,N_14002);
and U17209 (N_17209,N_14921,N_14126);
or U17210 (N_17210,N_15024,N_14635);
xnor U17211 (N_17211,N_15135,N_15013);
and U17212 (N_17212,N_15658,N_15994);
nand U17213 (N_17213,N_15785,N_15368);
or U17214 (N_17214,N_14318,N_15740);
nand U17215 (N_17215,N_15122,N_15738);
nand U17216 (N_17216,N_14848,N_15561);
nand U17217 (N_17217,N_14208,N_15040);
and U17218 (N_17218,N_14672,N_14408);
and U17219 (N_17219,N_15773,N_15963);
nor U17220 (N_17220,N_15262,N_15141);
nor U17221 (N_17221,N_15818,N_15389);
nor U17222 (N_17222,N_14702,N_15160);
and U17223 (N_17223,N_15444,N_15151);
or U17224 (N_17224,N_14317,N_14849);
nand U17225 (N_17225,N_15656,N_14595);
nor U17226 (N_17226,N_14181,N_15365);
nor U17227 (N_17227,N_15618,N_15295);
nor U17228 (N_17228,N_15304,N_15835);
or U17229 (N_17229,N_14572,N_15395);
and U17230 (N_17230,N_15798,N_14808);
and U17231 (N_17231,N_15488,N_14697);
or U17232 (N_17232,N_14142,N_14981);
nand U17233 (N_17233,N_14587,N_14536);
or U17234 (N_17234,N_14331,N_14494);
nor U17235 (N_17235,N_14827,N_15883);
nand U17236 (N_17236,N_15245,N_15342);
and U17237 (N_17237,N_14556,N_14203);
and U17238 (N_17238,N_15129,N_15355);
and U17239 (N_17239,N_14017,N_14918);
and U17240 (N_17240,N_14763,N_15933);
nor U17241 (N_17241,N_15053,N_15961);
nand U17242 (N_17242,N_14312,N_15663);
or U17243 (N_17243,N_15091,N_15842);
nand U17244 (N_17244,N_15490,N_15824);
nor U17245 (N_17245,N_14690,N_14080);
nor U17246 (N_17246,N_14586,N_15577);
and U17247 (N_17247,N_15800,N_15690);
nor U17248 (N_17248,N_14754,N_14049);
nand U17249 (N_17249,N_14522,N_15699);
and U17250 (N_17250,N_15757,N_14517);
xnor U17251 (N_17251,N_15167,N_14865);
nor U17252 (N_17252,N_15692,N_14034);
and U17253 (N_17253,N_14371,N_15023);
nor U17254 (N_17254,N_14344,N_14999);
nand U17255 (N_17255,N_14307,N_15356);
or U17256 (N_17256,N_15234,N_14125);
and U17257 (N_17257,N_14046,N_15373);
nor U17258 (N_17258,N_15919,N_15283);
nor U17259 (N_17259,N_15841,N_14686);
nor U17260 (N_17260,N_15685,N_15488);
nand U17261 (N_17261,N_14809,N_15070);
nor U17262 (N_17262,N_14209,N_14325);
and U17263 (N_17263,N_14568,N_15281);
or U17264 (N_17264,N_15322,N_14703);
and U17265 (N_17265,N_14385,N_14593);
nor U17266 (N_17266,N_14860,N_14332);
xnor U17267 (N_17267,N_15733,N_15888);
or U17268 (N_17268,N_14810,N_14374);
or U17269 (N_17269,N_15236,N_14891);
xor U17270 (N_17270,N_14573,N_14177);
nand U17271 (N_17271,N_14885,N_15893);
nor U17272 (N_17272,N_15882,N_15723);
and U17273 (N_17273,N_15713,N_15478);
or U17274 (N_17274,N_15055,N_15968);
xnor U17275 (N_17275,N_15409,N_14296);
xnor U17276 (N_17276,N_15618,N_15837);
and U17277 (N_17277,N_14257,N_15011);
or U17278 (N_17278,N_14250,N_14108);
nand U17279 (N_17279,N_14158,N_15873);
nand U17280 (N_17280,N_15868,N_14092);
and U17281 (N_17281,N_15568,N_14242);
and U17282 (N_17282,N_14853,N_14052);
nor U17283 (N_17283,N_14717,N_15800);
and U17284 (N_17284,N_14916,N_14660);
nor U17285 (N_17285,N_15841,N_15498);
nor U17286 (N_17286,N_15804,N_15024);
or U17287 (N_17287,N_14794,N_14631);
or U17288 (N_17288,N_15074,N_15520);
or U17289 (N_17289,N_14135,N_15095);
and U17290 (N_17290,N_14393,N_14706);
and U17291 (N_17291,N_14757,N_15912);
or U17292 (N_17292,N_14784,N_15370);
and U17293 (N_17293,N_14216,N_15637);
nand U17294 (N_17294,N_14405,N_15099);
nor U17295 (N_17295,N_14139,N_14715);
or U17296 (N_17296,N_14843,N_15366);
and U17297 (N_17297,N_15834,N_15775);
or U17298 (N_17298,N_14417,N_14318);
and U17299 (N_17299,N_14812,N_15142);
nor U17300 (N_17300,N_15224,N_15958);
nor U17301 (N_17301,N_14050,N_14959);
nand U17302 (N_17302,N_14733,N_14224);
or U17303 (N_17303,N_14886,N_14974);
nor U17304 (N_17304,N_14230,N_14878);
nor U17305 (N_17305,N_15226,N_15900);
nand U17306 (N_17306,N_15347,N_15824);
or U17307 (N_17307,N_15922,N_15410);
or U17308 (N_17308,N_14796,N_15428);
and U17309 (N_17309,N_15711,N_15152);
or U17310 (N_17310,N_14900,N_14364);
and U17311 (N_17311,N_15083,N_14779);
and U17312 (N_17312,N_15287,N_15666);
nor U17313 (N_17313,N_15371,N_15993);
or U17314 (N_17314,N_15214,N_14025);
or U17315 (N_17315,N_14413,N_14598);
or U17316 (N_17316,N_14285,N_14205);
nand U17317 (N_17317,N_15408,N_14765);
nand U17318 (N_17318,N_14488,N_14138);
and U17319 (N_17319,N_14054,N_15733);
nand U17320 (N_17320,N_14382,N_14697);
xnor U17321 (N_17321,N_15748,N_15689);
nand U17322 (N_17322,N_14401,N_14472);
nand U17323 (N_17323,N_15688,N_14266);
and U17324 (N_17324,N_15584,N_14286);
xnor U17325 (N_17325,N_14056,N_15029);
and U17326 (N_17326,N_15261,N_15157);
and U17327 (N_17327,N_15423,N_14816);
or U17328 (N_17328,N_15101,N_14538);
nor U17329 (N_17329,N_14780,N_14012);
nor U17330 (N_17330,N_14580,N_14243);
and U17331 (N_17331,N_14177,N_15537);
nand U17332 (N_17332,N_15365,N_15235);
nor U17333 (N_17333,N_14558,N_14426);
and U17334 (N_17334,N_14639,N_15642);
and U17335 (N_17335,N_15801,N_14094);
nand U17336 (N_17336,N_15082,N_14100);
or U17337 (N_17337,N_14476,N_15504);
nand U17338 (N_17338,N_14713,N_15937);
and U17339 (N_17339,N_15528,N_15291);
or U17340 (N_17340,N_14504,N_15831);
nor U17341 (N_17341,N_14111,N_14291);
and U17342 (N_17342,N_14404,N_14874);
nor U17343 (N_17343,N_14653,N_15900);
nand U17344 (N_17344,N_15040,N_14943);
nand U17345 (N_17345,N_15958,N_15183);
and U17346 (N_17346,N_14390,N_15497);
nand U17347 (N_17347,N_14653,N_14495);
and U17348 (N_17348,N_15136,N_15660);
xor U17349 (N_17349,N_14887,N_14445);
nand U17350 (N_17350,N_15155,N_15245);
and U17351 (N_17351,N_15842,N_14993);
nor U17352 (N_17352,N_15364,N_15057);
and U17353 (N_17353,N_14398,N_14410);
nand U17354 (N_17354,N_14499,N_15246);
or U17355 (N_17355,N_14186,N_14626);
nand U17356 (N_17356,N_14099,N_14538);
nand U17357 (N_17357,N_15294,N_15491);
and U17358 (N_17358,N_14404,N_14670);
or U17359 (N_17359,N_14300,N_15774);
or U17360 (N_17360,N_14276,N_15419);
nor U17361 (N_17361,N_14373,N_14166);
nand U17362 (N_17362,N_14060,N_14539);
or U17363 (N_17363,N_14699,N_14440);
xor U17364 (N_17364,N_14885,N_15202);
nor U17365 (N_17365,N_15356,N_15059);
nand U17366 (N_17366,N_15061,N_14621);
nand U17367 (N_17367,N_15352,N_14037);
nor U17368 (N_17368,N_14176,N_15531);
and U17369 (N_17369,N_14343,N_14630);
nor U17370 (N_17370,N_15406,N_15766);
or U17371 (N_17371,N_14064,N_14291);
nor U17372 (N_17372,N_15733,N_15637);
nor U17373 (N_17373,N_15666,N_15774);
nor U17374 (N_17374,N_14887,N_15994);
and U17375 (N_17375,N_15036,N_14732);
nor U17376 (N_17376,N_14560,N_15830);
nand U17377 (N_17377,N_14094,N_14122);
nor U17378 (N_17378,N_14772,N_14811);
nor U17379 (N_17379,N_15045,N_14197);
and U17380 (N_17380,N_14308,N_15878);
and U17381 (N_17381,N_15964,N_15126);
xor U17382 (N_17382,N_14987,N_14725);
nor U17383 (N_17383,N_14615,N_15290);
and U17384 (N_17384,N_14517,N_14975);
or U17385 (N_17385,N_14774,N_14060);
or U17386 (N_17386,N_15968,N_15154);
nor U17387 (N_17387,N_14867,N_15829);
nor U17388 (N_17388,N_15969,N_15252);
xnor U17389 (N_17389,N_15504,N_14457);
xor U17390 (N_17390,N_14684,N_14766);
and U17391 (N_17391,N_15210,N_15490);
and U17392 (N_17392,N_14798,N_15482);
or U17393 (N_17393,N_15329,N_14726);
and U17394 (N_17394,N_15100,N_15030);
or U17395 (N_17395,N_15882,N_14013);
or U17396 (N_17396,N_14348,N_15024);
and U17397 (N_17397,N_14917,N_15011);
nor U17398 (N_17398,N_15247,N_15706);
nand U17399 (N_17399,N_14339,N_14845);
xor U17400 (N_17400,N_15590,N_15478);
nand U17401 (N_17401,N_15333,N_14379);
xnor U17402 (N_17402,N_15568,N_14267);
or U17403 (N_17403,N_14731,N_15090);
xor U17404 (N_17404,N_15500,N_14408);
or U17405 (N_17405,N_15248,N_14817);
and U17406 (N_17406,N_14907,N_14440);
and U17407 (N_17407,N_14965,N_14651);
or U17408 (N_17408,N_15178,N_14659);
nand U17409 (N_17409,N_14266,N_14029);
nand U17410 (N_17410,N_15505,N_14968);
nor U17411 (N_17411,N_14591,N_15867);
and U17412 (N_17412,N_15863,N_15893);
nand U17413 (N_17413,N_15084,N_15033);
and U17414 (N_17414,N_15242,N_14731);
xnor U17415 (N_17415,N_15116,N_15326);
or U17416 (N_17416,N_14963,N_14502);
nand U17417 (N_17417,N_14940,N_14034);
or U17418 (N_17418,N_14119,N_15025);
and U17419 (N_17419,N_15075,N_14368);
nand U17420 (N_17420,N_15024,N_14054);
nand U17421 (N_17421,N_14010,N_15305);
or U17422 (N_17422,N_14910,N_15985);
nor U17423 (N_17423,N_14299,N_14483);
nand U17424 (N_17424,N_14187,N_15472);
nor U17425 (N_17425,N_15509,N_15105);
nor U17426 (N_17426,N_14076,N_14520);
nor U17427 (N_17427,N_14524,N_15548);
nand U17428 (N_17428,N_15253,N_15587);
xor U17429 (N_17429,N_14394,N_15315);
nand U17430 (N_17430,N_14259,N_15809);
nand U17431 (N_17431,N_15876,N_15332);
xnor U17432 (N_17432,N_15536,N_14768);
and U17433 (N_17433,N_15121,N_15308);
and U17434 (N_17434,N_14146,N_15403);
xnor U17435 (N_17435,N_15832,N_15495);
nand U17436 (N_17436,N_15768,N_15660);
nor U17437 (N_17437,N_14551,N_14154);
or U17438 (N_17438,N_14427,N_15692);
or U17439 (N_17439,N_15715,N_14956);
and U17440 (N_17440,N_15496,N_14087);
and U17441 (N_17441,N_14942,N_14110);
nand U17442 (N_17442,N_14555,N_14081);
nor U17443 (N_17443,N_14315,N_14147);
xnor U17444 (N_17444,N_15947,N_14080);
and U17445 (N_17445,N_14414,N_15909);
nand U17446 (N_17446,N_14859,N_14096);
or U17447 (N_17447,N_15355,N_14066);
nor U17448 (N_17448,N_15439,N_14063);
nor U17449 (N_17449,N_14173,N_15288);
and U17450 (N_17450,N_14500,N_14694);
nor U17451 (N_17451,N_14085,N_14307);
nor U17452 (N_17452,N_15431,N_14668);
and U17453 (N_17453,N_15153,N_14164);
nand U17454 (N_17454,N_15607,N_15657);
nor U17455 (N_17455,N_15145,N_15413);
or U17456 (N_17456,N_14198,N_15667);
or U17457 (N_17457,N_15481,N_15168);
nor U17458 (N_17458,N_15156,N_15041);
and U17459 (N_17459,N_14230,N_14000);
xor U17460 (N_17460,N_15280,N_14216);
xnor U17461 (N_17461,N_15251,N_15761);
or U17462 (N_17462,N_14405,N_14656);
and U17463 (N_17463,N_15527,N_14446);
nand U17464 (N_17464,N_15194,N_14367);
and U17465 (N_17465,N_14104,N_15683);
or U17466 (N_17466,N_15588,N_15161);
nand U17467 (N_17467,N_15504,N_14242);
or U17468 (N_17468,N_15865,N_14440);
and U17469 (N_17469,N_14587,N_15922);
and U17470 (N_17470,N_15169,N_15874);
xnor U17471 (N_17471,N_15562,N_14700);
and U17472 (N_17472,N_15137,N_15178);
and U17473 (N_17473,N_15445,N_14524);
xnor U17474 (N_17474,N_14914,N_14932);
nand U17475 (N_17475,N_14478,N_15054);
xnor U17476 (N_17476,N_15764,N_15998);
xnor U17477 (N_17477,N_14489,N_15465);
and U17478 (N_17478,N_15646,N_15291);
xnor U17479 (N_17479,N_15004,N_14526);
and U17480 (N_17480,N_15148,N_14700);
nand U17481 (N_17481,N_15863,N_14259);
nand U17482 (N_17482,N_15501,N_14524);
nand U17483 (N_17483,N_14372,N_15449);
and U17484 (N_17484,N_14111,N_14589);
nor U17485 (N_17485,N_14813,N_15646);
or U17486 (N_17486,N_14961,N_14107);
nand U17487 (N_17487,N_14656,N_14787);
and U17488 (N_17488,N_15852,N_14824);
nand U17489 (N_17489,N_15420,N_14535);
nor U17490 (N_17490,N_15944,N_14602);
nand U17491 (N_17491,N_14516,N_14683);
xor U17492 (N_17492,N_14440,N_14484);
and U17493 (N_17493,N_14837,N_15635);
nand U17494 (N_17494,N_15928,N_15737);
or U17495 (N_17495,N_15362,N_14731);
and U17496 (N_17496,N_14209,N_14065);
xnor U17497 (N_17497,N_15399,N_15357);
nor U17498 (N_17498,N_14642,N_15191);
and U17499 (N_17499,N_15861,N_14384);
nand U17500 (N_17500,N_15051,N_15783);
nor U17501 (N_17501,N_14364,N_14877);
or U17502 (N_17502,N_14974,N_15015);
nand U17503 (N_17503,N_14230,N_15129);
nand U17504 (N_17504,N_15559,N_15783);
or U17505 (N_17505,N_14674,N_15295);
nor U17506 (N_17506,N_15836,N_15309);
or U17507 (N_17507,N_15024,N_15692);
nand U17508 (N_17508,N_14471,N_15645);
or U17509 (N_17509,N_14398,N_14826);
and U17510 (N_17510,N_14707,N_14107);
or U17511 (N_17511,N_15232,N_14330);
and U17512 (N_17512,N_15666,N_14059);
and U17513 (N_17513,N_14826,N_14376);
and U17514 (N_17514,N_15994,N_14998);
nor U17515 (N_17515,N_14911,N_14891);
or U17516 (N_17516,N_14104,N_15013);
nand U17517 (N_17517,N_15468,N_15109);
nor U17518 (N_17518,N_14012,N_15998);
xnor U17519 (N_17519,N_14225,N_14744);
and U17520 (N_17520,N_15360,N_14297);
and U17521 (N_17521,N_14666,N_14155);
nand U17522 (N_17522,N_14507,N_15590);
and U17523 (N_17523,N_14595,N_15942);
xnor U17524 (N_17524,N_15392,N_15054);
and U17525 (N_17525,N_15455,N_15746);
and U17526 (N_17526,N_14848,N_15805);
nor U17527 (N_17527,N_15009,N_15340);
nor U17528 (N_17528,N_14150,N_15359);
nor U17529 (N_17529,N_15634,N_15515);
or U17530 (N_17530,N_15516,N_14999);
nand U17531 (N_17531,N_15359,N_14719);
or U17532 (N_17532,N_15170,N_14582);
nand U17533 (N_17533,N_14448,N_14933);
nor U17534 (N_17534,N_15846,N_15082);
and U17535 (N_17535,N_15745,N_15914);
nor U17536 (N_17536,N_15171,N_14940);
nand U17537 (N_17537,N_15681,N_14868);
nand U17538 (N_17538,N_14338,N_15757);
nor U17539 (N_17539,N_15070,N_14561);
nor U17540 (N_17540,N_14882,N_15361);
nor U17541 (N_17541,N_14063,N_14219);
and U17542 (N_17542,N_14598,N_14950);
nand U17543 (N_17543,N_15893,N_14631);
xnor U17544 (N_17544,N_14147,N_14960);
or U17545 (N_17545,N_15613,N_15096);
and U17546 (N_17546,N_14829,N_14675);
nor U17547 (N_17547,N_15522,N_14937);
or U17548 (N_17548,N_15121,N_15958);
nand U17549 (N_17549,N_15015,N_14973);
xnor U17550 (N_17550,N_15469,N_14606);
xor U17551 (N_17551,N_14712,N_15155);
nor U17552 (N_17552,N_15630,N_15102);
and U17553 (N_17553,N_14347,N_14969);
or U17554 (N_17554,N_14576,N_15158);
xor U17555 (N_17555,N_15275,N_14478);
nand U17556 (N_17556,N_15368,N_14035);
and U17557 (N_17557,N_14549,N_15681);
nand U17558 (N_17558,N_15151,N_14964);
xor U17559 (N_17559,N_15371,N_14741);
or U17560 (N_17560,N_15283,N_15536);
nor U17561 (N_17561,N_15197,N_15914);
and U17562 (N_17562,N_14116,N_15358);
and U17563 (N_17563,N_14487,N_15283);
nand U17564 (N_17564,N_15812,N_15079);
nor U17565 (N_17565,N_14094,N_14113);
nand U17566 (N_17566,N_15330,N_15604);
nor U17567 (N_17567,N_14084,N_15310);
nand U17568 (N_17568,N_14183,N_14500);
nand U17569 (N_17569,N_15243,N_15503);
nor U17570 (N_17570,N_15225,N_15853);
xnor U17571 (N_17571,N_14738,N_15721);
nand U17572 (N_17572,N_15331,N_15732);
nand U17573 (N_17573,N_15885,N_14132);
nand U17574 (N_17574,N_15156,N_15741);
or U17575 (N_17575,N_15480,N_14908);
nand U17576 (N_17576,N_14298,N_15385);
and U17577 (N_17577,N_15147,N_14548);
or U17578 (N_17578,N_14436,N_15672);
or U17579 (N_17579,N_15399,N_14447);
nor U17580 (N_17580,N_14482,N_15177);
nor U17581 (N_17581,N_14225,N_14056);
nor U17582 (N_17582,N_15555,N_14482);
or U17583 (N_17583,N_15093,N_15042);
xnor U17584 (N_17584,N_15750,N_14607);
nor U17585 (N_17585,N_15990,N_15328);
and U17586 (N_17586,N_14080,N_14064);
nor U17587 (N_17587,N_15669,N_14403);
and U17588 (N_17588,N_14971,N_15327);
nand U17589 (N_17589,N_14526,N_14251);
xnor U17590 (N_17590,N_14293,N_15303);
or U17591 (N_17591,N_14483,N_15975);
and U17592 (N_17592,N_14813,N_14918);
nor U17593 (N_17593,N_15675,N_15799);
and U17594 (N_17594,N_14460,N_14782);
and U17595 (N_17595,N_15503,N_15420);
nor U17596 (N_17596,N_15618,N_15654);
and U17597 (N_17597,N_15742,N_14550);
nor U17598 (N_17598,N_14518,N_14468);
and U17599 (N_17599,N_15018,N_14809);
nand U17600 (N_17600,N_15054,N_15119);
xnor U17601 (N_17601,N_14082,N_14455);
and U17602 (N_17602,N_15864,N_14934);
or U17603 (N_17603,N_14150,N_15301);
nor U17604 (N_17604,N_15966,N_15237);
nand U17605 (N_17605,N_15358,N_15956);
or U17606 (N_17606,N_15475,N_15124);
and U17607 (N_17607,N_14928,N_15414);
or U17608 (N_17608,N_15378,N_14522);
nand U17609 (N_17609,N_15209,N_14303);
nand U17610 (N_17610,N_15813,N_14252);
nand U17611 (N_17611,N_15567,N_15931);
nor U17612 (N_17612,N_14105,N_14553);
and U17613 (N_17613,N_15910,N_15548);
or U17614 (N_17614,N_15615,N_15312);
or U17615 (N_17615,N_14994,N_14610);
and U17616 (N_17616,N_14780,N_15684);
and U17617 (N_17617,N_14889,N_15516);
xnor U17618 (N_17618,N_14026,N_15418);
xor U17619 (N_17619,N_14835,N_14270);
nor U17620 (N_17620,N_15475,N_14272);
or U17621 (N_17621,N_14549,N_15234);
and U17622 (N_17622,N_15466,N_14348);
and U17623 (N_17623,N_14049,N_14375);
nand U17624 (N_17624,N_14176,N_15692);
nor U17625 (N_17625,N_15784,N_14035);
xnor U17626 (N_17626,N_15952,N_15955);
or U17627 (N_17627,N_14830,N_14870);
xnor U17628 (N_17628,N_14052,N_15426);
or U17629 (N_17629,N_14929,N_15622);
and U17630 (N_17630,N_14286,N_15247);
and U17631 (N_17631,N_14008,N_15199);
xnor U17632 (N_17632,N_15250,N_14658);
nand U17633 (N_17633,N_15177,N_14798);
and U17634 (N_17634,N_14266,N_15860);
nor U17635 (N_17635,N_15688,N_14334);
nand U17636 (N_17636,N_14895,N_15117);
or U17637 (N_17637,N_14811,N_15515);
xor U17638 (N_17638,N_14022,N_14328);
nor U17639 (N_17639,N_15106,N_14577);
nand U17640 (N_17640,N_15507,N_14539);
nand U17641 (N_17641,N_14561,N_14746);
or U17642 (N_17642,N_15441,N_15237);
nor U17643 (N_17643,N_14995,N_15574);
nor U17644 (N_17644,N_15306,N_15038);
and U17645 (N_17645,N_14882,N_15339);
or U17646 (N_17646,N_14450,N_14556);
nor U17647 (N_17647,N_15623,N_14292);
and U17648 (N_17648,N_15294,N_15710);
nor U17649 (N_17649,N_14544,N_15323);
and U17650 (N_17650,N_15442,N_15106);
nand U17651 (N_17651,N_14968,N_15804);
and U17652 (N_17652,N_14754,N_15259);
or U17653 (N_17653,N_14167,N_15226);
and U17654 (N_17654,N_15464,N_14138);
nor U17655 (N_17655,N_15587,N_14220);
or U17656 (N_17656,N_15424,N_15869);
xnor U17657 (N_17657,N_15585,N_14777);
nor U17658 (N_17658,N_14893,N_15389);
nand U17659 (N_17659,N_15978,N_15590);
nor U17660 (N_17660,N_14329,N_14317);
or U17661 (N_17661,N_15132,N_14805);
and U17662 (N_17662,N_15189,N_15280);
nand U17663 (N_17663,N_15833,N_14461);
xnor U17664 (N_17664,N_14980,N_15974);
nor U17665 (N_17665,N_15492,N_15166);
and U17666 (N_17666,N_14735,N_15958);
and U17667 (N_17667,N_15468,N_14198);
nor U17668 (N_17668,N_15262,N_15395);
xnor U17669 (N_17669,N_15960,N_14247);
or U17670 (N_17670,N_14363,N_14434);
or U17671 (N_17671,N_15071,N_14186);
nand U17672 (N_17672,N_14753,N_15799);
xnor U17673 (N_17673,N_14837,N_15693);
nor U17674 (N_17674,N_15413,N_14227);
nand U17675 (N_17675,N_15810,N_14094);
nor U17676 (N_17676,N_14543,N_14237);
xor U17677 (N_17677,N_14221,N_15251);
nor U17678 (N_17678,N_14774,N_14935);
nor U17679 (N_17679,N_14884,N_15747);
xor U17680 (N_17680,N_15537,N_14309);
and U17681 (N_17681,N_15447,N_14122);
and U17682 (N_17682,N_15217,N_14322);
and U17683 (N_17683,N_14651,N_15008);
and U17684 (N_17684,N_14084,N_15212);
and U17685 (N_17685,N_15080,N_15036);
and U17686 (N_17686,N_15036,N_14569);
and U17687 (N_17687,N_14239,N_15910);
nor U17688 (N_17688,N_14475,N_15084);
nand U17689 (N_17689,N_14140,N_14344);
and U17690 (N_17690,N_15460,N_14495);
or U17691 (N_17691,N_15444,N_14901);
nand U17692 (N_17692,N_14458,N_15398);
xor U17693 (N_17693,N_15191,N_14973);
nand U17694 (N_17694,N_14090,N_14683);
or U17695 (N_17695,N_15866,N_14151);
nand U17696 (N_17696,N_14032,N_15097);
nand U17697 (N_17697,N_15194,N_15067);
and U17698 (N_17698,N_14029,N_14207);
and U17699 (N_17699,N_15469,N_14003);
and U17700 (N_17700,N_15338,N_15072);
nand U17701 (N_17701,N_14923,N_15179);
nor U17702 (N_17702,N_15919,N_14897);
or U17703 (N_17703,N_15836,N_15577);
and U17704 (N_17704,N_15227,N_14296);
and U17705 (N_17705,N_15537,N_15418);
nand U17706 (N_17706,N_15874,N_14574);
or U17707 (N_17707,N_15132,N_15264);
nand U17708 (N_17708,N_15866,N_15542);
or U17709 (N_17709,N_14134,N_14488);
xnor U17710 (N_17710,N_15564,N_15126);
and U17711 (N_17711,N_15850,N_15589);
or U17712 (N_17712,N_15398,N_14204);
and U17713 (N_17713,N_15095,N_15643);
nor U17714 (N_17714,N_15042,N_14059);
nor U17715 (N_17715,N_15862,N_14224);
or U17716 (N_17716,N_14728,N_14118);
nand U17717 (N_17717,N_14619,N_15335);
nor U17718 (N_17718,N_15062,N_14051);
or U17719 (N_17719,N_15390,N_14472);
and U17720 (N_17720,N_14523,N_15754);
or U17721 (N_17721,N_15344,N_15136);
and U17722 (N_17722,N_15415,N_15574);
xnor U17723 (N_17723,N_14073,N_15689);
xor U17724 (N_17724,N_15256,N_14081);
or U17725 (N_17725,N_14455,N_14431);
nand U17726 (N_17726,N_15196,N_15502);
nor U17727 (N_17727,N_14514,N_15679);
nor U17728 (N_17728,N_14930,N_15507);
or U17729 (N_17729,N_14696,N_15616);
nor U17730 (N_17730,N_14986,N_15813);
nand U17731 (N_17731,N_14752,N_14196);
or U17732 (N_17732,N_14808,N_15808);
nor U17733 (N_17733,N_14343,N_14534);
and U17734 (N_17734,N_15265,N_14102);
nor U17735 (N_17735,N_14469,N_14409);
nand U17736 (N_17736,N_14932,N_14895);
or U17737 (N_17737,N_14471,N_14296);
nand U17738 (N_17738,N_14305,N_15933);
nand U17739 (N_17739,N_14877,N_15504);
nor U17740 (N_17740,N_15004,N_14893);
or U17741 (N_17741,N_14934,N_15968);
and U17742 (N_17742,N_14608,N_14986);
and U17743 (N_17743,N_15069,N_15034);
nand U17744 (N_17744,N_15240,N_14417);
xnor U17745 (N_17745,N_14008,N_15429);
xor U17746 (N_17746,N_15305,N_15245);
or U17747 (N_17747,N_15785,N_15623);
and U17748 (N_17748,N_14606,N_15922);
or U17749 (N_17749,N_15741,N_15011);
xor U17750 (N_17750,N_15410,N_15270);
nand U17751 (N_17751,N_14260,N_15796);
xnor U17752 (N_17752,N_15901,N_15017);
and U17753 (N_17753,N_14905,N_15885);
nand U17754 (N_17754,N_14790,N_14105);
nand U17755 (N_17755,N_14176,N_14139);
nand U17756 (N_17756,N_15800,N_14068);
nand U17757 (N_17757,N_14785,N_14052);
and U17758 (N_17758,N_14181,N_14587);
nor U17759 (N_17759,N_15385,N_14586);
or U17760 (N_17760,N_15571,N_15406);
or U17761 (N_17761,N_14107,N_14302);
or U17762 (N_17762,N_14711,N_15142);
xor U17763 (N_17763,N_15675,N_15850);
and U17764 (N_17764,N_14639,N_15267);
nor U17765 (N_17765,N_14567,N_15990);
nor U17766 (N_17766,N_14682,N_14385);
and U17767 (N_17767,N_14157,N_14542);
or U17768 (N_17768,N_14231,N_14294);
or U17769 (N_17769,N_15968,N_14936);
nand U17770 (N_17770,N_15227,N_15375);
nand U17771 (N_17771,N_15511,N_14267);
nand U17772 (N_17772,N_15188,N_15656);
and U17773 (N_17773,N_15915,N_14119);
nand U17774 (N_17774,N_15152,N_14806);
nand U17775 (N_17775,N_15083,N_14363);
nand U17776 (N_17776,N_14374,N_14306);
and U17777 (N_17777,N_14936,N_14610);
nand U17778 (N_17778,N_14451,N_15278);
nand U17779 (N_17779,N_15924,N_15032);
or U17780 (N_17780,N_15811,N_14451);
nor U17781 (N_17781,N_15137,N_14089);
nand U17782 (N_17782,N_14975,N_15624);
nor U17783 (N_17783,N_15376,N_14756);
nor U17784 (N_17784,N_14656,N_15988);
and U17785 (N_17785,N_15379,N_15737);
and U17786 (N_17786,N_14401,N_15130);
nor U17787 (N_17787,N_15900,N_14068);
or U17788 (N_17788,N_15528,N_15774);
or U17789 (N_17789,N_15060,N_15047);
xnor U17790 (N_17790,N_15067,N_15639);
or U17791 (N_17791,N_15475,N_15044);
and U17792 (N_17792,N_14161,N_14606);
nand U17793 (N_17793,N_15626,N_14866);
nor U17794 (N_17794,N_14797,N_14208);
and U17795 (N_17795,N_14791,N_14884);
xnor U17796 (N_17796,N_14574,N_14969);
nand U17797 (N_17797,N_14770,N_14563);
or U17798 (N_17798,N_14514,N_15751);
or U17799 (N_17799,N_15430,N_15828);
or U17800 (N_17800,N_15078,N_15757);
xnor U17801 (N_17801,N_15178,N_14736);
nor U17802 (N_17802,N_15461,N_14977);
or U17803 (N_17803,N_15886,N_15964);
nor U17804 (N_17804,N_14333,N_14446);
nand U17805 (N_17805,N_15455,N_14102);
and U17806 (N_17806,N_15464,N_15426);
or U17807 (N_17807,N_15420,N_14616);
nor U17808 (N_17808,N_15737,N_14681);
nand U17809 (N_17809,N_14869,N_15383);
and U17810 (N_17810,N_14310,N_14152);
nand U17811 (N_17811,N_15784,N_15966);
nor U17812 (N_17812,N_15696,N_15670);
and U17813 (N_17813,N_14382,N_14102);
nor U17814 (N_17814,N_14606,N_15142);
and U17815 (N_17815,N_14330,N_14263);
or U17816 (N_17816,N_15382,N_15228);
nor U17817 (N_17817,N_15564,N_14222);
xnor U17818 (N_17818,N_14034,N_14283);
nor U17819 (N_17819,N_14636,N_14038);
or U17820 (N_17820,N_14431,N_14243);
and U17821 (N_17821,N_15131,N_15073);
and U17822 (N_17822,N_14373,N_15645);
nor U17823 (N_17823,N_14164,N_14092);
xor U17824 (N_17824,N_14998,N_14145);
nor U17825 (N_17825,N_14187,N_15654);
or U17826 (N_17826,N_15251,N_14915);
nand U17827 (N_17827,N_14436,N_14131);
and U17828 (N_17828,N_14336,N_15316);
nand U17829 (N_17829,N_14305,N_15214);
nand U17830 (N_17830,N_14968,N_15734);
nor U17831 (N_17831,N_15831,N_15027);
or U17832 (N_17832,N_14903,N_15688);
or U17833 (N_17833,N_14025,N_15507);
or U17834 (N_17834,N_14129,N_15496);
and U17835 (N_17835,N_15330,N_15166);
and U17836 (N_17836,N_14098,N_15132);
nand U17837 (N_17837,N_15377,N_14681);
nor U17838 (N_17838,N_14836,N_15303);
nor U17839 (N_17839,N_15790,N_15365);
or U17840 (N_17840,N_14114,N_15388);
and U17841 (N_17841,N_14682,N_14843);
and U17842 (N_17842,N_14923,N_15195);
nor U17843 (N_17843,N_15828,N_14746);
nor U17844 (N_17844,N_15045,N_14583);
nand U17845 (N_17845,N_14397,N_14676);
nand U17846 (N_17846,N_15754,N_15617);
nand U17847 (N_17847,N_14592,N_15780);
and U17848 (N_17848,N_14696,N_14467);
or U17849 (N_17849,N_14764,N_14538);
nand U17850 (N_17850,N_15999,N_14684);
and U17851 (N_17851,N_15531,N_14005);
and U17852 (N_17852,N_14656,N_14582);
or U17853 (N_17853,N_14002,N_15724);
nand U17854 (N_17854,N_14362,N_14445);
and U17855 (N_17855,N_14871,N_14131);
nand U17856 (N_17856,N_14190,N_15074);
nor U17857 (N_17857,N_15059,N_15451);
nand U17858 (N_17858,N_14792,N_15431);
and U17859 (N_17859,N_14305,N_14642);
nand U17860 (N_17860,N_15038,N_14050);
xnor U17861 (N_17861,N_14161,N_15819);
or U17862 (N_17862,N_14187,N_15423);
or U17863 (N_17863,N_14975,N_15039);
nand U17864 (N_17864,N_14372,N_14870);
and U17865 (N_17865,N_14765,N_14172);
nand U17866 (N_17866,N_15895,N_15410);
nand U17867 (N_17867,N_15953,N_15202);
xnor U17868 (N_17868,N_15038,N_14670);
and U17869 (N_17869,N_15793,N_14542);
nand U17870 (N_17870,N_15272,N_15885);
nand U17871 (N_17871,N_15519,N_14097);
nor U17872 (N_17872,N_15982,N_14704);
and U17873 (N_17873,N_14460,N_14822);
and U17874 (N_17874,N_15180,N_14515);
or U17875 (N_17875,N_14076,N_15228);
or U17876 (N_17876,N_14946,N_15891);
or U17877 (N_17877,N_14647,N_14200);
nand U17878 (N_17878,N_14297,N_15835);
nand U17879 (N_17879,N_15209,N_14706);
nand U17880 (N_17880,N_15970,N_14840);
nor U17881 (N_17881,N_14455,N_15881);
nand U17882 (N_17882,N_15839,N_14244);
nor U17883 (N_17883,N_15829,N_14751);
and U17884 (N_17884,N_14098,N_15589);
nor U17885 (N_17885,N_15151,N_15707);
or U17886 (N_17886,N_14514,N_14508);
or U17887 (N_17887,N_15729,N_15976);
or U17888 (N_17888,N_15993,N_14874);
xnor U17889 (N_17889,N_14646,N_14351);
nor U17890 (N_17890,N_14499,N_15488);
nand U17891 (N_17891,N_14876,N_15378);
and U17892 (N_17892,N_14795,N_15585);
nand U17893 (N_17893,N_14304,N_14558);
and U17894 (N_17894,N_14060,N_14619);
xor U17895 (N_17895,N_15055,N_15730);
or U17896 (N_17896,N_14428,N_15388);
nand U17897 (N_17897,N_15870,N_14128);
or U17898 (N_17898,N_15363,N_14245);
or U17899 (N_17899,N_15866,N_14361);
and U17900 (N_17900,N_14327,N_14554);
or U17901 (N_17901,N_14700,N_15564);
or U17902 (N_17902,N_14431,N_14118);
xor U17903 (N_17903,N_14192,N_15510);
or U17904 (N_17904,N_14601,N_14625);
nand U17905 (N_17905,N_15341,N_14943);
nor U17906 (N_17906,N_15656,N_15437);
and U17907 (N_17907,N_15069,N_14031);
nand U17908 (N_17908,N_14864,N_15606);
nand U17909 (N_17909,N_15473,N_15164);
and U17910 (N_17910,N_14820,N_14007);
nor U17911 (N_17911,N_15753,N_14206);
xor U17912 (N_17912,N_14192,N_14801);
nand U17913 (N_17913,N_14635,N_14560);
or U17914 (N_17914,N_14944,N_15590);
and U17915 (N_17915,N_14360,N_14765);
and U17916 (N_17916,N_15497,N_15676);
nand U17917 (N_17917,N_15356,N_14664);
or U17918 (N_17918,N_14381,N_14046);
nand U17919 (N_17919,N_15124,N_14507);
or U17920 (N_17920,N_14594,N_14312);
and U17921 (N_17921,N_14119,N_14619);
or U17922 (N_17922,N_14823,N_15275);
xnor U17923 (N_17923,N_14205,N_15636);
nor U17924 (N_17924,N_15516,N_14372);
xnor U17925 (N_17925,N_14871,N_14053);
and U17926 (N_17926,N_14489,N_14456);
or U17927 (N_17927,N_15838,N_15583);
xnor U17928 (N_17928,N_15884,N_15749);
and U17929 (N_17929,N_14272,N_15078);
nand U17930 (N_17930,N_15338,N_14932);
and U17931 (N_17931,N_15834,N_14076);
nor U17932 (N_17932,N_15924,N_14585);
or U17933 (N_17933,N_14454,N_14809);
or U17934 (N_17934,N_14393,N_15538);
or U17935 (N_17935,N_15882,N_14355);
nand U17936 (N_17936,N_14127,N_15206);
nor U17937 (N_17937,N_15053,N_14428);
and U17938 (N_17938,N_14794,N_15811);
and U17939 (N_17939,N_15830,N_15995);
or U17940 (N_17940,N_14953,N_14519);
nor U17941 (N_17941,N_15331,N_14222);
and U17942 (N_17942,N_14395,N_14417);
and U17943 (N_17943,N_15291,N_14927);
and U17944 (N_17944,N_15187,N_15304);
xnor U17945 (N_17945,N_15940,N_15955);
or U17946 (N_17946,N_15632,N_14731);
or U17947 (N_17947,N_14963,N_15470);
nand U17948 (N_17948,N_15122,N_14176);
nand U17949 (N_17949,N_14679,N_15859);
and U17950 (N_17950,N_14422,N_15154);
and U17951 (N_17951,N_14443,N_15896);
nor U17952 (N_17952,N_14014,N_15696);
nand U17953 (N_17953,N_15238,N_14392);
nor U17954 (N_17954,N_14489,N_14067);
nand U17955 (N_17955,N_14363,N_14673);
nor U17956 (N_17956,N_14254,N_15589);
nand U17957 (N_17957,N_14247,N_14728);
or U17958 (N_17958,N_15228,N_15942);
and U17959 (N_17959,N_15719,N_14909);
or U17960 (N_17960,N_15899,N_15508);
nor U17961 (N_17961,N_15686,N_15873);
and U17962 (N_17962,N_15345,N_15929);
nand U17963 (N_17963,N_15237,N_15503);
and U17964 (N_17964,N_15604,N_15446);
nor U17965 (N_17965,N_15909,N_14574);
or U17966 (N_17966,N_14773,N_14642);
or U17967 (N_17967,N_15030,N_14959);
xnor U17968 (N_17968,N_15952,N_15227);
or U17969 (N_17969,N_15020,N_14423);
nor U17970 (N_17970,N_14983,N_15979);
or U17971 (N_17971,N_14340,N_14183);
nand U17972 (N_17972,N_14864,N_14678);
nand U17973 (N_17973,N_15900,N_15366);
or U17974 (N_17974,N_14854,N_15289);
xor U17975 (N_17975,N_14286,N_14544);
and U17976 (N_17976,N_15522,N_15572);
nand U17977 (N_17977,N_15120,N_14144);
and U17978 (N_17978,N_15177,N_14320);
nand U17979 (N_17979,N_15289,N_15928);
and U17980 (N_17980,N_15126,N_15468);
xor U17981 (N_17981,N_14539,N_15861);
nor U17982 (N_17982,N_15269,N_14095);
nand U17983 (N_17983,N_15357,N_15968);
nand U17984 (N_17984,N_14429,N_14656);
nor U17985 (N_17985,N_14097,N_14608);
and U17986 (N_17986,N_14240,N_14753);
or U17987 (N_17987,N_15812,N_14854);
or U17988 (N_17988,N_15845,N_15920);
or U17989 (N_17989,N_15972,N_15183);
xnor U17990 (N_17990,N_15153,N_15647);
nor U17991 (N_17991,N_15920,N_14149);
and U17992 (N_17992,N_14017,N_14304);
nor U17993 (N_17993,N_15123,N_14466);
nand U17994 (N_17994,N_14748,N_14243);
nand U17995 (N_17995,N_15513,N_15607);
and U17996 (N_17996,N_15429,N_14626);
or U17997 (N_17997,N_14724,N_14013);
or U17998 (N_17998,N_14403,N_14415);
nor U17999 (N_17999,N_14946,N_14331);
nor U18000 (N_18000,N_17467,N_16433);
and U18001 (N_18001,N_17252,N_16525);
xnor U18002 (N_18002,N_16959,N_16415);
nand U18003 (N_18003,N_17801,N_16252);
and U18004 (N_18004,N_16444,N_17631);
nand U18005 (N_18005,N_16485,N_17530);
nor U18006 (N_18006,N_17385,N_17743);
xnor U18007 (N_18007,N_17687,N_16610);
and U18008 (N_18008,N_16777,N_16609);
nor U18009 (N_18009,N_17606,N_17830);
nand U18010 (N_18010,N_16545,N_16864);
or U18011 (N_18011,N_16233,N_16483);
or U18012 (N_18012,N_16672,N_17785);
nand U18013 (N_18013,N_16816,N_17675);
nand U18014 (N_18014,N_17454,N_17704);
and U18015 (N_18015,N_17726,N_17384);
and U18016 (N_18016,N_16073,N_17962);
nor U18017 (N_18017,N_17664,N_17236);
or U18018 (N_18018,N_17949,N_16400);
nor U18019 (N_18019,N_17635,N_17988);
or U18020 (N_18020,N_17678,N_17740);
nor U18021 (N_18021,N_17238,N_17413);
and U18022 (N_18022,N_16602,N_16068);
nand U18023 (N_18023,N_16318,N_16999);
xnor U18024 (N_18024,N_16008,N_16133);
nand U18025 (N_18025,N_16773,N_16786);
or U18026 (N_18026,N_16766,N_17973);
or U18027 (N_18027,N_16280,N_16847);
or U18028 (N_18028,N_17355,N_17322);
nand U18029 (N_18029,N_16587,N_17284);
nor U18030 (N_18030,N_17438,N_16467);
or U18031 (N_18031,N_17208,N_16599);
or U18032 (N_18032,N_17417,N_16331);
nand U18033 (N_18033,N_16244,N_16770);
or U18034 (N_18034,N_16633,N_17045);
nand U18035 (N_18035,N_17489,N_17897);
nor U18036 (N_18036,N_16995,N_17829);
nand U18037 (N_18037,N_16882,N_17207);
nand U18038 (N_18038,N_16040,N_16496);
nor U18039 (N_18039,N_16692,N_16705);
nand U18040 (N_18040,N_16982,N_17237);
nor U18041 (N_18041,N_16029,N_16978);
nand U18042 (N_18042,N_17856,N_16527);
or U18043 (N_18043,N_17433,N_17057);
and U18044 (N_18044,N_16071,N_16511);
xnor U18045 (N_18045,N_16498,N_17947);
xnor U18046 (N_18046,N_16658,N_17012);
nor U18047 (N_18047,N_16323,N_17182);
or U18048 (N_18048,N_16696,N_17789);
and U18049 (N_18049,N_17483,N_16649);
nand U18050 (N_18050,N_17734,N_16750);
nor U18051 (N_18051,N_17604,N_17472);
nor U18052 (N_18052,N_16870,N_17493);
and U18053 (N_18053,N_17071,N_17085);
or U18054 (N_18054,N_17172,N_16470);
nand U18055 (N_18055,N_16435,N_17531);
nand U18056 (N_18056,N_16583,N_16905);
or U18057 (N_18057,N_17439,N_17568);
nor U18058 (N_18058,N_16574,N_16184);
nand U18059 (N_18059,N_17721,N_17100);
or U18060 (N_18060,N_16768,N_17837);
or U18061 (N_18061,N_17533,N_16440);
nand U18062 (N_18062,N_16389,N_16034);
or U18063 (N_18063,N_17958,N_17637);
nor U18064 (N_18064,N_17692,N_16542);
and U18065 (N_18065,N_17399,N_16053);
or U18066 (N_18066,N_16550,N_16829);
nor U18067 (N_18067,N_17563,N_17333);
nor U18068 (N_18068,N_16675,N_17550);
nand U18069 (N_18069,N_17719,N_17266);
nor U18070 (N_18070,N_16226,N_17915);
and U18071 (N_18071,N_16501,N_16359);
nand U18072 (N_18072,N_17885,N_17598);
nand U18073 (N_18073,N_17034,N_16160);
nand U18074 (N_18074,N_17951,N_17326);
and U18075 (N_18075,N_16484,N_16432);
xnor U18076 (N_18076,N_17440,N_16590);
nor U18077 (N_18077,N_17123,N_16354);
or U18078 (N_18078,N_17392,N_17083);
and U18079 (N_18079,N_16579,N_17039);
nand U18080 (N_18080,N_16812,N_17044);
or U18081 (N_18081,N_16948,N_17360);
and U18082 (N_18082,N_17356,N_16411);
nor U18083 (N_18083,N_16544,N_16463);
and U18084 (N_18084,N_17193,N_16946);
or U18085 (N_18085,N_17168,N_17736);
or U18086 (N_18086,N_16756,N_16437);
and U18087 (N_18087,N_17338,N_17090);
nor U18088 (N_18088,N_17371,N_16606);
and U18089 (N_18089,N_16563,N_17127);
nor U18090 (N_18090,N_17735,N_16351);
nand U18091 (N_18091,N_16936,N_16297);
xnor U18092 (N_18092,N_17893,N_17633);
and U18093 (N_18093,N_16600,N_17321);
and U18094 (N_18094,N_16622,N_17254);
and U18095 (N_18095,N_17742,N_17724);
nor U18096 (N_18096,N_17184,N_17672);
nand U18097 (N_18097,N_17889,N_16255);
nor U18098 (N_18098,N_16837,N_16130);
nor U18099 (N_18099,N_17043,N_17288);
and U18100 (N_18100,N_16258,N_16871);
and U18101 (N_18101,N_17005,N_16186);
nand U18102 (N_18102,N_16933,N_16794);
nor U18103 (N_18103,N_16030,N_16753);
and U18104 (N_18104,N_16980,N_17854);
nand U18105 (N_18105,N_16701,N_16549);
or U18106 (N_18106,N_17777,N_16385);
nor U18107 (N_18107,N_16395,N_16124);
nand U18108 (N_18108,N_16059,N_16648);
or U18109 (N_18109,N_16589,N_16761);
and U18110 (N_18110,N_17283,N_17569);
xor U18111 (N_18111,N_17370,N_16222);
or U18112 (N_18112,N_16094,N_16854);
or U18113 (N_18113,N_16358,N_17747);
nand U18114 (N_18114,N_17708,N_16302);
nand U18115 (N_18115,N_17296,N_16971);
nor U18116 (N_18116,N_17901,N_17479);
and U18117 (N_18117,N_16588,N_16063);
and U18118 (N_18118,N_16047,N_16067);
or U18119 (N_18119,N_16977,N_17019);
xor U18120 (N_18120,N_17883,N_17394);
nor U18121 (N_18121,N_16779,N_16076);
nor U18122 (N_18122,N_16678,N_16253);
or U18123 (N_18123,N_17871,N_16451);
or U18124 (N_18124,N_17335,N_16056);
nor U18125 (N_18125,N_17778,N_17315);
nand U18126 (N_18126,N_16452,N_17122);
nand U18127 (N_18127,N_17359,N_16876);
and U18128 (N_18128,N_16901,N_16221);
and U18129 (N_18129,N_17106,N_16046);
xnor U18130 (N_18130,N_17874,N_16990);
nor U18131 (N_18131,N_16194,N_16249);
nand U18132 (N_18132,N_16725,N_16121);
nor U18133 (N_18133,N_17762,N_16548);
and U18134 (N_18134,N_16431,N_16401);
nor U18135 (N_18135,N_16507,N_16625);
or U18136 (N_18136,N_16667,N_16627);
nor U18137 (N_18137,N_16763,N_16007);
or U18138 (N_18138,N_16655,N_16394);
and U18139 (N_18139,N_17154,N_16185);
or U18140 (N_18140,N_17872,N_17389);
nand U18141 (N_18141,N_16099,N_17782);
nor U18142 (N_18142,N_16390,N_16552);
or U18143 (N_18143,N_16804,N_17485);
nand U18144 (N_18144,N_16917,N_17926);
xor U18145 (N_18145,N_16216,N_17727);
nand U18146 (N_18146,N_16488,N_16863);
and U18147 (N_18147,N_17764,N_16294);
and U18148 (N_18148,N_16897,N_17943);
nand U18149 (N_18149,N_17625,N_17132);
or U18150 (N_18150,N_16098,N_16232);
nor U18151 (N_18151,N_16833,N_16229);
nor U18152 (N_18152,N_16095,N_17136);
xor U18153 (N_18153,N_17999,N_17194);
and U18154 (N_18154,N_16708,N_17802);
and U18155 (N_18155,N_16145,N_17286);
and U18156 (N_18156,N_16840,N_17447);
and U18157 (N_18157,N_17673,N_16413);
nand U18158 (N_18158,N_17792,N_16754);
nor U18159 (N_18159,N_16581,N_17078);
nand U18160 (N_18160,N_17181,N_16962);
nand U18161 (N_18161,N_16744,N_16921);
nand U18162 (N_18162,N_17260,N_16427);
or U18163 (N_18163,N_16448,N_17310);
and U18164 (N_18164,N_16157,N_16514);
xnor U18165 (N_18165,N_16630,N_16953);
and U18166 (N_18166,N_16376,N_17632);
and U18167 (N_18167,N_16181,N_17676);
nand U18168 (N_18168,N_17639,N_17643);
nor U18169 (N_18169,N_16225,N_16814);
nand U18170 (N_18170,N_17804,N_16866);
nand U18171 (N_18171,N_17696,N_16717);
xor U18172 (N_18172,N_16577,N_17297);
nor U18173 (N_18173,N_16333,N_17537);
nand U18174 (N_18174,N_17161,N_16193);
or U18175 (N_18175,N_17173,N_16503);
nor U18176 (N_18176,N_17526,N_17985);
or U18177 (N_18177,N_17803,N_16805);
nor U18178 (N_18178,N_16096,N_17853);
nor U18179 (N_18179,N_17738,N_16139);
nor U18180 (N_18180,N_17822,N_17410);
or U18181 (N_18181,N_17574,N_16624);
or U18182 (N_18182,N_17120,N_16784);
and U18183 (N_18183,N_16582,N_17059);
or U18184 (N_18184,N_16983,N_17340);
nand U18185 (N_18185,N_16827,N_16832);
nor U18186 (N_18186,N_17810,N_17940);
nand U18187 (N_18187,N_17564,N_17027);
nor U18188 (N_18188,N_17124,N_16900);
and U18189 (N_18189,N_17709,N_17573);
nand U18190 (N_18190,N_16997,N_17627);
and U18191 (N_18191,N_16704,N_17102);
and U18192 (N_18192,N_16809,N_17066);
nor U18193 (N_18193,N_17987,N_17206);
xor U18194 (N_18194,N_17386,N_16557);
nor U18195 (N_18195,N_17784,N_16739);
nand U18196 (N_18196,N_16218,N_16656);
and U18197 (N_18197,N_16450,N_17797);
nand U18198 (N_18198,N_16453,N_16320);
and U18199 (N_18199,N_17199,N_17164);
nand U18200 (N_18200,N_16927,N_16154);
nand U18201 (N_18201,N_16994,N_17325);
and U18202 (N_18202,N_17904,N_16090);
or U18203 (N_18203,N_16706,N_16522);
or U18204 (N_18204,N_16815,N_16504);
and U18205 (N_18205,N_16668,N_16965);
or U18206 (N_18206,N_17244,N_17249);
and U18207 (N_18207,N_17151,N_17583);
and U18208 (N_18208,N_16623,N_17733);
xnor U18209 (N_18209,N_17409,N_17843);
nor U18210 (N_18210,N_16362,N_17587);
nor U18211 (N_18211,N_16074,N_16227);
or U18212 (N_18212,N_17271,N_16906);
and U18213 (N_18213,N_17428,N_17481);
nand U18214 (N_18214,N_17706,N_16884);
and U18215 (N_18215,N_17959,N_16165);
or U18216 (N_18216,N_17866,N_16373);
or U18217 (N_18217,N_17374,N_16004);
nand U18218 (N_18218,N_17349,N_17553);
and U18219 (N_18219,N_16263,N_17215);
or U18220 (N_18220,N_17524,N_17970);
nand U18221 (N_18221,N_16027,N_17556);
and U18222 (N_18222,N_16629,N_16239);
xnor U18223 (N_18223,N_17293,N_16170);
nor U18224 (N_18224,N_17723,N_17138);
nor U18225 (N_18225,N_17155,N_16443);
or U18226 (N_18226,N_17700,N_16019);
nand U18227 (N_18227,N_17307,N_17783);
or U18228 (N_18228,N_16638,N_17645);
and U18229 (N_18229,N_17536,N_17732);
and U18230 (N_18230,N_16474,N_17354);
nor U18231 (N_18231,N_16353,N_17836);
and U18232 (N_18232,N_16085,N_16825);
and U18233 (N_18233,N_16872,N_16778);
nand U18234 (N_18234,N_17174,N_17917);
and U18235 (N_18235,N_17697,N_16179);
nand U18236 (N_18236,N_16428,N_16892);
or U18237 (N_18237,N_17521,N_17179);
nand U18238 (N_18238,N_17010,N_17593);
or U18239 (N_18239,N_17660,N_17276);
nor U18240 (N_18240,N_17952,N_16920);
nand U18241 (N_18241,N_16259,N_17600);
and U18242 (N_18242,N_17757,N_16891);
and U18243 (N_18243,N_16989,N_16038);
nand U18244 (N_18244,N_17977,N_17093);
nand U18245 (N_18245,N_16231,N_17362);
nor U18246 (N_18246,N_16043,N_17111);
nor U18247 (N_18247,N_17157,N_16423);
nor U18248 (N_18248,N_17203,N_17220);
xnor U18249 (N_18249,N_16714,N_17539);
nor U18250 (N_18250,N_16486,N_17603);
xor U18251 (N_18251,N_17205,N_17147);
and U18252 (N_18252,N_17544,N_17729);
xnor U18253 (N_18253,N_16420,N_17329);
and U18254 (N_18254,N_17429,N_17135);
nand U18255 (N_18255,N_16340,N_16283);
nand U18256 (N_18256,N_17994,N_17101);
nor U18257 (N_18257,N_16643,N_17906);
nand U18258 (N_18258,N_16370,N_17636);
nor U18259 (N_18259,N_17806,N_16336);
and U18260 (N_18260,N_17444,N_16407);
nor U18261 (N_18261,N_16762,N_16277);
and U18262 (N_18262,N_16894,N_17975);
nor U18263 (N_18263,N_16585,N_16325);
nor U18264 (N_18264,N_16873,N_17339);
nor U18265 (N_18265,N_17759,N_17551);
nand U18266 (N_18266,N_17552,N_17163);
nand U18267 (N_18267,N_17300,N_16580);
nand U18268 (N_18268,N_17142,N_16841);
nor U18269 (N_18269,N_17016,N_17942);
or U18270 (N_18270,N_16908,N_16554);
nand U18271 (N_18271,N_16419,N_16970);
nand U18272 (N_18272,N_17169,N_17641);
nor U18273 (N_18273,N_17227,N_17056);
nand U18274 (N_18274,N_17980,N_17476);
nand U18275 (N_18275,N_17509,N_16541);
nor U18276 (N_18276,N_16939,N_17763);
and U18277 (N_18277,N_16080,N_17511);
nor U18278 (N_18278,N_16952,N_16724);
nor U18279 (N_18279,N_17838,N_16352);
or U18280 (N_18280,N_17013,N_17543);
xor U18281 (N_18281,N_17195,N_16693);
and U18282 (N_18282,N_17957,N_17277);
and U18283 (N_18283,N_17094,N_16149);
nor U18284 (N_18284,N_16575,N_16659);
nand U18285 (N_18285,N_17491,N_17855);
nor U18286 (N_18286,N_17525,N_16912);
nor U18287 (N_18287,N_17458,N_17150);
or U18288 (N_18288,N_16058,N_17542);
nor U18289 (N_18289,N_17964,N_17112);
and U18290 (N_18290,N_17914,N_17884);
nand U18291 (N_18291,N_17456,N_16381);
nor U18292 (N_18292,N_16048,N_17559);
and U18293 (N_18293,N_16597,N_16337);
nor U18294 (N_18294,N_16210,N_16663);
and U18295 (N_18295,N_16306,N_16572);
nand U18296 (N_18296,N_16640,N_16751);
nor U18297 (N_18297,N_17423,N_16887);
and U18298 (N_18298,N_17579,N_16288);
and U18299 (N_18299,N_17262,N_16788);
nor U18300 (N_18300,N_17756,N_17042);
nor U18301 (N_18301,N_16468,N_17597);
or U18302 (N_18302,N_16117,N_16935);
and U18303 (N_18303,N_17514,N_16309);
and U18304 (N_18304,N_16148,N_17594);
nand U18305 (N_18305,N_17047,N_17451);
and U18306 (N_18306,N_16310,N_17814);
nand U18307 (N_18307,N_16391,N_17891);
nand U18308 (N_18308,N_17176,N_16802);
or U18309 (N_18309,N_17912,N_17121);
and U18310 (N_18310,N_16881,N_16492);
and U18311 (N_18311,N_17412,N_16742);
and U18312 (N_18312,N_16964,N_17565);
nand U18313 (N_18313,N_17628,N_16520);
or U18314 (N_18314,N_17649,N_16430);
xor U18315 (N_18315,N_17946,N_17143);
nor U18316 (N_18316,N_17405,N_16016);
or U18317 (N_18317,N_17546,N_16931);
nor U18318 (N_18318,N_17555,N_17993);
or U18319 (N_18319,N_17484,N_16760);
or U18320 (N_18320,N_16457,N_17074);
nand U18321 (N_18321,N_17538,N_17812);
or U18322 (N_18322,N_16300,N_16162);
nor U18323 (N_18323,N_16902,N_16202);
xor U18324 (N_18324,N_16329,N_16533);
and U18325 (N_18325,N_16250,N_17463);
xor U18326 (N_18326,N_16026,N_16101);
nand U18327 (N_18327,N_17713,N_17584);
and U18328 (N_18328,N_16566,N_16114);
or U18329 (N_18329,N_16031,N_17372);
or U18330 (N_18330,N_17611,N_16267);
nor U18331 (N_18331,N_17768,N_17670);
xor U18332 (N_18332,N_17183,N_16679);
or U18333 (N_18333,N_16846,N_16772);
xor U18334 (N_18334,N_17684,N_16680);
and U18335 (N_18335,N_17907,N_17925);
or U18336 (N_18336,N_17613,N_16558);
nand U18337 (N_18337,N_17911,N_16199);
and U18338 (N_18338,N_16383,N_16543);
or U18339 (N_18339,N_16203,N_16562);
nand U18340 (N_18340,N_16726,N_16743);
and U18341 (N_18341,N_17629,N_17730);
nor U18342 (N_18342,N_17790,N_17879);
nor U18343 (N_18343,N_17069,N_17368);
nor U18344 (N_18344,N_17968,N_16850);
or U18345 (N_18345,N_16348,N_17092);
nor U18346 (N_18346,N_17818,N_17769);
nand U18347 (N_18347,N_16516,N_17459);
and U18348 (N_18348,N_17892,N_17848);
nand U18349 (N_18349,N_16112,N_16645);
nor U18350 (N_18350,N_17578,N_16746);
xor U18351 (N_18351,N_17400,N_17246);
nor U18352 (N_18352,N_17710,N_16228);
xnor U18353 (N_18353,N_17860,N_16619);
nand U18354 (N_18354,N_17001,N_16929);
or U18355 (N_18355,N_16111,N_17849);
nand U18356 (N_18356,N_16843,N_16561);
or U18357 (N_18357,N_17139,N_16050);
or U18358 (N_18358,N_16088,N_16918);
or U18359 (N_18359,N_17502,N_17327);
nor U18360 (N_18360,N_16108,N_17888);
and U18361 (N_18361,N_16867,N_17920);
or U18362 (N_18362,N_16044,N_17520);
or U18363 (N_18363,N_16895,N_17337);
xnor U18364 (N_18364,N_16510,N_16270);
nor U18365 (N_18365,N_16810,N_17470);
xor U18366 (N_18366,N_16072,N_16472);
xnor U18367 (N_18367,N_16342,N_16652);
or U18368 (N_18368,N_17041,N_16555);
or U18369 (N_18369,N_16538,N_16266);
xor U18370 (N_18370,N_16839,N_16269);
nor U18371 (N_18371,N_17928,N_17638);
or U18372 (N_18372,N_17406,N_16365);
nand U18373 (N_18373,N_17876,N_16276);
or U18374 (N_18374,N_16508,N_17712);
nor U18375 (N_18375,N_17334,N_17268);
or U18376 (N_18376,N_16289,N_16366);
or U18377 (N_18377,N_16321,N_16445);
or U18378 (N_18378,N_17863,N_17647);
nor U18379 (N_18379,N_17773,N_17937);
nand U18380 (N_18380,N_16404,N_17667);
nor U18381 (N_18381,N_16107,N_16860);
nor U18382 (N_18382,N_16398,N_17226);
or U18383 (N_18383,N_16106,N_17250);
and U18384 (N_18384,N_16618,N_17395);
or U18385 (N_18385,N_17365,N_17029);
and U18386 (N_18386,N_16967,N_17725);
and U18387 (N_18387,N_17351,N_17137);
and U18388 (N_18388,N_17414,N_17469);
nand U18389 (N_18389,N_16945,N_16326);
or U18390 (N_18390,N_17217,N_16776);
nor U18391 (N_18391,N_17835,N_17053);
xor U18392 (N_18392,N_17381,N_16402);
nor U18393 (N_18393,N_16120,N_16519);
or U18394 (N_18394,N_17075,N_17105);
nor U18395 (N_18395,N_17648,N_17634);
nor U18396 (N_18396,N_16922,N_17845);
nor U18397 (N_18397,N_16890,N_16877);
and U18398 (N_18398,N_17130,N_16204);
or U18399 (N_18399,N_17851,N_17323);
nor U18400 (N_18400,N_16314,N_16615);
xor U18401 (N_18401,N_16715,N_16426);
nand U18402 (N_18402,N_17180,N_17131);
and U18403 (N_18403,N_17930,N_17328);
or U18404 (N_18404,N_17082,N_17828);
nor U18405 (N_18405,N_17877,N_17366);
nand U18406 (N_18406,N_16368,N_16070);
or U18407 (N_18407,N_16338,N_17929);
or U18408 (N_18408,N_17443,N_16482);
and U18409 (N_18409,N_16175,N_16834);
xor U18410 (N_18410,N_16968,N_16273);
nand U18411 (N_18411,N_16916,N_17976);
nand U18412 (N_18412,N_17390,N_16925);
nor U18413 (N_18413,N_16205,N_17497);
nand U18414 (N_18414,N_16010,N_17997);
and U18415 (N_18415,N_16075,N_17982);
nor U18416 (N_18416,N_16360,N_16350);
and U18417 (N_18417,N_16690,N_16975);
and U18418 (N_18418,N_16764,N_16093);
and U18419 (N_18419,N_17701,N_16741);
or U18420 (N_18420,N_17809,N_16844);
xor U18421 (N_18421,N_17640,N_16898);
xnor U18422 (N_18422,N_17765,N_17022);
or U18423 (N_18423,N_16611,N_16178);
or U18424 (N_18424,N_17460,N_17677);
nor U18425 (N_18425,N_16686,N_16893);
and U18426 (N_18426,N_17817,N_17160);
or U18427 (N_18427,N_17890,N_16568);
or U18428 (N_18428,N_16985,N_16617);
nor U18429 (N_18429,N_16988,N_17963);
nor U18430 (N_18430,N_16196,N_16691);
nor U18431 (N_18431,N_16694,N_16189);
and U18432 (N_18432,N_16279,N_16045);
xnor U18433 (N_18433,N_16796,N_16003);
or U18434 (N_18434,N_17188,N_17508);
xor U18435 (N_18435,N_16459,N_16635);
and U18436 (N_18436,N_16681,N_17496);
and U18437 (N_18437,N_17654,N_16713);
nand U18438 (N_18438,N_16752,N_16261);
xnor U18439 (N_18439,N_16158,N_16446);
or U18440 (N_18440,N_17201,N_17050);
or U18441 (N_18441,N_17548,N_17465);
and U18442 (N_18442,N_17495,N_17886);
nor U18443 (N_18443,N_17210,N_16384);
or U18444 (N_18444,N_17519,N_17342);
nand U18445 (N_18445,N_16355,N_16116);
xor U18446 (N_18446,N_17055,N_16677);
nor U18447 (N_18447,N_16710,N_16981);
or U18448 (N_18448,N_16344,N_16238);
and U18449 (N_18449,N_16857,N_16291);
and U18450 (N_18450,N_16826,N_17916);
nor U18451 (N_18451,N_17619,N_17858);
and U18452 (N_18452,N_17245,N_17404);
or U18453 (N_18453,N_17791,N_17067);
nor U18454 (N_18454,N_16260,N_17223);
or U18455 (N_18455,N_17159,N_17504);
nor U18456 (N_18456,N_17718,N_16782);
and U18457 (N_18457,N_16002,N_17534);
nand U18458 (N_18458,N_17590,N_17623);
nor U18459 (N_18459,N_16209,N_17149);
nand U18460 (N_18460,N_17265,N_16792);
nor U18461 (N_18461,N_17477,N_17089);
or U18462 (N_18462,N_16128,N_16969);
or U18463 (N_18463,N_17774,N_17330);
and U18464 (N_18464,N_16268,N_16180);
nand U18465 (N_18465,N_17243,N_16497);
xor U18466 (N_18466,N_17566,N_17602);
xnor U18467 (N_18467,N_16246,N_16378);
and U18468 (N_18468,N_17331,N_17388);
and U18469 (N_18469,N_16438,N_16702);
or U18470 (N_18470,N_16041,N_17668);
xor U18471 (N_18471,N_17003,N_17343);
nor U18472 (N_18472,N_17024,N_16198);
nor U18473 (N_18473,N_17545,N_16439);
or U18474 (N_18474,N_16941,N_16405);
nand U18475 (N_18475,N_16214,N_16334);
or U18476 (N_18476,N_17974,N_16274);
nor U18477 (N_18477,N_17852,N_17680);
and U18478 (N_18478,N_16118,N_16565);
and U18479 (N_18479,N_16613,N_17948);
or U18480 (N_18480,N_16206,N_16220);
and U18481 (N_18481,N_17026,N_17475);
and U18482 (N_18482,N_17086,N_16992);
nor U18483 (N_18483,N_16505,N_16212);
nand U18484 (N_18484,N_17133,N_17786);
and U18485 (N_18485,N_16082,N_17017);
or U18486 (N_18486,N_16914,N_17189);
and U18487 (N_18487,N_17516,N_17685);
and U18488 (N_18488,N_17978,N_17666);
and U18489 (N_18489,N_17585,N_17811);
nor U18490 (N_18490,N_16547,N_17595);
or U18491 (N_18491,N_16343,N_17153);
nor U18492 (N_18492,N_16005,N_16998);
xnor U18493 (N_18493,N_17316,N_17880);
and U18494 (N_18494,N_17787,N_17054);
nor U18495 (N_18495,N_17224,N_16241);
nor U18496 (N_18496,N_16092,N_17760);
nand U18497 (N_18497,N_17607,N_16639);
or U18498 (N_18498,N_17927,N_17450);
nor U18499 (N_18499,N_17049,N_17287);
or U18500 (N_18500,N_16243,N_17900);
xor U18501 (N_18501,N_17767,N_17006);
or U18502 (N_18502,N_17332,N_17229);
nand U18503 (N_18503,N_17966,N_16765);
and U18504 (N_18504,N_17347,N_16907);
xnor U18505 (N_18505,N_17308,N_17312);
nand U18506 (N_18506,N_17267,N_16406);
or U18507 (N_18507,N_17945,N_16324);
nand U18508 (N_18508,N_16251,N_16529);
nor U18509 (N_18509,N_17617,N_17058);
and U18510 (N_18510,N_16163,N_16682);
nor U18511 (N_18511,N_17273,N_17609);
and U18512 (N_18512,N_16836,N_16614);
nand U18513 (N_18513,N_17644,N_17235);
nor U18514 (N_18514,N_16208,N_16396);
nor U18515 (N_18515,N_17198,N_16375);
nand U18516 (N_18516,N_16173,N_17256);
or U18517 (N_18517,N_16215,N_17936);
and U18518 (N_18518,N_17731,N_17068);
nor U18519 (N_18519,N_16584,N_17376);
or U18520 (N_18520,N_16595,N_17992);
or U18521 (N_18521,N_16661,N_17831);
and U18522 (N_18522,N_16831,N_17717);
nor U18523 (N_18523,N_16166,N_16966);
nand U18524 (N_18524,N_16471,N_17291);
nand U18525 (N_18525,N_16183,N_16055);
and U18526 (N_18526,N_17020,N_16357);
nor U18527 (N_18527,N_17186,N_16303);
nand U18528 (N_18528,N_16025,N_17522);
nand U18529 (N_18529,N_17748,N_16789);
or U18530 (N_18530,N_16033,N_17571);
nor U18531 (N_18531,N_16626,N_17052);
or U18532 (N_18532,N_17302,N_17166);
nand U18533 (N_18533,N_17861,N_17486);
or U18534 (N_18534,N_17560,N_17847);
or U18535 (N_18535,N_16716,N_16409);
nor U18536 (N_18536,N_16201,N_17040);
xor U18537 (N_18537,N_17499,N_17490);
xnor U18538 (N_18538,N_17228,N_16122);
or U18539 (N_18539,N_17191,N_16188);
nor U18540 (N_18540,N_17025,N_16849);
nor U18541 (N_18541,N_17346,N_16113);
nand U18542 (N_18542,N_17558,N_16697);
nor U18543 (N_18543,N_17088,N_17218);
or U18544 (N_18544,N_17113,N_17253);
nor U18545 (N_18545,N_16245,N_16475);
nand U18546 (N_18546,N_16732,N_16254);
and U18547 (N_18547,N_16851,N_17209);
and U18548 (N_18548,N_17715,N_16880);
or U18549 (N_18549,N_17918,N_17577);
and U18550 (N_18550,N_17589,N_17826);
xnor U18551 (N_18551,N_17141,N_17233);
and U18552 (N_18552,N_17859,N_17699);
nor U18553 (N_18553,N_16213,N_17682);
or U18554 (N_18554,N_16769,N_17705);
or U18555 (N_18555,N_16436,N_16512);
and U18556 (N_18556,N_17722,N_17698);
nand U18557 (N_18557,N_16926,N_16069);
or U18558 (N_18558,N_17369,N_17028);
or U18559 (N_18559,N_16421,N_17931);
nand U18560 (N_18560,N_17995,N_16687);
or U18561 (N_18561,N_17320,N_16379);
nand U18562 (N_18562,N_16319,N_16028);
and U18563 (N_18563,N_17819,N_17562);
and U18564 (N_18564,N_17015,N_16888);
and U18565 (N_18565,N_17391,N_17313);
nand U18566 (N_18566,N_16377,N_17294);
nand U18567 (N_18567,N_16822,N_17115);
and U18568 (N_18568,N_16006,N_17196);
nor U18569 (N_18569,N_17510,N_16703);
and U18570 (N_18570,N_17857,N_17527);
nand U18571 (N_18571,N_16593,N_16883);
nor U18572 (N_18572,N_16911,N_17116);
and U18573 (N_18573,N_16086,N_16608);
xor U18574 (N_18574,N_17905,N_16553);
nand U18575 (N_18575,N_16190,N_17983);
and U18576 (N_18576,N_17239,N_17221);
or U18577 (N_18577,N_16418,N_16560);
or U18578 (N_18578,N_17367,N_16944);
xor U18579 (N_18579,N_17834,N_16885);
or U18580 (N_18580,N_17816,N_16177);
nand U18581 (N_18581,N_16958,N_17398);
and U18582 (N_18582,N_17998,N_16248);
and U18583 (N_18583,N_16830,N_16119);
nand U18584 (N_18584,N_16546,N_16748);
nand U18585 (N_18585,N_16151,N_17110);
nor U18586 (N_18586,N_16479,N_16060);
and U18587 (N_18587,N_17924,N_16960);
or U18588 (N_18588,N_16509,N_16570);
nor U18589 (N_18589,N_16996,N_16862);
nand U18590 (N_18590,N_16084,N_17187);
nand U18591 (N_18591,N_17798,N_16878);
xor U18592 (N_18592,N_17941,N_17986);
nand U18593 (N_18593,N_16603,N_17990);
or U18594 (N_18594,N_17776,N_16530);
nor U18595 (N_18595,N_16612,N_17832);
nand U18596 (N_18596,N_16528,N_17301);
or U18597 (N_18597,N_17842,N_16757);
and U18598 (N_18598,N_17263,N_16211);
nor U18599 (N_18599,N_16144,N_16087);
nand U18600 (N_18600,N_16089,N_16904);
and U18601 (N_18601,N_17018,N_16292);
nor U18602 (N_18602,N_17653,N_16012);
nand U18603 (N_18603,N_17062,N_16293);
or U18604 (N_18604,N_16035,N_17601);
nand U18605 (N_18605,N_16097,N_17383);
nor U18606 (N_18606,N_17661,N_17944);
nand U18607 (N_18607,N_17387,N_16657);
and U18608 (N_18608,N_17379,N_17167);
nor U18609 (N_18609,N_16408,N_17934);
or U18610 (N_18610,N_16287,N_16388);
nor U18611 (N_18611,N_17211,N_16078);
and U18612 (N_18612,N_17908,N_16416);
or U18613 (N_18613,N_16410,N_16125);
nor U18614 (N_18614,N_16596,N_16749);
and U18615 (N_18615,N_17532,N_17036);
nand U18616 (N_18616,N_17422,N_17482);
xor U18617 (N_18617,N_16755,N_16707);
or U18618 (N_18618,N_16709,N_17658);
nand U18619 (N_18619,N_16349,N_16730);
or U18620 (N_18620,N_16057,N_16791);
or U18621 (N_18621,N_17165,N_16955);
and U18622 (N_18622,N_17506,N_17431);
or U18623 (N_18623,N_16081,N_17753);
nand U18624 (N_18624,N_16367,N_17471);
and U18625 (N_18625,N_16984,N_16110);
nor U18626 (N_18626,N_17204,N_17932);
or U18627 (N_18627,N_16874,N_17197);
nor U18628 (N_18628,N_17796,N_16335);
nor U18629 (N_18629,N_17575,N_16875);
or U18630 (N_18630,N_16676,N_16718);
nor U18631 (N_18631,N_17669,N_17004);
nand U18632 (N_18632,N_17126,N_17494);
and U18633 (N_18633,N_16372,N_16032);
and U18634 (N_18634,N_17586,N_17453);
or U18635 (N_18635,N_16973,N_16062);
and U18636 (N_18636,N_16976,N_17011);
and U18637 (N_18637,N_16065,N_16654);
nor U18638 (N_18638,N_16793,N_17171);
and U18639 (N_18639,N_17570,N_17505);
nor U18640 (N_18640,N_16685,N_16631);
xor U18641 (N_18641,N_17939,N_16064);
nor U18642 (N_18642,N_16799,N_17382);
or U18643 (N_18643,N_16466,N_16140);
nand U18644 (N_18644,N_16771,N_17192);
or U18645 (N_18645,N_17114,N_16734);
nand U18646 (N_18646,N_16156,N_17060);
and U18647 (N_18647,N_17077,N_17938);
xor U18648 (N_18648,N_16729,N_16738);
nor U18649 (N_18649,N_16759,N_16924);
nand U18650 (N_18650,N_16785,N_17008);
nand U18651 (N_18651,N_17305,N_16780);
nor U18652 (N_18652,N_16535,N_17626);
and U18653 (N_18653,N_17345,N_16465);
nand U18654 (N_18654,N_16131,N_17878);
and U18655 (N_18655,N_16733,N_17823);
or U18656 (N_18656,N_16666,N_16928);
nor U18657 (N_18657,N_16434,N_17689);
and U18658 (N_18658,N_16961,N_16899);
nor U18659 (N_18659,N_16022,N_16172);
or U18660 (N_18660,N_16559,N_17108);
nand U18661 (N_18661,N_16299,N_16795);
nand U18662 (N_18662,N_17984,N_16695);
or U18663 (N_18663,N_17825,N_17190);
xnor U18664 (N_18664,N_16700,N_16774);
and U18665 (N_18665,N_16282,N_17259);
nor U18666 (N_18666,N_16257,N_17251);
and U18667 (N_18667,N_17933,N_16013);
nand U18668 (N_18668,N_16747,N_17989);
nor U18669 (N_18669,N_16569,N_17841);
or U18670 (N_18670,N_17624,N_17616);
and U18671 (N_18671,N_16515,N_17278);
nor U18672 (N_18672,N_17591,N_17178);
or U18673 (N_18673,N_16767,N_16937);
or U18674 (N_18674,N_16842,N_17037);
nor U18675 (N_18675,N_17257,N_17258);
xor U18676 (N_18676,N_16499,N_17032);
or U18677 (N_18677,N_17352,N_16731);
nand U18678 (N_18678,N_16374,N_17754);
or U18679 (N_18679,N_16711,N_16195);
nor U18680 (N_18680,N_16200,N_16102);
nand U18681 (N_18681,N_16477,N_17474);
or U18682 (N_18682,N_16576,N_17899);
or U18683 (N_18683,N_17683,N_17702);
or U18684 (N_18684,N_16020,N_16858);
xnor U18685 (N_18685,N_16942,N_16489);
xor U18686 (N_18686,N_16422,N_17850);
nor U18687 (N_18687,N_17214,N_16403);
or U18688 (N_18688,N_16536,N_17377);
nor U18689 (N_18689,N_17073,N_17681);
nand U18690 (N_18690,N_17350,N_17038);
or U18691 (N_18691,N_16000,N_17292);
or U18692 (N_18692,N_17839,N_16049);
and U18693 (N_18693,N_17314,N_16821);
and U18694 (N_18694,N_16913,N_16230);
xnor U18695 (N_18695,N_17441,N_17547);
nand U18696 (N_18696,N_16182,N_16736);
xor U18697 (N_18697,N_16387,N_16651);
or U18698 (N_18698,N_16147,N_16517);
or U18699 (N_18699,N_17231,N_16015);
nor U18700 (N_18700,N_16290,N_17076);
nand U18701 (N_18701,N_16219,N_17270);
nand U18702 (N_18702,N_17299,N_17580);
nor U18703 (N_18703,N_17107,N_16819);
and U18704 (N_18704,N_17739,N_17679);
nand U18705 (N_18705,N_16594,N_17833);
nor U18706 (N_18706,N_16910,N_16264);
and U18707 (N_18707,N_17674,N_16328);
or U18708 (N_18708,N_17411,N_16856);
or U18709 (N_18709,N_17225,N_17622);
xor U18710 (N_18710,N_17408,N_17275);
xnor U18711 (N_18711,N_16932,N_17222);
nor U18712 (N_18712,N_17662,N_17303);
and U18713 (N_18713,N_17466,N_17554);
or U18714 (N_18714,N_16478,N_16628);
and U18715 (N_18715,N_16153,N_17344);
nor U18716 (N_18716,N_17129,N_17247);
or U18717 (N_18717,N_16393,N_16146);
or U18718 (N_18718,N_17185,N_16284);
nand U18719 (N_18719,N_16449,N_16604);
and U18720 (N_18720,N_16458,N_17758);
and U18721 (N_18721,N_16721,N_16083);
nand U18722 (N_18722,N_17448,N_16424);
or U18723 (N_18723,N_17030,N_17894);
and U18724 (N_18724,N_16103,N_17118);
and U18725 (N_18725,N_16425,N_17761);
and U18726 (N_18726,N_16513,N_17824);
nand U18727 (N_18727,N_16524,N_16644);
nor U18728 (N_18728,N_16295,N_16462);
nand U18729 (N_18729,N_17541,N_17099);
or U18730 (N_18730,N_16647,N_16115);
nand U18731 (N_18731,N_16024,N_17960);
and U18732 (N_18732,N_16235,N_17087);
or U18733 (N_18733,N_17200,N_16311);
xor U18734 (N_18734,N_17535,N_17844);
and U18735 (N_18735,N_17426,N_16852);
and U18736 (N_18736,N_16143,N_16142);
and U18737 (N_18737,N_16991,N_17864);
and U18738 (N_18738,N_16502,N_17478);
nand U18739 (N_18739,N_17419,N_16735);
or U18740 (N_18740,N_16564,N_16813);
nor U18741 (N_18741,N_17140,N_16313);
and U18742 (N_18742,N_16859,N_16129);
and U18743 (N_18743,N_17002,N_16781);
or U18744 (N_18744,N_17457,N_17396);
nand U18745 (N_18745,N_17714,N_17280);
nor U18746 (N_18746,N_17358,N_17128);
or U18747 (N_18747,N_17771,N_17353);
or U18748 (N_18748,N_16669,N_17436);
or U18749 (N_18749,N_16972,N_16168);
or U18750 (N_18750,N_17630,N_16934);
and U18751 (N_18751,N_16371,N_16152);
or U18752 (N_18752,N_16957,N_17576);
xnor U18753 (N_18753,N_17896,N_16494);
or U18754 (N_18754,N_17146,N_17744);
nor U18755 (N_18755,N_16414,N_17415);
nor U18756 (N_18756,N_16109,N_16493);
and U18757 (N_18757,N_17903,N_16347);
and U18758 (N_18758,N_16345,N_16473);
or U18759 (N_18759,N_16174,N_16281);
and U18760 (N_18760,N_16018,N_17290);
or U18761 (N_18761,N_17498,N_16077);
nand U18762 (N_18762,N_17750,N_16417);
xor U18763 (N_18763,N_16828,N_17961);
or U18764 (N_18764,N_16327,N_17656);
nor U18765 (N_18765,N_17234,N_16469);
xor U18766 (N_18766,N_16683,N_16664);
xor U18767 (N_18767,N_17655,N_16823);
xor U18768 (N_18768,N_17881,N_16316);
nor U18769 (N_18769,N_17781,N_16476);
or U18770 (N_18770,N_16464,N_17703);
or U18771 (N_18771,N_17909,N_17051);
nand U18772 (N_18772,N_17954,N_17882);
nand U18773 (N_18773,N_16356,N_17652);
nor U18774 (N_18774,N_16341,N_16317);
nor U18775 (N_18775,N_16531,N_17503);
and U18776 (N_18776,N_16369,N_16460);
and U18777 (N_18777,N_16919,N_17979);
or U18778 (N_18778,N_17695,N_17870);
nand U18779 (N_18779,N_17033,N_17540);
xor U18780 (N_18780,N_16775,N_16286);
nand U18781 (N_18781,N_16551,N_17035);
or U18782 (N_18782,N_16506,N_17523);
nor U18783 (N_18783,N_17775,N_17561);
nand U18784 (N_18784,N_17202,N_16688);
or U18785 (N_18785,N_16386,N_16207);
nor U18786 (N_18786,N_17298,N_17427);
nor U18787 (N_18787,N_16061,N_16521);
or U18788 (N_18788,N_17375,N_16155);
and U18789 (N_18789,N_16567,N_16650);
nor U18790 (N_18790,N_16066,N_17728);
or U18791 (N_18791,N_16540,N_16674);
nand U18792 (N_18792,N_17445,N_17079);
nor U18793 (N_18793,N_17464,N_17592);
nand U18794 (N_18794,N_16879,N_16171);
nand U18795 (N_18795,N_17996,N_17808);
or U18796 (N_18796,N_16855,N_16301);
nor U18797 (N_18797,N_17119,N_16673);
nand U18798 (N_18798,N_17373,N_17935);
and U18799 (N_18799,N_16023,N_17827);
nand U18800 (N_18800,N_17690,N_17862);
nand U18801 (N_18801,N_16001,N_16720);
nor U18802 (N_18802,N_17021,N_17642);
or U18803 (N_18803,N_16526,N_17755);
nor U18804 (N_18804,N_17156,N_17711);
nand U18805 (N_18805,N_17588,N_17418);
and U18806 (N_18806,N_16322,N_16036);
nor U18807 (N_18807,N_17401,N_17452);
nand U18808 (N_18808,N_17965,N_16938);
nand U18809 (N_18809,N_17425,N_16454);
xnor U18810 (N_18810,N_17795,N_17449);
or U18811 (N_18811,N_17407,N_16429);
or U18812 (N_18812,N_17091,N_17061);
or U18813 (N_18813,N_16456,N_16632);
and U18814 (N_18814,N_16480,N_16719);
nor U18815 (N_18815,N_16330,N_17615);
nor U18816 (N_18816,N_17746,N_17096);
nor U18817 (N_18817,N_17869,N_16265);
nor U18818 (N_18818,N_16132,N_17610);
or U18819 (N_18819,N_17317,N_17612);
and U18820 (N_18820,N_17364,N_17513);
nand U18821 (N_18821,N_17549,N_17581);
xnor U18822 (N_18822,N_16712,N_16797);
xor U18823 (N_18823,N_17688,N_16954);
and U18824 (N_18824,N_16865,N_17380);
nand U18825 (N_18825,N_17922,N_17152);
nand U18826 (N_18826,N_17693,N_16915);
and U18827 (N_18827,N_17799,N_17492);
nand U18828 (N_18828,N_17023,N_16308);
nor U18829 (N_18829,N_16646,N_16262);
and U18830 (N_18830,N_16950,N_16399);
xor U18831 (N_18831,N_17887,N_17311);
or U18832 (N_18832,N_16167,N_16021);
nand U18833 (N_18833,N_16382,N_16943);
xor U18834 (N_18834,N_16491,N_16346);
nor U18835 (N_18835,N_16137,N_16141);
nand U18836 (N_18836,N_16304,N_17772);
or U18837 (N_18837,N_16490,N_16660);
or U18838 (N_18838,N_17324,N_16296);
or U18839 (N_18839,N_17517,N_17745);
or U18840 (N_18840,N_17752,N_17000);
nand U18841 (N_18841,N_16192,N_16820);
nand U18842 (N_18842,N_17582,N_16312);
nor U18843 (N_18843,N_16234,N_16237);
or U18844 (N_18844,N_16392,N_16271);
xor U18845 (N_18845,N_17065,N_16363);
or U18846 (N_18846,N_16256,N_17432);
xnor U18847 (N_18847,N_17898,N_17357);
and U18848 (N_18848,N_17650,N_17274);
or U18849 (N_18849,N_17109,N_17219);
nor U18850 (N_18850,N_16723,N_16105);
or U18851 (N_18851,N_16079,N_17424);
nor U18852 (N_18852,N_16798,N_17014);
nor U18853 (N_18853,N_17403,N_16930);
and U18854 (N_18854,N_17095,N_17104);
nor U18855 (N_18855,N_17304,N_16787);
nor U18856 (N_18856,N_16240,N_16412);
xnor U18857 (N_18857,N_17865,N_17397);
nand U18858 (N_18858,N_16665,N_17815);
and U18859 (N_18859,N_17981,N_17420);
nand U18860 (N_18860,N_17518,N_16191);
nor U18861 (N_18861,N_17255,N_17318);
nand U18862 (N_18862,N_17269,N_17950);
or U18863 (N_18863,N_17605,N_16790);
nand U18864 (N_18864,N_17780,N_16949);
and U18865 (N_18865,N_17991,N_17820);
and U18866 (N_18866,N_17261,N_17098);
or U18867 (N_18867,N_16903,N_17468);
nand U18868 (N_18868,N_16727,N_17868);
nor U18869 (N_18869,N_16495,N_16305);
or U18870 (N_18870,N_16993,N_17162);
and U18871 (N_18871,N_17117,N_16698);
nor U18872 (N_18872,N_16285,N_17435);
xnor U18873 (N_18873,N_17272,N_16889);
xnor U18874 (N_18874,N_17800,N_17840);
nand U18875 (N_18875,N_16699,N_16951);
and U18876 (N_18876,N_17248,N_16224);
and U18877 (N_18877,N_17751,N_17421);
or U18878 (N_18878,N_17007,N_16653);
nor U18879 (N_18879,N_17282,N_17148);
nand U18880 (N_18880,N_17671,N_16811);
and U18881 (N_18881,N_16176,N_17501);
nand U18882 (N_18882,N_16722,N_16556);
xor U18883 (N_18883,N_16817,N_17103);
and U18884 (N_18884,N_16161,N_16298);
nand U18885 (N_18885,N_17213,N_16728);
nor U18886 (N_18886,N_16104,N_16616);
or U18887 (N_18887,N_16051,N_17500);
nor U18888 (N_18888,N_16364,N_16621);
nand U18889 (N_18889,N_16740,N_16974);
nor U18890 (N_18890,N_17621,N_16963);
xnor U18891 (N_18891,N_17216,N_17793);
nor U18892 (N_18892,N_17956,N_16242);
and U18893 (N_18893,N_17572,N_17770);
nand U18894 (N_18894,N_16909,N_17955);
or U18895 (N_18895,N_16591,N_16986);
or U18896 (N_18896,N_16523,N_17240);
or U18897 (N_18897,N_16824,N_16380);
or U18898 (N_18898,N_17608,N_17821);
nand U18899 (N_18899,N_16518,N_17528);
xor U18900 (N_18900,N_16868,N_16126);
nand U18901 (N_18901,N_17063,N_17665);
and U18902 (N_18902,N_16662,N_17969);
or U18903 (N_18903,N_17529,N_16979);
and U18904 (N_18904,N_16278,N_17910);
and U18905 (N_18905,N_16014,N_16315);
or U18906 (N_18906,N_17242,N_16197);
or U18907 (N_18907,N_16745,N_17741);
nand U18908 (N_18908,N_17134,N_17659);
nand U18909 (N_18909,N_17341,N_16642);
nor U18910 (N_18910,N_16223,N_17953);
nand U18911 (N_18911,N_17657,N_17557);
nand U18912 (N_18912,N_17319,N_16803);
or U18913 (N_18913,N_16987,N_16332);
nand U18914 (N_18914,N_16573,N_17279);
nand U18915 (N_18915,N_17009,N_17766);
xnor U18916 (N_18916,N_16684,N_17923);
nor U18917 (N_18917,N_16940,N_17971);
nand U18918 (N_18918,N_16169,N_16150);
nor U18919 (N_18919,N_16861,N_16634);
or U18920 (N_18920,N_17599,N_16620);
nand U18921 (N_18921,N_17596,N_17462);
nor U18922 (N_18922,N_17031,N_17416);
and U18923 (N_18923,N_16127,N_16689);
nor U18924 (N_18924,N_16134,N_16136);
nor U18925 (N_18925,N_16947,N_17170);
nand U18926 (N_18926,N_16039,N_17084);
and U18927 (N_18927,N_17437,N_16100);
nor U18928 (N_18928,N_16598,N_16236);
nand U18929 (N_18929,N_16853,N_16758);
nor U18930 (N_18930,N_17473,N_17873);
or U18931 (N_18931,N_17614,N_17212);
or U18932 (N_18932,N_16307,N_16818);
nand U18933 (N_18933,N_16848,N_17921);
and U18934 (N_18934,N_16956,N_16011);
nor U18935 (N_18935,N_17080,N_16641);
nand U18936 (N_18936,N_17064,N_17306);
or U18937 (N_18937,N_17618,N_17158);
nor U18938 (N_18938,N_17309,N_16017);
nor U18939 (N_18939,N_16442,N_17480);
and U18940 (N_18940,N_17686,N_17175);
and U18941 (N_18941,N_17716,N_16135);
xor U18942 (N_18942,N_16737,N_16808);
nand U18943 (N_18943,N_17046,N_16923);
or U18944 (N_18944,N_17363,N_16339);
nand U18945 (N_18945,N_16532,N_17972);
and U18946 (N_18946,N_16272,N_17442);
and U18947 (N_18947,N_16481,N_16670);
or U18948 (N_18948,N_16447,N_17446);
and U18949 (N_18949,N_17902,N_17281);
and U18950 (N_18950,N_16247,N_16886);
or U18951 (N_18951,N_17620,N_16441);
or U18952 (N_18952,N_17378,N_17048);
or U18953 (N_18953,N_16807,N_17737);
nor U18954 (N_18954,N_16845,N_16896);
and U18955 (N_18955,N_16571,N_16275);
nand U18956 (N_18956,N_16138,N_16091);
or U18957 (N_18957,N_17794,N_16455);
and U18958 (N_18958,N_16009,N_16164);
or U18959 (N_18959,N_17097,N_16636);
and U18960 (N_18960,N_16500,N_17691);
and U18961 (N_18961,N_17788,N_17295);
xnor U18962 (N_18962,N_17461,N_16592);
and U18963 (N_18963,N_17707,N_17805);
nor U18964 (N_18964,N_16578,N_17512);
nand U18965 (N_18965,N_17289,N_17913);
xor U18966 (N_18966,N_17651,N_16487);
xnor U18967 (N_18967,N_17895,N_16539);
and U18968 (N_18968,N_17402,N_17070);
or U18969 (N_18969,N_17393,N_16534);
nand U18970 (N_18970,N_17144,N_16123);
or U18971 (N_18971,N_17488,N_17694);
nor U18972 (N_18972,N_16054,N_16586);
nor U18973 (N_18973,N_17241,N_16838);
nand U18974 (N_18974,N_16605,N_16607);
nand U18975 (N_18975,N_16806,N_17807);
or U18976 (N_18976,N_17846,N_17264);
and U18977 (N_18977,N_16637,N_16217);
nor U18978 (N_18978,N_17177,N_16671);
or U18979 (N_18979,N_17813,N_17515);
or U18980 (N_18980,N_16052,N_17567);
or U18981 (N_18981,N_17720,N_17663);
or U18982 (N_18982,N_17081,N_16037);
nand U18983 (N_18983,N_16801,N_16042);
and U18984 (N_18984,N_16397,N_17507);
and U18985 (N_18985,N_17430,N_17336);
nand U18986 (N_18986,N_16361,N_16159);
and U18987 (N_18987,N_17230,N_17875);
or U18988 (N_18988,N_17232,N_17646);
nor U18989 (N_18989,N_16783,N_16869);
nor U18990 (N_18990,N_16835,N_17919);
and U18991 (N_18991,N_17867,N_17967);
xor U18992 (N_18992,N_16187,N_17779);
or U18993 (N_18993,N_16461,N_16537);
and U18994 (N_18994,N_16800,N_17749);
nand U18995 (N_18995,N_17348,N_17434);
nor U18996 (N_18996,N_17455,N_17145);
nor U18997 (N_18997,N_17125,N_17487);
and U18998 (N_18998,N_17361,N_16601);
or U18999 (N_18999,N_17072,N_17285);
nor U19000 (N_19000,N_16346,N_16841);
and U19001 (N_19001,N_16557,N_17877);
nand U19002 (N_19002,N_16400,N_17549);
and U19003 (N_19003,N_16608,N_16392);
xnor U19004 (N_19004,N_17860,N_17854);
xor U19005 (N_19005,N_17644,N_16264);
or U19006 (N_19006,N_16048,N_17354);
xnor U19007 (N_19007,N_16603,N_16321);
or U19008 (N_19008,N_16410,N_17017);
and U19009 (N_19009,N_16676,N_17590);
and U19010 (N_19010,N_16207,N_16097);
nor U19011 (N_19011,N_16148,N_17208);
or U19012 (N_19012,N_16166,N_17362);
nand U19013 (N_19013,N_17082,N_16915);
nand U19014 (N_19014,N_16356,N_17949);
or U19015 (N_19015,N_16464,N_17300);
nor U19016 (N_19016,N_16583,N_16712);
nor U19017 (N_19017,N_16982,N_17035);
nand U19018 (N_19018,N_17524,N_16758);
nand U19019 (N_19019,N_16205,N_16034);
xnor U19020 (N_19020,N_17635,N_17326);
nor U19021 (N_19021,N_16820,N_17269);
nand U19022 (N_19022,N_17889,N_17603);
xor U19023 (N_19023,N_17823,N_16201);
nor U19024 (N_19024,N_16050,N_17430);
nor U19025 (N_19025,N_17377,N_17852);
or U19026 (N_19026,N_17170,N_16792);
nor U19027 (N_19027,N_16267,N_16450);
and U19028 (N_19028,N_17777,N_16647);
and U19029 (N_19029,N_16004,N_17620);
and U19030 (N_19030,N_17206,N_16825);
or U19031 (N_19031,N_17435,N_16798);
xor U19032 (N_19032,N_16098,N_16487);
or U19033 (N_19033,N_17652,N_17620);
nor U19034 (N_19034,N_17434,N_16444);
nand U19035 (N_19035,N_17162,N_16790);
and U19036 (N_19036,N_16129,N_17109);
nor U19037 (N_19037,N_16436,N_16355);
nand U19038 (N_19038,N_17543,N_16377);
nand U19039 (N_19039,N_17160,N_17970);
or U19040 (N_19040,N_17732,N_17956);
or U19041 (N_19041,N_16416,N_17788);
or U19042 (N_19042,N_17849,N_16326);
nor U19043 (N_19043,N_17519,N_17119);
or U19044 (N_19044,N_17115,N_16423);
nand U19045 (N_19045,N_16540,N_17778);
and U19046 (N_19046,N_16293,N_17425);
and U19047 (N_19047,N_17359,N_17238);
and U19048 (N_19048,N_16738,N_17086);
and U19049 (N_19049,N_17307,N_16372);
nand U19050 (N_19050,N_16344,N_16554);
nor U19051 (N_19051,N_16946,N_16812);
and U19052 (N_19052,N_17636,N_17274);
and U19053 (N_19053,N_17720,N_17759);
or U19054 (N_19054,N_17477,N_16369);
nand U19055 (N_19055,N_16221,N_17200);
and U19056 (N_19056,N_16681,N_16830);
nor U19057 (N_19057,N_17728,N_16349);
nand U19058 (N_19058,N_16031,N_16370);
nor U19059 (N_19059,N_16087,N_16865);
nand U19060 (N_19060,N_17049,N_16774);
nand U19061 (N_19061,N_17278,N_17090);
nor U19062 (N_19062,N_16636,N_16816);
and U19063 (N_19063,N_16359,N_16519);
xor U19064 (N_19064,N_17631,N_17743);
nand U19065 (N_19065,N_17584,N_16048);
nor U19066 (N_19066,N_17656,N_16350);
nand U19067 (N_19067,N_16831,N_16347);
or U19068 (N_19068,N_17018,N_16164);
nor U19069 (N_19069,N_17782,N_16306);
and U19070 (N_19070,N_16713,N_17661);
or U19071 (N_19071,N_16475,N_16242);
nand U19072 (N_19072,N_16234,N_16949);
nand U19073 (N_19073,N_16205,N_16791);
and U19074 (N_19074,N_16672,N_17565);
xor U19075 (N_19075,N_16490,N_17904);
or U19076 (N_19076,N_17586,N_16005);
nor U19077 (N_19077,N_16076,N_17446);
xnor U19078 (N_19078,N_16897,N_17067);
nand U19079 (N_19079,N_17543,N_17685);
nor U19080 (N_19080,N_17636,N_16034);
nand U19081 (N_19081,N_17224,N_17180);
nand U19082 (N_19082,N_16433,N_17017);
or U19083 (N_19083,N_17060,N_16800);
and U19084 (N_19084,N_17466,N_17500);
nor U19085 (N_19085,N_17591,N_17589);
or U19086 (N_19086,N_16921,N_16272);
xor U19087 (N_19087,N_17100,N_16879);
xor U19088 (N_19088,N_16031,N_16217);
and U19089 (N_19089,N_16980,N_16570);
nand U19090 (N_19090,N_16192,N_17539);
and U19091 (N_19091,N_16012,N_17298);
or U19092 (N_19092,N_17813,N_17448);
nand U19093 (N_19093,N_16020,N_16617);
nand U19094 (N_19094,N_17811,N_16169);
nand U19095 (N_19095,N_16036,N_16429);
nor U19096 (N_19096,N_17303,N_17233);
xnor U19097 (N_19097,N_17308,N_17749);
or U19098 (N_19098,N_16061,N_16898);
and U19099 (N_19099,N_16274,N_16381);
nor U19100 (N_19100,N_16807,N_16150);
xor U19101 (N_19101,N_16855,N_17228);
xor U19102 (N_19102,N_16024,N_17170);
nand U19103 (N_19103,N_16042,N_17613);
or U19104 (N_19104,N_16204,N_16831);
and U19105 (N_19105,N_16796,N_17123);
or U19106 (N_19106,N_17741,N_16442);
nor U19107 (N_19107,N_16270,N_16602);
nand U19108 (N_19108,N_17482,N_16597);
or U19109 (N_19109,N_17210,N_16693);
nand U19110 (N_19110,N_17119,N_17576);
or U19111 (N_19111,N_17925,N_16217);
nor U19112 (N_19112,N_16878,N_17244);
nand U19113 (N_19113,N_17796,N_17705);
nand U19114 (N_19114,N_17103,N_17901);
and U19115 (N_19115,N_16539,N_17482);
xor U19116 (N_19116,N_17788,N_16175);
or U19117 (N_19117,N_16696,N_17717);
or U19118 (N_19118,N_16871,N_16616);
xnor U19119 (N_19119,N_16654,N_17893);
and U19120 (N_19120,N_16211,N_16942);
nand U19121 (N_19121,N_16423,N_17000);
and U19122 (N_19122,N_16400,N_17432);
nor U19123 (N_19123,N_16370,N_17078);
nor U19124 (N_19124,N_17354,N_17232);
or U19125 (N_19125,N_16665,N_16788);
and U19126 (N_19126,N_17307,N_17800);
nor U19127 (N_19127,N_17423,N_17381);
nand U19128 (N_19128,N_17777,N_16714);
or U19129 (N_19129,N_17933,N_16452);
and U19130 (N_19130,N_17136,N_16358);
nand U19131 (N_19131,N_16112,N_16920);
nor U19132 (N_19132,N_17125,N_16621);
nand U19133 (N_19133,N_17467,N_17170);
nor U19134 (N_19134,N_17846,N_16298);
nor U19135 (N_19135,N_16513,N_16745);
nand U19136 (N_19136,N_17829,N_16788);
nand U19137 (N_19137,N_17995,N_17136);
xor U19138 (N_19138,N_16864,N_17752);
or U19139 (N_19139,N_16039,N_17736);
xor U19140 (N_19140,N_17426,N_16030);
or U19141 (N_19141,N_17081,N_16442);
nor U19142 (N_19142,N_16533,N_17607);
xor U19143 (N_19143,N_16718,N_17960);
or U19144 (N_19144,N_17732,N_16453);
nor U19145 (N_19145,N_17648,N_16276);
or U19146 (N_19146,N_16512,N_17392);
nor U19147 (N_19147,N_17823,N_17426);
nor U19148 (N_19148,N_17620,N_16096);
and U19149 (N_19149,N_17623,N_16151);
xor U19150 (N_19150,N_16381,N_17995);
nand U19151 (N_19151,N_16264,N_17554);
nand U19152 (N_19152,N_16510,N_17689);
xor U19153 (N_19153,N_16502,N_17782);
or U19154 (N_19154,N_17348,N_17734);
and U19155 (N_19155,N_16657,N_16958);
or U19156 (N_19156,N_17648,N_16391);
and U19157 (N_19157,N_16734,N_17647);
and U19158 (N_19158,N_17055,N_17570);
and U19159 (N_19159,N_16741,N_17686);
nand U19160 (N_19160,N_17115,N_16217);
and U19161 (N_19161,N_17957,N_17588);
or U19162 (N_19162,N_16421,N_17383);
nand U19163 (N_19163,N_17808,N_16608);
nor U19164 (N_19164,N_16382,N_17029);
or U19165 (N_19165,N_17893,N_16336);
or U19166 (N_19166,N_16452,N_17510);
or U19167 (N_19167,N_17467,N_16584);
nand U19168 (N_19168,N_17362,N_16045);
nand U19169 (N_19169,N_16571,N_16584);
nand U19170 (N_19170,N_17989,N_17224);
or U19171 (N_19171,N_17861,N_17969);
nand U19172 (N_19172,N_16124,N_16615);
nor U19173 (N_19173,N_17664,N_16090);
and U19174 (N_19174,N_16653,N_16315);
or U19175 (N_19175,N_16629,N_17545);
and U19176 (N_19176,N_16952,N_17389);
nand U19177 (N_19177,N_17151,N_16700);
and U19178 (N_19178,N_16770,N_16182);
and U19179 (N_19179,N_17766,N_17745);
nand U19180 (N_19180,N_16501,N_16250);
nor U19181 (N_19181,N_16610,N_16370);
nand U19182 (N_19182,N_17332,N_16525);
or U19183 (N_19183,N_16915,N_16788);
and U19184 (N_19184,N_16123,N_16899);
and U19185 (N_19185,N_16433,N_16510);
xor U19186 (N_19186,N_17321,N_16723);
nand U19187 (N_19187,N_16374,N_17902);
xnor U19188 (N_19188,N_16765,N_16320);
nor U19189 (N_19189,N_17408,N_16795);
or U19190 (N_19190,N_16807,N_17558);
nand U19191 (N_19191,N_17429,N_16249);
nand U19192 (N_19192,N_16076,N_16894);
or U19193 (N_19193,N_16894,N_17094);
nor U19194 (N_19194,N_17596,N_17260);
nand U19195 (N_19195,N_16159,N_16955);
xnor U19196 (N_19196,N_16388,N_17811);
nand U19197 (N_19197,N_16062,N_16664);
nor U19198 (N_19198,N_16127,N_17077);
nor U19199 (N_19199,N_16746,N_16552);
or U19200 (N_19200,N_17378,N_16007);
and U19201 (N_19201,N_17621,N_16248);
and U19202 (N_19202,N_16499,N_17115);
nor U19203 (N_19203,N_17075,N_17607);
nor U19204 (N_19204,N_17860,N_16285);
or U19205 (N_19205,N_16330,N_17775);
and U19206 (N_19206,N_17425,N_17282);
and U19207 (N_19207,N_17567,N_16497);
xor U19208 (N_19208,N_16081,N_16029);
or U19209 (N_19209,N_17013,N_16724);
nand U19210 (N_19210,N_17403,N_17551);
and U19211 (N_19211,N_17883,N_17885);
or U19212 (N_19212,N_16504,N_17346);
nor U19213 (N_19213,N_16538,N_16294);
xnor U19214 (N_19214,N_17507,N_17706);
nand U19215 (N_19215,N_17560,N_16775);
or U19216 (N_19216,N_16356,N_17776);
nor U19217 (N_19217,N_16063,N_17232);
xnor U19218 (N_19218,N_16597,N_17810);
and U19219 (N_19219,N_17118,N_17839);
and U19220 (N_19220,N_17141,N_17751);
nor U19221 (N_19221,N_16687,N_16456);
nor U19222 (N_19222,N_16930,N_17213);
nor U19223 (N_19223,N_17091,N_16244);
or U19224 (N_19224,N_16544,N_16360);
xor U19225 (N_19225,N_17155,N_17012);
or U19226 (N_19226,N_17360,N_16103);
xor U19227 (N_19227,N_17819,N_17687);
or U19228 (N_19228,N_17402,N_17215);
xor U19229 (N_19229,N_17623,N_16255);
nor U19230 (N_19230,N_16407,N_16091);
and U19231 (N_19231,N_16924,N_16401);
nand U19232 (N_19232,N_16832,N_16288);
or U19233 (N_19233,N_17804,N_16373);
nor U19234 (N_19234,N_16822,N_17590);
nand U19235 (N_19235,N_16273,N_16228);
and U19236 (N_19236,N_16193,N_16552);
xor U19237 (N_19237,N_17359,N_16402);
nor U19238 (N_19238,N_17959,N_17601);
or U19239 (N_19239,N_16636,N_16373);
nor U19240 (N_19240,N_16028,N_16193);
nor U19241 (N_19241,N_17891,N_16543);
nand U19242 (N_19242,N_16566,N_17579);
or U19243 (N_19243,N_17752,N_17955);
nor U19244 (N_19244,N_17556,N_16223);
or U19245 (N_19245,N_16438,N_17648);
nand U19246 (N_19246,N_17848,N_17619);
or U19247 (N_19247,N_17908,N_17835);
nand U19248 (N_19248,N_17904,N_16507);
xnor U19249 (N_19249,N_17602,N_16287);
xor U19250 (N_19250,N_16205,N_16629);
nand U19251 (N_19251,N_17193,N_16522);
or U19252 (N_19252,N_17060,N_17229);
and U19253 (N_19253,N_16419,N_16738);
xor U19254 (N_19254,N_17909,N_16231);
nor U19255 (N_19255,N_16684,N_17197);
nor U19256 (N_19256,N_17147,N_17562);
nand U19257 (N_19257,N_17041,N_16994);
nor U19258 (N_19258,N_16629,N_16429);
or U19259 (N_19259,N_17081,N_17038);
and U19260 (N_19260,N_16237,N_16226);
nor U19261 (N_19261,N_16508,N_17460);
nor U19262 (N_19262,N_16855,N_16529);
nor U19263 (N_19263,N_17160,N_17476);
nand U19264 (N_19264,N_17962,N_16821);
nor U19265 (N_19265,N_16260,N_16024);
nor U19266 (N_19266,N_16542,N_16872);
and U19267 (N_19267,N_17382,N_17229);
nand U19268 (N_19268,N_17376,N_17757);
nand U19269 (N_19269,N_16138,N_16418);
or U19270 (N_19270,N_17021,N_17506);
nor U19271 (N_19271,N_16328,N_16534);
nand U19272 (N_19272,N_17727,N_16642);
nand U19273 (N_19273,N_16251,N_17120);
nor U19274 (N_19274,N_16060,N_17548);
or U19275 (N_19275,N_16023,N_16679);
nor U19276 (N_19276,N_17299,N_17047);
nor U19277 (N_19277,N_16626,N_17207);
nor U19278 (N_19278,N_17568,N_17697);
or U19279 (N_19279,N_16749,N_16032);
and U19280 (N_19280,N_17205,N_17619);
nor U19281 (N_19281,N_16686,N_17699);
nor U19282 (N_19282,N_17552,N_17806);
nand U19283 (N_19283,N_17351,N_16084);
or U19284 (N_19284,N_16728,N_16720);
nor U19285 (N_19285,N_16274,N_16062);
nand U19286 (N_19286,N_16270,N_17180);
nor U19287 (N_19287,N_17345,N_17623);
nand U19288 (N_19288,N_17807,N_16402);
nor U19289 (N_19289,N_17424,N_17889);
and U19290 (N_19290,N_16289,N_17185);
xnor U19291 (N_19291,N_17158,N_17996);
and U19292 (N_19292,N_16147,N_16208);
or U19293 (N_19293,N_17902,N_17899);
and U19294 (N_19294,N_17030,N_16000);
xor U19295 (N_19295,N_17120,N_17484);
and U19296 (N_19296,N_16765,N_17484);
and U19297 (N_19297,N_17985,N_16172);
nand U19298 (N_19298,N_17224,N_16346);
and U19299 (N_19299,N_17041,N_17819);
or U19300 (N_19300,N_16919,N_17281);
xnor U19301 (N_19301,N_17860,N_17817);
or U19302 (N_19302,N_16278,N_16077);
or U19303 (N_19303,N_16377,N_17568);
and U19304 (N_19304,N_17041,N_17940);
or U19305 (N_19305,N_16610,N_16555);
nor U19306 (N_19306,N_17738,N_16386);
or U19307 (N_19307,N_17968,N_17474);
and U19308 (N_19308,N_17944,N_16350);
or U19309 (N_19309,N_16583,N_17501);
xnor U19310 (N_19310,N_16545,N_17513);
or U19311 (N_19311,N_17962,N_16905);
and U19312 (N_19312,N_17098,N_17002);
nand U19313 (N_19313,N_16364,N_17649);
xnor U19314 (N_19314,N_16712,N_16143);
nor U19315 (N_19315,N_17244,N_16754);
nand U19316 (N_19316,N_16944,N_17473);
nand U19317 (N_19317,N_17809,N_17437);
nand U19318 (N_19318,N_16512,N_17725);
nor U19319 (N_19319,N_17428,N_16204);
nor U19320 (N_19320,N_16977,N_16899);
nand U19321 (N_19321,N_17319,N_17698);
xnor U19322 (N_19322,N_17868,N_17837);
nand U19323 (N_19323,N_16149,N_16500);
or U19324 (N_19324,N_17515,N_16664);
and U19325 (N_19325,N_16695,N_16843);
and U19326 (N_19326,N_16359,N_16937);
and U19327 (N_19327,N_17554,N_16300);
and U19328 (N_19328,N_17137,N_17391);
nor U19329 (N_19329,N_16433,N_17420);
or U19330 (N_19330,N_17251,N_16358);
nand U19331 (N_19331,N_17239,N_17932);
and U19332 (N_19332,N_16806,N_16734);
and U19333 (N_19333,N_17178,N_17736);
or U19334 (N_19334,N_17085,N_16137);
nor U19335 (N_19335,N_16064,N_16418);
xnor U19336 (N_19336,N_17654,N_17960);
or U19337 (N_19337,N_16028,N_17211);
or U19338 (N_19338,N_16266,N_16809);
nor U19339 (N_19339,N_17188,N_16378);
nand U19340 (N_19340,N_16540,N_17032);
nor U19341 (N_19341,N_17934,N_16833);
nand U19342 (N_19342,N_16676,N_17885);
nor U19343 (N_19343,N_16217,N_16140);
or U19344 (N_19344,N_17212,N_17618);
nand U19345 (N_19345,N_17014,N_17585);
nand U19346 (N_19346,N_16647,N_16826);
and U19347 (N_19347,N_17543,N_17609);
nand U19348 (N_19348,N_16559,N_17805);
nand U19349 (N_19349,N_17196,N_17617);
nor U19350 (N_19350,N_16529,N_17895);
nor U19351 (N_19351,N_17299,N_17553);
nor U19352 (N_19352,N_17691,N_16158);
nand U19353 (N_19353,N_17333,N_16405);
and U19354 (N_19354,N_17557,N_17997);
nor U19355 (N_19355,N_16338,N_17844);
nor U19356 (N_19356,N_16697,N_17389);
or U19357 (N_19357,N_17524,N_16833);
nand U19358 (N_19358,N_16771,N_16751);
nand U19359 (N_19359,N_17995,N_16714);
nand U19360 (N_19360,N_16009,N_16135);
nor U19361 (N_19361,N_16691,N_17438);
and U19362 (N_19362,N_17573,N_17393);
and U19363 (N_19363,N_16667,N_17516);
nor U19364 (N_19364,N_17795,N_17346);
nor U19365 (N_19365,N_17321,N_17689);
and U19366 (N_19366,N_17348,N_17731);
xor U19367 (N_19367,N_16657,N_17393);
nand U19368 (N_19368,N_16723,N_16140);
or U19369 (N_19369,N_16932,N_16382);
xor U19370 (N_19370,N_17294,N_16340);
nor U19371 (N_19371,N_16789,N_16706);
and U19372 (N_19372,N_17524,N_16834);
and U19373 (N_19373,N_16745,N_17704);
or U19374 (N_19374,N_16353,N_17624);
nor U19375 (N_19375,N_16060,N_16797);
and U19376 (N_19376,N_17147,N_16282);
or U19377 (N_19377,N_16767,N_16517);
and U19378 (N_19378,N_17059,N_16794);
or U19379 (N_19379,N_16191,N_17229);
nor U19380 (N_19380,N_16907,N_17348);
or U19381 (N_19381,N_17004,N_16677);
nand U19382 (N_19382,N_17986,N_16353);
or U19383 (N_19383,N_17367,N_16492);
nor U19384 (N_19384,N_16436,N_16610);
nand U19385 (N_19385,N_16258,N_17419);
nor U19386 (N_19386,N_16298,N_17125);
and U19387 (N_19387,N_16256,N_16650);
nand U19388 (N_19388,N_16594,N_16924);
nor U19389 (N_19389,N_16599,N_16580);
nand U19390 (N_19390,N_17905,N_17971);
nand U19391 (N_19391,N_16404,N_17585);
and U19392 (N_19392,N_17156,N_16748);
or U19393 (N_19393,N_17000,N_16455);
nor U19394 (N_19394,N_17453,N_17246);
nor U19395 (N_19395,N_17190,N_17397);
and U19396 (N_19396,N_17928,N_17214);
nor U19397 (N_19397,N_17580,N_17060);
and U19398 (N_19398,N_17137,N_17986);
nand U19399 (N_19399,N_16566,N_17407);
xor U19400 (N_19400,N_16860,N_17214);
nor U19401 (N_19401,N_16526,N_16321);
xnor U19402 (N_19402,N_17265,N_16192);
nand U19403 (N_19403,N_16984,N_16980);
and U19404 (N_19404,N_16640,N_16846);
and U19405 (N_19405,N_17009,N_17625);
nand U19406 (N_19406,N_16777,N_17601);
or U19407 (N_19407,N_16177,N_16305);
and U19408 (N_19408,N_16847,N_17731);
xnor U19409 (N_19409,N_17056,N_16197);
nor U19410 (N_19410,N_17654,N_17501);
nand U19411 (N_19411,N_17387,N_17578);
nand U19412 (N_19412,N_17807,N_16943);
xor U19413 (N_19413,N_17715,N_17924);
and U19414 (N_19414,N_17001,N_16677);
and U19415 (N_19415,N_17466,N_16027);
or U19416 (N_19416,N_16658,N_17831);
and U19417 (N_19417,N_16513,N_16541);
nor U19418 (N_19418,N_17300,N_16097);
nor U19419 (N_19419,N_17224,N_16629);
and U19420 (N_19420,N_17262,N_16683);
and U19421 (N_19421,N_16613,N_17091);
nor U19422 (N_19422,N_17406,N_17153);
and U19423 (N_19423,N_17884,N_16123);
and U19424 (N_19424,N_16722,N_17768);
and U19425 (N_19425,N_17991,N_16962);
and U19426 (N_19426,N_17572,N_17359);
and U19427 (N_19427,N_16262,N_16559);
xnor U19428 (N_19428,N_17809,N_16542);
nor U19429 (N_19429,N_17975,N_16497);
or U19430 (N_19430,N_16700,N_16862);
nand U19431 (N_19431,N_16345,N_16059);
or U19432 (N_19432,N_17539,N_16526);
and U19433 (N_19433,N_16511,N_17737);
nor U19434 (N_19434,N_16343,N_17812);
nand U19435 (N_19435,N_17220,N_16108);
or U19436 (N_19436,N_16947,N_16360);
xor U19437 (N_19437,N_16258,N_16777);
nor U19438 (N_19438,N_17559,N_17595);
nand U19439 (N_19439,N_16635,N_17522);
nor U19440 (N_19440,N_16104,N_16095);
and U19441 (N_19441,N_17427,N_16286);
xor U19442 (N_19442,N_17938,N_16095);
or U19443 (N_19443,N_17963,N_17585);
nor U19444 (N_19444,N_16703,N_16562);
or U19445 (N_19445,N_17376,N_17266);
and U19446 (N_19446,N_17194,N_16320);
nor U19447 (N_19447,N_16462,N_16973);
nor U19448 (N_19448,N_16696,N_17256);
nor U19449 (N_19449,N_16017,N_17999);
and U19450 (N_19450,N_16878,N_16948);
or U19451 (N_19451,N_16524,N_16349);
and U19452 (N_19452,N_17268,N_17190);
nor U19453 (N_19453,N_17988,N_17528);
and U19454 (N_19454,N_17599,N_16049);
nor U19455 (N_19455,N_17298,N_17410);
and U19456 (N_19456,N_17929,N_17225);
nor U19457 (N_19457,N_16193,N_17554);
nor U19458 (N_19458,N_17757,N_17805);
nand U19459 (N_19459,N_17765,N_16486);
nor U19460 (N_19460,N_17199,N_16845);
nand U19461 (N_19461,N_17296,N_17028);
nand U19462 (N_19462,N_16217,N_17082);
and U19463 (N_19463,N_17736,N_16798);
and U19464 (N_19464,N_16105,N_16322);
or U19465 (N_19465,N_17948,N_16743);
or U19466 (N_19466,N_17355,N_16029);
and U19467 (N_19467,N_17739,N_16150);
or U19468 (N_19468,N_17798,N_16832);
nor U19469 (N_19469,N_17008,N_16190);
nor U19470 (N_19470,N_16111,N_17324);
and U19471 (N_19471,N_16895,N_16625);
or U19472 (N_19472,N_17915,N_16623);
and U19473 (N_19473,N_17836,N_17418);
or U19474 (N_19474,N_17016,N_16352);
and U19475 (N_19475,N_16232,N_16477);
and U19476 (N_19476,N_16577,N_16850);
or U19477 (N_19477,N_17045,N_16040);
nor U19478 (N_19478,N_17251,N_16450);
or U19479 (N_19479,N_16854,N_16730);
and U19480 (N_19480,N_16733,N_17366);
xnor U19481 (N_19481,N_17223,N_17089);
xor U19482 (N_19482,N_17897,N_17639);
xnor U19483 (N_19483,N_16106,N_16496);
xnor U19484 (N_19484,N_17644,N_17353);
or U19485 (N_19485,N_17112,N_17997);
or U19486 (N_19486,N_16979,N_16530);
or U19487 (N_19487,N_17056,N_17789);
nor U19488 (N_19488,N_16089,N_16380);
and U19489 (N_19489,N_17631,N_16657);
nand U19490 (N_19490,N_16649,N_16520);
nor U19491 (N_19491,N_16187,N_16022);
nor U19492 (N_19492,N_16540,N_16597);
nor U19493 (N_19493,N_16950,N_16442);
nor U19494 (N_19494,N_17503,N_17968);
nand U19495 (N_19495,N_17978,N_17470);
nand U19496 (N_19496,N_16386,N_16556);
and U19497 (N_19497,N_16443,N_17964);
nor U19498 (N_19498,N_16718,N_16180);
xor U19499 (N_19499,N_17834,N_17019);
nor U19500 (N_19500,N_16539,N_17480);
nand U19501 (N_19501,N_17780,N_17192);
and U19502 (N_19502,N_16594,N_17338);
nand U19503 (N_19503,N_17559,N_17085);
nand U19504 (N_19504,N_17770,N_16025);
nand U19505 (N_19505,N_17971,N_17322);
nand U19506 (N_19506,N_16773,N_16237);
or U19507 (N_19507,N_17003,N_17710);
nand U19508 (N_19508,N_17170,N_16890);
or U19509 (N_19509,N_17951,N_17437);
or U19510 (N_19510,N_16407,N_17318);
nor U19511 (N_19511,N_17913,N_17047);
or U19512 (N_19512,N_17347,N_16678);
nand U19513 (N_19513,N_17058,N_17211);
and U19514 (N_19514,N_16101,N_16700);
xnor U19515 (N_19515,N_16141,N_17924);
and U19516 (N_19516,N_16624,N_17090);
and U19517 (N_19517,N_16924,N_17557);
nor U19518 (N_19518,N_16331,N_16211);
and U19519 (N_19519,N_17517,N_17722);
nor U19520 (N_19520,N_17094,N_17229);
or U19521 (N_19521,N_17792,N_17054);
and U19522 (N_19522,N_16175,N_17154);
and U19523 (N_19523,N_16515,N_16143);
and U19524 (N_19524,N_17758,N_17674);
and U19525 (N_19525,N_16703,N_17045);
or U19526 (N_19526,N_17293,N_16062);
and U19527 (N_19527,N_16370,N_16132);
or U19528 (N_19528,N_17055,N_16318);
xor U19529 (N_19529,N_16109,N_16747);
and U19530 (N_19530,N_16802,N_17841);
nor U19531 (N_19531,N_17982,N_17866);
or U19532 (N_19532,N_17335,N_17225);
nor U19533 (N_19533,N_16334,N_16245);
and U19534 (N_19534,N_17166,N_17817);
and U19535 (N_19535,N_16271,N_16427);
or U19536 (N_19536,N_17401,N_17590);
and U19537 (N_19537,N_16958,N_17637);
and U19538 (N_19538,N_16804,N_16272);
and U19539 (N_19539,N_17132,N_17275);
nand U19540 (N_19540,N_17556,N_17085);
nand U19541 (N_19541,N_17279,N_17910);
or U19542 (N_19542,N_16586,N_16250);
nor U19543 (N_19543,N_16074,N_17956);
nor U19544 (N_19544,N_17533,N_16052);
xor U19545 (N_19545,N_16711,N_16477);
and U19546 (N_19546,N_17215,N_17743);
or U19547 (N_19547,N_17468,N_16539);
xor U19548 (N_19548,N_16347,N_17662);
or U19549 (N_19549,N_16006,N_16492);
or U19550 (N_19550,N_16118,N_17138);
and U19551 (N_19551,N_17224,N_16048);
and U19552 (N_19552,N_16671,N_16049);
and U19553 (N_19553,N_17025,N_16909);
and U19554 (N_19554,N_16956,N_17367);
xor U19555 (N_19555,N_16050,N_16291);
or U19556 (N_19556,N_16579,N_16601);
or U19557 (N_19557,N_17037,N_17427);
or U19558 (N_19558,N_16151,N_17166);
xnor U19559 (N_19559,N_16517,N_16770);
nor U19560 (N_19560,N_16446,N_17373);
xnor U19561 (N_19561,N_16153,N_16019);
and U19562 (N_19562,N_17741,N_17165);
or U19563 (N_19563,N_17539,N_17834);
nand U19564 (N_19564,N_17051,N_17841);
and U19565 (N_19565,N_16957,N_16175);
or U19566 (N_19566,N_17138,N_16441);
and U19567 (N_19567,N_16595,N_17758);
or U19568 (N_19568,N_17735,N_17679);
or U19569 (N_19569,N_17278,N_17308);
and U19570 (N_19570,N_17755,N_16416);
or U19571 (N_19571,N_17341,N_16419);
nand U19572 (N_19572,N_16497,N_17067);
nand U19573 (N_19573,N_17335,N_16920);
nand U19574 (N_19574,N_17238,N_17225);
nor U19575 (N_19575,N_17901,N_16662);
nor U19576 (N_19576,N_16943,N_17798);
or U19577 (N_19577,N_16054,N_17538);
xor U19578 (N_19578,N_17924,N_17914);
nand U19579 (N_19579,N_16356,N_17435);
or U19580 (N_19580,N_17600,N_17338);
and U19581 (N_19581,N_17830,N_17646);
or U19582 (N_19582,N_17689,N_16046);
and U19583 (N_19583,N_17453,N_17228);
nor U19584 (N_19584,N_17516,N_17241);
and U19585 (N_19585,N_17479,N_16484);
nor U19586 (N_19586,N_16394,N_16199);
and U19587 (N_19587,N_16542,N_17957);
nand U19588 (N_19588,N_16692,N_17366);
nor U19589 (N_19589,N_17576,N_17350);
or U19590 (N_19590,N_16571,N_16479);
and U19591 (N_19591,N_16720,N_16188);
and U19592 (N_19592,N_16956,N_16224);
and U19593 (N_19593,N_16687,N_17429);
or U19594 (N_19594,N_17073,N_16390);
nand U19595 (N_19595,N_17529,N_16992);
and U19596 (N_19596,N_16288,N_16132);
nand U19597 (N_19597,N_16002,N_17103);
xnor U19598 (N_19598,N_17080,N_16266);
nor U19599 (N_19599,N_17251,N_16673);
or U19600 (N_19600,N_16138,N_17709);
or U19601 (N_19601,N_17814,N_17800);
xnor U19602 (N_19602,N_16054,N_16652);
nand U19603 (N_19603,N_17797,N_17196);
nand U19604 (N_19604,N_16345,N_16482);
nand U19605 (N_19605,N_17318,N_17232);
and U19606 (N_19606,N_17376,N_17986);
nand U19607 (N_19607,N_16070,N_16308);
nor U19608 (N_19608,N_16736,N_17826);
and U19609 (N_19609,N_17236,N_17138);
or U19610 (N_19610,N_16012,N_16344);
xor U19611 (N_19611,N_16835,N_16941);
nor U19612 (N_19612,N_16266,N_17812);
and U19613 (N_19613,N_16079,N_17709);
nor U19614 (N_19614,N_17833,N_17573);
nor U19615 (N_19615,N_16772,N_16803);
and U19616 (N_19616,N_16799,N_17023);
or U19617 (N_19617,N_16934,N_17276);
nor U19618 (N_19618,N_17949,N_16934);
nor U19619 (N_19619,N_16285,N_17913);
nor U19620 (N_19620,N_17702,N_16791);
nand U19621 (N_19621,N_16331,N_17542);
nand U19622 (N_19622,N_17515,N_16653);
nor U19623 (N_19623,N_17214,N_17133);
or U19624 (N_19624,N_16837,N_17274);
nand U19625 (N_19625,N_16699,N_17888);
xnor U19626 (N_19626,N_16491,N_17051);
nand U19627 (N_19627,N_17965,N_17068);
nand U19628 (N_19628,N_17567,N_16393);
xnor U19629 (N_19629,N_16206,N_16321);
nand U19630 (N_19630,N_17115,N_16412);
and U19631 (N_19631,N_17100,N_17728);
or U19632 (N_19632,N_17159,N_16052);
nand U19633 (N_19633,N_17827,N_17445);
or U19634 (N_19634,N_17478,N_17673);
and U19635 (N_19635,N_17481,N_16925);
nor U19636 (N_19636,N_17571,N_16975);
or U19637 (N_19637,N_17885,N_16173);
and U19638 (N_19638,N_17811,N_16787);
nand U19639 (N_19639,N_16465,N_17060);
and U19640 (N_19640,N_16755,N_16613);
nand U19641 (N_19641,N_16708,N_16911);
nand U19642 (N_19642,N_16285,N_16539);
nand U19643 (N_19643,N_16970,N_16858);
nor U19644 (N_19644,N_16773,N_17812);
xor U19645 (N_19645,N_17471,N_16133);
nor U19646 (N_19646,N_16997,N_17779);
or U19647 (N_19647,N_17883,N_16635);
nand U19648 (N_19648,N_17749,N_17586);
nor U19649 (N_19649,N_16823,N_17002);
nand U19650 (N_19650,N_17656,N_16266);
or U19651 (N_19651,N_17191,N_16790);
xor U19652 (N_19652,N_16181,N_16984);
or U19653 (N_19653,N_17814,N_16005);
nand U19654 (N_19654,N_16805,N_17374);
and U19655 (N_19655,N_17844,N_16108);
nand U19656 (N_19656,N_16550,N_16862);
nor U19657 (N_19657,N_16676,N_17811);
nand U19658 (N_19658,N_16814,N_17895);
or U19659 (N_19659,N_17499,N_17446);
or U19660 (N_19660,N_16055,N_16727);
and U19661 (N_19661,N_16307,N_17691);
and U19662 (N_19662,N_16769,N_16626);
nor U19663 (N_19663,N_17971,N_17923);
nor U19664 (N_19664,N_17654,N_17087);
and U19665 (N_19665,N_17792,N_16202);
nor U19666 (N_19666,N_17538,N_17661);
and U19667 (N_19667,N_16158,N_17250);
or U19668 (N_19668,N_16467,N_16350);
nand U19669 (N_19669,N_16954,N_17343);
nor U19670 (N_19670,N_17371,N_16005);
nand U19671 (N_19671,N_16142,N_17739);
nor U19672 (N_19672,N_16180,N_16291);
and U19673 (N_19673,N_17625,N_17809);
or U19674 (N_19674,N_17128,N_17335);
xnor U19675 (N_19675,N_16096,N_16831);
nor U19676 (N_19676,N_17448,N_17687);
and U19677 (N_19677,N_16387,N_16578);
or U19678 (N_19678,N_16390,N_16443);
xor U19679 (N_19679,N_16562,N_16181);
or U19680 (N_19680,N_17895,N_17040);
and U19681 (N_19681,N_17298,N_17513);
or U19682 (N_19682,N_17086,N_16626);
xnor U19683 (N_19683,N_16915,N_16851);
nand U19684 (N_19684,N_17718,N_16606);
nor U19685 (N_19685,N_17209,N_16844);
xnor U19686 (N_19686,N_17468,N_17546);
xor U19687 (N_19687,N_16525,N_16836);
or U19688 (N_19688,N_17101,N_17540);
or U19689 (N_19689,N_16907,N_16799);
nor U19690 (N_19690,N_16513,N_17360);
and U19691 (N_19691,N_16879,N_16082);
nor U19692 (N_19692,N_17530,N_16248);
or U19693 (N_19693,N_17378,N_17229);
nand U19694 (N_19694,N_17031,N_16065);
or U19695 (N_19695,N_16975,N_16452);
nand U19696 (N_19696,N_16641,N_16883);
nor U19697 (N_19697,N_16044,N_17759);
nor U19698 (N_19698,N_16937,N_17165);
nand U19699 (N_19699,N_17329,N_16254);
nand U19700 (N_19700,N_17300,N_17426);
nand U19701 (N_19701,N_16648,N_16159);
and U19702 (N_19702,N_16645,N_16985);
nor U19703 (N_19703,N_17782,N_17159);
nand U19704 (N_19704,N_17311,N_16517);
or U19705 (N_19705,N_17374,N_17854);
nor U19706 (N_19706,N_17316,N_16601);
and U19707 (N_19707,N_16288,N_17585);
or U19708 (N_19708,N_16467,N_17973);
and U19709 (N_19709,N_16889,N_17284);
or U19710 (N_19710,N_17583,N_17337);
and U19711 (N_19711,N_16497,N_17186);
or U19712 (N_19712,N_17406,N_16395);
nor U19713 (N_19713,N_17927,N_16131);
xor U19714 (N_19714,N_16399,N_17854);
nand U19715 (N_19715,N_17765,N_16015);
or U19716 (N_19716,N_17937,N_17663);
nor U19717 (N_19717,N_17695,N_16534);
nor U19718 (N_19718,N_17551,N_16913);
or U19719 (N_19719,N_16403,N_17379);
or U19720 (N_19720,N_17073,N_17228);
nand U19721 (N_19721,N_16488,N_16027);
or U19722 (N_19722,N_17234,N_17725);
nor U19723 (N_19723,N_16752,N_16494);
or U19724 (N_19724,N_17716,N_17125);
and U19725 (N_19725,N_16454,N_16919);
or U19726 (N_19726,N_17916,N_17482);
and U19727 (N_19727,N_16763,N_16290);
nand U19728 (N_19728,N_17464,N_17717);
nor U19729 (N_19729,N_17999,N_17384);
xor U19730 (N_19730,N_16655,N_17117);
nand U19731 (N_19731,N_16829,N_16910);
xnor U19732 (N_19732,N_17713,N_17384);
nand U19733 (N_19733,N_16247,N_16234);
nor U19734 (N_19734,N_17214,N_16087);
nand U19735 (N_19735,N_17453,N_16392);
or U19736 (N_19736,N_17734,N_16049);
or U19737 (N_19737,N_17339,N_16455);
nor U19738 (N_19738,N_16457,N_17494);
or U19739 (N_19739,N_17699,N_16831);
nand U19740 (N_19740,N_16737,N_17012);
and U19741 (N_19741,N_16449,N_16515);
and U19742 (N_19742,N_16586,N_16521);
nor U19743 (N_19743,N_16952,N_16239);
and U19744 (N_19744,N_16938,N_16963);
and U19745 (N_19745,N_17739,N_16856);
or U19746 (N_19746,N_17718,N_16380);
nand U19747 (N_19747,N_16430,N_16859);
xnor U19748 (N_19748,N_17755,N_16879);
nor U19749 (N_19749,N_17468,N_16905);
nor U19750 (N_19750,N_17201,N_16224);
or U19751 (N_19751,N_17803,N_16587);
nor U19752 (N_19752,N_17691,N_17894);
nand U19753 (N_19753,N_16974,N_17812);
or U19754 (N_19754,N_16709,N_16209);
or U19755 (N_19755,N_16279,N_17353);
and U19756 (N_19756,N_16716,N_17217);
nor U19757 (N_19757,N_17403,N_16866);
and U19758 (N_19758,N_16968,N_16002);
or U19759 (N_19759,N_16287,N_17883);
nor U19760 (N_19760,N_16381,N_16407);
nor U19761 (N_19761,N_17212,N_17590);
nand U19762 (N_19762,N_16842,N_16712);
or U19763 (N_19763,N_17808,N_16653);
nor U19764 (N_19764,N_17456,N_16453);
nor U19765 (N_19765,N_16718,N_16517);
nand U19766 (N_19766,N_17530,N_16206);
or U19767 (N_19767,N_16275,N_17961);
or U19768 (N_19768,N_17849,N_17546);
and U19769 (N_19769,N_17978,N_17428);
and U19770 (N_19770,N_17329,N_17065);
nand U19771 (N_19771,N_16519,N_16387);
or U19772 (N_19772,N_16115,N_16398);
nand U19773 (N_19773,N_17401,N_17316);
or U19774 (N_19774,N_16703,N_17467);
nand U19775 (N_19775,N_16523,N_16285);
or U19776 (N_19776,N_17196,N_17811);
nor U19777 (N_19777,N_16954,N_16556);
or U19778 (N_19778,N_17012,N_16219);
nor U19779 (N_19779,N_17902,N_16440);
nand U19780 (N_19780,N_16505,N_17437);
nor U19781 (N_19781,N_17785,N_17004);
nand U19782 (N_19782,N_16573,N_16567);
or U19783 (N_19783,N_16581,N_17877);
nor U19784 (N_19784,N_16163,N_17250);
and U19785 (N_19785,N_16454,N_17393);
nand U19786 (N_19786,N_16059,N_16313);
nor U19787 (N_19787,N_16285,N_16244);
xnor U19788 (N_19788,N_16571,N_16812);
nand U19789 (N_19789,N_16476,N_16930);
nand U19790 (N_19790,N_16067,N_16615);
nor U19791 (N_19791,N_16271,N_17261);
or U19792 (N_19792,N_16120,N_17387);
and U19793 (N_19793,N_17410,N_16338);
xor U19794 (N_19794,N_16006,N_17249);
nor U19795 (N_19795,N_17970,N_17858);
and U19796 (N_19796,N_17202,N_16889);
or U19797 (N_19797,N_16914,N_16463);
or U19798 (N_19798,N_16936,N_17038);
and U19799 (N_19799,N_16395,N_17753);
and U19800 (N_19800,N_17648,N_16602);
or U19801 (N_19801,N_17567,N_16819);
and U19802 (N_19802,N_17260,N_17507);
nand U19803 (N_19803,N_16425,N_16159);
and U19804 (N_19804,N_17768,N_17252);
or U19805 (N_19805,N_16070,N_16515);
xor U19806 (N_19806,N_16336,N_17218);
nand U19807 (N_19807,N_17416,N_16662);
or U19808 (N_19808,N_16658,N_16639);
and U19809 (N_19809,N_16884,N_17315);
xnor U19810 (N_19810,N_16765,N_17493);
nand U19811 (N_19811,N_16679,N_17135);
or U19812 (N_19812,N_17202,N_16495);
nor U19813 (N_19813,N_16557,N_16152);
or U19814 (N_19814,N_16189,N_16098);
nand U19815 (N_19815,N_17472,N_16735);
xor U19816 (N_19816,N_16463,N_16102);
or U19817 (N_19817,N_16047,N_16084);
or U19818 (N_19818,N_17340,N_16441);
or U19819 (N_19819,N_17616,N_16168);
nor U19820 (N_19820,N_16127,N_17357);
and U19821 (N_19821,N_16434,N_17489);
nand U19822 (N_19822,N_17753,N_17226);
xor U19823 (N_19823,N_16377,N_17531);
or U19824 (N_19824,N_17887,N_16895);
or U19825 (N_19825,N_17523,N_16102);
nor U19826 (N_19826,N_16005,N_16908);
or U19827 (N_19827,N_17117,N_17384);
and U19828 (N_19828,N_16006,N_17724);
xor U19829 (N_19829,N_16628,N_16943);
nand U19830 (N_19830,N_17634,N_17899);
nand U19831 (N_19831,N_17479,N_17537);
nand U19832 (N_19832,N_16323,N_17824);
or U19833 (N_19833,N_17360,N_16403);
nand U19834 (N_19834,N_17049,N_17566);
nand U19835 (N_19835,N_17019,N_17688);
or U19836 (N_19836,N_17793,N_16364);
and U19837 (N_19837,N_16796,N_17446);
nor U19838 (N_19838,N_16284,N_16133);
nor U19839 (N_19839,N_16924,N_17375);
and U19840 (N_19840,N_16697,N_17567);
and U19841 (N_19841,N_17633,N_16692);
nor U19842 (N_19842,N_17983,N_16563);
and U19843 (N_19843,N_17167,N_17285);
and U19844 (N_19844,N_17635,N_17725);
and U19845 (N_19845,N_16525,N_16392);
nor U19846 (N_19846,N_17552,N_16652);
xor U19847 (N_19847,N_17892,N_16344);
or U19848 (N_19848,N_16808,N_16520);
or U19849 (N_19849,N_16206,N_16773);
xor U19850 (N_19850,N_16679,N_17767);
xor U19851 (N_19851,N_17151,N_17019);
nor U19852 (N_19852,N_17903,N_16092);
and U19853 (N_19853,N_17148,N_17240);
nand U19854 (N_19854,N_17119,N_16657);
xnor U19855 (N_19855,N_16504,N_17341);
xnor U19856 (N_19856,N_17936,N_17490);
nand U19857 (N_19857,N_16065,N_16669);
and U19858 (N_19858,N_16984,N_16650);
xnor U19859 (N_19859,N_16734,N_17824);
or U19860 (N_19860,N_16095,N_17243);
nor U19861 (N_19861,N_17044,N_17526);
xnor U19862 (N_19862,N_16865,N_17149);
xnor U19863 (N_19863,N_16042,N_17633);
nand U19864 (N_19864,N_17083,N_17470);
and U19865 (N_19865,N_17000,N_16162);
or U19866 (N_19866,N_17244,N_16122);
xnor U19867 (N_19867,N_16697,N_17790);
and U19868 (N_19868,N_16649,N_16849);
nor U19869 (N_19869,N_17545,N_16257);
or U19870 (N_19870,N_16049,N_17736);
nor U19871 (N_19871,N_16034,N_16386);
nand U19872 (N_19872,N_16227,N_16042);
nand U19873 (N_19873,N_17839,N_17714);
or U19874 (N_19874,N_16228,N_17629);
nand U19875 (N_19875,N_16727,N_17022);
and U19876 (N_19876,N_16996,N_17886);
and U19877 (N_19877,N_17930,N_16223);
and U19878 (N_19878,N_17725,N_17549);
nor U19879 (N_19879,N_16621,N_16790);
or U19880 (N_19880,N_17198,N_16546);
or U19881 (N_19881,N_17883,N_17938);
or U19882 (N_19882,N_16573,N_16615);
or U19883 (N_19883,N_17569,N_16749);
and U19884 (N_19884,N_17039,N_16209);
nand U19885 (N_19885,N_16510,N_17351);
or U19886 (N_19886,N_17372,N_16211);
and U19887 (N_19887,N_16293,N_16753);
nand U19888 (N_19888,N_16995,N_17458);
nor U19889 (N_19889,N_17752,N_16627);
and U19890 (N_19890,N_16499,N_16620);
and U19891 (N_19891,N_16842,N_16159);
and U19892 (N_19892,N_16129,N_16243);
nand U19893 (N_19893,N_17792,N_16437);
and U19894 (N_19894,N_16871,N_16122);
or U19895 (N_19895,N_16657,N_17822);
and U19896 (N_19896,N_16266,N_16664);
nor U19897 (N_19897,N_16735,N_17598);
and U19898 (N_19898,N_16417,N_17873);
and U19899 (N_19899,N_17170,N_17410);
and U19900 (N_19900,N_16664,N_16396);
nor U19901 (N_19901,N_16972,N_16371);
or U19902 (N_19902,N_16463,N_16669);
and U19903 (N_19903,N_17102,N_16485);
nand U19904 (N_19904,N_17789,N_17199);
or U19905 (N_19905,N_16657,N_17937);
nand U19906 (N_19906,N_16181,N_17141);
and U19907 (N_19907,N_17176,N_17438);
or U19908 (N_19908,N_17346,N_17782);
and U19909 (N_19909,N_17838,N_16430);
xor U19910 (N_19910,N_16319,N_17196);
or U19911 (N_19911,N_16568,N_16207);
xor U19912 (N_19912,N_16165,N_16947);
xnor U19913 (N_19913,N_16490,N_16445);
or U19914 (N_19914,N_17676,N_16863);
nor U19915 (N_19915,N_16001,N_17932);
or U19916 (N_19916,N_17172,N_16573);
nand U19917 (N_19917,N_16258,N_17456);
and U19918 (N_19918,N_17285,N_17923);
xnor U19919 (N_19919,N_16521,N_17161);
and U19920 (N_19920,N_16892,N_17685);
and U19921 (N_19921,N_16740,N_17612);
and U19922 (N_19922,N_17521,N_17724);
or U19923 (N_19923,N_17104,N_16646);
nor U19924 (N_19924,N_16378,N_16499);
nor U19925 (N_19925,N_16009,N_16146);
or U19926 (N_19926,N_16247,N_17771);
or U19927 (N_19927,N_17934,N_16549);
nand U19928 (N_19928,N_16959,N_16259);
nand U19929 (N_19929,N_16570,N_16947);
nand U19930 (N_19930,N_17103,N_17426);
nor U19931 (N_19931,N_17056,N_16848);
or U19932 (N_19932,N_17155,N_16631);
xnor U19933 (N_19933,N_17650,N_17384);
nand U19934 (N_19934,N_16251,N_17631);
or U19935 (N_19935,N_16570,N_16023);
or U19936 (N_19936,N_17336,N_16827);
and U19937 (N_19937,N_16209,N_17944);
nor U19938 (N_19938,N_17929,N_17916);
and U19939 (N_19939,N_16800,N_17768);
or U19940 (N_19940,N_16457,N_17289);
nor U19941 (N_19941,N_17705,N_17850);
and U19942 (N_19942,N_16970,N_16539);
nor U19943 (N_19943,N_16421,N_17653);
nor U19944 (N_19944,N_16456,N_16529);
nand U19945 (N_19945,N_17818,N_17138);
or U19946 (N_19946,N_17028,N_17939);
nand U19947 (N_19947,N_16027,N_17965);
and U19948 (N_19948,N_16056,N_16641);
or U19949 (N_19949,N_16108,N_16430);
nor U19950 (N_19950,N_16062,N_17498);
and U19951 (N_19951,N_17189,N_16621);
or U19952 (N_19952,N_17675,N_16213);
nor U19953 (N_19953,N_17179,N_16975);
nor U19954 (N_19954,N_16694,N_16013);
or U19955 (N_19955,N_17646,N_16763);
or U19956 (N_19956,N_17125,N_17288);
nor U19957 (N_19957,N_16677,N_16020);
and U19958 (N_19958,N_16917,N_17118);
and U19959 (N_19959,N_16937,N_16350);
and U19960 (N_19960,N_16968,N_16167);
or U19961 (N_19961,N_17472,N_16353);
and U19962 (N_19962,N_16066,N_17371);
nor U19963 (N_19963,N_17283,N_16190);
and U19964 (N_19964,N_16313,N_17563);
xnor U19965 (N_19965,N_17137,N_16674);
nand U19966 (N_19966,N_17829,N_17774);
xnor U19967 (N_19967,N_16033,N_17427);
and U19968 (N_19968,N_17238,N_16736);
or U19969 (N_19969,N_16146,N_16560);
nand U19970 (N_19970,N_16302,N_16345);
and U19971 (N_19971,N_17411,N_16746);
nand U19972 (N_19972,N_16582,N_16579);
or U19973 (N_19973,N_17470,N_17126);
nor U19974 (N_19974,N_16604,N_17458);
and U19975 (N_19975,N_16730,N_16600);
or U19976 (N_19976,N_17770,N_17283);
nand U19977 (N_19977,N_17950,N_16237);
and U19978 (N_19978,N_17394,N_16897);
nand U19979 (N_19979,N_17305,N_17582);
and U19980 (N_19980,N_17352,N_16420);
nand U19981 (N_19981,N_16508,N_16406);
nor U19982 (N_19982,N_16667,N_16811);
nor U19983 (N_19983,N_17350,N_16597);
xor U19984 (N_19984,N_16077,N_16436);
nor U19985 (N_19985,N_16304,N_16611);
and U19986 (N_19986,N_17057,N_16195);
nor U19987 (N_19987,N_17113,N_16368);
and U19988 (N_19988,N_17847,N_16835);
or U19989 (N_19989,N_17769,N_16404);
or U19990 (N_19990,N_17347,N_17105);
nand U19991 (N_19991,N_16031,N_17855);
nand U19992 (N_19992,N_16155,N_17913);
nand U19993 (N_19993,N_17687,N_17604);
and U19994 (N_19994,N_16314,N_17235);
or U19995 (N_19995,N_16950,N_17578);
and U19996 (N_19996,N_17596,N_16635);
and U19997 (N_19997,N_17707,N_16251);
or U19998 (N_19998,N_17031,N_17944);
or U19999 (N_19999,N_17647,N_17344);
and UO_0 (O_0,N_19471,N_19692);
nand UO_1 (O_1,N_18207,N_19448);
nor UO_2 (O_2,N_18395,N_19890);
nor UO_3 (O_3,N_19341,N_18143);
xor UO_4 (O_4,N_18345,N_19667);
nor UO_5 (O_5,N_19846,N_19856);
or UO_6 (O_6,N_18217,N_18170);
and UO_7 (O_7,N_19336,N_19808);
and UO_8 (O_8,N_19902,N_19151);
nor UO_9 (O_9,N_18500,N_18433);
and UO_10 (O_10,N_18499,N_18942);
or UO_11 (O_11,N_19748,N_19609);
nand UO_12 (O_12,N_18090,N_19826);
and UO_13 (O_13,N_19941,N_18921);
and UO_14 (O_14,N_18107,N_19348);
or UO_15 (O_15,N_19176,N_19604);
or UO_16 (O_16,N_19555,N_18900);
or UO_17 (O_17,N_18160,N_19451);
nand UO_18 (O_18,N_18163,N_18834);
nor UO_19 (O_19,N_18463,N_18864);
nor UO_20 (O_20,N_18050,N_18914);
or UO_21 (O_21,N_18064,N_19861);
nor UO_22 (O_22,N_18047,N_18669);
xnor UO_23 (O_23,N_19293,N_18147);
nand UO_24 (O_24,N_19880,N_19346);
and UO_25 (O_25,N_18387,N_18067);
and UO_26 (O_26,N_18861,N_18294);
and UO_27 (O_27,N_18762,N_18338);
nor UO_28 (O_28,N_19875,N_18240);
or UO_29 (O_29,N_18645,N_19558);
nand UO_30 (O_30,N_18046,N_18181);
and UO_31 (O_31,N_19047,N_18928);
nor UO_32 (O_32,N_18597,N_18990);
nand UO_33 (O_33,N_18568,N_18326);
nor UO_34 (O_34,N_19574,N_18808);
nor UO_35 (O_35,N_18201,N_18825);
xnor UO_36 (O_36,N_19459,N_19479);
and UO_37 (O_37,N_18048,N_19515);
and UO_38 (O_38,N_18954,N_19951);
nand UO_39 (O_39,N_19911,N_18153);
nor UO_40 (O_40,N_18709,N_19076);
nor UO_41 (O_41,N_18906,N_18695);
nor UO_42 (O_42,N_19419,N_18770);
or UO_43 (O_43,N_18646,N_18078);
nor UO_44 (O_44,N_19651,N_18394);
nor UO_45 (O_45,N_18037,N_18949);
or UO_46 (O_46,N_19550,N_19921);
and UO_47 (O_47,N_19625,N_19982);
nor UO_48 (O_48,N_19843,N_19330);
nor UO_49 (O_49,N_18295,N_19088);
nand UO_50 (O_50,N_19691,N_18741);
or UO_51 (O_51,N_18927,N_19187);
and UO_52 (O_52,N_18104,N_18337);
and UO_53 (O_53,N_19876,N_19791);
nand UO_54 (O_54,N_19482,N_19647);
nand UO_55 (O_55,N_19792,N_19731);
nor UO_56 (O_56,N_18472,N_19567);
and UO_57 (O_57,N_19130,N_18800);
or UO_58 (O_58,N_18363,N_19732);
nor UO_59 (O_59,N_18149,N_18911);
nand UO_60 (O_60,N_19081,N_19660);
and UO_61 (O_61,N_18456,N_19623);
nor UO_62 (O_62,N_18358,N_19458);
xnor UO_63 (O_63,N_19372,N_18252);
and UO_64 (O_64,N_18847,N_19117);
and UO_65 (O_65,N_19620,N_19136);
and UO_66 (O_66,N_18120,N_19583);
or UO_67 (O_67,N_19619,N_18421);
nand UO_68 (O_68,N_19484,N_18154);
or UO_69 (O_69,N_18397,N_18029);
nor UO_70 (O_70,N_19265,N_18871);
nor UO_71 (O_71,N_19971,N_19444);
nor UO_72 (O_72,N_18944,N_18846);
or UO_73 (O_73,N_19377,N_18687);
and UO_74 (O_74,N_19927,N_18359);
nor UO_75 (O_75,N_18164,N_19290);
and UO_76 (O_76,N_18373,N_19492);
nor UO_77 (O_77,N_18905,N_19511);
and UO_78 (O_78,N_19554,N_18309);
or UO_79 (O_79,N_19184,N_18554);
or UO_80 (O_80,N_18842,N_18079);
and UO_81 (O_81,N_19154,N_19928);
nand UO_82 (O_82,N_19199,N_19464);
nand UO_83 (O_83,N_19203,N_19235);
nor UO_84 (O_84,N_19910,N_18671);
or UO_85 (O_85,N_18253,N_19282);
or UO_86 (O_86,N_19475,N_19469);
and UO_87 (O_87,N_18276,N_18857);
xor UO_88 (O_88,N_19763,N_18895);
and UO_89 (O_89,N_19103,N_18013);
nand UO_90 (O_90,N_19837,N_18100);
or UO_91 (O_91,N_19391,N_18109);
nor UO_92 (O_92,N_19592,N_19612);
or UO_93 (O_93,N_19367,N_19799);
and UO_94 (O_94,N_19283,N_18964);
or UO_95 (O_95,N_19460,N_19998);
and UO_96 (O_96,N_19153,N_18971);
nor UO_97 (O_97,N_19305,N_18015);
nor UO_98 (O_98,N_19593,N_18083);
nand UO_99 (O_99,N_18166,N_19828);
nand UO_100 (O_100,N_18859,N_19576);
xor UO_101 (O_101,N_18904,N_18427);
or UO_102 (O_102,N_19427,N_18116);
and UO_103 (O_103,N_18579,N_19406);
or UO_104 (O_104,N_19727,N_19288);
and UO_105 (O_105,N_18182,N_18136);
nor UO_106 (O_106,N_19805,N_18784);
and UO_107 (O_107,N_19543,N_19125);
and UO_108 (O_108,N_19237,N_18729);
nand UO_109 (O_109,N_18768,N_18250);
nor UO_110 (O_110,N_19708,N_19816);
nand UO_111 (O_111,N_19734,N_19559);
nor UO_112 (O_112,N_18619,N_18888);
and UO_113 (O_113,N_18993,N_19466);
nor UO_114 (O_114,N_19289,N_18551);
nand UO_115 (O_115,N_18756,N_18573);
or UO_116 (O_116,N_19128,N_19725);
or UO_117 (O_117,N_18916,N_19110);
nor UO_118 (O_118,N_18113,N_18165);
and UO_119 (O_119,N_18434,N_19663);
nand UO_120 (O_120,N_19895,N_18214);
or UO_121 (O_121,N_19924,N_19967);
nand UO_122 (O_122,N_19877,N_18161);
nand UO_123 (O_123,N_18608,N_18103);
xnor UO_124 (O_124,N_18985,N_19312);
or UO_125 (O_125,N_18706,N_19353);
nor UO_126 (O_126,N_19859,N_18351);
xnor UO_127 (O_127,N_18522,N_19785);
nor UO_128 (O_128,N_19741,N_19351);
nand UO_129 (O_129,N_18416,N_19032);
or UO_130 (O_130,N_19066,N_19955);
and UO_131 (O_131,N_18679,N_19950);
or UO_132 (O_132,N_19806,N_19143);
nand UO_133 (O_133,N_19292,N_19820);
nand UO_134 (O_134,N_18076,N_18091);
nor UO_135 (O_135,N_18736,N_18773);
nand UO_136 (O_136,N_18099,N_18431);
nand UO_137 (O_137,N_19487,N_18176);
nand UO_138 (O_138,N_19997,N_19425);
and UO_139 (O_139,N_19524,N_18465);
and UO_140 (O_140,N_19940,N_18391);
and UO_141 (O_141,N_19468,N_18393);
or UO_142 (O_142,N_18682,N_18313);
and UO_143 (O_143,N_19380,N_18966);
nand UO_144 (O_144,N_19481,N_19229);
nand UO_145 (O_145,N_19914,N_19214);
and UO_146 (O_146,N_18915,N_18887);
nor UO_147 (O_147,N_19578,N_19362);
nor UO_148 (O_148,N_18812,N_18383);
or UO_149 (O_149,N_18350,N_19019);
xor UO_150 (O_150,N_19234,N_19587);
nand UO_151 (O_151,N_19139,N_19095);
or UO_152 (O_152,N_19707,N_19122);
or UO_153 (O_153,N_18901,N_18260);
nand UO_154 (O_154,N_18066,N_19375);
or UO_155 (O_155,N_18772,N_19602);
or UO_156 (O_156,N_19839,N_18005);
or UO_157 (O_157,N_19302,N_18848);
nand UO_158 (O_158,N_19945,N_19414);
nand UO_159 (O_159,N_18323,N_18955);
or UO_160 (O_160,N_19886,N_19493);
or UO_161 (O_161,N_18519,N_18419);
nor UO_162 (O_162,N_19055,N_19190);
nor UO_163 (O_163,N_18854,N_18200);
and UO_164 (O_164,N_19992,N_19486);
nor UO_165 (O_165,N_18445,N_18024);
and UO_166 (O_166,N_18304,N_18508);
nand UO_167 (O_167,N_19022,N_19938);
and UO_168 (O_168,N_18845,N_19831);
nor UO_169 (O_169,N_18466,N_18407);
and UO_170 (O_170,N_18012,N_18852);
and UO_171 (O_171,N_18720,N_18585);
nand UO_172 (O_172,N_18035,N_18697);
and UO_173 (O_173,N_19590,N_19909);
and UO_174 (O_174,N_18259,N_18491);
xnor UO_175 (O_175,N_18725,N_19401);
or UO_176 (O_176,N_19495,N_18837);
and UO_177 (O_177,N_19571,N_18674);
and UO_178 (O_178,N_19287,N_18584);
xnor UO_179 (O_179,N_18867,N_19045);
or UO_180 (O_180,N_19108,N_19607);
or UO_181 (O_181,N_18953,N_18685);
nand UO_182 (O_182,N_19106,N_19853);
nand UO_183 (O_183,N_18603,N_19254);
and UO_184 (O_184,N_19112,N_18467);
nand UO_185 (O_185,N_18544,N_18839);
nor UO_186 (O_186,N_19294,N_19390);
or UO_187 (O_187,N_18251,N_18778);
nand UO_188 (O_188,N_18622,N_18931);
nor UO_189 (O_189,N_19788,N_18314);
and UO_190 (O_190,N_19251,N_19855);
nor UO_191 (O_191,N_19564,N_18275);
nor UO_192 (O_192,N_18636,N_18560);
or UO_193 (O_193,N_18436,N_19669);
nor UO_194 (O_194,N_18423,N_19327);
or UO_195 (O_195,N_19304,N_19916);
nor UO_196 (O_196,N_18926,N_18368);
or UO_197 (O_197,N_18643,N_19256);
nor UO_198 (O_198,N_18405,N_19407);
or UO_199 (O_199,N_18833,N_19243);
and UO_200 (O_200,N_19438,N_18001);
xnor UO_201 (O_201,N_18714,N_19031);
nor UO_202 (O_202,N_18771,N_18678);
and UO_203 (O_203,N_18936,N_18530);
nor UO_204 (O_204,N_18607,N_19894);
nand UO_205 (O_205,N_18257,N_18219);
and UO_206 (O_206,N_19197,N_18003);
or UO_207 (O_207,N_18683,N_18392);
and UO_208 (O_208,N_18339,N_19422);
nor UO_209 (O_209,N_19568,N_19092);
or UO_210 (O_210,N_19617,N_19522);
and UO_211 (O_211,N_18045,N_19907);
nand UO_212 (O_212,N_19321,N_19549);
nor UO_213 (O_213,N_19978,N_18305);
nand UO_214 (O_214,N_19347,N_18513);
nor UO_215 (O_215,N_18101,N_19067);
or UO_216 (O_216,N_19518,N_18095);
nor UO_217 (O_217,N_18520,N_18177);
or UO_218 (O_218,N_18476,N_19838);
nand UO_219 (O_219,N_18733,N_18468);
nand UO_220 (O_220,N_19309,N_19827);
and UO_221 (O_221,N_19675,N_19646);
nor UO_222 (O_222,N_18816,N_18269);
and UO_223 (O_223,N_18475,N_18000);
nand UO_224 (O_224,N_18142,N_18652);
nor UO_225 (O_225,N_18981,N_19610);
nor UO_226 (O_226,N_19316,N_18899);
nor UO_227 (O_227,N_19400,N_18016);
nor UO_228 (O_228,N_18370,N_18810);
nor UO_229 (O_229,N_19410,N_18195);
nor UO_230 (O_230,N_18289,N_18126);
or UO_231 (O_231,N_18092,N_19996);
nand UO_232 (O_232,N_19478,N_19324);
nand UO_233 (O_233,N_19714,N_18247);
nor UO_234 (O_234,N_18032,N_19948);
or UO_235 (O_235,N_19929,N_19865);
nand UO_236 (O_236,N_18183,N_19424);
or UO_237 (O_237,N_19453,N_19360);
or UO_238 (O_238,N_18737,N_19537);
nand UO_239 (O_239,N_18922,N_19934);
and UO_240 (O_240,N_19253,N_19188);
nor UO_241 (O_241,N_19250,N_19171);
and UO_242 (O_242,N_18105,N_19811);
and UO_243 (O_243,N_18420,N_18742);
and UO_244 (O_244,N_18938,N_18794);
or UO_245 (O_245,N_19120,N_18543);
nor UO_246 (O_246,N_18084,N_18357);
and UO_247 (O_247,N_19392,N_18451);
and UO_248 (O_248,N_19278,N_19599);
and UO_249 (O_249,N_18157,N_18186);
or UO_250 (O_250,N_18399,N_19769);
or UO_251 (O_251,N_19442,N_19363);
and UO_252 (O_252,N_19228,N_19064);
nand UO_253 (O_253,N_19965,N_19946);
or UO_254 (O_254,N_19025,N_19246);
or UO_255 (O_255,N_18849,N_19848);
or UO_256 (O_256,N_18902,N_19091);
xor UO_257 (O_257,N_19062,N_18447);
xor UO_258 (O_258,N_18462,N_18667);
nand UO_259 (O_259,N_18984,N_19926);
xor UO_260 (O_260,N_18612,N_18583);
and UO_261 (O_261,N_19193,N_19157);
nor UO_262 (O_262,N_19519,N_19913);
nand UO_263 (O_263,N_19005,N_18759);
xor UO_264 (O_264,N_19661,N_19042);
or UO_265 (O_265,N_18965,N_18750);
nor UO_266 (O_266,N_18972,N_19648);
or UO_267 (O_267,N_19465,N_19535);
xor UO_268 (O_268,N_19654,N_19206);
and UO_269 (O_269,N_19695,N_19381);
and UO_270 (O_270,N_19098,N_19701);
or UO_271 (O_271,N_18366,N_18209);
or UO_272 (O_272,N_19795,N_18141);
xor UO_273 (O_273,N_18482,N_19009);
and UO_274 (O_274,N_19758,N_18428);
and UO_275 (O_275,N_18448,N_19165);
nor UO_276 (O_276,N_18497,N_18486);
nand UO_277 (O_277,N_19298,N_19454);
nor UO_278 (O_278,N_19595,N_19566);
xor UO_279 (O_279,N_19631,N_18234);
nand UO_280 (O_280,N_18912,N_19908);
nand UO_281 (O_281,N_19705,N_18469);
and UO_282 (O_282,N_19455,N_18115);
nand UO_283 (O_283,N_18571,N_18702);
or UO_284 (O_284,N_19674,N_19185);
nand UO_285 (O_285,N_19709,N_19704);
and UO_286 (O_286,N_19656,N_18039);
and UO_287 (O_287,N_19447,N_18461);
nor UO_288 (O_288,N_19477,N_19517);
xnor UO_289 (O_289,N_18668,N_19494);
nor UO_290 (O_290,N_19783,N_18995);
or UO_291 (O_291,N_19553,N_19061);
and UO_292 (O_292,N_18121,N_18131);
or UO_293 (O_293,N_19205,N_19776);
xnor UO_294 (O_294,N_19010,N_18306);
nand UO_295 (O_295,N_18701,N_18268);
nand UO_296 (O_296,N_18509,N_18470);
nand UO_297 (O_297,N_19984,N_18376);
xor UO_298 (O_298,N_18510,N_18890);
or UO_299 (O_299,N_19762,N_18892);
and UO_300 (O_300,N_19462,N_18650);
or UO_301 (O_301,N_19684,N_18030);
and UO_302 (O_302,N_18492,N_18239);
and UO_303 (O_303,N_19624,N_19408);
xor UO_304 (O_304,N_18820,N_18069);
or UO_305 (O_305,N_18686,N_19717);
nand UO_306 (O_306,N_19833,N_18072);
and UO_307 (O_307,N_18460,N_18379);
nor UO_308 (O_308,N_19233,N_18865);
nand UO_309 (O_309,N_19129,N_18213);
nor UO_310 (O_310,N_19020,N_18992);
and UO_311 (O_311,N_19079,N_19993);
nand UO_312 (O_312,N_18190,N_19276);
nor UO_313 (O_313,N_18644,N_19073);
and UO_314 (O_314,N_18883,N_19664);
or UO_315 (O_315,N_19071,N_18249);
or UO_316 (O_316,N_19150,N_19085);
nand UO_317 (O_317,N_18442,N_19166);
nor UO_318 (O_318,N_19627,N_19178);
xnor UO_319 (O_319,N_19683,N_19087);
and UO_320 (O_320,N_18384,N_18137);
nor UO_321 (O_321,N_19207,N_19093);
nor UO_322 (O_322,N_19029,N_19077);
xnor UO_323 (O_323,N_18653,N_19249);
nor UO_324 (O_324,N_19747,N_19300);
nand UO_325 (O_325,N_19140,N_18606);
nand UO_326 (O_326,N_19480,N_18353);
and UO_327 (O_327,N_19680,N_18982);
and UO_328 (O_328,N_18027,N_18707);
xor UO_329 (O_329,N_18792,N_19258);
nor UO_330 (O_330,N_19641,N_19275);
nor UO_331 (O_331,N_19433,N_18605);
and UO_332 (O_332,N_18025,N_18506);
and UO_333 (O_333,N_19794,N_18630);
nor UO_334 (O_334,N_19121,N_19474);
and UO_335 (O_335,N_18986,N_19441);
and UO_336 (O_336,N_18098,N_18588);
nand UO_337 (O_337,N_18557,N_19114);
nand UO_338 (O_338,N_18390,N_19883);
nand UO_339 (O_339,N_19919,N_18380);
and UO_340 (O_340,N_19039,N_18057);
nor UO_341 (O_341,N_18807,N_19461);
nand UO_342 (O_342,N_18913,N_18563);
xnor UO_343 (O_343,N_19803,N_19393);
or UO_344 (O_344,N_18934,N_18324);
xor UO_345 (O_345,N_19182,N_19232);
xor UO_346 (O_346,N_19196,N_18272);
and UO_347 (O_347,N_18429,N_19416);
nor UO_348 (O_348,N_18377,N_19180);
or UO_349 (O_349,N_18385,N_18087);
xor UO_350 (O_350,N_19923,N_19386);
or UO_351 (O_351,N_18918,N_18699);
nor UO_352 (O_352,N_18657,N_19516);
or UO_353 (O_353,N_19509,N_18220);
and UO_354 (O_354,N_18757,N_18321);
nand UO_355 (O_355,N_19850,N_19751);
or UO_356 (O_356,N_18322,N_18375);
xor UO_357 (O_357,N_19937,N_18937);
nand UO_358 (O_358,N_18724,N_18818);
or UO_359 (O_359,N_18531,N_18626);
xor UO_360 (O_360,N_19070,N_19152);
or UO_361 (O_361,N_18286,N_19622);
nor UO_362 (O_362,N_18415,N_19297);
nand UO_363 (O_363,N_18263,N_19529);
or UO_364 (O_364,N_19847,N_19450);
or UO_365 (O_365,N_18396,N_19616);
and UO_366 (O_366,N_19059,N_19954);
or UO_367 (O_367,N_18718,N_18962);
nand UO_368 (O_368,N_18340,N_19815);
nand UO_369 (O_369,N_19018,N_18941);
xor UO_370 (O_370,N_18320,N_18801);
or UO_371 (O_371,N_19830,N_19867);
and UO_372 (O_372,N_18178,N_18018);
nand UO_373 (O_373,N_19134,N_19215);
xnor UO_374 (O_374,N_19614,N_19065);
xnor UO_375 (O_375,N_19819,N_18226);
or UO_376 (O_376,N_19696,N_18863);
nor UO_377 (O_377,N_19635,N_18829);
or UO_378 (O_378,N_18898,N_18404);
and UO_379 (O_379,N_18593,N_19693);
or UO_380 (O_380,N_18655,N_18400);
nand UO_381 (O_381,N_19063,N_18071);
or UO_382 (O_382,N_18331,N_19269);
nor UO_383 (O_383,N_18617,N_19995);
and UO_384 (O_384,N_18139,N_19716);
or UO_385 (O_385,N_18872,N_18961);
or UO_386 (O_386,N_19456,N_19655);
and UO_387 (O_387,N_19262,N_19817);
nand UO_388 (O_388,N_19645,N_18075);
or UO_389 (O_389,N_19099,N_19713);
nor UO_390 (O_390,N_19457,N_19037);
nor UO_391 (O_391,N_18978,N_18490);
nand UO_392 (O_392,N_19733,N_18145);
and UO_393 (O_393,N_18274,N_19024);
nor UO_394 (O_394,N_18374,N_18204);
nand UO_395 (O_395,N_19502,N_18049);
nor UO_396 (O_396,N_18664,N_19332);
xor UO_397 (O_397,N_18805,N_18424);
and UO_398 (O_398,N_19813,N_18019);
nand UO_399 (O_399,N_18059,N_19962);
nand UO_400 (O_400,N_18281,N_18279);
nand UO_401 (O_401,N_18208,N_19183);
and UO_402 (O_402,N_18346,N_19489);
and UO_403 (O_403,N_18894,N_18273);
nand UO_404 (O_404,N_19968,N_18577);
nor UO_405 (O_405,N_19303,N_19488);
xor UO_406 (O_406,N_19740,N_19672);
nor UO_407 (O_407,N_19739,N_19328);
or UO_408 (O_408,N_18923,N_19584);
nor UO_409 (O_409,N_18648,N_18766);
and UO_410 (O_410,N_19086,N_19679);
or UO_411 (O_411,N_19649,N_18717);
nor UO_412 (O_412,N_19871,N_18360);
and UO_413 (O_413,N_19643,N_19580);
or UO_414 (O_414,N_18719,N_18782);
or UO_415 (O_415,N_19318,N_19706);
nand UO_416 (O_416,N_18675,N_18746);
and UO_417 (O_417,N_19560,N_18793);
nor UO_418 (O_418,N_18844,N_18547);
or UO_419 (O_419,N_19389,N_18879);
and UO_420 (O_420,N_18205,N_18457);
and UO_421 (O_421,N_19331,N_19286);
nor UO_422 (O_422,N_18666,N_19111);
and UO_423 (O_423,N_18110,N_18658);
xor UO_424 (O_424,N_19131,N_19531);
nor UO_425 (O_425,N_19896,N_18093);
or UO_426 (O_426,N_19893,N_18056);
and UO_427 (O_427,N_19688,N_18033);
nor UO_428 (O_428,N_19082,N_18372);
nor UO_429 (O_429,N_19388,N_19026);
nand UO_430 (O_430,N_19023,N_18038);
or UO_431 (O_431,N_19075,N_18525);
xor UO_432 (O_432,N_19510,N_19078);
or UO_433 (O_433,N_19825,N_18540);
and UO_434 (O_434,N_19223,N_18378);
xor UO_435 (O_435,N_18173,N_19528);
nor UO_436 (O_436,N_18505,N_18999);
and UO_437 (O_437,N_18007,N_18712);
nor UO_438 (O_438,N_19809,N_18210);
nand UO_439 (O_439,N_19439,N_18227);
nor UO_440 (O_440,N_18527,N_18755);
or UO_441 (O_441,N_19116,N_19930);
xnor UO_442 (O_442,N_18300,N_19015);
nor UO_443 (O_443,N_18485,N_19943);
nand UO_444 (O_444,N_18187,N_18172);
or UO_445 (O_445,N_18053,N_18297);
nor UO_446 (O_446,N_19273,N_18748);
nor UO_447 (O_447,N_19775,N_18809);
xor UO_448 (O_448,N_18371,N_19426);
nor UO_449 (O_449,N_19473,N_18271);
or UO_450 (O_450,N_18691,N_19773);
nand UO_451 (O_451,N_19359,N_18052);
nor UO_452 (O_452,N_18073,N_19857);
nand UO_453 (O_453,N_18601,N_18973);
or UO_454 (O_454,N_18988,N_18672);
nand UO_455 (O_455,N_19854,N_19244);
nor UO_456 (O_456,N_18815,N_18814);
nand UO_457 (O_457,N_18721,N_19581);
or UO_458 (O_458,N_18327,N_19350);
and UO_459 (O_459,N_19842,N_18361);
nand UO_460 (O_460,N_19284,N_19490);
and UO_461 (O_461,N_19659,N_19365);
and UO_462 (O_462,N_19034,N_19906);
nand UO_463 (O_463,N_19142,N_19340);
or UO_464 (O_464,N_18040,N_19772);
nor UO_465 (O_465,N_18676,N_19508);
or UO_466 (O_466,N_19311,N_19217);
or UO_467 (O_467,N_18493,N_18696);
or UO_468 (O_468,N_18502,N_19296);
xor UO_469 (O_469,N_18343,N_19821);
or UO_470 (O_470,N_18088,N_18726);
nand UO_471 (O_471,N_18501,N_19004);
nor UO_472 (O_472,N_18663,N_18111);
or UO_473 (O_473,N_18488,N_18980);
nor UO_474 (O_474,N_18882,N_19851);
or UO_475 (O_475,N_19405,N_18118);
nand UO_476 (O_476,N_18444,N_19252);
and UO_477 (O_477,N_18947,N_19885);
or UO_478 (O_478,N_19124,N_19089);
xnor UO_479 (O_479,N_19718,N_19200);
xor UO_480 (O_480,N_19366,N_18489);
and UO_481 (O_481,N_18715,N_19102);
xnor UO_482 (O_482,N_19858,N_18237);
nand UO_483 (O_483,N_19991,N_19172);
or UO_484 (O_484,N_18797,N_19383);
nand UO_485 (O_485,N_19723,N_18189);
or UO_486 (O_486,N_18117,N_19133);
nand UO_487 (O_487,N_19011,N_18997);
nand UO_488 (O_488,N_19364,N_18575);
and UO_489 (O_489,N_18856,N_18945);
and UO_490 (O_490,N_18296,N_19272);
xnor UO_491 (O_491,N_18564,N_18957);
and UO_492 (O_492,N_19887,N_18449);
nor UO_493 (O_493,N_19814,N_19526);
xnor UO_494 (O_494,N_18920,N_19041);
nor UO_495 (O_495,N_18680,N_19323);
and UO_496 (O_496,N_18783,N_19900);
nor UO_497 (O_497,N_18108,N_18775);
and UO_498 (O_498,N_19467,N_18621);
nand UO_499 (O_499,N_18511,N_19137);
nand UO_500 (O_500,N_18751,N_18452);
or UO_501 (O_501,N_18140,N_19548);
or UO_502 (O_502,N_18526,N_19744);
xnor UO_503 (O_503,N_18963,N_19192);
nor UO_504 (O_504,N_19306,N_19983);
and UO_505 (O_505,N_19742,N_18179);
nor UO_506 (O_506,N_18823,N_19356);
and UO_507 (O_507,N_18261,N_19449);
or UO_508 (O_508,N_19335,N_19376);
nor UO_509 (O_509,N_18412,N_18341);
or UO_510 (O_510,N_18329,N_19325);
nand UO_511 (O_511,N_19682,N_19191);
or UO_512 (O_512,N_18684,N_19613);
nand UO_513 (O_513,N_18730,N_19822);
and UO_514 (O_514,N_18020,N_18749);
or UO_515 (O_515,N_19195,N_18132);
xnor UO_516 (O_516,N_18285,N_19852);
xnor UO_517 (O_517,N_18570,N_19677);
nand UO_518 (O_518,N_18512,N_18763);
and UO_519 (O_519,N_18362,N_18026);
nand UO_520 (O_520,N_19503,N_18352);
or UO_521 (O_521,N_19644,N_19586);
and UO_522 (O_522,N_18835,N_19936);
nand UO_523 (O_523,N_19337,N_18194);
nor UO_524 (O_524,N_18665,N_18532);
nor UO_525 (O_525,N_19209,N_18009);
and UO_526 (O_526,N_18168,N_19634);
nor UO_527 (O_527,N_18828,N_18058);
xnor UO_528 (O_528,N_18455,N_18097);
nand UO_529 (O_529,N_18060,N_19226);
and UO_530 (O_530,N_18536,N_19245);
nand UO_531 (O_531,N_19764,N_19957);
xnor UO_532 (O_532,N_18910,N_18336);
xor UO_533 (O_533,N_19428,N_19033);
and UO_534 (O_534,N_18175,N_18481);
and UO_535 (O_535,N_18446,N_19002);
nor UO_536 (O_536,N_18077,N_18158);
nand UO_537 (O_537,N_19329,N_19437);
or UO_538 (O_538,N_18125,N_19212);
nor UO_539 (O_539,N_19729,N_18803);
xnor UO_540 (O_540,N_18382,N_18515);
nand UO_541 (O_541,N_19175,N_19975);
or UO_542 (O_542,N_19291,N_19673);
or UO_543 (O_543,N_19790,N_18318);
and UO_544 (O_544,N_19000,N_19241);
or UO_545 (O_545,N_18146,N_18080);
nand UO_546 (O_546,N_18881,N_19720);
or UO_547 (O_547,N_19499,N_18230);
or UO_548 (O_548,N_18698,N_18851);
and UO_549 (O_549,N_19903,N_18787);
and UO_550 (O_550,N_18364,N_19638);
nor UO_551 (O_551,N_18708,N_18681);
nand UO_552 (O_552,N_19219,N_18550);
nand UO_553 (O_553,N_18312,N_19615);
xnor UO_554 (O_554,N_18191,N_19096);
or UO_555 (O_555,N_19765,N_19657);
nand UO_556 (O_556,N_18723,N_18595);
or UO_557 (O_557,N_19403,N_19959);
nand UO_558 (O_558,N_18600,N_19892);
and UO_559 (O_559,N_18283,N_18114);
xor UO_560 (O_560,N_18123,N_19710);
nand UO_561 (O_561,N_19618,N_18255);
and UO_562 (O_562,N_19213,N_18441);
nand UO_563 (O_563,N_19897,N_19104);
or UO_564 (O_564,N_19561,N_18477);
nor UO_565 (O_565,N_18558,N_19686);
or UO_566 (O_566,N_19222,N_18832);
nand UO_567 (O_567,N_19642,N_19504);
or UO_568 (O_568,N_19307,N_19653);
nand UO_569 (O_569,N_18034,N_18974);
nor UO_570 (O_570,N_19712,N_19774);
nand UO_571 (O_571,N_19382,N_18602);
or UO_572 (O_572,N_18632,N_19281);
and UO_573 (O_573,N_19202,N_18781);
and UO_574 (O_574,N_19904,N_19038);
nor UO_575 (O_575,N_18537,N_19242);
and UO_576 (O_576,N_18553,N_18642);
or UO_577 (O_577,N_19247,N_19231);
nand UO_578 (O_578,N_18827,N_18909);
nand UO_579 (O_579,N_19141,N_18689);
or UO_580 (O_580,N_18414,N_18552);
nand UO_581 (O_581,N_18156,N_19148);
nand UO_582 (O_582,N_18656,N_19752);
nand UO_583 (O_583,N_19514,N_19779);
and UO_584 (O_584,N_19849,N_18635);
and UO_585 (O_585,N_18754,N_19161);
xor UO_586 (O_586,N_18991,N_18785);
nand UO_587 (O_587,N_19628,N_19429);
and UO_588 (O_588,N_18555,N_18235);
or UO_589 (O_589,N_18979,N_19882);
nor UO_590 (O_590,N_19563,N_19314);
and UO_591 (O_591,N_19520,N_19884);
or UO_592 (O_592,N_18041,N_19546);
or UO_593 (O_593,N_19582,N_18740);
nand UO_594 (O_594,N_18598,N_18494);
nor UO_595 (O_595,N_19703,N_18567);
nor UO_596 (O_596,N_18507,N_18349);
nand UO_597 (O_597,N_19046,N_19626);
nor UO_598 (O_598,N_19387,N_19260);
or UO_599 (O_599,N_18229,N_19976);
nand UO_600 (O_600,N_19844,N_19698);
or UO_601 (O_601,N_19052,N_19804);
or UO_602 (O_602,N_19413,N_19016);
nor UO_603 (O_603,N_19523,N_19221);
xnor UO_604 (O_604,N_19721,N_18504);
or UO_605 (O_605,N_19452,N_19497);
nor UO_606 (O_606,N_18796,N_18514);
xor UO_607 (O_607,N_18948,N_19915);
xor UO_608 (O_608,N_19204,N_18458);
nor UO_609 (O_609,N_18054,N_18549);
nand UO_610 (O_610,N_19700,N_18315);
nor UO_611 (O_611,N_18211,N_19953);
and UO_612 (O_612,N_18188,N_18703);
and UO_613 (O_613,N_19263,N_18243);
nor UO_614 (O_614,N_18869,N_19920);
xor UO_615 (O_615,N_18638,N_19711);
nor UO_616 (O_616,N_19798,N_18611);
and UO_617 (O_617,N_18908,N_19174);
nor UO_618 (O_618,N_19463,N_19874);
xor UO_619 (O_619,N_19181,N_18649);
and UO_620 (O_620,N_19402,N_19652);
or UO_621 (O_621,N_18659,N_18956);
xor UO_622 (O_622,N_19354,N_19823);
nor UO_623 (O_623,N_18150,N_19898);
or UO_624 (O_624,N_18831,N_19753);
and UO_625 (O_625,N_18960,N_18538);
nor UO_626 (O_626,N_18824,N_18242);
nor UO_627 (O_627,N_18690,N_19639);
or UO_628 (O_628,N_19891,N_18022);
or UO_629 (O_629,N_18589,N_19745);
and UO_630 (O_630,N_18710,N_18802);
nand UO_631 (O_631,N_19123,N_18969);
or UO_632 (O_632,N_18853,N_18641);
or UO_633 (O_633,N_19869,N_18236);
nor UO_634 (O_634,N_19603,N_18907);
and UO_635 (O_635,N_19800,N_18604);
nand UO_636 (O_636,N_18225,N_18238);
and UO_637 (O_637,N_18128,N_19605);
xnor UO_638 (O_638,N_18119,N_19771);
nand UO_639 (O_639,N_18002,N_18633);
or UO_640 (O_640,N_19008,N_18518);
and UO_641 (O_641,N_18129,N_19770);
nand UO_642 (O_642,N_19030,N_18996);
and UO_643 (O_643,N_19044,N_18480);
nor UO_644 (O_644,N_18330,N_19598);
nand UO_645 (O_645,N_19069,N_19735);
xnor UO_646 (O_646,N_18609,N_19371);
nand UO_647 (O_647,N_19802,N_19418);
xor UO_648 (O_648,N_19094,N_19933);
and UO_649 (O_649,N_19594,N_19343);
or UO_650 (O_650,N_19862,N_19218);
nand UO_651 (O_651,N_18998,N_18094);
nand UO_652 (O_652,N_19358,N_19236);
or UO_653 (O_653,N_18402,N_18479);
and UO_654 (O_654,N_18333,N_18293);
nand UO_655 (O_655,N_19107,N_18334);
nand UO_656 (O_656,N_18086,N_19440);
or UO_657 (O_657,N_18840,N_18791);
and UO_658 (O_658,N_19159,N_18732);
nor UO_659 (O_659,N_18062,N_18651);
and UO_660 (O_660,N_18627,N_19074);
xnor UO_661 (O_661,N_19778,N_19496);
and UO_662 (O_662,N_19777,N_19227);
and UO_663 (O_663,N_19267,N_18155);
nand UO_664 (O_664,N_18310,N_19956);
and UO_665 (O_665,N_19738,N_18171);
nor UO_666 (O_666,N_18959,N_19759);
nor UO_667 (O_667,N_18616,N_19591);
or UO_668 (O_668,N_18629,N_18198);
nor UO_669 (O_669,N_19845,N_19670);
and UO_670 (O_670,N_18342,N_19981);
or UO_671 (O_671,N_18231,N_19146);
or UO_672 (O_672,N_19541,N_18432);
xor UO_673 (O_673,N_19868,N_19060);
nor UO_674 (O_674,N_18769,N_18929);
or UO_675 (O_675,N_19322,N_18976);
or UO_676 (O_676,N_19931,N_18798);
nand UO_677 (O_677,N_19342,N_18152);
or UO_678 (O_678,N_19485,N_18752);
or UO_679 (O_679,N_18303,N_19872);
or UO_680 (O_680,N_19889,N_18212);
or UO_681 (O_681,N_18042,N_19538);
nand UO_682 (O_682,N_19606,N_19551);
or UO_683 (O_683,N_18278,N_19421);
or UO_684 (O_684,N_18222,N_18747);
and UO_685 (O_685,N_19969,N_19378);
or UO_686 (O_686,N_19266,N_18843);
or UO_687 (O_687,N_18135,N_18821);
xor UO_688 (O_688,N_18924,N_19863);
and UO_689 (O_689,N_19666,N_19100);
or UO_690 (O_690,N_19797,N_19264);
nand UO_691 (O_691,N_18369,N_19423);
or UO_692 (O_692,N_18264,N_19780);
or UO_693 (O_693,N_19918,N_18398);
nand UO_694 (O_694,N_19101,N_19979);
or UO_695 (O_695,N_19905,N_18862);
nor UO_696 (O_696,N_18408,N_18542);
nand UO_697 (O_697,N_19973,N_19577);
or UO_698 (O_698,N_19118,N_18919);
nor UO_699 (O_699,N_19370,N_19017);
nor UO_700 (O_700,N_19105,N_18613);
nor UO_701 (O_701,N_18031,N_18946);
nor UO_702 (O_702,N_19912,N_19155);
nor UO_703 (O_703,N_19169,N_19170);
nand UO_704 (O_704,N_18224,N_19565);
nor UO_705 (O_705,N_18266,N_18566);
xor UO_706 (O_706,N_18081,N_18411);
xor UO_707 (O_707,N_18471,N_18051);
or UO_708 (O_708,N_18348,N_19310);
or UO_709 (O_709,N_19840,N_19665);
nor UO_710 (O_710,N_18779,N_19633);
or UO_711 (O_711,N_18292,N_19295);
or UO_712 (O_712,N_18925,N_18716);
nand UO_713 (O_713,N_19958,N_18082);
and UO_714 (O_714,N_18070,N_18561);
or UO_715 (O_715,N_19368,N_19966);
and UO_716 (O_716,N_18106,N_19728);
nor UO_717 (O_717,N_19225,N_19083);
or UO_718 (O_718,N_18764,N_19841);
and UO_719 (O_719,N_19319,N_18221);
nor UO_720 (O_720,N_19164,N_18065);
and UO_721 (O_721,N_18006,N_19271);
or UO_722 (O_722,N_19483,N_18640);
nor UO_723 (O_723,N_18216,N_18738);
nor UO_724 (O_724,N_18478,N_18162);
or UO_725 (O_725,N_18192,N_18705);
and UO_726 (O_726,N_19766,N_18244);
or UO_727 (O_727,N_18893,N_19014);
and UO_728 (O_728,N_19601,N_18958);
nor UO_729 (O_729,N_18885,N_19836);
xor UO_730 (O_730,N_18562,N_19881);
or UO_731 (O_731,N_19630,N_18774);
nand UO_732 (O_732,N_19575,N_18896);
and UO_733 (O_733,N_18728,N_18004);
xor UO_734 (O_734,N_18590,N_19873);
xor UO_735 (O_735,N_19687,N_19530);
nor UO_736 (O_736,N_19162,N_19949);
nand UO_737 (O_737,N_18417,N_18386);
nand UO_738 (O_738,N_19239,N_18693);
xor UO_739 (O_739,N_19569,N_19261);
nor UO_740 (O_740,N_18265,N_19621);
or UO_741 (O_741,N_18533,N_19431);
and UO_742 (O_742,N_19277,N_18347);
and UO_743 (O_743,N_18951,N_19013);
nor UO_744 (O_744,N_19507,N_18634);
nand UO_745 (O_745,N_19274,N_19573);
or UO_746 (O_746,N_18933,N_18112);
and UO_747 (O_747,N_19999,N_19796);
nand UO_748 (O_748,N_18811,N_18233);
nand UO_749 (O_749,N_18647,N_18381);
nor UO_750 (O_750,N_19198,N_18804);
and UO_751 (O_751,N_18299,N_19781);
and UO_752 (O_752,N_18694,N_19917);
or UO_753 (O_753,N_19498,N_18767);
or UO_754 (O_754,N_19589,N_18055);
nand UO_755 (O_755,N_19126,N_19051);
and UO_756 (O_756,N_19629,N_18496);
and UO_757 (O_757,N_19285,N_18254);
nand UO_758 (O_758,N_19818,N_19048);
nand UO_759 (O_759,N_19384,N_18483);
or UO_760 (O_760,N_18677,N_19006);
or UO_761 (O_761,N_19007,N_18438);
nand UO_762 (O_762,N_19719,N_19379);
and UO_763 (O_763,N_18939,N_19156);
xnor UO_764 (O_764,N_19301,N_18631);
or UO_765 (O_765,N_19757,N_18365);
or UO_766 (O_766,N_19409,N_18830);
nand UO_767 (O_767,N_18068,N_19690);
or UO_768 (O_768,N_19724,N_18826);
nor UO_769 (O_769,N_19658,N_19746);
and UO_770 (O_770,N_18354,N_18484);
and UO_771 (O_771,N_19257,N_18435);
or UO_772 (O_772,N_18967,N_18130);
and UO_773 (O_773,N_18897,N_19552);
nor UO_774 (O_774,N_18317,N_18661);
and UO_775 (O_775,N_18874,N_18148);
and UO_776 (O_776,N_19420,N_19534);
or UO_777 (O_777,N_18989,N_19259);
or UO_778 (O_778,N_18975,N_19115);
nor UO_779 (O_779,N_18765,N_18692);
and UO_780 (O_780,N_18521,N_19147);
or UO_781 (O_781,N_18930,N_19570);
and UO_782 (O_782,N_19835,N_18535);
or UO_783 (O_783,N_19167,N_18267);
and UO_784 (O_784,N_18017,N_18403);
nor UO_785 (O_785,N_18388,N_18426);
or UO_786 (O_786,N_18970,N_19542);
or UO_787 (O_787,N_18256,N_19944);
and UO_788 (O_788,N_18594,N_18529);
and UO_789 (O_789,N_19505,N_19210);
or UO_790 (O_790,N_18795,N_19935);
nand UO_791 (O_791,N_19650,N_19678);
nor UO_792 (O_792,N_18744,N_19866);
nor UO_793 (O_793,N_18277,N_19749);
xor UO_794 (O_794,N_19313,N_19545);
and UO_795 (O_795,N_19961,N_18319);
or UO_796 (O_796,N_18880,N_18180);
nand UO_797 (O_797,N_18670,N_19097);
nor UO_798 (O_798,N_19500,N_18301);
and UO_799 (O_799,N_19832,N_18952);
nor UO_800 (O_800,N_19901,N_18850);
or UO_801 (O_801,N_19001,N_18335);
and UO_802 (O_802,N_19600,N_19829);
nor UO_803 (O_803,N_19334,N_18443);
xnor UO_804 (O_804,N_19211,N_18819);
xor UO_805 (O_805,N_18618,N_19394);
nor UO_806 (O_806,N_19544,N_19540);
nand UO_807 (O_807,N_18624,N_18258);
or UO_808 (O_808,N_19434,N_18889);
or UO_809 (O_809,N_18891,N_18822);
nand UO_810 (O_810,N_18576,N_18572);
and UO_811 (O_811,N_18790,N_18556);
nand UO_812 (O_812,N_19352,N_19476);
xor UO_813 (O_813,N_18169,N_19501);
nor UO_814 (O_814,N_18977,N_18541);
nand UO_815 (O_815,N_18498,N_19715);
nand UO_816 (O_816,N_19119,N_18524);
xor UO_817 (O_817,N_19299,N_19160);
nand UO_818 (O_818,N_18806,N_18788);
nor UO_819 (O_819,N_18565,N_18096);
and UO_820 (O_820,N_19824,N_19280);
and UO_821 (O_821,N_18903,N_19990);
nand UO_822 (O_822,N_18623,N_18875);
and UO_823 (O_823,N_18425,N_19068);
xnor UO_824 (O_824,N_18011,N_18459);
or UO_825 (O_825,N_18401,N_19596);
nand UO_826 (O_826,N_19396,N_18102);
nand UO_827 (O_827,N_18203,N_18873);
or UO_828 (O_828,N_18043,N_18409);
or UO_829 (O_829,N_19238,N_19585);
or UO_830 (O_830,N_19547,N_19512);
or UO_831 (O_831,N_18487,N_18586);
or UO_832 (O_832,N_18184,N_19694);
or UO_833 (O_833,N_19611,N_18185);
nand UO_834 (O_834,N_18582,N_19588);
xnor UO_835 (O_835,N_18817,N_18620);
or UO_836 (O_836,N_19177,N_19668);
and UO_837 (O_837,N_18202,N_19435);
or UO_838 (O_838,N_18610,N_18578);
and UO_839 (O_839,N_18218,N_19697);
or UO_840 (O_840,N_18878,N_19194);
or UO_841 (O_841,N_19922,N_19768);
nor UO_842 (O_842,N_19925,N_19109);
or UO_843 (O_843,N_18418,N_18776);
or UO_844 (O_844,N_19135,N_18503);
xor UO_845 (O_845,N_19754,N_19786);
xor UO_846 (O_846,N_19986,N_19964);
nand UO_847 (O_847,N_18780,N_19472);
or UO_848 (O_848,N_18474,N_19689);
or UO_849 (O_849,N_18711,N_19339);
nor UO_850 (O_850,N_19899,N_18546);
or UO_851 (O_851,N_19793,N_18328);
nor UO_852 (O_852,N_19240,N_19415);
and UO_853 (O_853,N_19608,N_18464);
or UO_854 (O_854,N_19446,N_19988);
nor UO_855 (O_855,N_18355,N_19049);
nor UO_856 (O_856,N_19224,N_19436);
xnor UO_857 (O_857,N_19870,N_19344);
or UO_858 (O_858,N_18356,N_19970);
xnor UO_859 (O_859,N_18727,N_19149);
nand UO_860 (O_860,N_18994,N_19399);
or UO_861 (O_861,N_18245,N_19636);
or UO_862 (O_862,N_19807,N_19736);
nor UO_863 (O_863,N_19801,N_19417);
nand UO_864 (O_864,N_19572,N_19760);
nand UO_865 (O_865,N_19201,N_19662);
xnor UO_866 (O_866,N_18223,N_19597);
and UO_867 (O_867,N_19338,N_18591);
nor UO_868 (O_868,N_18950,N_18287);
xnor UO_869 (O_869,N_18439,N_18367);
or UO_870 (O_870,N_18138,N_19527);
nor UO_871 (O_871,N_19040,N_18596);
and UO_872 (O_872,N_19506,N_18581);
nand UO_873 (O_873,N_18280,N_18614);
nand UO_874 (O_874,N_18430,N_18777);
nand UO_875 (O_875,N_19726,N_18545);
nand UO_876 (O_876,N_18298,N_18592);
nand UO_877 (O_877,N_18332,N_18215);
nor UO_878 (O_878,N_19179,N_18437);
nand UO_879 (O_879,N_18063,N_18876);
nand UO_880 (O_880,N_19787,N_19521);
and UO_881 (O_881,N_18450,N_19080);
nand UO_882 (O_882,N_19279,N_18786);
or UO_883 (O_883,N_19132,N_18021);
and UO_884 (O_884,N_18983,N_18159);
xor UO_885 (O_885,N_19144,N_19761);
nor UO_886 (O_886,N_18841,N_18799);
nand UO_887 (O_887,N_18639,N_19145);
nor UO_888 (O_888,N_19972,N_18134);
xnor UO_889 (O_889,N_18528,N_19989);
xor UO_890 (O_890,N_18886,N_18284);
and UO_891 (O_891,N_18167,N_19539);
and UO_892 (O_892,N_18232,N_19987);
nor UO_893 (O_893,N_19208,N_18308);
and UO_894 (O_894,N_19864,N_19879);
nor UO_895 (O_895,N_19947,N_18122);
and UO_896 (O_896,N_18124,N_19345);
xnor UO_897 (O_897,N_18523,N_19756);
or UO_898 (O_898,N_19963,N_18660);
or UO_899 (O_899,N_19525,N_18196);
nor UO_900 (O_900,N_19127,N_18760);
and UO_901 (O_901,N_19671,N_19317);
and UO_902 (O_902,N_18085,N_19361);
and UO_903 (O_903,N_19810,N_19268);
or UO_904 (O_904,N_19533,N_18206);
nor UO_905 (O_905,N_18722,N_19784);
and UO_906 (O_906,N_19374,N_19878);
nand UO_907 (O_907,N_19443,N_19942);
or UO_908 (O_908,N_19385,N_19058);
or UO_909 (O_909,N_19397,N_18291);
and UO_910 (O_910,N_19681,N_19113);
or UO_911 (O_911,N_18241,N_18010);
or UO_912 (O_912,N_19398,N_18410);
and UO_913 (O_913,N_18133,N_18932);
nand UO_914 (O_914,N_18548,N_18516);
xnor UO_915 (O_915,N_19750,N_18868);
or UO_916 (O_916,N_18943,N_18539);
nand UO_917 (O_917,N_19186,N_19021);
nand UO_918 (O_918,N_19743,N_19168);
xor UO_919 (O_919,N_19834,N_19812);
nand UO_920 (O_920,N_19355,N_19036);
xor UO_921 (O_921,N_19470,N_18789);
or UO_922 (O_922,N_18290,N_18758);
nor UO_923 (O_923,N_18197,N_19369);
xor UO_924 (O_924,N_18968,N_18440);
and UO_925 (O_925,N_18855,N_19035);
and UO_926 (O_926,N_18089,N_19027);
nor UO_927 (O_927,N_18174,N_18061);
nand UO_928 (O_928,N_19888,N_19430);
xnor UO_929 (O_929,N_19320,N_19072);
nor UO_930 (O_930,N_18413,N_18735);
and UO_931 (O_931,N_19163,N_19270);
and UO_932 (O_932,N_18688,N_18743);
nor UO_933 (O_933,N_19637,N_19491);
or UO_934 (O_934,N_19932,N_18940);
nand UO_935 (O_935,N_18288,N_18325);
nand UO_936 (O_936,N_18044,N_18248);
nand UO_937 (O_937,N_19057,N_18144);
or UO_938 (O_938,N_19248,N_18628);
and UO_939 (O_939,N_18127,N_18731);
nand UO_940 (O_940,N_18023,N_18014);
nand UO_941 (O_941,N_18704,N_18344);
and UO_942 (O_942,N_18587,N_18008);
nand UO_943 (O_943,N_19230,N_19084);
nor UO_944 (O_944,N_19939,N_19189);
or UO_945 (O_945,N_19308,N_18199);
nand UO_946 (O_946,N_19994,N_19216);
nor UO_947 (O_947,N_18495,N_18739);
nand UO_948 (O_948,N_18574,N_19640);
nand UO_949 (O_949,N_18987,N_18870);
and UO_950 (O_950,N_19395,N_18917);
xnor UO_951 (O_951,N_19737,N_18262);
xnor UO_952 (O_952,N_18858,N_19357);
or UO_953 (O_953,N_19012,N_18389);
and UO_954 (O_954,N_18877,N_19054);
xnor UO_955 (O_955,N_18713,N_18454);
nand UO_956 (O_956,N_18836,N_18860);
and UO_957 (O_957,N_18302,N_19028);
or UO_958 (O_958,N_18813,N_18935);
nor UO_959 (O_959,N_19977,N_18700);
nor UO_960 (O_960,N_18228,N_19676);
nand UO_961 (O_961,N_19980,N_19043);
xor UO_962 (O_962,N_18615,N_19003);
nor UO_963 (O_963,N_19782,N_19412);
nand UO_964 (O_964,N_19220,N_18534);
or UO_965 (O_965,N_19789,N_19056);
xnor UO_966 (O_966,N_19090,N_19411);
nand UO_967 (O_967,N_18884,N_18637);
nand UO_968 (O_968,N_19315,N_18662);
nand UO_969 (O_969,N_18761,N_19333);
and UO_970 (O_970,N_19050,N_19173);
or UO_971 (O_971,N_19138,N_18473);
or UO_972 (O_972,N_19255,N_18753);
or UO_973 (O_973,N_19404,N_19755);
xor UO_974 (O_974,N_18406,N_18734);
nand UO_975 (O_975,N_19532,N_19685);
or UO_976 (O_976,N_19536,N_19730);
or UO_977 (O_977,N_18838,N_19632);
xor UO_978 (O_978,N_19562,N_18307);
nor UO_979 (O_979,N_19699,N_19432);
nand UO_980 (O_980,N_19326,N_19556);
nor UO_981 (O_981,N_18422,N_19960);
nand UO_982 (O_982,N_18866,N_19974);
nand UO_983 (O_983,N_18599,N_18246);
nor UO_984 (O_984,N_19860,N_18316);
and UO_985 (O_985,N_18517,N_18625);
nand UO_986 (O_986,N_19952,N_18193);
nand UO_987 (O_987,N_19349,N_19579);
nor UO_988 (O_988,N_19767,N_18654);
nand UO_989 (O_989,N_19702,N_19985);
and UO_990 (O_990,N_18673,N_19722);
xor UO_991 (O_991,N_19557,N_18036);
and UO_992 (O_992,N_18569,N_19158);
xor UO_993 (O_993,N_19445,N_19053);
and UO_994 (O_994,N_18074,N_18151);
and UO_995 (O_995,N_18270,N_18028);
or UO_996 (O_996,N_19513,N_18559);
or UO_997 (O_997,N_18745,N_19373);
xor UO_998 (O_998,N_18282,N_18580);
or UO_999 (O_999,N_18311,N_18453);
and UO_1000 (O_1000,N_19128,N_18998);
nand UO_1001 (O_1001,N_18904,N_18031);
and UO_1002 (O_1002,N_19263,N_19471);
nor UO_1003 (O_1003,N_18135,N_19439);
nor UO_1004 (O_1004,N_19638,N_18343);
nor UO_1005 (O_1005,N_19521,N_18500);
or UO_1006 (O_1006,N_18267,N_19747);
or UO_1007 (O_1007,N_19938,N_18728);
or UO_1008 (O_1008,N_19459,N_19359);
and UO_1009 (O_1009,N_18120,N_18849);
and UO_1010 (O_1010,N_19951,N_18020);
nand UO_1011 (O_1011,N_19828,N_18855);
and UO_1012 (O_1012,N_18654,N_18977);
or UO_1013 (O_1013,N_18993,N_19777);
nand UO_1014 (O_1014,N_19178,N_19109);
xnor UO_1015 (O_1015,N_19778,N_19292);
nand UO_1016 (O_1016,N_19541,N_19978);
nor UO_1017 (O_1017,N_18815,N_18282);
or UO_1018 (O_1018,N_19227,N_18263);
xor UO_1019 (O_1019,N_19318,N_18833);
and UO_1020 (O_1020,N_18042,N_19041);
nor UO_1021 (O_1021,N_19079,N_18089);
nor UO_1022 (O_1022,N_18902,N_19862);
and UO_1023 (O_1023,N_18822,N_18296);
and UO_1024 (O_1024,N_18894,N_19688);
nand UO_1025 (O_1025,N_19085,N_19268);
xor UO_1026 (O_1026,N_18191,N_18250);
nor UO_1027 (O_1027,N_18952,N_18186);
nor UO_1028 (O_1028,N_19078,N_19923);
nor UO_1029 (O_1029,N_19741,N_19816);
xnor UO_1030 (O_1030,N_19321,N_19570);
and UO_1031 (O_1031,N_19407,N_19410);
or UO_1032 (O_1032,N_18398,N_19646);
nand UO_1033 (O_1033,N_18575,N_19672);
nor UO_1034 (O_1034,N_18327,N_18387);
or UO_1035 (O_1035,N_19214,N_19736);
or UO_1036 (O_1036,N_19962,N_18081);
xnor UO_1037 (O_1037,N_19588,N_18904);
nand UO_1038 (O_1038,N_18413,N_19737);
or UO_1039 (O_1039,N_19695,N_18518);
nand UO_1040 (O_1040,N_18289,N_18964);
and UO_1041 (O_1041,N_19564,N_18044);
and UO_1042 (O_1042,N_18753,N_18937);
or UO_1043 (O_1043,N_19004,N_19935);
nor UO_1044 (O_1044,N_19380,N_19779);
nor UO_1045 (O_1045,N_19132,N_18361);
nor UO_1046 (O_1046,N_19240,N_19170);
and UO_1047 (O_1047,N_19496,N_19580);
xor UO_1048 (O_1048,N_19419,N_19269);
and UO_1049 (O_1049,N_19140,N_18270);
xor UO_1050 (O_1050,N_19061,N_19307);
nand UO_1051 (O_1051,N_19605,N_19891);
or UO_1052 (O_1052,N_19448,N_18944);
nand UO_1053 (O_1053,N_18426,N_18687);
xnor UO_1054 (O_1054,N_19139,N_18176);
or UO_1055 (O_1055,N_19939,N_19605);
or UO_1056 (O_1056,N_18426,N_18145);
nor UO_1057 (O_1057,N_19781,N_19481);
and UO_1058 (O_1058,N_19364,N_18475);
nor UO_1059 (O_1059,N_19969,N_18866);
nand UO_1060 (O_1060,N_18567,N_18360);
or UO_1061 (O_1061,N_18359,N_18622);
or UO_1062 (O_1062,N_18295,N_19439);
nor UO_1063 (O_1063,N_18852,N_18602);
nand UO_1064 (O_1064,N_19490,N_19580);
or UO_1065 (O_1065,N_18578,N_19606);
nand UO_1066 (O_1066,N_19023,N_19487);
xnor UO_1067 (O_1067,N_18744,N_19948);
xor UO_1068 (O_1068,N_19853,N_18890);
xnor UO_1069 (O_1069,N_18846,N_19373);
nand UO_1070 (O_1070,N_18652,N_19256);
and UO_1071 (O_1071,N_18099,N_18969);
nand UO_1072 (O_1072,N_19147,N_19169);
or UO_1073 (O_1073,N_19051,N_19390);
nor UO_1074 (O_1074,N_19958,N_18060);
and UO_1075 (O_1075,N_18230,N_18893);
nor UO_1076 (O_1076,N_19096,N_18783);
and UO_1077 (O_1077,N_19077,N_19956);
and UO_1078 (O_1078,N_18488,N_19845);
nand UO_1079 (O_1079,N_18748,N_18261);
or UO_1080 (O_1080,N_18392,N_18320);
nor UO_1081 (O_1081,N_18591,N_19594);
or UO_1082 (O_1082,N_18058,N_19336);
nor UO_1083 (O_1083,N_19240,N_18785);
or UO_1084 (O_1084,N_19502,N_19553);
or UO_1085 (O_1085,N_18294,N_19473);
or UO_1086 (O_1086,N_19311,N_19317);
or UO_1087 (O_1087,N_19711,N_18562);
nor UO_1088 (O_1088,N_18966,N_19328);
nor UO_1089 (O_1089,N_18151,N_18529);
nand UO_1090 (O_1090,N_18541,N_19418);
nor UO_1091 (O_1091,N_19848,N_19866);
or UO_1092 (O_1092,N_19615,N_19887);
nand UO_1093 (O_1093,N_18776,N_19483);
or UO_1094 (O_1094,N_18586,N_18359);
or UO_1095 (O_1095,N_19344,N_19637);
or UO_1096 (O_1096,N_18117,N_19073);
and UO_1097 (O_1097,N_19415,N_19197);
and UO_1098 (O_1098,N_19718,N_18465);
or UO_1099 (O_1099,N_19284,N_19082);
and UO_1100 (O_1100,N_19858,N_18266);
nand UO_1101 (O_1101,N_19528,N_19531);
nand UO_1102 (O_1102,N_19760,N_18654);
nand UO_1103 (O_1103,N_19943,N_18357);
or UO_1104 (O_1104,N_18887,N_18762);
nor UO_1105 (O_1105,N_19178,N_19017);
xor UO_1106 (O_1106,N_18629,N_18768);
nor UO_1107 (O_1107,N_18614,N_18980);
or UO_1108 (O_1108,N_19456,N_18700);
nand UO_1109 (O_1109,N_18661,N_18173);
or UO_1110 (O_1110,N_18037,N_18401);
nand UO_1111 (O_1111,N_19626,N_19455);
nand UO_1112 (O_1112,N_19949,N_18754);
and UO_1113 (O_1113,N_18355,N_19446);
and UO_1114 (O_1114,N_18013,N_19963);
nor UO_1115 (O_1115,N_19417,N_18930);
or UO_1116 (O_1116,N_19894,N_19969);
and UO_1117 (O_1117,N_19232,N_18295);
nand UO_1118 (O_1118,N_19795,N_18504);
nand UO_1119 (O_1119,N_19430,N_19482);
nor UO_1120 (O_1120,N_19750,N_18215);
and UO_1121 (O_1121,N_19932,N_18305);
nand UO_1122 (O_1122,N_18689,N_19431);
nor UO_1123 (O_1123,N_18555,N_18536);
nand UO_1124 (O_1124,N_18858,N_18850);
nor UO_1125 (O_1125,N_19719,N_19238);
nor UO_1126 (O_1126,N_18105,N_19996);
xnor UO_1127 (O_1127,N_19949,N_18215);
or UO_1128 (O_1128,N_19496,N_18975);
and UO_1129 (O_1129,N_19357,N_19551);
or UO_1130 (O_1130,N_19835,N_18358);
nand UO_1131 (O_1131,N_18519,N_18364);
nand UO_1132 (O_1132,N_18580,N_18850);
and UO_1133 (O_1133,N_18998,N_19013);
nand UO_1134 (O_1134,N_19905,N_19913);
nand UO_1135 (O_1135,N_18144,N_18209);
nor UO_1136 (O_1136,N_19173,N_18315);
nand UO_1137 (O_1137,N_18407,N_18665);
or UO_1138 (O_1138,N_18865,N_19262);
and UO_1139 (O_1139,N_18159,N_19595);
xor UO_1140 (O_1140,N_18596,N_18751);
nand UO_1141 (O_1141,N_19537,N_19738);
and UO_1142 (O_1142,N_18326,N_18896);
nor UO_1143 (O_1143,N_19665,N_18675);
and UO_1144 (O_1144,N_18765,N_19834);
nor UO_1145 (O_1145,N_19475,N_19256);
or UO_1146 (O_1146,N_19730,N_18443);
nor UO_1147 (O_1147,N_18656,N_18935);
or UO_1148 (O_1148,N_19268,N_18409);
and UO_1149 (O_1149,N_18189,N_18791);
and UO_1150 (O_1150,N_19068,N_18694);
nor UO_1151 (O_1151,N_19090,N_19364);
nor UO_1152 (O_1152,N_18027,N_18908);
xnor UO_1153 (O_1153,N_18924,N_18267);
nand UO_1154 (O_1154,N_18896,N_19265);
and UO_1155 (O_1155,N_19087,N_19307);
or UO_1156 (O_1156,N_18116,N_19594);
nor UO_1157 (O_1157,N_19023,N_19826);
nand UO_1158 (O_1158,N_19523,N_18860);
and UO_1159 (O_1159,N_19417,N_18166);
nor UO_1160 (O_1160,N_18275,N_19015);
nand UO_1161 (O_1161,N_18944,N_19824);
nor UO_1162 (O_1162,N_19113,N_19929);
or UO_1163 (O_1163,N_19882,N_18697);
and UO_1164 (O_1164,N_18265,N_18685);
and UO_1165 (O_1165,N_19056,N_18729);
nor UO_1166 (O_1166,N_18474,N_18639);
or UO_1167 (O_1167,N_19488,N_19033);
xor UO_1168 (O_1168,N_18528,N_19985);
nor UO_1169 (O_1169,N_18406,N_19802);
and UO_1170 (O_1170,N_18457,N_19075);
nand UO_1171 (O_1171,N_18021,N_19325);
nor UO_1172 (O_1172,N_19360,N_18991);
nor UO_1173 (O_1173,N_19923,N_19470);
nand UO_1174 (O_1174,N_18626,N_19175);
nor UO_1175 (O_1175,N_19885,N_19605);
nor UO_1176 (O_1176,N_19979,N_18610);
nand UO_1177 (O_1177,N_19098,N_19966);
or UO_1178 (O_1178,N_18101,N_19849);
or UO_1179 (O_1179,N_18553,N_18405);
nand UO_1180 (O_1180,N_19890,N_18912);
nor UO_1181 (O_1181,N_19804,N_18111);
nor UO_1182 (O_1182,N_19507,N_18798);
nand UO_1183 (O_1183,N_19668,N_19436);
nand UO_1184 (O_1184,N_19976,N_19372);
or UO_1185 (O_1185,N_19562,N_19950);
nand UO_1186 (O_1186,N_19915,N_19970);
nor UO_1187 (O_1187,N_18016,N_18292);
nand UO_1188 (O_1188,N_19299,N_19956);
xor UO_1189 (O_1189,N_18470,N_19524);
or UO_1190 (O_1190,N_18500,N_18712);
and UO_1191 (O_1191,N_19827,N_19065);
nor UO_1192 (O_1192,N_19579,N_18217);
or UO_1193 (O_1193,N_19806,N_19310);
nand UO_1194 (O_1194,N_19142,N_19528);
nand UO_1195 (O_1195,N_18159,N_18331);
xnor UO_1196 (O_1196,N_18311,N_18463);
nor UO_1197 (O_1197,N_18524,N_19794);
nor UO_1198 (O_1198,N_19440,N_19657);
nor UO_1199 (O_1199,N_19964,N_18893);
nor UO_1200 (O_1200,N_19324,N_18127);
nand UO_1201 (O_1201,N_19120,N_19003);
and UO_1202 (O_1202,N_18065,N_19477);
xnor UO_1203 (O_1203,N_19199,N_18417);
nor UO_1204 (O_1204,N_18914,N_18217);
nand UO_1205 (O_1205,N_19074,N_18426);
nor UO_1206 (O_1206,N_19186,N_19430);
and UO_1207 (O_1207,N_18209,N_18262);
nand UO_1208 (O_1208,N_18984,N_19697);
nor UO_1209 (O_1209,N_19916,N_19792);
nor UO_1210 (O_1210,N_18096,N_18815);
and UO_1211 (O_1211,N_18193,N_19878);
and UO_1212 (O_1212,N_18373,N_18721);
nand UO_1213 (O_1213,N_18576,N_18114);
xnor UO_1214 (O_1214,N_18566,N_19486);
nand UO_1215 (O_1215,N_18666,N_18742);
nor UO_1216 (O_1216,N_19151,N_19250);
and UO_1217 (O_1217,N_18054,N_18308);
or UO_1218 (O_1218,N_18634,N_19696);
and UO_1219 (O_1219,N_19058,N_18404);
or UO_1220 (O_1220,N_18117,N_19205);
nand UO_1221 (O_1221,N_18277,N_18321);
or UO_1222 (O_1222,N_19423,N_18550);
and UO_1223 (O_1223,N_19723,N_19255);
nor UO_1224 (O_1224,N_18302,N_19539);
or UO_1225 (O_1225,N_19048,N_19137);
or UO_1226 (O_1226,N_19967,N_19072);
and UO_1227 (O_1227,N_18261,N_19361);
and UO_1228 (O_1228,N_18462,N_18142);
xor UO_1229 (O_1229,N_19825,N_19328);
nand UO_1230 (O_1230,N_19258,N_18914);
nor UO_1231 (O_1231,N_18003,N_19124);
or UO_1232 (O_1232,N_18731,N_18732);
or UO_1233 (O_1233,N_18597,N_18193);
or UO_1234 (O_1234,N_19078,N_19920);
and UO_1235 (O_1235,N_18422,N_19240);
nor UO_1236 (O_1236,N_18132,N_18937);
nor UO_1237 (O_1237,N_19082,N_19243);
and UO_1238 (O_1238,N_18635,N_19040);
nand UO_1239 (O_1239,N_18498,N_18080);
and UO_1240 (O_1240,N_18710,N_18095);
or UO_1241 (O_1241,N_18645,N_18021);
nand UO_1242 (O_1242,N_18303,N_19839);
nor UO_1243 (O_1243,N_18559,N_18877);
xor UO_1244 (O_1244,N_19542,N_19016);
xor UO_1245 (O_1245,N_18213,N_19797);
nor UO_1246 (O_1246,N_18972,N_18169);
or UO_1247 (O_1247,N_19706,N_19548);
nand UO_1248 (O_1248,N_18049,N_18396);
nor UO_1249 (O_1249,N_19386,N_19891);
nor UO_1250 (O_1250,N_19431,N_18188);
nor UO_1251 (O_1251,N_19801,N_18095);
and UO_1252 (O_1252,N_18776,N_19288);
or UO_1253 (O_1253,N_18708,N_18503);
and UO_1254 (O_1254,N_19705,N_19202);
and UO_1255 (O_1255,N_18644,N_18716);
xnor UO_1256 (O_1256,N_19147,N_19607);
nor UO_1257 (O_1257,N_18326,N_19587);
and UO_1258 (O_1258,N_18207,N_19019);
or UO_1259 (O_1259,N_19306,N_19193);
or UO_1260 (O_1260,N_18850,N_19624);
nand UO_1261 (O_1261,N_19987,N_18858);
nand UO_1262 (O_1262,N_19061,N_19276);
nor UO_1263 (O_1263,N_18392,N_18598);
nor UO_1264 (O_1264,N_18357,N_19753);
nand UO_1265 (O_1265,N_19631,N_19988);
and UO_1266 (O_1266,N_18022,N_18538);
xor UO_1267 (O_1267,N_18689,N_19555);
nand UO_1268 (O_1268,N_18317,N_18580);
or UO_1269 (O_1269,N_19950,N_18038);
nand UO_1270 (O_1270,N_19448,N_18865);
or UO_1271 (O_1271,N_18250,N_19088);
nand UO_1272 (O_1272,N_18724,N_19768);
and UO_1273 (O_1273,N_19264,N_18684);
and UO_1274 (O_1274,N_19212,N_18295);
and UO_1275 (O_1275,N_19216,N_18230);
and UO_1276 (O_1276,N_18394,N_19344);
nand UO_1277 (O_1277,N_19508,N_19169);
nor UO_1278 (O_1278,N_18270,N_18351);
nor UO_1279 (O_1279,N_18695,N_18328);
and UO_1280 (O_1280,N_19644,N_18715);
nor UO_1281 (O_1281,N_19306,N_19175);
and UO_1282 (O_1282,N_18011,N_19317);
nand UO_1283 (O_1283,N_19773,N_18884);
nand UO_1284 (O_1284,N_19758,N_19736);
and UO_1285 (O_1285,N_18148,N_19758);
xor UO_1286 (O_1286,N_19435,N_18739);
or UO_1287 (O_1287,N_18284,N_18190);
nand UO_1288 (O_1288,N_19036,N_18142);
nor UO_1289 (O_1289,N_19628,N_18500);
nand UO_1290 (O_1290,N_18829,N_18229);
or UO_1291 (O_1291,N_19281,N_19192);
nor UO_1292 (O_1292,N_18053,N_18283);
nor UO_1293 (O_1293,N_19388,N_18682);
nor UO_1294 (O_1294,N_18768,N_18897);
nor UO_1295 (O_1295,N_18429,N_18239);
and UO_1296 (O_1296,N_19854,N_19039);
nor UO_1297 (O_1297,N_19004,N_18121);
and UO_1298 (O_1298,N_18003,N_18811);
and UO_1299 (O_1299,N_19297,N_18760);
and UO_1300 (O_1300,N_18951,N_19490);
nor UO_1301 (O_1301,N_18055,N_18968);
and UO_1302 (O_1302,N_19842,N_18251);
nor UO_1303 (O_1303,N_18337,N_18972);
nand UO_1304 (O_1304,N_19853,N_18285);
and UO_1305 (O_1305,N_19637,N_19295);
or UO_1306 (O_1306,N_18351,N_19307);
and UO_1307 (O_1307,N_18181,N_18798);
and UO_1308 (O_1308,N_19797,N_19615);
nand UO_1309 (O_1309,N_18817,N_19238);
nor UO_1310 (O_1310,N_19483,N_18593);
nand UO_1311 (O_1311,N_18615,N_19187);
and UO_1312 (O_1312,N_18299,N_18060);
and UO_1313 (O_1313,N_18713,N_18574);
and UO_1314 (O_1314,N_18042,N_19200);
or UO_1315 (O_1315,N_18137,N_18105);
and UO_1316 (O_1316,N_19407,N_18592);
or UO_1317 (O_1317,N_18170,N_19495);
or UO_1318 (O_1318,N_19711,N_18031);
or UO_1319 (O_1319,N_19097,N_19986);
nand UO_1320 (O_1320,N_18251,N_18781);
nand UO_1321 (O_1321,N_18669,N_19253);
nand UO_1322 (O_1322,N_19642,N_18548);
nor UO_1323 (O_1323,N_18701,N_18467);
nor UO_1324 (O_1324,N_19031,N_19108);
nor UO_1325 (O_1325,N_18433,N_18597);
nor UO_1326 (O_1326,N_18252,N_18557);
nand UO_1327 (O_1327,N_19056,N_19571);
and UO_1328 (O_1328,N_19307,N_18721);
and UO_1329 (O_1329,N_19486,N_18053);
and UO_1330 (O_1330,N_19300,N_18816);
nand UO_1331 (O_1331,N_19016,N_18706);
or UO_1332 (O_1332,N_18406,N_19550);
nand UO_1333 (O_1333,N_18510,N_18484);
or UO_1334 (O_1334,N_18291,N_18479);
and UO_1335 (O_1335,N_19403,N_18495);
nand UO_1336 (O_1336,N_18628,N_19090);
and UO_1337 (O_1337,N_19056,N_18471);
or UO_1338 (O_1338,N_18885,N_18168);
nor UO_1339 (O_1339,N_19312,N_19586);
nor UO_1340 (O_1340,N_19696,N_19059);
or UO_1341 (O_1341,N_19382,N_18893);
nor UO_1342 (O_1342,N_19056,N_18163);
nor UO_1343 (O_1343,N_18402,N_18999);
and UO_1344 (O_1344,N_19595,N_18191);
or UO_1345 (O_1345,N_18062,N_19994);
xor UO_1346 (O_1346,N_19490,N_19235);
nor UO_1347 (O_1347,N_19386,N_19736);
and UO_1348 (O_1348,N_19930,N_18001);
or UO_1349 (O_1349,N_18059,N_18803);
nor UO_1350 (O_1350,N_18046,N_18707);
nand UO_1351 (O_1351,N_19586,N_19791);
and UO_1352 (O_1352,N_18895,N_19182);
nor UO_1353 (O_1353,N_19060,N_19804);
xnor UO_1354 (O_1354,N_18026,N_19875);
nand UO_1355 (O_1355,N_18685,N_19051);
xor UO_1356 (O_1356,N_19524,N_18677);
and UO_1357 (O_1357,N_19671,N_19844);
nor UO_1358 (O_1358,N_18656,N_18683);
nand UO_1359 (O_1359,N_19581,N_19000);
nor UO_1360 (O_1360,N_19724,N_19295);
or UO_1361 (O_1361,N_19192,N_18137);
and UO_1362 (O_1362,N_18739,N_18045);
nor UO_1363 (O_1363,N_18597,N_18879);
nor UO_1364 (O_1364,N_18370,N_18288);
or UO_1365 (O_1365,N_19970,N_19665);
xor UO_1366 (O_1366,N_18753,N_19663);
nor UO_1367 (O_1367,N_18345,N_18551);
or UO_1368 (O_1368,N_18930,N_19458);
xnor UO_1369 (O_1369,N_19581,N_18999);
nand UO_1370 (O_1370,N_18730,N_19998);
and UO_1371 (O_1371,N_18777,N_18362);
nand UO_1372 (O_1372,N_19760,N_18814);
xor UO_1373 (O_1373,N_18319,N_19754);
or UO_1374 (O_1374,N_18657,N_18939);
nor UO_1375 (O_1375,N_18331,N_19225);
or UO_1376 (O_1376,N_19321,N_19014);
nand UO_1377 (O_1377,N_19249,N_19821);
nand UO_1378 (O_1378,N_18251,N_19837);
xnor UO_1379 (O_1379,N_18931,N_18449);
nor UO_1380 (O_1380,N_19439,N_18913);
nand UO_1381 (O_1381,N_18762,N_19496);
and UO_1382 (O_1382,N_18472,N_19533);
xnor UO_1383 (O_1383,N_18202,N_19155);
and UO_1384 (O_1384,N_18962,N_19570);
and UO_1385 (O_1385,N_19469,N_19785);
or UO_1386 (O_1386,N_18623,N_18899);
and UO_1387 (O_1387,N_19484,N_18625);
or UO_1388 (O_1388,N_18011,N_19420);
xnor UO_1389 (O_1389,N_19760,N_18723);
nand UO_1390 (O_1390,N_18228,N_19942);
nor UO_1391 (O_1391,N_18318,N_18113);
nand UO_1392 (O_1392,N_19931,N_19555);
nor UO_1393 (O_1393,N_18229,N_19145);
nor UO_1394 (O_1394,N_18426,N_18129);
and UO_1395 (O_1395,N_18498,N_18760);
nand UO_1396 (O_1396,N_19809,N_18239);
nand UO_1397 (O_1397,N_18304,N_19291);
or UO_1398 (O_1398,N_18310,N_18483);
and UO_1399 (O_1399,N_19234,N_19091);
nand UO_1400 (O_1400,N_19324,N_18577);
nand UO_1401 (O_1401,N_18248,N_18144);
nor UO_1402 (O_1402,N_19048,N_18285);
nand UO_1403 (O_1403,N_18121,N_19751);
nand UO_1404 (O_1404,N_19845,N_18876);
nand UO_1405 (O_1405,N_18747,N_19111);
nor UO_1406 (O_1406,N_18595,N_19477);
nand UO_1407 (O_1407,N_19870,N_18564);
nor UO_1408 (O_1408,N_18626,N_18700);
and UO_1409 (O_1409,N_18800,N_18005);
nand UO_1410 (O_1410,N_18897,N_18156);
or UO_1411 (O_1411,N_19773,N_19688);
nor UO_1412 (O_1412,N_18791,N_19583);
xnor UO_1413 (O_1413,N_19102,N_19052);
and UO_1414 (O_1414,N_18082,N_18472);
and UO_1415 (O_1415,N_18420,N_18579);
nor UO_1416 (O_1416,N_19302,N_18924);
and UO_1417 (O_1417,N_19227,N_18782);
nor UO_1418 (O_1418,N_18239,N_18921);
nor UO_1419 (O_1419,N_19047,N_19408);
and UO_1420 (O_1420,N_19914,N_19599);
nand UO_1421 (O_1421,N_18040,N_19674);
and UO_1422 (O_1422,N_18845,N_18531);
nand UO_1423 (O_1423,N_18443,N_18948);
nor UO_1424 (O_1424,N_19982,N_19656);
or UO_1425 (O_1425,N_18841,N_19281);
or UO_1426 (O_1426,N_19273,N_19891);
nor UO_1427 (O_1427,N_19373,N_18767);
and UO_1428 (O_1428,N_19768,N_18784);
nand UO_1429 (O_1429,N_18109,N_18358);
nor UO_1430 (O_1430,N_18820,N_19113);
nor UO_1431 (O_1431,N_18023,N_18496);
and UO_1432 (O_1432,N_19829,N_18242);
nand UO_1433 (O_1433,N_18904,N_19027);
and UO_1434 (O_1434,N_19946,N_19527);
nor UO_1435 (O_1435,N_18051,N_19664);
and UO_1436 (O_1436,N_18906,N_18326);
nor UO_1437 (O_1437,N_19056,N_19059);
and UO_1438 (O_1438,N_18534,N_18065);
and UO_1439 (O_1439,N_18646,N_19329);
nand UO_1440 (O_1440,N_19694,N_19324);
nand UO_1441 (O_1441,N_18611,N_19725);
and UO_1442 (O_1442,N_19923,N_18975);
xor UO_1443 (O_1443,N_19535,N_18614);
nand UO_1444 (O_1444,N_18385,N_19245);
nand UO_1445 (O_1445,N_19877,N_19481);
nand UO_1446 (O_1446,N_19147,N_19383);
nand UO_1447 (O_1447,N_18137,N_19625);
or UO_1448 (O_1448,N_19597,N_18512);
or UO_1449 (O_1449,N_18983,N_18527);
and UO_1450 (O_1450,N_19381,N_19440);
xor UO_1451 (O_1451,N_18458,N_19655);
or UO_1452 (O_1452,N_18972,N_18700);
nand UO_1453 (O_1453,N_19085,N_18185);
nand UO_1454 (O_1454,N_18940,N_19519);
nand UO_1455 (O_1455,N_19393,N_18952);
nor UO_1456 (O_1456,N_18892,N_18377);
or UO_1457 (O_1457,N_18180,N_19186);
nand UO_1458 (O_1458,N_18027,N_19830);
or UO_1459 (O_1459,N_18973,N_19491);
nor UO_1460 (O_1460,N_18403,N_18346);
nor UO_1461 (O_1461,N_19339,N_18737);
nor UO_1462 (O_1462,N_18859,N_19073);
and UO_1463 (O_1463,N_18420,N_18068);
and UO_1464 (O_1464,N_18283,N_18551);
nor UO_1465 (O_1465,N_19678,N_18332);
and UO_1466 (O_1466,N_18698,N_18048);
nand UO_1467 (O_1467,N_19704,N_18975);
nand UO_1468 (O_1468,N_18190,N_18409);
or UO_1469 (O_1469,N_18245,N_19117);
nand UO_1470 (O_1470,N_19944,N_18069);
and UO_1471 (O_1471,N_18605,N_18586);
nor UO_1472 (O_1472,N_19377,N_19119);
or UO_1473 (O_1473,N_19140,N_19468);
xnor UO_1474 (O_1474,N_19505,N_18626);
and UO_1475 (O_1475,N_18403,N_18781);
and UO_1476 (O_1476,N_19257,N_18375);
nand UO_1477 (O_1477,N_18489,N_19023);
or UO_1478 (O_1478,N_19860,N_19655);
nand UO_1479 (O_1479,N_18503,N_19834);
or UO_1480 (O_1480,N_18401,N_18741);
or UO_1481 (O_1481,N_19056,N_19454);
and UO_1482 (O_1482,N_19280,N_19779);
and UO_1483 (O_1483,N_18143,N_18000);
and UO_1484 (O_1484,N_18178,N_18967);
or UO_1485 (O_1485,N_18637,N_19721);
or UO_1486 (O_1486,N_18464,N_18520);
xor UO_1487 (O_1487,N_19157,N_18438);
nor UO_1488 (O_1488,N_19876,N_18855);
nand UO_1489 (O_1489,N_18745,N_18466);
nor UO_1490 (O_1490,N_18246,N_18643);
xnor UO_1491 (O_1491,N_19229,N_18314);
and UO_1492 (O_1492,N_18074,N_19309);
nand UO_1493 (O_1493,N_19872,N_19283);
and UO_1494 (O_1494,N_19862,N_19319);
and UO_1495 (O_1495,N_18631,N_19690);
or UO_1496 (O_1496,N_18816,N_18561);
xor UO_1497 (O_1497,N_18210,N_19435);
nand UO_1498 (O_1498,N_19314,N_18017);
or UO_1499 (O_1499,N_19428,N_18950);
and UO_1500 (O_1500,N_19230,N_19193);
and UO_1501 (O_1501,N_19615,N_19755);
nand UO_1502 (O_1502,N_18000,N_19627);
and UO_1503 (O_1503,N_19270,N_18921);
nand UO_1504 (O_1504,N_19248,N_18545);
xor UO_1505 (O_1505,N_19762,N_19883);
nor UO_1506 (O_1506,N_19974,N_19672);
nor UO_1507 (O_1507,N_19525,N_18564);
and UO_1508 (O_1508,N_18592,N_19679);
nor UO_1509 (O_1509,N_19927,N_18142);
or UO_1510 (O_1510,N_19473,N_18556);
nand UO_1511 (O_1511,N_19505,N_19924);
or UO_1512 (O_1512,N_19572,N_18327);
nor UO_1513 (O_1513,N_19090,N_19521);
nand UO_1514 (O_1514,N_18234,N_19694);
and UO_1515 (O_1515,N_19775,N_18186);
or UO_1516 (O_1516,N_19360,N_18318);
or UO_1517 (O_1517,N_19804,N_19242);
nand UO_1518 (O_1518,N_18972,N_19842);
nand UO_1519 (O_1519,N_18589,N_19924);
and UO_1520 (O_1520,N_19854,N_18184);
nand UO_1521 (O_1521,N_18496,N_19879);
xnor UO_1522 (O_1522,N_19720,N_18125);
and UO_1523 (O_1523,N_18781,N_19195);
nand UO_1524 (O_1524,N_19256,N_19794);
and UO_1525 (O_1525,N_18450,N_18271);
and UO_1526 (O_1526,N_18018,N_19322);
or UO_1527 (O_1527,N_18223,N_18845);
or UO_1528 (O_1528,N_19784,N_18170);
or UO_1529 (O_1529,N_19208,N_18038);
and UO_1530 (O_1530,N_19236,N_19191);
or UO_1531 (O_1531,N_18672,N_18839);
nor UO_1532 (O_1532,N_19458,N_18811);
or UO_1533 (O_1533,N_18798,N_19776);
xnor UO_1534 (O_1534,N_18808,N_19547);
nor UO_1535 (O_1535,N_19322,N_19569);
or UO_1536 (O_1536,N_18348,N_19268);
and UO_1537 (O_1537,N_19230,N_18647);
nand UO_1538 (O_1538,N_19050,N_19742);
or UO_1539 (O_1539,N_19214,N_19837);
or UO_1540 (O_1540,N_19080,N_19752);
and UO_1541 (O_1541,N_19399,N_18495);
xor UO_1542 (O_1542,N_18287,N_18441);
or UO_1543 (O_1543,N_19106,N_19394);
nor UO_1544 (O_1544,N_19053,N_18222);
nor UO_1545 (O_1545,N_18082,N_19419);
xor UO_1546 (O_1546,N_19121,N_18321);
xnor UO_1547 (O_1547,N_19727,N_18266);
nand UO_1548 (O_1548,N_19037,N_18889);
nor UO_1549 (O_1549,N_18265,N_18491);
nand UO_1550 (O_1550,N_18176,N_18203);
or UO_1551 (O_1551,N_18899,N_19824);
nor UO_1552 (O_1552,N_19556,N_18552);
and UO_1553 (O_1553,N_19370,N_18718);
and UO_1554 (O_1554,N_19715,N_18390);
nor UO_1555 (O_1555,N_18196,N_19721);
nor UO_1556 (O_1556,N_18472,N_19328);
nand UO_1557 (O_1557,N_18516,N_18608);
and UO_1558 (O_1558,N_18504,N_18947);
nand UO_1559 (O_1559,N_18459,N_18730);
nor UO_1560 (O_1560,N_18422,N_18699);
xnor UO_1561 (O_1561,N_18909,N_18964);
or UO_1562 (O_1562,N_18273,N_19547);
and UO_1563 (O_1563,N_19067,N_19686);
or UO_1564 (O_1564,N_18188,N_18566);
nand UO_1565 (O_1565,N_19610,N_19387);
or UO_1566 (O_1566,N_19091,N_18154);
and UO_1567 (O_1567,N_18225,N_18916);
xor UO_1568 (O_1568,N_18180,N_18693);
xnor UO_1569 (O_1569,N_18280,N_19518);
nand UO_1570 (O_1570,N_18426,N_19912);
or UO_1571 (O_1571,N_19128,N_19852);
or UO_1572 (O_1572,N_18647,N_18736);
and UO_1573 (O_1573,N_19839,N_19549);
xnor UO_1574 (O_1574,N_18847,N_18372);
xnor UO_1575 (O_1575,N_19444,N_19229);
or UO_1576 (O_1576,N_18909,N_18025);
nor UO_1577 (O_1577,N_18195,N_18916);
or UO_1578 (O_1578,N_19518,N_18888);
nor UO_1579 (O_1579,N_18680,N_19164);
or UO_1580 (O_1580,N_19891,N_19363);
xnor UO_1581 (O_1581,N_18400,N_19802);
and UO_1582 (O_1582,N_18289,N_18612);
nor UO_1583 (O_1583,N_19619,N_19375);
nor UO_1584 (O_1584,N_18757,N_18807);
nand UO_1585 (O_1585,N_18991,N_18100);
nand UO_1586 (O_1586,N_19596,N_18359);
nand UO_1587 (O_1587,N_18584,N_19360);
nor UO_1588 (O_1588,N_18843,N_18516);
xor UO_1589 (O_1589,N_19348,N_18514);
or UO_1590 (O_1590,N_18777,N_19657);
nor UO_1591 (O_1591,N_18257,N_18302);
or UO_1592 (O_1592,N_19907,N_19025);
nor UO_1593 (O_1593,N_19304,N_18547);
and UO_1594 (O_1594,N_19850,N_19636);
nor UO_1595 (O_1595,N_18049,N_18782);
and UO_1596 (O_1596,N_18056,N_19169);
nand UO_1597 (O_1597,N_19347,N_18837);
nand UO_1598 (O_1598,N_18390,N_18755);
nor UO_1599 (O_1599,N_18834,N_18668);
nand UO_1600 (O_1600,N_19173,N_18297);
nor UO_1601 (O_1601,N_18942,N_18387);
or UO_1602 (O_1602,N_19513,N_19528);
nor UO_1603 (O_1603,N_18418,N_18247);
nand UO_1604 (O_1604,N_18649,N_19008);
xnor UO_1605 (O_1605,N_19174,N_19841);
nor UO_1606 (O_1606,N_19719,N_19871);
nand UO_1607 (O_1607,N_18021,N_19568);
xnor UO_1608 (O_1608,N_19919,N_19226);
nor UO_1609 (O_1609,N_19929,N_18640);
nand UO_1610 (O_1610,N_19807,N_19870);
xor UO_1611 (O_1611,N_18010,N_18528);
and UO_1612 (O_1612,N_18550,N_18421);
nor UO_1613 (O_1613,N_18491,N_18165);
nand UO_1614 (O_1614,N_18929,N_18510);
nand UO_1615 (O_1615,N_18234,N_18540);
nand UO_1616 (O_1616,N_19271,N_18604);
or UO_1617 (O_1617,N_19808,N_19271);
xor UO_1618 (O_1618,N_18302,N_19046);
xor UO_1619 (O_1619,N_19859,N_18968);
nor UO_1620 (O_1620,N_18211,N_18196);
and UO_1621 (O_1621,N_18659,N_18207);
nor UO_1622 (O_1622,N_19975,N_19499);
nand UO_1623 (O_1623,N_18510,N_19705);
or UO_1624 (O_1624,N_19332,N_19983);
or UO_1625 (O_1625,N_18563,N_19995);
or UO_1626 (O_1626,N_19488,N_19868);
and UO_1627 (O_1627,N_19924,N_18921);
xnor UO_1628 (O_1628,N_19359,N_18941);
and UO_1629 (O_1629,N_18261,N_18382);
nor UO_1630 (O_1630,N_18100,N_18193);
nor UO_1631 (O_1631,N_19970,N_18018);
and UO_1632 (O_1632,N_18583,N_18905);
or UO_1633 (O_1633,N_18328,N_18507);
nor UO_1634 (O_1634,N_18785,N_19290);
xnor UO_1635 (O_1635,N_19010,N_19907);
nand UO_1636 (O_1636,N_19346,N_19515);
nand UO_1637 (O_1637,N_18258,N_19335);
or UO_1638 (O_1638,N_19536,N_18327);
nand UO_1639 (O_1639,N_19616,N_19660);
or UO_1640 (O_1640,N_18192,N_19339);
xor UO_1641 (O_1641,N_18530,N_18049);
nand UO_1642 (O_1642,N_19775,N_19921);
nor UO_1643 (O_1643,N_18998,N_18066);
nor UO_1644 (O_1644,N_18749,N_18009);
and UO_1645 (O_1645,N_18785,N_19518);
and UO_1646 (O_1646,N_18687,N_19564);
nand UO_1647 (O_1647,N_19470,N_18353);
nand UO_1648 (O_1648,N_18913,N_18320);
nand UO_1649 (O_1649,N_19428,N_19266);
xnor UO_1650 (O_1650,N_18046,N_19233);
nor UO_1651 (O_1651,N_19554,N_18812);
nand UO_1652 (O_1652,N_19872,N_18260);
or UO_1653 (O_1653,N_18226,N_18115);
or UO_1654 (O_1654,N_19116,N_19617);
nor UO_1655 (O_1655,N_18314,N_18049);
and UO_1656 (O_1656,N_19622,N_18348);
or UO_1657 (O_1657,N_18232,N_19262);
nor UO_1658 (O_1658,N_18956,N_18923);
or UO_1659 (O_1659,N_19064,N_18273);
nor UO_1660 (O_1660,N_19989,N_18022);
nor UO_1661 (O_1661,N_18270,N_19116);
and UO_1662 (O_1662,N_18760,N_19111);
xnor UO_1663 (O_1663,N_18328,N_18122);
or UO_1664 (O_1664,N_19979,N_18505);
and UO_1665 (O_1665,N_18045,N_18225);
nand UO_1666 (O_1666,N_19765,N_19641);
nor UO_1667 (O_1667,N_19894,N_19934);
or UO_1668 (O_1668,N_18366,N_19706);
or UO_1669 (O_1669,N_18459,N_18038);
nor UO_1670 (O_1670,N_19153,N_18666);
and UO_1671 (O_1671,N_19725,N_18983);
or UO_1672 (O_1672,N_18028,N_18761);
and UO_1673 (O_1673,N_19774,N_19225);
or UO_1674 (O_1674,N_18878,N_19569);
nand UO_1675 (O_1675,N_18259,N_19539);
or UO_1676 (O_1676,N_18674,N_18893);
nand UO_1677 (O_1677,N_18349,N_18029);
or UO_1678 (O_1678,N_18370,N_19487);
and UO_1679 (O_1679,N_18459,N_18112);
nor UO_1680 (O_1680,N_19242,N_19370);
nor UO_1681 (O_1681,N_19148,N_18893);
or UO_1682 (O_1682,N_18539,N_19323);
nand UO_1683 (O_1683,N_19077,N_18600);
and UO_1684 (O_1684,N_19928,N_18771);
nand UO_1685 (O_1685,N_19143,N_19254);
and UO_1686 (O_1686,N_18388,N_18902);
and UO_1687 (O_1687,N_18791,N_18528);
or UO_1688 (O_1688,N_19079,N_19509);
xor UO_1689 (O_1689,N_19781,N_19247);
and UO_1690 (O_1690,N_19777,N_19957);
nand UO_1691 (O_1691,N_19148,N_19858);
nor UO_1692 (O_1692,N_19058,N_18231);
and UO_1693 (O_1693,N_19609,N_19873);
nor UO_1694 (O_1694,N_18281,N_19622);
or UO_1695 (O_1695,N_19753,N_18249);
nor UO_1696 (O_1696,N_18232,N_19506);
and UO_1697 (O_1697,N_18726,N_18400);
xnor UO_1698 (O_1698,N_19950,N_19322);
or UO_1699 (O_1699,N_18686,N_18151);
nand UO_1700 (O_1700,N_19906,N_19651);
and UO_1701 (O_1701,N_19440,N_18281);
xor UO_1702 (O_1702,N_19694,N_18542);
or UO_1703 (O_1703,N_18752,N_18821);
xor UO_1704 (O_1704,N_18594,N_18916);
nor UO_1705 (O_1705,N_19868,N_18963);
or UO_1706 (O_1706,N_19869,N_19675);
or UO_1707 (O_1707,N_19868,N_18054);
xor UO_1708 (O_1708,N_19575,N_19418);
nand UO_1709 (O_1709,N_18594,N_19187);
or UO_1710 (O_1710,N_18146,N_18612);
or UO_1711 (O_1711,N_18663,N_18787);
nand UO_1712 (O_1712,N_19933,N_18446);
nor UO_1713 (O_1713,N_18837,N_18494);
nor UO_1714 (O_1714,N_19004,N_19009);
and UO_1715 (O_1715,N_19531,N_18060);
nor UO_1716 (O_1716,N_19920,N_18237);
and UO_1717 (O_1717,N_18282,N_18768);
xnor UO_1718 (O_1718,N_19206,N_18461);
or UO_1719 (O_1719,N_19201,N_19419);
nand UO_1720 (O_1720,N_18713,N_19412);
nand UO_1721 (O_1721,N_19737,N_19705);
or UO_1722 (O_1722,N_18264,N_18906);
and UO_1723 (O_1723,N_19579,N_19316);
nor UO_1724 (O_1724,N_19398,N_18708);
xnor UO_1725 (O_1725,N_18938,N_19543);
nand UO_1726 (O_1726,N_19964,N_19156);
nor UO_1727 (O_1727,N_19092,N_18877);
nor UO_1728 (O_1728,N_18180,N_18984);
nand UO_1729 (O_1729,N_19979,N_19026);
and UO_1730 (O_1730,N_19649,N_18434);
and UO_1731 (O_1731,N_19549,N_18194);
nor UO_1732 (O_1732,N_18991,N_19648);
or UO_1733 (O_1733,N_19085,N_19972);
nor UO_1734 (O_1734,N_19680,N_19482);
nand UO_1735 (O_1735,N_18255,N_19635);
nand UO_1736 (O_1736,N_18440,N_19939);
or UO_1737 (O_1737,N_19140,N_19546);
or UO_1738 (O_1738,N_19656,N_18694);
xnor UO_1739 (O_1739,N_19580,N_19136);
nor UO_1740 (O_1740,N_19915,N_18366);
xnor UO_1741 (O_1741,N_19374,N_19502);
nor UO_1742 (O_1742,N_19847,N_18872);
nand UO_1743 (O_1743,N_19323,N_19594);
and UO_1744 (O_1744,N_18704,N_19360);
nor UO_1745 (O_1745,N_19077,N_19627);
nand UO_1746 (O_1746,N_19147,N_19585);
nor UO_1747 (O_1747,N_19191,N_19385);
and UO_1748 (O_1748,N_18015,N_18301);
and UO_1749 (O_1749,N_18820,N_19232);
nor UO_1750 (O_1750,N_18370,N_18320);
nor UO_1751 (O_1751,N_18451,N_18098);
xnor UO_1752 (O_1752,N_19910,N_19288);
nand UO_1753 (O_1753,N_19805,N_18688);
nand UO_1754 (O_1754,N_18894,N_19739);
and UO_1755 (O_1755,N_19700,N_19688);
xor UO_1756 (O_1756,N_18929,N_19679);
nor UO_1757 (O_1757,N_19740,N_19173);
or UO_1758 (O_1758,N_19322,N_19208);
nand UO_1759 (O_1759,N_18657,N_18741);
or UO_1760 (O_1760,N_18969,N_18436);
and UO_1761 (O_1761,N_18111,N_19630);
nor UO_1762 (O_1762,N_19998,N_18840);
xor UO_1763 (O_1763,N_19055,N_19720);
and UO_1764 (O_1764,N_19842,N_18104);
nand UO_1765 (O_1765,N_19908,N_18610);
nand UO_1766 (O_1766,N_19797,N_19292);
and UO_1767 (O_1767,N_18225,N_19436);
and UO_1768 (O_1768,N_18457,N_18912);
and UO_1769 (O_1769,N_18504,N_19055);
or UO_1770 (O_1770,N_19234,N_18557);
and UO_1771 (O_1771,N_19565,N_19174);
or UO_1772 (O_1772,N_19896,N_19173);
or UO_1773 (O_1773,N_18380,N_19615);
and UO_1774 (O_1774,N_18387,N_18738);
and UO_1775 (O_1775,N_19006,N_19646);
nor UO_1776 (O_1776,N_18820,N_18865);
and UO_1777 (O_1777,N_18663,N_18831);
nand UO_1778 (O_1778,N_18548,N_18930);
and UO_1779 (O_1779,N_18749,N_19604);
and UO_1780 (O_1780,N_18567,N_19956);
nor UO_1781 (O_1781,N_19593,N_19222);
and UO_1782 (O_1782,N_19990,N_19323);
and UO_1783 (O_1783,N_19703,N_19176);
nor UO_1784 (O_1784,N_18652,N_18668);
or UO_1785 (O_1785,N_18371,N_18817);
nand UO_1786 (O_1786,N_18670,N_18488);
nor UO_1787 (O_1787,N_19107,N_19480);
nand UO_1788 (O_1788,N_18801,N_18277);
nand UO_1789 (O_1789,N_19221,N_19853);
nor UO_1790 (O_1790,N_18000,N_18054);
or UO_1791 (O_1791,N_18341,N_18073);
nor UO_1792 (O_1792,N_18938,N_19754);
nand UO_1793 (O_1793,N_19993,N_18503);
nor UO_1794 (O_1794,N_18342,N_18130);
or UO_1795 (O_1795,N_18255,N_19851);
nand UO_1796 (O_1796,N_18244,N_18587);
and UO_1797 (O_1797,N_18353,N_19851);
and UO_1798 (O_1798,N_18284,N_18315);
and UO_1799 (O_1799,N_19949,N_18944);
nand UO_1800 (O_1800,N_18671,N_18119);
nor UO_1801 (O_1801,N_18466,N_19237);
and UO_1802 (O_1802,N_19024,N_19195);
nand UO_1803 (O_1803,N_18837,N_19392);
nand UO_1804 (O_1804,N_19713,N_19029);
or UO_1805 (O_1805,N_18415,N_19456);
or UO_1806 (O_1806,N_19275,N_19910);
nand UO_1807 (O_1807,N_18889,N_19444);
nor UO_1808 (O_1808,N_19968,N_19982);
nand UO_1809 (O_1809,N_18609,N_18389);
nand UO_1810 (O_1810,N_18994,N_19166);
nor UO_1811 (O_1811,N_19493,N_19181);
nor UO_1812 (O_1812,N_19697,N_19310);
or UO_1813 (O_1813,N_18523,N_18516);
xor UO_1814 (O_1814,N_19166,N_19133);
nor UO_1815 (O_1815,N_19142,N_18861);
nor UO_1816 (O_1816,N_18988,N_18435);
nand UO_1817 (O_1817,N_18658,N_18223);
or UO_1818 (O_1818,N_19210,N_18079);
and UO_1819 (O_1819,N_18286,N_19496);
nor UO_1820 (O_1820,N_18580,N_18125);
xor UO_1821 (O_1821,N_19584,N_18971);
and UO_1822 (O_1822,N_19342,N_18766);
nor UO_1823 (O_1823,N_18233,N_18352);
or UO_1824 (O_1824,N_18383,N_19821);
and UO_1825 (O_1825,N_18919,N_19329);
nor UO_1826 (O_1826,N_19066,N_18147);
nand UO_1827 (O_1827,N_19823,N_18755);
or UO_1828 (O_1828,N_19151,N_18381);
nand UO_1829 (O_1829,N_18924,N_19872);
nand UO_1830 (O_1830,N_19209,N_18259);
and UO_1831 (O_1831,N_18036,N_18609);
or UO_1832 (O_1832,N_18812,N_19578);
nand UO_1833 (O_1833,N_18970,N_19669);
nor UO_1834 (O_1834,N_19520,N_19097);
nor UO_1835 (O_1835,N_18384,N_18080);
nor UO_1836 (O_1836,N_19017,N_18115);
or UO_1837 (O_1837,N_19231,N_18371);
and UO_1838 (O_1838,N_19331,N_18961);
nor UO_1839 (O_1839,N_19908,N_19413);
nor UO_1840 (O_1840,N_18643,N_18811);
xnor UO_1841 (O_1841,N_19140,N_19021);
nor UO_1842 (O_1842,N_18195,N_18877);
xor UO_1843 (O_1843,N_18019,N_19592);
nor UO_1844 (O_1844,N_19290,N_19020);
and UO_1845 (O_1845,N_19312,N_19719);
or UO_1846 (O_1846,N_19769,N_19876);
and UO_1847 (O_1847,N_19199,N_18133);
nand UO_1848 (O_1848,N_19370,N_18702);
and UO_1849 (O_1849,N_19243,N_18234);
nand UO_1850 (O_1850,N_18432,N_19504);
nor UO_1851 (O_1851,N_18040,N_19363);
or UO_1852 (O_1852,N_18591,N_19924);
and UO_1853 (O_1853,N_19045,N_18454);
xnor UO_1854 (O_1854,N_19422,N_19800);
nand UO_1855 (O_1855,N_18801,N_18642);
or UO_1856 (O_1856,N_18075,N_19833);
nand UO_1857 (O_1857,N_19078,N_19153);
nand UO_1858 (O_1858,N_19596,N_18596);
nor UO_1859 (O_1859,N_19352,N_18616);
and UO_1860 (O_1860,N_18006,N_18150);
xnor UO_1861 (O_1861,N_18328,N_19276);
nor UO_1862 (O_1862,N_18364,N_18305);
nor UO_1863 (O_1863,N_19803,N_18281);
and UO_1864 (O_1864,N_18085,N_18747);
nor UO_1865 (O_1865,N_19613,N_18752);
or UO_1866 (O_1866,N_18395,N_18351);
and UO_1867 (O_1867,N_19319,N_18739);
or UO_1868 (O_1868,N_19125,N_18712);
and UO_1869 (O_1869,N_19303,N_18073);
nand UO_1870 (O_1870,N_18203,N_18199);
and UO_1871 (O_1871,N_18751,N_18378);
nor UO_1872 (O_1872,N_19989,N_19108);
or UO_1873 (O_1873,N_18222,N_18422);
and UO_1874 (O_1874,N_19575,N_18174);
xor UO_1875 (O_1875,N_18700,N_19975);
or UO_1876 (O_1876,N_19951,N_19188);
and UO_1877 (O_1877,N_19425,N_18095);
nand UO_1878 (O_1878,N_18925,N_18321);
nor UO_1879 (O_1879,N_19124,N_19284);
nor UO_1880 (O_1880,N_19103,N_18828);
and UO_1881 (O_1881,N_18455,N_19648);
nand UO_1882 (O_1882,N_19567,N_18277);
or UO_1883 (O_1883,N_18704,N_19458);
or UO_1884 (O_1884,N_18558,N_19651);
nor UO_1885 (O_1885,N_18041,N_19866);
nor UO_1886 (O_1886,N_18053,N_18807);
nand UO_1887 (O_1887,N_19749,N_19417);
nor UO_1888 (O_1888,N_19363,N_19893);
nand UO_1889 (O_1889,N_19327,N_18214);
nor UO_1890 (O_1890,N_18714,N_18307);
nor UO_1891 (O_1891,N_18220,N_18900);
xor UO_1892 (O_1892,N_19197,N_18033);
and UO_1893 (O_1893,N_18182,N_18418);
nor UO_1894 (O_1894,N_18053,N_19344);
nand UO_1895 (O_1895,N_19524,N_18260);
or UO_1896 (O_1896,N_19069,N_18311);
or UO_1897 (O_1897,N_18536,N_18112);
nor UO_1898 (O_1898,N_19605,N_18964);
nand UO_1899 (O_1899,N_18865,N_19053);
and UO_1900 (O_1900,N_18372,N_19054);
or UO_1901 (O_1901,N_19766,N_18749);
xnor UO_1902 (O_1902,N_19741,N_19749);
nor UO_1903 (O_1903,N_19170,N_18941);
or UO_1904 (O_1904,N_18002,N_19317);
xnor UO_1905 (O_1905,N_18963,N_18622);
and UO_1906 (O_1906,N_18523,N_18759);
and UO_1907 (O_1907,N_18286,N_18732);
nor UO_1908 (O_1908,N_19155,N_19369);
nor UO_1909 (O_1909,N_19648,N_19431);
and UO_1910 (O_1910,N_19311,N_19012);
or UO_1911 (O_1911,N_19146,N_19627);
or UO_1912 (O_1912,N_18622,N_19369);
or UO_1913 (O_1913,N_18551,N_19626);
and UO_1914 (O_1914,N_19377,N_18571);
nor UO_1915 (O_1915,N_18486,N_18989);
nor UO_1916 (O_1916,N_18595,N_18275);
and UO_1917 (O_1917,N_19336,N_18698);
or UO_1918 (O_1918,N_18490,N_18107);
nor UO_1919 (O_1919,N_18241,N_19476);
nor UO_1920 (O_1920,N_18456,N_18321);
nand UO_1921 (O_1921,N_18918,N_19996);
xnor UO_1922 (O_1922,N_19768,N_19902);
and UO_1923 (O_1923,N_18520,N_18610);
nor UO_1924 (O_1924,N_18784,N_19679);
nand UO_1925 (O_1925,N_19171,N_18926);
or UO_1926 (O_1926,N_18960,N_18523);
and UO_1927 (O_1927,N_18941,N_19070);
and UO_1928 (O_1928,N_19906,N_19484);
or UO_1929 (O_1929,N_18723,N_19172);
nand UO_1930 (O_1930,N_18732,N_19360);
or UO_1931 (O_1931,N_18898,N_19354);
or UO_1932 (O_1932,N_19442,N_18180);
nand UO_1933 (O_1933,N_19715,N_18657);
nor UO_1934 (O_1934,N_18324,N_19774);
nor UO_1935 (O_1935,N_19034,N_19122);
or UO_1936 (O_1936,N_19162,N_19371);
or UO_1937 (O_1937,N_18059,N_19586);
and UO_1938 (O_1938,N_18094,N_19903);
xor UO_1939 (O_1939,N_19294,N_18180);
nand UO_1940 (O_1940,N_19135,N_18058);
or UO_1941 (O_1941,N_18352,N_19252);
nor UO_1942 (O_1942,N_19076,N_18983);
and UO_1943 (O_1943,N_18943,N_19827);
nand UO_1944 (O_1944,N_18602,N_19884);
or UO_1945 (O_1945,N_18191,N_19694);
nor UO_1946 (O_1946,N_19773,N_19395);
xor UO_1947 (O_1947,N_19521,N_18606);
nand UO_1948 (O_1948,N_18183,N_18145);
nand UO_1949 (O_1949,N_18862,N_19569);
nor UO_1950 (O_1950,N_19648,N_18793);
or UO_1951 (O_1951,N_18863,N_19073);
and UO_1952 (O_1952,N_18613,N_19090);
nor UO_1953 (O_1953,N_18934,N_18088);
nand UO_1954 (O_1954,N_18076,N_19864);
nand UO_1955 (O_1955,N_19335,N_18729);
or UO_1956 (O_1956,N_19596,N_18876);
and UO_1957 (O_1957,N_19935,N_18435);
or UO_1958 (O_1958,N_19317,N_19146);
nor UO_1959 (O_1959,N_18064,N_18977);
nand UO_1960 (O_1960,N_18840,N_18634);
nand UO_1961 (O_1961,N_18453,N_18379);
nand UO_1962 (O_1962,N_18840,N_19173);
and UO_1963 (O_1963,N_18605,N_19823);
and UO_1964 (O_1964,N_19036,N_18971);
nand UO_1965 (O_1965,N_19459,N_19243);
or UO_1966 (O_1966,N_18757,N_19177);
nand UO_1967 (O_1967,N_19157,N_18104);
nand UO_1968 (O_1968,N_19893,N_19026);
or UO_1969 (O_1969,N_19286,N_18690);
nand UO_1970 (O_1970,N_18952,N_19193);
and UO_1971 (O_1971,N_19624,N_18653);
nor UO_1972 (O_1972,N_18170,N_19352);
nor UO_1973 (O_1973,N_18832,N_19068);
xor UO_1974 (O_1974,N_19879,N_19995);
and UO_1975 (O_1975,N_18902,N_18041);
and UO_1976 (O_1976,N_18166,N_18483);
nor UO_1977 (O_1977,N_19548,N_19844);
or UO_1978 (O_1978,N_18449,N_18770);
nand UO_1979 (O_1979,N_18176,N_19663);
or UO_1980 (O_1980,N_19481,N_19506);
or UO_1981 (O_1981,N_19883,N_18757);
and UO_1982 (O_1982,N_18898,N_18865);
nand UO_1983 (O_1983,N_19230,N_18325);
xor UO_1984 (O_1984,N_19819,N_19313);
and UO_1985 (O_1985,N_19248,N_19465);
or UO_1986 (O_1986,N_19040,N_18709);
and UO_1987 (O_1987,N_19036,N_18298);
nor UO_1988 (O_1988,N_18210,N_18582);
nand UO_1989 (O_1989,N_19251,N_19833);
or UO_1990 (O_1990,N_18722,N_19013);
nor UO_1991 (O_1991,N_18861,N_19227);
and UO_1992 (O_1992,N_18914,N_19051);
or UO_1993 (O_1993,N_18496,N_18846);
nand UO_1994 (O_1994,N_19853,N_18696);
nand UO_1995 (O_1995,N_19596,N_18086);
and UO_1996 (O_1996,N_19474,N_19651);
and UO_1997 (O_1997,N_18535,N_19733);
or UO_1998 (O_1998,N_18751,N_19490);
and UO_1999 (O_1999,N_19347,N_18345);
nand UO_2000 (O_2000,N_18733,N_18725);
or UO_2001 (O_2001,N_18111,N_19039);
nor UO_2002 (O_2002,N_18615,N_18369);
and UO_2003 (O_2003,N_18189,N_18997);
or UO_2004 (O_2004,N_18021,N_18053);
nand UO_2005 (O_2005,N_18938,N_19351);
or UO_2006 (O_2006,N_19400,N_18715);
and UO_2007 (O_2007,N_18863,N_18026);
and UO_2008 (O_2008,N_18062,N_19136);
xor UO_2009 (O_2009,N_19348,N_19645);
nand UO_2010 (O_2010,N_18341,N_19215);
or UO_2011 (O_2011,N_19599,N_18173);
or UO_2012 (O_2012,N_18722,N_19468);
and UO_2013 (O_2013,N_18420,N_19684);
and UO_2014 (O_2014,N_18151,N_18450);
nand UO_2015 (O_2015,N_18716,N_18940);
nor UO_2016 (O_2016,N_19316,N_18903);
or UO_2017 (O_2017,N_18091,N_19227);
and UO_2018 (O_2018,N_19056,N_19342);
nand UO_2019 (O_2019,N_18882,N_19726);
xnor UO_2020 (O_2020,N_18063,N_19391);
or UO_2021 (O_2021,N_18332,N_19964);
nor UO_2022 (O_2022,N_19020,N_19450);
and UO_2023 (O_2023,N_18646,N_19664);
nand UO_2024 (O_2024,N_19742,N_18612);
xor UO_2025 (O_2025,N_19759,N_19234);
and UO_2026 (O_2026,N_18701,N_18055);
nor UO_2027 (O_2027,N_18325,N_19987);
or UO_2028 (O_2028,N_19471,N_18661);
nor UO_2029 (O_2029,N_18235,N_18685);
nor UO_2030 (O_2030,N_18798,N_19301);
nand UO_2031 (O_2031,N_18263,N_18028);
nor UO_2032 (O_2032,N_19592,N_19596);
and UO_2033 (O_2033,N_19458,N_19678);
or UO_2034 (O_2034,N_19091,N_19248);
and UO_2035 (O_2035,N_18502,N_18627);
and UO_2036 (O_2036,N_18936,N_19855);
xor UO_2037 (O_2037,N_18089,N_19579);
nand UO_2038 (O_2038,N_19415,N_18686);
and UO_2039 (O_2039,N_19999,N_18221);
and UO_2040 (O_2040,N_19950,N_18281);
or UO_2041 (O_2041,N_18953,N_18601);
and UO_2042 (O_2042,N_18543,N_19166);
and UO_2043 (O_2043,N_19570,N_18852);
nand UO_2044 (O_2044,N_18284,N_18152);
nor UO_2045 (O_2045,N_18054,N_19344);
or UO_2046 (O_2046,N_18169,N_18990);
nand UO_2047 (O_2047,N_19664,N_19643);
or UO_2048 (O_2048,N_18870,N_19367);
nor UO_2049 (O_2049,N_19089,N_19766);
or UO_2050 (O_2050,N_19989,N_18802);
nand UO_2051 (O_2051,N_19945,N_18350);
and UO_2052 (O_2052,N_19282,N_18242);
nor UO_2053 (O_2053,N_18824,N_19604);
nand UO_2054 (O_2054,N_19402,N_19214);
and UO_2055 (O_2055,N_18627,N_19757);
or UO_2056 (O_2056,N_19380,N_19723);
nand UO_2057 (O_2057,N_19646,N_18503);
nand UO_2058 (O_2058,N_18531,N_19105);
nand UO_2059 (O_2059,N_19424,N_19923);
and UO_2060 (O_2060,N_19507,N_18051);
or UO_2061 (O_2061,N_18573,N_19725);
and UO_2062 (O_2062,N_18408,N_19292);
nand UO_2063 (O_2063,N_19249,N_18204);
nand UO_2064 (O_2064,N_18319,N_19832);
and UO_2065 (O_2065,N_19565,N_19201);
or UO_2066 (O_2066,N_19793,N_19389);
xnor UO_2067 (O_2067,N_18606,N_19478);
or UO_2068 (O_2068,N_19630,N_18251);
nor UO_2069 (O_2069,N_18055,N_19030);
nand UO_2070 (O_2070,N_18716,N_18070);
nor UO_2071 (O_2071,N_19917,N_18215);
or UO_2072 (O_2072,N_19261,N_18204);
or UO_2073 (O_2073,N_19773,N_18162);
nor UO_2074 (O_2074,N_18075,N_18724);
nor UO_2075 (O_2075,N_19922,N_19009);
nand UO_2076 (O_2076,N_19874,N_19760);
or UO_2077 (O_2077,N_19678,N_19904);
and UO_2078 (O_2078,N_19472,N_18785);
nor UO_2079 (O_2079,N_19651,N_18427);
or UO_2080 (O_2080,N_19096,N_19059);
and UO_2081 (O_2081,N_19541,N_18512);
nor UO_2082 (O_2082,N_19477,N_19117);
xor UO_2083 (O_2083,N_18279,N_19384);
xor UO_2084 (O_2084,N_19712,N_18318);
or UO_2085 (O_2085,N_18396,N_18450);
nor UO_2086 (O_2086,N_19105,N_18611);
or UO_2087 (O_2087,N_18088,N_19785);
and UO_2088 (O_2088,N_19814,N_19813);
nand UO_2089 (O_2089,N_18643,N_19746);
nand UO_2090 (O_2090,N_19152,N_19227);
nor UO_2091 (O_2091,N_19498,N_19319);
nor UO_2092 (O_2092,N_18811,N_19589);
nor UO_2093 (O_2093,N_18094,N_19600);
nand UO_2094 (O_2094,N_19748,N_18854);
nand UO_2095 (O_2095,N_19554,N_18739);
and UO_2096 (O_2096,N_18547,N_19712);
or UO_2097 (O_2097,N_18159,N_18200);
and UO_2098 (O_2098,N_18165,N_18621);
or UO_2099 (O_2099,N_18723,N_19613);
nor UO_2100 (O_2100,N_18804,N_19539);
nand UO_2101 (O_2101,N_18458,N_19191);
nand UO_2102 (O_2102,N_18324,N_18227);
or UO_2103 (O_2103,N_19907,N_18054);
or UO_2104 (O_2104,N_18168,N_18196);
or UO_2105 (O_2105,N_19329,N_19416);
xor UO_2106 (O_2106,N_18948,N_19910);
or UO_2107 (O_2107,N_18548,N_19937);
nor UO_2108 (O_2108,N_19434,N_19435);
xnor UO_2109 (O_2109,N_19522,N_18983);
and UO_2110 (O_2110,N_18755,N_18909);
nor UO_2111 (O_2111,N_18024,N_19729);
and UO_2112 (O_2112,N_19474,N_19743);
or UO_2113 (O_2113,N_18185,N_19675);
nor UO_2114 (O_2114,N_18207,N_18389);
or UO_2115 (O_2115,N_19394,N_18249);
nand UO_2116 (O_2116,N_19303,N_19990);
nor UO_2117 (O_2117,N_18874,N_18936);
nor UO_2118 (O_2118,N_18201,N_19300);
or UO_2119 (O_2119,N_19400,N_18221);
nor UO_2120 (O_2120,N_19452,N_18667);
or UO_2121 (O_2121,N_18144,N_19159);
or UO_2122 (O_2122,N_18752,N_18619);
xor UO_2123 (O_2123,N_19942,N_19951);
nand UO_2124 (O_2124,N_19037,N_18412);
xnor UO_2125 (O_2125,N_18543,N_18629);
nor UO_2126 (O_2126,N_18201,N_19861);
or UO_2127 (O_2127,N_19301,N_19458);
and UO_2128 (O_2128,N_19495,N_19583);
nand UO_2129 (O_2129,N_19026,N_19624);
nor UO_2130 (O_2130,N_19109,N_18299);
or UO_2131 (O_2131,N_19170,N_18922);
or UO_2132 (O_2132,N_19606,N_19983);
nand UO_2133 (O_2133,N_18706,N_18502);
or UO_2134 (O_2134,N_18947,N_19168);
or UO_2135 (O_2135,N_19385,N_18060);
or UO_2136 (O_2136,N_18579,N_19306);
nor UO_2137 (O_2137,N_18329,N_19777);
nand UO_2138 (O_2138,N_18497,N_19465);
and UO_2139 (O_2139,N_18314,N_18172);
and UO_2140 (O_2140,N_19629,N_19552);
nor UO_2141 (O_2141,N_19765,N_19793);
nor UO_2142 (O_2142,N_19597,N_19845);
xnor UO_2143 (O_2143,N_19250,N_18877);
nor UO_2144 (O_2144,N_19185,N_19187);
xor UO_2145 (O_2145,N_19617,N_18406);
and UO_2146 (O_2146,N_19215,N_19479);
and UO_2147 (O_2147,N_19309,N_19529);
nand UO_2148 (O_2148,N_18340,N_19762);
and UO_2149 (O_2149,N_19808,N_18226);
xnor UO_2150 (O_2150,N_18607,N_19037);
nand UO_2151 (O_2151,N_18585,N_18426);
nor UO_2152 (O_2152,N_18706,N_18682);
nand UO_2153 (O_2153,N_19807,N_19367);
and UO_2154 (O_2154,N_18143,N_19216);
and UO_2155 (O_2155,N_18081,N_18354);
and UO_2156 (O_2156,N_18093,N_18005);
or UO_2157 (O_2157,N_18391,N_18945);
or UO_2158 (O_2158,N_19461,N_18948);
or UO_2159 (O_2159,N_18934,N_19121);
and UO_2160 (O_2160,N_19347,N_18263);
or UO_2161 (O_2161,N_18665,N_19826);
or UO_2162 (O_2162,N_19819,N_18037);
and UO_2163 (O_2163,N_19790,N_19590);
xor UO_2164 (O_2164,N_18460,N_18938);
nand UO_2165 (O_2165,N_19453,N_19836);
and UO_2166 (O_2166,N_19578,N_18852);
and UO_2167 (O_2167,N_19638,N_19577);
and UO_2168 (O_2168,N_19255,N_18455);
xor UO_2169 (O_2169,N_18890,N_18024);
and UO_2170 (O_2170,N_18020,N_18411);
and UO_2171 (O_2171,N_18440,N_19001);
or UO_2172 (O_2172,N_19974,N_18380);
and UO_2173 (O_2173,N_19717,N_19980);
or UO_2174 (O_2174,N_19159,N_19465);
xnor UO_2175 (O_2175,N_19227,N_19762);
and UO_2176 (O_2176,N_18890,N_18975);
or UO_2177 (O_2177,N_18654,N_19415);
nor UO_2178 (O_2178,N_18954,N_18617);
nor UO_2179 (O_2179,N_19961,N_18451);
nand UO_2180 (O_2180,N_19998,N_18963);
nor UO_2181 (O_2181,N_18889,N_19724);
or UO_2182 (O_2182,N_18537,N_18705);
nand UO_2183 (O_2183,N_18018,N_19107);
xor UO_2184 (O_2184,N_18021,N_19437);
nand UO_2185 (O_2185,N_18636,N_18362);
and UO_2186 (O_2186,N_19474,N_18464);
nand UO_2187 (O_2187,N_18576,N_19998);
nor UO_2188 (O_2188,N_19689,N_18991);
or UO_2189 (O_2189,N_18667,N_19066);
nor UO_2190 (O_2190,N_19862,N_19183);
or UO_2191 (O_2191,N_19532,N_19036);
and UO_2192 (O_2192,N_18841,N_19138);
or UO_2193 (O_2193,N_18535,N_18428);
and UO_2194 (O_2194,N_18608,N_19078);
nor UO_2195 (O_2195,N_19483,N_18968);
xor UO_2196 (O_2196,N_19080,N_19474);
nand UO_2197 (O_2197,N_18319,N_19449);
nor UO_2198 (O_2198,N_19893,N_18042);
nor UO_2199 (O_2199,N_19161,N_18729);
xnor UO_2200 (O_2200,N_19874,N_18645);
nor UO_2201 (O_2201,N_18839,N_18780);
nand UO_2202 (O_2202,N_18151,N_19761);
nand UO_2203 (O_2203,N_18151,N_19021);
nand UO_2204 (O_2204,N_19648,N_19785);
and UO_2205 (O_2205,N_18550,N_19967);
nand UO_2206 (O_2206,N_19017,N_19650);
nand UO_2207 (O_2207,N_19824,N_18077);
nand UO_2208 (O_2208,N_18557,N_18291);
nand UO_2209 (O_2209,N_18003,N_18431);
nand UO_2210 (O_2210,N_18454,N_19815);
or UO_2211 (O_2211,N_19837,N_19169);
or UO_2212 (O_2212,N_19120,N_19599);
or UO_2213 (O_2213,N_19160,N_19917);
nor UO_2214 (O_2214,N_19167,N_18013);
or UO_2215 (O_2215,N_19087,N_19278);
nor UO_2216 (O_2216,N_18991,N_19207);
or UO_2217 (O_2217,N_19034,N_18397);
nand UO_2218 (O_2218,N_19747,N_19334);
nand UO_2219 (O_2219,N_18168,N_18295);
and UO_2220 (O_2220,N_18310,N_18217);
and UO_2221 (O_2221,N_19907,N_18668);
nor UO_2222 (O_2222,N_19125,N_19366);
and UO_2223 (O_2223,N_19116,N_18490);
nand UO_2224 (O_2224,N_18771,N_19701);
and UO_2225 (O_2225,N_18778,N_18237);
or UO_2226 (O_2226,N_18716,N_18870);
nand UO_2227 (O_2227,N_19193,N_19959);
nor UO_2228 (O_2228,N_19144,N_19045);
nand UO_2229 (O_2229,N_19409,N_18963);
xnor UO_2230 (O_2230,N_18297,N_18617);
and UO_2231 (O_2231,N_19735,N_18223);
xor UO_2232 (O_2232,N_19364,N_18729);
and UO_2233 (O_2233,N_19100,N_19299);
and UO_2234 (O_2234,N_18121,N_18644);
and UO_2235 (O_2235,N_19918,N_19783);
or UO_2236 (O_2236,N_19079,N_19716);
and UO_2237 (O_2237,N_19552,N_19548);
nor UO_2238 (O_2238,N_19606,N_18234);
nand UO_2239 (O_2239,N_18338,N_19408);
and UO_2240 (O_2240,N_19320,N_19991);
and UO_2241 (O_2241,N_18943,N_18534);
xor UO_2242 (O_2242,N_19142,N_19699);
xor UO_2243 (O_2243,N_18388,N_18264);
or UO_2244 (O_2244,N_19258,N_19829);
nor UO_2245 (O_2245,N_19007,N_18735);
nor UO_2246 (O_2246,N_18129,N_19044);
or UO_2247 (O_2247,N_19398,N_19140);
and UO_2248 (O_2248,N_19812,N_18610);
nor UO_2249 (O_2249,N_19451,N_19322);
nand UO_2250 (O_2250,N_18763,N_18908);
or UO_2251 (O_2251,N_18881,N_18330);
nand UO_2252 (O_2252,N_18928,N_19426);
or UO_2253 (O_2253,N_19955,N_18441);
nand UO_2254 (O_2254,N_18172,N_18111);
nor UO_2255 (O_2255,N_18068,N_18469);
and UO_2256 (O_2256,N_18368,N_18875);
and UO_2257 (O_2257,N_18791,N_18496);
or UO_2258 (O_2258,N_18918,N_19818);
nor UO_2259 (O_2259,N_19597,N_19342);
and UO_2260 (O_2260,N_18172,N_19181);
nand UO_2261 (O_2261,N_19211,N_18138);
and UO_2262 (O_2262,N_19399,N_19881);
nand UO_2263 (O_2263,N_19129,N_19440);
or UO_2264 (O_2264,N_18681,N_19086);
and UO_2265 (O_2265,N_18691,N_19946);
or UO_2266 (O_2266,N_18154,N_19011);
nor UO_2267 (O_2267,N_18375,N_18948);
and UO_2268 (O_2268,N_18167,N_19556);
or UO_2269 (O_2269,N_19129,N_18499);
or UO_2270 (O_2270,N_18976,N_18423);
or UO_2271 (O_2271,N_18145,N_18615);
or UO_2272 (O_2272,N_19323,N_19400);
or UO_2273 (O_2273,N_18736,N_18972);
or UO_2274 (O_2274,N_19862,N_18308);
or UO_2275 (O_2275,N_19902,N_18210);
and UO_2276 (O_2276,N_18806,N_18479);
and UO_2277 (O_2277,N_18578,N_19637);
or UO_2278 (O_2278,N_18866,N_19499);
nor UO_2279 (O_2279,N_19529,N_18538);
nand UO_2280 (O_2280,N_19073,N_18962);
nand UO_2281 (O_2281,N_19877,N_18401);
nand UO_2282 (O_2282,N_19252,N_18930);
and UO_2283 (O_2283,N_18914,N_19559);
and UO_2284 (O_2284,N_18656,N_18404);
nand UO_2285 (O_2285,N_19832,N_19477);
or UO_2286 (O_2286,N_18977,N_18692);
or UO_2287 (O_2287,N_18087,N_19221);
or UO_2288 (O_2288,N_19396,N_18907);
or UO_2289 (O_2289,N_18852,N_19799);
nor UO_2290 (O_2290,N_19297,N_19671);
nand UO_2291 (O_2291,N_19955,N_18537);
and UO_2292 (O_2292,N_18963,N_19849);
and UO_2293 (O_2293,N_18514,N_19058);
and UO_2294 (O_2294,N_19804,N_18035);
nor UO_2295 (O_2295,N_18585,N_18605);
nand UO_2296 (O_2296,N_18161,N_19778);
and UO_2297 (O_2297,N_18387,N_19572);
or UO_2298 (O_2298,N_18025,N_18527);
xor UO_2299 (O_2299,N_19679,N_19752);
nor UO_2300 (O_2300,N_19242,N_19880);
or UO_2301 (O_2301,N_18013,N_18729);
nand UO_2302 (O_2302,N_19098,N_18609);
nand UO_2303 (O_2303,N_18891,N_18719);
and UO_2304 (O_2304,N_19645,N_18814);
and UO_2305 (O_2305,N_18136,N_19141);
nand UO_2306 (O_2306,N_19412,N_19095);
nor UO_2307 (O_2307,N_19570,N_18298);
or UO_2308 (O_2308,N_19954,N_19887);
and UO_2309 (O_2309,N_18487,N_19971);
xor UO_2310 (O_2310,N_19933,N_18783);
nor UO_2311 (O_2311,N_19519,N_19483);
xnor UO_2312 (O_2312,N_18520,N_19275);
nor UO_2313 (O_2313,N_18130,N_19006);
nand UO_2314 (O_2314,N_18831,N_18883);
nor UO_2315 (O_2315,N_19795,N_19229);
and UO_2316 (O_2316,N_19088,N_19971);
or UO_2317 (O_2317,N_19950,N_19917);
xor UO_2318 (O_2318,N_19748,N_19578);
or UO_2319 (O_2319,N_18263,N_19777);
xnor UO_2320 (O_2320,N_18655,N_19611);
or UO_2321 (O_2321,N_19420,N_18504);
xnor UO_2322 (O_2322,N_19992,N_19348);
nor UO_2323 (O_2323,N_18483,N_19862);
nor UO_2324 (O_2324,N_18872,N_18248);
nor UO_2325 (O_2325,N_18357,N_18701);
xnor UO_2326 (O_2326,N_18704,N_18522);
nor UO_2327 (O_2327,N_19492,N_19624);
or UO_2328 (O_2328,N_19581,N_19874);
or UO_2329 (O_2329,N_18072,N_19473);
xnor UO_2330 (O_2330,N_19952,N_19159);
nand UO_2331 (O_2331,N_18191,N_19598);
xnor UO_2332 (O_2332,N_18807,N_19126);
nand UO_2333 (O_2333,N_19240,N_18752);
nor UO_2334 (O_2334,N_19203,N_18291);
nor UO_2335 (O_2335,N_18832,N_18513);
nand UO_2336 (O_2336,N_18750,N_19253);
nand UO_2337 (O_2337,N_18963,N_18676);
or UO_2338 (O_2338,N_18495,N_18752);
or UO_2339 (O_2339,N_18123,N_18641);
xnor UO_2340 (O_2340,N_19645,N_19094);
nand UO_2341 (O_2341,N_18695,N_19918);
nand UO_2342 (O_2342,N_19518,N_18515);
xnor UO_2343 (O_2343,N_18760,N_18399);
nor UO_2344 (O_2344,N_19373,N_19800);
nor UO_2345 (O_2345,N_19690,N_18243);
or UO_2346 (O_2346,N_18258,N_19240);
nor UO_2347 (O_2347,N_18713,N_19861);
and UO_2348 (O_2348,N_19139,N_19578);
and UO_2349 (O_2349,N_18351,N_18306);
or UO_2350 (O_2350,N_19562,N_19225);
or UO_2351 (O_2351,N_18938,N_18398);
xnor UO_2352 (O_2352,N_19367,N_19978);
nor UO_2353 (O_2353,N_19482,N_18752);
xnor UO_2354 (O_2354,N_19279,N_18167);
nor UO_2355 (O_2355,N_18234,N_19203);
and UO_2356 (O_2356,N_19207,N_18940);
and UO_2357 (O_2357,N_18211,N_19272);
nand UO_2358 (O_2358,N_19472,N_18180);
or UO_2359 (O_2359,N_19911,N_18492);
nor UO_2360 (O_2360,N_18467,N_18815);
xor UO_2361 (O_2361,N_19830,N_19329);
or UO_2362 (O_2362,N_19257,N_19353);
nand UO_2363 (O_2363,N_18427,N_19799);
nand UO_2364 (O_2364,N_19200,N_19602);
or UO_2365 (O_2365,N_19314,N_19957);
or UO_2366 (O_2366,N_18887,N_18107);
nor UO_2367 (O_2367,N_18889,N_18665);
nand UO_2368 (O_2368,N_19510,N_19622);
nor UO_2369 (O_2369,N_18626,N_19697);
or UO_2370 (O_2370,N_18665,N_18323);
nor UO_2371 (O_2371,N_19184,N_19406);
nand UO_2372 (O_2372,N_18894,N_18706);
nand UO_2373 (O_2373,N_18971,N_18962);
or UO_2374 (O_2374,N_19518,N_19443);
nand UO_2375 (O_2375,N_18079,N_18826);
xor UO_2376 (O_2376,N_19034,N_19059);
nand UO_2377 (O_2377,N_19697,N_18473);
and UO_2378 (O_2378,N_19749,N_19993);
nand UO_2379 (O_2379,N_18563,N_18883);
and UO_2380 (O_2380,N_18867,N_19354);
nand UO_2381 (O_2381,N_18906,N_18297);
and UO_2382 (O_2382,N_19090,N_19014);
nor UO_2383 (O_2383,N_18343,N_19335);
nand UO_2384 (O_2384,N_18914,N_19300);
or UO_2385 (O_2385,N_19869,N_18997);
nand UO_2386 (O_2386,N_19037,N_18803);
or UO_2387 (O_2387,N_18586,N_18485);
nand UO_2388 (O_2388,N_18195,N_19166);
or UO_2389 (O_2389,N_19581,N_19082);
or UO_2390 (O_2390,N_19995,N_18165);
and UO_2391 (O_2391,N_19249,N_18504);
and UO_2392 (O_2392,N_19157,N_19857);
nand UO_2393 (O_2393,N_19786,N_18571);
or UO_2394 (O_2394,N_18463,N_18820);
nor UO_2395 (O_2395,N_18426,N_18171);
nand UO_2396 (O_2396,N_18598,N_18364);
and UO_2397 (O_2397,N_19451,N_18666);
nor UO_2398 (O_2398,N_19637,N_19984);
nand UO_2399 (O_2399,N_18945,N_19632);
xor UO_2400 (O_2400,N_19029,N_19682);
or UO_2401 (O_2401,N_19570,N_18056);
nand UO_2402 (O_2402,N_19432,N_18668);
nor UO_2403 (O_2403,N_18022,N_19981);
nor UO_2404 (O_2404,N_19211,N_18226);
nand UO_2405 (O_2405,N_19228,N_18189);
and UO_2406 (O_2406,N_19278,N_18683);
or UO_2407 (O_2407,N_18053,N_18253);
and UO_2408 (O_2408,N_18712,N_18805);
nand UO_2409 (O_2409,N_19053,N_18165);
or UO_2410 (O_2410,N_19127,N_18676);
nand UO_2411 (O_2411,N_18859,N_19612);
nor UO_2412 (O_2412,N_19670,N_19069);
or UO_2413 (O_2413,N_19014,N_18828);
xor UO_2414 (O_2414,N_18934,N_19651);
nor UO_2415 (O_2415,N_18087,N_19262);
and UO_2416 (O_2416,N_19426,N_19142);
or UO_2417 (O_2417,N_19613,N_19186);
xnor UO_2418 (O_2418,N_19379,N_19541);
nor UO_2419 (O_2419,N_18791,N_19515);
or UO_2420 (O_2420,N_19329,N_19800);
and UO_2421 (O_2421,N_18963,N_19662);
nand UO_2422 (O_2422,N_18475,N_19537);
nor UO_2423 (O_2423,N_18078,N_18246);
and UO_2424 (O_2424,N_19653,N_19105);
nor UO_2425 (O_2425,N_19862,N_18194);
nor UO_2426 (O_2426,N_18092,N_19155);
or UO_2427 (O_2427,N_18057,N_19331);
nor UO_2428 (O_2428,N_18166,N_19594);
nand UO_2429 (O_2429,N_18585,N_19948);
nor UO_2430 (O_2430,N_19610,N_19899);
nand UO_2431 (O_2431,N_18673,N_18966);
and UO_2432 (O_2432,N_19277,N_18827);
or UO_2433 (O_2433,N_18753,N_18158);
nor UO_2434 (O_2434,N_18305,N_19557);
xnor UO_2435 (O_2435,N_18828,N_19336);
nor UO_2436 (O_2436,N_19465,N_19545);
nand UO_2437 (O_2437,N_18431,N_18130);
nor UO_2438 (O_2438,N_19315,N_18125);
nor UO_2439 (O_2439,N_18119,N_18589);
nand UO_2440 (O_2440,N_18320,N_19425);
nand UO_2441 (O_2441,N_19489,N_18817);
and UO_2442 (O_2442,N_19893,N_18251);
and UO_2443 (O_2443,N_19161,N_18273);
nor UO_2444 (O_2444,N_19011,N_18538);
and UO_2445 (O_2445,N_18488,N_19399);
nand UO_2446 (O_2446,N_19250,N_18046);
or UO_2447 (O_2447,N_18177,N_18743);
nand UO_2448 (O_2448,N_18355,N_19450);
or UO_2449 (O_2449,N_19578,N_18796);
nor UO_2450 (O_2450,N_19205,N_18540);
and UO_2451 (O_2451,N_18964,N_18897);
and UO_2452 (O_2452,N_18250,N_19349);
nand UO_2453 (O_2453,N_19135,N_18253);
or UO_2454 (O_2454,N_19663,N_18383);
xor UO_2455 (O_2455,N_18742,N_18676);
xor UO_2456 (O_2456,N_19922,N_19167);
and UO_2457 (O_2457,N_19022,N_18428);
or UO_2458 (O_2458,N_18355,N_18541);
nor UO_2459 (O_2459,N_18191,N_18488);
nor UO_2460 (O_2460,N_18492,N_18125);
and UO_2461 (O_2461,N_18506,N_19096);
nand UO_2462 (O_2462,N_19743,N_19811);
nor UO_2463 (O_2463,N_19412,N_18826);
or UO_2464 (O_2464,N_18214,N_19565);
nand UO_2465 (O_2465,N_18231,N_19030);
or UO_2466 (O_2466,N_19123,N_19665);
or UO_2467 (O_2467,N_18016,N_19861);
nor UO_2468 (O_2468,N_18128,N_19707);
or UO_2469 (O_2469,N_18486,N_19683);
or UO_2470 (O_2470,N_19375,N_19820);
nand UO_2471 (O_2471,N_18681,N_19509);
nand UO_2472 (O_2472,N_19500,N_19362);
and UO_2473 (O_2473,N_18709,N_19555);
xor UO_2474 (O_2474,N_19390,N_18530);
nor UO_2475 (O_2475,N_19456,N_19513);
nor UO_2476 (O_2476,N_19707,N_18933);
and UO_2477 (O_2477,N_18356,N_18777);
xor UO_2478 (O_2478,N_18423,N_18087);
nand UO_2479 (O_2479,N_18105,N_19050);
nand UO_2480 (O_2480,N_19615,N_19414);
nor UO_2481 (O_2481,N_19117,N_19547);
and UO_2482 (O_2482,N_19357,N_18240);
nand UO_2483 (O_2483,N_19106,N_18053);
nor UO_2484 (O_2484,N_19046,N_19507);
and UO_2485 (O_2485,N_18596,N_18687);
or UO_2486 (O_2486,N_19351,N_19502);
nor UO_2487 (O_2487,N_19266,N_19185);
nor UO_2488 (O_2488,N_19084,N_18555);
xor UO_2489 (O_2489,N_18309,N_18667);
or UO_2490 (O_2490,N_19835,N_18428);
nand UO_2491 (O_2491,N_18228,N_19006);
nand UO_2492 (O_2492,N_19377,N_18734);
nor UO_2493 (O_2493,N_19928,N_19265);
nor UO_2494 (O_2494,N_19918,N_18716);
nor UO_2495 (O_2495,N_18771,N_19899);
and UO_2496 (O_2496,N_19984,N_18610);
and UO_2497 (O_2497,N_18320,N_18969);
and UO_2498 (O_2498,N_19253,N_19082);
xor UO_2499 (O_2499,N_19456,N_18886);
endmodule