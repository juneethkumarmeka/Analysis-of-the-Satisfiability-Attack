module basic_500_3000_500_5_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_465,In_13);
nor U1 (N_1,In_85,In_422);
or U2 (N_2,In_136,In_378);
nand U3 (N_3,In_10,In_284);
nor U4 (N_4,In_434,In_257);
and U5 (N_5,In_183,In_387);
or U6 (N_6,In_247,In_52);
xnor U7 (N_7,In_189,In_101);
xor U8 (N_8,In_373,In_285);
xnor U9 (N_9,In_231,In_230);
nand U10 (N_10,In_154,In_335);
or U11 (N_11,In_164,In_473);
nor U12 (N_12,In_60,In_433);
nor U13 (N_13,In_315,In_471);
or U14 (N_14,In_296,In_447);
xor U15 (N_15,In_334,In_3);
and U16 (N_16,In_385,In_307);
or U17 (N_17,In_356,In_32);
nand U18 (N_18,In_12,In_144);
nand U19 (N_19,In_347,In_94);
xnor U20 (N_20,In_421,In_71);
nand U21 (N_21,In_475,In_439);
xor U22 (N_22,In_424,In_401);
or U23 (N_23,In_236,In_223);
nor U24 (N_24,In_483,In_117);
nand U25 (N_25,In_30,In_448);
and U26 (N_26,In_429,In_279);
and U27 (N_27,In_330,In_66);
nor U28 (N_28,In_54,In_179);
and U29 (N_29,In_338,In_415);
xor U30 (N_30,In_46,In_109);
nand U31 (N_31,In_391,In_187);
or U32 (N_32,In_93,In_392);
nand U33 (N_33,In_84,In_262);
nor U34 (N_34,In_331,In_360);
nand U35 (N_35,In_72,In_274);
xor U36 (N_36,In_132,In_463);
or U37 (N_37,In_478,In_1);
xnor U38 (N_38,In_177,In_402);
and U39 (N_39,In_290,In_68);
nand U40 (N_40,In_18,In_370);
and U41 (N_41,In_282,In_413);
and U42 (N_42,In_135,In_488);
nor U43 (N_43,In_88,In_355);
xor U44 (N_44,In_299,In_376);
nand U45 (N_45,In_14,In_114);
nand U46 (N_46,In_38,In_65);
and U47 (N_47,In_270,In_408);
nand U48 (N_48,In_192,In_344);
xnor U49 (N_49,In_237,In_70);
and U50 (N_50,In_169,In_363);
and U51 (N_51,In_210,In_375);
or U52 (N_52,In_23,In_322);
and U53 (N_53,In_56,In_388);
nand U54 (N_54,In_219,In_267);
nor U55 (N_55,In_220,In_277);
and U56 (N_56,In_466,In_254);
nand U57 (N_57,In_116,In_368);
xnor U58 (N_58,In_453,In_286);
or U59 (N_59,In_235,In_126);
or U60 (N_60,In_228,In_98);
or U61 (N_61,In_359,In_497);
nor U62 (N_62,In_61,In_321);
or U63 (N_63,In_134,In_437);
nand U64 (N_64,In_140,In_108);
nor U65 (N_65,In_460,In_40);
xnor U66 (N_66,In_310,In_265);
xor U67 (N_67,In_246,In_455);
or U68 (N_68,In_245,In_420);
and U69 (N_69,In_248,In_317);
or U70 (N_70,In_167,In_159);
and U71 (N_71,In_252,In_351);
nor U72 (N_72,In_324,In_59);
or U73 (N_73,In_211,In_441);
and U74 (N_74,In_367,In_481);
xor U75 (N_75,In_339,In_444);
nand U76 (N_76,In_173,In_250);
nand U77 (N_77,In_328,In_125);
xor U78 (N_78,In_291,In_272);
or U79 (N_79,In_452,In_89);
nand U80 (N_80,In_152,In_316);
nand U81 (N_81,In_435,In_107);
xnor U82 (N_82,In_258,In_194);
nor U83 (N_83,In_24,In_498);
nor U84 (N_84,In_329,In_5);
and U85 (N_85,In_303,In_416);
nor U86 (N_86,In_490,In_242);
or U87 (N_87,In_7,In_480);
xnor U88 (N_88,In_142,In_207);
nor U89 (N_89,In_81,In_352);
or U90 (N_90,In_137,In_288);
xor U91 (N_91,In_349,In_346);
and U92 (N_92,In_249,In_449);
nor U93 (N_93,In_423,In_275);
or U94 (N_94,In_42,In_193);
xor U95 (N_95,In_232,In_384);
xnor U96 (N_96,In_305,In_234);
xor U97 (N_97,In_182,In_157);
xor U98 (N_98,In_263,In_199);
and U99 (N_99,In_302,In_204);
nand U100 (N_100,In_15,In_468);
xnor U101 (N_101,In_119,In_106);
and U102 (N_102,In_259,In_405);
xnor U103 (N_103,In_105,In_149);
nor U104 (N_104,In_225,In_464);
xor U105 (N_105,In_362,In_165);
nor U106 (N_106,In_319,In_8);
nor U107 (N_107,In_425,In_342);
nor U108 (N_108,In_426,In_227);
nor U109 (N_109,In_412,In_146);
and U110 (N_110,In_418,In_369);
nor U111 (N_111,In_95,In_97);
nand U112 (N_112,In_19,In_361);
or U113 (N_113,In_160,In_158);
xor U114 (N_114,In_340,In_382);
xnor U115 (N_115,In_47,In_29);
xor U116 (N_116,In_394,In_364);
nand U117 (N_117,In_264,In_371);
or U118 (N_118,In_80,In_256);
nand U119 (N_119,In_380,In_278);
nor U120 (N_120,In_176,In_241);
nand U121 (N_121,In_196,In_202);
nand U122 (N_122,In_233,In_399);
xor U123 (N_123,In_240,In_57);
xnor U124 (N_124,In_404,In_104);
xnor U125 (N_125,In_37,In_477);
nand U126 (N_126,In_406,In_11);
nand U127 (N_127,In_386,In_201);
nand U128 (N_128,In_120,In_92);
nand U129 (N_129,In_485,In_431);
nor U130 (N_130,In_209,In_34);
xnor U131 (N_131,In_96,In_69);
and U132 (N_132,In_45,In_489);
xnor U133 (N_133,In_295,In_381);
or U134 (N_134,In_49,In_161);
or U135 (N_135,In_205,In_450);
xnor U136 (N_136,In_287,In_398);
and U137 (N_137,In_461,In_343);
xor U138 (N_138,In_221,In_229);
nand U139 (N_139,In_99,In_311);
or U140 (N_140,In_292,In_493);
nor U141 (N_141,In_320,In_358);
or U142 (N_142,In_175,In_58);
nand U143 (N_143,In_472,In_162);
nor U144 (N_144,In_396,In_467);
and U145 (N_145,In_130,In_4);
nor U146 (N_146,In_300,In_442);
and U147 (N_147,In_20,In_314);
nand U148 (N_148,In_39,In_222);
xnor U149 (N_149,In_112,In_26);
xnor U150 (N_150,In_118,In_186);
nor U151 (N_151,In_28,In_337);
xor U152 (N_152,In_353,In_393);
xnor U153 (N_153,In_326,In_341);
or U154 (N_154,In_150,In_403);
nand U155 (N_155,In_494,In_180);
or U156 (N_156,In_390,In_21);
xnor U157 (N_157,In_178,In_147);
and U158 (N_158,In_276,In_327);
xor U159 (N_159,In_430,In_16);
and U160 (N_160,In_128,In_499);
xnor U161 (N_161,In_332,In_436);
nor U162 (N_162,In_87,In_172);
and U163 (N_163,In_255,In_377);
xnor U164 (N_164,In_366,In_103);
nand U165 (N_165,In_27,In_357);
xnor U166 (N_166,In_44,In_309);
and U167 (N_167,In_197,In_151);
or U168 (N_168,In_409,In_43);
nor U169 (N_169,In_451,In_83);
or U170 (N_170,In_289,In_123);
and U171 (N_171,In_9,In_389);
nor U172 (N_172,In_208,In_491);
and U173 (N_173,In_200,In_62);
nor U174 (N_174,In_244,In_170);
xnor U175 (N_175,In_458,In_438);
xnor U176 (N_176,In_411,In_479);
and U177 (N_177,In_428,In_261);
nor U178 (N_178,In_31,In_462);
and U179 (N_179,In_239,In_459);
nor U180 (N_180,In_446,In_226);
nor U181 (N_181,In_171,In_496);
xnor U182 (N_182,In_102,In_163);
nor U183 (N_183,In_407,In_454);
xnor U184 (N_184,In_218,In_298);
nand U185 (N_185,In_492,In_139);
nand U186 (N_186,In_206,In_443);
nand U187 (N_187,In_111,In_195);
xnor U188 (N_188,In_414,In_203);
and U189 (N_189,In_74,In_133);
or U190 (N_190,In_50,In_145);
nor U191 (N_191,In_383,In_484);
or U192 (N_192,In_121,In_432);
nand U193 (N_193,In_2,In_457);
nand U194 (N_194,In_91,In_79);
nor U195 (N_195,In_323,In_336);
and U196 (N_196,In_6,In_86);
xor U197 (N_197,In_36,In_417);
and U198 (N_198,In_372,In_184);
nand U199 (N_199,In_419,In_410);
and U200 (N_200,In_400,In_76);
or U201 (N_201,In_476,In_138);
xor U202 (N_202,In_395,In_188);
nor U203 (N_203,In_260,In_122);
and U204 (N_204,In_191,In_440);
xnor U205 (N_205,In_214,In_190);
xnor U206 (N_206,In_141,In_64);
nand U207 (N_207,In_33,In_113);
nand U208 (N_208,In_354,In_63);
nand U209 (N_209,In_75,In_156);
and U210 (N_210,In_212,In_90);
or U211 (N_211,In_168,In_41);
nor U212 (N_212,In_280,In_127);
xnor U213 (N_213,In_487,In_313);
xor U214 (N_214,In_397,In_374);
and U215 (N_215,In_469,In_213);
and U216 (N_216,In_294,In_100);
nor U217 (N_217,In_181,In_297);
nor U218 (N_218,In_55,In_148);
or U219 (N_219,In_253,In_115);
and U220 (N_220,In_22,In_0);
and U221 (N_221,In_243,In_486);
or U222 (N_222,In_17,In_268);
xnor U223 (N_223,In_379,In_308);
and U224 (N_224,In_266,In_129);
xor U225 (N_225,In_131,In_174);
nand U226 (N_226,In_474,In_53);
and U227 (N_227,In_124,In_217);
and U228 (N_228,In_350,In_185);
and U229 (N_229,In_318,In_304);
and U230 (N_230,In_216,In_283);
or U231 (N_231,In_482,In_281);
xnor U232 (N_232,In_445,In_166);
nand U233 (N_233,In_251,In_110);
nor U234 (N_234,In_238,In_273);
or U235 (N_235,In_365,In_215);
or U236 (N_236,In_224,In_77);
or U237 (N_237,In_306,In_78);
xnor U238 (N_238,In_198,In_73);
nand U239 (N_239,In_271,In_67);
and U240 (N_240,In_333,In_82);
xor U241 (N_241,In_293,In_25);
nand U242 (N_242,In_427,In_325);
nor U243 (N_243,In_48,In_153);
and U244 (N_244,In_35,In_470);
and U245 (N_245,In_345,In_456);
or U246 (N_246,In_269,In_348);
and U247 (N_247,In_155,In_143);
nand U248 (N_248,In_495,In_312);
nand U249 (N_249,In_301,In_51);
and U250 (N_250,In_313,In_123);
or U251 (N_251,In_449,In_93);
and U252 (N_252,In_107,In_43);
and U253 (N_253,In_188,In_310);
and U254 (N_254,In_280,In_480);
nand U255 (N_255,In_247,In_77);
xor U256 (N_256,In_482,In_88);
nand U257 (N_257,In_247,In_91);
and U258 (N_258,In_137,In_221);
or U259 (N_259,In_226,In_353);
or U260 (N_260,In_322,In_329);
nand U261 (N_261,In_187,In_23);
nand U262 (N_262,In_304,In_475);
and U263 (N_263,In_452,In_19);
and U264 (N_264,In_267,In_304);
and U265 (N_265,In_444,In_56);
and U266 (N_266,In_391,In_417);
xnor U267 (N_267,In_174,In_13);
or U268 (N_268,In_488,In_383);
and U269 (N_269,In_492,In_101);
or U270 (N_270,In_133,In_212);
nand U271 (N_271,In_19,In_48);
nor U272 (N_272,In_88,In_31);
xor U273 (N_273,In_96,In_468);
and U274 (N_274,In_127,In_453);
nor U275 (N_275,In_185,In_356);
nand U276 (N_276,In_495,In_481);
nand U277 (N_277,In_98,In_149);
or U278 (N_278,In_88,In_463);
xnor U279 (N_279,In_182,In_23);
and U280 (N_280,In_361,In_399);
nor U281 (N_281,In_26,In_322);
xnor U282 (N_282,In_23,In_488);
or U283 (N_283,In_113,In_110);
nor U284 (N_284,In_373,In_303);
xor U285 (N_285,In_111,In_434);
xor U286 (N_286,In_56,In_121);
and U287 (N_287,In_74,In_285);
or U288 (N_288,In_406,In_324);
xor U289 (N_289,In_456,In_498);
nand U290 (N_290,In_140,In_204);
xnor U291 (N_291,In_477,In_53);
nor U292 (N_292,In_361,In_358);
and U293 (N_293,In_245,In_352);
nor U294 (N_294,In_457,In_240);
and U295 (N_295,In_375,In_331);
nor U296 (N_296,In_415,In_96);
nand U297 (N_297,In_125,In_263);
or U298 (N_298,In_112,In_392);
or U299 (N_299,In_23,In_84);
xnor U300 (N_300,In_164,In_327);
nand U301 (N_301,In_339,In_56);
or U302 (N_302,In_375,In_288);
nand U303 (N_303,In_352,In_170);
or U304 (N_304,In_233,In_104);
or U305 (N_305,In_331,In_299);
or U306 (N_306,In_23,In_492);
nand U307 (N_307,In_139,In_194);
nand U308 (N_308,In_54,In_293);
and U309 (N_309,In_439,In_418);
nor U310 (N_310,In_123,In_199);
xnor U311 (N_311,In_275,In_403);
or U312 (N_312,In_382,In_330);
nor U313 (N_313,In_141,In_123);
or U314 (N_314,In_241,In_129);
and U315 (N_315,In_264,In_86);
nor U316 (N_316,In_85,In_425);
or U317 (N_317,In_278,In_484);
and U318 (N_318,In_363,In_100);
nand U319 (N_319,In_380,In_430);
and U320 (N_320,In_492,In_116);
xor U321 (N_321,In_471,In_449);
xnor U322 (N_322,In_341,In_71);
or U323 (N_323,In_363,In_10);
nor U324 (N_324,In_234,In_245);
or U325 (N_325,In_76,In_414);
nand U326 (N_326,In_459,In_404);
nor U327 (N_327,In_383,In_252);
nor U328 (N_328,In_461,In_437);
or U329 (N_329,In_112,In_480);
nor U330 (N_330,In_331,In_392);
xor U331 (N_331,In_345,In_440);
and U332 (N_332,In_15,In_206);
and U333 (N_333,In_7,In_125);
and U334 (N_334,In_186,In_47);
xnor U335 (N_335,In_336,In_41);
and U336 (N_336,In_348,In_362);
nand U337 (N_337,In_221,In_389);
and U338 (N_338,In_66,In_160);
or U339 (N_339,In_410,In_33);
nor U340 (N_340,In_438,In_122);
and U341 (N_341,In_472,In_155);
nand U342 (N_342,In_247,In_265);
nand U343 (N_343,In_249,In_362);
xor U344 (N_344,In_411,In_234);
nand U345 (N_345,In_414,In_390);
or U346 (N_346,In_351,In_157);
or U347 (N_347,In_53,In_457);
xnor U348 (N_348,In_452,In_440);
nor U349 (N_349,In_119,In_70);
xor U350 (N_350,In_230,In_105);
and U351 (N_351,In_197,In_81);
or U352 (N_352,In_344,In_301);
nand U353 (N_353,In_236,In_267);
or U354 (N_354,In_229,In_100);
xnor U355 (N_355,In_274,In_149);
xnor U356 (N_356,In_395,In_335);
or U357 (N_357,In_470,In_29);
xnor U358 (N_358,In_486,In_202);
and U359 (N_359,In_188,In_372);
nand U360 (N_360,In_222,In_18);
xor U361 (N_361,In_416,In_118);
xor U362 (N_362,In_316,In_408);
xor U363 (N_363,In_346,In_399);
or U364 (N_364,In_2,In_365);
nor U365 (N_365,In_494,In_111);
nor U366 (N_366,In_307,In_82);
xnor U367 (N_367,In_27,In_284);
and U368 (N_368,In_326,In_389);
or U369 (N_369,In_351,In_143);
and U370 (N_370,In_459,In_75);
or U371 (N_371,In_326,In_89);
or U372 (N_372,In_369,In_173);
and U373 (N_373,In_143,In_320);
xnor U374 (N_374,In_74,In_219);
xor U375 (N_375,In_54,In_172);
nor U376 (N_376,In_484,In_343);
nor U377 (N_377,In_112,In_466);
or U378 (N_378,In_112,In_115);
nor U379 (N_379,In_94,In_375);
xnor U380 (N_380,In_140,In_132);
and U381 (N_381,In_136,In_325);
xnor U382 (N_382,In_365,In_433);
nand U383 (N_383,In_68,In_59);
xnor U384 (N_384,In_139,In_323);
and U385 (N_385,In_110,In_114);
nor U386 (N_386,In_243,In_4);
and U387 (N_387,In_66,In_294);
xor U388 (N_388,In_47,In_383);
xor U389 (N_389,In_23,In_276);
or U390 (N_390,In_239,In_363);
or U391 (N_391,In_138,In_258);
nand U392 (N_392,In_317,In_431);
xnor U393 (N_393,In_374,In_341);
nor U394 (N_394,In_38,In_141);
or U395 (N_395,In_480,In_476);
nand U396 (N_396,In_288,In_1);
xor U397 (N_397,In_267,In_10);
or U398 (N_398,In_105,In_428);
or U399 (N_399,In_475,In_332);
xnor U400 (N_400,In_96,In_478);
xnor U401 (N_401,In_19,In_40);
nor U402 (N_402,In_34,In_356);
or U403 (N_403,In_452,In_198);
nand U404 (N_404,In_427,In_457);
xor U405 (N_405,In_68,In_289);
and U406 (N_406,In_402,In_277);
nand U407 (N_407,In_443,In_191);
or U408 (N_408,In_28,In_178);
and U409 (N_409,In_499,In_248);
nand U410 (N_410,In_21,In_167);
or U411 (N_411,In_155,In_174);
nand U412 (N_412,In_142,In_382);
and U413 (N_413,In_245,In_178);
nor U414 (N_414,In_164,In_237);
nand U415 (N_415,In_166,In_318);
or U416 (N_416,In_183,In_19);
and U417 (N_417,In_326,In_445);
nor U418 (N_418,In_9,In_106);
or U419 (N_419,In_410,In_359);
and U420 (N_420,In_406,In_346);
nor U421 (N_421,In_247,In_246);
xnor U422 (N_422,In_337,In_125);
and U423 (N_423,In_358,In_388);
nor U424 (N_424,In_48,In_357);
xnor U425 (N_425,In_480,In_262);
or U426 (N_426,In_473,In_46);
nor U427 (N_427,In_152,In_371);
xnor U428 (N_428,In_294,In_307);
nand U429 (N_429,In_460,In_248);
nand U430 (N_430,In_156,In_297);
nor U431 (N_431,In_441,In_41);
and U432 (N_432,In_199,In_211);
and U433 (N_433,In_170,In_149);
nor U434 (N_434,In_86,In_383);
nor U435 (N_435,In_22,In_230);
nor U436 (N_436,In_157,In_150);
xor U437 (N_437,In_70,In_445);
and U438 (N_438,In_230,In_399);
and U439 (N_439,In_119,In_309);
nor U440 (N_440,In_140,In_329);
or U441 (N_441,In_441,In_11);
or U442 (N_442,In_290,In_490);
nand U443 (N_443,In_164,In_491);
nor U444 (N_444,In_114,In_155);
xnor U445 (N_445,In_32,In_144);
or U446 (N_446,In_9,In_160);
nand U447 (N_447,In_253,In_112);
nand U448 (N_448,In_135,In_363);
and U449 (N_449,In_0,In_381);
or U450 (N_450,In_23,In_280);
or U451 (N_451,In_151,In_58);
nor U452 (N_452,In_178,In_229);
xnor U453 (N_453,In_20,In_48);
nor U454 (N_454,In_397,In_49);
and U455 (N_455,In_352,In_87);
or U456 (N_456,In_336,In_8);
xnor U457 (N_457,In_299,In_404);
nor U458 (N_458,In_422,In_358);
nor U459 (N_459,In_185,In_469);
and U460 (N_460,In_37,In_465);
nor U461 (N_461,In_236,In_245);
and U462 (N_462,In_424,In_337);
nor U463 (N_463,In_274,In_231);
nor U464 (N_464,In_459,In_82);
nand U465 (N_465,In_248,In_44);
nor U466 (N_466,In_98,In_18);
xnor U467 (N_467,In_27,In_294);
or U468 (N_468,In_110,In_457);
and U469 (N_469,In_142,In_117);
xor U470 (N_470,In_299,In_388);
nand U471 (N_471,In_155,In_411);
and U472 (N_472,In_355,In_63);
nor U473 (N_473,In_268,In_378);
xnor U474 (N_474,In_498,In_430);
nand U475 (N_475,In_407,In_335);
xor U476 (N_476,In_260,In_341);
nand U477 (N_477,In_273,In_35);
xnor U478 (N_478,In_42,In_135);
and U479 (N_479,In_286,In_278);
xnor U480 (N_480,In_489,In_37);
nand U481 (N_481,In_319,In_103);
xnor U482 (N_482,In_332,In_117);
nor U483 (N_483,In_283,In_403);
nor U484 (N_484,In_495,In_232);
and U485 (N_485,In_292,In_441);
or U486 (N_486,In_426,In_378);
or U487 (N_487,In_149,In_50);
nor U488 (N_488,In_152,In_3);
nor U489 (N_489,In_397,In_473);
and U490 (N_490,In_354,In_124);
and U491 (N_491,In_55,In_294);
nand U492 (N_492,In_10,In_13);
nand U493 (N_493,In_82,In_178);
nand U494 (N_494,In_119,In_98);
nand U495 (N_495,In_316,In_302);
or U496 (N_496,In_95,In_448);
nand U497 (N_497,In_43,In_452);
nor U498 (N_498,In_278,In_361);
nor U499 (N_499,In_330,In_348);
or U500 (N_500,In_472,In_329);
nand U501 (N_501,In_395,In_336);
nand U502 (N_502,In_264,In_56);
xor U503 (N_503,In_48,In_41);
xor U504 (N_504,In_94,In_302);
or U505 (N_505,In_470,In_484);
or U506 (N_506,In_335,In_224);
xor U507 (N_507,In_23,In_142);
nand U508 (N_508,In_378,In_302);
xnor U509 (N_509,In_149,In_479);
xor U510 (N_510,In_97,In_279);
nand U511 (N_511,In_111,In_64);
nand U512 (N_512,In_455,In_413);
nor U513 (N_513,In_40,In_395);
and U514 (N_514,In_256,In_442);
nand U515 (N_515,In_337,In_182);
and U516 (N_516,In_64,In_349);
nand U517 (N_517,In_211,In_401);
xnor U518 (N_518,In_111,In_132);
xor U519 (N_519,In_176,In_328);
and U520 (N_520,In_316,In_20);
nor U521 (N_521,In_100,In_122);
nor U522 (N_522,In_84,In_390);
xor U523 (N_523,In_166,In_176);
or U524 (N_524,In_271,In_335);
xnor U525 (N_525,In_76,In_84);
and U526 (N_526,In_253,In_315);
nand U527 (N_527,In_218,In_340);
xor U528 (N_528,In_459,In_188);
nor U529 (N_529,In_203,In_347);
xor U530 (N_530,In_228,In_420);
nor U531 (N_531,In_109,In_14);
or U532 (N_532,In_447,In_431);
nand U533 (N_533,In_453,In_380);
and U534 (N_534,In_267,In_153);
and U535 (N_535,In_162,In_45);
xor U536 (N_536,In_329,In_93);
and U537 (N_537,In_156,In_428);
nor U538 (N_538,In_9,In_289);
xor U539 (N_539,In_308,In_361);
nand U540 (N_540,In_134,In_171);
nand U541 (N_541,In_80,In_108);
or U542 (N_542,In_436,In_475);
and U543 (N_543,In_347,In_492);
nand U544 (N_544,In_164,In_411);
and U545 (N_545,In_4,In_431);
nand U546 (N_546,In_150,In_53);
or U547 (N_547,In_336,In_134);
nand U548 (N_548,In_427,In_258);
xnor U549 (N_549,In_482,In_278);
or U550 (N_550,In_302,In_411);
xor U551 (N_551,In_349,In_253);
nor U552 (N_552,In_296,In_430);
and U553 (N_553,In_444,In_95);
nand U554 (N_554,In_243,In_347);
or U555 (N_555,In_458,In_97);
xnor U556 (N_556,In_236,In_292);
and U557 (N_557,In_34,In_433);
and U558 (N_558,In_443,In_12);
and U559 (N_559,In_58,In_7);
and U560 (N_560,In_287,In_103);
or U561 (N_561,In_290,In_197);
nor U562 (N_562,In_451,In_261);
xnor U563 (N_563,In_74,In_58);
nand U564 (N_564,In_238,In_39);
and U565 (N_565,In_227,In_216);
and U566 (N_566,In_281,In_431);
nor U567 (N_567,In_396,In_26);
nand U568 (N_568,In_247,In_140);
nand U569 (N_569,In_333,In_182);
nor U570 (N_570,In_461,In_389);
and U571 (N_571,In_244,In_209);
nand U572 (N_572,In_126,In_260);
nand U573 (N_573,In_274,In_205);
xor U574 (N_574,In_55,In_135);
nor U575 (N_575,In_310,In_288);
or U576 (N_576,In_222,In_372);
nor U577 (N_577,In_186,In_408);
and U578 (N_578,In_159,In_314);
nor U579 (N_579,In_64,In_332);
nor U580 (N_580,In_482,In_271);
nand U581 (N_581,In_470,In_174);
and U582 (N_582,In_46,In_215);
and U583 (N_583,In_215,In_225);
nor U584 (N_584,In_319,In_412);
or U585 (N_585,In_492,In_230);
nand U586 (N_586,In_305,In_393);
or U587 (N_587,In_445,In_478);
nand U588 (N_588,In_158,In_299);
nand U589 (N_589,In_104,In_333);
xnor U590 (N_590,In_93,In_403);
nand U591 (N_591,In_416,In_23);
nor U592 (N_592,In_417,In_179);
xor U593 (N_593,In_258,In_197);
and U594 (N_594,In_101,In_384);
nand U595 (N_595,In_25,In_36);
and U596 (N_596,In_422,In_378);
nor U597 (N_597,In_77,In_29);
nand U598 (N_598,In_426,In_422);
xnor U599 (N_599,In_409,In_89);
nor U600 (N_600,N_253,N_452);
and U601 (N_601,N_94,N_507);
and U602 (N_602,N_30,N_86);
or U603 (N_603,N_549,N_584);
or U604 (N_604,N_392,N_235);
or U605 (N_605,N_117,N_27);
nor U606 (N_606,N_98,N_487);
or U607 (N_607,N_156,N_343);
xnor U608 (N_608,N_573,N_334);
or U609 (N_609,N_345,N_543);
xnor U610 (N_610,N_361,N_150);
or U611 (N_611,N_404,N_365);
xor U612 (N_612,N_537,N_285);
nand U613 (N_613,N_476,N_562);
or U614 (N_614,N_576,N_242);
or U615 (N_615,N_388,N_384);
xor U616 (N_616,N_493,N_508);
xnor U617 (N_617,N_199,N_319);
and U618 (N_618,N_478,N_520);
and U619 (N_619,N_44,N_233);
and U620 (N_620,N_312,N_48);
nand U621 (N_621,N_479,N_275);
nor U622 (N_622,N_77,N_100);
or U623 (N_623,N_169,N_350);
xor U624 (N_624,N_225,N_95);
and U625 (N_625,N_542,N_454);
xnor U626 (N_626,N_243,N_380);
nand U627 (N_627,N_0,N_214);
xor U628 (N_628,N_567,N_24);
or U629 (N_629,N_208,N_218);
or U630 (N_630,N_455,N_265);
and U631 (N_631,N_333,N_582);
nor U632 (N_632,N_194,N_284);
or U633 (N_633,N_359,N_278);
nor U634 (N_634,N_468,N_399);
or U635 (N_635,N_126,N_205);
or U636 (N_636,N_534,N_357);
xnor U637 (N_637,N_344,N_2);
nor U638 (N_638,N_230,N_29);
nor U639 (N_639,N_481,N_73);
nand U640 (N_640,N_129,N_165);
or U641 (N_641,N_32,N_207);
nor U642 (N_642,N_456,N_341);
nand U643 (N_643,N_535,N_189);
and U644 (N_644,N_459,N_463);
xor U645 (N_645,N_66,N_244);
nor U646 (N_646,N_441,N_439);
xnor U647 (N_647,N_526,N_367);
and U648 (N_648,N_458,N_234);
and U649 (N_649,N_41,N_35);
nand U650 (N_650,N_81,N_197);
xor U651 (N_651,N_201,N_179);
nor U652 (N_652,N_354,N_310);
nor U653 (N_653,N_587,N_503);
xor U654 (N_654,N_346,N_482);
nor U655 (N_655,N_352,N_162);
xor U656 (N_656,N_449,N_295);
nand U657 (N_657,N_202,N_203);
and U658 (N_658,N_200,N_134);
or U659 (N_659,N_375,N_421);
or U660 (N_660,N_288,N_530);
or U661 (N_661,N_475,N_241);
nand U662 (N_662,N_324,N_464);
or U663 (N_663,N_236,N_595);
or U664 (N_664,N_377,N_17);
xnor U665 (N_665,N_239,N_405);
nor U666 (N_666,N_364,N_93);
nor U667 (N_667,N_237,N_510);
or U668 (N_668,N_566,N_320);
xnor U669 (N_669,N_213,N_220);
nand U670 (N_670,N_215,N_61);
xnor U671 (N_671,N_308,N_4);
or U672 (N_672,N_461,N_67);
nor U673 (N_673,N_137,N_436);
nand U674 (N_674,N_206,N_188);
or U675 (N_675,N_484,N_120);
xor U676 (N_676,N_3,N_490);
and U677 (N_677,N_163,N_415);
nand U678 (N_678,N_321,N_460);
or U679 (N_679,N_114,N_280);
nor U680 (N_680,N_374,N_25);
or U681 (N_681,N_57,N_523);
xnor U682 (N_682,N_572,N_416);
nand U683 (N_683,N_512,N_267);
or U684 (N_684,N_276,N_140);
xor U685 (N_685,N_531,N_467);
or U686 (N_686,N_286,N_72);
and U687 (N_687,N_574,N_528);
xnor U688 (N_688,N_492,N_389);
and U689 (N_689,N_58,N_433);
or U690 (N_690,N_485,N_80);
nor U691 (N_691,N_131,N_107);
nor U692 (N_692,N_103,N_581);
nor U693 (N_693,N_578,N_159);
or U694 (N_694,N_119,N_178);
nor U695 (N_695,N_160,N_408);
and U696 (N_696,N_465,N_403);
nor U697 (N_697,N_297,N_106);
nand U698 (N_698,N_412,N_154);
nand U699 (N_699,N_173,N_586);
xnor U700 (N_700,N_296,N_217);
or U701 (N_701,N_125,N_486);
nor U702 (N_702,N_446,N_168);
and U703 (N_703,N_51,N_184);
xnor U704 (N_704,N_229,N_84);
nor U705 (N_705,N_246,N_74);
xor U706 (N_706,N_317,N_351);
or U707 (N_707,N_39,N_26);
xor U708 (N_708,N_315,N_327);
and U709 (N_709,N_87,N_366);
and U710 (N_710,N_6,N_282);
and U711 (N_711,N_360,N_538);
or U712 (N_712,N_391,N_142);
xnor U713 (N_713,N_264,N_124);
nor U714 (N_714,N_298,N_394);
and U715 (N_715,N_473,N_385);
and U716 (N_716,N_151,N_55);
nor U717 (N_717,N_420,N_422);
nor U718 (N_718,N_429,N_301);
nor U719 (N_719,N_330,N_291);
or U720 (N_720,N_338,N_325);
or U721 (N_721,N_593,N_382);
xor U722 (N_722,N_248,N_60);
xor U723 (N_723,N_33,N_191);
nand U724 (N_724,N_316,N_506);
and U725 (N_725,N_299,N_251);
or U726 (N_726,N_488,N_349);
nand U727 (N_727,N_190,N_513);
or U728 (N_728,N_470,N_555);
and U729 (N_729,N_548,N_147);
nand U730 (N_730,N_294,N_303);
or U731 (N_731,N_209,N_430);
nor U732 (N_732,N_469,N_347);
nor U733 (N_733,N_270,N_193);
or U734 (N_734,N_505,N_522);
xnor U735 (N_735,N_21,N_115);
nand U736 (N_736,N_116,N_560);
xnor U737 (N_737,N_172,N_434);
or U738 (N_738,N_28,N_544);
xnor U739 (N_739,N_509,N_34);
or U740 (N_740,N_552,N_588);
xor U741 (N_741,N_182,N_292);
or U742 (N_742,N_450,N_356);
and U743 (N_743,N_328,N_226);
nor U744 (N_744,N_307,N_49);
nor U745 (N_745,N_164,N_414);
nand U746 (N_746,N_501,N_227);
and U747 (N_747,N_397,N_348);
xor U748 (N_748,N_211,N_323);
or U749 (N_749,N_79,N_254);
nand U750 (N_750,N_198,N_171);
nor U751 (N_751,N_504,N_157);
nand U752 (N_752,N_259,N_314);
xnor U753 (N_753,N_546,N_551);
nand U754 (N_754,N_266,N_570);
nand U755 (N_755,N_144,N_186);
and U756 (N_756,N_402,N_263);
xnor U757 (N_757,N_466,N_440);
nand U758 (N_758,N_91,N_594);
or U759 (N_759,N_149,N_500);
and U760 (N_760,N_68,N_136);
and U761 (N_761,N_498,N_395);
and U762 (N_762,N_104,N_224);
or U763 (N_763,N_425,N_532);
nor U764 (N_764,N_138,N_212);
nor U765 (N_765,N_54,N_483);
nor U766 (N_766,N_272,N_499);
nor U767 (N_767,N_599,N_502);
nor U768 (N_768,N_378,N_53);
xor U769 (N_769,N_45,N_5);
and U770 (N_770,N_180,N_568);
nand U771 (N_771,N_269,N_10);
nor U772 (N_772,N_477,N_20);
nor U773 (N_773,N_101,N_557);
or U774 (N_774,N_153,N_155);
xor U775 (N_775,N_38,N_219);
nand U776 (N_776,N_368,N_148);
or U777 (N_777,N_290,N_221);
xnor U778 (N_778,N_443,N_70);
nand U779 (N_779,N_491,N_556);
and U780 (N_780,N_398,N_424);
or U781 (N_781,N_279,N_268);
xnor U782 (N_782,N_71,N_515);
nand U783 (N_783,N_418,N_442);
or U784 (N_784,N_335,N_431);
xnor U785 (N_785,N_69,N_255);
nand U786 (N_786,N_139,N_192);
and U787 (N_787,N_92,N_579);
and U788 (N_788,N_447,N_400);
nor U789 (N_789,N_277,N_252);
nand U790 (N_790,N_43,N_222);
xor U791 (N_791,N_65,N_133);
nand U792 (N_792,N_262,N_31);
nand U793 (N_793,N_448,N_362);
xor U794 (N_794,N_260,N_426);
xor U795 (N_795,N_337,N_231);
or U796 (N_796,N_339,N_527);
xnor U797 (N_797,N_540,N_113);
nor U798 (N_798,N_300,N_177);
and U799 (N_799,N_210,N_99);
nand U800 (N_800,N_132,N_363);
nor U801 (N_801,N_118,N_406);
or U802 (N_802,N_519,N_529);
nor U803 (N_803,N_474,N_283);
xnor U804 (N_804,N_161,N_302);
nor U805 (N_805,N_97,N_281);
nor U806 (N_806,N_564,N_386);
and U807 (N_807,N_89,N_112);
xor U808 (N_808,N_240,N_121);
xor U809 (N_809,N_273,N_517);
xor U810 (N_810,N_353,N_575);
nand U811 (N_811,N_417,N_289);
nand U812 (N_812,N_216,N_340);
or U813 (N_813,N_533,N_390);
or U814 (N_814,N_18,N_561);
xor U815 (N_815,N_381,N_511);
or U816 (N_816,N_247,N_471);
and U817 (N_817,N_46,N_590);
xnor U818 (N_818,N_451,N_419);
nand U819 (N_819,N_536,N_596);
or U820 (N_820,N_598,N_40);
xor U821 (N_821,N_583,N_8);
or U822 (N_822,N_409,N_445);
or U823 (N_823,N_83,N_196);
nor U824 (N_824,N_514,N_411);
or U825 (N_825,N_176,N_185);
nor U826 (N_826,N_85,N_571);
or U827 (N_827,N_332,N_12);
nand U828 (N_828,N_245,N_372);
nor U829 (N_829,N_183,N_521);
nand U830 (N_830,N_167,N_379);
xnor U831 (N_831,N_105,N_195);
nor U832 (N_832,N_591,N_545);
nand U833 (N_833,N_274,N_494);
and U834 (N_834,N_370,N_518);
xnor U835 (N_835,N_1,N_96);
and U836 (N_836,N_52,N_64);
and U837 (N_837,N_539,N_497);
xnor U838 (N_838,N_82,N_228);
xnor U839 (N_839,N_293,N_427);
nand U840 (N_840,N_50,N_158);
nand U841 (N_841,N_62,N_313);
nor U842 (N_842,N_187,N_558);
and U843 (N_843,N_271,N_597);
nand U844 (N_844,N_524,N_232);
nand U845 (N_845,N_146,N_435);
and U846 (N_846,N_525,N_453);
nand U847 (N_847,N_496,N_145);
nor U848 (N_848,N_437,N_135);
and U849 (N_849,N_580,N_309);
nand U850 (N_850,N_428,N_410);
nand U851 (N_851,N_128,N_108);
or U852 (N_852,N_553,N_122);
and U853 (N_853,N_13,N_250);
or U854 (N_854,N_109,N_371);
and U855 (N_855,N_123,N_170);
nor U856 (N_856,N_401,N_305);
nor U857 (N_857,N_369,N_329);
and U858 (N_858,N_287,N_589);
and U859 (N_859,N_9,N_102);
and U860 (N_860,N_238,N_110);
nor U861 (N_861,N_376,N_585);
and U862 (N_862,N_326,N_516);
and U863 (N_863,N_358,N_355);
xor U864 (N_864,N_489,N_423);
nand U865 (N_865,N_127,N_322);
nand U866 (N_866,N_37,N_342);
and U867 (N_867,N_257,N_56);
or U868 (N_868,N_541,N_336);
nor U869 (N_869,N_16,N_258);
xnor U870 (N_870,N_75,N_7);
nor U871 (N_871,N_174,N_76);
and U872 (N_872,N_166,N_256);
or U873 (N_873,N_495,N_331);
and U874 (N_874,N_111,N_181);
or U875 (N_875,N_152,N_90);
or U876 (N_876,N_432,N_23);
and U877 (N_877,N_318,N_472);
xnor U878 (N_878,N_63,N_373);
nor U879 (N_879,N_143,N_462);
xnor U880 (N_880,N_393,N_11);
xnor U881 (N_881,N_554,N_444);
and U882 (N_882,N_223,N_457);
nor U883 (N_883,N_175,N_559);
or U884 (N_884,N_59,N_577);
nor U885 (N_885,N_383,N_387);
nor U886 (N_886,N_311,N_130);
nand U887 (N_887,N_141,N_407);
nor U888 (N_888,N_569,N_592);
xnor U889 (N_889,N_88,N_563);
nand U890 (N_890,N_14,N_306);
nor U891 (N_891,N_22,N_47);
xor U892 (N_892,N_413,N_78);
and U893 (N_893,N_438,N_565);
xnor U894 (N_894,N_547,N_42);
or U895 (N_895,N_396,N_249);
nor U896 (N_896,N_15,N_304);
or U897 (N_897,N_36,N_204);
and U898 (N_898,N_261,N_19);
or U899 (N_899,N_480,N_550);
xnor U900 (N_900,N_410,N_422);
nor U901 (N_901,N_281,N_47);
and U902 (N_902,N_540,N_225);
xor U903 (N_903,N_48,N_183);
nor U904 (N_904,N_203,N_451);
xor U905 (N_905,N_592,N_555);
xor U906 (N_906,N_226,N_178);
and U907 (N_907,N_440,N_176);
xor U908 (N_908,N_590,N_521);
and U909 (N_909,N_276,N_106);
xnor U910 (N_910,N_55,N_457);
nor U911 (N_911,N_394,N_81);
or U912 (N_912,N_581,N_547);
nor U913 (N_913,N_278,N_577);
and U914 (N_914,N_587,N_105);
or U915 (N_915,N_445,N_69);
xor U916 (N_916,N_79,N_534);
and U917 (N_917,N_564,N_531);
nor U918 (N_918,N_156,N_223);
xor U919 (N_919,N_444,N_246);
nor U920 (N_920,N_524,N_151);
xor U921 (N_921,N_79,N_581);
nor U922 (N_922,N_33,N_399);
or U923 (N_923,N_321,N_381);
or U924 (N_924,N_553,N_212);
xor U925 (N_925,N_229,N_565);
or U926 (N_926,N_282,N_416);
nand U927 (N_927,N_362,N_61);
xor U928 (N_928,N_305,N_353);
and U929 (N_929,N_324,N_60);
or U930 (N_930,N_234,N_470);
and U931 (N_931,N_527,N_374);
and U932 (N_932,N_375,N_58);
and U933 (N_933,N_251,N_7);
nor U934 (N_934,N_118,N_324);
xnor U935 (N_935,N_530,N_4);
xor U936 (N_936,N_454,N_569);
xnor U937 (N_937,N_124,N_396);
nor U938 (N_938,N_203,N_395);
xnor U939 (N_939,N_290,N_550);
nor U940 (N_940,N_108,N_414);
nor U941 (N_941,N_315,N_352);
nor U942 (N_942,N_347,N_245);
nand U943 (N_943,N_245,N_577);
xnor U944 (N_944,N_537,N_136);
nor U945 (N_945,N_66,N_405);
or U946 (N_946,N_117,N_468);
and U947 (N_947,N_118,N_232);
and U948 (N_948,N_165,N_218);
or U949 (N_949,N_361,N_463);
nand U950 (N_950,N_373,N_268);
xnor U951 (N_951,N_408,N_574);
nor U952 (N_952,N_223,N_118);
nand U953 (N_953,N_303,N_58);
and U954 (N_954,N_292,N_234);
nor U955 (N_955,N_247,N_23);
nand U956 (N_956,N_543,N_412);
and U957 (N_957,N_454,N_279);
xnor U958 (N_958,N_414,N_26);
xnor U959 (N_959,N_467,N_356);
xnor U960 (N_960,N_489,N_377);
nor U961 (N_961,N_516,N_170);
xor U962 (N_962,N_87,N_456);
and U963 (N_963,N_194,N_376);
xor U964 (N_964,N_360,N_116);
nor U965 (N_965,N_359,N_507);
and U966 (N_966,N_200,N_2);
nor U967 (N_967,N_378,N_242);
nor U968 (N_968,N_376,N_406);
or U969 (N_969,N_300,N_423);
and U970 (N_970,N_359,N_12);
or U971 (N_971,N_548,N_178);
and U972 (N_972,N_81,N_184);
xor U973 (N_973,N_23,N_559);
nor U974 (N_974,N_477,N_422);
nand U975 (N_975,N_401,N_513);
nand U976 (N_976,N_484,N_582);
xnor U977 (N_977,N_443,N_383);
nor U978 (N_978,N_27,N_160);
nor U979 (N_979,N_418,N_120);
xnor U980 (N_980,N_72,N_308);
xor U981 (N_981,N_210,N_260);
xnor U982 (N_982,N_280,N_310);
or U983 (N_983,N_390,N_123);
nor U984 (N_984,N_241,N_366);
and U985 (N_985,N_415,N_211);
nand U986 (N_986,N_62,N_433);
nor U987 (N_987,N_155,N_325);
nand U988 (N_988,N_76,N_527);
or U989 (N_989,N_56,N_311);
xor U990 (N_990,N_445,N_348);
xor U991 (N_991,N_261,N_476);
or U992 (N_992,N_26,N_138);
and U993 (N_993,N_332,N_351);
or U994 (N_994,N_499,N_550);
xnor U995 (N_995,N_419,N_474);
or U996 (N_996,N_57,N_457);
nor U997 (N_997,N_125,N_243);
xor U998 (N_998,N_192,N_100);
and U999 (N_999,N_182,N_184);
nor U1000 (N_1000,N_232,N_448);
and U1001 (N_1001,N_279,N_504);
xor U1002 (N_1002,N_475,N_421);
xor U1003 (N_1003,N_577,N_252);
or U1004 (N_1004,N_36,N_325);
and U1005 (N_1005,N_94,N_326);
and U1006 (N_1006,N_72,N_448);
nand U1007 (N_1007,N_415,N_226);
nand U1008 (N_1008,N_589,N_86);
nor U1009 (N_1009,N_413,N_396);
and U1010 (N_1010,N_236,N_414);
and U1011 (N_1011,N_243,N_104);
or U1012 (N_1012,N_204,N_45);
nor U1013 (N_1013,N_143,N_271);
or U1014 (N_1014,N_583,N_124);
and U1015 (N_1015,N_159,N_404);
nor U1016 (N_1016,N_165,N_159);
nand U1017 (N_1017,N_311,N_529);
and U1018 (N_1018,N_573,N_597);
nand U1019 (N_1019,N_456,N_283);
and U1020 (N_1020,N_162,N_19);
nand U1021 (N_1021,N_251,N_416);
nand U1022 (N_1022,N_296,N_149);
and U1023 (N_1023,N_437,N_274);
or U1024 (N_1024,N_360,N_421);
and U1025 (N_1025,N_511,N_541);
nand U1026 (N_1026,N_166,N_550);
or U1027 (N_1027,N_242,N_210);
or U1028 (N_1028,N_112,N_265);
xnor U1029 (N_1029,N_564,N_67);
nor U1030 (N_1030,N_509,N_317);
and U1031 (N_1031,N_24,N_365);
nand U1032 (N_1032,N_0,N_207);
xor U1033 (N_1033,N_337,N_192);
or U1034 (N_1034,N_158,N_224);
xnor U1035 (N_1035,N_214,N_293);
xor U1036 (N_1036,N_347,N_590);
or U1037 (N_1037,N_439,N_165);
nand U1038 (N_1038,N_142,N_382);
or U1039 (N_1039,N_371,N_224);
nand U1040 (N_1040,N_430,N_269);
nand U1041 (N_1041,N_114,N_137);
nor U1042 (N_1042,N_143,N_540);
nor U1043 (N_1043,N_565,N_543);
and U1044 (N_1044,N_500,N_537);
and U1045 (N_1045,N_216,N_176);
and U1046 (N_1046,N_494,N_92);
nor U1047 (N_1047,N_445,N_541);
nor U1048 (N_1048,N_39,N_190);
or U1049 (N_1049,N_514,N_507);
nor U1050 (N_1050,N_384,N_353);
nand U1051 (N_1051,N_228,N_407);
nand U1052 (N_1052,N_191,N_431);
nand U1053 (N_1053,N_480,N_53);
nor U1054 (N_1054,N_57,N_520);
nand U1055 (N_1055,N_429,N_113);
and U1056 (N_1056,N_349,N_387);
xnor U1057 (N_1057,N_514,N_337);
and U1058 (N_1058,N_37,N_473);
nor U1059 (N_1059,N_582,N_238);
and U1060 (N_1060,N_110,N_555);
and U1061 (N_1061,N_174,N_351);
nand U1062 (N_1062,N_461,N_4);
and U1063 (N_1063,N_37,N_210);
nor U1064 (N_1064,N_562,N_549);
or U1065 (N_1065,N_340,N_439);
nor U1066 (N_1066,N_30,N_450);
and U1067 (N_1067,N_428,N_486);
or U1068 (N_1068,N_48,N_53);
nand U1069 (N_1069,N_99,N_374);
nand U1070 (N_1070,N_154,N_315);
nor U1071 (N_1071,N_208,N_387);
and U1072 (N_1072,N_561,N_127);
nor U1073 (N_1073,N_431,N_398);
or U1074 (N_1074,N_225,N_327);
and U1075 (N_1075,N_142,N_541);
nand U1076 (N_1076,N_122,N_269);
xnor U1077 (N_1077,N_153,N_345);
nor U1078 (N_1078,N_16,N_128);
or U1079 (N_1079,N_280,N_561);
nand U1080 (N_1080,N_121,N_450);
and U1081 (N_1081,N_432,N_130);
xor U1082 (N_1082,N_75,N_336);
xnor U1083 (N_1083,N_166,N_409);
or U1084 (N_1084,N_304,N_462);
nand U1085 (N_1085,N_142,N_169);
and U1086 (N_1086,N_184,N_497);
xnor U1087 (N_1087,N_175,N_122);
nand U1088 (N_1088,N_568,N_440);
nand U1089 (N_1089,N_190,N_352);
and U1090 (N_1090,N_89,N_295);
and U1091 (N_1091,N_452,N_522);
nand U1092 (N_1092,N_392,N_240);
nor U1093 (N_1093,N_306,N_592);
nor U1094 (N_1094,N_80,N_446);
nor U1095 (N_1095,N_234,N_148);
xor U1096 (N_1096,N_273,N_310);
xnor U1097 (N_1097,N_445,N_592);
and U1098 (N_1098,N_148,N_142);
nor U1099 (N_1099,N_577,N_447);
nor U1100 (N_1100,N_511,N_539);
or U1101 (N_1101,N_64,N_3);
nand U1102 (N_1102,N_105,N_417);
nor U1103 (N_1103,N_29,N_129);
and U1104 (N_1104,N_379,N_62);
or U1105 (N_1105,N_513,N_421);
and U1106 (N_1106,N_133,N_442);
or U1107 (N_1107,N_74,N_196);
nand U1108 (N_1108,N_549,N_487);
and U1109 (N_1109,N_246,N_307);
nor U1110 (N_1110,N_593,N_292);
or U1111 (N_1111,N_77,N_581);
xor U1112 (N_1112,N_581,N_312);
and U1113 (N_1113,N_509,N_48);
and U1114 (N_1114,N_58,N_79);
nand U1115 (N_1115,N_457,N_86);
and U1116 (N_1116,N_346,N_400);
nand U1117 (N_1117,N_126,N_490);
xor U1118 (N_1118,N_1,N_411);
xnor U1119 (N_1119,N_285,N_457);
nand U1120 (N_1120,N_27,N_412);
nand U1121 (N_1121,N_462,N_486);
or U1122 (N_1122,N_364,N_571);
nor U1123 (N_1123,N_379,N_392);
or U1124 (N_1124,N_579,N_563);
nor U1125 (N_1125,N_302,N_89);
and U1126 (N_1126,N_403,N_494);
and U1127 (N_1127,N_64,N_15);
nand U1128 (N_1128,N_532,N_12);
nor U1129 (N_1129,N_332,N_83);
xnor U1130 (N_1130,N_187,N_474);
nand U1131 (N_1131,N_452,N_13);
and U1132 (N_1132,N_226,N_7);
or U1133 (N_1133,N_90,N_374);
and U1134 (N_1134,N_119,N_459);
nand U1135 (N_1135,N_556,N_212);
or U1136 (N_1136,N_421,N_580);
or U1137 (N_1137,N_175,N_395);
nor U1138 (N_1138,N_261,N_71);
xnor U1139 (N_1139,N_354,N_233);
or U1140 (N_1140,N_501,N_340);
nor U1141 (N_1141,N_516,N_438);
nand U1142 (N_1142,N_342,N_162);
nor U1143 (N_1143,N_588,N_110);
or U1144 (N_1144,N_525,N_292);
nor U1145 (N_1145,N_91,N_412);
and U1146 (N_1146,N_425,N_588);
or U1147 (N_1147,N_443,N_280);
and U1148 (N_1148,N_339,N_590);
or U1149 (N_1149,N_357,N_321);
and U1150 (N_1150,N_524,N_159);
and U1151 (N_1151,N_558,N_200);
nand U1152 (N_1152,N_302,N_496);
xnor U1153 (N_1153,N_483,N_504);
nand U1154 (N_1154,N_46,N_349);
nand U1155 (N_1155,N_181,N_32);
nand U1156 (N_1156,N_406,N_306);
nor U1157 (N_1157,N_154,N_585);
xor U1158 (N_1158,N_502,N_287);
nand U1159 (N_1159,N_251,N_263);
xor U1160 (N_1160,N_598,N_71);
or U1161 (N_1161,N_307,N_116);
xnor U1162 (N_1162,N_109,N_174);
nor U1163 (N_1163,N_534,N_557);
and U1164 (N_1164,N_59,N_393);
and U1165 (N_1165,N_561,N_567);
or U1166 (N_1166,N_469,N_4);
nand U1167 (N_1167,N_492,N_134);
xor U1168 (N_1168,N_98,N_453);
and U1169 (N_1169,N_189,N_237);
or U1170 (N_1170,N_416,N_360);
or U1171 (N_1171,N_144,N_526);
and U1172 (N_1172,N_581,N_590);
or U1173 (N_1173,N_95,N_495);
nor U1174 (N_1174,N_569,N_438);
or U1175 (N_1175,N_274,N_128);
nand U1176 (N_1176,N_145,N_338);
xnor U1177 (N_1177,N_79,N_125);
xor U1178 (N_1178,N_96,N_138);
or U1179 (N_1179,N_112,N_131);
or U1180 (N_1180,N_363,N_71);
nor U1181 (N_1181,N_368,N_433);
nand U1182 (N_1182,N_564,N_450);
and U1183 (N_1183,N_466,N_596);
nor U1184 (N_1184,N_420,N_105);
nor U1185 (N_1185,N_535,N_5);
and U1186 (N_1186,N_50,N_390);
and U1187 (N_1187,N_125,N_53);
or U1188 (N_1188,N_372,N_480);
xor U1189 (N_1189,N_544,N_73);
nor U1190 (N_1190,N_236,N_551);
xor U1191 (N_1191,N_560,N_146);
xor U1192 (N_1192,N_212,N_162);
nor U1193 (N_1193,N_582,N_259);
nor U1194 (N_1194,N_359,N_230);
and U1195 (N_1195,N_271,N_322);
and U1196 (N_1196,N_346,N_267);
or U1197 (N_1197,N_87,N_383);
xnor U1198 (N_1198,N_433,N_21);
nand U1199 (N_1199,N_93,N_378);
xnor U1200 (N_1200,N_963,N_962);
xor U1201 (N_1201,N_631,N_958);
nand U1202 (N_1202,N_619,N_1016);
and U1203 (N_1203,N_1005,N_763);
and U1204 (N_1204,N_1108,N_764);
or U1205 (N_1205,N_924,N_901);
and U1206 (N_1206,N_702,N_1123);
or U1207 (N_1207,N_1019,N_951);
xor U1208 (N_1208,N_1192,N_605);
and U1209 (N_1209,N_933,N_711);
nand U1210 (N_1210,N_770,N_860);
and U1211 (N_1211,N_882,N_1105);
xor U1212 (N_1212,N_894,N_768);
or U1213 (N_1213,N_1059,N_613);
or U1214 (N_1214,N_1190,N_993);
xor U1215 (N_1215,N_1037,N_736);
or U1216 (N_1216,N_1022,N_1101);
nor U1217 (N_1217,N_706,N_828);
nor U1218 (N_1218,N_831,N_1011);
nor U1219 (N_1219,N_733,N_809);
or U1220 (N_1220,N_853,N_786);
nand U1221 (N_1221,N_1099,N_723);
xnor U1222 (N_1222,N_679,N_648);
nor U1223 (N_1223,N_720,N_1013);
and U1224 (N_1224,N_703,N_666);
and U1225 (N_1225,N_801,N_713);
nor U1226 (N_1226,N_681,N_928);
nand U1227 (N_1227,N_628,N_603);
xnor U1228 (N_1228,N_1077,N_966);
nand U1229 (N_1229,N_745,N_779);
and U1230 (N_1230,N_717,N_1183);
and U1231 (N_1231,N_908,N_865);
nand U1232 (N_1232,N_1128,N_674);
nand U1233 (N_1233,N_823,N_769);
and U1234 (N_1234,N_1088,N_880);
nor U1235 (N_1235,N_952,N_761);
or U1236 (N_1236,N_1141,N_1159);
nand U1237 (N_1237,N_795,N_610);
and U1238 (N_1238,N_746,N_1180);
xor U1239 (N_1239,N_1142,N_740);
xor U1240 (N_1240,N_800,N_998);
xor U1241 (N_1241,N_689,N_879);
nand U1242 (N_1242,N_615,N_682);
and U1243 (N_1243,N_859,N_1081);
and U1244 (N_1244,N_874,N_611);
nand U1245 (N_1245,N_1127,N_1071);
or U1246 (N_1246,N_930,N_1155);
and U1247 (N_1247,N_1057,N_949);
nand U1248 (N_1248,N_1018,N_622);
nor U1249 (N_1249,N_983,N_917);
nor U1250 (N_1250,N_1032,N_772);
or U1251 (N_1251,N_688,N_721);
nand U1252 (N_1252,N_735,N_905);
and U1253 (N_1253,N_1116,N_939);
and U1254 (N_1254,N_612,N_929);
nand U1255 (N_1255,N_1026,N_766);
nand U1256 (N_1256,N_849,N_1066);
nand U1257 (N_1257,N_658,N_781);
nand U1258 (N_1258,N_1186,N_1198);
xor U1259 (N_1259,N_1104,N_1178);
xnor U1260 (N_1260,N_1028,N_896);
nand U1261 (N_1261,N_953,N_821);
or U1262 (N_1262,N_1034,N_1001);
and U1263 (N_1263,N_1040,N_1045);
or U1264 (N_1264,N_700,N_1119);
nor U1265 (N_1265,N_685,N_1007);
and U1266 (N_1266,N_785,N_1014);
nor U1267 (N_1267,N_641,N_881);
nor U1268 (N_1268,N_707,N_926);
or U1269 (N_1269,N_1134,N_1000);
xnor U1270 (N_1270,N_1164,N_927);
and U1271 (N_1271,N_832,N_1184);
xnor U1272 (N_1272,N_1015,N_1024);
xor U1273 (N_1273,N_1165,N_1096);
nand U1274 (N_1274,N_1163,N_1181);
nor U1275 (N_1275,N_669,N_737);
and U1276 (N_1276,N_825,N_794);
and U1277 (N_1277,N_730,N_1076);
or U1278 (N_1278,N_835,N_959);
or U1279 (N_1279,N_699,N_996);
nor U1280 (N_1280,N_639,N_805);
xor U1281 (N_1281,N_625,N_1038);
nand U1282 (N_1282,N_742,N_784);
or U1283 (N_1283,N_743,N_977);
nand U1284 (N_1284,N_695,N_826);
and U1285 (N_1285,N_891,N_990);
and U1286 (N_1286,N_1167,N_1158);
nand U1287 (N_1287,N_797,N_1130);
nand U1288 (N_1288,N_1042,N_630);
or U1289 (N_1289,N_878,N_1020);
nor U1290 (N_1290,N_969,N_808);
or U1291 (N_1291,N_877,N_621);
or U1292 (N_1292,N_812,N_655);
nor U1293 (N_1293,N_854,N_1097);
xnor U1294 (N_1294,N_637,N_672);
xor U1295 (N_1295,N_961,N_1073);
nand U1296 (N_1296,N_701,N_851);
nand U1297 (N_1297,N_697,N_898);
nor U1298 (N_1298,N_873,N_796);
nor U1299 (N_1299,N_1199,N_943);
and U1300 (N_1300,N_1176,N_845);
or U1301 (N_1301,N_1061,N_938);
or U1302 (N_1302,N_1002,N_614);
nor U1303 (N_1303,N_676,N_843);
or U1304 (N_1304,N_1110,N_607);
or U1305 (N_1305,N_725,N_806);
nand U1306 (N_1306,N_978,N_935);
xnor U1307 (N_1307,N_980,N_678);
nand U1308 (N_1308,N_1033,N_1177);
or U1309 (N_1309,N_753,N_1062);
nor U1310 (N_1310,N_841,N_696);
nand U1311 (N_1311,N_709,N_1052);
nand U1312 (N_1312,N_751,N_1129);
or U1313 (N_1313,N_897,N_1175);
xor U1314 (N_1314,N_632,N_687);
xnor U1315 (N_1315,N_862,N_654);
or U1316 (N_1316,N_955,N_1182);
and U1317 (N_1317,N_757,N_652);
nand U1318 (N_1318,N_738,N_1078);
nand U1319 (N_1319,N_810,N_694);
nand U1320 (N_1320,N_921,N_1030);
and U1321 (N_1321,N_1115,N_1075);
xnor U1322 (N_1322,N_829,N_904);
or U1323 (N_1323,N_732,N_985);
nor U1324 (N_1324,N_778,N_661);
xor U1325 (N_1325,N_762,N_712);
nand U1326 (N_1326,N_1084,N_675);
xnor U1327 (N_1327,N_1055,N_1048);
and U1328 (N_1328,N_1068,N_1072);
and U1329 (N_1329,N_1189,N_1193);
nor U1330 (N_1330,N_923,N_957);
nand U1331 (N_1331,N_680,N_1107);
nand U1332 (N_1332,N_1191,N_657);
or U1333 (N_1333,N_1150,N_686);
or U1334 (N_1334,N_836,N_945);
xor U1335 (N_1335,N_856,N_846);
nand U1336 (N_1336,N_642,N_988);
or U1337 (N_1337,N_665,N_649);
nor U1338 (N_1338,N_1023,N_1169);
or U1339 (N_1339,N_1140,N_1044);
nand U1340 (N_1340,N_1118,N_1010);
nand U1341 (N_1341,N_1122,N_872);
xor U1342 (N_1342,N_914,N_875);
or U1343 (N_1343,N_1195,N_827);
nor U1344 (N_1344,N_1166,N_997);
nand U1345 (N_1345,N_724,N_1079);
nor U1346 (N_1346,N_931,N_1156);
and U1347 (N_1347,N_1106,N_972);
xnor U1348 (N_1348,N_1171,N_1113);
nand U1349 (N_1349,N_774,N_1069);
or U1350 (N_1350,N_602,N_1082);
nor U1351 (N_1351,N_918,N_604);
or U1352 (N_1352,N_729,N_866);
nand U1353 (N_1353,N_705,N_989);
nor U1354 (N_1354,N_1058,N_600);
nand U1355 (N_1355,N_667,N_964);
or U1356 (N_1356,N_822,N_792);
nand U1357 (N_1357,N_671,N_876);
or U1358 (N_1358,N_967,N_660);
nor U1359 (N_1359,N_787,N_1070);
and U1360 (N_1360,N_965,N_635);
nand U1361 (N_1361,N_1021,N_818);
nand U1362 (N_1362,N_920,N_902);
xor U1363 (N_1363,N_1086,N_1132);
nand U1364 (N_1364,N_889,N_1196);
xor U1365 (N_1365,N_858,N_728);
or U1366 (N_1366,N_870,N_793);
xnor U1367 (N_1367,N_861,N_645);
and U1368 (N_1368,N_994,N_1157);
nand U1369 (N_1369,N_925,N_1187);
and U1370 (N_1370,N_629,N_995);
and U1371 (N_1371,N_884,N_1065);
nand U1372 (N_1372,N_1095,N_773);
nand U1373 (N_1373,N_906,N_1102);
nor U1374 (N_1374,N_814,N_932);
and U1375 (N_1375,N_1039,N_704);
or U1376 (N_1376,N_815,N_819);
nor U1377 (N_1377,N_1146,N_775);
or U1378 (N_1378,N_886,N_1036);
nand U1379 (N_1379,N_782,N_1089);
nor U1380 (N_1380,N_1139,N_971);
nor U1381 (N_1381,N_1017,N_948);
and U1382 (N_1382,N_1053,N_783);
xnor U1383 (N_1383,N_893,N_895);
or U1384 (N_1384,N_1092,N_1025);
and U1385 (N_1385,N_734,N_767);
and U1386 (N_1386,N_677,N_760);
nor U1387 (N_1387,N_907,N_912);
and U1388 (N_1388,N_991,N_747);
nor U1389 (N_1389,N_1029,N_754);
nand U1390 (N_1390,N_975,N_1083);
nor U1391 (N_1391,N_864,N_950);
xnor U1392 (N_1392,N_651,N_1056);
xnor U1393 (N_1393,N_739,N_617);
nand U1394 (N_1394,N_911,N_976);
nand U1395 (N_1395,N_840,N_1094);
nand U1396 (N_1396,N_634,N_1136);
xor U1397 (N_1397,N_1012,N_620);
and U1398 (N_1398,N_834,N_662);
nor U1399 (N_1399,N_922,N_1074);
xor U1400 (N_1400,N_776,N_1063);
xnor U1401 (N_1401,N_1148,N_718);
nand U1402 (N_1402,N_1172,N_1145);
nor U1403 (N_1403,N_839,N_656);
nor U1404 (N_1404,N_863,N_1137);
nand U1405 (N_1405,N_1047,N_616);
nand U1406 (N_1406,N_624,N_608);
nor U1407 (N_1407,N_892,N_1133);
nand U1408 (N_1408,N_986,N_788);
nor U1409 (N_1409,N_716,N_982);
and U1410 (N_1410,N_744,N_749);
xnor U1411 (N_1411,N_1009,N_1138);
xnor U1412 (N_1412,N_992,N_1046);
and U1413 (N_1413,N_946,N_643);
and U1414 (N_1414,N_811,N_1160);
nand U1415 (N_1415,N_693,N_979);
nand U1416 (N_1416,N_910,N_1008);
nand U1417 (N_1417,N_1147,N_1185);
nand U1418 (N_1418,N_623,N_937);
or U1419 (N_1419,N_1112,N_1173);
and U1420 (N_1420,N_683,N_1091);
nand U1421 (N_1421,N_941,N_719);
nand U1422 (N_1422,N_1087,N_999);
nor U1423 (N_1423,N_1174,N_606);
xor U1424 (N_1424,N_844,N_981);
or U1425 (N_1425,N_817,N_903);
and U1426 (N_1426,N_802,N_653);
nor U1427 (N_1427,N_644,N_640);
nor U1428 (N_1428,N_633,N_916);
or U1429 (N_1429,N_942,N_1135);
nand U1430 (N_1430,N_636,N_867);
and U1431 (N_1431,N_650,N_1170);
nor U1432 (N_1432,N_900,N_714);
nand U1433 (N_1433,N_838,N_627);
or U1434 (N_1434,N_1114,N_816);
nand U1435 (N_1435,N_1064,N_771);
nand U1436 (N_1436,N_1050,N_890);
and U1437 (N_1437,N_1080,N_847);
nand U1438 (N_1438,N_1149,N_944);
or U1439 (N_1439,N_791,N_1197);
and U1440 (N_1440,N_752,N_710);
and U1441 (N_1441,N_885,N_765);
nand U1442 (N_1442,N_837,N_698);
xnor U1443 (N_1443,N_1124,N_807);
nand U1444 (N_1444,N_646,N_915);
nand U1445 (N_1445,N_813,N_690);
nand U1446 (N_1446,N_1098,N_647);
and U1447 (N_1447,N_974,N_601);
and U1448 (N_1448,N_868,N_1111);
nand U1449 (N_1449,N_1162,N_855);
and U1450 (N_1450,N_970,N_1093);
nor U1451 (N_1451,N_1194,N_715);
xor U1452 (N_1452,N_684,N_798);
xnor U1453 (N_1453,N_842,N_947);
or U1454 (N_1454,N_618,N_659);
nand U1455 (N_1455,N_1003,N_799);
nand U1456 (N_1456,N_1043,N_850);
nand U1457 (N_1457,N_987,N_664);
and U1458 (N_1458,N_1027,N_824);
and U1459 (N_1459,N_750,N_759);
or U1460 (N_1460,N_1161,N_869);
and U1461 (N_1461,N_1085,N_833);
nand U1462 (N_1462,N_954,N_899);
and U1463 (N_1463,N_984,N_804);
and U1464 (N_1464,N_726,N_848);
xnor U1465 (N_1465,N_1126,N_1188);
xnor U1466 (N_1466,N_727,N_609);
or U1467 (N_1467,N_1131,N_871);
nand U1468 (N_1468,N_692,N_1153);
xor U1469 (N_1469,N_968,N_909);
nand U1470 (N_1470,N_820,N_1006);
and U1471 (N_1471,N_790,N_780);
xor U1472 (N_1472,N_626,N_960);
xnor U1473 (N_1473,N_670,N_956);
or U1474 (N_1474,N_1100,N_1067);
nor U1475 (N_1475,N_1143,N_1121);
nand U1476 (N_1476,N_722,N_852);
and U1477 (N_1477,N_1090,N_731);
and U1478 (N_1478,N_973,N_1120);
nand U1479 (N_1479,N_1151,N_673);
nand U1480 (N_1480,N_1035,N_638);
nand U1481 (N_1481,N_748,N_741);
nand U1482 (N_1482,N_936,N_1103);
nand U1483 (N_1483,N_1041,N_883);
and U1484 (N_1484,N_1049,N_1125);
and U1485 (N_1485,N_1054,N_755);
and U1486 (N_1486,N_777,N_1154);
nor U1487 (N_1487,N_758,N_663);
nand U1488 (N_1488,N_934,N_1051);
nor U1489 (N_1489,N_1004,N_888);
nand U1490 (N_1490,N_691,N_1179);
or U1491 (N_1491,N_708,N_668);
or U1492 (N_1492,N_1144,N_940);
and U1493 (N_1493,N_803,N_830);
xor U1494 (N_1494,N_913,N_1109);
and U1495 (N_1495,N_1031,N_789);
and U1496 (N_1496,N_756,N_1060);
xnor U1497 (N_1497,N_1152,N_919);
or U1498 (N_1498,N_887,N_1168);
or U1499 (N_1499,N_857,N_1117);
and U1500 (N_1500,N_1072,N_952);
nand U1501 (N_1501,N_1133,N_601);
nand U1502 (N_1502,N_1034,N_875);
nor U1503 (N_1503,N_840,N_985);
and U1504 (N_1504,N_1188,N_1166);
nand U1505 (N_1505,N_979,N_733);
nand U1506 (N_1506,N_708,N_805);
xnor U1507 (N_1507,N_916,N_919);
or U1508 (N_1508,N_640,N_1119);
or U1509 (N_1509,N_1135,N_636);
nand U1510 (N_1510,N_1028,N_882);
or U1511 (N_1511,N_656,N_637);
or U1512 (N_1512,N_986,N_963);
xor U1513 (N_1513,N_918,N_755);
and U1514 (N_1514,N_653,N_801);
xor U1515 (N_1515,N_620,N_838);
or U1516 (N_1516,N_1110,N_1174);
nor U1517 (N_1517,N_978,N_966);
nor U1518 (N_1518,N_1150,N_1159);
nor U1519 (N_1519,N_625,N_617);
nand U1520 (N_1520,N_1105,N_845);
or U1521 (N_1521,N_1101,N_805);
xor U1522 (N_1522,N_955,N_871);
nand U1523 (N_1523,N_831,N_1013);
nand U1524 (N_1524,N_904,N_1182);
nor U1525 (N_1525,N_1106,N_1122);
xor U1526 (N_1526,N_898,N_1101);
nor U1527 (N_1527,N_807,N_611);
nand U1528 (N_1528,N_976,N_603);
or U1529 (N_1529,N_802,N_1098);
nand U1530 (N_1530,N_707,N_1007);
xor U1531 (N_1531,N_1007,N_961);
nor U1532 (N_1532,N_621,N_745);
nand U1533 (N_1533,N_877,N_1168);
and U1534 (N_1534,N_1029,N_876);
or U1535 (N_1535,N_785,N_667);
nor U1536 (N_1536,N_981,N_1148);
nand U1537 (N_1537,N_941,N_671);
or U1538 (N_1538,N_984,N_664);
or U1539 (N_1539,N_758,N_678);
and U1540 (N_1540,N_1058,N_764);
and U1541 (N_1541,N_650,N_880);
xnor U1542 (N_1542,N_882,N_819);
and U1543 (N_1543,N_753,N_719);
and U1544 (N_1544,N_1018,N_865);
or U1545 (N_1545,N_998,N_731);
nand U1546 (N_1546,N_951,N_843);
xor U1547 (N_1547,N_831,N_994);
or U1548 (N_1548,N_812,N_605);
and U1549 (N_1549,N_1115,N_776);
nor U1550 (N_1550,N_769,N_709);
xor U1551 (N_1551,N_956,N_1103);
nor U1552 (N_1552,N_702,N_928);
xor U1553 (N_1553,N_614,N_1022);
nor U1554 (N_1554,N_762,N_778);
and U1555 (N_1555,N_638,N_1021);
and U1556 (N_1556,N_948,N_865);
or U1557 (N_1557,N_601,N_867);
or U1558 (N_1558,N_873,N_1173);
xor U1559 (N_1559,N_698,N_1195);
nor U1560 (N_1560,N_706,N_848);
xnor U1561 (N_1561,N_992,N_1088);
nor U1562 (N_1562,N_1061,N_779);
and U1563 (N_1563,N_1157,N_823);
xor U1564 (N_1564,N_1007,N_855);
nor U1565 (N_1565,N_1111,N_1105);
xnor U1566 (N_1566,N_1005,N_982);
or U1567 (N_1567,N_664,N_1184);
and U1568 (N_1568,N_978,N_883);
and U1569 (N_1569,N_687,N_1107);
and U1570 (N_1570,N_1005,N_837);
or U1571 (N_1571,N_635,N_608);
xnor U1572 (N_1572,N_1028,N_1171);
or U1573 (N_1573,N_614,N_848);
nand U1574 (N_1574,N_956,N_925);
nor U1575 (N_1575,N_1024,N_798);
nor U1576 (N_1576,N_1154,N_680);
nor U1577 (N_1577,N_1058,N_1018);
xnor U1578 (N_1578,N_741,N_607);
and U1579 (N_1579,N_749,N_1043);
and U1580 (N_1580,N_1177,N_768);
xor U1581 (N_1581,N_767,N_714);
xnor U1582 (N_1582,N_1008,N_626);
nor U1583 (N_1583,N_975,N_755);
and U1584 (N_1584,N_653,N_780);
and U1585 (N_1585,N_1196,N_745);
xnor U1586 (N_1586,N_1118,N_634);
nor U1587 (N_1587,N_862,N_765);
xor U1588 (N_1588,N_887,N_1033);
or U1589 (N_1589,N_1012,N_780);
nand U1590 (N_1590,N_1174,N_629);
nand U1591 (N_1591,N_758,N_1183);
xnor U1592 (N_1592,N_1015,N_627);
xnor U1593 (N_1593,N_1141,N_618);
and U1594 (N_1594,N_672,N_924);
xor U1595 (N_1595,N_1083,N_755);
nor U1596 (N_1596,N_825,N_1115);
xnor U1597 (N_1597,N_1194,N_1117);
or U1598 (N_1598,N_1192,N_763);
or U1599 (N_1599,N_638,N_976);
xnor U1600 (N_1600,N_1199,N_693);
nor U1601 (N_1601,N_681,N_722);
xnor U1602 (N_1602,N_885,N_817);
nand U1603 (N_1603,N_1102,N_691);
or U1604 (N_1604,N_1052,N_937);
nor U1605 (N_1605,N_1103,N_919);
or U1606 (N_1606,N_887,N_777);
xnor U1607 (N_1607,N_741,N_743);
nand U1608 (N_1608,N_1111,N_976);
nor U1609 (N_1609,N_720,N_768);
nand U1610 (N_1610,N_1170,N_1114);
nor U1611 (N_1611,N_838,N_1012);
and U1612 (N_1612,N_835,N_825);
nand U1613 (N_1613,N_807,N_1044);
nor U1614 (N_1614,N_639,N_750);
and U1615 (N_1615,N_649,N_882);
nor U1616 (N_1616,N_1116,N_733);
and U1617 (N_1617,N_895,N_766);
and U1618 (N_1618,N_896,N_808);
or U1619 (N_1619,N_1160,N_746);
or U1620 (N_1620,N_1196,N_1042);
nor U1621 (N_1621,N_1088,N_1041);
xnor U1622 (N_1622,N_1134,N_616);
or U1623 (N_1623,N_1140,N_1068);
nand U1624 (N_1624,N_777,N_1172);
nor U1625 (N_1625,N_1092,N_600);
nand U1626 (N_1626,N_794,N_987);
or U1627 (N_1627,N_868,N_1156);
and U1628 (N_1628,N_738,N_782);
nor U1629 (N_1629,N_621,N_759);
nor U1630 (N_1630,N_658,N_627);
xor U1631 (N_1631,N_940,N_1107);
xor U1632 (N_1632,N_815,N_625);
nor U1633 (N_1633,N_1122,N_909);
nor U1634 (N_1634,N_1018,N_1022);
nor U1635 (N_1635,N_685,N_774);
nor U1636 (N_1636,N_710,N_1136);
and U1637 (N_1637,N_742,N_659);
nor U1638 (N_1638,N_990,N_926);
nor U1639 (N_1639,N_1009,N_795);
xor U1640 (N_1640,N_927,N_931);
and U1641 (N_1641,N_847,N_783);
nor U1642 (N_1642,N_1153,N_1053);
or U1643 (N_1643,N_786,N_1044);
nand U1644 (N_1644,N_936,N_827);
nand U1645 (N_1645,N_1193,N_1058);
or U1646 (N_1646,N_797,N_650);
nor U1647 (N_1647,N_1142,N_973);
and U1648 (N_1648,N_968,N_623);
nor U1649 (N_1649,N_1063,N_1075);
and U1650 (N_1650,N_956,N_732);
nor U1651 (N_1651,N_919,N_796);
xnor U1652 (N_1652,N_752,N_1010);
xor U1653 (N_1653,N_1061,N_827);
and U1654 (N_1654,N_1012,N_662);
nor U1655 (N_1655,N_984,N_848);
and U1656 (N_1656,N_745,N_927);
and U1657 (N_1657,N_1093,N_868);
nand U1658 (N_1658,N_1023,N_741);
or U1659 (N_1659,N_694,N_1189);
and U1660 (N_1660,N_875,N_953);
and U1661 (N_1661,N_789,N_754);
nand U1662 (N_1662,N_663,N_1027);
or U1663 (N_1663,N_1011,N_1156);
and U1664 (N_1664,N_713,N_737);
nor U1665 (N_1665,N_1195,N_1103);
or U1666 (N_1666,N_914,N_926);
xnor U1667 (N_1667,N_978,N_1104);
and U1668 (N_1668,N_961,N_789);
nor U1669 (N_1669,N_881,N_817);
or U1670 (N_1670,N_828,N_1156);
xor U1671 (N_1671,N_660,N_1193);
and U1672 (N_1672,N_1122,N_608);
nor U1673 (N_1673,N_1009,N_895);
or U1674 (N_1674,N_828,N_912);
and U1675 (N_1675,N_1029,N_843);
nor U1676 (N_1676,N_967,N_1106);
and U1677 (N_1677,N_920,N_997);
nand U1678 (N_1678,N_1054,N_611);
or U1679 (N_1679,N_610,N_986);
nand U1680 (N_1680,N_1199,N_1022);
nor U1681 (N_1681,N_1036,N_606);
or U1682 (N_1682,N_695,N_999);
xnor U1683 (N_1683,N_663,N_878);
nor U1684 (N_1684,N_905,N_771);
xnor U1685 (N_1685,N_821,N_1167);
nor U1686 (N_1686,N_803,N_952);
nor U1687 (N_1687,N_952,N_1034);
xnor U1688 (N_1688,N_828,N_897);
nand U1689 (N_1689,N_1044,N_994);
nand U1690 (N_1690,N_798,N_781);
nand U1691 (N_1691,N_797,N_759);
and U1692 (N_1692,N_715,N_703);
xor U1693 (N_1693,N_738,N_741);
nand U1694 (N_1694,N_861,N_1059);
nor U1695 (N_1695,N_1155,N_1041);
xnor U1696 (N_1696,N_788,N_859);
xnor U1697 (N_1697,N_999,N_1105);
and U1698 (N_1698,N_633,N_864);
or U1699 (N_1699,N_924,N_680);
and U1700 (N_1700,N_1183,N_870);
nand U1701 (N_1701,N_953,N_608);
nand U1702 (N_1702,N_987,N_818);
nor U1703 (N_1703,N_962,N_1010);
nand U1704 (N_1704,N_1074,N_764);
and U1705 (N_1705,N_1068,N_1059);
and U1706 (N_1706,N_733,N_1169);
xnor U1707 (N_1707,N_979,N_838);
nor U1708 (N_1708,N_849,N_631);
or U1709 (N_1709,N_1008,N_875);
and U1710 (N_1710,N_844,N_890);
and U1711 (N_1711,N_940,N_772);
and U1712 (N_1712,N_878,N_631);
or U1713 (N_1713,N_685,N_1110);
and U1714 (N_1714,N_906,N_704);
or U1715 (N_1715,N_1000,N_938);
nand U1716 (N_1716,N_986,N_1182);
and U1717 (N_1717,N_1082,N_1070);
nand U1718 (N_1718,N_774,N_907);
and U1719 (N_1719,N_1021,N_789);
nor U1720 (N_1720,N_1019,N_1013);
and U1721 (N_1721,N_1099,N_609);
nor U1722 (N_1722,N_993,N_900);
or U1723 (N_1723,N_971,N_867);
nor U1724 (N_1724,N_937,N_959);
nand U1725 (N_1725,N_1141,N_788);
and U1726 (N_1726,N_621,N_1106);
or U1727 (N_1727,N_1005,N_1023);
and U1728 (N_1728,N_885,N_1039);
or U1729 (N_1729,N_1033,N_891);
xor U1730 (N_1730,N_925,N_1018);
nor U1731 (N_1731,N_732,N_687);
nor U1732 (N_1732,N_1032,N_771);
xnor U1733 (N_1733,N_637,N_634);
xor U1734 (N_1734,N_956,N_623);
nor U1735 (N_1735,N_673,N_952);
xor U1736 (N_1736,N_1017,N_1127);
and U1737 (N_1737,N_1083,N_988);
nand U1738 (N_1738,N_636,N_914);
nor U1739 (N_1739,N_1140,N_1186);
nand U1740 (N_1740,N_727,N_785);
and U1741 (N_1741,N_693,N_708);
nor U1742 (N_1742,N_1175,N_996);
xor U1743 (N_1743,N_772,N_962);
nand U1744 (N_1744,N_1092,N_614);
or U1745 (N_1745,N_1114,N_821);
xnor U1746 (N_1746,N_709,N_976);
nand U1747 (N_1747,N_779,N_905);
nand U1748 (N_1748,N_1134,N_891);
nand U1749 (N_1749,N_1152,N_760);
nor U1750 (N_1750,N_784,N_981);
xnor U1751 (N_1751,N_1168,N_736);
or U1752 (N_1752,N_1056,N_900);
and U1753 (N_1753,N_734,N_897);
or U1754 (N_1754,N_956,N_937);
nor U1755 (N_1755,N_688,N_880);
nand U1756 (N_1756,N_1050,N_1154);
nand U1757 (N_1757,N_920,N_667);
xnor U1758 (N_1758,N_946,N_790);
and U1759 (N_1759,N_1151,N_1082);
nor U1760 (N_1760,N_1055,N_696);
xnor U1761 (N_1761,N_1073,N_1037);
xor U1762 (N_1762,N_620,N_942);
or U1763 (N_1763,N_915,N_1170);
nor U1764 (N_1764,N_1073,N_794);
nand U1765 (N_1765,N_649,N_694);
and U1766 (N_1766,N_979,N_803);
xor U1767 (N_1767,N_880,N_1175);
or U1768 (N_1768,N_1029,N_878);
nand U1769 (N_1769,N_882,N_1038);
xor U1770 (N_1770,N_1185,N_1011);
nor U1771 (N_1771,N_802,N_851);
nor U1772 (N_1772,N_751,N_644);
or U1773 (N_1773,N_1054,N_1047);
and U1774 (N_1774,N_803,N_727);
and U1775 (N_1775,N_746,N_806);
nor U1776 (N_1776,N_831,N_1078);
and U1777 (N_1777,N_868,N_882);
xor U1778 (N_1778,N_1111,N_895);
and U1779 (N_1779,N_839,N_971);
xnor U1780 (N_1780,N_911,N_865);
nor U1781 (N_1781,N_861,N_1084);
and U1782 (N_1782,N_1173,N_1120);
xor U1783 (N_1783,N_1062,N_1067);
nand U1784 (N_1784,N_1195,N_648);
or U1785 (N_1785,N_1017,N_997);
nor U1786 (N_1786,N_643,N_1121);
or U1787 (N_1787,N_615,N_964);
or U1788 (N_1788,N_1128,N_894);
or U1789 (N_1789,N_994,N_735);
xor U1790 (N_1790,N_1016,N_753);
or U1791 (N_1791,N_841,N_1043);
nand U1792 (N_1792,N_993,N_1171);
nand U1793 (N_1793,N_865,N_625);
nand U1794 (N_1794,N_1075,N_654);
xnor U1795 (N_1795,N_1119,N_917);
or U1796 (N_1796,N_1064,N_758);
and U1797 (N_1797,N_701,N_629);
nor U1798 (N_1798,N_1124,N_761);
and U1799 (N_1799,N_965,N_1034);
nor U1800 (N_1800,N_1783,N_1581);
xor U1801 (N_1801,N_1537,N_1530);
xor U1802 (N_1802,N_1413,N_1732);
xor U1803 (N_1803,N_1524,N_1308);
xnor U1804 (N_1804,N_1664,N_1327);
and U1805 (N_1805,N_1686,N_1291);
or U1806 (N_1806,N_1543,N_1339);
and U1807 (N_1807,N_1427,N_1400);
nand U1808 (N_1808,N_1222,N_1466);
and U1809 (N_1809,N_1408,N_1425);
nand U1810 (N_1810,N_1301,N_1557);
nor U1811 (N_1811,N_1628,N_1292);
xnor U1812 (N_1812,N_1217,N_1658);
or U1813 (N_1813,N_1283,N_1406);
and U1814 (N_1814,N_1680,N_1617);
xnor U1815 (N_1815,N_1395,N_1643);
and U1816 (N_1816,N_1439,N_1546);
xnor U1817 (N_1817,N_1312,N_1355);
nor U1818 (N_1818,N_1679,N_1706);
xor U1819 (N_1819,N_1422,N_1349);
and U1820 (N_1820,N_1377,N_1755);
nand U1821 (N_1821,N_1527,N_1762);
nor U1822 (N_1822,N_1372,N_1363);
nor U1823 (N_1823,N_1616,N_1502);
or U1824 (N_1824,N_1671,N_1402);
and U1825 (N_1825,N_1214,N_1249);
and U1826 (N_1826,N_1510,N_1490);
or U1827 (N_1827,N_1766,N_1500);
or U1828 (N_1828,N_1273,N_1541);
nor U1829 (N_1829,N_1626,N_1412);
or U1830 (N_1830,N_1202,N_1397);
or U1831 (N_1831,N_1352,N_1242);
nor U1832 (N_1832,N_1236,N_1358);
xor U1833 (N_1833,N_1704,N_1648);
xor U1834 (N_1834,N_1277,N_1208);
nand U1835 (N_1835,N_1653,N_1730);
nand U1836 (N_1836,N_1369,N_1305);
nor U1837 (N_1837,N_1359,N_1348);
nor U1838 (N_1838,N_1434,N_1216);
nand U1839 (N_1839,N_1230,N_1205);
nand U1840 (N_1840,N_1670,N_1209);
xor U1841 (N_1841,N_1331,N_1615);
nand U1842 (N_1842,N_1651,N_1266);
nand U1843 (N_1843,N_1503,N_1523);
xor U1844 (N_1844,N_1221,N_1442);
nand U1845 (N_1845,N_1765,N_1746);
xor U1846 (N_1846,N_1380,N_1280);
or U1847 (N_1847,N_1409,N_1711);
and U1848 (N_1848,N_1593,N_1575);
xor U1849 (N_1849,N_1788,N_1685);
xor U1850 (N_1850,N_1640,N_1271);
or U1851 (N_1851,N_1346,N_1726);
nor U1852 (N_1852,N_1549,N_1660);
nand U1853 (N_1853,N_1274,N_1411);
or U1854 (N_1854,N_1340,N_1754);
xor U1855 (N_1855,N_1389,N_1529);
nand U1856 (N_1856,N_1451,N_1764);
xnor U1857 (N_1857,N_1513,N_1716);
or U1858 (N_1858,N_1356,N_1384);
nand U1859 (N_1859,N_1371,N_1600);
and U1860 (N_1860,N_1335,N_1319);
or U1861 (N_1861,N_1775,N_1342);
or U1862 (N_1862,N_1784,N_1579);
xor U1863 (N_1863,N_1486,N_1370);
nor U1864 (N_1864,N_1611,N_1360);
or U1865 (N_1865,N_1731,N_1646);
xnor U1866 (N_1866,N_1692,N_1580);
xor U1867 (N_1867,N_1298,N_1394);
or U1868 (N_1868,N_1390,N_1769);
xor U1869 (N_1869,N_1760,N_1487);
nand U1870 (N_1870,N_1578,N_1694);
and U1871 (N_1871,N_1554,N_1744);
nor U1872 (N_1872,N_1213,N_1588);
or U1873 (N_1873,N_1225,N_1777);
xnor U1874 (N_1874,N_1673,N_1666);
nor U1875 (N_1875,N_1376,N_1753);
nor U1876 (N_1876,N_1682,N_1337);
and U1877 (N_1877,N_1304,N_1798);
or U1878 (N_1878,N_1248,N_1668);
nand U1879 (N_1879,N_1599,N_1404);
and U1880 (N_1880,N_1498,N_1226);
nor U1881 (N_1881,N_1459,N_1388);
nor U1882 (N_1882,N_1343,N_1489);
nor U1883 (N_1883,N_1696,N_1661);
xor U1884 (N_1884,N_1284,N_1454);
xor U1885 (N_1885,N_1734,N_1574);
nor U1886 (N_1886,N_1620,N_1756);
nor U1887 (N_1887,N_1547,N_1642);
xor U1888 (N_1888,N_1624,N_1234);
nor U1889 (N_1889,N_1576,N_1649);
xnor U1890 (N_1890,N_1258,N_1470);
and U1891 (N_1891,N_1430,N_1573);
or U1892 (N_1892,N_1458,N_1311);
or U1893 (N_1893,N_1598,N_1220);
xnor U1894 (N_1894,N_1597,N_1505);
nor U1895 (N_1895,N_1351,N_1431);
xor U1896 (N_1896,N_1545,N_1347);
nor U1897 (N_1897,N_1508,N_1595);
nand U1898 (N_1898,N_1367,N_1307);
and U1899 (N_1899,N_1636,N_1594);
nand U1900 (N_1900,N_1771,N_1428);
and U1901 (N_1901,N_1210,N_1296);
xor U1902 (N_1902,N_1718,N_1251);
nand U1903 (N_1903,N_1647,N_1203);
xor U1904 (N_1904,N_1538,N_1279);
xor U1905 (N_1905,N_1644,N_1794);
nand U1906 (N_1906,N_1715,N_1577);
xor U1907 (N_1907,N_1767,N_1678);
nand U1908 (N_1908,N_1344,N_1714);
and U1909 (N_1909,N_1478,N_1219);
nor U1910 (N_1910,N_1385,N_1691);
nand U1911 (N_1911,N_1269,N_1460);
nor U1912 (N_1912,N_1623,N_1495);
nor U1913 (N_1913,N_1420,N_1447);
nand U1914 (N_1914,N_1432,N_1608);
and U1915 (N_1915,N_1776,N_1528);
nand U1916 (N_1916,N_1603,N_1584);
and U1917 (N_1917,N_1382,N_1561);
nor U1918 (N_1918,N_1614,N_1493);
xor U1919 (N_1919,N_1381,N_1281);
nor U1920 (N_1920,N_1733,N_1695);
nor U1921 (N_1921,N_1738,N_1638);
nor U1922 (N_1922,N_1383,N_1270);
nor U1923 (N_1923,N_1552,N_1619);
and U1924 (N_1924,N_1635,N_1585);
and U1925 (N_1925,N_1727,N_1795);
nand U1926 (N_1926,N_1450,N_1627);
xnor U1927 (N_1927,N_1229,N_1419);
and U1928 (N_1928,N_1609,N_1272);
and U1929 (N_1929,N_1789,N_1562);
or U1930 (N_1930,N_1496,N_1659);
nand U1931 (N_1931,N_1227,N_1247);
nand U1932 (N_1932,N_1294,N_1749);
nor U1933 (N_1933,N_1278,N_1518);
or U1934 (N_1934,N_1309,N_1268);
xor U1935 (N_1935,N_1590,N_1736);
xnor U1936 (N_1936,N_1472,N_1433);
and U1937 (N_1937,N_1793,N_1375);
or U1938 (N_1938,N_1534,N_1318);
nor U1939 (N_1939,N_1414,N_1260);
or U1940 (N_1940,N_1297,N_1633);
nor U1941 (N_1941,N_1519,N_1778);
and U1942 (N_1942,N_1437,N_1449);
nor U1943 (N_1943,N_1515,N_1607);
or U1944 (N_1944,N_1403,N_1483);
and U1945 (N_1945,N_1672,N_1630);
nand U1946 (N_1946,N_1265,N_1699);
xor U1947 (N_1947,N_1206,N_1322);
and U1948 (N_1948,N_1768,N_1740);
and U1949 (N_1949,N_1444,N_1326);
nor U1950 (N_1950,N_1758,N_1463);
xnor U1951 (N_1951,N_1315,N_1462);
xor U1952 (N_1952,N_1485,N_1325);
xor U1953 (N_1953,N_1737,N_1641);
nor U1954 (N_1954,N_1548,N_1407);
nand U1955 (N_1955,N_1567,N_1338);
nor U1956 (N_1956,N_1742,N_1401);
nand U1957 (N_1957,N_1482,N_1316);
or U1958 (N_1958,N_1332,N_1514);
and U1959 (N_1959,N_1566,N_1448);
xnor U1960 (N_1960,N_1512,N_1453);
nand U1961 (N_1961,N_1417,N_1424);
nand U1962 (N_1962,N_1582,N_1314);
nand U1963 (N_1963,N_1473,N_1681);
nor U1964 (N_1964,N_1479,N_1387);
or U1965 (N_1965,N_1386,N_1378);
and U1966 (N_1966,N_1440,N_1725);
xor U1967 (N_1967,N_1781,N_1701);
xor U1968 (N_1968,N_1465,N_1204);
nand U1969 (N_1969,N_1717,N_1622);
nand U1970 (N_1970,N_1361,N_1257);
and U1971 (N_1971,N_1405,N_1264);
and U1972 (N_1972,N_1583,N_1320);
nor U1973 (N_1973,N_1750,N_1586);
xor U1974 (N_1974,N_1262,N_1475);
nand U1975 (N_1975,N_1391,N_1558);
or U1976 (N_1976,N_1520,N_1739);
xor U1977 (N_1977,N_1511,N_1263);
nand U1978 (N_1978,N_1488,N_1243);
and U1979 (N_1979,N_1572,N_1504);
nor U1980 (N_1980,N_1313,N_1341);
and U1981 (N_1981,N_1521,N_1244);
nor U1982 (N_1982,N_1667,N_1569);
nor U1983 (N_1983,N_1565,N_1729);
nor U1984 (N_1984,N_1741,N_1452);
or U1985 (N_1985,N_1759,N_1790);
or U1986 (N_1986,N_1366,N_1613);
nand U1987 (N_1987,N_1492,N_1555);
or U1988 (N_1988,N_1791,N_1568);
nor U1989 (N_1989,N_1350,N_1751);
nor U1990 (N_1990,N_1589,N_1663);
or U1991 (N_1991,N_1396,N_1207);
nor U1992 (N_1992,N_1445,N_1708);
or U1993 (N_1993,N_1772,N_1542);
or U1994 (N_1994,N_1656,N_1215);
nand U1995 (N_1995,N_1329,N_1373);
or U1996 (N_1996,N_1393,N_1665);
and U1997 (N_1997,N_1255,N_1621);
xor U1998 (N_1998,N_1480,N_1532);
xnor U1999 (N_1999,N_1392,N_1398);
or U2000 (N_2000,N_1233,N_1293);
nor U2001 (N_2001,N_1299,N_1774);
nor U2002 (N_2002,N_1645,N_1629);
xnor U2003 (N_2003,N_1232,N_1639);
and U2004 (N_2004,N_1415,N_1353);
nand U2005 (N_2005,N_1700,N_1256);
xor U2006 (N_2006,N_1357,N_1559);
xor U2007 (N_2007,N_1724,N_1416);
or U2008 (N_2008,N_1709,N_1719);
or U2009 (N_2009,N_1650,N_1362);
and U2010 (N_2010,N_1522,N_1735);
or U2011 (N_2011,N_1379,N_1334);
nor U2012 (N_2012,N_1637,N_1275);
nor U2013 (N_2013,N_1787,N_1757);
xor U2014 (N_2014,N_1231,N_1752);
or U2015 (N_2015,N_1295,N_1779);
and U2016 (N_2016,N_1517,N_1228);
or U2017 (N_2017,N_1245,N_1618);
nor U2018 (N_2018,N_1720,N_1797);
and U2019 (N_2019,N_1687,N_1596);
nand U2020 (N_2020,N_1556,N_1745);
nand U2021 (N_2021,N_1282,N_1276);
nand U2022 (N_2022,N_1604,N_1662);
or U2023 (N_2023,N_1399,N_1410);
and U2024 (N_2024,N_1421,N_1728);
or U2025 (N_2025,N_1368,N_1551);
nand U2026 (N_2026,N_1698,N_1300);
or U2027 (N_2027,N_1476,N_1669);
xor U2028 (N_2028,N_1443,N_1455);
xnor U2029 (N_2029,N_1484,N_1799);
nand U2030 (N_2030,N_1655,N_1782);
and U2031 (N_2031,N_1238,N_1286);
or U2032 (N_2032,N_1654,N_1336);
xnor U2033 (N_2033,N_1501,N_1533);
xor U2034 (N_2034,N_1212,N_1634);
xor U2035 (N_2035,N_1710,N_1693);
xor U2036 (N_2036,N_1536,N_1345);
or U2037 (N_2037,N_1702,N_1540);
nor U2038 (N_2038,N_1683,N_1539);
or U2039 (N_2039,N_1571,N_1535);
or U2040 (N_2040,N_1306,N_1241);
nand U2041 (N_2041,N_1606,N_1526);
or U2042 (N_2042,N_1288,N_1773);
nand U2043 (N_2043,N_1516,N_1761);
nand U2044 (N_2044,N_1612,N_1235);
xor U2045 (N_2045,N_1200,N_1324);
and U2046 (N_2046,N_1441,N_1748);
nand U2047 (N_2047,N_1677,N_1477);
xnor U2048 (N_2048,N_1457,N_1317);
nand U2049 (N_2049,N_1328,N_1261);
nand U2050 (N_2050,N_1509,N_1223);
and U2051 (N_2051,N_1446,N_1239);
nor U2052 (N_2052,N_1330,N_1497);
xnor U2053 (N_2053,N_1438,N_1252);
or U2054 (N_2054,N_1610,N_1246);
or U2055 (N_2055,N_1747,N_1770);
and U2056 (N_2056,N_1436,N_1707);
xor U2057 (N_2057,N_1550,N_1601);
and U2058 (N_2058,N_1254,N_1560);
and U2059 (N_2059,N_1602,N_1285);
xnor U2060 (N_2060,N_1786,N_1652);
xnor U2061 (N_2061,N_1570,N_1302);
nand U2062 (N_2062,N_1250,N_1464);
or U2063 (N_2063,N_1723,N_1625);
nand U2064 (N_2064,N_1657,N_1310);
nor U2065 (N_2065,N_1321,N_1267);
and U2066 (N_2066,N_1674,N_1237);
xnor U2067 (N_2067,N_1323,N_1333);
xnor U2068 (N_2068,N_1697,N_1763);
or U2069 (N_2069,N_1364,N_1259);
nor U2070 (N_2070,N_1494,N_1531);
and U2071 (N_2071,N_1544,N_1469);
nand U2072 (N_2072,N_1743,N_1564);
and U2073 (N_2073,N_1632,N_1365);
xor U2074 (N_2074,N_1592,N_1499);
nand U2075 (N_2075,N_1481,N_1418);
and U2076 (N_2076,N_1461,N_1224);
nand U2077 (N_2077,N_1553,N_1506);
and U2078 (N_2078,N_1423,N_1525);
and U2079 (N_2079,N_1240,N_1796);
nand U2080 (N_2080,N_1675,N_1491);
or U2081 (N_2081,N_1201,N_1435);
and U2082 (N_2082,N_1605,N_1705);
nand U2083 (N_2083,N_1631,N_1703);
nor U2084 (N_2084,N_1471,N_1689);
nand U2085 (N_2085,N_1303,N_1374);
nor U2086 (N_2086,N_1429,N_1289);
xor U2087 (N_2087,N_1467,N_1780);
nand U2088 (N_2088,N_1785,N_1591);
or U2089 (N_2089,N_1690,N_1792);
or U2090 (N_2090,N_1456,N_1721);
xor U2091 (N_2091,N_1218,N_1563);
and U2092 (N_2092,N_1287,N_1684);
xor U2093 (N_2093,N_1468,N_1507);
or U2094 (N_2094,N_1426,N_1713);
or U2095 (N_2095,N_1474,N_1211);
xnor U2096 (N_2096,N_1722,N_1290);
nor U2097 (N_2097,N_1587,N_1712);
and U2098 (N_2098,N_1676,N_1354);
or U2099 (N_2099,N_1688,N_1253);
and U2100 (N_2100,N_1397,N_1639);
nor U2101 (N_2101,N_1581,N_1227);
xnor U2102 (N_2102,N_1365,N_1246);
or U2103 (N_2103,N_1521,N_1559);
nor U2104 (N_2104,N_1208,N_1461);
nand U2105 (N_2105,N_1544,N_1626);
nor U2106 (N_2106,N_1496,N_1572);
and U2107 (N_2107,N_1678,N_1358);
xnor U2108 (N_2108,N_1614,N_1223);
nand U2109 (N_2109,N_1607,N_1567);
and U2110 (N_2110,N_1309,N_1495);
or U2111 (N_2111,N_1218,N_1437);
nand U2112 (N_2112,N_1668,N_1647);
nor U2113 (N_2113,N_1697,N_1240);
nand U2114 (N_2114,N_1389,N_1613);
or U2115 (N_2115,N_1541,N_1526);
nor U2116 (N_2116,N_1270,N_1726);
or U2117 (N_2117,N_1227,N_1213);
nand U2118 (N_2118,N_1474,N_1677);
xnor U2119 (N_2119,N_1464,N_1215);
xor U2120 (N_2120,N_1730,N_1536);
nor U2121 (N_2121,N_1673,N_1541);
nand U2122 (N_2122,N_1577,N_1542);
or U2123 (N_2123,N_1377,N_1381);
nand U2124 (N_2124,N_1430,N_1368);
xor U2125 (N_2125,N_1508,N_1753);
nor U2126 (N_2126,N_1643,N_1501);
xor U2127 (N_2127,N_1378,N_1208);
nand U2128 (N_2128,N_1415,N_1476);
nand U2129 (N_2129,N_1556,N_1333);
or U2130 (N_2130,N_1523,N_1530);
nor U2131 (N_2131,N_1556,N_1431);
nor U2132 (N_2132,N_1353,N_1239);
nor U2133 (N_2133,N_1379,N_1244);
and U2134 (N_2134,N_1392,N_1786);
xnor U2135 (N_2135,N_1754,N_1418);
xor U2136 (N_2136,N_1788,N_1724);
nand U2137 (N_2137,N_1713,N_1370);
and U2138 (N_2138,N_1238,N_1246);
xor U2139 (N_2139,N_1478,N_1207);
xnor U2140 (N_2140,N_1726,N_1333);
nor U2141 (N_2141,N_1431,N_1318);
and U2142 (N_2142,N_1761,N_1591);
nor U2143 (N_2143,N_1213,N_1513);
or U2144 (N_2144,N_1551,N_1515);
nand U2145 (N_2145,N_1760,N_1522);
and U2146 (N_2146,N_1641,N_1608);
or U2147 (N_2147,N_1507,N_1435);
or U2148 (N_2148,N_1735,N_1567);
or U2149 (N_2149,N_1423,N_1455);
nor U2150 (N_2150,N_1645,N_1510);
nand U2151 (N_2151,N_1471,N_1778);
xnor U2152 (N_2152,N_1480,N_1257);
nor U2153 (N_2153,N_1322,N_1620);
and U2154 (N_2154,N_1492,N_1232);
xor U2155 (N_2155,N_1608,N_1393);
or U2156 (N_2156,N_1408,N_1570);
or U2157 (N_2157,N_1350,N_1609);
xnor U2158 (N_2158,N_1546,N_1443);
nand U2159 (N_2159,N_1683,N_1205);
nor U2160 (N_2160,N_1752,N_1255);
or U2161 (N_2161,N_1635,N_1777);
xnor U2162 (N_2162,N_1308,N_1316);
nand U2163 (N_2163,N_1593,N_1578);
and U2164 (N_2164,N_1332,N_1680);
and U2165 (N_2165,N_1525,N_1739);
or U2166 (N_2166,N_1589,N_1465);
or U2167 (N_2167,N_1487,N_1354);
or U2168 (N_2168,N_1463,N_1764);
or U2169 (N_2169,N_1464,N_1558);
or U2170 (N_2170,N_1732,N_1375);
nor U2171 (N_2171,N_1428,N_1358);
nand U2172 (N_2172,N_1574,N_1413);
and U2173 (N_2173,N_1615,N_1323);
or U2174 (N_2174,N_1762,N_1582);
xnor U2175 (N_2175,N_1556,N_1280);
or U2176 (N_2176,N_1477,N_1618);
xor U2177 (N_2177,N_1704,N_1250);
or U2178 (N_2178,N_1285,N_1283);
nor U2179 (N_2179,N_1373,N_1512);
xor U2180 (N_2180,N_1426,N_1648);
and U2181 (N_2181,N_1692,N_1223);
and U2182 (N_2182,N_1336,N_1728);
nand U2183 (N_2183,N_1318,N_1774);
nor U2184 (N_2184,N_1409,N_1210);
nand U2185 (N_2185,N_1426,N_1441);
nor U2186 (N_2186,N_1420,N_1377);
or U2187 (N_2187,N_1393,N_1246);
xor U2188 (N_2188,N_1234,N_1687);
and U2189 (N_2189,N_1460,N_1329);
nand U2190 (N_2190,N_1308,N_1385);
and U2191 (N_2191,N_1591,N_1297);
xnor U2192 (N_2192,N_1691,N_1425);
nand U2193 (N_2193,N_1687,N_1645);
nand U2194 (N_2194,N_1605,N_1527);
and U2195 (N_2195,N_1594,N_1360);
or U2196 (N_2196,N_1776,N_1590);
or U2197 (N_2197,N_1288,N_1543);
xor U2198 (N_2198,N_1575,N_1403);
and U2199 (N_2199,N_1630,N_1539);
nor U2200 (N_2200,N_1765,N_1469);
and U2201 (N_2201,N_1491,N_1259);
nor U2202 (N_2202,N_1297,N_1597);
and U2203 (N_2203,N_1352,N_1699);
nor U2204 (N_2204,N_1516,N_1694);
xor U2205 (N_2205,N_1259,N_1422);
nor U2206 (N_2206,N_1755,N_1257);
and U2207 (N_2207,N_1709,N_1735);
or U2208 (N_2208,N_1540,N_1271);
xnor U2209 (N_2209,N_1748,N_1699);
nor U2210 (N_2210,N_1650,N_1351);
nor U2211 (N_2211,N_1218,N_1450);
nand U2212 (N_2212,N_1726,N_1379);
nand U2213 (N_2213,N_1739,N_1284);
xnor U2214 (N_2214,N_1670,N_1607);
or U2215 (N_2215,N_1597,N_1716);
nor U2216 (N_2216,N_1550,N_1673);
nand U2217 (N_2217,N_1744,N_1508);
or U2218 (N_2218,N_1277,N_1702);
xnor U2219 (N_2219,N_1226,N_1319);
and U2220 (N_2220,N_1349,N_1370);
nand U2221 (N_2221,N_1326,N_1743);
nor U2222 (N_2222,N_1281,N_1495);
nor U2223 (N_2223,N_1351,N_1691);
or U2224 (N_2224,N_1547,N_1717);
xnor U2225 (N_2225,N_1478,N_1281);
xnor U2226 (N_2226,N_1652,N_1208);
or U2227 (N_2227,N_1577,N_1794);
nor U2228 (N_2228,N_1643,N_1635);
or U2229 (N_2229,N_1259,N_1609);
xnor U2230 (N_2230,N_1249,N_1672);
and U2231 (N_2231,N_1454,N_1351);
nor U2232 (N_2232,N_1535,N_1598);
nand U2233 (N_2233,N_1368,N_1582);
nand U2234 (N_2234,N_1281,N_1244);
nand U2235 (N_2235,N_1623,N_1731);
nor U2236 (N_2236,N_1754,N_1795);
xor U2237 (N_2237,N_1524,N_1715);
nor U2238 (N_2238,N_1788,N_1252);
nand U2239 (N_2239,N_1285,N_1353);
and U2240 (N_2240,N_1766,N_1450);
xor U2241 (N_2241,N_1445,N_1752);
or U2242 (N_2242,N_1595,N_1247);
and U2243 (N_2243,N_1699,N_1353);
or U2244 (N_2244,N_1797,N_1686);
and U2245 (N_2245,N_1419,N_1408);
nor U2246 (N_2246,N_1442,N_1710);
nand U2247 (N_2247,N_1649,N_1375);
nor U2248 (N_2248,N_1768,N_1405);
nand U2249 (N_2249,N_1558,N_1675);
and U2250 (N_2250,N_1767,N_1446);
nand U2251 (N_2251,N_1558,N_1322);
nand U2252 (N_2252,N_1656,N_1373);
and U2253 (N_2253,N_1787,N_1575);
and U2254 (N_2254,N_1673,N_1774);
xor U2255 (N_2255,N_1714,N_1630);
nand U2256 (N_2256,N_1561,N_1542);
nor U2257 (N_2257,N_1544,N_1740);
nor U2258 (N_2258,N_1501,N_1611);
or U2259 (N_2259,N_1605,N_1430);
xnor U2260 (N_2260,N_1203,N_1429);
or U2261 (N_2261,N_1770,N_1614);
or U2262 (N_2262,N_1470,N_1396);
nand U2263 (N_2263,N_1595,N_1473);
nand U2264 (N_2264,N_1444,N_1396);
nand U2265 (N_2265,N_1578,N_1498);
or U2266 (N_2266,N_1539,N_1295);
or U2267 (N_2267,N_1734,N_1354);
and U2268 (N_2268,N_1367,N_1610);
nand U2269 (N_2269,N_1616,N_1310);
and U2270 (N_2270,N_1311,N_1393);
and U2271 (N_2271,N_1623,N_1642);
nand U2272 (N_2272,N_1485,N_1529);
nand U2273 (N_2273,N_1360,N_1636);
or U2274 (N_2274,N_1561,N_1461);
nor U2275 (N_2275,N_1770,N_1606);
nand U2276 (N_2276,N_1582,N_1655);
nand U2277 (N_2277,N_1507,N_1362);
xnor U2278 (N_2278,N_1418,N_1769);
nand U2279 (N_2279,N_1739,N_1524);
or U2280 (N_2280,N_1326,N_1399);
or U2281 (N_2281,N_1670,N_1603);
xnor U2282 (N_2282,N_1547,N_1208);
nor U2283 (N_2283,N_1641,N_1291);
nand U2284 (N_2284,N_1420,N_1384);
nand U2285 (N_2285,N_1560,N_1344);
and U2286 (N_2286,N_1663,N_1312);
nand U2287 (N_2287,N_1744,N_1252);
and U2288 (N_2288,N_1681,N_1365);
nand U2289 (N_2289,N_1328,N_1619);
xnor U2290 (N_2290,N_1575,N_1376);
nand U2291 (N_2291,N_1594,N_1211);
or U2292 (N_2292,N_1221,N_1794);
xnor U2293 (N_2293,N_1600,N_1308);
and U2294 (N_2294,N_1338,N_1598);
or U2295 (N_2295,N_1238,N_1394);
or U2296 (N_2296,N_1279,N_1601);
and U2297 (N_2297,N_1238,N_1362);
nor U2298 (N_2298,N_1525,N_1412);
or U2299 (N_2299,N_1670,N_1694);
xnor U2300 (N_2300,N_1533,N_1646);
xor U2301 (N_2301,N_1677,N_1285);
xnor U2302 (N_2302,N_1652,N_1381);
or U2303 (N_2303,N_1601,N_1620);
and U2304 (N_2304,N_1379,N_1262);
nor U2305 (N_2305,N_1286,N_1614);
nand U2306 (N_2306,N_1359,N_1672);
nand U2307 (N_2307,N_1578,N_1336);
or U2308 (N_2308,N_1771,N_1249);
and U2309 (N_2309,N_1360,N_1430);
or U2310 (N_2310,N_1670,N_1424);
or U2311 (N_2311,N_1408,N_1515);
or U2312 (N_2312,N_1738,N_1407);
or U2313 (N_2313,N_1268,N_1609);
or U2314 (N_2314,N_1284,N_1403);
and U2315 (N_2315,N_1480,N_1445);
or U2316 (N_2316,N_1384,N_1628);
nor U2317 (N_2317,N_1407,N_1744);
nor U2318 (N_2318,N_1763,N_1773);
xor U2319 (N_2319,N_1221,N_1679);
or U2320 (N_2320,N_1771,N_1415);
and U2321 (N_2321,N_1781,N_1201);
nand U2322 (N_2322,N_1389,N_1351);
nand U2323 (N_2323,N_1712,N_1663);
xor U2324 (N_2324,N_1354,N_1520);
xnor U2325 (N_2325,N_1761,N_1609);
nor U2326 (N_2326,N_1433,N_1417);
nor U2327 (N_2327,N_1372,N_1234);
nor U2328 (N_2328,N_1402,N_1689);
or U2329 (N_2329,N_1729,N_1568);
and U2330 (N_2330,N_1400,N_1653);
nor U2331 (N_2331,N_1559,N_1712);
xor U2332 (N_2332,N_1439,N_1529);
or U2333 (N_2333,N_1728,N_1314);
xor U2334 (N_2334,N_1504,N_1380);
nor U2335 (N_2335,N_1766,N_1461);
nor U2336 (N_2336,N_1564,N_1445);
and U2337 (N_2337,N_1611,N_1544);
or U2338 (N_2338,N_1372,N_1750);
and U2339 (N_2339,N_1510,N_1479);
and U2340 (N_2340,N_1299,N_1542);
and U2341 (N_2341,N_1237,N_1578);
xor U2342 (N_2342,N_1747,N_1776);
and U2343 (N_2343,N_1756,N_1472);
nand U2344 (N_2344,N_1697,N_1521);
and U2345 (N_2345,N_1695,N_1475);
or U2346 (N_2346,N_1544,N_1273);
nand U2347 (N_2347,N_1766,N_1287);
nand U2348 (N_2348,N_1258,N_1602);
and U2349 (N_2349,N_1775,N_1694);
nand U2350 (N_2350,N_1210,N_1523);
and U2351 (N_2351,N_1446,N_1280);
nand U2352 (N_2352,N_1629,N_1560);
or U2353 (N_2353,N_1614,N_1553);
and U2354 (N_2354,N_1347,N_1273);
and U2355 (N_2355,N_1284,N_1636);
and U2356 (N_2356,N_1795,N_1213);
nor U2357 (N_2357,N_1420,N_1307);
or U2358 (N_2358,N_1627,N_1535);
or U2359 (N_2359,N_1209,N_1493);
xor U2360 (N_2360,N_1421,N_1629);
nor U2361 (N_2361,N_1698,N_1289);
nand U2362 (N_2362,N_1284,N_1763);
and U2363 (N_2363,N_1219,N_1389);
nor U2364 (N_2364,N_1786,N_1653);
xor U2365 (N_2365,N_1396,N_1244);
nand U2366 (N_2366,N_1401,N_1657);
xnor U2367 (N_2367,N_1756,N_1776);
nand U2368 (N_2368,N_1525,N_1795);
xnor U2369 (N_2369,N_1679,N_1307);
nand U2370 (N_2370,N_1615,N_1375);
nor U2371 (N_2371,N_1313,N_1703);
or U2372 (N_2372,N_1316,N_1611);
xor U2373 (N_2373,N_1488,N_1212);
nand U2374 (N_2374,N_1378,N_1337);
nand U2375 (N_2375,N_1204,N_1623);
nand U2376 (N_2376,N_1371,N_1277);
nand U2377 (N_2377,N_1592,N_1793);
nor U2378 (N_2378,N_1425,N_1579);
or U2379 (N_2379,N_1491,N_1742);
nand U2380 (N_2380,N_1653,N_1475);
or U2381 (N_2381,N_1612,N_1597);
xor U2382 (N_2382,N_1256,N_1240);
or U2383 (N_2383,N_1289,N_1335);
xnor U2384 (N_2384,N_1774,N_1524);
nor U2385 (N_2385,N_1379,N_1695);
nor U2386 (N_2386,N_1553,N_1775);
or U2387 (N_2387,N_1701,N_1648);
xnor U2388 (N_2388,N_1555,N_1244);
or U2389 (N_2389,N_1233,N_1492);
or U2390 (N_2390,N_1325,N_1611);
xor U2391 (N_2391,N_1555,N_1506);
xnor U2392 (N_2392,N_1532,N_1719);
or U2393 (N_2393,N_1420,N_1327);
or U2394 (N_2394,N_1291,N_1231);
xnor U2395 (N_2395,N_1596,N_1528);
xor U2396 (N_2396,N_1366,N_1660);
xor U2397 (N_2397,N_1548,N_1453);
nor U2398 (N_2398,N_1316,N_1703);
and U2399 (N_2399,N_1668,N_1797);
and U2400 (N_2400,N_2009,N_2076);
nor U2401 (N_2401,N_1978,N_2291);
or U2402 (N_2402,N_2176,N_2221);
or U2403 (N_2403,N_1962,N_2129);
or U2404 (N_2404,N_2103,N_1965);
or U2405 (N_2405,N_2100,N_2010);
nor U2406 (N_2406,N_2254,N_2226);
nand U2407 (N_2407,N_2243,N_2182);
nor U2408 (N_2408,N_1901,N_2029);
and U2409 (N_2409,N_2138,N_1808);
or U2410 (N_2410,N_2204,N_1864);
and U2411 (N_2411,N_2005,N_2345);
nand U2412 (N_2412,N_2365,N_2230);
or U2413 (N_2413,N_1963,N_2329);
nor U2414 (N_2414,N_2355,N_2283);
nor U2415 (N_2415,N_2250,N_2170);
or U2416 (N_2416,N_2036,N_1974);
nand U2417 (N_2417,N_2099,N_2341);
nand U2418 (N_2418,N_2232,N_1831);
nand U2419 (N_2419,N_2276,N_2030);
and U2420 (N_2420,N_1926,N_2108);
nor U2421 (N_2421,N_2094,N_2300);
nor U2422 (N_2422,N_2262,N_2368);
or U2423 (N_2423,N_1935,N_2095);
and U2424 (N_2424,N_1896,N_2119);
nor U2425 (N_2425,N_2390,N_1853);
and U2426 (N_2426,N_2375,N_1815);
nor U2427 (N_2427,N_2132,N_2309);
nand U2428 (N_2428,N_2122,N_2091);
or U2429 (N_2429,N_2396,N_2180);
nor U2430 (N_2430,N_2214,N_1918);
nand U2431 (N_2431,N_1872,N_2111);
and U2432 (N_2432,N_2159,N_2225);
nor U2433 (N_2433,N_2001,N_1940);
xnor U2434 (N_2434,N_1929,N_1994);
xor U2435 (N_2435,N_2236,N_2019);
xnor U2436 (N_2436,N_2387,N_2187);
or U2437 (N_2437,N_2231,N_2340);
xnor U2438 (N_2438,N_2248,N_2245);
xor U2439 (N_2439,N_2002,N_1908);
nor U2440 (N_2440,N_2391,N_1984);
nor U2441 (N_2441,N_1989,N_1819);
and U2442 (N_2442,N_2241,N_1813);
and U2443 (N_2443,N_2376,N_2017);
or U2444 (N_2444,N_2163,N_2144);
nor U2445 (N_2445,N_2145,N_1820);
or U2446 (N_2446,N_2217,N_1850);
nor U2447 (N_2447,N_2346,N_2025);
xnor U2448 (N_2448,N_1863,N_2284);
xor U2449 (N_2449,N_1919,N_2066);
nor U2450 (N_2450,N_1964,N_2059);
and U2451 (N_2451,N_2270,N_1828);
nor U2452 (N_2452,N_2125,N_2085);
nand U2453 (N_2453,N_2312,N_1955);
xnor U2454 (N_2454,N_2367,N_1802);
and U2455 (N_2455,N_2344,N_2388);
and U2456 (N_2456,N_2084,N_2318);
nand U2457 (N_2457,N_2303,N_1975);
and U2458 (N_2458,N_1969,N_2165);
nor U2459 (N_2459,N_2149,N_2104);
xnor U2460 (N_2460,N_2354,N_2304);
nand U2461 (N_2461,N_1999,N_2275);
xor U2462 (N_2462,N_2353,N_1959);
xnor U2463 (N_2463,N_2317,N_1846);
or U2464 (N_2464,N_1824,N_1939);
nor U2465 (N_2465,N_1986,N_2299);
nor U2466 (N_2466,N_2126,N_2332);
nor U2467 (N_2467,N_2333,N_2127);
nor U2468 (N_2468,N_2193,N_2361);
or U2469 (N_2469,N_2358,N_1877);
or U2470 (N_2470,N_1875,N_2201);
nand U2471 (N_2471,N_2118,N_1980);
nand U2472 (N_2472,N_2326,N_1928);
nor U2473 (N_2473,N_2296,N_2016);
nor U2474 (N_2474,N_1920,N_1804);
nor U2475 (N_2475,N_2237,N_2351);
nor U2476 (N_2476,N_2208,N_2281);
and U2477 (N_2477,N_1834,N_2142);
or U2478 (N_2478,N_2362,N_2087);
or U2479 (N_2479,N_1899,N_1990);
and U2480 (N_2480,N_2373,N_2280);
nand U2481 (N_2481,N_2013,N_1985);
or U2482 (N_2482,N_1871,N_2392);
nand U2483 (N_2483,N_1858,N_1966);
xor U2484 (N_2484,N_1817,N_1868);
and U2485 (N_2485,N_2377,N_2229);
or U2486 (N_2486,N_2315,N_2020);
nor U2487 (N_2487,N_1997,N_2027);
or U2488 (N_2488,N_2200,N_2109);
nand U2489 (N_2489,N_2289,N_2056);
or U2490 (N_2490,N_2028,N_1810);
or U2491 (N_2491,N_2188,N_2024);
and U2492 (N_2492,N_2181,N_2047);
nand U2493 (N_2493,N_2397,N_1805);
nor U2494 (N_2494,N_2252,N_1952);
nor U2495 (N_2495,N_2139,N_2175);
nor U2496 (N_2496,N_1803,N_1968);
and U2497 (N_2497,N_1931,N_2107);
and U2498 (N_2498,N_1845,N_2324);
and U2499 (N_2499,N_2061,N_1890);
xor U2500 (N_2500,N_2383,N_2366);
or U2501 (N_2501,N_2224,N_2057);
nand U2502 (N_2502,N_2360,N_1888);
or U2503 (N_2503,N_1916,N_1905);
or U2504 (N_2504,N_2342,N_2169);
nand U2505 (N_2505,N_2320,N_2081);
nor U2506 (N_2506,N_1860,N_1891);
xor U2507 (N_2507,N_2302,N_2325);
and U2508 (N_2508,N_2060,N_1949);
nand U2509 (N_2509,N_2082,N_1878);
and U2510 (N_2510,N_2038,N_2316);
nor U2511 (N_2511,N_2268,N_2073);
and U2512 (N_2512,N_2386,N_1937);
and U2513 (N_2513,N_2008,N_1854);
nand U2514 (N_2514,N_2372,N_2018);
and U2515 (N_2515,N_2363,N_2135);
nor U2516 (N_2516,N_1809,N_1900);
xor U2517 (N_2517,N_2247,N_2389);
xnor U2518 (N_2518,N_2161,N_2253);
nand U2519 (N_2519,N_1944,N_2246);
and U2520 (N_2520,N_1814,N_2274);
nor U2521 (N_2521,N_2140,N_2006);
and U2522 (N_2522,N_2301,N_2042);
or U2523 (N_2523,N_2211,N_2065);
or U2524 (N_2524,N_1923,N_1898);
nor U2525 (N_2525,N_2322,N_2216);
or U2526 (N_2526,N_1925,N_2235);
nor U2527 (N_2527,N_2096,N_2157);
nand U2528 (N_2528,N_2278,N_2128);
nand U2529 (N_2529,N_2249,N_2271);
and U2530 (N_2530,N_2151,N_2210);
and U2531 (N_2531,N_2293,N_2043);
xor U2532 (N_2532,N_1822,N_1998);
and U2533 (N_2533,N_2213,N_1823);
and U2534 (N_2534,N_2160,N_1895);
or U2535 (N_2535,N_2046,N_2359);
nor U2536 (N_2536,N_2168,N_1988);
xnor U2537 (N_2537,N_1913,N_1909);
xor U2538 (N_2538,N_2219,N_1880);
and U2539 (N_2539,N_2092,N_1870);
xor U2540 (N_2540,N_1833,N_2032);
and U2541 (N_2541,N_1855,N_1948);
and U2542 (N_2542,N_2069,N_1979);
xor U2543 (N_2543,N_2080,N_2189);
xnor U2544 (N_2544,N_2063,N_1907);
nand U2545 (N_2545,N_1910,N_1865);
nand U2546 (N_2546,N_1973,N_2378);
or U2547 (N_2547,N_1947,N_1945);
nor U2548 (N_2548,N_2053,N_2222);
xor U2549 (N_2549,N_1859,N_1876);
nand U2550 (N_2550,N_1827,N_2295);
nor U2551 (N_2551,N_1861,N_1970);
nand U2552 (N_2552,N_2112,N_2071);
nor U2553 (N_2553,N_2070,N_2348);
xor U2554 (N_2554,N_1921,N_2218);
or U2555 (N_2555,N_2379,N_2220);
or U2556 (N_2556,N_1971,N_2190);
nor U2557 (N_2557,N_2141,N_2055);
nand U2558 (N_2558,N_2259,N_1991);
nor U2559 (N_2559,N_1837,N_2078);
and U2560 (N_2560,N_1912,N_2093);
nor U2561 (N_2561,N_2048,N_2088);
nand U2562 (N_2562,N_2179,N_1933);
or U2563 (N_2563,N_1879,N_2357);
nor U2564 (N_2564,N_2212,N_2338);
and U2565 (N_2565,N_1836,N_2195);
and U2566 (N_2566,N_2285,N_1903);
xor U2567 (N_2567,N_2374,N_1934);
and U2568 (N_2568,N_2121,N_2305);
and U2569 (N_2569,N_2062,N_1839);
and U2570 (N_2570,N_1904,N_2155);
xor U2571 (N_2571,N_2106,N_1960);
nand U2572 (N_2572,N_1930,N_2239);
or U2573 (N_2573,N_2167,N_1862);
xor U2574 (N_2574,N_2177,N_1844);
nand U2575 (N_2575,N_2371,N_1902);
xnor U2576 (N_2576,N_1911,N_1826);
xor U2577 (N_2577,N_2313,N_2294);
and U2578 (N_2578,N_2136,N_1936);
nand U2579 (N_2579,N_2045,N_2244);
nand U2580 (N_2580,N_1866,N_1806);
or U2581 (N_2581,N_2044,N_1847);
nand U2582 (N_2582,N_2227,N_2335);
and U2583 (N_2583,N_1982,N_2185);
and U2584 (N_2584,N_2031,N_1835);
xor U2585 (N_2585,N_2297,N_2004);
or U2586 (N_2586,N_1927,N_2086);
nor U2587 (N_2587,N_2037,N_2288);
nand U2588 (N_2588,N_2194,N_1981);
nand U2589 (N_2589,N_2343,N_2015);
or U2590 (N_2590,N_1829,N_2072);
nand U2591 (N_2591,N_2395,N_2166);
nor U2592 (N_2592,N_2382,N_2064);
nand U2593 (N_2593,N_2183,N_1857);
or U2594 (N_2594,N_2120,N_2058);
xnor U2595 (N_2595,N_2173,N_2321);
nand U2596 (N_2596,N_2101,N_2079);
or U2597 (N_2597,N_2394,N_2398);
nand U2598 (N_2598,N_1852,N_2223);
xnor U2599 (N_2599,N_1886,N_1874);
nor U2600 (N_2600,N_1884,N_1856);
nor U2601 (N_2601,N_1924,N_2007);
xnor U2602 (N_2602,N_2114,N_2310);
xor U2603 (N_2603,N_2124,N_1954);
and U2604 (N_2604,N_2090,N_1922);
nand U2605 (N_2605,N_1894,N_2369);
xor U2606 (N_2606,N_1977,N_2233);
and U2607 (N_2607,N_2186,N_2147);
or U2608 (N_2608,N_2040,N_2323);
or U2609 (N_2609,N_2207,N_2134);
nand U2610 (N_2610,N_1849,N_2265);
xor U2611 (N_2611,N_1818,N_2308);
xor U2612 (N_2612,N_2143,N_2393);
nor U2613 (N_2613,N_2350,N_2349);
or U2614 (N_2614,N_1946,N_2021);
nor U2615 (N_2615,N_1842,N_2202);
nand U2616 (N_2616,N_2196,N_2282);
or U2617 (N_2617,N_1995,N_2307);
and U2618 (N_2618,N_1915,N_1807);
nand U2619 (N_2619,N_2327,N_2003);
nor U2620 (N_2620,N_2067,N_1993);
nand U2621 (N_2621,N_2337,N_1976);
xnor U2622 (N_2622,N_2116,N_1906);
nor U2623 (N_2623,N_1841,N_1893);
and U2624 (N_2624,N_2026,N_2334);
and U2625 (N_2625,N_2206,N_1897);
and U2626 (N_2626,N_1996,N_2191);
and U2627 (N_2627,N_2256,N_2172);
or U2628 (N_2628,N_1958,N_1812);
nand U2629 (N_2629,N_1883,N_2035);
nand U2630 (N_2630,N_1892,N_2384);
or U2631 (N_2631,N_1887,N_2154);
or U2632 (N_2632,N_1972,N_2215);
xnor U2633 (N_2633,N_1889,N_2385);
nand U2634 (N_2634,N_1882,N_2330);
nand U2635 (N_2635,N_1951,N_2171);
nor U2636 (N_2636,N_1873,N_2153);
and U2637 (N_2637,N_1941,N_1851);
and U2638 (N_2638,N_2331,N_1800);
and U2639 (N_2639,N_1987,N_2261);
nor U2640 (N_2640,N_1885,N_2000);
or U2641 (N_2641,N_2105,N_2089);
xnor U2642 (N_2642,N_1938,N_2033);
and U2643 (N_2643,N_1967,N_1950);
or U2644 (N_2644,N_1983,N_1943);
nand U2645 (N_2645,N_1848,N_2130);
xnor U2646 (N_2646,N_2364,N_2098);
or U2647 (N_2647,N_2314,N_1825);
nor U2648 (N_2648,N_2292,N_1957);
nor U2649 (N_2649,N_2290,N_2054);
nand U2650 (N_2650,N_2075,N_2205);
nor U2651 (N_2651,N_1961,N_2381);
nor U2652 (N_2652,N_2150,N_2198);
nor U2653 (N_2653,N_2148,N_2034);
xnor U2654 (N_2654,N_1956,N_2117);
and U2655 (N_2655,N_2257,N_2110);
or U2656 (N_2656,N_1838,N_2162);
xor U2657 (N_2657,N_1932,N_2164);
nand U2658 (N_2658,N_1992,N_2102);
nand U2659 (N_2659,N_1942,N_2251);
or U2660 (N_2660,N_2049,N_2266);
or U2661 (N_2661,N_1914,N_1869);
and U2662 (N_2662,N_2269,N_1953);
and U2663 (N_2663,N_1832,N_2356);
nand U2664 (N_2664,N_1811,N_2260);
and U2665 (N_2665,N_2258,N_2298);
nand U2666 (N_2666,N_2286,N_1881);
and U2667 (N_2667,N_2083,N_2192);
and U2668 (N_2668,N_2399,N_2199);
xnor U2669 (N_2669,N_2352,N_2041);
nand U2670 (N_2670,N_2050,N_2234);
or U2671 (N_2671,N_2115,N_2077);
nor U2672 (N_2672,N_1801,N_2123);
or U2673 (N_2673,N_2174,N_2068);
and U2674 (N_2674,N_2306,N_2328);
nor U2675 (N_2675,N_2279,N_2267);
nor U2676 (N_2676,N_1867,N_2228);
nand U2677 (N_2677,N_2133,N_2370);
nor U2678 (N_2678,N_2263,N_2264);
nor U2679 (N_2679,N_2014,N_2242);
and U2680 (N_2680,N_2336,N_2152);
nand U2681 (N_2681,N_2039,N_2287);
nor U2682 (N_2682,N_1821,N_2272);
xor U2683 (N_2683,N_2178,N_2012);
xnor U2684 (N_2684,N_2131,N_2052);
nand U2685 (N_2685,N_2097,N_2347);
or U2686 (N_2686,N_2074,N_2240);
and U2687 (N_2687,N_2197,N_2023);
nor U2688 (N_2688,N_2255,N_2238);
nor U2689 (N_2689,N_2022,N_2146);
nor U2690 (N_2690,N_1843,N_2113);
nand U2691 (N_2691,N_1917,N_2158);
nor U2692 (N_2692,N_1816,N_2277);
nand U2693 (N_2693,N_2011,N_2311);
and U2694 (N_2694,N_1840,N_2380);
or U2695 (N_2695,N_2156,N_2273);
or U2696 (N_2696,N_2339,N_2051);
xnor U2697 (N_2697,N_2184,N_1830);
nor U2698 (N_2698,N_2319,N_2203);
nor U2699 (N_2699,N_2209,N_2137);
xnor U2700 (N_2700,N_2052,N_1964);
or U2701 (N_2701,N_2271,N_2051);
nor U2702 (N_2702,N_1823,N_2268);
or U2703 (N_2703,N_2237,N_2396);
xnor U2704 (N_2704,N_2281,N_2038);
nor U2705 (N_2705,N_2335,N_2338);
xnor U2706 (N_2706,N_2329,N_1947);
xor U2707 (N_2707,N_1816,N_2050);
nor U2708 (N_2708,N_1926,N_1948);
nor U2709 (N_2709,N_2012,N_1948);
nand U2710 (N_2710,N_1834,N_1836);
xnor U2711 (N_2711,N_2369,N_1919);
xor U2712 (N_2712,N_2394,N_1887);
nor U2713 (N_2713,N_2042,N_1995);
nor U2714 (N_2714,N_2200,N_2162);
nor U2715 (N_2715,N_1859,N_2314);
or U2716 (N_2716,N_2281,N_1994);
or U2717 (N_2717,N_2014,N_2282);
xor U2718 (N_2718,N_2252,N_2234);
or U2719 (N_2719,N_2318,N_2078);
and U2720 (N_2720,N_2150,N_1901);
nor U2721 (N_2721,N_1838,N_2384);
xor U2722 (N_2722,N_2216,N_1888);
nand U2723 (N_2723,N_2260,N_2237);
and U2724 (N_2724,N_2236,N_2368);
or U2725 (N_2725,N_2019,N_2037);
nor U2726 (N_2726,N_1925,N_1969);
xor U2727 (N_2727,N_1818,N_1806);
and U2728 (N_2728,N_2236,N_2311);
or U2729 (N_2729,N_2214,N_2386);
xnor U2730 (N_2730,N_1876,N_1936);
or U2731 (N_2731,N_2301,N_2277);
nand U2732 (N_2732,N_2001,N_2274);
and U2733 (N_2733,N_2000,N_2134);
xor U2734 (N_2734,N_2366,N_1891);
nor U2735 (N_2735,N_2159,N_2100);
nand U2736 (N_2736,N_2104,N_2085);
and U2737 (N_2737,N_1804,N_2265);
or U2738 (N_2738,N_2275,N_2332);
xnor U2739 (N_2739,N_1848,N_1837);
xnor U2740 (N_2740,N_2027,N_2242);
and U2741 (N_2741,N_2210,N_2165);
and U2742 (N_2742,N_2119,N_2160);
nor U2743 (N_2743,N_2109,N_2100);
nand U2744 (N_2744,N_1956,N_2317);
nor U2745 (N_2745,N_2097,N_1857);
nand U2746 (N_2746,N_2373,N_1986);
nor U2747 (N_2747,N_1886,N_1996);
nand U2748 (N_2748,N_2344,N_2105);
or U2749 (N_2749,N_1801,N_1852);
nand U2750 (N_2750,N_2314,N_1818);
and U2751 (N_2751,N_1902,N_2340);
and U2752 (N_2752,N_2377,N_2171);
and U2753 (N_2753,N_2315,N_2080);
or U2754 (N_2754,N_2205,N_2132);
nand U2755 (N_2755,N_1806,N_1896);
xnor U2756 (N_2756,N_1973,N_2390);
nor U2757 (N_2757,N_2206,N_1988);
or U2758 (N_2758,N_2352,N_1934);
nand U2759 (N_2759,N_2037,N_2026);
or U2760 (N_2760,N_2191,N_1949);
xnor U2761 (N_2761,N_1939,N_2194);
or U2762 (N_2762,N_1820,N_2019);
and U2763 (N_2763,N_2231,N_1917);
or U2764 (N_2764,N_2334,N_1971);
xor U2765 (N_2765,N_1924,N_2394);
xnor U2766 (N_2766,N_2115,N_1855);
nor U2767 (N_2767,N_1852,N_2335);
or U2768 (N_2768,N_1959,N_2116);
and U2769 (N_2769,N_2277,N_1995);
and U2770 (N_2770,N_1929,N_2315);
or U2771 (N_2771,N_2307,N_2187);
nor U2772 (N_2772,N_2163,N_2169);
and U2773 (N_2773,N_2100,N_2144);
nor U2774 (N_2774,N_2298,N_1879);
xor U2775 (N_2775,N_2014,N_2195);
nand U2776 (N_2776,N_2174,N_2262);
or U2777 (N_2777,N_2182,N_2147);
nor U2778 (N_2778,N_2151,N_2018);
and U2779 (N_2779,N_1868,N_1967);
nand U2780 (N_2780,N_2288,N_2345);
nand U2781 (N_2781,N_1994,N_2337);
and U2782 (N_2782,N_1988,N_2219);
or U2783 (N_2783,N_2094,N_2370);
xnor U2784 (N_2784,N_1859,N_1810);
xnor U2785 (N_2785,N_2174,N_1852);
or U2786 (N_2786,N_1825,N_1815);
xor U2787 (N_2787,N_2300,N_1987);
nor U2788 (N_2788,N_2352,N_2208);
nand U2789 (N_2789,N_1984,N_1947);
or U2790 (N_2790,N_1813,N_1903);
or U2791 (N_2791,N_2370,N_2122);
nand U2792 (N_2792,N_2073,N_2299);
nand U2793 (N_2793,N_2236,N_2040);
xor U2794 (N_2794,N_2206,N_1924);
or U2795 (N_2795,N_1869,N_2015);
nand U2796 (N_2796,N_2145,N_2370);
and U2797 (N_2797,N_1931,N_2228);
or U2798 (N_2798,N_1822,N_2161);
xor U2799 (N_2799,N_1805,N_2279);
nor U2800 (N_2800,N_1857,N_2120);
xnor U2801 (N_2801,N_2230,N_2280);
and U2802 (N_2802,N_2128,N_2076);
and U2803 (N_2803,N_2129,N_2061);
xnor U2804 (N_2804,N_1883,N_2188);
and U2805 (N_2805,N_2051,N_2216);
xor U2806 (N_2806,N_1887,N_2111);
or U2807 (N_2807,N_1887,N_2073);
and U2808 (N_2808,N_2307,N_2155);
nand U2809 (N_2809,N_2083,N_2255);
or U2810 (N_2810,N_2079,N_1969);
xor U2811 (N_2811,N_1999,N_1814);
and U2812 (N_2812,N_2137,N_2109);
nor U2813 (N_2813,N_2041,N_2257);
nand U2814 (N_2814,N_1873,N_1928);
and U2815 (N_2815,N_2049,N_2201);
nand U2816 (N_2816,N_2186,N_2124);
nand U2817 (N_2817,N_2297,N_1986);
or U2818 (N_2818,N_1869,N_1938);
nand U2819 (N_2819,N_1875,N_1942);
nor U2820 (N_2820,N_1920,N_2287);
and U2821 (N_2821,N_1991,N_2090);
xnor U2822 (N_2822,N_1861,N_1998);
nor U2823 (N_2823,N_2297,N_2024);
xor U2824 (N_2824,N_2226,N_1858);
nor U2825 (N_2825,N_2170,N_1925);
and U2826 (N_2826,N_2095,N_1939);
xnor U2827 (N_2827,N_2030,N_2169);
and U2828 (N_2828,N_2025,N_1981);
and U2829 (N_2829,N_1916,N_2164);
xnor U2830 (N_2830,N_1989,N_1864);
nor U2831 (N_2831,N_2077,N_2248);
xnor U2832 (N_2832,N_2108,N_2036);
nand U2833 (N_2833,N_2093,N_1932);
xor U2834 (N_2834,N_1958,N_2167);
nor U2835 (N_2835,N_1820,N_2310);
nor U2836 (N_2836,N_2191,N_2094);
nand U2837 (N_2837,N_2086,N_1888);
and U2838 (N_2838,N_1812,N_2199);
nand U2839 (N_2839,N_1882,N_2126);
or U2840 (N_2840,N_2254,N_2221);
or U2841 (N_2841,N_2115,N_1842);
and U2842 (N_2842,N_2017,N_2130);
and U2843 (N_2843,N_2388,N_2011);
nor U2844 (N_2844,N_2351,N_2051);
xor U2845 (N_2845,N_2333,N_2160);
xnor U2846 (N_2846,N_2038,N_2396);
nor U2847 (N_2847,N_2278,N_2330);
or U2848 (N_2848,N_2274,N_1982);
or U2849 (N_2849,N_1947,N_2311);
or U2850 (N_2850,N_2169,N_2053);
and U2851 (N_2851,N_1848,N_1884);
nand U2852 (N_2852,N_2203,N_2045);
nor U2853 (N_2853,N_2089,N_1943);
and U2854 (N_2854,N_1966,N_2047);
xor U2855 (N_2855,N_2225,N_2066);
and U2856 (N_2856,N_1818,N_1946);
xor U2857 (N_2857,N_1816,N_2266);
or U2858 (N_2858,N_2362,N_2386);
nor U2859 (N_2859,N_1859,N_1885);
xnor U2860 (N_2860,N_2395,N_2059);
and U2861 (N_2861,N_1903,N_2099);
xnor U2862 (N_2862,N_2061,N_2256);
and U2863 (N_2863,N_2209,N_2174);
and U2864 (N_2864,N_2066,N_1878);
or U2865 (N_2865,N_2298,N_2315);
nor U2866 (N_2866,N_1934,N_2099);
nand U2867 (N_2867,N_2209,N_2033);
xnor U2868 (N_2868,N_2363,N_1864);
nand U2869 (N_2869,N_1800,N_2073);
and U2870 (N_2870,N_1908,N_2057);
xnor U2871 (N_2871,N_2184,N_1912);
nand U2872 (N_2872,N_1907,N_1894);
nand U2873 (N_2873,N_1951,N_2382);
xor U2874 (N_2874,N_2056,N_1824);
nand U2875 (N_2875,N_2384,N_2197);
xor U2876 (N_2876,N_2207,N_2096);
or U2877 (N_2877,N_1848,N_2212);
nand U2878 (N_2878,N_2371,N_2142);
xor U2879 (N_2879,N_2236,N_2399);
xnor U2880 (N_2880,N_2051,N_1887);
nor U2881 (N_2881,N_2184,N_2132);
and U2882 (N_2882,N_1927,N_2202);
or U2883 (N_2883,N_1928,N_1880);
nor U2884 (N_2884,N_2387,N_2174);
nand U2885 (N_2885,N_2291,N_2359);
and U2886 (N_2886,N_2329,N_2215);
and U2887 (N_2887,N_2212,N_2199);
and U2888 (N_2888,N_2283,N_2263);
nand U2889 (N_2889,N_1952,N_2097);
or U2890 (N_2890,N_2351,N_2377);
nor U2891 (N_2891,N_2201,N_1987);
xnor U2892 (N_2892,N_2241,N_1918);
or U2893 (N_2893,N_2073,N_2374);
nand U2894 (N_2894,N_2083,N_1961);
nand U2895 (N_2895,N_2024,N_2163);
or U2896 (N_2896,N_2100,N_2310);
nand U2897 (N_2897,N_2382,N_2293);
or U2898 (N_2898,N_2385,N_2374);
xnor U2899 (N_2899,N_1872,N_2189);
nand U2900 (N_2900,N_2154,N_1958);
and U2901 (N_2901,N_1939,N_1885);
nand U2902 (N_2902,N_1851,N_1899);
and U2903 (N_2903,N_1945,N_2017);
and U2904 (N_2904,N_2251,N_2040);
nand U2905 (N_2905,N_2031,N_2201);
or U2906 (N_2906,N_2092,N_2324);
or U2907 (N_2907,N_1975,N_1834);
or U2908 (N_2908,N_2150,N_1945);
nand U2909 (N_2909,N_2261,N_1889);
xor U2910 (N_2910,N_2333,N_1935);
nor U2911 (N_2911,N_2295,N_2179);
xor U2912 (N_2912,N_2152,N_1948);
and U2913 (N_2913,N_1982,N_2113);
nand U2914 (N_2914,N_2282,N_1960);
or U2915 (N_2915,N_2327,N_2250);
or U2916 (N_2916,N_2295,N_1813);
nor U2917 (N_2917,N_1804,N_2197);
xnor U2918 (N_2918,N_2162,N_2269);
xnor U2919 (N_2919,N_1968,N_2097);
nand U2920 (N_2920,N_1993,N_2157);
and U2921 (N_2921,N_2389,N_2234);
xnor U2922 (N_2922,N_1827,N_2059);
nand U2923 (N_2923,N_2295,N_1895);
and U2924 (N_2924,N_2082,N_2261);
or U2925 (N_2925,N_2026,N_2324);
and U2926 (N_2926,N_1875,N_1910);
nor U2927 (N_2927,N_2334,N_1857);
nor U2928 (N_2928,N_2301,N_2341);
nand U2929 (N_2929,N_2073,N_2130);
and U2930 (N_2930,N_2398,N_2249);
nor U2931 (N_2931,N_2341,N_1866);
xnor U2932 (N_2932,N_2259,N_2092);
and U2933 (N_2933,N_2032,N_2006);
and U2934 (N_2934,N_2322,N_1950);
nand U2935 (N_2935,N_1856,N_1824);
nand U2936 (N_2936,N_2243,N_2027);
and U2937 (N_2937,N_1819,N_2301);
or U2938 (N_2938,N_1997,N_2382);
xnor U2939 (N_2939,N_2262,N_1888);
and U2940 (N_2940,N_2160,N_2027);
xnor U2941 (N_2941,N_2386,N_1978);
and U2942 (N_2942,N_2330,N_2189);
xnor U2943 (N_2943,N_2244,N_1855);
or U2944 (N_2944,N_2361,N_2144);
xnor U2945 (N_2945,N_2344,N_2251);
xnor U2946 (N_2946,N_2099,N_1898);
nand U2947 (N_2947,N_2367,N_2352);
and U2948 (N_2948,N_1964,N_2135);
nor U2949 (N_2949,N_1852,N_2007);
nand U2950 (N_2950,N_2173,N_2284);
xor U2951 (N_2951,N_2030,N_2349);
nand U2952 (N_2952,N_2162,N_1832);
or U2953 (N_2953,N_1995,N_1801);
or U2954 (N_2954,N_2327,N_1911);
nand U2955 (N_2955,N_2384,N_2155);
nor U2956 (N_2956,N_2329,N_2336);
xor U2957 (N_2957,N_2056,N_1817);
nand U2958 (N_2958,N_2288,N_2147);
xor U2959 (N_2959,N_2135,N_1858);
and U2960 (N_2960,N_1863,N_2133);
xor U2961 (N_2961,N_2147,N_2220);
nand U2962 (N_2962,N_2116,N_2092);
or U2963 (N_2963,N_2279,N_2276);
nand U2964 (N_2964,N_2281,N_2051);
or U2965 (N_2965,N_2346,N_1818);
and U2966 (N_2966,N_1931,N_1946);
and U2967 (N_2967,N_1965,N_2145);
nor U2968 (N_2968,N_2095,N_2288);
nor U2969 (N_2969,N_2066,N_2381);
xnor U2970 (N_2970,N_2376,N_1915);
or U2971 (N_2971,N_2119,N_2075);
nand U2972 (N_2972,N_2200,N_2296);
or U2973 (N_2973,N_2371,N_2385);
xor U2974 (N_2974,N_2177,N_2001);
or U2975 (N_2975,N_2300,N_1961);
xor U2976 (N_2976,N_1889,N_1926);
xnor U2977 (N_2977,N_2350,N_2072);
and U2978 (N_2978,N_2273,N_2059);
and U2979 (N_2979,N_2274,N_2003);
and U2980 (N_2980,N_2356,N_1981);
and U2981 (N_2981,N_2355,N_1842);
xor U2982 (N_2982,N_2020,N_2047);
xnor U2983 (N_2983,N_1993,N_2194);
and U2984 (N_2984,N_2060,N_2293);
xor U2985 (N_2985,N_1892,N_2097);
and U2986 (N_2986,N_2273,N_2243);
nand U2987 (N_2987,N_2106,N_2056);
nor U2988 (N_2988,N_1914,N_2189);
and U2989 (N_2989,N_2193,N_1967);
or U2990 (N_2990,N_2004,N_1862);
and U2991 (N_2991,N_1832,N_1902);
nor U2992 (N_2992,N_2380,N_2398);
nor U2993 (N_2993,N_2229,N_2162);
and U2994 (N_2994,N_2144,N_2009);
and U2995 (N_2995,N_2074,N_1913);
xor U2996 (N_2996,N_2040,N_2348);
and U2997 (N_2997,N_2263,N_2312);
nand U2998 (N_2998,N_2356,N_2208);
nand U2999 (N_2999,N_2311,N_1917);
nand UO_0 (O_0,N_2425,N_2928);
xor UO_1 (O_1,N_2614,N_2704);
nor UO_2 (O_2,N_2635,N_2974);
or UO_3 (O_3,N_2547,N_2806);
nand UO_4 (O_4,N_2636,N_2588);
nand UO_5 (O_5,N_2837,N_2793);
xnor UO_6 (O_6,N_2613,N_2758);
nand UO_7 (O_7,N_2930,N_2722);
nor UO_8 (O_8,N_2553,N_2535);
xor UO_9 (O_9,N_2851,N_2477);
nor UO_10 (O_10,N_2436,N_2498);
nand UO_11 (O_11,N_2988,N_2420);
nand UO_12 (O_12,N_2752,N_2743);
xnor UO_13 (O_13,N_2830,N_2602);
and UO_14 (O_14,N_2737,N_2880);
xnor UO_15 (O_15,N_2802,N_2805);
and UO_16 (O_16,N_2662,N_2583);
or UO_17 (O_17,N_2609,N_2560);
and UO_18 (O_18,N_2824,N_2685);
or UO_19 (O_19,N_2856,N_2652);
xor UO_20 (O_20,N_2571,N_2782);
nor UO_21 (O_21,N_2697,N_2512);
nand UO_22 (O_22,N_2649,N_2688);
and UO_23 (O_23,N_2631,N_2478);
xnor UO_24 (O_24,N_2927,N_2825);
or UO_25 (O_25,N_2965,N_2634);
xnor UO_26 (O_26,N_2770,N_2552);
xor UO_27 (O_27,N_2513,N_2711);
or UO_28 (O_28,N_2980,N_2731);
and UO_29 (O_29,N_2807,N_2754);
xnor UO_30 (O_30,N_2587,N_2959);
or UO_31 (O_31,N_2681,N_2709);
and UO_32 (O_32,N_2895,N_2667);
and UO_33 (O_33,N_2774,N_2616);
nand UO_34 (O_34,N_2505,N_2577);
xor UO_35 (O_35,N_2867,N_2556);
nor UO_36 (O_36,N_2536,N_2475);
and UO_37 (O_37,N_2934,N_2760);
nor UO_38 (O_38,N_2675,N_2818);
nor UO_39 (O_39,N_2444,N_2844);
or UO_40 (O_40,N_2518,N_2708);
nor UO_41 (O_41,N_2692,N_2558);
nand UO_42 (O_42,N_2843,N_2592);
nand UO_43 (O_43,N_2516,N_2911);
or UO_44 (O_44,N_2719,N_2869);
and UO_45 (O_45,N_2773,N_2854);
or UO_46 (O_46,N_2620,N_2463);
nor UO_47 (O_47,N_2501,N_2973);
or UO_48 (O_48,N_2790,N_2985);
nand UO_49 (O_49,N_2705,N_2575);
nand UO_50 (O_50,N_2909,N_2646);
xor UO_51 (O_51,N_2661,N_2725);
xnor UO_52 (O_52,N_2751,N_2544);
nor UO_53 (O_53,N_2918,N_2929);
xor UO_54 (O_54,N_2640,N_2991);
or UO_55 (O_55,N_2455,N_2716);
and UO_56 (O_56,N_2581,N_2739);
nand UO_57 (O_57,N_2561,N_2625);
nand UO_58 (O_58,N_2890,N_2441);
nor UO_59 (O_59,N_2670,N_2559);
and UO_60 (O_60,N_2721,N_2448);
nand UO_61 (O_61,N_2892,N_2611);
or UO_62 (O_62,N_2992,N_2821);
xor UO_63 (O_63,N_2827,N_2914);
or UO_64 (O_64,N_2957,N_2701);
xnor UO_65 (O_65,N_2771,N_2666);
nand UO_66 (O_66,N_2888,N_2971);
and UO_67 (O_67,N_2960,N_2589);
and UO_68 (O_68,N_2462,N_2833);
and UO_69 (O_69,N_2452,N_2781);
xor UO_70 (O_70,N_2522,N_2735);
or UO_71 (O_71,N_2578,N_2794);
and UO_72 (O_72,N_2700,N_2761);
and UO_73 (O_73,N_2698,N_2996);
and UO_74 (O_74,N_2434,N_2894);
nor UO_75 (O_75,N_2972,N_2726);
or UO_76 (O_76,N_2686,N_2415);
nor UO_77 (O_77,N_2526,N_2445);
nor UO_78 (O_78,N_2920,N_2683);
nor UO_79 (O_79,N_2956,N_2846);
xnor UO_80 (O_80,N_2795,N_2473);
nor UO_81 (O_81,N_2669,N_2955);
or UO_82 (O_82,N_2570,N_2476);
nor UO_83 (O_83,N_2595,N_2608);
nand UO_84 (O_84,N_2472,N_2762);
nand UO_85 (O_85,N_2881,N_2426);
or UO_86 (O_86,N_2940,N_2968);
and UO_87 (O_87,N_2878,N_2404);
nor UO_88 (O_88,N_2785,N_2826);
nand UO_89 (O_89,N_2569,N_2599);
nor UO_90 (O_90,N_2995,N_2532);
nand UO_91 (O_91,N_2531,N_2413);
nand UO_92 (O_92,N_2823,N_2598);
or UO_93 (O_93,N_2953,N_2772);
xnor UO_94 (O_94,N_2615,N_2885);
and UO_95 (O_95,N_2811,N_2515);
or UO_96 (O_96,N_2730,N_2554);
or UO_97 (O_97,N_2917,N_2423);
or UO_98 (O_98,N_2769,N_2586);
or UO_99 (O_99,N_2479,N_2813);
xor UO_100 (O_100,N_2766,N_2746);
and UO_101 (O_101,N_2567,N_2873);
nor UO_102 (O_102,N_2411,N_2502);
nor UO_103 (O_103,N_2984,N_2836);
or UO_104 (O_104,N_2506,N_2490);
and UO_105 (O_105,N_2639,N_2677);
xor UO_106 (O_106,N_2779,N_2954);
and UO_107 (O_107,N_2446,N_2563);
or UO_108 (O_108,N_2975,N_2939);
nor UO_109 (O_109,N_2753,N_2948);
and UO_110 (O_110,N_2978,N_2514);
nor UO_111 (O_111,N_2924,N_2495);
nand UO_112 (O_112,N_2799,N_2458);
or UO_113 (O_113,N_2745,N_2842);
xor UO_114 (O_114,N_2907,N_2707);
xnor UO_115 (O_115,N_2864,N_2810);
nor UO_116 (O_116,N_2757,N_2494);
nand UO_117 (O_117,N_2528,N_2576);
xor UO_118 (O_118,N_2933,N_2913);
and UO_119 (O_119,N_2682,N_2428);
and UO_120 (O_120,N_2520,N_2962);
xor UO_121 (O_121,N_2884,N_2606);
nand UO_122 (O_122,N_2470,N_2564);
xnor UO_123 (O_123,N_2565,N_2938);
or UO_124 (O_124,N_2853,N_2672);
and UO_125 (O_125,N_2660,N_2454);
nor UO_126 (O_126,N_2604,N_2926);
nand UO_127 (O_127,N_2936,N_2442);
and UO_128 (O_128,N_2733,N_2819);
and UO_129 (O_129,N_2429,N_2642);
and UO_130 (O_130,N_2488,N_2555);
xor UO_131 (O_131,N_2741,N_2847);
and UO_132 (O_132,N_2724,N_2841);
and UO_133 (O_133,N_2852,N_2944);
nand UO_134 (O_134,N_2814,N_2659);
nand UO_135 (O_135,N_2568,N_2950);
nor UO_136 (O_136,N_2767,N_2879);
xnor UO_137 (O_137,N_2792,N_2902);
or UO_138 (O_138,N_2803,N_2966);
nand UO_139 (O_139,N_2922,N_2783);
and UO_140 (O_140,N_2828,N_2572);
xor UO_141 (O_141,N_2456,N_2776);
xnor UO_142 (O_142,N_2573,N_2712);
nand UO_143 (O_143,N_2937,N_2848);
or UO_144 (O_144,N_2676,N_2644);
nor UO_145 (O_145,N_2416,N_2400);
or UO_146 (O_146,N_2627,N_2775);
nand UO_147 (O_147,N_2401,N_2650);
nand UO_148 (O_148,N_2756,N_2906);
xor UO_149 (O_149,N_2656,N_2808);
nor UO_150 (O_150,N_2874,N_2893);
or UO_151 (O_151,N_2862,N_2622);
xnor UO_152 (O_152,N_2632,N_2983);
and UO_153 (O_153,N_2875,N_2403);
or UO_154 (O_154,N_2469,N_2947);
nand UO_155 (O_155,N_2863,N_2877);
and UO_156 (O_156,N_2464,N_2859);
and UO_157 (O_157,N_2418,N_2804);
nand UO_158 (O_158,N_2921,N_2839);
or UO_159 (O_159,N_2500,N_2607);
or UO_160 (O_160,N_2925,N_2527);
nor UO_161 (O_161,N_2543,N_2480);
nand UO_162 (O_162,N_2524,N_2503);
xor UO_163 (O_163,N_2610,N_2507);
and UO_164 (O_164,N_2896,N_2858);
nand UO_165 (O_165,N_2800,N_2633);
and UO_166 (O_166,N_2409,N_2549);
nand UO_167 (O_167,N_2812,N_2597);
nand UO_168 (O_168,N_2433,N_2798);
and UO_169 (O_169,N_2424,N_2637);
xnor UO_170 (O_170,N_2489,N_2601);
nand UO_171 (O_171,N_2687,N_2579);
nor UO_172 (O_172,N_2990,N_2816);
nand UO_173 (O_173,N_2900,N_2663);
nor UO_174 (O_174,N_2986,N_2923);
xnor UO_175 (O_175,N_2786,N_2414);
and UO_176 (O_176,N_2829,N_2749);
nor UO_177 (O_177,N_2529,N_2694);
nand UO_178 (O_178,N_2468,N_2600);
or UO_179 (O_179,N_2887,N_2467);
xnor UO_180 (O_180,N_2497,N_2658);
nand UO_181 (O_181,N_2747,N_2419);
nand UO_182 (O_182,N_2742,N_2443);
xnor UO_183 (O_183,N_2860,N_2897);
nand UO_184 (O_184,N_2696,N_2715);
or UO_185 (O_185,N_2801,N_2643);
nand UO_186 (O_186,N_2402,N_2674);
xor UO_187 (O_187,N_2417,N_2693);
nor UO_188 (O_188,N_2673,N_2574);
or UO_189 (O_189,N_2484,N_2540);
or UO_190 (O_190,N_2872,N_2439);
nand UO_191 (O_191,N_2407,N_2450);
or UO_192 (O_192,N_2967,N_2777);
nand UO_193 (O_193,N_2457,N_2408);
nor UO_194 (O_194,N_2509,N_2738);
and UO_195 (O_195,N_2499,N_2908);
nand UO_196 (O_196,N_2734,N_2870);
and UO_197 (O_197,N_2732,N_2679);
xor UO_198 (O_198,N_2551,N_2998);
nor UO_199 (O_199,N_2740,N_2621);
and UO_200 (O_200,N_2657,N_2580);
or UO_201 (O_201,N_2618,N_2727);
xor UO_202 (O_202,N_2504,N_2822);
nand UO_203 (O_203,N_2412,N_2593);
or UO_204 (O_204,N_2750,N_2710);
nor UO_205 (O_205,N_2461,N_2427);
or UO_206 (O_206,N_2630,N_2493);
or UO_207 (O_207,N_2713,N_2788);
nor UO_208 (O_208,N_2511,N_2849);
nor UO_209 (O_209,N_2706,N_2838);
xnor UO_210 (O_210,N_2834,N_2942);
nand UO_211 (O_211,N_2951,N_2459);
or UO_212 (O_212,N_2865,N_2820);
and UO_213 (O_213,N_2945,N_2961);
xor UO_214 (O_214,N_2728,N_2997);
xnor UO_215 (O_215,N_2958,N_2703);
xnor UO_216 (O_216,N_2508,N_2562);
nand UO_217 (O_217,N_2530,N_2964);
nor UO_218 (O_218,N_2465,N_2868);
and UO_219 (O_219,N_2437,N_2979);
or UO_220 (O_220,N_2678,N_2585);
xnor UO_221 (O_221,N_2596,N_2612);
xor UO_222 (O_222,N_2695,N_2915);
xnor UO_223 (O_223,N_2410,N_2590);
xor UO_224 (O_224,N_2898,N_2668);
nand UO_225 (O_225,N_2582,N_2717);
xor UO_226 (O_226,N_2482,N_2691);
nand UO_227 (O_227,N_2970,N_2748);
or UO_228 (O_228,N_2671,N_2491);
and UO_229 (O_229,N_2545,N_2720);
xnor UO_230 (O_230,N_2645,N_2949);
xnor UO_231 (O_231,N_2431,N_2541);
and UO_232 (O_232,N_2629,N_2550);
and UO_233 (O_233,N_2519,N_2664);
xor UO_234 (O_234,N_2438,N_2421);
and UO_235 (O_235,N_2977,N_2689);
and UO_236 (O_236,N_2537,N_2916);
or UO_237 (O_237,N_2594,N_2603);
nor UO_238 (O_238,N_2883,N_2755);
or UO_239 (O_239,N_2729,N_2989);
and UO_240 (O_240,N_2882,N_2487);
xnor UO_241 (O_241,N_2886,N_2523);
nand UO_242 (O_242,N_2647,N_2447);
and UO_243 (O_243,N_2866,N_2993);
nor UO_244 (O_244,N_2486,N_2744);
and UO_245 (O_245,N_2542,N_2901);
or UO_246 (O_246,N_2903,N_2517);
and UO_247 (O_247,N_2876,N_2778);
nor UO_248 (O_248,N_2406,N_2440);
or UO_249 (O_249,N_2525,N_2453);
or UO_250 (O_250,N_2605,N_2699);
and UO_251 (O_251,N_2904,N_2976);
nor UO_252 (O_252,N_2449,N_2655);
nor UO_253 (O_253,N_2815,N_2943);
xor UO_254 (O_254,N_2809,N_2474);
nor UO_255 (O_255,N_2931,N_2764);
nand UO_256 (O_256,N_2641,N_2768);
nand UO_257 (O_257,N_2763,N_2905);
and UO_258 (O_258,N_2619,N_2432);
nand UO_259 (O_259,N_2591,N_2485);
xor UO_260 (O_260,N_2665,N_2584);
nand UO_261 (O_261,N_2451,N_2999);
xnor UO_262 (O_262,N_2981,N_2483);
or UO_263 (O_263,N_2496,N_2684);
and UO_264 (O_264,N_2702,N_2736);
nor UO_265 (O_265,N_2405,N_2946);
xnor UO_266 (O_266,N_2987,N_2835);
nand UO_267 (O_267,N_2935,N_2680);
xor UO_268 (O_268,N_2963,N_2850);
nand UO_269 (O_269,N_2994,N_2617);
or UO_270 (O_270,N_2952,N_2857);
nand UO_271 (O_271,N_2831,N_2628);
nor UO_272 (O_272,N_2919,N_2638);
nand UO_273 (O_273,N_2714,N_2521);
and UO_274 (O_274,N_2466,N_2780);
xor UO_275 (O_275,N_2623,N_2789);
and UO_276 (O_276,N_2891,N_2651);
nor UO_277 (O_277,N_2969,N_2941);
and UO_278 (O_278,N_2435,N_2787);
xor UO_279 (O_279,N_2899,N_2653);
nor UO_280 (O_280,N_2982,N_2626);
and UO_281 (O_281,N_2832,N_2534);
or UO_282 (O_282,N_2538,N_2861);
or UO_283 (O_283,N_2654,N_2460);
and UO_284 (O_284,N_2539,N_2422);
and UO_285 (O_285,N_2791,N_2566);
nand UO_286 (O_286,N_2510,N_2889);
nand UO_287 (O_287,N_2759,N_2765);
or UO_288 (O_288,N_2855,N_2481);
or UO_289 (O_289,N_2557,N_2546);
xor UO_290 (O_290,N_2723,N_2533);
nand UO_291 (O_291,N_2797,N_2624);
nand UO_292 (O_292,N_2690,N_2840);
and UO_293 (O_293,N_2932,N_2912);
nor UO_294 (O_294,N_2910,N_2548);
xnor UO_295 (O_295,N_2784,N_2492);
nand UO_296 (O_296,N_2817,N_2471);
nor UO_297 (O_297,N_2648,N_2796);
nand UO_298 (O_298,N_2430,N_2845);
xnor UO_299 (O_299,N_2718,N_2871);
and UO_300 (O_300,N_2561,N_2409);
xor UO_301 (O_301,N_2948,N_2831);
nor UO_302 (O_302,N_2430,N_2895);
or UO_303 (O_303,N_2714,N_2527);
nand UO_304 (O_304,N_2568,N_2687);
nand UO_305 (O_305,N_2799,N_2976);
or UO_306 (O_306,N_2792,N_2767);
and UO_307 (O_307,N_2559,N_2557);
xor UO_308 (O_308,N_2666,N_2452);
and UO_309 (O_309,N_2735,N_2743);
and UO_310 (O_310,N_2401,N_2446);
xnor UO_311 (O_311,N_2935,N_2420);
xor UO_312 (O_312,N_2828,N_2669);
and UO_313 (O_313,N_2786,N_2811);
and UO_314 (O_314,N_2863,N_2770);
or UO_315 (O_315,N_2805,N_2430);
nor UO_316 (O_316,N_2795,N_2645);
or UO_317 (O_317,N_2415,N_2601);
and UO_318 (O_318,N_2954,N_2433);
nor UO_319 (O_319,N_2577,N_2885);
xor UO_320 (O_320,N_2454,N_2418);
nand UO_321 (O_321,N_2444,N_2792);
and UO_322 (O_322,N_2698,N_2911);
nand UO_323 (O_323,N_2945,N_2718);
nor UO_324 (O_324,N_2647,N_2542);
nor UO_325 (O_325,N_2588,N_2567);
or UO_326 (O_326,N_2474,N_2977);
and UO_327 (O_327,N_2885,N_2738);
nor UO_328 (O_328,N_2400,N_2432);
xnor UO_329 (O_329,N_2615,N_2614);
xor UO_330 (O_330,N_2639,N_2457);
and UO_331 (O_331,N_2746,N_2628);
or UO_332 (O_332,N_2838,N_2911);
and UO_333 (O_333,N_2450,N_2934);
or UO_334 (O_334,N_2768,N_2404);
nor UO_335 (O_335,N_2833,N_2996);
nand UO_336 (O_336,N_2405,N_2422);
and UO_337 (O_337,N_2617,N_2559);
and UO_338 (O_338,N_2531,N_2450);
nand UO_339 (O_339,N_2618,N_2678);
nand UO_340 (O_340,N_2592,N_2898);
and UO_341 (O_341,N_2892,N_2563);
and UO_342 (O_342,N_2859,N_2664);
nor UO_343 (O_343,N_2804,N_2932);
xor UO_344 (O_344,N_2993,N_2659);
xor UO_345 (O_345,N_2404,N_2434);
and UO_346 (O_346,N_2606,N_2766);
or UO_347 (O_347,N_2933,N_2416);
xor UO_348 (O_348,N_2461,N_2878);
nand UO_349 (O_349,N_2904,N_2723);
and UO_350 (O_350,N_2426,N_2731);
and UO_351 (O_351,N_2826,N_2842);
and UO_352 (O_352,N_2749,N_2712);
or UO_353 (O_353,N_2757,N_2907);
or UO_354 (O_354,N_2965,N_2955);
or UO_355 (O_355,N_2670,N_2686);
or UO_356 (O_356,N_2666,N_2749);
or UO_357 (O_357,N_2600,N_2509);
xnor UO_358 (O_358,N_2902,N_2933);
and UO_359 (O_359,N_2404,N_2972);
and UO_360 (O_360,N_2699,N_2493);
nand UO_361 (O_361,N_2650,N_2783);
xnor UO_362 (O_362,N_2557,N_2416);
nor UO_363 (O_363,N_2707,N_2706);
or UO_364 (O_364,N_2655,N_2822);
and UO_365 (O_365,N_2795,N_2768);
xnor UO_366 (O_366,N_2938,N_2579);
xnor UO_367 (O_367,N_2865,N_2461);
or UO_368 (O_368,N_2830,N_2763);
or UO_369 (O_369,N_2767,N_2954);
nor UO_370 (O_370,N_2602,N_2403);
and UO_371 (O_371,N_2810,N_2736);
xor UO_372 (O_372,N_2810,N_2759);
or UO_373 (O_373,N_2546,N_2718);
nor UO_374 (O_374,N_2848,N_2941);
xnor UO_375 (O_375,N_2953,N_2653);
xnor UO_376 (O_376,N_2700,N_2970);
nand UO_377 (O_377,N_2809,N_2939);
xnor UO_378 (O_378,N_2893,N_2919);
nor UO_379 (O_379,N_2848,N_2833);
xnor UO_380 (O_380,N_2709,N_2963);
xor UO_381 (O_381,N_2926,N_2814);
nor UO_382 (O_382,N_2935,N_2570);
nand UO_383 (O_383,N_2986,N_2511);
nor UO_384 (O_384,N_2749,N_2583);
and UO_385 (O_385,N_2689,N_2443);
xnor UO_386 (O_386,N_2477,N_2777);
or UO_387 (O_387,N_2763,N_2694);
nand UO_388 (O_388,N_2446,N_2816);
and UO_389 (O_389,N_2613,N_2517);
or UO_390 (O_390,N_2467,N_2491);
nor UO_391 (O_391,N_2618,N_2486);
xnor UO_392 (O_392,N_2604,N_2828);
and UO_393 (O_393,N_2459,N_2500);
nor UO_394 (O_394,N_2742,N_2696);
or UO_395 (O_395,N_2402,N_2719);
nand UO_396 (O_396,N_2850,N_2843);
nand UO_397 (O_397,N_2402,N_2423);
nand UO_398 (O_398,N_2639,N_2436);
or UO_399 (O_399,N_2810,N_2499);
xor UO_400 (O_400,N_2977,N_2639);
xor UO_401 (O_401,N_2502,N_2728);
or UO_402 (O_402,N_2544,N_2672);
or UO_403 (O_403,N_2823,N_2721);
and UO_404 (O_404,N_2661,N_2458);
or UO_405 (O_405,N_2951,N_2919);
xnor UO_406 (O_406,N_2984,N_2593);
nand UO_407 (O_407,N_2711,N_2575);
xnor UO_408 (O_408,N_2873,N_2808);
nor UO_409 (O_409,N_2803,N_2633);
nor UO_410 (O_410,N_2511,N_2889);
nand UO_411 (O_411,N_2669,N_2451);
or UO_412 (O_412,N_2816,N_2979);
nor UO_413 (O_413,N_2467,N_2601);
and UO_414 (O_414,N_2934,N_2689);
nor UO_415 (O_415,N_2974,N_2675);
nor UO_416 (O_416,N_2662,N_2822);
or UO_417 (O_417,N_2988,N_2604);
nor UO_418 (O_418,N_2529,N_2759);
nor UO_419 (O_419,N_2446,N_2627);
xor UO_420 (O_420,N_2605,N_2594);
or UO_421 (O_421,N_2936,N_2842);
nor UO_422 (O_422,N_2496,N_2670);
or UO_423 (O_423,N_2631,N_2571);
nor UO_424 (O_424,N_2577,N_2751);
and UO_425 (O_425,N_2466,N_2417);
nand UO_426 (O_426,N_2952,N_2592);
nand UO_427 (O_427,N_2680,N_2442);
nand UO_428 (O_428,N_2501,N_2933);
or UO_429 (O_429,N_2515,N_2539);
nand UO_430 (O_430,N_2800,N_2915);
xor UO_431 (O_431,N_2614,N_2765);
nor UO_432 (O_432,N_2963,N_2976);
or UO_433 (O_433,N_2949,N_2771);
nand UO_434 (O_434,N_2984,N_2988);
nand UO_435 (O_435,N_2947,N_2728);
nor UO_436 (O_436,N_2428,N_2567);
or UO_437 (O_437,N_2549,N_2515);
nor UO_438 (O_438,N_2504,N_2541);
nor UO_439 (O_439,N_2746,N_2902);
or UO_440 (O_440,N_2889,N_2816);
and UO_441 (O_441,N_2497,N_2548);
nor UO_442 (O_442,N_2855,N_2535);
and UO_443 (O_443,N_2980,N_2897);
or UO_444 (O_444,N_2933,N_2818);
or UO_445 (O_445,N_2976,N_2686);
xor UO_446 (O_446,N_2719,N_2598);
nand UO_447 (O_447,N_2958,N_2791);
or UO_448 (O_448,N_2406,N_2567);
or UO_449 (O_449,N_2913,N_2660);
nor UO_450 (O_450,N_2635,N_2580);
nor UO_451 (O_451,N_2493,N_2422);
nor UO_452 (O_452,N_2722,N_2832);
nor UO_453 (O_453,N_2918,N_2401);
nor UO_454 (O_454,N_2996,N_2661);
and UO_455 (O_455,N_2877,N_2967);
and UO_456 (O_456,N_2509,N_2766);
nor UO_457 (O_457,N_2847,N_2904);
xor UO_458 (O_458,N_2694,N_2606);
and UO_459 (O_459,N_2950,N_2496);
or UO_460 (O_460,N_2760,N_2528);
nand UO_461 (O_461,N_2943,N_2848);
or UO_462 (O_462,N_2700,N_2671);
xor UO_463 (O_463,N_2763,N_2945);
xnor UO_464 (O_464,N_2740,N_2840);
nor UO_465 (O_465,N_2439,N_2991);
nor UO_466 (O_466,N_2814,N_2872);
xor UO_467 (O_467,N_2683,N_2526);
nand UO_468 (O_468,N_2948,N_2604);
and UO_469 (O_469,N_2572,N_2496);
xnor UO_470 (O_470,N_2997,N_2614);
and UO_471 (O_471,N_2666,N_2454);
xor UO_472 (O_472,N_2651,N_2473);
and UO_473 (O_473,N_2494,N_2547);
and UO_474 (O_474,N_2648,N_2977);
xnor UO_475 (O_475,N_2542,N_2638);
nand UO_476 (O_476,N_2951,N_2848);
nor UO_477 (O_477,N_2598,N_2521);
nor UO_478 (O_478,N_2560,N_2887);
or UO_479 (O_479,N_2577,N_2410);
nor UO_480 (O_480,N_2412,N_2953);
nor UO_481 (O_481,N_2765,N_2917);
nand UO_482 (O_482,N_2868,N_2601);
xnor UO_483 (O_483,N_2662,N_2684);
nor UO_484 (O_484,N_2685,N_2605);
nand UO_485 (O_485,N_2892,N_2738);
xnor UO_486 (O_486,N_2779,N_2999);
or UO_487 (O_487,N_2472,N_2601);
nor UO_488 (O_488,N_2491,N_2781);
nand UO_489 (O_489,N_2751,N_2443);
and UO_490 (O_490,N_2925,N_2711);
or UO_491 (O_491,N_2904,N_2630);
nand UO_492 (O_492,N_2732,N_2565);
and UO_493 (O_493,N_2481,N_2572);
or UO_494 (O_494,N_2426,N_2983);
or UO_495 (O_495,N_2775,N_2745);
xnor UO_496 (O_496,N_2991,N_2428);
xnor UO_497 (O_497,N_2474,N_2591);
and UO_498 (O_498,N_2820,N_2967);
nand UO_499 (O_499,N_2863,N_2586);
endmodule