module basic_3000_30000_3500_15_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2742,In_2709);
or U1 (N_1,In_1311,In_1858);
nor U2 (N_2,In_2365,In_482);
and U3 (N_3,In_2129,In_2763);
nor U4 (N_4,In_2225,In_2432);
nor U5 (N_5,In_1652,In_2778);
and U6 (N_6,In_1116,In_2822);
nor U7 (N_7,In_2592,In_1004);
nand U8 (N_8,In_39,In_1265);
nor U9 (N_9,In_442,In_381);
or U10 (N_10,In_2274,In_1670);
xnor U11 (N_11,In_2916,In_171);
or U12 (N_12,In_887,In_2550);
xnor U13 (N_13,In_2114,In_2152);
nor U14 (N_14,In_684,In_450);
xor U15 (N_15,In_704,In_2044);
and U16 (N_16,In_2836,In_1573);
nor U17 (N_17,In_844,In_1275);
nor U18 (N_18,In_2919,In_1182);
and U19 (N_19,In_1046,In_2173);
nor U20 (N_20,In_2459,In_837);
or U21 (N_21,In_2242,In_106);
xnor U22 (N_22,In_2257,In_2039);
xor U23 (N_23,In_1944,In_2259);
and U24 (N_24,In_1132,In_1536);
or U25 (N_25,In_2815,In_453);
xor U26 (N_26,In_307,In_937);
nand U27 (N_27,In_1624,In_2617);
xnor U28 (N_28,In_1263,In_2800);
and U29 (N_29,In_170,In_361);
or U30 (N_30,In_695,In_2794);
nor U31 (N_31,In_1135,In_510);
and U32 (N_32,In_1916,In_2947);
xor U33 (N_33,In_2549,In_2726);
or U34 (N_34,In_1097,In_1225);
nand U35 (N_35,In_920,In_2767);
or U36 (N_36,In_479,In_2308);
nand U37 (N_37,In_2123,In_2573);
nand U38 (N_38,In_228,In_444);
xnor U39 (N_39,In_2803,In_2509);
nor U40 (N_40,In_260,In_2854);
xor U41 (N_41,In_600,In_817);
xnor U42 (N_42,In_2807,In_338);
xnor U43 (N_43,In_2570,In_185);
nand U44 (N_44,In_1114,In_498);
or U45 (N_45,In_1505,In_878);
or U46 (N_46,In_2302,In_1098);
nand U47 (N_47,In_1503,In_1433);
or U48 (N_48,In_1615,In_733);
nand U49 (N_49,In_2915,In_757);
nand U50 (N_50,In_980,In_1320);
nand U51 (N_51,In_1224,In_590);
nand U52 (N_52,In_1024,In_2736);
or U53 (N_53,In_2166,In_2183);
and U54 (N_54,In_693,In_2994);
and U55 (N_55,In_2099,In_2370);
and U56 (N_56,In_1887,In_2018);
nor U57 (N_57,In_1565,In_2766);
xor U58 (N_58,In_1129,In_1680);
or U59 (N_59,In_666,In_364);
nor U60 (N_60,In_2126,In_720);
xnor U61 (N_61,In_233,In_2989);
xnor U62 (N_62,In_2619,In_2175);
nor U63 (N_63,In_2250,In_1165);
or U64 (N_64,In_212,In_858);
or U65 (N_65,In_2016,In_280);
nor U66 (N_66,In_794,In_1648);
and U67 (N_67,In_2507,In_595);
and U68 (N_68,In_682,In_490);
and U69 (N_69,In_1429,In_1612);
or U70 (N_70,In_1830,In_759);
nor U71 (N_71,In_2019,In_2817);
nand U72 (N_72,In_2725,In_2596);
nand U73 (N_73,In_2160,In_2150);
nand U74 (N_74,In_2377,In_1529);
nand U75 (N_75,In_1507,In_2856);
nand U76 (N_76,In_1253,In_897);
and U77 (N_77,In_2329,In_1439);
xor U78 (N_78,In_321,In_82);
xor U79 (N_79,In_2748,In_2829);
or U80 (N_80,In_612,In_1298);
and U81 (N_81,In_1806,In_1119);
and U82 (N_82,In_2482,In_2546);
or U83 (N_83,In_1818,In_300);
nor U84 (N_84,In_1942,In_2988);
nand U85 (N_85,In_1519,In_1362);
and U86 (N_86,In_1158,In_2946);
or U87 (N_87,In_964,In_1594);
or U88 (N_88,In_2936,In_2973);
nor U89 (N_89,In_1658,In_2091);
xor U90 (N_90,In_545,In_1629);
nand U91 (N_91,In_1662,In_1401);
and U92 (N_92,In_972,In_2562);
nor U93 (N_93,In_1866,In_2314);
nand U94 (N_94,In_353,In_1299);
xor U95 (N_95,In_2035,In_1956);
xor U96 (N_96,In_1560,In_2072);
nor U97 (N_97,In_77,In_830);
or U98 (N_98,In_2650,In_81);
nand U99 (N_99,In_445,In_2640);
xor U100 (N_100,In_2900,In_1886);
or U101 (N_101,In_1077,In_588);
or U102 (N_102,In_2880,In_2122);
or U103 (N_103,In_1581,In_2034);
or U104 (N_104,In_274,In_1240);
nor U105 (N_105,In_1894,In_2013);
nand U106 (N_106,In_134,In_2764);
and U107 (N_107,In_1738,In_2165);
xnor U108 (N_108,In_2738,In_121);
or U109 (N_109,In_2228,In_1504);
and U110 (N_110,In_1526,In_2474);
and U111 (N_111,In_304,In_857);
xnor U112 (N_112,In_2073,In_107);
xor U113 (N_113,In_213,In_1788);
xor U114 (N_114,In_2821,In_2442);
nand U115 (N_115,In_2323,In_2876);
nor U116 (N_116,In_494,In_2426);
nor U117 (N_117,In_509,In_1909);
nor U118 (N_118,In_1527,In_644);
and U119 (N_119,In_2361,In_1235);
xnor U120 (N_120,In_614,In_1996);
and U121 (N_121,In_2059,In_1405);
nor U122 (N_122,In_72,In_68);
or U123 (N_123,In_2548,In_615);
nor U124 (N_124,In_2326,In_1568);
xor U125 (N_125,In_2237,In_1248);
xor U126 (N_126,In_1793,In_2369);
nor U127 (N_127,In_2222,In_2655);
or U128 (N_128,In_489,In_1141);
nor U129 (N_129,In_1923,In_492);
nor U130 (N_130,In_1451,In_696);
nand U131 (N_131,In_895,In_192);
nand U132 (N_132,In_2454,In_2083);
nand U133 (N_133,In_1705,In_366);
nor U134 (N_134,In_1908,In_1812);
nand U135 (N_135,In_15,In_2608);
xnor U136 (N_136,In_423,In_252);
and U137 (N_137,In_2098,In_2568);
nand U138 (N_138,In_815,In_1930);
or U139 (N_139,In_2848,In_1206);
and U140 (N_140,In_2158,In_853);
xor U141 (N_141,In_825,In_385);
nand U142 (N_142,In_1399,In_2477);
and U143 (N_143,In_784,In_390);
xnor U144 (N_144,In_698,In_2125);
and U145 (N_145,In_318,In_1359);
nor U146 (N_146,In_1563,In_149);
and U147 (N_147,In_1000,In_2851);
and U148 (N_148,In_1307,In_1369);
and U149 (N_149,In_2344,In_2716);
xor U150 (N_150,In_1234,In_427);
xnor U151 (N_151,In_1659,In_380);
or U152 (N_152,In_2681,In_652);
nand U153 (N_153,In_1875,In_1572);
or U154 (N_154,In_2127,In_1628);
xor U155 (N_155,In_675,In_363);
nor U156 (N_156,In_2440,In_2676);
and U157 (N_157,In_2462,In_2627);
nor U158 (N_158,In_276,In_9);
nor U159 (N_159,In_371,In_2008);
nand U160 (N_160,In_1425,In_1569);
and U161 (N_161,In_2248,In_1796);
nor U162 (N_162,In_1809,In_502);
nand U163 (N_163,In_1692,In_1543);
nor U164 (N_164,In_351,In_557);
nand U165 (N_165,In_443,In_995);
nor U166 (N_166,In_1623,In_2980);
xnor U167 (N_167,In_1846,In_1105);
or U168 (N_168,In_2423,In_2061);
and U169 (N_169,In_629,In_2223);
nor U170 (N_170,In_102,In_616);
nor U171 (N_171,In_2296,In_1333);
nor U172 (N_172,In_246,In_1213);
nand U173 (N_173,In_796,In_2428);
xor U174 (N_174,In_2969,In_1103);
nor U175 (N_175,In_250,In_1361);
nand U176 (N_176,In_866,In_2322);
nand U177 (N_177,In_2054,In_2720);
xor U178 (N_178,In_2846,In_2868);
nor U179 (N_179,In_219,In_2399);
nand U180 (N_180,In_352,In_1233);
or U181 (N_181,In_648,In_840);
nand U182 (N_182,In_1990,In_1166);
xor U183 (N_183,In_864,In_1099);
xor U184 (N_184,In_926,In_2917);
nand U185 (N_185,In_2106,In_1920);
nor U186 (N_186,In_922,In_1445);
nor U187 (N_187,In_1063,In_1372);
and U188 (N_188,In_1202,In_969);
nor U189 (N_189,In_2712,In_2699);
nand U190 (N_190,In_2170,In_67);
nor U191 (N_191,In_2662,In_2384);
or U192 (N_192,In_1833,In_162);
nor U193 (N_193,In_2189,In_2710);
or U194 (N_194,In_663,In_2045);
and U195 (N_195,In_2508,In_2262);
nor U196 (N_196,In_2398,In_347);
xor U197 (N_197,In_1417,In_235);
xor U198 (N_198,In_767,In_810);
and U199 (N_199,In_310,In_1477);
and U200 (N_200,In_2280,In_2372);
xor U201 (N_201,In_789,In_271);
nand U202 (N_202,In_1021,In_284);
or U203 (N_203,In_2694,In_683);
or U204 (N_204,In_195,In_1023);
xnor U205 (N_205,In_2700,In_2648);
or U206 (N_206,In_2221,In_1610);
nand U207 (N_207,In_2678,In_2882);
nand U208 (N_208,In_2185,In_2258);
xor U209 (N_209,In_8,In_916);
xnor U210 (N_210,In_1330,In_2254);
nand U211 (N_211,In_1819,In_1229);
or U212 (N_212,In_2719,In_1939);
or U213 (N_213,In_947,In_326);
and U214 (N_214,In_92,In_591);
xor U215 (N_215,In_1962,In_2537);
or U216 (N_216,In_737,In_2362);
nand U217 (N_217,In_2793,In_524);
or U218 (N_218,In_1285,In_1409);
nand U219 (N_219,In_2132,In_2538);
nand U220 (N_220,In_440,In_2058);
or U221 (N_221,In_1602,In_475);
xor U222 (N_222,In_1423,In_362);
nand U223 (N_223,In_1332,In_254);
nor U224 (N_224,In_691,In_2360);
nand U225 (N_225,In_2465,In_1597);
nor U226 (N_226,In_1755,In_2757);
or U227 (N_227,In_1885,In_1955);
or U228 (N_228,In_1431,In_2139);
xor U229 (N_229,In_2151,In_738);
and U230 (N_230,In_1384,In_1749);
xnor U231 (N_231,In_151,In_1513);
nand U232 (N_232,In_2415,In_177);
xnor U233 (N_233,In_473,In_1901);
nand U234 (N_234,In_1559,In_431);
or U235 (N_235,In_278,In_838);
nand U236 (N_236,In_286,In_2288);
xnor U237 (N_237,In_2871,In_236);
and U238 (N_238,In_2079,In_376);
or U239 (N_239,In_1247,In_37);
xor U240 (N_240,In_807,In_2553);
and U241 (N_241,In_1344,In_323);
and U242 (N_242,In_1546,In_1252);
nor U243 (N_243,In_2046,In_1821);
nor U244 (N_244,In_716,In_273);
nor U245 (N_245,In_2481,In_1036);
xnor U246 (N_246,In_802,In_90);
or U247 (N_247,In_1801,In_205);
xor U248 (N_248,In_1254,In_1470);
or U249 (N_249,In_2751,In_899);
nor U250 (N_250,In_646,In_2557);
nand U251 (N_251,In_1111,In_2765);
nor U252 (N_252,In_2999,In_2480);
xor U253 (N_253,In_435,In_2402);
xnor U254 (N_254,In_2930,In_1989);
nand U255 (N_255,In_499,In_1030);
nor U256 (N_256,In_1317,In_1269);
or U257 (N_257,In_468,In_4);
nand U258 (N_258,In_2172,In_1195);
or U259 (N_259,In_2450,In_199);
or U260 (N_260,In_1140,In_1732);
nand U261 (N_261,In_2976,In_670);
nand U262 (N_262,In_2804,In_1981);
and U263 (N_263,In_2032,In_110);
nand U264 (N_264,In_2746,In_1701);
or U265 (N_265,In_950,In_2923);
or U266 (N_266,In_214,In_2327);
and U267 (N_267,In_2485,In_2967);
or U268 (N_268,In_230,In_2138);
and U269 (N_269,In_1204,In_143);
nor U270 (N_270,In_181,In_2893);
or U271 (N_271,In_350,In_2914);
or U272 (N_272,In_239,In_1758);
xnor U273 (N_273,In_21,In_2001);
or U274 (N_274,In_2587,In_2241);
and U275 (N_275,In_2230,In_2203);
or U276 (N_276,In_30,In_1667);
or U277 (N_277,In_2554,In_2526);
nor U278 (N_278,In_1056,In_1378);
or U279 (N_279,In_229,In_1906);
xor U280 (N_280,In_888,In_2272);
nand U281 (N_281,In_579,In_1294);
nand U282 (N_282,In_2421,In_823);
nand U283 (N_283,In_681,In_983);
or U284 (N_284,In_240,In_1003);
nand U285 (N_285,In_1697,In_661);
and U286 (N_286,In_2156,In_534);
xnor U287 (N_287,In_1198,In_799);
or U288 (N_288,In_1197,In_2981);
nand U289 (N_289,In_2847,In_1574);
nand U290 (N_290,In_1131,In_1139);
nand U291 (N_291,In_1205,In_2453);
and U292 (N_292,In_2962,In_2888);
nand U293 (N_293,In_703,In_1595);
xor U294 (N_294,In_1743,In_2735);
or U295 (N_295,In_1452,In_2469);
nor U296 (N_296,In_2569,In_2333);
or U297 (N_297,In_505,In_126);
nand U298 (N_298,In_1741,In_848);
xnor U299 (N_299,In_2579,In_624);
or U300 (N_300,In_1564,In_256);
and U301 (N_301,In_593,In_1357);
and U302 (N_302,In_2779,In_415);
or U303 (N_303,In_1426,In_2612);
nor U304 (N_304,In_2464,In_1538);
xor U305 (N_305,In_1408,In_2993);
or U306 (N_306,In_1406,In_464);
nor U307 (N_307,In_1193,In_583);
nand U308 (N_308,In_1292,In_798);
or U309 (N_309,In_2721,In_605);
or U310 (N_310,In_2996,In_2795);
or U311 (N_311,In_989,In_2238);
or U312 (N_312,In_2468,In_2202);
xnor U313 (N_313,In_2910,In_748);
xor U314 (N_314,In_609,In_986);
or U315 (N_315,In_1570,In_1187);
or U316 (N_316,In_1067,In_1499);
nor U317 (N_317,In_1746,In_1411);
or U318 (N_318,In_454,In_265);
and U319 (N_319,In_736,In_610);
nor U320 (N_320,In_211,In_2245);
nor U321 (N_321,In_2522,In_111);
xor U322 (N_322,In_1789,In_2680);
and U323 (N_323,In_1338,In_2862);
xor U324 (N_324,In_2486,In_159);
or U325 (N_325,In_1102,In_458);
nor U326 (N_326,In_835,In_651);
nor U327 (N_327,In_2055,In_598);
xnor U328 (N_328,In_1432,In_2084);
xor U329 (N_329,In_867,In_1185);
xor U330 (N_330,In_1551,In_2603);
nor U331 (N_331,In_2063,In_1925);
or U332 (N_332,In_1555,In_91);
and U333 (N_333,In_2000,In_1528);
and U334 (N_334,In_702,In_2886);
xor U335 (N_335,In_1770,In_1778);
nand U336 (N_336,In_1241,In_701);
or U337 (N_337,In_2441,In_2275);
nand U338 (N_338,In_1808,In_1161);
xor U339 (N_339,In_168,In_144);
nand U340 (N_340,In_174,In_1700);
xnor U341 (N_341,In_432,In_224);
or U342 (N_342,In_1237,In_1373);
nor U343 (N_343,In_1037,In_2216);
and U344 (N_344,In_2503,In_1396);
nand U345 (N_345,In_1723,In_1002);
xor U346 (N_346,In_2443,In_2797);
and U347 (N_347,In_951,In_1080);
nand U348 (N_348,In_1386,In_147);
xnor U349 (N_349,In_2331,In_2635);
and U350 (N_350,In_558,In_2708);
xnor U351 (N_351,In_935,In_1759);
or U352 (N_352,In_1826,In_1175);
xor U353 (N_353,In_1126,In_1022);
xor U354 (N_354,In_542,In_2843);
or U355 (N_355,In_1929,In_2731);
nor U356 (N_356,In_2925,In_688);
nor U357 (N_357,In_1676,In_617);
nor U358 (N_358,In_2641,In_1088);
or U359 (N_359,In_2665,In_1486);
or U360 (N_360,In_2392,In_2492);
xor U361 (N_361,In_2075,In_160);
xor U362 (N_362,In_541,In_2071);
xor U363 (N_363,In_1553,In_1853);
and U364 (N_364,In_2535,In_484);
nand U365 (N_365,In_1876,In_657);
xor U366 (N_366,In_34,In_1954);
and U367 (N_367,In_2651,In_1941);
and U368 (N_368,In_2430,In_142);
nand U369 (N_369,In_846,In_2358);
nand U370 (N_370,In_1609,In_1588);
or U371 (N_371,In_2545,In_868);
or U372 (N_372,In_1711,In_52);
and U373 (N_373,In_944,In_1008);
nand U374 (N_374,In_1694,In_1825);
nand U375 (N_375,In_1071,In_1270);
nor U376 (N_376,In_2645,In_2633);
or U377 (N_377,In_2532,In_6);
and U378 (N_378,In_1403,In_533);
nand U379 (N_379,In_1867,In_1835);
nor U380 (N_380,In_1054,In_2559);
xnor U381 (N_381,In_2877,In_2544);
nand U382 (N_382,In_901,In_2286);
xor U383 (N_383,In_741,In_2412);
and U384 (N_384,In_1390,In_2698);
nand U385 (N_385,In_1964,In_2502);
or U386 (N_386,In_329,In_1306);
and U387 (N_387,In_613,In_1837);
or U388 (N_388,In_140,In_360);
and U389 (N_389,In_1502,In_1295);
or U390 (N_390,In_225,In_1548);
nor U391 (N_391,In_2819,In_1707);
nand U392 (N_392,In_1841,In_1839);
and U393 (N_393,In_495,In_2838);
nor U394 (N_394,In_2496,In_299);
and U395 (N_395,In_2425,In_2281);
nand U396 (N_396,In_1893,In_2770);
and U397 (N_397,In_2755,In_826);
and U398 (N_398,In_2869,In_1168);
or U399 (N_399,In_2661,In_1634);
and U400 (N_400,In_637,In_2310);
and U401 (N_401,In_2670,In_708);
or U402 (N_402,In_1180,In_369);
nor U403 (N_403,In_686,In_190);
or U404 (N_404,In_1687,In_1614);
nand U405 (N_405,In_724,In_387);
and U406 (N_406,In_2108,In_2600);
xor U407 (N_407,In_2111,In_1582);
or U408 (N_408,In_1441,In_19);
nand U409 (N_409,In_1675,In_1038);
and U410 (N_410,In_2932,In_36);
or U411 (N_411,In_1783,In_1978);
and U412 (N_412,In_1249,In_845);
or U413 (N_413,In_860,In_2005);
nand U414 (N_414,In_1065,In_2639);
xor U415 (N_415,In_56,In_1508);
xor U416 (N_416,In_43,In_2849);
xor U417 (N_417,In_422,In_2895);
nor U418 (N_418,In_1276,In_2445);
and U419 (N_419,In_973,In_1974);
and U420 (N_420,In_1660,In_215);
xnor U421 (N_421,In_514,In_831);
and U422 (N_422,In_936,In_1767);
nand U423 (N_423,In_2839,In_992);
and U424 (N_424,In_2208,In_2205);
nand U425 (N_425,In_2169,In_2263);
and U426 (N_426,In_86,In_1151);
nor U427 (N_427,In_1931,In_1945);
nor U428 (N_428,In_2253,In_83);
xnor U429 (N_429,In_154,In_234);
or U430 (N_430,In_653,In_1869);
nor U431 (N_431,In_1771,In_957);
xnor U432 (N_432,In_1490,In_2604);
or U433 (N_433,In_2162,In_1048);
and U434 (N_434,In_386,In_555);
nor U435 (N_435,In_426,In_1027);
xor U436 (N_436,In_641,In_1972);
and U437 (N_437,In_374,In_2656);
xnor U438 (N_438,In_1475,In_76);
xor U439 (N_439,In_2312,In_721);
nand U440 (N_440,In_180,In_2984);
nor U441 (N_441,In_999,In_306);
xnor U442 (N_442,In_2217,In_2476);
nor U443 (N_443,In_549,In_75);
or U444 (N_444,In_1,In_2186);
xnor U445 (N_445,In_2558,In_576);
nor U446 (N_446,In_1683,In_2664);
nand U447 (N_447,In_2632,In_1855);
or U448 (N_448,In_822,In_2531);
nor U449 (N_449,In_1245,In_1476);
or U450 (N_450,In_204,In_419);
xnor U451 (N_451,In_328,In_2338);
and U452 (N_452,In_1184,In_64);
xor U453 (N_453,In_2479,In_373);
or U454 (N_454,In_1852,In_988);
xor U455 (N_455,In_1443,In_1636);
nor U456 (N_456,In_66,In_1820);
nor U457 (N_457,In_2438,In_2626);
and U458 (N_458,In_312,In_2772);
xor U459 (N_459,In_395,In_1091);
xnor U460 (N_460,In_2715,In_2193);
nand U461 (N_461,In_2093,In_2422);
nor U462 (N_462,In_1115,In_1335);
nor U463 (N_463,In_2313,In_2926);
nand U464 (N_464,In_1874,In_332);
or U465 (N_465,In_2806,In_2504);
nand U466 (N_466,In_625,In_2686);
or U467 (N_467,In_792,In_827);
nand U468 (N_468,In_335,In_1765);
nand U469 (N_469,In_1699,In_2137);
nor U470 (N_470,In_2840,In_187);
nand U471 (N_471,In_2148,In_2857);
nor U472 (N_472,In_2157,In_2841);
and U473 (N_473,In_2041,In_1671);
nand U474 (N_474,In_1289,In_967);
and U475 (N_475,In_1340,In_2337);
or U476 (N_476,In_1217,In_1488);
xor U477 (N_477,In_809,In_565);
nand U478 (N_478,In_1096,In_2828);
or U479 (N_479,In_890,In_2867);
and U480 (N_480,In_730,In_886);
or U481 (N_481,In_33,In_2799);
nand U482 (N_482,In_2825,In_849);
xnor U483 (N_483,In_1961,In_2760);
or U484 (N_484,In_585,In_1688);
and U485 (N_485,In_2178,In_1147);
nand U486 (N_486,In_2644,In_782);
or U487 (N_487,In_1169,In_780);
nand U488 (N_488,In_1152,In_949);
and U489 (N_489,In_1109,In_2273);
and U490 (N_490,In_1100,In_2420);
and U491 (N_491,In_631,In_2214);
or U492 (N_492,In_1542,In_1993);
and U493 (N_493,In_2017,In_806);
xnor U494 (N_494,In_163,In_668);
nand U495 (N_495,In_903,In_2565);
xnor U496 (N_496,In_481,In_803);
nor U497 (N_497,In_808,In_2845);
nand U498 (N_498,In_889,In_153);
nor U499 (N_499,In_786,In_1640);
nand U500 (N_500,In_659,In_311);
nor U501 (N_501,In_2693,In_2730);
nand U502 (N_502,In_1834,In_1447);
xnor U503 (N_503,In_2667,In_818);
and U504 (N_504,In_1379,In_2117);
or U505 (N_505,In_2740,In_1400);
and U506 (N_506,In_2620,In_2523);
and U507 (N_507,In_998,In_1807);
nor U508 (N_508,In_383,In_1654);
nor U509 (N_509,In_1580,In_1734);
xor U510 (N_510,In_1509,In_216);
xor U511 (N_511,In_301,In_2260);
or U512 (N_512,In_877,In_2832);
and U513 (N_513,In_813,In_1155);
nor U514 (N_514,In_87,In_17);
or U515 (N_515,In_1984,In_1315);
nand U516 (N_516,In_25,In_1829);
nand U517 (N_517,In_2024,In_14);
or U518 (N_518,In_2575,In_131);
and U519 (N_519,In_27,In_167);
nor U520 (N_520,In_2964,In_1463);
or U521 (N_521,In_1638,In_1286);
and U522 (N_522,In_1354,In_1625);
nor U523 (N_523,In_1626,In_275);
or U524 (N_524,In_1673,In_483);
nor U525 (N_525,In_1033,In_7);
xnor U526 (N_526,In_1051,In_649);
nand U527 (N_527,In_1523,In_2340);
xor U528 (N_528,In_1584,In_635);
nand U529 (N_529,In_2473,In_393);
nor U530 (N_530,In_207,In_2417);
nor U531 (N_531,In_2295,In_2153);
xor U532 (N_532,In_2437,In_1226);
and U533 (N_533,In_1014,In_2227);
and U534 (N_534,In_31,In_1236);
nor U535 (N_535,In_2931,In_1342);
and U536 (N_536,In_2818,In_1062);
nand U537 (N_537,In_2395,In_768);
nor U538 (N_538,In_1935,In_963);
nor U539 (N_539,In_1677,In_1888);
nand U540 (N_540,In_714,In_173);
nand U541 (N_541,In_1231,In_2311);
nor U542 (N_542,In_2505,In_723);
xor U543 (N_543,In_2394,In_2863);
and U544 (N_544,In_1992,In_1618);
xor U545 (N_545,In_1907,In_863);
and U546 (N_546,In_781,In_424);
and U547 (N_547,In_1637,In_2210);
xnor U548 (N_548,In_1428,In_2324);
nand U549 (N_549,In_706,In_2247);
and U550 (N_550,In_2961,In_2671);
nor U551 (N_551,In_722,In_921);
or U552 (N_552,In_705,In_1437);
nor U553 (N_553,In_2714,In_1693);
xor U554 (N_554,In_2585,In_1167);
xor U555 (N_555,In_537,In_2777);
xor U556 (N_556,In_2121,In_2339);
xor U557 (N_557,In_209,In_2524);
xnor U558 (N_558,In_2050,In_1606);
and U559 (N_559,In_115,In_297);
and U560 (N_560,In_1078,In_1018);
nor U561 (N_561,In_573,In_2012);
and U562 (N_562,In_279,In_2787);
nor U563 (N_563,In_1520,In_1442);
nand U564 (N_564,In_2334,In_78);
and U565 (N_565,In_2357,In_2741);
or U566 (N_566,In_725,In_1412);
or U567 (N_567,In_2085,In_596);
nand U568 (N_568,In_1814,In_1813);
or U569 (N_569,In_769,In_1632);
or U570 (N_570,In_1782,In_2534);
xor U571 (N_571,In_1822,In_2220);
or U572 (N_572,In_1076,In_289);
nand U573 (N_573,In_1419,In_2341);
or U574 (N_574,In_2624,In_2033);
and U575 (N_575,In_1243,In_2375);
or U576 (N_576,In_563,In_2977);
or U577 (N_577,In_522,In_487);
xnor U578 (N_578,In_1421,In_24);
nor U579 (N_579,In_948,In_2673);
and U580 (N_580,In_754,In_302);
nand U581 (N_581,In_2419,In_337);
xor U582 (N_582,In_98,In_493);
xnor U583 (N_583,In_2728,In_905);
xnor U584 (N_584,In_2536,In_2879);
and U585 (N_585,In_447,In_1681);
nor U586 (N_586,In_1776,In_377);
xor U587 (N_587,In_508,In_1159);
and U588 (N_588,In_114,In_859);
nand U589 (N_589,In_1032,In_1352);
or U590 (N_590,In_788,In_438);
or U591 (N_591,In_2615,In_1657);
nor U592 (N_592,In_1260,In_2727);
xnor U593 (N_593,In_623,In_2675);
xor U594 (N_594,In_1424,In_1034);
or U595 (N_595,In_1957,In_416);
nand U596 (N_596,In_2386,In_2351);
or U597 (N_597,In_1744,In_1190);
or U598 (N_598,In_1556,In_1300);
xor U599 (N_599,In_1762,In_2147);
xnor U600 (N_600,In_811,In_1084);
xor U601 (N_601,In_2343,In_1722);
nand U602 (N_602,In_1924,In_1157);
nand U603 (N_603,In_2628,In_917);
and U604 (N_604,In_1110,In_1087);
and U605 (N_605,In_1450,In_1323);
and U606 (N_606,In_941,In_2128);
and U607 (N_607,In_1891,In_1267);
and U608 (N_608,In_71,In_1873);
and U609 (N_609,In_1312,In_1053);
xnor U610 (N_610,In_2820,In_251);
nand U611 (N_611,In_257,In_1261);
nand U612 (N_612,In_1073,In_2048);
nor U613 (N_613,In_169,In_46);
or U614 (N_614,In_650,In_1122);
nor U615 (N_615,In_1708,In_2878);
or U616 (N_616,In_959,In_2436);
nor U617 (N_617,In_2992,In_2411);
and U618 (N_618,In_1188,In_762);
and U619 (N_619,In_1238,In_463);
and U620 (N_620,In_2448,In_1532);
nand U621 (N_621,In_2685,In_1838);
nand U622 (N_622,In_923,In_452);
xor U623 (N_623,In_2060,In_927);
and U624 (N_624,In_567,In_2243);
and U625 (N_625,In_288,In_778);
nor U626 (N_626,In_1766,In_2892);
and U627 (N_627,In_2037,In_296);
nand U628 (N_628,In_2576,In_2197);
nand U629 (N_629,In_1622,In_2100);
nand U630 (N_630,In_2950,In_2572);
or U631 (N_631,In_2781,In_1446);
or U632 (N_632,In_2416,In_750);
and U633 (N_633,In_1112,In_2403);
nand U634 (N_634,In_2542,In_2623);
xor U635 (N_635,In_2021,In_2616);
nor U636 (N_636,In_1039,In_1162);
and U637 (N_637,In_2177,In_1547);
and U638 (N_638,In_2218,In_2875);
and U639 (N_639,In_457,In_146);
and U640 (N_640,In_2555,In_2953);
nand U641 (N_641,In_2373,In_1578);
and U642 (N_642,In_60,In_1879);
or U643 (N_643,In_2107,In_2958);
nand U644 (N_644,In_1516,In_2938);
nor U645 (N_645,In_2115,In_2229);
nor U646 (N_646,In_2928,In_2102);
or U647 (N_647,In_2870,In_1427);
xor U648 (N_648,In_2552,In_178);
and U649 (N_649,In_99,In_1514);
or U650 (N_650,In_2903,In_562);
nand U651 (N_651,In_2244,In_2219);
and U652 (N_652,In_1768,In_1971);
or U653 (N_653,In_469,In_2830);
xor U654 (N_654,In_2991,In_2088);
and U655 (N_655,In_1650,In_1836);
nor U656 (N_656,In_2471,In_2894);
nor U657 (N_657,In_1163,In_1304);
and U658 (N_658,In_372,In_317);
and U659 (N_659,In_2683,In_2135);
xor U660 (N_660,In_938,In_1518);
and U661 (N_661,In_84,In_2692);
xnor U662 (N_662,In_420,In_1787);
or U663 (N_663,In_990,In_1562);
and U664 (N_664,In_2883,In_925);
and U665 (N_665,In_2743,In_1868);
or U666 (N_666,In_2998,In_1794);
nor U667 (N_667,In_2458,In_1932);
nor U668 (N_668,In_1557,In_2861);
nand U669 (N_669,In_29,In_1533);
xor U670 (N_670,In_1377,In_528);
or U671 (N_671,In_1620,In_2759);
or U672 (N_672,In_2261,In_117);
xor U673 (N_673,In_2199,In_552);
nand U674 (N_674,In_2586,In_587);
and U675 (N_675,In_2264,In_2750);
or U676 (N_676,In_1878,In_1890);
nand U677 (N_677,In_2499,In_1136);
nor U678 (N_678,In_2816,In_914);
xor U679 (N_679,In_2494,In_1196);
nor U680 (N_680,In_2609,In_2409);
or U681 (N_681,In_208,In_1074);
and U682 (N_682,In_2090,In_2734);
nor U683 (N_683,In_35,In_564);
or U684 (N_684,In_1257,In_2391);
nand U685 (N_685,In_881,In_2927);
xor U686 (N_686,In_2077,In_1724);
or U687 (N_687,In_1715,In_2352);
and U688 (N_688,In_2691,In_2801);
nor U689 (N_689,In_883,In_1194);
and U690 (N_690,In_915,In_1271);
nand U691 (N_691,In_2574,In_1160);
or U692 (N_692,In_2707,In_2541);
or U693 (N_693,In_1402,In_470);
or U694 (N_694,In_934,In_1422);
nor U695 (N_695,In_1521,In_100);
nor U696 (N_696,In_89,In_1760);
xnor U697 (N_697,In_1960,In_448);
nor U698 (N_698,In_2364,In_1720);
xnor U699 (N_699,In_871,In_1847);
or U700 (N_700,In_2271,In_1991);
nand U701 (N_701,In_1537,In_10);
or U702 (N_702,In_729,In_680);
and U703 (N_703,In_1730,In_1466);
and U704 (N_704,In_2182,In_1389);
or U705 (N_705,In_2997,In_1395);
and U706 (N_706,In_2307,In_1571);
xor U707 (N_707,In_1713,In_382);
nand U708 (N_708,In_2028,In_862);
xnor U709 (N_709,In_305,In_2461);
nand U710 (N_710,In_314,In_32);
nor U711 (N_711,In_413,In_1259);
xnor U712 (N_712,In_23,In_1164);
or U713 (N_713,In_497,In_2256);
nor U714 (N_714,In_1430,In_389);
and U715 (N_715,In_2749,In_388);
nor U716 (N_716,In_1726,In_1337);
nor U717 (N_717,In_546,In_18);
or U718 (N_718,In_2874,In_2563);
and U719 (N_719,In_186,In_2161);
nand U720 (N_720,In_1973,In_960);
nor U721 (N_721,In_238,In_2081);
nor U722 (N_722,In_566,In_548);
nand U723 (N_723,In_270,In_157);
xor U724 (N_724,In_2056,In_1118);
nor U725 (N_725,In_2922,In_1994);
nor U726 (N_726,In_2780,In_135);
nor U727 (N_727,In_1860,In_1436);
nor U728 (N_728,In_2140,In_94);
and U729 (N_729,In_2495,In_2722);
nand U730 (N_730,In_2940,In_2912);
nand U731 (N_731,In_2109,In_2621);
xnor U732 (N_732,In_1605,In_1346);
nand U733 (N_733,In_896,In_774);
xnor U734 (N_734,In_2239,In_1884);
nor U735 (N_735,In_902,In_1393);
nand U736 (N_736,In_804,In_96);
nand U737 (N_737,In_295,In_1558);
nand U738 (N_738,In_2887,In_1001);
nand U739 (N_739,In_2789,In_1322);
xor U740 (N_740,In_1012,In_232);
nor U741 (N_741,In_1290,In_268);
nand U742 (N_742,In_755,In_1685);
nor U743 (N_743,In_2995,In_2393);
nor U744 (N_744,In_1501,In_262);
or U745 (N_745,In_2378,In_2663);
nand U746 (N_746,In_1716,In_2521);
nand U747 (N_747,In_2305,In_2297);
nor U748 (N_748,In_471,In_336);
xor U749 (N_749,In_2094,In_1915);
xor U750 (N_750,In_503,In_1242);
nand U751 (N_751,In_197,In_113);
nand U752 (N_752,In_910,In_1007);
nor U753 (N_753,In_2007,In_2190);
or U754 (N_754,In_928,In_206);
xnor U755 (N_755,In_412,In_734);
xnor U756 (N_756,In_2483,In_1011);
nor U757 (N_757,In_660,In_1856);
or U758 (N_758,In_2226,In_569);
or U759 (N_759,In_2527,In_188);
nand U760 (N_760,In_16,In_1481);
nor U761 (N_761,In_54,In_2920);
nor U762 (N_762,In_2610,In_1999);
nand U763 (N_763,In_1214,In_331);
nor U764 (N_764,In_2941,In_47);
and U765 (N_765,In_2567,In_290);
xnor U766 (N_766,In_2282,In_1052);
nand U767 (N_767,In_1266,In_2885);
or U768 (N_768,In_820,In_132);
xor U769 (N_769,In_242,In_261);
nor U770 (N_770,In_2737,In_2860);
nor U771 (N_771,In_2865,In_520);
nor U772 (N_772,In_2149,In_2512);
nand U773 (N_773,In_2318,In_2733);
nand U774 (N_774,In_1207,In_744);
nor U775 (N_775,In_1060,In_184);
xor U776 (N_776,In_2269,In_183);
nor U777 (N_777,In_2515,In_2466);
nor U778 (N_778,In_1952,In_2618);
xor U779 (N_779,In_2601,In_2301);
nand U780 (N_780,In_689,In_1353);
xnor U781 (N_781,In_1709,In_367);
nand U782 (N_782,In_2396,In_854);
and U783 (N_783,In_1222,In_1799);
nand U784 (N_784,In_1388,In_855);
and U785 (N_785,In_1805,In_870);
or U786 (N_786,In_1383,In_865);
or U787 (N_787,In_2711,In_194);
and U788 (N_788,In_1517,In_2187);
or U789 (N_789,In_1823,In_407);
and U790 (N_790,In_606,In_2937);
xnor U791 (N_791,In_1391,In_1535);
or U792 (N_792,In_88,In_2959);
or U793 (N_793,In_2703,In_2660);
nor U794 (N_794,In_525,In_2606);
xnor U795 (N_795,In_955,In_108);
xnor U796 (N_796,In_1418,In_1599);
and U797 (N_797,In_324,In_795);
or U798 (N_798,In_1742,In_1020);
nor U799 (N_799,In_1510,In_529);
and U800 (N_800,In_1210,In_1449);
or U801 (N_801,In_776,In_2408);
xnor U802 (N_802,In_264,In_2983);
xnor U803 (N_803,In_2401,In_2376);
and U804 (N_804,In_1220,In_742);
nand U805 (N_805,In_53,In_292);
and U806 (N_806,In_1444,In_2506);
xnor U807 (N_807,In_267,In_2433);
or U808 (N_808,In_1668,In_123);
nor U809 (N_809,In_480,In_2184);
nor U810 (N_810,In_685,In_1392);
or U811 (N_811,In_467,In_2688);
nand U812 (N_812,In_2834,In_2934);
and U813 (N_813,In_384,In_2584);
xor U814 (N_814,In_417,In_907);
or U815 (N_815,In_2796,In_764);
nor U816 (N_816,In_2594,In_220);
xnor U817 (N_817,In_1448,In_1414);
nor U818 (N_818,In_1754,In_636);
xor U819 (N_819,In_2598,In_436);
nor U820 (N_820,In_141,In_783);
or U821 (N_821,In_69,In_1044);
or U822 (N_822,In_1892,In_2292);
nor U823 (N_823,In_2890,In_952);
nor U824 (N_824,In_1604,In_2629);
nor U825 (N_825,In_189,In_1462);
nor U826 (N_826,In_1977,In_1567);
and U827 (N_827,In_713,In_1986);
or U828 (N_828,In_2844,In_2276);
and U829 (N_829,In_1321,In_1534);
nor U830 (N_830,In_1385,In_11);
nor U831 (N_831,In_130,In_488);
nand U832 (N_832,In_1649,In_638);
or U833 (N_833,In_1142,In_504);
nor U834 (N_834,In_2303,In_991);
nor U835 (N_835,In_1987,In_1079);
nand U836 (N_836,In_2478,In_2978);
or U837 (N_837,In_1848,In_2697);
nor U838 (N_838,In_2255,In_2346);
nand U839 (N_839,In_202,In_2811);
and U840 (N_840,In_2520,In_898);
xor U841 (N_841,In_2933,In_370);
nor U842 (N_842,In_1644,In_2968);
xor U843 (N_843,In_2891,In_2823);
xor U844 (N_844,In_2188,In_904);
or U845 (N_845,In_1949,In_2540);
and U846 (N_846,In_2490,In_1703);
nor U847 (N_847,In_2913,In_578);
and U848 (N_848,In_179,In_1301);
nor U849 (N_849,In_414,In_1524);
xnor U850 (N_850,In_626,In_1045);
and U851 (N_851,In_1747,In_472);
xor U852 (N_852,In_391,In_344);
or U853 (N_853,In_718,In_592);
or U854 (N_854,In_2444,In_2516);
xnor U855 (N_855,In_1937,In_1174);
nor U856 (N_856,In_57,In_175);
xnor U857 (N_857,In_961,In_103);
xnor U858 (N_858,In_334,In_551);
or U859 (N_859,In_1872,In_553);
and U860 (N_860,In_2385,In_599);
xnor U861 (N_861,In_2096,In_128);
xnor U862 (N_862,In_731,In_378);
xor U863 (N_863,In_287,In_1903);
nor U864 (N_864,In_409,In_577);
nor U865 (N_865,In_1211,In_45);
nand U866 (N_866,In_531,In_1729);
nand U867 (N_867,In_3,In_2602);
xnor U868 (N_868,In_2201,In_1308);
and U869 (N_869,In_1998,In_622);
xor U870 (N_870,In_1576,In_93);
xor U871 (N_871,In_2582,In_793);
and U872 (N_872,In_2131,In_150);
nand U873 (N_873,In_2457,In_2036);
nor U874 (N_874,In_2631,In_1976);
nand U875 (N_875,In_832,In_970);
xnor U876 (N_876,In_2270,In_1951);
xnor U877 (N_877,In_2952,In_1779);
nand U878 (N_878,In_1108,In_2069);
or U879 (N_879,In_2449,In_747);
or U880 (N_880,In_1922,In_687);
and U881 (N_881,In_2350,In_2808);
or U882 (N_882,In_2589,In_1368);
or U883 (N_883,In_954,In_1928);
nor U884 (N_884,In_2167,In_1227);
and U885 (N_885,In_2897,In_1143);
nand U886 (N_886,In_2277,In_1455);
nand U887 (N_887,In_398,In_410);
nand U888 (N_888,In_1850,In_1579);
nor U889 (N_889,In_1137,In_2911);
nor U890 (N_890,In_1740,In_1305);
xnor U891 (N_891,In_1094,In_2853);
and U892 (N_892,In_2942,In_1262);
nand U893 (N_893,In_1364,In_2500);
and U894 (N_894,In_2407,In_1068);
and U895 (N_895,In_1282,In_2404);
xor U896 (N_896,In_1075,In_1603);
or U897 (N_897,In_1183,In_1669);
xnor U898 (N_898,In_2080,In_2397);
nor U899 (N_899,In_842,In_892);
xor U900 (N_900,In_2191,In_2679);
xnor U901 (N_901,In_1593,In_1970);
nand U902 (N_902,In_1495,In_2636);
or U903 (N_903,In_281,In_441);
xnor U904 (N_904,In_1031,In_341);
and U905 (N_905,In_1512,In_2595);
nand U906 (N_906,In_1343,In_2674);
nand U907 (N_907,In_1531,In_247);
and U908 (N_908,In_2975,In_2798);
and U909 (N_909,In_339,In_2379);
or U910 (N_910,In_1064,In_1479);
xor U911 (N_911,In_451,In_2511);
nand U912 (N_912,In_1348,In_2652);
nand U913 (N_913,In_1756,In_1704);
nor U914 (N_914,In_2701,In_1566);
and U915 (N_915,In_282,In_2291);
nor U916 (N_916,In_699,In_2824);
nand U917 (N_917,In_2982,In_2905);
xnor U918 (N_918,In_1492,In_1712);
nand U919 (N_919,In_2510,In_2452);
or U920 (N_920,In_1786,In_2439);
and U921 (N_921,In_630,In_1358);
nor U922 (N_922,In_1381,In_589);
or U923 (N_923,In_425,In_359);
or U924 (N_924,In_1661,In_523);
nor U925 (N_925,In_603,In_166);
nand U926 (N_926,In_1631,In_95);
or U927 (N_927,In_1696,In_2484);
nand U928 (N_928,In_2064,In_2336);
nor U929 (N_929,In_707,In_2043);
and U930 (N_930,In_501,In_2990);
nand U931 (N_931,In_1347,In_2400);
or U932 (N_932,In_2918,In_379);
nor U933 (N_933,In_1101,In_913);
nor U934 (N_934,In_226,In_726);
nor U935 (N_935,In_979,In_773);
or U936 (N_936,In_2943,In_619);
nor U937 (N_937,In_203,In_1969);
nor U938 (N_938,In_1124,In_2224);
or U939 (N_939,In_2003,In_2951);
xnor U940 (N_940,In_519,In_1251);
or U941 (N_941,In_253,In_1472);
nor U942 (N_942,In_316,In_61);
or U943 (N_943,In_2957,In_1281);
xor U944 (N_944,In_719,In_1963);
or U945 (N_945,In_2002,In_2026);
xnor U946 (N_946,In_2785,In_1844);
and U947 (N_947,In_1328,In_1690);
or U948 (N_948,In_1982,In_958);
nand U949 (N_949,In_1178,In_1651);
nor U950 (N_950,In_2110,In_2590);
xnor U951 (N_951,In_2049,In_1367);
nand U952 (N_952,In_164,In_1058);
nand U953 (N_953,In_58,In_2833);
xnor U954 (N_954,In_2015,In_1917);
and U955 (N_955,In_1491,In_1686);
nand U956 (N_956,In_1154,In_2119);
or U957 (N_957,In_1777,In_2299);
nand U958 (N_958,In_1679,In_1946);
xor U959 (N_959,In_2752,In_594);
xnor U960 (N_960,In_28,In_2827);
and U961 (N_961,In_1228,In_1127);
nor U962 (N_962,In_349,In_2038);
nand U963 (N_963,In_1324,In_1736);
nand U964 (N_964,In_2164,In_571);
nor U965 (N_965,In_1775,In_1072);
or U966 (N_966,In_277,In_269);
nor U967 (N_967,In_1177,In_2622);
nor U968 (N_968,In_856,In_434);
and U969 (N_969,In_491,In_1727);
or U970 (N_970,In_2368,In_2501);
nand U971 (N_971,In_222,In_1375);
nor U972 (N_972,In_138,In_2802);
nand U973 (N_973,In_2533,In_1313);
or U974 (N_974,In_746,In_1948);
or U975 (N_975,In_258,In_2014);
xor U976 (N_976,In_2791,In_1280);
nor U977 (N_977,In_2155,In_403);
nand U978 (N_978,In_437,In_2380);
xor U979 (N_979,In_874,In_2431);
nand U980 (N_980,In_2006,In_2062);
and U981 (N_981,In_456,In_1090);
xor U982 (N_982,In_582,In_643);
nand U983 (N_983,In_245,In_2613);
and U984 (N_984,In_44,In_1057);
or U985 (N_985,In_2176,In_1334);
xnor U986 (N_986,In_1587,In_906);
or U987 (N_987,In_418,In_2543);
nand U988 (N_988,In_2593,In_2200);
and U989 (N_989,In_2530,In_2427);
or U990 (N_990,In_1769,In_2124);
xnor U991 (N_991,In_787,In_2835);
xnor U992 (N_992,In_2235,In_2642);
and U993 (N_993,In_1153,In_2814);
nand U994 (N_994,In_2643,In_953);
nor U995 (N_995,In_1735,In_770);
xor U996 (N_996,In_2116,In_2383);
nand U997 (N_997,In_672,In_893);
nand U998 (N_998,In_2316,In_2788);
and U999 (N_999,In_1473,In_879);
or U1000 (N_1000,In_2491,In_1218);
and U1001 (N_1001,In_1682,In_1751);
nor U1002 (N_1002,In_2614,In_1750);
and U1003 (N_1003,In_671,In_2103);
or U1004 (N_1004,In_1691,In_2672);
xor U1005 (N_1005,In_2142,In_1043);
xor U1006 (N_1006,In_1134,In_692);
and U1007 (N_1007,In_217,In_805);
nand U1008 (N_1008,In_715,In_1522);
nor U1009 (N_1009,In_2762,In_2097);
and U1010 (N_1010,In_740,In_446);
or U1011 (N_1011,In_538,In_1904);
or U1012 (N_1012,In_2390,In_1714);
xor U1013 (N_1013,In_2289,In_1404);
nand U1014 (N_1014,In_2517,In_517);
xnor U1015 (N_1015,In_1474,In_2287);
and U1016 (N_1016,In_124,In_1042);
nand U1017 (N_1017,In_13,In_2924);
or U1018 (N_1018,In_2290,In_48);
and U1019 (N_1019,In_2657,In_2095);
nor U1020 (N_1020,In_1047,In_1200);
nand U1021 (N_1021,In_1545,In_1913);
xor U1022 (N_1022,In_2240,In_2086);
nand U1023 (N_1023,In_2447,In_2355);
nand U1024 (N_1024,In_2366,In_2784);
nand U1025 (N_1025,In_2944,In_1710);
or U1026 (N_1026,In_109,In_839);
xor U1027 (N_1027,In_1017,In_574);
or U1028 (N_1028,In_1719,In_2813);
or U1029 (N_1029,In_1093,In_2192);
or U1030 (N_1030,In_2881,In_2966);
nor U1031 (N_1031,In_460,In_1958);
nor U1032 (N_1032,In_1525,In_2786);
xor U1033 (N_1033,In_836,In_966);
or U1034 (N_1034,In_2315,In_547);
nand U1035 (N_1035,In_342,In_320);
and U1036 (N_1036,In_2418,In_918);
nand U1037 (N_1037,In_1757,In_2004);
nor U1038 (N_1038,In_1465,In_932);
and U1039 (N_1039,In_476,In_496);
nand U1040 (N_1040,In_1360,In_873);
or U1041 (N_1041,In_1309,In_634);
nor U1042 (N_1042,In_1049,In_1370);
xor U1043 (N_1043,In_2866,In_1684);
nand U1044 (N_1044,In_2718,In_2371);
nor U1045 (N_1045,In_544,In_2267);
nor U1046 (N_1046,In_981,In_2057);
nor U1047 (N_1047,In_2266,In_1706);
and U1048 (N_1048,In_2406,In_127);
and U1049 (N_1049,In_291,In_728);
nor U1050 (N_1050,In_891,In_2181);
or U1051 (N_1051,In_801,In_521);
and U1052 (N_1052,In_1861,In_327);
and U1053 (N_1053,In_931,In_618);
and U1054 (N_1054,In_1059,In_462);
or U1055 (N_1055,In_248,In_1927);
nand U1056 (N_1056,In_2031,In_1831);
and U1057 (N_1057,In_956,In_1416);
and U1058 (N_1058,In_632,In_679);
and U1059 (N_1059,In_2771,In_2174);
xor U1060 (N_1060,In_1296,In_1288);
xnor U1061 (N_1061,In_1208,In_193);
xnor U1062 (N_1062,In_1239,In_2904);
and U1063 (N_1063,In_1464,In_2556);
xor U1064 (N_1064,In_2194,In_1798);
or U1065 (N_1065,In_1171,In_554);
or U1066 (N_1066,In_399,In_1041);
and U1067 (N_1067,In_700,In_1149);
nor U1068 (N_1068,In_872,In_1672);
or U1069 (N_1069,In_2739,In_1106);
or U1070 (N_1070,In_1146,In_1781);
or U1071 (N_1071,In_2335,In_1828);
nand U1072 (N_1072,In_2252,In_402);
xnor U1073 (N_1073,In_2213,In_1376);
nor U1074 (N_1074,In_1790,In_1480);
xnor U1075 (N_1075,In_392,In_709);
and U1076 (N_1076,In_241,In_850);
nand U1077 (N_1077,In_2022,In_2234);
and U1078 (N_1078,In_758,In_2965);
nand U1079 (N_1079,In_2134,In_79);
nand U1080 (N_1080,In_2405,In_2089);
or U1081 (N_1081,In_2529,In_145);
nor U1082 (N_1082,In_191,In_559);
nand U1083 (N_1083,In_2705,In_116);
and U1084 (N_1084,In_2159,In_2306);
and U1085 (N_1085,In_2195,In_1902);
nand U1086 (N_1086,In_1601,In_294);
or U1087 (N_1087,In_2319,In_678);
nand U1088 (N_1088,In_532,In_1215);
nand U1089 (N_1089,In_2294,In_543);
nor U1090 (N_1090,In_1763,In_2070);
nand U1091 (N_1091,In_161,In_1851);
nand U1092 (N_1092,In_1627,In_971);
or U1093 (N_1093,In_1484,In_1647);
nor U1094 (N_1094,In_2330,In_2758);
xor U1095 (N_1095,In_1478,In_74);
nand U1096 (N_1096,In_710,In_771);
nand U1097 (N_1097,In_1026,In_2974);
nor U1098 (N_1098,In_340,In_1113);
xor U1099 (N_1099,In_1363,In_1104);
or U1100 (N_1100,In_2960,In_1351);
and U1101 (N_1101,In_2677,In_1540);
and U1102 (N_1102,In_2498,In_940);
nor U1103 (N_1103,In_2872,In_2145);
and U1104 (N_1104,In_1203,In_2144);
and U1105 (N_1105,In_263,In_1244);
xor U1106 (N_1106,In_1413,In_790);
and U1107 (N_1107,In_2011,In_1857);
xnor U1108 (N_1108,In_994,In_2435);
or U1109 (N_1109,In_1725,In_1689);
xnor U1110 (N_1110,In_2717,In_2754);
nand U1111 (N_1111,In_2896,In_200);
or U1112 (N_1112,In_1019,In_2723);
nand U1113 (N_1113,In_1028,In_1515);
xnor U1114 (N_1114,In_223,In_2899);
and U1115 (N_1115,In_1434,In_2010);
nor U1116 (N_1116,In_2087,In_1232);
nor U1117 (N_1117,In_1832,In_1223);
or U1118 (N_1118,In_2902,In_293);
nor U1119 (N_1119,In_1784,In_712);
and U1120 (N_1120,In_1985,In_1483);
and U1121 (N_1121,In_2637,In_1349);
and U1122 (N_1122,In_2206,In_2774);
and U1123 (N_1123,In_639,In_2551);
nor U1124 (N_1124,In_1273,In_1055);
nand U1125 (N_1125,In_1410,In_1356);
or U1126 (N_1126,In_1840,In_673);
nand U1127 (N_1127,In_1458,In_1914);
or U1128 (N_1128,In_2898,In_2381);
xnor U1129 (N_1129,In_1250,In_120);
or U1130 (N_1130,In_1938,In_1621);
or U1131 (N_1131,In_122,In_2497);
nand U1132 (N_1132,In_1979,In_1082);
xor U1133 (N_1133,In_1219,In_852);
xnor U1134 (N_1134,In_664,In_2769);
and U1135 (N_1135,In_945,In_2463);
or U1136 (N_1136,In_1965,In_1302);
nor U1137 (N_1137,In_1382,In_1291);
nor U1138 (N_1138,In_2424,In_2970);
xnor U1139 (N_1139,In_1635,In_1761);
xnor U1140 (N_1140,In_139,In_1881);
nand U1141 (N_1141,In_2761,In_2065);
and U1142 (N_1142,In_1642,In_1496);
xor U1143 (N_1143,In_539,In_1345);
xor U1144 (N_1144,In_2790,In_2171);
or U1145 (N_1145,In_924,In_2979);
nand U1146 (N_1146,In_1586,In_763);
or U1147 (N_1147,In_1493,In_1824);
or U1148 (N_1148,In_1350,In_1845);
nand U1149 (N_1149,In_1221,In_1069);
nor U1150 (N_1150,In_1731,In_1590);
nand U1151 (N_1151,In_1871,In_2907);
xor U1152 (N_1152,In_1804,In_2689);
nor U1153 (N_1153,In_516,In_1591);
or U1154 (N_1154,In_1577,In_2105);
nor U1155 (N_1155,In_125,In_2092);
nand U1156 (N_1156,In_73,In_285);
nor U1157 (N_1157,In_2493,In_1589);
and U1158 (N_1158,In_1061,In_401);
xnor U1159 (N_1159,In_50,In_1617);
nand U1160 (N_1160,In_2285,In_1374);
xnor U1161 (N_1161,In_1575,In_760);
xnor U1162 (N_1162,In_1897,In_2168);
and U1163 (N_1163,In_2309,In_1355);
or U1164 (N_1164,In_656,In_1081);
nand U1165 (N_1165,In_2118,In_500);
nor U1166 (N_1166,In_2042,In_2580);
xnor U1167 (N_1167,In_919,In_1561);
and U1168 (N_1168,In_1800,In_908);
nand U1169 (N_1169,In_1156,In_2625);
or U1170 (N_1170,In_775,In_1666);
nor U1171 (N_1171,In_2347,In_751);
and U1172 (N_1172,In_231,In_1268);
nand U1173 (N_1173,In_570,In_2354);
or U1174 (N_1174,In_2724,In_319);
nand U1175 (N_1175,In_22,In_1918);
nand U1176 (N_1176,In_2597,In_1117);
nand U1177 (N_1177,In_735,In_12);
and U1178 (N_1178,In_674,In_356);
nor U1179 (N_1179,In_1085,In_1125);
xor U1180 (N_1180,In_2826,In_2810);
xnor U1181 (N_1181,In_1148,In_2209);
nand U1182 (N_1182,In_1645,In_930);
and U1183 (N_1183,In_507,In_1435);
xnor U1184 (N_1184,In_2279,In_2101);
or U1185 (N_1185,In_1284,In_2146);
nand U1186 (N_1186,In_355,In_1150);
xor U1187 (N_1187,In_1864,In_2232);
nand U1188 (N_1188,In_1753,In_308);
nor U1189 (N_1189,In_1803,In_739);
or U1190 (N_1190,In_1029,In_2320);
or U1191 (N_1191,In_1698,In_1310);
or U1192 (N_1192,In_2133,In_49);
or U1193 (N_1193,In_1967,In_1489);
nor U1194 (N_1194,In_2812,In_1511);
xnor U1195 (N_1195,In_2864,In_2388);
nor U1196 (N_1196,In_1066,In_621);
xor U1197 (N_1197,In_1619,In_2342);
and U1198 (N_1198,In_2539,In_1083);
nand U1199 (N_1199,In_430,In_2231);
nand U1200 (N_1200,In_1176,In_1264);
and U1201 (N_1201,In_2414,In_977);
nand U1202 (N_1202,In_1678,In_2389);
and U1203 (N_1203,In_829,In_1795);
and U1204 (N_1204,In_1608,In_512);
or U1205 (N_1205,In_2850,In_1186);
nor U1206 (N_1206,In_1469,In_1940);
nor U1207 (N_1207,In_1201,In_1331);
nand U1208 (N_1208,In_2249,In_513);
nand U1209 (N_1209,In_2963,In_2460);
and U1210 (N_1210,In_2475,In_2858);
or U1211 (N_1211,In_1966,In_1643);
nand U1212 (N_1212,In_511,In_711);
or U1213 (N_1213,In_461,In_1810);
and U1214 (N_1214,In_1983,In_156);
and U1215 (N_1215,In_5,In_1095);
nor U1216 (N_1216,In_933,In_2198);
nand U1217 (N_1217,In_1780,In_824);
nand U1218 (N_1218,In_80,In_978);
xor U1219 (N_1219,In_1272,In_929);
nor U1220 (N_1220,In_2246,In_357);
and U1221 (N_1221,In_2668,In_1453);
or U1222 (N_1222,In_1748,In_1341);
or U1223 (N_1223,In_819,In_997);
xor U1224 (N_1224,In_408,In_584);
nor U1225 (N_1225,In_1145,In_2696);
xnor U1226 (N_1226,In_1138,In_1468);
nor U1227 (N_1227,In_1130,In_218);
or U1228 (N_1228,In_2488,In_2948);
and U1229 (N_1229,In_2387,In_1882);
or U1230 (N_1230,In_568,In_1013);
xor U1231 (N_1231,In_0,In_1230);
nand U1232 (N_1232,In_1544,In_1733);
or U1233 (N_1233,In_1854,In_1739);
or U1234 (N_1234,In_51,In_105);
nor U1235 (N_1235,In_1006,In_1718);
nand U1236 (N_1236,In_346,In_2052);
or U1237 (N_1237,In_2030,In_1633);
or U1238 (N_1238,In_2363,In_97);
nor U1239 (N_1239,In_1870,In_1639);
nand U1240 (N_1240,In_1471,In_2317);
nor U1241 (N_1241,In_1934,In_2180);
xnor U1242 (N_1242,In_1900,In_2104);
xor U1243 (N_1243,In_2265,In_669);
xnor U1244 (N_1244,In_1025,In_259);
and U1245 (N_1245,In_2514,In_2591);
or U1246 (N_1246,In_1613,In_1494);
nand U1247 (N_1247,In_1336,In_885);
nor U1248 (N_1248,In_816,In_2078);
nor U1249 (N_1249,In_1009,In_833);
nor U1250 (N_1250,In_642,In_1592);
nand U1251 (N_1251,In_727,In_1943);
nor U1252 (N_1252,In_982,In_2112);
nor U1253 (N_1253,In_861,In_2298);
and U1254 (N_1254,In_1123,In_2113);
nand U1255 (N_1255,In_2583,In_2768);
nand U1256 (N_1256,In_965,In_942);
or U1257 (N_1257,In_63,In_298);
or U1258 (N_1258,In_2163,In_2356);
nor U1259 (N_1259,In_640,In_2020);
nor U1260 (N_1260,In_158,In_315);
xor U1261 (N_1261,In_118,In_2909);
or U1262 (N_1262,In_2154,In_345);
nor U1263 (N_1263,In_2,In_2809);
xor U1264 (N_1264,In_2470,In_1326);
nor U1265 (N_1265,In_1842,In_2283);
nor U1266 (N_1266,In_2196,In_2669);
xor U1267 (N_1267,In_1883,In_2776);
or U1268 (N_1268,In_2519,In_2141);
or U1269 (N_1269,In_428,In_869);
xnor U1270 (N_1270,In_1816,In_785);
and U1271 (N_1271,In_766,In_717);
nor U1272 (N_1272,In_2935,In_2434);
nor U1273 (N_1273,In_2842,In_2349);
xor U1274 (N_1274,In_266,In_1173);
nand U1275 (N_1275,In_322,In_2207);
xor U1276 (N_1276,In_2653,In_1255);
xor U1277 (N_1277,In_1530,In_2658);
and U1278 (N_1278,In_396,In_2528);
nor U1279 (N_1279,In_761,In_1936);
or U1280 (N_1280,In_2873,In_2945);
or U1281 (N_1281,In_527,In_1487);
nor U1282 (N_1282,In_2702,In_2792);
nand U1283 (N_1283,In_1170,In_1297);
nor U1284 (N_1284,In_2605,In_112);
or U1285 (N_1285,In_772,In_2634);
nor U1286 (N_1286,In_478,In_55);
and U1287 (N_1287,In_572,In_2578);
nand U1288 (N_1288,In_993,In_975);
and U1289 (N_1289,In_1283,In_2353);
nand U1290 (N_1290,In_779,In_1016);
nand U1291 (N_1291,In_2956,In_474);
nor U1292 (N_1292,In_2560,In_1933);
or U1293 (N_1293,In_397,In_676);
or U1294 (N_1294,In_1950,In_2348);
or U1295 (N_1295,In_984,In_690);
or U1296 (N_1296,In_987,In_2009);
nand U1297 (N_1297,In_1209,In_2837);
and U1298 (N_1298,In_404,In_655);
xor U1299 (N_1299,In_1339,In_882);
and U1300 (N_1300,In_1460,In_2472);
and U1301 (N_1301,In_20,In_152);
xor U1302 (N_1302,In_38,In_1600);
or U1303 (N_1303,In_749,In_880);
xor U1304 (N_1304,In_2564,In_1880);
xnor U1305 (N_1305,In_2704,In_560);
nor U1306 (N_1306,In_2638,In_1611);
nand U1307 (N_1307,In_1802,In_309);
xor U1308 (N_1308,In_628,In_1905);
or U1309 (N_1309,In_2805,In_133);
nor U1310 (N_1310,In_597,In_400);
nand U1311 (N_1311,In_1461,In_909);
and U1312 (N_1312,In_485,In_2630);
xnor U1313 (N_1313,In_1456,In_1665);
or U1314 (N_1314,In_2136,In_946);
nand U1315 (N_1315,In_255,In_1005);
nand U1316 (N_1316,In_875,In_2690);
nor U1317 (N_1317,In_1910,In_1674);
xor U1318 (N_1318,In_465,In_421);
nand U1319 (N_1319,In_119,In_40);
nand U1320 (N_1320,In_2025,In_1898);
and U1321 (N_1321,In_1318,In_1420);
nor U1322 (N_1322,In_1407,In_1959);
nand U1323 (N_1323,In_59,In_221);
nor U1324 (N_1324,In_198,In_2756);
and U1325 (N_1325,In_2278,In_1550);
nor U1326 (N_1326,In_2855,In_2332);
nor U1327 (N_1327,In_2706,In_1764);
or U1328 (N_1328,In_821,In_912);
or U1329 (N_1329,In_2212,In_449);
nor U1330 (N_1330,In_814,In_2852);
nor U1331 (N_1331,In_2588,In_2284);
or U1332 (N_1332,In_2066,In_1035);
or U1333 (N_1333,In_939,In_1980);
nand U1334 (N_1334,In_466,In_42);
xnor U1335 (N_1335,In_1092,In_2571);
or U1336 (N_1336,In_1919,In_243);
xnor U1337 (N_1337,In_1258,In_101);
xor U1338 (N_1338,In_1968,In_2649);
or U1339 (N_1339,In_1616,In_348);
and U1340 (N_1340,In_2687,In_1366);
and U1341 (N_1341,In_2293,In_325);
and U1342 (N_1342,In_2328,In_752);
nor U1343 (N_1343,In_1752,In_1988);
nor U1344 (N_1344,In_2732,In_2143);
nand U1345 (N_1345,In_2654,In_1717);
or U1346 (N_1346,In_976,In_2429);
nor U1347 (N_1347,In_196,In_1721);
nand U1348 (N_1348,In_620,In_2525);
and U1349 (N_1349,In_2345,In_2987);
nand U1350 (N_1350,In_2647,In_2889);
xor U1351 (N_1351,In_1128,In_394);
or U1352 (N_1352,In_611,In_581);
and U1353 (N_1353,In_2646,In_1863);
nor U1354 (N_1354,In_2456,In_1482);
xnor U1355 (N_1355,In_633,In_536);
and U1356 (N_1356,In_1050,In_2747);
xor U1357 (N_1357,In_1191,In_2040);
and U1358 (N_1358,In_433,In_343);
or U1359 (N_1359,In_1394,In_1827);
or U1360 (N_1360,In_1552,In_894);
nand U1361 (N_1361,In_1911,In_1316);
or U1362 (N_1362,In_1303,In_851);
xor U1363 (N_1363,In_354,In_580);
nor U1364 (N_1364,In_365,In_26);
nand U1365 (N_1365,In_586,In_1815);
nand U1366 (N_1366,In_550,In_1371);
or U1367 (N_1367,In_2744,In_2179);
and U1368 (N_1368,In_2775,In_2027);
xor U1369 (N_1369,In_1862,In_486);
and U1370 (N_1370,In_1438,In_834);
xnor U1371 (N_1371,In_2611,In_405);
and U1372 (N_1372,In_1655,In_985);
nand U1373 (N_1373,In_530,In_968);
and U1374 (N_1374,In_477,In_2082);
or U1375 (N_1375,In_227,In_2921);
and U1376 (N_1376,In_2986,In_677);
and U1377 (N_1377,In_667,In_201);
nor U1378 (N_1378,In_2304,In_1877);
nand U1379 (N_1379,In_2972,In_1653);
xnor U1380 (N_1380,In_1607,In_996);
xnor U1381 (N_1381,In_1497,In_743);
nor U1382 (N_1382,In_1797,In_1583);
nand U1383 (N_1383,In_2906,In_455);
nand U1384 (N_1384,In_1121,In_1997);
or U1385 (N_1385,In_1415,In_1785);
nor U1386 (N_1386,In_1549,In_962);
nand U1387 (N_1387,In_2745,In_283);
or U1388 (N_1388,In_2233,In_1274);
nor U1389 (N_1389,In_1107,In_1975);
nor U1390 (N_1390,In_2251,In_1596);
nor U1391 (N_1391,In_1278,In_104);
nor U1392 (N_1392,In_176,In_1953);
nand U1393 (N_1393,In_1896,In_1500);
or U1394 (N_1394,In_607,In_604);
or U1395 (N_1395,In_1397,In_1314);
and U1396 (N_1396,In_515,In_1467);
xnor U1397 (N_1397,In_1387,In_526);
and U1398 (N_1398,In_1246,In_797);
xnor U1399 (N_1399,In_1181,In_561);
nand U1400 (N_1400,In_602,In_575);
xnor U1401 (N_1401,In_2713,In_974);
and U1402 (N_1402,In_358,In_244);
nand U1403 (N_1403,In_647,In_1745);
or U1404 (N_1404,In_1541,In_439);
nor U1405 (N_1405,In_1192,In_1398);
nor U1406 (N_1406,In_2682,In_1774);
and U1407 (N_1407,In_2753,In_753);
and U1408 (N_1408,In_85,In_1811);
nor U1409 (N_1409,In_1070,In_182);
and U1410 (N_1410,In_1995,In_1947);
and U1411 (N_1411,In_148,In_1040);
and U1412 (N_1412,In_2547,In_2268);
nand U1413 (N_1413,In_791,In_2513);
nand U1414 (N_1414,In_2300,In_2783);
xor U1415 (N_1415,In_2321,In_313);
or U1416 (N_1416,In_847,In_165);
xnor U1417 (N_1417,In_1772,In_876);
or U1418 (N_1418,In_172,In_1641);
nor U1419 (N_1419,In_62,In_800);
nor U1420 (N_1420,In_1702,In_2884);
or U1421 (N_1421,In_2325,In_1293);
and U1422 (N_1422,In_658,In_1172);
nor U1423 (N_1423,In_1506,In_2029);
and U1424 (N_1424,In_1646,In_70);
nor U1425 (N_1425,In_2489,In_1179);
nor U1426 (N_1426,In_2782,In_1144);
and U1427 (N_1427,In_2607,In_2413);
xor U1428 (N_1428,In_694,In_1325);
or U1429 (N_1429,In_1440,In_2695);
and U1430 (N_1430,In_2410,In_2047);
xnor U1431 (N_1431,In_2053,In_411);
and U1432 (N_1432,In_2374,In_1454);
nand U1433 (N_1433,In_1792,In_765);
or U1434 (N_1434,In_2067,In_601);
nor U1435 (N_1435,In_2729,In_1865);
xor U1436 (N_1436,In_1554,In_1889);
xnor U1437 (N_1437,In_1457,In_2023);
xor U1438 (N_1438,In_1895,In_1329);
or U1439 (N_1439,In_2367,In_2130);
and U1440 (N_1440,In_627,In_841);
nor U1441 (N_1441,In_2566,In_2929);
nor U1442 (N_1442,In_506,In_1664);
nor U1443 (N_1443,In_1485,In_2955);
and U1444 (N_1444,In_368,In_662);
xnor U1445 (N_1445,In_1380,In_540);
or U1446 (N_1446,In_900,In_2487);
nand U1447 (N_1447,In_1663,In_1327);
xnor U1448 (N_1448,In_1212,In_812);
xor U1449 (N_1449,In_249,In_2581);
and U1450 (N_1450,In_2120,In_697);
and U1451 (N_1451,In_1256,In_1912);
nand U1452 (N_1452,In_129,In_745);
nand U1453 (N_1453,In_654,In_330);
nor U1454 (N_1454,In_911,In_2659);
nor U1455 (N_1455,In_1585,In_2451);
nor U1456 (N_1456,In_303,In_2359);
nor U1457 (N_1457,In_608,In_1216);
nor U1458 (N_1458,In_1086,In_1737);
nand U1459 (N_1459,In_1459,In_1287);
nand U1460 (N_1460,In_2561,In_828);
and U1461 (N_1461,In_1843,In_2215);
nand U1462 (N_1462,In_1539,In_2446);
nor U1463 (N_1463,In_272,In_65);
xnor U1464 (N_1464,In_2949,In_1791);
or U1465 (N_1465,In_1656,In_2599);
xnor U1466 (N_1466,In_2455,In_2684);
nand U1467 (N_1467,In_2971,In_843);
nor U1468 (N_1468,In_2051,In_1189);
xnor U1469 (N_1469,In_375,In_210);
xor U1470 (N_1470,In_1010,In_884);
nor U1471 (N_1471,In_2985,In_2382);
and U1472 (N_1472,In_1849,In_2074);
nand U1473 (N_1473,In_1695,In_1817);
nor U1474 (N_1474,In_429,In_1015);
xnor U1475 (N_1475,In_2773,In_1498);
xor U1476 (N_1476,In_645,In_943);
nor U1477 (N_1477,In_2939,In_155);
nor U1478 (N_1478,In_1089,In_2831);
nor U1479 (N_1479,In_2211,In_2518);
xnor U1480 (N_1480,In_1921,In_333);
nor U1481 (N_1481,In_1199,In_41);
nand U1482 (N_1482,In_2577,In_2204);
nor U1483 (N_1483,In_1859,In_665);
and U1484 (N_1484,In_2467,In_732);
and U1485 (N_1485,In_1728,In_459);
xor U1486 (N_1486,In_1365,In_1133);
nor U1487 (N_1487,In_1926,In_518);
and U1488 (N_1488,In_777,In_1277);
xor U1489 (N_1489,In_535,In_1279);
nor U1490 (N_1490,In_2901,In_237);
and U1491 (N_1491,In_2068,In_1899);
nand U1492 (N_1492,In_1319,In_2236);
xor U1493 (N_1493,In_2954,In_556);
nor U1494 (N_1494,In_136,In_2076);
or U1495 (N_1495,In_137,In_2859);
or U1496 (N_1496,In_2908,In_1630);
or U1497 (N_1497,In_1120,In_2666);
nor U1498 (N_1498,In_1598,In_406);
xnor U1499 (N_1499,In_1773,In_756);
and U1500 (N_1500,In_2384,In_1865);
xnor U1501 (N_1501,In_2516,In_532);
nor U1502 (N_1502,In_2553,In_2358);
or U1503 (N_1503,In_1090,In_2105);
nor U1504 (N_1504,In_2702,In_1601);
or U1505 (N_1505,In_2085,In_2536);
nand U1506 (N_1506,In_577,In_418);
xor U1507 (N_1507,In_2261,In_1426);
and U1508 (N_1508,In_2644,In_1993);
xor U1509 (N_1509,In_731,In_904);
nand U1510 (N_1510,In_935,In_823);
or U1511 (N_1511,In_510,In_802);
nand U1512 (N_1512,In_1541,In_2518);
or U1513 (N_1513,In_2457,In_2326);
nand U1514 (N_1514,In_1067,In_2499);
nor U1515 (N_1515,In_708,In_1786);
and U1516 (N_1516,In_1054,In_1799);
nor U1517 (N_1517,In_756,In_1969);
nand U1518 (N_1518,In_0,In_2405);
or U1519 (N_1519,In_2749,In_1493);
nand U1520 (N_1520,In_2640,In_462);
and U1521 (N_1521,In_272,In_717);
or U1522 (N_1522,In_2999,In_1147);
or U1523 (N_1523,In_2966,In_2917);
nor U1524 (N_1524,In_2531,In_2853);
or U1525 (N_1525,In_1937,In_1744);
or U1526 (N_1526,In_818,In_2651);
or U1527 (N_1527,In_318,In_2832);
and U1528 (N_1528,In_2666,In_1323);
xnor U1529 (N_1529,In_2045,In_2411);
and U1530 (N_1530,In_1583,In_97);
xor U1531 (N_1531,In_1131,In_2280);
or U1532 (N_1532,In_1310,In_373);
or U1533 (N_1533,In_1641,In_602);
xor U1534 (N_1534,In_819,In_2881);
xnor U1535 (N_1535,In_565,In_1998);
nor U1536 (N_1536,In_2156,In_2819);
and U1537 (N_1537,In_2790,In_1700);
xnor U1538 (N_1538,In_1381,In_1281);
or U1539 (N_1539,In_314,In_958);
nor U1540 (N_1540,In_1438,In_2086);
or U1541 (N_1541,In_844,In_2191);
or U1542 (N_1542,In_2639,In_303);
or U1543 (N_1543,In_1602,In_686);
or U1544 (N_1544,In_2059,In_1979);
or U1545 (N_1545,In_1825,In_1197);
nor U1546 (N_1546,In_265,In_1719);
nand U1547 (N_1547,In_1710,In_2657);
nand U1548 (N_1548,In_1149,In_2179);
xnor U1549 (N_1549,In_2148,In_1378);
or U1550 (N_1550,In_1334,In_2359);
xor U1551 (N_1551,In_1578,In_437);
and U1552 (N_1552,In_992,In_356);
nand U1553 (N_1553,In_1625,In_125);
nand U1554 (N_1554,In_198,In_1643);
nand U1555 (N_1555,In_915,In_1082);
xnor U1556 (N_1556,In_296,In_298);
nand U1557 (N_1557,In_2724,In_544);
xnor U1558 (N_1558,In_419,In_2886);
or U1559 (N_1559,In_1182,In_397);
or U1560 (N_1560,In_2554,In_2040);
nor U1561 (N_1561,In_185,In_970);
nand U1562 (N_1562,In_2295,In_867);
or U1563 (N_1563,In_1834,In_1666);
xnor U1564 (N_1564,In_218,In_2851);
nor U1565 (N_1565,In_1046,In_485);
xnor U1566 (N_1566,In_310,In_1069);
nor U1567 (N_1567,In_2821,In_533);
nor U1568 (N_1568,In_2008,In_2949);
nor U1569 (N_1569,In_1180,In_308);
nor U1570 (N_1570,In_951,In_930);
xnor U1571 (N_1571,In_1457,In_2544);
and U1572 (N_1572,In_201,In_1369);
and U1573 (N_1573,In_1878,In_1699);
nor U1574 (N_1574,In_1628,In_1785);
and U1575 (N_1575,In_2137,In_282);
xor U1576 (N_1576,In_587,In_1289);
nor U1577 (N_1577,In_1349,In_1779);
nand U1578 (N_1578,In_620,In_2600);
xor U1579 (N_1579,In_2245,In_1238);
nand U1580 (N_1580,In_97,In_1460);
nor U1581 (N_1581,In_1707,In_1391);
nand U1582 (N_1582,In_731,In_1053);
nand U1583 (N_1583,In_2482,In_751);
xor U1584 (N_1584,In_2071,In_1294);
or U1585 (N_1585,In_2140,In_1912);
nand U1586 (N_1586,In_424,In_2935);
xor U1587 (N_1587,In_411,In_2614);
xor U1588 (N_1588,In_1789,In_1343);
nor U1589 (N_1589,In_1352,In_1012);
xor U1590 (N_1590,In_1763,In_2748);
or U1591 (N_1591,In_1497,In_2466);
nor U1592 (N_1592,In_107,In_18);
xnor U1593 (N_1593,In_1518,In_2692);
and U1594 (N_1594,In_926,In_1326);
and U1595 (N_1595,In_2396,In_2516);
xor U1596 (N_1596,In_712,In_1172);
nor U1597 (N_1597,In_1731,In_1703);
xnor U1598 (N_1598,In_707,In_1545);
xor U1599 (N_1599,In_1559,In_1831);
or U1600 (N_1600,In_2913,In_727);
xnor U1601 (N_1601,In_2689,In_764);
nand U1602 (N_1602,In_497,In_352);
or U1603 (N_1603,In_239,In_327);
xor U1604 (N_1604,In_1658,In_2721);
nand U1605 (N_1605,In_2330,In_2499);
or U1606 (N_1606,In_617,In_311);
nor U1607 (N_1607,In_2323,In_65);
nand U1608 (N_1608,In_840,In_5);
xnor U1609 (N_1609,In_2228,In_1632);
nor U1610 (N_1610,In_49,In_2399);
and U1611 (N_1611,In_1129,In_1199);
nor U1612 (N_1612,In_2374,In_2140);
xor U1613 (N_1613,In_593,In_754);
or U1614 (N_1614,In_236,In_2636);
nand U1615 (N_1615,In_680,In_1543);
nor U1616 (N_1616,In_532,In_1390);
nand U1617 (N_1617,In_587,In_1187);
nor U1618 (N_1618,In_1289,In_557);
and U1619 (N_1619,In_2574,In_1860);
or U1620 (N_1620,In_2061,In_178);
and U1621 (N_1621,In_17,In_352);
nand U1622 (N_1622,In_2643,In_2144);
or U1623 (N_1623,In_1458,In_2183);
nor U1624 (N_1624,In_1877,In_1195);
or U1625 (N_1625,In_1855,In_1894);
or U1626 (N_1626,In_5,In_1415);
or U1627 (N_1627,In_1354,In_399);
xnor U1628 (N_1628,In_1192,In_2944);
xor U1629 (N_1629,In_1180,In_889);
nor U1630 (N_1630,In_2717,In_2427);
or U1631 (N_1631,In_2534,In_1914);
or U1632 (N_1632,In_942,In_2763);
xnor U1633 (N_1633,In_1551,In_1377);
and U1634 (N_1634,In_2432,In_141);
xnor U1635 (N_1635,In_619,In_1417);
and U1636 (N_1636,In_743,In_1318);
nand U1637 (N_1637,In_1057,In_1706);
and U1638 (N_1638,In_934,In_897);
nor U1639 (N_1639,In_1171,In_208);
xor U1640 (N_1640,In_2476,In_264);
nor U1641 (N_1641,In_31,In_2198);
nand U1642 (N_1642,In_2600,In_1688);
xnor U1643 (N_1643,In_499,In_1980);
and U1644 (N_1644,In_1339,In_2916);
and U1645 (N_1645,In_2481,In_2123);
nand U1646 (N_1646,In_2891,In_1512);
xnor U1647 (N_1647,In_260,In_1784);
xnor U1648 (N_1648,In_118,In_2562);
or U1649 (N_1649,In_2138,In_1970);
nor U1650 (N_1650,In_2046,In_44);
nor U1651 (N_1651,In_2260,In_2133);
nand U1652 (N_1652,In_1080,In_1469);
nand U1653 (N_1653,In_262,In_2683);
nor U1654 (N_1654,In_2228,In_2317);
or U1655 (N_1655,In_2062,In_848);
and U1656 (N_1656,In_2685,In_2738);
xor U1657 (N_1657,In_532,In_2014);
nor U1658 (N_1658,In_190,In_829);
xor U1659 (N_1659,In_1329,In_2790);
xnor U1660 (N_1660,In_321,In_1685);
or U1661 (N_1661,In_158,In_2734);
nor U1662 (N_1662,In_56,In_274);
nor U1663 (N_1663,In_1124,In_2262);
or U1664 (N_1664,In_492,In_1981);
or U1665 (N_1665,In_486,In_663);
or U1666 (N_1666,In_1820,In_1231);
and U1667 (N_1667,In_233,In_194);
and U1668 (N_1668,In_1999,In_1594);
nand U1669 (N_1669,In_1779,In_549);
or U1670 (N_1670,In_2040,In_1009);
and U1671 (N_1671,In_562,In_1321);
nand U1672 (N_1672,In_750,In_2612);
and U1673 (N_1673,In_1501,In_888);
and U1674 (N_1674,In_2885,In_1960);
or U1675 (N_1675,In_2442,In_1224);
and U1676 (N_1676,In_1572,In_2593);
nor U1677 (N_1677,In_1701,In_1734);
or U1678 (N_1678,In_997,In_2982);
and U1679 (N_1679,In_1578,In_167);
and U1680 (N_1680,In_1649,In_1299);
xnor U1681 (N_1681,In_99,In_1242);
xor U1682 (N_1682,In_2625,In_1313);
nand U1683 (N_1683,In_1099,In_2851);
nand U1684 (N_1684,In_958,In_2282);
or U1685 (N_1685,In_1199,In_1717);
and U1686 (N_1686,In_842,In_1835);
xnor U1687 (N_1687,In_2082,In_99);
nor U1688 (N_1688,In_417,In_2634);
or U1689 (N_1689,In_198,In_2625);
or U1690 (N_1690,In_2550,In_2192);
nand U1691 (N_1691,In_1762,In_176);
and U1692 (N_1692,In_2847,In_2037);
and U1693 (N_1693,In_2221,In_1669);
nor U1694 (N_1694,In_1714,In_1845);
or U1695 (N_1695,In_73,In_974);
nor U1696 (N_1696,In_865,In_853);
xnor U1697 (N_1697,In_1352,In_1626);
xor U1698 (N_1698,In_818,In_1025);
nor U1699 (N_1699,In_951,In_2857);
and U1700 (N_1700,In_2619,In_2744);
nand U1701 (N_1701,In_53,In_1890);
and U1702 (N_1702,In_1461,In_35);
xor U1703 (N_1703,In_93,In_77);
nor U1704 (N_1704,In_1429,In_133);
nand U1705 (N_1705,In_1138,In_2448);
or U1706 (N_1706,In_2708,In_307);
and U1707 (N_1707,In_2647,In_1686);
or U1708 (N_1708,In_1351,In_12);
and U1709 (N_1709,In_782,In_2282);
xnor U1710 (N_1710,In_713,In_42);
nor U1711 (N_1711,In_990,In_180);
and U1712 (N_1712,In_1592,In_1239);
xnor U1713 (N_1713,In_837,In_762);
xnor U1714 (N_1714,In_2922,In_1331);
or U1715 (N_1715,In_2680,In_1691);
and U1716 (N_1716,In_863,In_1288);
nor U1717 (N_1717,In_503,In_2419);
nand U1718 (N_1718,In_2748,In_1851);
or U1719 (N_1719,In_2375,In_2022);
nor U1720 (N_1720,In_1511,In_1776);
nor U1721 (N_1721,In_273,In_2884);
and U1722 (N_1722,In_299,In_334);
or U1723 (N_1723,In_246,In_2939);
and U1724 (N_1724,In_2801,In_314);
nor U1725 (N_1725,In_2605,In_2296);
nor U1726 (N_1726,In_1477,In_2238);
xnor U1727 (N_1727,In_1591,In_2617);
nor U1728 (N_1728,In_2044,In_2478);
xnor U1729 (N_1729,In_50,In_2279);
nand U1730 (N_1730,In_878,In_48);
nor U1731 (N_1731,In_1523,In_1749);
nand U1732 (N_1732,In_163,In_1865);
and U1733 (N_1733,In_56,In_2067);
xor U1734 (N_1734,In_2229,In_439);
or U1735 (N_1735,In_2854,In_877);
nand U1736 (N_1736,In_2759,In_674);
nand U1737 (N_1737,In_1622,In_2015);
and U1738 (N_1738,In_249,In_227);
and U1739 (N_1739,In_98,In_277);
or U1740 (N_1740,In_1231,In_1963);
or U1741 (N_1741,In_2969,In_613);
or U1742 (N_1742,In_94,In_2100);
nor U1743 (N_1743,In_699,In_1278);
and U1744 (N_1744,In_2733,In_2605);
nor U1745 (N_1745,In_737,In_790);
nor U1746 (N_1746,In_760,In_2432);
nand U1747 (N_1747,In_806,In_563);
nor U1748 (N_1748,In_1518,In_2723);
nor U1749 (N_1749,In_1994,In_2141);
nor U1750 (N_1750,In_2346,In_1877);
nor U1751 (N_1751,In_2841,In_2831);
and U1752 (N_1752,In_2953,In_55);
or U1753 (N_1753,In_1061,In_2165);
nor U1754 (N_1754,In_488,In_2051);
xor U1755 (N_1755,In_519,In_2511);
nor U1756 (N_1756,In_1570,In_349);
and U1757 (N_1757,In_1412,In_37);
or U1758 (N_1758,In_2343,In_989);
nand U1759 (N_1759,In_69,In_1042);
xor U1760 (N_1760,In_1149,In_2242);
xor U1761 (N_1761,In_113,In_2022);
nand U1762 (N_1762,In_134,In_2944);
xor U1763 (N_1763,In_1906,In_1639);
and U1764 (N_1764,In_2266,In_1068);
and U1765 (N_1765,In_811,In_667);
nor U1766 (N_1766,In_786,In_1949);
and U1767 (N_1767,In_876,In_969);
nand U1768 (N_1768,In_511,In_2982);
or U1769 (N_1769,In_1851,In_1957);
and U1770 (N_1770,In_263,In_2639);
nor U1771 (N_1771,In_1212,In_2804);
nor U1772 (N_1772,In_2749,In_1753);
xor U1773 (N_1773,In_2078,In_1509);
xor U1774 (N_1774,In_2298,In_1421);
and U1775 (N_1775,In_1845,In_968);
nand U1776 (N_1776,In_1177,In_4);
nand U1777 (N_1777,In_1869,In_931);
nand U1778 (N_1778,In_2145,In_2688);
xnor U1779 (N_1779,In_2784,In_687);
xor U1780 (N_1780,In_1884,In_259);
xnor U1781 (N_1781,In_1553,In_64);
or U1782 (N_1782,In_1343,In_729);
and U1783 (N_1783,In_2883,In_2507);
and U1784 (N_1784,In_1969,In_1549);
xor U1785 (N_1785,In_2229,In_11);
and U1786 (N_1786,In_2877,In_1713);
and U1787 (N_1787,In_657,In_2544);
nand U1788 (N_1788,In_1977,In_2769);
xnor U1789 (N_1789,In_1261,In_2363);
nor U1790 (N_1790,In_2295,In_1697);
nand U1791 (N_1791,In_1711,In_2544);
or U1792 (N_1792,In_1155,In_1036);
or U1793 (N_1793,In_1409,In_1886);
or U1794 (N_1794,In_423,In_1192);
and U1795 (N_1795,In_361,In_2891);
or U1796 (N_1796,In_794,In_700);
or U1797 (N_1797,In_99,In_834);
nor U1798 (N_1798,In_2209,In_2885);
or U1799 (N_1799,In_2245,In_1610);
and U1800 (N_1800,In_2721,In_1021);
or U1801 (N_1801,In_1356,In_886);
nor U1802 (N_1802,In_1940,In_2125);
nand U1803 (N_1803,In_1815,In_1652);
or U1804 (N_1804,In_142,In_2686);
nand U1805 (N_1805,In_1012,In_1807);
and U1806 (N_1806,In_1316,In_331);
nor U1807 (N_1807,In_840,In_2665);
nor U1808 (N_1808,In_1204,In_2631);
nor U1809 (N_1809,In_178,In_990);
or U1810 (N_1810,In_1513,In_2439);
nand U1811 (N_1811,In_2894,In_1415);
and U1812 (N_1812,In_2593,In_2451);
xor U1813 (N_1813,In_1170,In_1477);
and U1814 (N_1814,In_937,In_1175);
xor U1815 (N_1815,In_2166,In_1054);
xor U1816 (N_1816,In_833,In_587);
xor U1817 (N_1817,In_881,In_573);
xor U1818 (N_1818,In_1348,In_1000);
nor U1819 (N_1819,In_2443,In_782);
or U1820 (N_1820,In_2509,In_2777);
xor U1821 (N_1821,In_892,In_1581);
or U1822 (N_1822,In_1108,In_1497);
xor U1823 (N_1823,In_810,In_400);
and U1824 (N_1824,In_1053,In_781);
and U1825 (N_1825,In_232,In_2794);
nor U1826 (N_1826,In_1014,In_1037);
or U1827 (N_1827,In_2923,In_985);
and U1828 (N_1828,In_1944,In_2752);
or U1829 (N_1829,In_2701,In_1930);
nor U1830 (N_1830,In_2893,In_2699);
xor U1831 (N_1831,In_1630,In_551);
and U1832 (N_1832,In_2953,In_1663);
nand U1833 (N_1833,In_1374,In_1250);
and U1834 (N_1834,In_2303,In_2873);
xor U1835 (N_1835,In_2844,In_2391);
nor U1836 (N_1836,In_301,In_2028);
nand U1837 (N_1837,In_2613,In_2882);
or U1838 (N_1838,In_2745,In_1524);
nor U1839 (N_1839,In_2784,In_394);
or U1840 (N_1840,In_2217,In_2475);
and U1841 (N_1841,In_2840,In_2286);
xnor U1842 (N_1842,In_2690,In_1562);
and U1843 (N_1843,In_1160,In_2086);
nor U1844 (N_1844,In_583,In_360);
nand U1845 (N_1845,In_1969,In_1253);
nor U1846 (N_1846,In_1034,In_737);
nand U1847 (N_1847,In_2731,In_1079);
nand U1848 (N_1848,In_1331,In_1405);
and U1849 (N_1849,In_2001,In_455);
nor U1850 (N_1850,In_1716,In_469);
xor U1851 (N_1851,In_1000,In_1902);
and U1852 (N_1852,In_557,In_779);
nor U1853 (N_1853,In_1884,In_2951);
and U1854 (N_1854,In_158,In_2221);
nor U1855 (N_1855,In_902,In_2859);
or U1856 (N_1856,In_2654,In_1427);
and U1857 (N_1857,In_312,In_2430);
xnor U1858 (N_1858,In_1747,In_1688);
nand U1859 (N_1859,In_2965,In_599);
or U1860 (N_1860,In_1887,In_2843);
and U1861 (N_1861,In_39,In_608);
and U1862 (N_1862,In_2048,In_1860);
nand U1863 (N_1863,In_1730,In_2496);
and U1864 (N_1864,In_1820,In_1066);
nand U1865 (N_1865,In_1176,In_657);
nor U1866 (N_1866,In_544,In_2199);
xnor U1867 (N_1867,In_312,In_1576);
xor U1868 (N_1868,In_1633,In_2059);
nor U1869 (N_1869,In_1082,In_2070);
or U1870 (N_1870,In_2195,In_864);
xor U1871 (N_1871,In_2850,In_1258);
and U1872 (N_1872,In_2176,In_2962);
nor U1873 (N_1873,In_1589,In_294);
and U1874 (N_1874,In_1308,In_1861);
or U1875 (N_1875,In_2521,In_1840);
xor U1876 (N_1876,In_2543,In_1092);
xor U1877 (N_1877,In_241,In_426);
nor U1878 (N_1878,In_154,In_694);
xnor U1879 (N_1879,In_719,In_1646);
nand U1880 (N_1880,In_177,In_1089);
nand U1881 (N_1881,In_1287,In_2494);
and U1882 (N_1882,In_250,In_1835);
and U1883 (N_1883,In_2096,In_1915);
nor U1884 (N_1884,In_585,In_633);
xnor U1885 (N_1885,In_432,In_495);
and U1886 (N_1886,In_1549,In_2498);
nor U1887 (N_1887,In_49,In_1747);
nor U1888 (N_1888,In_150,In_2077);
and U1889 (N_1889,In_2821,In_2335);
or U1890 (N_1890,In_801,In_2514);
or U1891 (N_1891,In_1234,In_1616);
or U1892 (N_1892,In_1537,In_2514);
nor U1893 (N_1893,In_196,In_1714);
nand U1894 (N_1894,In_2547,In_2427);
or U1895 (N_1895,In_383,In_994);
nand U1896 (N_1896,In_2576,In_2182);
or U1897 (N_1897,In_2067,In_1991);
nand U1898 (N_1898,In_1624,In_1775);
and U1899 (N_1899,In_1736,In_1016);
nand U1900 (N_1900,In_318,In_2841);
or U1901 (N_1901,In_137,In_1922);
xor U1902 (N_1902,In_824,In_774);
or U1903 (N_1903,In_1060,In_648);
nand U1904 (N_1904,In_2489,In_239);
xor U1905 (N_1905,In_1705,In_1846);
and U1906 (N_1906,In_522,In_428);
and U1907 (N_1907,In_859,In_925);
nand U1908 (N_1908,In_2489,In_2590);
or U1909 (N_1909,In_2154,In_2866);
and U1910 (N_1910,In_1577,In_1992);
or U1911 (N_1911,In_300,In_332);
and U1912 (N_1912,In_242,In_2574);
nand U1913 (N_1913,In_2114,In_1540);
nand U1914 (N_1914,In_345,In_1857);
or U1915 (N_1915,In_1861,In_1974);
and U1916 (N_1916,In_2947,In_2843);
nand U1917 (N_1917,In_818,In_2994);
and U1918 (N_1918,In_2457,In_2861);
nor U1919 (N_1919,In_2462,In_2025);
nand U1920 (N_1920,In_2620,In_1581);
xor U1921 (N_1921,In_2341,In_1283);
nand U1922 (N_1922,In_2951,In_1071);
xnor U1923 (N_1923,In_2962,In_1579);
or U1924 (N_1924,In_1493,In_494);
xor U1925 (N_1925,In_2689,In_442);
or U1926 (N_1926,In_1583,In_2613);
nand U1927 (N_1927,In_889,In_1704);
nor U1928 (N_1928,In_2671,In_2979);
nor U1929 (N_1929,In_2303,In_2014);
xnor U1930 (N_1930,In_1415,In_1485);
or U1931 (N_1931,In_2393,In_673);
xor U1932 (N_1932,In_1445,In_2557);
and U1933 (N_1933,In_1362,In_1184);
xor U1934 (N_1934,In_519,In_1843);
nor U1935 (N_1935,In_1722,In_2748);
nor U1936 (N_1936,In_2486,In_605);
xnor U1937 (N_1937,In_1209,In_2871);
xnor U1938 (N_1938,In_1928,In_2781);
and U1939 (N_1939,In_812,In_1701);
nor U1940 (N_1940,In_2364,In_869);
and U1941 (N_1941,In_566,In_1688);
nand U1942 (N_1942,In_2597,In_2261);
or U1943 (N_1943,In_2226,In_1740);
xnor U1944 (N_1944,In_2947,In_1850);
xnor U1945 (N_1945,In_969,In_353);
nand U1946 (N_1946,In_2687,In_2666);
or U1947 (N_1947,In_341,In_2703);
and U1948 (N_1948,In_1641,In_2232);
nor U1949 (N_1949,In_1583,In_809);
or U1950 (N_1950,In_1771,In_2182);
or U1951 (N_1951,In_935,In_2720);
nor U1952 (N_1952,In_1679,In_446);
or U1953 (N_1953,In_423,In_327);
nor U1954 (N_1954,In_2997,In_1055);
and U1955 (N_1955,In_882,In_2508);
or U1956 (N_1956,In_505,In_1173);
xnor U1957 (N_1957,In_661,In_1804);
nor U1958 (N_1958,In_786,In_746);
nand U1959 (N_1959,In_1462,In_1125);
or U1960 (N_1960,In_1343,In_1972);
nand U1961 (N_1961,In_2388,In_2421);
and U1962 (N_1962,In_2402,In_2160);
xor U1963 (N_1963,In_152,In_424);
nor U1964 (N_1964,In_1753,In_737);
nor U1965 (N_1965,In_2605,In_283);
nand U1966 (N_1966,In_1970,In_2216);
and U1967 (N_1967,In_2849,In_685);
and U1968 (N_1968,In_2285,In_2125);
or U1969 (N_1969,In_2099,In_1801);
or U1970 (N_1970,In_2773,In_1377);
xor U1971 (N_1971,In_448,In_496);
nor U1972 (N_1972,In_98,In_799);
nor U1973 (N_1973,In_185,In_2468);
and U1974 (N_1974,In_1167,In_2982);
nor U1975 (N_1975,In_1702,In_1692);
and U1976 (N_1976,In_968,In_2117);
xnor U1977 (N_1977,In_1469,In_1);
nor U1978 (N_1978,In_320,In_958);
and U1979 (N_1979,In_2200,In_1245);
nor U1980 (N_1980,In_2270,In_2478);
xnor U1981 (N_1981,In_700,In_2339);
nor U1982 (N_1982,In_677,In_1414);
and U1983 (N_1983,In_1280,In_619);
or U1984 (N_1984,In_139,In_1076);
or U1985 (N_1985,In_263,In_2662);
or U1986 (N_1986,In_1957,In_2098);
xnor U1987 (N_1987,In_2369,In_632);
and U1988 (N_1988,In_2108,In_2462);
and U1989 (N_1989,In_334,In_1354);
nand U1990 (N_1990,In_281,In_2111);
or U1991 (N_1991,In_998,In_2957);
and U1992 (N_1992,In_1186,In_1192);
and U1993 (N_1993,In_331,In_2902);
nor U1994 (N_1994,In_215,In_334);
and U1995 (N_1995,In_2789,In_2067);
nand U1996 (N_1996,In_2908,In_1900);
or U1997 (N_1997,In_2413,In_1793);
xnor U1998 (N_1998,In_1720,In_2460);
or U1999 (N_1999,In_2780,In_216);
xor U2000 (N_2000,N_1368,N_339);
xnor U2001 (N_2001,N_633,N_1756);
nand U2002 (N_2002,N_406,N_1301);
and U2003 (N_2003,N_180,N_936);
and U2004 (N_2004,N_739,N_539);
or U2005 (N_2005,N_258,N_632);
or U2006 (N_2006,N_1440,N_660);
and U2007 (N_2007,N_404,N_1192);
xnor U2008 (N_2008,N_728,N_84);
xor U2009 (N_2009,N_1814,N_400);
xor U2010 (N_2010,N_1680,N_1429);
nor U2011 (N_2011,N_1097,N_336);
xnor U2012 (N_2012,N_1416,N_1057);
nor U2013 (N_2013,N_1553,N_668);
or U2014 (N_2014,N_1664,N_1707);
or U2015 (N_2015,N_1089,N_424);
nor U2016 (N_2016,N_118,N_1373);
xor U2017 (N_2017,N_1527,N_1919);
or U2018 (N_2018,N_691,N_1968);
xnor U2019 (N_2019,N_486,N_109);
and U2020 (N_2020,N_1980,N_1138);
nor U2021 (N_2021,N_412,N_1374);
nand U2022 (N_2022,N_452,N_387);
nand U2023 (N_2023,N_1034,N_549);
or U2024 (N_2024,N_1069,N_1472);
and U2025 (N_2025,N_781,N_1334);
and U2026 (N_2026,N_1582,N_927);
or U2027 (N_2027,N_815,N_498);
nor U2028 (N_2028,N_88,N_651);
xor U2029 (N_2029,N_1139,N_630);
nand U2030 (N_2030,N_1446,N_391);
nand U2031 (N_2031,N_475,N_300);
or U2032 (N_2032,N_1515,N_553);
or U2033 (N_2033,N_59,N_1130);
xor U2034 (N_2034,N_1335,N_1914);
nand U2035 (N_2035,N_35,N_1865);
nand U2036 (N_2036,N_908,N_352);
and U2037 (N_2037,N_1918,N_705);
nand U2038 (N_2038,N_717,N_996);
xnor U2039 (N_2039,N_1183,N_157);
or U2040 (N_2040,N_494,N_642);
and U2041 (N_2041,N_1890,N_1819);
and U2042 (N_2042,N_817,N_1381);
or U2043 (N_2043,N_69,N_1260);
nand U2044 (N_2044,N_1251,N_372);
and U2045 (N_2045,N_402,N_800);
nand U2046 (N_2046,N_145,N_1344);
nor U2047 (N_2047,N_1889,N_426);
nor U2048 (N_2048,N_445,N_1128);
nand U2049 (N_2049,N_945,N_1289);
and U2050 (N_2050,N_1888,N_499);
xnor U2051 (N_2051,N_286,N_86);
or U2052 (N_2052,N_467,N_1573);
or U2053 (N_2053,N_1233,N_461);
xor U2054 (N_2054,N_357,N_2);
nor U2055 (N_2055,N_1385,N_137);
and U2056 (N_2056,N_1551,N_281);
nor U2057 (N_2057,N_918,N_305);
xor U2058 (N_2058,N_1349,N_673);
xor U2059 (N_2059,N_1807,N_155);
nand U2060 (N_2060,N_704,N_291);
nand U2061 (N_2061,N_221,N_1786);
and U2062 (N_2062,N_360,N_1867);
nand U2063 (N_2063,N_1801,N_714);
xnor U2064 (N_2064,N_1592,N_287);
nor U2065 (N_2065,N_451,N_220);
xnor U2066 (N_2066,N_558,N_1279);
xnor U2067 (N_2067,N_1228,N_1875);
and U2068 (N_2068,N_480,N_1105);
or U2069 (N_2069,N_34,N_1015);
xnor U2070 (N_2070,N_677,N_359);
nand U2071 (N_2071,N_1578,N_1845);
nand U2072 (N_2072,N_179,N_1424);
nand U2073 (N_2073,N_1376,N_1896);
or U2074 (N_2074,N_1821,N_1148);
or U2075 (N_2075,N_1397,N_1058);
and U2076 (N_2076,N_1309,N_1943);
nor U2077 (N_2077,N_1156,N_1092);
or U2078 (N_2078,N_1250,N_909);
nor U2079 (N_2079,N_610,N_522);
xnor U2080 (N_2080,N_333,N_682);
xnor U2081 (N_2081,N_36,N_1455);
and U2082 (N_2082,N_1163,N_548);
and U2083 (N_2083,N_1957,N_1825);
or U2084 (N_2084,N_1784,N_485);
xor U2085 (N_2085,N_174,N_1616);
xnor U2086 (N_2086,N_363,N_1478);
xnor U2087 (N_2087,N_506,N_367);
and U2088 (N_2088,N_913,N_857);
xnor U2089 (N_2089,N_591,N_1731);
and U2090 (N_2090,N_1188,N_707);
nor U2091 (N_2091,N_310,N_314);
and U2092 (N_2092,N_955,N_1257);
nand U2093 (N_2093,N_1065,N_1240);
nor U2094 (N_2094,N_162,N_1283);
and U2095 (N_2095,N_1815,N_1569);
or U2096 (N_2096,N_809,N_1432);
xnor U2097 (N_2097,N_1848,N_1360);
or U2098 (N_2098,N_1362,N_1262);
nor U2099 (N_2099,N_659,N_460);
xor U2100 (N_2100,N_1215,N_1496);
nand U2101 (N_2101,N_628,N_82);
nand U2102 (N_2102,N_1259,N_415);
nand U2103 (N_2103,N_743,N_702);
and U2104 (N_2104,N_1874,N_1794);
nand U2105 (N_2105,N_738,N_319);
and U2106 (N_2106,N_1558,N_289);
nand U2107 (N_2107,N_184,N_75);
or U2108 (N_2108,N_520,N_940);
nor U2109 (N_2109,N_556,N_317);
or U2110 (N_2110,N_1217,N_55);
xor U2111 (N_2111,N_928,N_1161);
nand U2112 (N_2112,N_1605,N_1054);
or U2113 (N_2113,N_427,N_134);
nor U2114 (N_2114,N_330,N_1729);
and U2115 (N_2115,N_1641,N_1944);
or U2116 (N_2116,N_661,N_1282);
or U2117 (N_2117,N_1086,N_700);
nand U2118 (N_2118,N_599,N_1727);
nand U2119 (N_2119,N_1434,N_1333);
nor U2120 (N_2120,N_483,N_890);
and U2121 (N_2121,N_1849,N_1683);
and U2122 (N_2122,N_1532,N_1290);
nand U2123 (N_2123,N_51,N_422);
and U2124 (N_2124,N_441,N_1909);
nand U2125 (N_2125,N_1415,N_942);
nand U2126 (N_2126,N_850,N_1823);
xnor U2127 (N_2127,N_1467,N_1066);
xor U2128 (N_2128,N_311,N_253);
xnor U2129 (N_2129,N_583,N_361);
and U2130 (N_2130,N_1614,N_1631);
xor U2131 (N_2131,N_1886,N_1375);
nand U2132 (N_2132,N_303,N_1928);
xnor U2133 (N_2133,N_735,N_1642);
or U2134 (N_2134,N_1407,N_616);
nand U2135 (N_2135,N_1648,N_188);
nand U2136 (N_2136,N_77,N_897);
nand U2137 (N_2137,N_411,N_984);
or U2138 (N_2138,N_212,N_1760);
nand U2139 (N_2139,N_368,N_1880);
nand U2140 (N_2140,N_295,N_378);
and U2141 (N_2141,N_1911,N_48);
nand U2142 (N_2142,N_1678,N_1717);
nor U2143 (N_2143,N_876,N_1535);
nand U2144 (N_2144,N_256,N_1125);
or U2145 (N_2145,N_1091,N_41);
or U2146 (N_2146,N_560,N_1607);
xor U2147 (N_2147,N_1844,N_1639);
and U2148 (N_2148,N_933,N_95);
xor U2149 (N_2149,N_135,N_1857);
and U2150 (N_2150,N_237,N_1212);
nor U2151 (N_2151,N_623,N_1908);
nor U2152 (N_2152,N_1129,N_773);
or U2153 (N_2153,N_1358,N_67);
nand U2154 (N_2154,N_1094,N_294);
or U2155 (N_2155,N_1339,N_1820);
nor U2156 (N_2156,N_1140,N_1363);
and U2157 (N_2157,N_1056,N_248);
nand U2158 (N_2158,N_1953,N_1936);
and U2159 (N_2159,N_489,N_1107);
or U2160 (N_2160,N_1489,N_154);
nor U2161 (N_2161,N_730,N_1068);
nand U2162 (N_2162,N_1955,N_748);
or U2163 (N_2163,N_1136,N_686);
xnor U2164 (N_2164,N_986,N_1511);
or U2165 (N_2165,N_1394,N_1617);
nor U2166 (N_2166,N_1585,N_1754);
and U2167 (N_2167,N_566,N_1321);
nand U2168 (N_2168,N_1750,N_637);
or U2169 (N_2169,N_1554,N_1032);
and U2170 (N_2170,N_1546,N_1693);
xor U2171 (N_2171,N_1116,N_403);
or U2172 (N_2172,N_1995,N_1651);
or U2173 (N_2173,N_769,N_1555);
xor U2174 (N_2174,N_1121,N_1584);
nand U2175 (N_2175,N_584,N_24);
or U2176 (N_2176,N_1133,N_103);
nor U2177 (N_2177,N_1347,N_172);
or U2178 (N_2178,N_195,N_1197);
xnor U2179 (N_2179,N_196,N_123);
or U2180 (N_2180,N_143,N_471);
and U2181 (N_2181,N_1010,N_678);
and U2182 (N_2182,N_657,N_274);
or U2183 (N_2183,N_930,N_1304);
nand U2184 (N_2184,N_1146,N_1168);
xnor U2185 (N_2185,N_1508,N_1268);
nor U2186 (N_2186,N_1012,N_1808);
nand U2187 (N_2187,N_233,N_354);
and U2188 (N_2188,N_521,N_226);
and U2189 (N_2189,N_1882,N_1166);
nor U2190 (N_2190,N_852,N_569);
nand U2191 (N_2191,N_1493,N_316);
nand U2192 (N_2192,N_1529,N_146);
or U2193 (N_2193,N_901,N_1969);
xnor U2194 (N_2194,N_249,N_62);
nor U2195 (N_2195,N_1494,N_987);
or U2196 (N_2196,N_15,N_1594);
nor U2197 (N_2197,N_1462,N_371);
nand U2198 (N_2198,N_239,N_1236);
and U2199 (N_2199,N_52,N_1986);
or U2200 (N_2200,N_32,N_1803);
nand U2201 (N_2201,N_1587,N_1738);
and U2202 (N_2202,N_57,N_1414);
and U2203 (N_2203,N_667,N_1158);
or U2204 (N_2204,N_1719,N_1963);
or U2205 (N_2205,N_979,N_11);
xnor U2206 (N_2206,N_470,N_43);
or U2207 (N_2207,N_581,N_453);
or U2208 (N_2208,N_1650,N_429);
xor U2209 (N_2209,N_1281,N_1636);
or U2210 (N_2210,N_1959,N_1016);
nor U2211 (N_2211,N_1923,N_1436);
and U2212 (N_2212,N_243,N_73);
nand U2213 (N_2213,N_366,N_491);
nor U2214 (N_2214,N_210,N_1190);
nor U2215 (N_2215,N_1761,N_1187);
nor U2216 (N_2216,N_1061,N_1145);
and U2217 (N_2217,N_92,N_640);
xnor U2218 (N_2218,N_802,N_312);
and U2219 (N_2219,N_1070,N_1332);
or U2220 (N_2220,N_13,N_1448);
and U2221 (N_2221,N_978,N_690);
or U2222 (N_2222,N_956,N_1396);
nor U2223 (N_2223,N_1318,N_607);
and U2224 (N_2224,N_1829,N_1095);
xnor U2225 (N_2225,N_373,N_167);
xor U2226 (N_2226,N_457,N_1682);
nand U2227 (N_2227,N_1975,N_1755);
xnor U2228 (N_2228,N_1624,N_1903);
nand U2229 (N_2229,N_843,N_663);
and U2230 (N_2230,N_495,N_752);
and U2231 (N_2231,N_1470,N_1151);
nor U2232 (N_2232,N_1739,N_125);
xnor U2233 (N_2233,N_797,N_806);
nand U2234 (N_2234,N_1457,N_711);
xor U2235 (N_2235,N_329,N_688);
nand U2236 (N_2236,N_1476,N_302);
nand U2237 (N_2237,N_1430,N_621);
and U2238 (N_2238,N_418,N_1037);
nor U2239 (N_2239,N_1053,N_216);
xnor U2240 (N_2240,N_536,N_1380);
or U2241 (N_2241,N_1917,N_1169);
or U2242 (N_2242,N_594,N_207);
nand U2243 (N_2243,N_1996,N_428);
nand U2244 (N_2244,N_1479,N_1635);
nor U2245 (N_2245,N_1762,N_1830);
nor U2246 (N_2246,N_171,N_810);
and U2247 (N_2247,N_638,N_1818);
or U2248 (N_2248,N_1063,N_440);
nand U2249 (N_2249,N_1518,N_879);
and U2250 (N_2250,N_1506,N_1400);
nor U2251 (N_2251,N_511,N_1713);
nand U2252 (N_2252,N_1783,N_983);
xor U2253 (N_2253,N_723,N_1672);
or U2254 (N_2254,N_947,N_1714);
and U2255 (N_2255,N_1435,N_782);
or U2256 (N_2256,N_1954,N_247);
nor U2257 (N_2257,N_27,N_794);
xor U2258 (N_2258,N_296,N_726);
nand U2259 (N_2259,N_1547,N_1920);
and U2260 (N_2260,N_261,N_1938);
nor U2261 (N_2261,N_1926,N_318);
or U2262 (N_2262,N_1278,N_350);
xor U2263 (N_2263,N_1297,N_1777);
or U2264 (N_2264,N_679,N_1778);
nand U2265 (N_2265,N_1742,N_156);
or U2266 (N_2266,N_1202,N_1235);
and U2267 (N_2267,N_907,N_1442);
xnor U2268 (N_2268,N_148,N_1177);
and U2269 (N_2269,N_292,N_1203);
or U2270 (N_2270,N_1471,N_1602);
nor U2271 (N_2271,N_535,N_1676);
and U2272 (N_2272,N_606,N_78);
xnor U2273 (N_2273,N_1412,N_1483);
and U2274 (N_2274,N_20,N_1409);
xnor U2275 (N_2275,N_859,N_1871);
or U2276 (N_2276,N_1486,N_814);
xor U2277 (N_2277,N_653,N_1907);
and U2278 (N_2278,N_1073,N_1785);
or U2279 (N_2279,N_846,N_1542);
and U2280 (N_2280,N_1770,N_202);
or U2281 (N_2281,N_772,N_1469);
and U2282 (N_2282,N_444,N_1157);
and U2283 (N_2283,N_1463,N_746);
and U2284 (N_2284,N_1930,N_1219);
xor U2285 (N_2285,N_503,N_1437);
nand U2286 (N_2286,N_1843,N_513);
or U2287 (N_2287,N_775,N_1473);
xnor U2288 (N_2288,N_1565,N_505);
nor U2289 (N_2289,N_254,N_1295);
nand U2290 (N_2290,N_379,N_946);
nor U2291 (N_2291,N_1254,N_492);
or U2292 (N_2292,N_1323,N_1286);
nand U2293 (N_2293,N_789,N_425);
nand U2294 (N_2294,N_356,N_874);
nor U2295 (N_2295,N_873,N_1790);
xnor U2296 (N_2296,N_635,N_1405);
xnor U2297 (N_2297,N_793,N_484);
nand U2298 (N_2298,N_858,N_937);
or U2299 (N_2299,N_1544,N_523);
and U2300 (N_2300,N_1608,N_380);
nand U2301 (N_2301,N_463,N_1221);
or U2302 (N_2302,N_563,N_1662);
nor U2303 (N_2303,N_435,N_1458);
or U2304 (N_2304,N_515,N_525);
nand U2305 (N_2305,N_699,N_266);
xnor U2306 (N_2306,N_1491,N_217);
nor U2307 (N_2307,N_1255,N_1075);
xor U2308 (N_2308,N_910,N_1645);
nor U2309 (N_2309,N_693,N_629);
nor U2310 (N_2310,N_935,N_919);
xnor U2311 (N_2311,N_1669,N_115);
xnor U2312 (N_2312,N_1237,N_1973);
nor U2313 (N_2313,N_602,N_309);
or U2314 (N_2314,N_416,N_614);
and U2315 (N_2315,N_1025,N_4);
or U2316 (N_2316,N_1560,N_332);
and U2317 (N_2317,N_995,N_1866);
and U2318 (N_2318,N_1732,N_1293);
and U2319 (N_2319,N_374,N_218);
or U2320 (N_2320,N_1444,N_899);
nor U2321 (N_2321,N_1526,N_1868);
nor U2322 (N_2322,N_410,N_830);
and U2323 (N_2323,N_1269,N_1900);
nand U2324 (N_2324,N_1378,N_1985);
nor U2325 (N_2325,N_1700,N_1654);
or U2326 (N_2326,N_1740,N_792);
nor U2327 (N_2327,N_1023,N_1661);
nor U2328 (N_2328,N_455,N_744);
or U2329 (N_2329,N_1505,N_669);
or U2330 (N_2330,N_1466,N_962);
xor U2331 (N_2331,N_169,N_975);
nand U2332 (N_2332,N_1940,N_308);
nand U2333 (N_2333,N_617,N_341);
xor U2334 (N_2334,N_1816,N_119);
nand U2335 (N_2335,N_1083,N_532);
nor U2336 (N_2336,N_1305,N_764);
xor U2337 (N_2337,N_1118,N_1325);
nor U2338 (N_2338,N_1241,N_1031);
or U2339 (N_2339,N_1499,N_1313);
and U2340 (N_2340,N_1984,N_1795);
xnor U2341 (N_2341,N_293,N_1319);
or U2342 (N_2342,N_545,N_1595);
nand U2343 (N_2343,N_821,N_790);
or U2344 (N_2344,N_770,N_219);
nand U2345 (N_2345,N_1512,N_1836);
nor U2346 (N_2346,N_1388,N_687);
xnor U2347 (N_2347,N_664,N_238);
xnor U2348 (N_2348,N_141,N_1842);
or U2349 (N_2349,N_454,N_534);
and U2350 (N_2350,N_1913,N_299);
nand U2351 (N_2351,N_1165,N_884);
and U2352 (N_2352,N_1200,N_1813);
or U2353 (N_2353,N_527,N_1620);
xnor U2354 (N_2354,N_47,N_829);
xnor U2355 (N_2355,N_1119,N_662);
nand U2356 (N_2356,N_776,N_1861);
xor U2357 (N_2357,N_1899,N_241);
nor U2358 (N_2358,N_1947,N_1211);
nand U2359 (N_2359,N_1082,N_1581);
xnor U2360 (N_2360,N_1503,N_337);
nor U2361 (N_2361,N_1199,N_376);
and U2362 (N_2362,N_1220,N_1538);
or U2363 (N_2363,N_820,N_1482);
or U2364 (N_2364,N_959,N_952);
nand U2365 (N_2365,N_853,N_1422);
nand U2366 (N_2366,N_509,N_777);
nand U2367 (N_2367,N_554,N_1180);
and U2368 (N_2368,N_209,N_698);
nand U2369 (N_2369,N_1055,N_1663);
nand U2370 (N_2370,N_1431,N_1461);
or U2371 (N_2371,N_466,N_812);
and U2372 (N_2372,N_1310,N_459);
nor U2373 (N_2373,N_1675,N_1149);
and U2374 (N_2374,N_600,N_1697);
nor U2375 (N_2375,N_370,N_1441);
xor U2376 (N_2376,N_3,N_795);
and U2377 (N_2377,N_1967,N_1150);
or U2378 (N_2378,N_1364,N_868);
and U2379 (N_2379,N_1657,N_231);
nand U2380 (N_2380,N_279,N_1111);
nand U2381 (N_2381,N_784,N_1179);
nor U2382 (N_2382,N_160,N_1428);
xnor U2383 (N_2383,N_1285,N_17);
nand U2384 (N_2384,N_578,N_1401);
xnor U2385 (N_2385,N_165,N_1264);
nor U2386 (N_2386,N_383,N_1182);
nor U2387 (N_2387,N_1124,N_465);
nor U2388 (N_2388,N_131,N_759);
or U2389 (N_2389,N_298,N_1287);
nor U2390 (N_2390,N_903,N_758);
or U2391 (N_2391,N_1487,N_304);
or U2392 (N_2392,N_482,N_906);
and U2393 (N_2393,N_375,N_358);
or U2394 (N_2394,N_1921,N_215);
xnor U2395 (N_2395,N_1859,N_1225);
nor U2396 (N_2396,N_1501,N_1591);
xor U2397 (N_2397,N_883,N_1193);
nor U2398 (N_2398,N_19,N_1854);
and U2399 (N_2399,N_436,N_1178);
or U2400 (N_2400,N_587,N_273);
nor U2401 (N_2401,N_1314,N_1109);
nor U2402 (N_2402,N_823,N_963);
nor U2403 (N_2403,N_1846,N_774);
nand U2404 (N_2404,N_1632,N_533);
nand U2405 (N_2405,N_263,N_30);
nand U2406 (N_2406,N_706,N_1925);
xnor U2407 (N_2407,N_1725,N_328);
and U2408 (N_2408,N_631,N_33);
nand U2409 (N_2409,N_1348,N_865);
or U2410 (N_2410,N_1093,N_1113);
xnor U2411 (N_2411,N_228,N_559);
xor U2412 (N_2412,N_16,N_497);
and U2413 (N_2413,N_306,N_147);
xnor U2414 (N_2414,N_1391,N_976);
xor U2415 (N_2415,N_1634,N_1234);
nor U2416 (N_2416,N_1929,N_14);
or U2417 (N_2417,N_1637,N_127);
and U2418 (N_2418,N_1835,N_1361);
nor U2419 (N_2419,N_1311,N_122);
or U2420 (N_2420,N_66,N_742);
and U2421 (N_2421,N_502,N_285);
nor U2422 (N_2422,N_65,N_791);
xor U2423 (N_2423,N_1593,N_761);
nand U2424 (N_2424,N_129,N_1110);
xnor U2425 (N_2425,N_710,N_516);
or U2426 (N_2426,N_1191,N_1956);
nor U2427 (N_2427,N_992,N_501);
nor U2428 (N_2428,N_528,N_1209);
and U2429 (N_2429,N_271,N_282);
nor U2430 (N_2430,N_1852,N_1329);
or U2431 (N_2431,N_922,N_245);
nand U2432 (N_2432,N_163,N_120);
or U2433 (N_2433,N_1590,N_1002);
nand U2434 (N_2434,N_604,N_1020);
or U2435 (N_2435,N_1974,N_275);
xor U2436 (N_2436,N_1265,N_1989);
or U2437 (N_2437,N_1753,N_1809);
nor U2438 (N_2438,N_1049,N_1224);
and U2439 (N_2439,N_595,N_778);
xor U2440 (N_2440,N_1863,N_1768);
nor U2441 (N_2441,N_44,N_194);
nand U2442 (N_2442,N_684,N_665);
or U2443 (N_2443,N_1115,N_1284);
nor U2444 (N_2444,N_1744,N_1811);
or U2445 (N_2445,N_283,N_1336);
nand U2446 (N_2446,N_1822,N_1640);
or U2447 (N_2447,N_1271,N_1556);
xnor U2448 (N_2448,N_1978,N_654);
nor U2449 (N_2449,N_537,N_694);
and U2450 (N_2450,N_1689,N_697);
xnor U2451 (N_2451,N_1104,N_1074);
nor U2452 (N_2452,N_827,N_736);
or U2453 (N_2453,N_1858,N_1748);
or U2454 (N_2454,N_1189,N_1312);
nand U2455 (N_2455,N_818,N_93);
or U2456 (N_2456,N_618,N_1781);
nand U2457 (N_2457,N_1612,N_917);
xnor U2458 (N_2458,N_397,N_825);
and U2459 (N_2459,N_572,N_552);
and U2460 (N_2460,N_622,N_1733);
nand U2461 (N_2461,N_181,N_26);
xor U2462 (N_2462,N_1142,N_1393);
nand U2463 (N_2463,N_849,N_1379);
nor U2464 (N_2464,N_620,N_1688);
and U2465 (N_2465,N_1656,N_1942);
nor U2466 (N_2466,N_571,N_1681);
and U2467 (N_2467,N_964,N_544);
and U2468 (N_2468,N_994,N_948);
xnor U2469 (N_2469,N_1144,N_1447);
or U2470 (N_2470,N_1005,N_588);
and U2471 (N_2471,N_1004,N_567);
nor U2472 (N_2472,N_1009,N_1824);
or U2473 (N_2473,N_1665,N_1932);
nor U2474 (N_2474,N_1961,N_201);
and U2475 (N_2475,N_882,N_313);
nand U2476 (N_2476,N_1272,N_0);
or U2477 (N_2477,N_938,N_1543);
and U2478 (N_2478,N_1051,N_1952);
nor U2479 (N_2479,N_50,N_944);
nand U2480 (N_2480,N_1481,N_168);
or U2481 (N_2481,N_139,N_1143);
and U2482 (N_2482,N_1706,N_1991);
nor U2483 (N_2483,N_1915,N_68);
xor U2484 (N_2484,N_1999,N_1270);
nor U2485 (N_2485,N_187,N_1885);
xor U2486 (N_2486,N_108,N_639);
xor U2487 (N_2487,N_1047,N_993);
and U2488 (N_2488,N_347,N_1630);
and U2489 (N_2489,N_1222,N_1566);
nor U2490 (N_2490,N_763,N_1490);
and U2491 (N_2491,N_916,N_1988);
xnor U2492 (N_2492,N_1562,N_1112);
nand U2493 (N_2493,N_510,N_625);
nor U2494 (N_2494,N_58,N_999);
and U2495 (N_2495,N_720,N_439);
nor U2496 (N_2496,N_891,N_985);
nand U2497 (N_2497,N_1692,N_70);
xor U2498 (N_2498,N_1300,N_1606);
and U2499 (N_2499,N_1519,N_178);
or U2500 (N_2500,N_481,N_1048);
xnor U2501 (N_2501,N_1343,N_1668);
and U2502 (N_2502,N_323,N_1797);
nor U2503 (N_2503,N_284,N_1085);
nand U2504 (N_2504,N_1106,N_1879);
and U2505 (N_2505,N_242,N_112);
nor U2506 (N_2506,N_950,N_89);
nor U2507 (N_2507,N_1402,N_1998);
xnor U2508 (N_2508,N_1017,N_681);
xor U2509 (N_2509,N_493,N_246);
or U2510 (N_2510,N_838,N_980);
xnor U2511 (N_2511,N_974,N_340);
xor U2512 (N_2512,N_819,N_1579);
nand U2513 (N_2513,N_107,N_325);
or U2514 (N_2514,N_1710,N_685);
nand U2515 (N_2515,N_941,N_1759);
or U2516 (N_2516,N_177,N_365);
nand U2517 (N_2517,N_582,N_703);
nand U2518 (N_2518,N_478,N_1296);
and U2519 (N_2519,N_56,N_796);
xor U2520 (N_2520,N_1734,N_561);
xor U2521 (N_2521,N_531,N_701);
nand U2522 (N_2522,N_1084,N_331);
and U2523 (N_2523,N_1114,N_130);
xor U2524 (N_2524,N_1772,N_1767);
or U2525 (N_2525,N_1800,N_1045);
nand U2526 (N_2526,N_788,N_161);
xor U2527 (N_2527,N_40,N_12);
xor U2528 (N_2528,N_267,N_342);
nand U2529 (N_2529,N_1390,N_437);
or U2530 (N_2530,N_1477,N_176);
xnor U2531 (N_2531,N_116,N_1924);
and U2532 (N_2532,N_98,N_1367);
and U2533 (N_2533,N_970,N_613);
nand U2534 (N_2534,N_960,N_345);
or U2535 (N_2535,N_1480,N_1175);
nor U2536 (N_2536,N_450,N_786);
or U2537 (N_2537,N_878,N_716);
and U2538 (N_2538,N_1370,N_1052);
nand U2539 (N_2539,N_1077,N_551);
xnor U2540 (N_2540,N_1600,N_1653);
nor U2541 (N_2541,N_392,N_1044);
xor U2542 (N_2542,N_756,N_854);
and U2543 (N_2543,N_1103,N_264);
nor U2544 (N_2544,N_783,N_1937);
xor U2545 (N_2545,N_1667,N_1787);
nor U2546 (N_2546,N_1793,N_1099);
and U2547 (N_2547,N_364,N_1539);
or U2548 (N_2548,N_1522,N_1965);
xor U2549 (N_2549,N_1320,N_1029);
xor U2550 (N_2550,N_1395,N_1894);
nor U2551 (N_2551,N_1805,N_288);
and U2552 (N_2552,N_1315,N_1207);
xnor U2553 (N_2553,N_1966,N_1766);
xor U2554 (N_2554,N_722,N_1080);
xnor U2555 (N_2555,N_1331,N_1059);
xnor U2556 (N_2556,N_1013,N_1897);
nand U2557 (N_2557,N_327,N_1389);
nor U2558 (N_2558,N_1071,N_1531);
or U2559 (N_2559,N_1383,N_401);
or U2560 (N_2560,N_346,N_731);
and U2561 (N_2561,N_1036,N_1574);
nor U2562 (N_2562,N_1342,N_97);
xnor U2563 (N_2563,N_230,N_641);
xnor U2564 (N_2564,N_490,N_79);
or U2565 (N_2565,N_1060,N_1007);
and U2566 (N_2566,N_476,N_733);
nand U2567 (N_2567,N_1774,N_826);
nor U2568 (N_2568,N_85,N_320);
nor U2569 (N_2569,N_270,N_1377);
nor U2570 (N_2570,N_1873,N_1126);
nor U2571 (N_2571,N_1108,N_1652);
xnor U2572 (N_2572,N_1277,N_255);
xnor U2573 (N_2573,N_747,N_1701);
xor U2574 (N_2574,N_530,N_526);
xnor U2575 (N_2575,N_236,N_1619);
xor U2576 (N_2576,N_737,N_1239);
and U2577 (N_2577,N_1231,N_1540);
xor U2578 (N_2578,N_1242,N_46);
nor U2579 (N_2579,N_257,N_1001);
nand U2580 (N_2580,N_1746,N_1273);
nand U2581 (N_2581,N_53,N_954);
nand U2582 (N_2582,N_1771,N_1382);
xor U2583 (N_2583,N_1420,N_1575);
or U2584 (N_2584,N_1576,N_1981);
nor U2585 (N_2585,N_1887,N_557);
nand U2586 (N_2586,N_1757,N_902);
and U2587 (N_2587,N_1723,N_579);
xor U2588 (N_2588,N_822,N_496);
xnor U2589 (N_2589,N_1263,N_1213);
nand U2590 (N_2590,N_969,N_1521);
xnor U2591 (N_2591,N_1184,N_477);
nor U2592 (N_2592,N_517,N_816);
and U2593 (N_2593,N_1950,N_875);
or U2594 (N_2594,N_718,N_106);
nand U2595 (N_2595,N_1365,N_1043);
and U2596 (N_2596,N_1516,N_251);
and U2597 (N_2597,N_804,N_1100);
nand U2598 (N_2598,N_507,N_1328);
nor U2599 (N_2599,N_1498,N_1421);
nor U2600 (N_2600,N_1454,N_423);
or U2601 (N_2601,N_1838,N_1561);
or U2602 (N_2602,N_1724,N_1949);
nand U2603 (N_2603,N_1948,N_750);
and U2604 (N_2604,N_1703,N_1465);
nor U2605 (N_2605,N_1445,N_973);
nand U2606 (N_2606,N_807,N_626);
or U2607 (N_2607,N_1041,N_1618);
xnor U2608 (N_2608,N_1101,N_1715);
or U2609 (N_2609,N_421,N_1552);
and U2610 (N_2610,N_771,N_1524);
or U2611 (N_2611,N_898,N_856);
or U2612 (N_2612,N_1528,N_1167);
nor U2613 (N_2613,N_1704,N_923);
or U2614 (N_2614,N_1763,N_1514);
xor U2615 (N_2615,N_1643,N_183);
and U2616 (N_2616,N_1570,N_395);
or U2617 (N_2617,N_9,N_1638);
nand U2618 (N_2618,N_1970,N_464);
xnor U2619 (N_2619,N_1366,N_1351);
nand U2620 (N_2620,N_1147,N_223);
nand U2621 (N_2621,N_1997,N_634);
or U2622 (N_2622,N_647,N_334);
nand U2623 (N_2623,N_1317,N_1306);
nor U2624 (N_2624,N_596,N_1536);
or U2625 (N_2625,N_1684,N_1853);
and U2626 (N_2626,N_1679,N_666);
nor U2627 (N_2627,N_813,N_798);
nor U2628 (N_2628,N_197,N_568);
xor U2629 (N_2629,N_1982,N_719);
nand U2630 (N_2630,N_1904,N_1204);
nor U2631 (N_2631,N_1568,N_1090);
nand U2632 (N_2632,N_1851,N_1945);
or U2633 (N_2633,N_1610,N_96);
xor U2634 (N_2634,N_696,N_468);
nor U2635 (N_2635,N_965,N_780);
and U2636 (N_2636,N_1438,N_91);
and U2637 (N_2637,N_892,N_753);
and U2638 (N_2638,N_855,N_575);
nand U2639 (N_2639,N_1245,N_1525);
nor U2640 (N_2640,N_1609,N_593);
nand U2641 (N_2641,N_912,N_1398);
nand U2642 (N_2642,N_1971,N_1884);
nand U2643 (N_2643,N_1171,N_1788);
nor U2644 (N_2644,N_1403,N_1862);
nand U2645 (N_2645,N_1261,N_1384);
nand U2646 (N_2646,N_713,N_1789);
xor U2647 (N_2647,N_1201,N_1338);
or U2648 (N_2648,N_1721,N_1572);
and U2649 (N_2649,N_190,N_414);
or U2650 (N_2650,N_61,N_1230);
xnor U2651 (N_2651,N_222,N_1408);
or U2652 (N_2652,N_864,N_1992);
or U2653 (N_2653,N_1659,N_1509);
xor U2654 (N_2654,N_1356,N_904);
nor U2655 (N_2655,N_905,N_1916);
nand U2656 (N_2656,N_741,N_1452);
nor U2657 (N_2657,N_692,N_1559);
xor U2658 (N_2658,N_646,N_114);
xnor U2659 (N_2659,N_695,N_586);
and U2660 (N_2660,N_1951,N_205);
and U2661 (N_2661,N_1799,N_1337);
and U2662 (N_2662,N_1804,N_1122);
and U2663 (N_2663,N_1464,N_1252);
nand U2664 (N_2664,N_895,N_1743);
nand U2665 (N_2665,N_644,N_408);
xor U2666 (N_2666,N_991,N_1625);
xor U2667 (N_2667,N_1728,N_1502);
nor U2668 (N_2668,N_541,N_1810);
and U2669 (N_2669,N_1773,N_863);
or U2670 (N_2670,N_446,N_915);
or U2671 (N_2671,N_1979,N_871);
xnor U2672 (N_2672,N_225,N_1837);
xnor U2673 (N_2673,N_1628,N_1702);
nor U2674 (N_2674,N_911,N_683);
nor U2675 (N_2675,N_519,N_1695);
xor U2676 (N_2676,N_1993,N_624);
and U2677 (N_2677,N_1006,N_1577);
or U2678 (N_2678,N_322,N_803);
nor U2679 (N_2679,N_1855,N_344);
nand U2680 (N_2680,N_837,N_1883);
nand U2681 (N_2681,N_1686,N_1266);
nor U2682 (N_2682,N_348,N_1324);
nor U2683 (N_2683,N_1040,N_893);
nand U2684 (N_2684,N_204,N_1359);
xnor U2685 (N_2685,N_419,N_1500);
nor U2686 (N_2686,N_573,N_712);
nor U2687 (N_2687,N_1549,N_1330);
xor U2688 (N_2688,N_1340,N_1386);
nand U2689 (N_2689,N_1798,N_1155);
nand U2690 (N_2690,N_159,N_488);
nor U2691 (N_2691,N_1802,N_1453);
xnor U2692 (N_2692,N_1046,N_932);
nand U2693 (N_2693,N_619,N_627);
xnor U2694 (N_2694,N_1316,N_474);
and U2695 (N_2695,N_1162,N_1198);
and U2696 (N_2696,N_831,N_1537);
nand U2697 (N_2697,N_540,N_894);
or U2698 (N_2698,N_199,N_149);
xor U2699 (N_2699,N_872,N_1633);
nor U2700 (N_2700,N_757,N_1218);
nand U2701 (N_2701,N_1708,N_1698);
or U2702 (N_2702,N_870,N_1583);
xnor U2703 (N_2703,N_326,N_1655);
nand U2704 (N_2704,N_997,N_888);
xor U2705 (N_2705,N_39,N_500);
or U2706 (N_2706,N_151,N_555);
or U2707 (N_2707,N_656,N_1096);
nand U2708 (N_2708,N_866,N_113);
or U2709 (N_2709,N_60,N_1417);
or U2710 (N_2710,N_1550,N_1);
nor U2711 (N_2711,N_1404,N_650);
or U2712 (N_2712,N_472,N_1427);
nand U2713 (N_2713,N_1831,N_87);
xnor U2714 (N_2714,N_1244,N_1291);
nor U2715 (N_2715,N_836,N_1327);
and U2716 (N_2716,N_989,N_734);
nand U2717 (N_2717,N_252,N_94);
and U2718 (N_2718,N_432,N_721);
or U2719 (N_2719,N_1775,N_1039);
or U2720 (N_2720,N_232,N_643);
nor U2721 (N_2721,N_45,N_150);
nor U2722 (N_2722,N_234,N_645);
or U2723 (N_2723,N_981,N_1035);
nor U2724 (N_2724,N_1792,N_1749);
and U2725 (N_2725,N_1026,N_1922);
nand U2726 (N_2726,N_768,N_1716);
nand U2727 (N_2727,N_1423,N_349);
or U2728 (N_2728,N_386,N_1172);
nor U2729 (N_2729,N_1983,N_192);
nor U2730 (N_2730,N_1877,N_529);
nor U2731 (N_2731,N_968,N_1062);
and U2732 (N_2732,N_1079,N_745);
or U2733 (N_2733,N_988,N_1492);
and U2734 (N_2734,N_443,N_1302);
and U2735 (N_2735,N_1745,N_589);
nor U2736 (N_2736,N_351,N_1164);
nor U2737 (N_2737,N_74,N_766);
xnor U2738 (N_2738,N_1711,N_1275);
xnor U2739 (N_2739,N_1927,N_900);
xor U2740 (N_2740,N_1495,N_1050);
and U2741 (N_2741,N_1796,N_1604);
or U2742 (N_2742,N_1839,N_867);
xnor U2743 (N_2743,N_1134,N_240);
nand U2744 (N_2744,N_10,N_29);
and U2745 (N_2745,N_1972,N_1449);
nand U2746 (N_2746,N_362,N_133);
or U2747 (N_2747,N_1298,N_1072);
and U2748 (N_2748,N_268,N_929);
or U2749 (N_2749,N_1307,N_448);
xnor U2750 (N_2750,N_1274,N_538);
or U2751 (N_2751,N_23,N_877);
nor U2752 (N_2752,N_676,N_1229);
nor U2753 (N_2753,N_1850,N_887);
xor U2754 (N_2754,N_132,N_417);
nor U2755 (N_2755,N_1350,N_547);
nor U2756 (N_2756,N_1910,N_1864);
and U2757 (N_2757,N_1170,N_725);
and U2758 (N_2758,N_1000,N_1735);
and U2759 (N_2759,N_1253,N_111);
or U2760 (N_2760,N_652,N_430);
and U2761 (N_2761,N_1812,N_1308);
and U2762 (N_2762,N_1137,N_546);
nor U2763 (N_2763,N_449,N_1720);
nor U2764 (N_2764,N_724,N_1159);
xnor U2765 (N_2765,N_1934,N_104);
and U2766 (N_2766,N_1288,N_504);
nor U2767 (N_2767,N_229,N_1174);
xor U2768 (N_2768,N_206,N_708);
nand U2769 (N_2769,N_1737,N_508);
nand U2770 (N_2770,N_1598,N_262);
xor U2771 (N_2771,N_1677,N_689);
or U2772 (N_2772,N_1523,N_1078);
nand U2773 (N_2773,N_1439,N_749);
nand U2774 (N_2774,N_580,N_1008);
nand U2775 (N_2775,N_861,N_1280);
nor U2776 (N_2776,N_399,N_524);
and U2777 (N_2777,N_1673,N_512);
nor U2778 (N_2778,N_211,N_603);
and U2779 (N_2779,N_1497,N_381);
xnor U2780 (N_2780,N_1326,N_982);
or U2781 (N_2781,N_1410,N_570);
or U2782 (N_2782,N_958,N_1413);
or U2783 (N_2783,N_173,N_208);
or U2784 (N_2784,N_1102,N_250);
and U2785 (N_2785,N_835,N_153);
or U2786 (N_2786,N_1752,N_1765);
or U2787 (N_2787,N_1387,N_609);
or U2788 (N_2788,N_1699,N_715);
nor U2789 (N_2789,N_1747,N_1649);
nor U2790 (N_2790,N_597,N_844);
nand U2791 (N_2791,N_100,N_1195);
and U2792 (N_2792,N_1088,N_203);
and U2793 (N_2793,N_1418,N_1131);
or U2794 (N_2794,N_840,N_542);
xnor U2795 (N_2795,N_1893,N_473);
nor U2796 (N_2796,N_740,N_124);
nand U2797 (N_2797,N_420,N_83);
nor U2798 (N_2798,N_8,N_1226);
xor U2799 (N_2799,N_860,N_1019);
xnor U2800 (N_2800,N_1357,N_433);
xor U2801 (N_2801,N_76,N_138);
and U2802 (N_2802,N_21,N_31);
xor U2803 (N_2803,N_801,N_272);
or U2804 (N_2804,N_1902,N_1127);
nand U2805 (N_2805,N_200,N_998);
xnor U2806 (N_2806,N_833,N_369);
nor U2807 (N_2807,N_920,N_385);
nor U2808 (N_2808,N_1345,N_1042);
xor U2809 (N_2809,N_442,N_565);
xor U2810 (N_2810,N_396,N_479);
or U2811 (N_2811,N_462,N_1589);
and U2812 (N_2812,N_1120,N_81);
xor U2813 (N_2813,N_577,N_1644);
nand U2814 (N_2814,N_117,N_1488);
and U2815 (N_2815,N_1870,N_7);
or U2816 (N_2816,N_1028,N_1806);
nand U2817 (N_2817,N_611,N_1621);
xor U2818 (N_2818,N_355,N_343);
xnor U2819 (N_2819,N_834,N_1081);
xor U2820 (N_2820,N_63,N_1828);
xor U2821 (N_2821,N_280,N_805);
nor U2822 (N_2822,N_1826,N_1541);
nor U2823 (N_2823,N_1647,N_1303);
or U2824 (N_2824,N_1504,N_1994);
xnor U2825 (N_2825,N_880,N_1694);
nand U2826 (N_2826,N_787,N_658);
or U2827 (N_2827,N_128,N_1216);
and U2828 (N_2828,N_649,N_278);
xnor U2829 (N_2829,N_1726,N_808);
nand U2830 (N_2830,N_1834,N_1660);
and U2831 (N_2831,N_842,N_896);
nor U2832 (N_2832,N_1869,N_727);
or U2833 (N_2833,N_1906,N_214);
nor U2834 (N_2834,N_25,N_1256);
xor U2835 (N_2835,N_1856,N_72);
xnor U2836 (N_2836,N_1718,N_1827);
and U2837 (N_2837,N_269,N_1658);
nor U2838 (N_2838,N_1580,N_1817);
nor U2839 (N_2839,N_1205,N_1722);
and U2840 (N_2840,N_1214,N_1173);
or U2841 (N_2841,N_675,N_388);
and U2842 (N_2842,N_54,N_785);
nor U2843 (N_2843,N_1769,N_42);
xor U2844 (N_2844,N_514,N_1962);
or U2845 (N_2845,N_405,N_1484);
nand U2846 (N_2846,N_22,N_1931);
xor U2847 (N_2847,N_1258,N_90);
nand U2848 (N_2848,N_1782,N_1758);
xnor U2849 (N_2849,N_828,N_1027);
or U2850 (N_2850,N_943,N_175);
xnor U2851 (N_2851,N_1411,N_166);
and U2852 (N_2852,N_848,N_1346);
xor U2853 (N_2853,N_767,N_1841);
and U2854 (N_2854,N_1687,N_1987);
nor U2855 (N_2855,N_1459,N_1141);
nor U2856 (N_2856,N_1196,N_307);
xor U2857 (N_2857,N_576,N_1341);
xor U2858 (N_2858,N_99,N_1764);
or U2859 (N_2859,N_321,N_170);
nand U2860 (N_2860,N_394,N_198);
xor U2861 (N_2861,N_967,N_1712);
or U2862 (N_2862,N_1627,N_382);
xor U2863 (N_2863,N_924,N_18);
nor U2864 (N_2864,N_1603,N_680);
xnor U2865 (N_2865,N_1276,N_990);
nand U2866 (N_2866,N_1941,N_37);
nor U2867 (N_2867,N_71,N_1690);
xnor U2868 (N_2868,N_926,N_1990);
and U2869 (N_2869,N_732,N_1878);
and U2870 (N_2870,N_1791,N_1935);
nor U2871 (N_2871,N_1152,N_1014);
or U2872 (N_2872,N_839,N_1939);
nor U2873 (N_2873,N_1433,N_458);
or U2874 (N_2874,N_324,N_1881);
or U2875 (N_2875,N_949,N_765);
nand U2876 (N_2876,N_1033,N_564);
or U2877 (N_2877,N_762,N_1671);
nand U2878 (N_2878,N_961,N_1599);
xnor U2879 (N_2879,N_64,N_914);
and U2880 (N_2880,N_615,N_1905);
and U2881 (N_2881,N_1294,N_1468);
and U2882 (N_2882,N_921,N_1087);
nor U2883 (N_2883,N_1696,N_1751);
xnor U2884 (N_2884,N_1946,N_389);
xor U2885 (N_2885,N_1534,N_290);
or U2886 (N_2886,N_1003,N_1030);
and U2887 (N_2887,N_1369,N_1736);
or U2888 (N_2888,N_934,N_1530);
nand U2889 (N_2889,N_1451,N_189);
nand U2890 (N_2890,N_1776,N_939);
xor U2891 (N_2891,N_80,N_1067);
nor U2892 (N_2892,N_709,N_1517);
nor U2893 (N_2893,N_384,N_182);
and U2894 (N_2894,N_832,N_1232);
and U2895 (N_2895,N_885,N_1024);
xor U2896 (N_2896,N_672,N_953);
nand U2897 (N_2897,N_152,N_636);
nand U2898 (N_2898,N_1958,N_1135);
or U2899 (N_2899,N_1615,N_1022);
nand U2900 (N_2900,N_1507,N_841);
or U2901 (N_2901,N_977,N_1392);
xnor U2902 (N_2902,N_438,N_1613);
nor U2903 (N_2903,N_755,N_1450);
or U2904 (N_2904,N_1246,N_1705);
or U2905 (N_2905,N_1960,N_1545);
nor U2906 (N_2906,N_1194,N_1372);
or U2907 (N_2907,N_1186,N_121);
xor U2908 (N_2908,N_297,N_1685);
or U2909 (N_2909,N_487,N_315);
xnor U2910 (N_2910,N_1181,N_543);
nand U2911 (N_2911,N_518,N_1018);
nand U2912 (N_2912,N_413,N_398);
nand U2913 (N_2913,N_1176,N_1353);
and U2914 (N_2914,N_193,N_1741);
xor U2915 (N_2915,N_1596,N_1011);
nand U2916 (N_2916,N_972,N_862);
xor U2917 (N_2917,N_605,N_1563);
and U2918 (N_2918,N_1626,N_409);
or U2919 (N_2919,N_1588,N_957);
or U2920 (N_2920,N_136,N_1322);
or U2921 (N_2921,N_1629,N_1132);
nor U2922 (N_2922,N_1208,N_1406);
nor U2923 (N_2923,N_1860,N_1586);
nor U2924 (N_2924,N_1443,N_185);
nand U2925 (N_2925,N_671,N_1892);
or U2926 (N_2926,N_1601,N_1292);
nand U2927 (N_2927,N_1976,N_1898);
nor U2928 (N_2928,N_655,N_259);
nor U2929 (N_2929,N_1872,N_1267);
nand U2930 (N_2930,N_847,N_28);
nor U2931 (N_2931,N_648,N_1299);
and U2932 (N_2932,N_1038,N_335);
nor U2933 (N_2933,N_1419,N_754);
nor U2934 (N_2934,N_1249,N_760);
nand U2935 (N_2935,N_235,N_469);
nor U2936 (N_2936,N_1895,N_1426);
xnor U2937 (N_2937,N_1611,N_1622);
xnor U2938 (N_2938,N_390,N_353);
nand U2939 (N_2939,N_144,N_779);
and U2940 (N_2940,N_1227,N_102);
xnor U2941 (N_2941,N_1154,N_1354);
or U2942 (N_2942,N_1456,N_869);
nor U2943 (N_2943,N_1891,N_1533);
xor U2944 (N_2944,N_751,N_191);
nor U2945 (N_2945,N_550,N_601);
and U2946 (N_2946,N_1730,N_456);
nor U2947 (N_2947,N_1474,N_1425);
xnor U2948 (N_2948,N_1564,N_971);
nand U2949 (N_2949,N_1548,N_1243);
nand U2950 (N_2950,N_612,N_608);
nand U2951 (N_2951,N_1597,N_562);
nand U2952 (N_2952,N_1571,N_277);
or U2953 (N_2953,N_585,N_1355);
and U2954 (N_2954,N_1557,N_276);
nor U2955 (N_2955,N_1964,N_931);
nor U2956 (N_2956,N_1153,N_1210);
and U2957 (N_2957,N_1510,N_1238);
xnor U2958 (N_2958,N_1833,N_1912);
nand U2959 (N_2959,N_811,N_1666);
nor U2960 (N_2960,N_105,N_164);
and U2961 (N_2961,N_1670,N_38);
or U2962 (N_2962,N_1876,N_431);
nand U2963 (N_2963,N_824,N_598);
xor U2964 (N_2964,N_1223,N_140);
and U2965 (N_2965,N_447,N_265);
nand U2966 (N_2966,N_393,N_49);
xor U2967 (N_2967,N_1123,N_1185);
xnor U2968 (N_2968,N_377,N_886);
nand U2969 (N_2969,N_213,N_101);
nand U2970 (N_2970,N_1206,N_1709);
or U2971 (N_2971,N_1780,N_729);
or U2972 (N_2972,N_1160,N_1691);
nor U2973 (N_2973,N_260,N_110);
xor U2974 (N_2974,N_1977,N_1901);
nor U2975 (N_2975,N_1117,N_338);
or U2976 (N_2976,N_186,N_574);
nand U2977 (N_2977,N_881,N_1064);
xnor U2978 (N_2978,N_925,N_1475);
and U2979 (N_2979,N_590,N_889);
xor U2980 (N_2980,N_6,N_1840);
nand U2981 (N_2981,N_1520,N_851);
xnor U2982 (N_2982,N_1098,N_407);
nand U2983 (N_2983,N_1485,N_1933);
or U2984 (N_2984,N_126,N_1076);
and U2985 (N_2985,N_142,N_1371);
xor U2986 (N_2986,N_674,N_1847);
nor U2987 (N_2987,N_1832,N_1674);
xnor U2988 (N_2988,N_951,N_1248);
nand U2989 (N_2989,N_845,N_592);
or U2990 (N_2990,N_1399,N_1567);
and U2991 (N_2991,N_227,N_1513);
xor U2992 (N_2992,N_158,N_5);
or U2993 (N_2993,N_301,N_1021);
and U2994 (N_2994,N_670,N_1460);
or U2995 (N_2995,N_799,N_1646);
xor U2996 (N_2996,N_1352,N_1779);
or U2997 (N_2997,N_966,N_1247);
and U2998 (N_2998,N_244,N_434);
nor U2999 (N_2999,N_1623,N_224);
nand U3000 (N_3000,N_1620,N_114);
nand U3001 (N_3001,N_1772,N_534);
xor U3002 (N_3002,N_705,N_138);
nor U3003 (N_3003,N_69,N_30);
nor U3004 (N_3004,N_1002,N_1589);
or U3005 (N_3005,N_1544,N_544);
or U3006 (N_3006,N_553,N_792);
and U3007 (N_3007,N_1938,N_1671);
xnor U3008 (N_3008,N_1126,N_1563);
and U3009 (N_3009,N_1821,N_476);
and U3010 (N_3010,N_226,N_818);
xor U3011 (N_3011,N_964,N_19);
and U3012 (N_3012,N_12,N_417);
or U3013 (N_3013,N_810,N_745);
nand U3014 (N_3014,N_1758,N_972);
or U3015 (N_3015,N_897,N_1932);
or U3016 (N_3016,N_1944,N_1234);
nor U3017 (N_3017,N_33,N_1441);
nor U3018 (N_3018,N_1917,N_1645);
or U3019 (N_3019,N_1603,N_1933);
xor U3020 (N_3020,N_441,N_100);
xnor U3021 (N_3021,N_523,N_1898);
nor U3022 (N_3022,N_1685,N_1687);
and U3023 (N_3023,N_1376,N_1115);
or U3024 (N_3024,N_124,N_330);
or U3025 (N_3025,N_914,N_864);
nor U3026 (N_3026,N_381,N_582);
and U3027 (N_3027,N_122,N_727);
nor U3028 (N_3028,N_1920,N_1969);
xor U3029 (N_3029,N_368,N_205);
xnor U3030 (N_3030,N_1507,N_314);
and U3031 (N_3031,N_373,N_1267);
and U3032 (N_3032,N_236,N_1697);
nor U3033 (N_3033,N_1933,N_1126);
nand U3034 (N_3034,N_1569,N_318);
or U3035 (N_3035,N_803,N_1823);
nor U3036 (N_3036,N_1339,N_134);
nor U3037 (N_3037,N_1174,N_300);
nor U3038 (N_3038,N_1647,N_1609);
nor U3039 (N_3039,N_1558,N_1457);
nor U3040 (N_3040,N_1063,N_928);
nand U3041 (N_3041,N_490,N_63);
nand U3042 (N_3042,N_295,N_520);
xnor U3043 (N_3043,N_1696,N_613);
xor U3044 (N_3044,N_428,N_898);
and U3045 (N_3045,N_1188,N_1218);
or U3046 (N_3046,N_1525,N_280);
nand U3047 (N_3047,N_1141,N_675);
nor U3048 (N_3048,N_1892,N_605);
xor U3049 (N_3049,N_1236,N_166);
nor U3050 (N_3050,N_1088,N_137);
nand U3051 (N_3051,N_186,N_54);
or U3052 (N_3052,N_964,N_904);
and U3053 (N_3053,N_1910,N_19);
nand U3054 (N_3054,N_554,N_421);
or U3055 (N_3055,N_118,N_1461);
nor U3056 (N_3056,N_1945,N_887);
and U3057 (N_3057,N_963,N_389);
nand U3058 (N_3058,N_937,N_929);
nor U3059 (N_3059,N_309,N_248);
xnor U3060 (N_3060,N_450,N_57);
xnor U3061 (N_3061,N_1896,N_1426);
nand U3062 (N_3062,N_1111,N_837);
nand U3063 (N_3063,N_1347,N_1988);
and U3064 (N_3064,N_559,N_1090);
nand U3065 (N_3065,N_393,N_1741);
nor U3066 (N_3066,N_1071,N_1627);
or U3067 (N_3067,N_38,N_133);
or U3068 (N_3068,N_580,N_366);
nand U3069 (N_3069,N_1774,N_317);
and U3070 (N_3070,N_382,N_1288);
nor U3071 (N_3071,N_479,N_505);
nor U3072 (N_3072,N_1648,N_38);
nor U3073 (N_3073,N_1671,N_237);
xnor U3074 (N_3074,N_1653,N_121);
xor U3075 (N_3075,N_1192,N_1805);
xnor U3076 (N_3076,N_1115,N_1089);
nand U3077 (N_3077,N_163,N_1870);
nand U3078 (N_3078,N_500,N_638);
and U3079 (N_3079,N_1960,N_1018);
xor U3080 (N_3080,N_1702,N_1640);
nor U3081 (N_3081,N_1881,N_698);
xor U3082 (N_3082,N_305,N_908);
xor U3083 (N_3083,N_1327,N_1505);
and U3084 (N_3084,N_525,N_141);
xnor U3085 (N_3085,N_877,N_1172);
and U3086 (N_3086,N_72,N_1074);
xnor U3087 (N_3087,N_1412,N_1671);
xor U3088 (N_3088,N_1094,N_1062);
nor U3089 (N_3089,N_1064,N_1804);
xor U3090 (N_3090,N_1855,N_876);
and U3091 (N_3091,N_1834,N_1954);
xor U3092 (N_3092,N_781,N_1084);
and U3093 (N_3093,N_1521,N_1383);
xor U3094 (N_3094,N_1376,N_549);
or U3095 (N_3095,N_1643,N_881);
or U3096 (N_3096,N_1064,N_1154);
nor U3097 (N_3097,N_1507,N_1975);
or U3098 (N_3098,N_506,N_1316);
or U3099 (N_3099,N_289,N_1842);
xor U3100 (N_3100,N_273,N_56);
xnor U3101 (N_3101,N_1812,N_400);
nand U3102 (N_3102,N_1858,N_205);
nor U3103 (N_3103,N_171,N_176);
or U3104 (N_3104,N_391,N_915);
nor U3105 (N_3105,N_296,N_286);
and U3106 (N_3106,N_628,N_1641);
nor U3107 (N_3107,N_1743,N_1018);
nor U3108 (N_3108,N_131,N_1122);
or U3109 (N_3109,N_422,N_47);
and U3110 (N_3110,N_538,N_619);
nand U3111 (N_3111,N_48,N_384);
nor U3112 (N_3112,N_274,N_641);
xor U3113 (N_3113,N_718,N_188);
or U3114 (N_3114,N_1356,N_1998);
nand U3115 (N_3115,N_1463,N_1533);
nand U3116 (N_3116,N_297,N_1125);
xnor U3117 (N_3117,N_649,N_1269);
and U3118 (N_3118,N_1667,N_1755);
xor U3119 (N_3119,N_341,N_710);
xnor U3120 (N_3120,N_503,N_1766);
nor U3121 (N_3121,N_1916,N_133);
xnor U3122 (N_3122,N_302,N_1737);
xor U3123 (N_3123,N_1662,N_1012);
and U3124 (N_3124,N_504,N_1977);
and U3125 (N_3125,N_1387,N_369);
or U3126 (N_3126,N_371,N_1311);
xor U3127 (N_3127,N_1484,N_151);
nand U3128 (N_3128,N_1424,N_2);
xor U3129 (N_3129,N_1841,N_95);
and U3130 (N_3130,N_648,N_1250);
or U3131 (N_3131,N_1111,N_486);
nand U3132 (N_3132,N_1545,N_79);
and U3133 (N_3133,N_80,N_278);
and U3134 (N_3134,N_1458,N_1656);
nor U3135 (N_3135,N_1694,N_1403);
xor U3136 (N_3136,N_1881,N_120);
nor U3137 (N_3137,N_250,N_1139);
and U3138 (N_3138,N_140,N_1892);
nand U3139 (N_3139,N_397,N_883);
nand U3140 (N_3140,N_153,N_1913);
nor U3141 (N_3141,N_1738,N_240);
or U3142 (N_3142,N_857,N_1349);
and U3143 (N_3143,N_1159,N_1365);
or U3144 (N_3144,N_196,N_1422);
nand U3145 (N_3145,N_1597,N_772);
nor U3146 (N_3146,N_1535,N_918);
or U3147 (N_3147,N_135,N_1798);
or U3148 (N_3148,N_118,N_797);
xnor U3149 (N_3149,N_467,N_824);
and U3150 (N_3150,N_89,N_1317);
and U3151 (N_3151,N_652,N_807);
xnor U3152 (N_3152,N_1770,N_374);
nor U3153 (N_3153,N_1371,N_1404);
and U3154 (N_3154,N_1632,N_940);
or U3155 (N_3155,N_489,N_1446);
nor U3156 (N_3156,N_1666,N_916);
xnor U3157 (N_3157,N_1955,N_304);
nor U3158 (N_3158,N_1982,N_1204);
nor U3159 (N_3159,N_1431,N_952);
nor U3160 (N_3160,N_1216,N_278);
or U3161 (N_3161,N_1005,N_317);
nor U3162 (N_3162,N_760,N_1551);
nor U3163 (N_3163,N_1247,N_1285);
and U3164 (N_3164,N_1267,N_1656);
nor U3165 (N_3165,N_14,N_1472);
or U3166 (N_3166,N_418,N_1350);
and U3167 (N_3167,N_1235,N_1427);
or U3168 (N_3168,N_1553,N_1336);
or U3169 (N_3169,N_1447,N_1485);
nor U3170 (N_3170,N_1370,N_1760);
or U3171 (N_3171,N_246,N_145);
nand U3172 (N_3172,N_45,N_1030);
and U3173 (N_3173,N_1977,N_1076);
xor U3174 (N_3174,N_1749,N_569);
nor U3175 (N_3175,N_1333,N_962);
xnor U3176 (N_3176,N_709,N_144);
or U3177 (N_3177,N_1874,N_1740);
and U3178 (N_3178,N_999,N_1856);
or U3179 (N_3179,N_359,N_1340);
nand U3180 (N_3180,N_1684,N_408);
or U3181 (N_3181,N_534,N_285);
nor U3182 (N_3182,N_334,N_1478);
nor U3183 (N_3183,N_1508,N_37);
or U3184 (N_3184,N_328,N_570);
and U3185 (N_3185,N_965,N_1222);
xor U3186 (N_3186,N_774,N_1387);
nor U3187 (N_3187,N_650,N_72);
nor U3188 (N_3188,N_392,N_1924);
nand U3189 (N_3189,N_1701,N_404);
nand U3190 (N_3190,N_1928,N_1792);
nor U3191 (N_3191,N_71,N_1748);
nand U3192 (N_3192,N_1466,N_1526);
xor U3193 (N_3193,N_1681,N_1403);
or U3194 (N_3194,N_1541,N_226);
xnor U3195 (N_3195,N_753,N_1907);
and U3196 (N_3196,N_1227,N_351);
nor U3197 (N_3197,N_929,N_1256);
nand U3198 (N_3198,N_1532,N_1243);
nor U3199 (N_3199,N_846,N_274);
and U3200 (N_3200,N_1481,N_1666);
nor U3201 (N_3201,N_361,N_1165);
nor U3202 (N_3202,N_1959,N_1516);
nand U3203 (N_3203,N_671,N_1783);
xnor U3204 (N_3204,N_562,N_462);
and U3205 (N_3205,N_1488,N_1417);
and U3206 (N_3206,N_959,N_1698);
xor U3207 (N_3207,N_1366,N_528);
and U3208 (N_3208,N_161,N_1329);
xnor U3209 (N_3209,N_411,N_100);
nand U3210 (N_3210,N_361,N_763);
and U3211 (N_3211,N_1146,N_1283);
nor U3212 (N_3212,N_900,N_1021);
nand U3213 (N_3213,N_378,N_951);
and U3214 (N_3214,N_614,N_1228);
nor U3215 (N_3215,N_1938,N_1);
nand U3216 (N_3216,N_1476,N_727);
or U3217 (N_3217,N_109,N_909);
or U3218 (N_3218,N_181,N_125);
nor U3219 (N_3219,N_1445,N_320);
nand U3220 (N_3220,N_1599,N_834);
and U3221 (N_3221,N_1849,N_1748);
or U3222 (N_3222,N_200,N_1454);
and U3223 (N_3223,N_1976,N_663);
nor U3224 (N_3224,N_786,N_104);
xnor U3225 (N_3225,N_1657,N_1604);
xor U3226 (N_3226,N_1308,N_582);
or U3227 (N_3227,N_72,N_1659);
and U3228 (N_3228,N_1030,N_250);
or U3229 (N_3229,N_909,N_166);
nor U3230 (N_3230,N_752,N_1405);
and U3231 (N_3231,N_1635,N_1497);
nor U3232 (N_3232,N_1003,N_1851);
xnor U3233 (N_3233,N_363,N_970);
and U3234 (N_3234,N_1313,N_875);
nor U3235 (N_3235,N_455,N_1040);
nand U3236 (N_3236,N_925,N_1834);
xor U3237 (N_3237,N_103,N_1022);
xnor U3238 (N_3238,N_645,N_1433);
nand U3239 (N_3239,N_613,N_1014);
and U3240 (N_3240,N_1258,N_1363);
or U3241 (N_3241,N_667,N_161);
or U3242 (N_3242,N_168,N_1231);
or U3243 (N_3243,N_306,N_1452);
xor U3244 (N_3244,N_1142,N_1425);
or U3245 (N_3245,N_1628,N_371);
nor U3246 (N_3246,N_927,N_391);
xnor U3247 (N_3247,N_1134,N_675);
nand U3248 (N_3248,N_344,N_362);
xor U3249 (N_3249,N_310,N_911);
and U3250 (N_3250,N_251,N_72);
nand U3251 (N_3251,N_477,N_1390);
and U3252 (N_3252,N_629,N_1879);
nand U3253 (N_3253,N_1015,N_1227);
or U3254 (N_3254,N_781,N_559);
and U3255 (N_3255,N_734,N_779);
or U3256 (N_3256,N_1080,N_1883);
and U3257 (N_3257,N_387,N_964);
and U3258 (N_3258,N_1318,N_1949);
or U3259 (N_3259,N_597,N_976);
nand U3260 (N_3260,N_1100,N_1528);
xor U3261 (N_3261,N_118,N_1056);
and U3262 (N_3262,N_1945,N_1174);
and U3263 (N_3263,N_1001,N_1553);
or U3264 (N_3264,N_485,N_219);
xor U3265 (N_3265,N_1089,N_453);
or U3266 (N_3266,N_1139,N_5);
nor U3267 (N_3267,N_596,N_1746);
nand U3268 (N_3268,N_580,N_1518);
nand U3269 (N_3269,N_53,N_297);
xor U3270 (N_3270,N_1358,N_1429);
nand U3271 (N_3271,N_1652,N_1424);
nor U3272 (N_3272,N_1482,N_219);
and U3273 (N_3273,N_541,N_1957);
xor U3274 (N_3274,N_97,N_1124);
xor U3275 (N_3275,N_697,N_1652);
xor U3276 (N_3276,N_707,N_316);
nor U3277 (N_3277,N_1698,N_1571);
nor U3278 (N_3278,N_1981,N_194);
and U3279 (N_3279,N_634,N_287);
nand U3280 (N_3280,N_1240,N_440);
or U3281 (N_3281,N_592,N_1316);
nand U3282 (N_3282,N_1491,N_1271);
nor U3283 (N_3283,N_1548,N_186);
and U3284 (N_3284,N_643,N_1575);
xor U3285 (N_3285,N_1030,N_1141);
nand U3286 (N_3286,N_1345,N_238);
nor U3287 (N_3287,N_1993,N_1709);
xor U3288 (N_3288,N_266,N_897);
xnor U3289 (N_3289,N_710,N_915);
or U3290 (N_3290,N_1323,N_202);
xor U3291 (N_3291,N_1823,N_1043);
nor U3292 (N_3292,N_1250,N_564);
xnor U3293 (N_3293,N_1807,N_963);
nand U3294 (N_3294,N_1432,N_1164);
nor U3295 (N_3295,N_1793,N_466);
and U3296 (N_3296,N_1633,N_177);
nand U3297 (N_3297,N_1804,N_288);
and U3298 (N_3298,N_321,N_963);
nand U3299 (N_3299,N_1388,N_1215);
nor U3300 (N_3300,N_1625,N_505);
xor U3301 (N_3301,N_377,N_1222);
or U3302 (N_3302,N_1401,N_714);
or U3303 (N_3303,N_1825,N_678);
nor U3304 (N_3304,N_1462,N_1873);
and U3305 (N_3305,N_1413,N_1379);
xor U3306 (N_3306,N_1784,N_102);
nor U3307 (N_3307,N_1618,N_1408);
nand U3308 (N_3308,N_1164,N_1316);
nand U3309 (N_3309,N_1110,N_357);
nand U3310 (N_3310,N_759,N_1305);
xor U3311 (N_3311,N_539,N_1708);
and U3312 (N_3312,N_119,N_593);
nor U3313 (N_3313,N_439,N_40);
and U3314 (N_3314,N_1755,N_1720);
nand U3315 (N_3315,N_1539,N_455);
xor U3316 (N_3316,N_1868,N_218);
xnor U3317 (N_3317,N_968,N_1037);
xor U3318 (N_3318,N_1944,N_1634);
and U3319 (N_3319,N_885,N_1878);
nor U3320 (N_3320,N_921,N_1948);
or U3321 (N_3321,N_244,N_1557);
and U3322 (N_3322,N_184,N_1781);
or U3323 (N_3323,N_840,N_74);
nor U3324 (N_3324,N_303,N_1985);
nand U3325 (N_3325,N_1664,N_587);
nor U3326 (N_3326,N_580,N_1043);
or U3327 (N_3327,N_1547,N_300);
xor U3328 (N_3328,N_1265,N_1214);
or U3329 (N_3329,N_1951,N_1313);
nand U3330 (N_3330,N_1870,N_1486);
xor U3331 (N_3331,N_965,N_1198);
nor U3332 (N_3332,N_190,N_1548);
and U3333 (N_3333,N_194,N_119);
xnor U3334 (N_3334,N_661,N_1113);
nor U3335 (N_3335,N_314,N_347);
nor U3336 (N_3336,N_289,N_1778);
and U3337 (N_3337,N_1529,N_271);
or U3338 (N_3338,N_1489,N_922);
or U3339 (N_3339,N_1489,N_1329);
or U3340 (N_3340,N_731,N_1392);
xnor U3341 (N_3341,N_1171,N_493);
nand U3342 (N_3342,N_385,N_543);
nand U3343 (N_3343,N_677,N_80);
xor U3344 (N_3344,N_1825,N_1820);
and U3345 (N_3345,N_1327,N_72);
xor U3346 (N_3346,N_698,N_1252);
xor U3347 (N_3347,N_1032,N_103);
nand U3348 (N_3348,N_159,N_117);
xnor U3349 (N_3349,N_108,N_1403);
and U3350 (N_3350,N_744,N_546);
and U3351 (N_3351,N_463,N_1272);
and U3352 (N_3352,N_316,N_502);
or U3353 (N_3353,N_1836,N_1869);
nand U3354 (N_3354,N_1796,N_385);
nand U3355 (N_3355,N_1906,N_400);
xor U3356 (N_3356,N_948,N_369);
nor U3357 (N_3357,N_1806,N_165);
or U3358 (N_3358,N_1738,N_1705);
xnor U3359 (N_3359,N_304,N_168);
or U3360 (N_3360,N_1465,N_542);
nor U3361 (N_3361,N_354,N_393);
xor U3362 (N_3362,N_1490,N_1345);
nor U3363 (N_3363,N_1581,N_1064);
and U3364 (N_3364,N_1499,N_1564);
or U3365 (N_3365,N_1367,N_1602);
xnor U3366 (N_3366,N_1365,N_1063);
nand U3367 (N_3367,N_530,N_1659);
nor U3368 (N_3368,N_767,N_1383);
and U3369 (N_3369,N_1287,N_1854);
nand U3370 (N_3370,N_1946,N_137);
nand U3371 (N_3371,N_489,N_1578);
xnor U3372 (N_3372,N_1973,N_156);
nand U3373 (N_3373,N_1336,N_1769);
nand U3374 (N_3374,N_1919,N_656);
nor U3375 (N_3375,N_1610,N_1511);
nor U3376 (N_3376,N_562,N_1836);
nor U3377 (N_3377,N_1087,N_605);
or U3378 (N_3378,N_1721,N_1531);
nor U3379 (N_3379,N_409,N_463);
nor U3380 (N_3380,N_977,N_1383);
nor U3381 (N_3381,N_840,N_1440);
nand U3382 (N_3382,N_880,N_270);
or U3383 (N_3383,N_450,N_1662);
nand U3384 (N_3384,N_869,N_1192);
or U3385 (N_3385,N_390,N_655);
or U3386 (N_3386,N_1472,N_657);
xnor U3387 (N_3387,N_34,N_559);
xnor U3388 (N_3388,N_108,N_584);
xor U3389 (N_3389,N_1223,N_102);
and U3390 (N_3390,N_1935,N_1802);
or U3391 (N_3391,N_321,N_157);
nand U3392 (N_3392,N_1825,N_264);
nand U3393 (N_3393,N_775,N_591);
nand U3394 (N_3394,N_520,N_832);
xor U3395 (N_3395,N_1219,N_1762);
xnor U3396 (N_3396,N_1057,N_1210);
and U3397 (N_3397,N_1351,N_1131);
and U3398 (N_3398,N_796,N_1803);
and U3399 (N_3399,N_245,N_626);
nand U3400 (N_3400,N_1475,N_352);
nor U3401 (N_3401,N_1259,N_1237);
xnor U3402 (N_3402,N_1025,N_1000);
nand U3403 (N_3403,N_1150,N_489);
xor U3404 (N_3404,N_1376,N_1413);
or U3405 (N_3405,N_1638,N_1421);
xor U3406 (N_3406,N_1552,N_1385);
xnor U3407 (N_3407,N_87,N_1105);
nand U3408 (N_3408,N_1352,N_1694);
nand U3409 (N_3409,N_1794,N_949);
xnor U3410 (N_3410,N_966,N_388);
or U3411 (N_3411,N_921,N_664);
or U3412 (N_3412,N_1108,N_1121);
or U3413 (N_3413,N_94,N_183);
nand U3414 (N_3414,N_1105,N_103);
or U3415 (N_3415,N_1894,N_1940);
nand U3416 (N_3416,N_1732,N_1932);
and U3417 (N_3417,N_706,N_1020);
or U3418 (N_3418,N_361,N_768);
nor U3419 (N_3419,N_754,N_387);
nand U3420 (N_3420,N_1626,N_42);
xor U3421 (N_3421,N_1122,N_612);
nand U3422 (N_3422,N_1339,N_1064);
xor U3423 (N_3423,N_169,N_1636);
and U3424 (N_3424,N_961,N_635);
xor U3425 (N_3425,N_487,N_547);
nand U3426 (N_3426,N_1647,N_1393);
xor U3427 (N_3427,N_1998,N_721);
xnor U3428 (N_3428,N_86,N_1087);
or U3429 (N_3429,N_424,N_1418);
nand U3430 (N_3430,N_463,N_1373);
nor U3431 (N_3431,N_13,N_968);
xnor U3432 (N_3432,N_1869,N_1816);
xnor U3433 (N_3433,N_1272,N_546);
or U3434 (N_3434,N_860,N_1389);
xnor U3435 (N_3435,N_1867,N_1604);
nand U3436 (N_3436,N_1393,N_1606);
xor U3437 (N_3437,N_810,N_1324);
nor U3438 (N_3438,N_767,N_1204);
xor U3439 (N_3439,N_931,N_874);
or U3440 (N_3440,N_1511,N_1645);
nand U3441 (N_3441,N_1136,N_233);
nand U3442 (N_3442,N_1399,N_357);
nor U3443 (N_3443,N_1873,N_620);
nand U3444 (N_3444,N_30,N_1841);
nor U3445 (N_3445,N_1591,N_1269);
nor U3446 (N_3446,N_863,N_1457);
nand U3447 (N_3447,N_439,N_621);
and U3448 (N_3448,N_1343,N_1040);
nor U3449 (N_3449,N_1160,N_318);
nor U3450 (N_3450,N_746,N_356);
nand U3451 (N_3451,N_1657,N_611);
and U3452 (N_3452,N_1359,N_1796);
and U3453 (N_3453,N_785,N_1069);
xnor U3454 (N_3454,N_790,N_1307);
nand U3455 (N_3455,N_1143,N_1592);
and U3456 (N_3456,N_696,N_1071);
xor U3457 (N_3457,N_1629,N_1001);
or U3458 (N_3458,N_1021,N_720);
xor U3459 (N_3459,N_1370,N_1201);
xnor U3460 (N_3460,N_946,N_500);
nor U3461 (N_3461,N_1679,N_1017);
xor U3462 (N_3462,N_178,N_1843);
nor U3463 (N_3463,N_266,N_1890);
and U3464 (N_3464,N_1310,N_1204);
xnor U3465 (N_3465,N_125,N_1319);
or U3466 (N_3466,N_212,N_1195);
nand U3467 (N_3467,N_623,N_987);
and U3468 (N_3468,N_474,N_1972);
nor U3469 (N_3469,N_795,N_109);
nand U3470 (N_3470,N_960,N_1294);
or U3471 (N_3471,N_1851,N_1193);
nor U3472 (N_3472,N_266,N_666);
nor U3473 (N_3473,N_796,N_1256);
nand U3474 (N_3474,N_674,N_167);
xnor U3475 (N_3475,N_169,N_1515);
nand U3476 (N_3476,N_532,N_973);
xnor U3477 (N_3477,N_1071,N_1564);
xor U3478 (N_3478,N_557,N_115);
and U3479 (N_3479,N_858,N_1345);
and U3480 (N_3480,N_1571,N_991);
nor U3481 (N_3481,N_503,N_707);
and U3482 (N_3482,N_723,N_1480);
and U3483 (N_3483,N_1503,N_459);
or U3484 (N_3484,N_545,N_36);
or U3485 (N_3485,N_1596,N_1518);
nor U3486 (N_3486,N_1711,N_1372);
nand U3487 (N_3487,N_1282,N_1173);
nor U3488 (N_3488,N_547,N_314);
nor U3489 (N_3489,N_421,N_957);
nor U3490 (N_3490,N_1387,N_1950);
and U3491 (N_3491,N_742,N_1785);
xnor U3492 (N_3492,N_177,N_689);
and U3493 (N_3493,N_1392,N_1757);
and U3494 (N_3494,N_1652,N_729);
nand U3495 (N_3495,N_1255,N_885);
nand U3496 (N_3496,N_231,N_991);
nor U3497 (N_3497,N_687,N_1147);
nor U3498 (N_3498,N_1410,N_1931);
nand U3499 (N_3499,N_1659,N_1491);
xnor U3500 (N_3500,N_1296,N_1746);
nand U3501 (N_3501,N_915,N_723);
nor U3502 (N_3502,N_1328,N_1643);
nand U3503 (N_3503,N_903,N_1786);
and U3504 (N_3504,N_931,N_677);
and U3505 (N_3505,N_1593,N_1706);
nand U3506 (N_3506,N_1946,N_642);
nor U3507 (N_3507,N_1773,N_1519);
and U3508 (N_3508,N_797,N_1146);
and U3509 (N_3509,N_640,N_863);
xnor U3510 (N_3510,N_1282,N_1775);
xor U3511 (N_3511,N_873,N_821);
or U3512 (N_3512,N_644,N_911);
and U3513 (N_3513,N_1186,N_506);
nand U3514 (N_3514,N_491,N_1591);
or U3515 (N_3515,N_1355,N_722);
nor U3516 (N_3516,N_962,N_1857);
xor U3517 (N_3517,N_1872,N_1996);
and U3518 (N_3518,N_225,N_1550);
nand U3519 (N_3519,N_1227,N_1652);
nand U3520 (N_3520,N_1260,N_158);
or U3521 (N_3521,N_811,N_1736);
nand U3522 (N_3522,N_117,N_1876);
and U3523 (N_3523,N_1937,N_1326);
xnor U3524 (N_3524,N_1387,N_353);
and U3525 (N_3525,N_1792,N_994);
or U3526 (N_3526,N_198,N_1322);
xor U3527 (N_3527,N_1051,N_82);
and U3528 (N_3528,N_183,N_194);
xor U3529 (N_3529,N_1747,N_866);
xnor U3530 (N_3530,N_1937,N_1704);
xnor U3531 (N_3531,N_322,N_270);
and U3532 (N_3532,N_1385,N_932);
and U3533 (N_3533,N_957,N_1733);
nor U3534 (N_3534,N_343,N_1284);
or U3535 (N_3535,N_826,N_1047);
nor U3536 (N_3536,N_1357,N_749);
or U3537 (N_3537,N_1264,N_1904);
and U3538 (N_3538,N_679,N_1578);
xnor U3539 (N_3539,N_1790,N_401);
nor U3540 (N_3540,N_93,N_690);
xnor U3541 (N_3541,N_1946,N_440);
and U3542 (N_3542,N_1776,N_172);
and U3543 (N_3543,N_1595,N_234);
nor U3544 (N_3544,N_1321,N_1831);
and U3545 (N_3545,N_1071,N_1604);
or U3546 (N_3546,N_1693,N_855);
or U3547 (N_3547,N_1818,N_1588);
or U3548 (N_3548,N_39,N_555);
nand U3549 (N_3549,N_63,N_1116);
and U3550 (N_3550,N_1475,N_11);
or U3551 (N_3551,N_1794,N_39);
nand U3552 (N_3552,N_561,N_584);
xor U3553 (N_3553,N_1313,N_593);
nor U3554 (N_3554,N_1042,N_870);
nor U3555 (N_3555,N_1673,N_916);
and U3556 (N_3556,N_888,N_1141);
nor U3557 (N_3557,N_709,N_341);
or U3558 (N_3558,N_1898,N_1505);
xor U3559 (N_3559,N_637,N_479);
xnor U3560 (N_3560,N_1094,N_1441);
and U3561 (N_3561,N_1729,N_1579);
or U3562 (N_3562,N_1428,N_1686);
nor U3563 (N_3563,N_191,N_993);
xor U3564 (N_3564,N_860,N_1269);
nor U3565 (N_3565,N_852,N_1805);
nand U3566 (N_3566,N_1615,N_424);
and U3567 (N_3567,N_1872,N_1051);
or U3568 (N_3568,N_1636,N_1003);
and U3569 (N_3569,N_894,N_905);
nor U3570 (N_3570,N_532,N_10);
or U3571 (N_3571,N_1418,N_1834);
nor U3572 (N_3572,N_418,N_1569);
or U3573 (N_3573,N_1269,N_737);
xor U3574 (N_3574,N_1159,N_1050);
or U3575 (N_3575,N_558,N_1014);
xor U3576 (N_3576,N_154,N_401);
or U3577 (N_3577,N_252,N_1974);
nand U3578 (N_3578,N_660,N_9);
xor U3579 (N_3579,N_1513,N_174);
xor U3580 (N_3580,N_1016,N_707);
xor U3581 (N_3581,N_413,N_377);
or U3582 (N_3582,N_700,N_440);
or U3583 (N_3583,N_1076,N_631);
nor U3584 (N_3584,N_523,N_1004);
xnor U3585 (N_3585,N_1142,N_1073);
or U3586 (N_3586,N_60,N_1659);
and U3587 (N_3587,N_798,N_487);
nand U3588 (N_3588,N_604,N_1384);
nor U3589 (N_3589,N_320,N_234);
nand U3590 (N_3590,N_507,N_268);
nand U3591 (N_3591,N_1501,N_934);
and U3592 (N_3592,N_214,N_29);
nor U3593 (N_3593,N_1476,N_853);
xnor U3594 (N_3594,N_609,N_280);
or U3595 (N_3595,N_631,N_1053);
nand U3596 (N_3596,N_83,N_581);
xor U3597 (N_3597,N_564,N_1961);
nand U3598 (N_3598,N_296,N_310);
and U3599 (N_3599,N_1080,N_1974);
or U3600 (N_3600,N_211,N_1984);
xor U3601 (N_3601,N_1980,N_893);
and U3602 (N_3602,N_1975,N_1059);
and U3603 (N_3603,N_1362,N_1302);
or U3604 (N_3604,N_1889,N_368);
xnor U3605 (N_3605,N_719,N_504);
nor U3606 (N_3606,N_1579,N_307);
nand U3607 (N_3607,N_1594,N_643);
xor U3608 (N_3608,N_931,N_1317);
nand U3609 (N_3609,N_124,N_1313);
nand U3610 (N_3610,N_1563,N_417);
xnor U3611 (N_3611,N_1239,N_997);
nor U3612 (N_3612,N_597,N_216);
and U3613 (N_3613,N_1425,N_1189);
nand U3614 (N_3614,N_1879,N_256);
or U3615 (N_3615,N_1292,N_462);
nand U3616 (N_3616,N_271,N_283);
xor U3617 (N_3617,N_364,N_1332);
nand U3618 (N_3618,N_981,N_1071);
nand U3619 (N_3619,N_537,N_214);
xor U3620 (N_3620,N_182,N_891);
xor U3621 (N_3621,N_709,N_1856);
or U3622 (N_3622,N_1800,N_559);
or U3623 (N_3623,N_1155,N_1018);
xnor U3624 (N_3624,N_161,N_99);
or U3625 (N_3625,N_679,N_323);
and U3626 (N_3626,N_610,N_1549);
or U3627 (N_3627,N_154,N_83);
nand U3628 (N_3628,N_431,N_1885);
nand U3629 (N_3629,N_1548,N_102);
and U3630 (N_3630,N_183,N_1225);
and U3631 (N_3631,N_1862,N_763);
nor U3632 (N_3632,N_1910,N_780);
nor U3633 (N_3633,N_1658,N_1797);
xor U3634 (N_3634,N_927,N_580);
nor U3635 (N_3635,N_1006,N_729);
nand U3636 (N_3636,N_845,N_223);
nor U3637 (N_3637,N_73,N_1247);
nand U3638 (N_3638,N_1289,N_1864);
nand U3639 (N_3639,N_791,N_1044);
nand U3640 (N_3640,N_253,N_458);
and U3641 (N_3641,N_1267,N_255);
and U3642 (N_3642,N_415,N_1860);
nand U3643 (N_3643,N_1292,N_1403);
xnor U3644 (N_3644,N_100,N_1713);
or U3645 (N_3645,N_355,N_1281);
or U3646 (N_3646,N_1973,N_842);
nand U3647 (N_3647,N_1967,N_1002);
nand U3648 (N_3648,N_1479,N_261);
nand U3649 (N_3649,N_1890,N_1290);
and U3650 (N_3650,N_1675,N_79);
xor U3651 (N_3651,N_1480,N_786);
xnor U3652 (N_3652,N_1136,N_759);
nor U3653 (N_3653,N_1108,N_1805);
and U3654 (N_3654,N_1849,N_1864);
nor U3655 (N_3655,N_1111,N_132);
and U3656 (N_3656,N_544,N_659);
and U3657 (N_3657,N_1021,N_1409);
nand U3658 (N_3658,N_988,N_299);
and U3659 (N_3659,N_822,N_468);
nand U3660 (N_3660,N_6,N_1993);
or U3661 (N_3661,N_973,N_1816);
or U3662 (N_3662,N_561,N_656);
xnor U3663 (N_3663,N_1179,N_1198);
or U3664 (N_3664,N_625,N_1499);
nor U3665 (N_3665,N_261,N_418);
and U3666 (N_3666,N_1753,N_1091);
xor U3667 (N_3667,N_319,N_306);
nor U3668 (N_3668,N_1867,N_1120);
or U3669 (N_3669,N_824,N_1044);
or U3670 (N_3670,N_1460,N_1902);
and U3671 (N_3671,N_155,N_1788);
or U3672 (N_3672,N_315,N_548);
xor U3673 (N_3673,N_1957,N_508);
xnor U3674 (N_3674,N_588,N_1534);
nor U3675 (N_3675,N_1406,N_570);
xor U3676 (N_3676,N_1936,N_576);
xnor U3677 (N_3677,N_1117,N_1239);
nor U3678 (N_3678,N_660,N_929);
xnor U3679 (N_3679,N_1482,N_1313);
and U3680 (N_3680,N_663,N_1826);
nor U3681 (N_3681,N_1208,N_150);
xnor U3682 (N_3682,N_1943,N_929);
or U3683 (N_3683,N_952,N_1053);
nor U3684 (N_3684,N_1046,N_1712);
or U3685 (N_3685,N_1198,N_656);
or U3686 (N_3686,N_1437,N_272);
nand U3687 (N_3687,N_1335,N_1828);
nor U3688 (N_3688,N_1453,N_1147);
nor U3689 (N_3689,N_30,N_473);
nand U3690 (N_3690,N_1201,N_435);
nand U3691 (N_3691,N_831,N_263);
nor U3692 (N_3692,N_1649,N_235);
and U3693 (N_3693,N_1366,N_1769);
and U3694 (N_3694,N_592,N_848);
xnor U3695 (N_3695,N_1992,N_501);
nor U3696 (N_3696,N_1616,N_219);
nor U3697 (N_3697,N_765,N_1268);
and U3698 (N_3698,N_1814,N_27);
nand U3699 (N_3699,N_759,N_1731);
nand U3700 (N_3700,N_1207,N_362);
nor U3701 (N_3701,N_1199,N_1319);
or U3702 (N_3702,N_1716,N_1710);
xor U3703 (N_3703,N_1183,N_543);
nor U3704 (N_3704,N_1763,N_781);
or U3705 (N_3705,N_1393,N_1030);
xor U3706 (N_3706,N_1674,N_915);
xnor U3707 (N_3707,N_628,N_1405);
nor U3708 (N_3708,N_1169,N_1932);
nand U3709 (N_3709,N_1826,N_943);
nand U3710 (N_3710,N_1704,N_566);
nand U3711 (N_3711,N_1927,N_296);
nand U3712 (N_3712,N_963,N_1666);
or U3713 (N_3713,N_1324,N_1366);
or U3714 (N_3714,N_1134,N_1033);
nand U3715 (N_3715,N_563,N_1136);
nor U3716 (N_3716,N_78,N_112);
nor U3717 (N_3717,N_52,N_824);
xnor U3718 (N_3718,N_694,N_284);
or U3719 (N_3719,N_1193,N_220);
xor U3720 (N_3720,N_1861,N_1637);
or U3721 (N_3721,N_1159,N_800);
xor U3722 (N_3722,N_1690,N_617);
and U3723 (N_3723,N_676,N_586);
nand U3724 (N_3724,N_1369,N_383);
and U3725 (N_3725,N_458,N_1498);
and U3726 (N_3726,N_185,N_577);
or U3727 (N_3727,N_1189,N_118);
nand U3728 (N_3728,N_1006,N_899);
nor U3729 (N_3729,N_1937,N_930);
nand U3730 (N_3730,N_671,N_1308);
and U3731 (N_3731,N_714,N_1411);
and U3732 (N_3732,N_442,N_453);
xor U3733 (N_3733,N_1267,N_1433);
nand U3734 (N_3734,N_383,N_237);
nor U3735 (N_3735,N_132,N_1341);
nor U3736 (N_3736,N_660,N_417);
nor U3737 (N_3737,N_921,N_1426);
xnor U3738 (N_3738,N_1404,N_1791);
and U3739 (N_3739,N_911,N_336);
nand U3740 (N_3740,N_1125,N_713);
nor U3741 (N_3741,N_806,N_1066);
nor U3742 (N_3742,N_1593,N_1740);
nor U3743 (N_3743,N_1205,N_1064);
and U3744 (N_3744,N_1307,N_1007);
xor U3745 (N_3745,N_182,N_1099);
or U3746 (N_3746,N_828,N_1474);
or U3747 (N_3747,N_339,N_887);
and U3748 (N_3748,N_1454,N_539);
nor U3749 (N_3749,N_679,N_907);
nor U3750 (N_3750,N_1097,N_73);
or U3751 (N_3751,N_1382,N_1442);
nand U3752 (N_3752,N_558,N_33);
nand U3753 (N_3753,N_1270,N_1230);
or U3754 (N_3754,N_847,N_1908);
nor U3755 (N_3755,N_1885,N_1781);
nand U3756 (N_3756,N_1778,N_582);
or U3757 (N_3757,N_998,N_1289);
or U3758 (N_3758,N_1903,N_1891);
nor U3759 (N_3759,N_1860,N_956);
nand U3760 (N_3760,N_632,N_809);
and U3761 (N_3761,N_1352,N_688);
nor U3762 (N_3762,N_1832,N_1273);
nor U3763 (N_3763,N_675,N_15);
xor U3764 (N_3764,N_1421,N_1832);
xnor U3765 (N_3765,N_1661,N_535);
xnor U3766 (N_3766,N_929,N_938);
or U3767 (N_3767,N_577,N_1960);
and U3768 (N_3768,N_30,N_201);
nor U3769 (N_3769,N_799,N_1715);
nand U3770 (N_3770,N_1583,N_920);
nor U3771 (N_3771,N_837,N_1933);
xor U3772 (N_3772,N_419,N_1371);
nand U3773 (N_3773,N_1618,N_50);
and U3774 (N_3774,N_745,N_540);
nor U3775 (N_3775,N_1692,N_1881);
nand U3776 (N_3776,N_42,N_498);
nand U3777 (N_3777,N_664,N_357);
nand U3778 (N_3778,N_292,N_719);
or U3779 (N_3779,N_1942,N_1180);
nand U3780 (N_3780,N_217,N_1889);
nand U3781 (N_3781,N_1823,N_1710);
and U3782 (N_3782,N_291,N_1346);
nand U3783 (N_3783,N_709,N_810);
nor U3784 (N_3784,N_1001,N_501);
xor U3785 (N_3785,N_1800,N_1473);
nor U3786 (N_3786,N_1032,N_484);
nor U3787 (N_3787,N_1490,N_706);
or U3788 (N_3788,N_1151,N_1967);
or U3789 (N_3789,N_224,N_1294);
xor U3790 (N_3790,N_1841,N_1738);
nor U3791 (N_3791,N_686,N_1444);
xor U3792 (N_3792,N_484,N_1317);
nor U3793 (N_3793,N_277,N_1995);
and U3794 (N_3794,N_236,N_849);
nand U3795 (N_3795,N_784,N_1951);
or U3796 (N_3796,N_880,N_969);
xnor U3797 (N_3797,N_1631,N_692);
and U3798 (N_3798,N_1148,N_983);
nand U3799 (N_3799,N_1686,N_646);
and U3800 (N_3800,N_347,N_842);
or U3801 (N_3801,N_952,N_559);
nor U3802 (N_3802,N_1231,N_1624);
nor U3803 (N_3803,N_402,N_187);
and U3804 (N_3804,N_699,N_506);
nor U3805 (N_3805,N_200,N_74);
nand U3806 (N_3806,N_961,N_170);
nor U3807 (N_3807,N_307,N_36);
or U3808 (N_3808,N_1004,N_1524);
nor U3809 (N_3809,N_1076,N_1260);
nor U3810 (N_3810,N_343,N_1366);
and U3811 (N_3811,N_1482,N_1243);
nand U3812 (N_3812,N_28,N_1870);
xor U3813 (N_3813,N_282,N_1918);
nor U3814 (N_3814,N_1631,N_1281);
or U3815 (N_3815,N_1204,N_988);
or U3816 (N_3816,N_1868,N_329);
and U3817 (N_3817,N_1569,N_1449);
nor U3818 (N_3818,N_1444,N_32);
xnor U3819 (N_3819,N_1883,N_905);
or U3820 (N_3820,N_1551,N_1293);
and U3821 (N_3821,N_1904,N_1061);
and U3822 (N_3822,N_931,N_1921);
nor U3823 (N_3823,N_1256,N_1831);
nand U3824 (N_3824,N_505,N_366);
nor U3825 (N_3825,N_1196,N_976);
nand U3826 (N_3826,N_1077,N_546);
nand U3827 (N_3827,N_1445,N_686);
nand U3828 (N_3828,N_1350,N_600);
nor U3829 (N_3829,N_1459,N_1956);
or U3830 (N_3830,N_1671,N_117);
nand U3831 (N_3831,N_814,N_1379);
nand U3832 (N_3832,N_482,N_1459);
or U3833 (N_3833,N_1524,N_1204);
nor U3834 (N_3834,N_1987,N_1936);
or U3835 (N_3835,N_1007,N_1510);
nor U3836 (N_3836,N_566,N_216);
and U3837 (N_3837,N_35,N_423);
nor U3838 (N_3838,N_1259,N_1007);
xor U3839 (N_3839,N_1641,N_1295);
xor U3840 (N_3840,N_1180,N_583);
or U3841 (N_3841,N_160,N_484);
and U3842 (N_3842,N_185,N_21);
nor U3843 (N_3843,N_1888,N_1969);
or U3844 (N_3844,N_1999,N_551);
nor U3845 (N_3845,N_1906,N_536);
nand U3846 (N_3846,N_1653,N_330);
nor U3847 (N_3847,N_631,N_1977);
xnor U3848 (N_3848,N_1110,N_1685);
nor U3849 (N_3849,N_1646,N_489);
nor U3850 (N_3850,N_924,N_1748);
or U3851 (N_3851,N_608,N_1437);
and U3852 (N_3852,N_544,N_578);
or U3853 (N_3853,N_25,N_1);
nand U3854 (N_3854,N_1338,N_916);
nor U3855 (N_3855,N_234,N_994);
xor U3856 (N_3856,N_1074,N_200);
nor U3857 (N_3857,N_1075,N_86);
or U3858 (N_3858,N_1779,N_357);
xor U3859 (N_3859,N_1073,N_1212);
and U3860 (N_3860,N_965,N_484);
nor U3861 (N_3861,N_588,N_1428);
xnor U3862 (N_3862,N_612,N_822);
or U3863 (N_3863,N_467,N_1178);
xor U3864 (N_3864,N_1728,N_688);
and U3865 (N_3865,N_838,N_1392);
nor U3866 (N_3866,N_269,N_724);
and U3867 (N_3867,N_726,N_1990);
xor U3868 (N_3868,N_475,N_1468);
nand U3869 (N_3869,N_916,N_331);
xnor U3870 (N_3870,N_1334,N_1620);
nor U3871 (N_3871,N_1849,N_780);
and U3872 (N_3872,N_26,N_1820);
nor U3873 (N_3873,N_1126,N_994);
nand U3874 (N_3874,N_1870,N_1575);
nor U3875 (N_3875,N_1244,N_267);
and U3876 (N_3876,N_42,N_976);
xnor U3877 (N_3877,N_974,N_824);
xor U3878 (N_3878,N_1668,N_1627);
nor U3879 (N_3879,N_124,N_1485);
xnor U3880 (N_3880,N_1922,N_395);
nand U3881 (N_3881,N_1636,N_5);
xnor U3882 (N_3882,N_687,N_1053);
and U3883 (N_3883,N_468,N_1790);
or U3884 (N_3884,N_1186,N_1655);
and U3885 (N_3885,N_1045,N_1926);
or U3886 (N_3886,N_1601,N_48);
xnor U3887 (N_3887,N_1435,N_814);
xnor U3888 (N_3888,N_618,N_1051);
xor U3889 (N_3889,N_1094,N_1569);
or U3890 (N_3890,N_1,N_1140);
or U3891 (N_3891,N_1201,N_821);
nand U3892 (N_3892,N_1863,N_703);
xnor U3893 (N_3893,N_1953,N_1811);
xor U3894 (N_3894,N_1893,N_643);
nand U3895 (N_3895,N_1541,N_520);
xnor U3896 (N_3896,N_968,N_1390);
nor U3897 (N_3897,N_1418,N_1656);
nand U3898 (N_3898,N_533,N_1130);
xnor U3899 (N_3899,N_852,N_901);
and U3900 (N_3900,N_687,N_479);
or U3901 (N_3901,N_1336,N_1984);
or U3902 (N_3902,N_1751,N_323);
or U3903 (N_3903,N_466,N_1172);
nand U3904 (N_3904,N_1670,N_1019);
and U3905 (N_3905,N_1565,N_387);
or U3906 (N_3906,N_931,N_646);
xor U3907 (N_3907,N_1634,N_1693);
nor U3908 (N_3908,N_1774,N_1303);
nand U3909 (N_3909,N_66,N_1603);
and U3910 (N_3910,N_1565,N_1846);
nor U3911 (N_3911,N_1366,N_198);
nand U3912 (N_3912,N_988,N_1977);
or U3913 (N_3913,N_321,N_1794);
xor U3914 (N_3914,N_310,N_1365);
nand U3915 (N_3915,N_1985,N_1449);
and U3916 (N_3916,N_667,N_771);
nor U3917 (N_3917,N_1269,N_1744);
xor U3918 (N_3918,N_1175,N_662);
and U3919 (N_3919,N_1812,N_1196);
xor U3920 (N_3920,N_7,N_661);
nor U3921 (N_3921,N_850,N_1039);
xnor U3922 (N_3922,N_1017,N_46);
nor U3923 (N_3923,N_1472,N_464);
and U3924 (N_3924,N_424,N_86);
xnor U3925 (N_3925,N_1902,N_1616);
or U3926 (N_3926,N_564,N_424);
nor U3927 (N_3927,N_1853,N_1815);
nand U3928 (N_3928,N_38,N_695);
nor U3929 (N_3929,N_1061,N_639);
nand U3930 (N_3930,N_1314,N_580);
xnor U3931 (N_3931,N_1672,N_1808);
or U3932 (N_3932,N_1673,N_947);
or U3933 (N_3933,N_54,N_1833);
nor U3934 (N_3934,N_982,N_1194);
nand U3935 (N_3935,N_449,N_906);
and U3936 (N_3936,N_4,N_1233);
nand U3937 (N_3937,N_248,N_553);
nand U3938 (N_3938,N_1105,N_1039);
and U3939 (N_3939,N_1167,N_247);
or U3940 (N_3940,N_816,N_1818);
nor U3941 (N_3941,N_1299,N_926);
nand U3942 (N_3942,N_1222,N_1484);
nor U3943 (N_3943,N_891,N_1139);
nand U3944 (N_3944,N_1260,N_1134);
and U3945 (N_3945,N_1015,N_1325);
nor U3946 (N_3946,N_1245,N_725);
xnor U3947 (N_3947,N_448,N_1518);
nand U3948 (N_3948,N_1009,N_1426);
xnor U3949 (N_3949,N_1785,N_767);
nand U3950 (N_3950,N_123,N_225);
or U3951 (N_3951,N_462,N_1976);
or U3952 (N_3952,N_1730,N_279);
xor U3953 (N_3953,N_1013,N_561);
and U3954 (N_3954,N_1589,N_1546);
nor U3955 (N_3955,N_356,N_1938);
and U3956 (N_3956,N_1716,N_1285);
xor U3957 (N_3957,N_1410,N_837);
xor U3958 (N_3958,N_887,N_1115);
or U3959 (N_3959,N_1478,N_1826);
and U3960 (N_3960,N_268,N_818);
nor U3961 (N_3961,N_1046,N_1393);
nand U3962 (N_3962,N_1688,N_1890);
nand U3963 (N_3963,N_1928,N_1426);
or U3964 (N_3964,N_437,N_1727);
xnor U3965 (N_3965,N_1378,N_1519);
or U3966 (N_3966,N_737,N_1);
nand U3967 (N_3967,N_1779,N_1669);
nand U3968 (N_3968,N_1066,N_786);
and U3969 (N_3969,N_280,N_1047);
xnor U3970 (N_3970,N_348,N_762);
xor U3971 (N_3971,N_192,N_882);
nor U3972 (N_3972,N_656,N_1246);
or U3973 (N_3973,N_1960,N_926);
nand U3974 (N_3974,N_1761,N_511);
nor U3975 (N_3975,N_480,N_1328);
or U3976 (N_3976,N_1083,N_1920);
xor U3977 (N_3977,N_509,N_1204);
nor U3978 (N_3978,N_503,N_32);
nand U3979 (N_3979,N_1150,N_446);
xor U3980 (N_3980,N_503,N_1279);
nor U3981 (N_3981,N_745,N_1933);
nand U3982 (N_3982,N_1357,N_1029);
nand U3983 (N_3983,N_1542,N_1877);
nand U3984 (N_3984,N_50,N_1234);
and U3985 (N_3985,N_1466,N_925);
nor U3986 (N_3986,N_992,N_879);
nand U3987 (N_3987,N_764,N_675);
nor U3988 (N_3988,N_1435,N_566);
nor U3989 (N_3989,N_535,N_645);
and U3990 (N_3990,N_740,N_774);
xnor U3991 (N_3991,N_1553,N_1230);
or U3992 (N_3992,N_1456,N_1213);
and U3993 (N_3993,N_578,N_1561);
nand U3994 (N_3994,N_1410,N_1526);
nand U3995 (N_3995,N_202,N_1537);
and U3996 (N_3996,N_502,N_204);
and U3997 (N_3997,N_1566,N_1071);
and U3998 (N_3998,N_293,N_1644);
nor U3999 (N_3999,N_454,N_580);
and U4000 (N_4000,N_2608,N_3582);
xnor U4001 (N_4001,N_3836,N_2520);
nand U4002 (N_4002,N_3954,N_3068);
nor U4003 (N_4003,N_2078,N_2507);
nand U4004 (N_4004,N_2181,N_2125);
nor U4005 (N_4005,N_2781,N_3653);
or U4006 (N_4006,N_2229,N_2142);
nand U4007 (N_4007,N_2892,N_2944);
and U4008 (N_4008,N_3554,N_2942);
and U4009 (N_4009,N_2138,N_2355);
and U4010 (N_4010,N_2332,N_3442);
xor U4011 (N_4011,N_2829,N_3595);
xor U4012 (N_4012,N_2688,N_3489);
xor U4013 (N_4013,N_3437,N_2272);
nor U4014 (N_4014,N_3285,N_3278);
nand U4015 (N_4015,N_2454,N_3759);
nand U4016 (N_4016,N_3073,N_2000);
or U4017 (N_4017,N_3923,N_2430);
or U4018 (N_4018,N_3668,N_3797);
and U4019 (N_4019,N_3784,N_2172);
and U4020 (N_4020,N_3288,N_3566);
xnor U4021 (N_4021,N_2906,N_3067);
and U4022 (N_4022,N_2686,N_3741);
or U4023 (N_4023,N_2136,N_3911);
and U4024 (N_4024,N_2976,N_2820);
xnor U4025 (N_4025,N_3903,N_3755);
and U4026 (N_4026,N_2305,N_3388);
nor U4027 (N_4027,N_3114,N_3482);
nor U4028 (N_4028,N_2995,N_2023);
xnor U4029 (N_4029,N_2870,N_3949);
and U4030 (N_4030,N_3147,N_3904);
and U4031 (N_4031,N_2844,N_2167);
xnor U4032 (N_4032,N_3453,N_2066);
and U4033 (N_4033,N_3166,N_2528);
xnor U4034 (N_4034,N_2220,N_2620);
xor U4035 (N_4035,N_2613,N_3933);
and U4036 (N_4036,N_2200,N_3985);
nand U4037 (N_4037,N_3555,N_3131);
nor U4038 (N_4038,N_3170,N_3485);
or U4039 (N_4039,N_2846,N_3331);
and U4040 (N_4040,N_3591,N_2910);
nor U4041 (N_4041,N_3488,N_3661);
xnor U4042 (N_4042,N_2329,N_3210);
and U4043 (N_4043,N_2012,N_3530);
xnor U4044 (N_4044,N_3999,N_2325);
xor U4045 (N_4045,N_2703,N_3828);
or U4046 (N_4046,N_3950,N_3586);
xor U4047 (N_4047,N_2750,N_3771);
xor U4048 (N_4048,N_2166,N_2529);
or U4049 (N_4049,N_3334,N_2415);
and U4050 (N_4050,N_3793,N_3520);
and U4051 (N_4051,N_3271,N_3409);
nor U4052 (N_4052,N_2720,N_2102);
and U4053 (N_4053,N_2130,N_3093);
xor U4054 (N_4054,N_3760,N_2572);
xnor U4055 (N_4055,N_3581,N_3357);
and U4056 (N_4056,N_3746,N_3136);
xor U4057 (N_4057,N_3924,N_2614);
nand U4058 (N_4058,N_3132,N_3328);
or U4059 (N_4059,N_2766,N_2684);
nor U4060 (N_4060,N_3543,N_2324);
xnor U4061 (N_4061,N_3994,N_2864);
and U4062 (N_4062,N_2773,N_2279);
and U4063 (N_4063,N_2231,N_3330);
nand U4064 (N_4064,N_2227,N_2994);
and U4065 (N_4065,N_3122,N_2112);
and U4066 (N_4066,N_3906,N_2095);
xor U4067 (N_4067,N_3153,N_2519);
nand U4068 (N_4068,N_3105,N_3426);
or U4069 (N_4069,N_3177,N_2506);
and U4070 (N_4070,N_3097,N_2396);
nor U4071 (N_4071,N_2353,N_3038);
nor U4072 (N_4072,N_3407,N_2173);
xnor U4073 (N_4073,N_2777,N_3648);
and U4074 (N_4074,N_3461,N_3667);
or U4075 (N_4075,N_2212,N_3229);
nand U4076 (N_4076,N_3321,N_2830);
xor U4077 (N_4077,N_2371,N_2639);
and U4078 (N_4078,N_3441,N_2103);
and U4079 (N_4079,N_2875,N_2425);
nor U4080 (N_4080,N_2246,N_2046);
and U4081 (N_4081,N_3925,N_3679);
nand U4082 (N_4082,N_3778,N_3524);
nor U4083 (N_4083,N_2216,N_2951);
nand U4084 (N_4084,N_2288,N_3724);
nor U4085 (N_4085,N_2729,N_2073);
nand U4086 (N_4086,N_2587,N_2185);
xnor U4087 (N_4087,N_3713,N_3029);
and U4088 (N_4088,N_2571,N_2453);
xnor U4089 (N_4089,N_2873,N_3474);
xnor U4090 (N_4090,N_3700,N_3337);
xnor U4091 (N_4091,N_3071,N_2561);
xor U4092 (N_4092,N_2874,N_2890);
xnor U4093 (N_4093,N_3308,N_3732);
xnor U4094 (N_4094,N_3935,N_2358);
nor U4095 (N_4095,N_3588,N_2017);
nor U4096 (N_4096,N_3421,N_3151);
and U4097 (N_4097,N_3777,N_3605);
or U4098 (N_4098,N_3881,N_3769);
nor U4099 (N_4099,N_2314,N_2597);
nand U4100 (N_4100,N_3203,N_3060);
xnor U4101 (N_4101,N_3310,N_2641);
and U4102 (N_4102,N_2949,N_2286);
nand U4103 (N_4103,N_2797,N_3876);
and U4104 (N_4104,N_2038,N_3459);
nand U4105 (N_4105,N_3841,N_2049);
or U4106 (N_4106,N_3155,N_2110);
and U4107 (N_4107,N_2492,N_2054);
and U4108 (N_4108,N_2786,N_2298);
or U4109 (N_4109,N_2232,N_2908);
nor U4110 (N_4110,N_2912,N_3557);
xnor U4111 (N_4111,N_2562,N_2438);
nor U4112 (N_4112,N_2512,N_3594);
nor U4113 (N_4113,N_3804,N_3230);
nand U4114 (N_4114,N_3291,N_2945);
nor U4115 (N_4115,N_3922,N_3625);
or U4116 (N_4116,N_3792,N_2582);
xnor U4117 (N_4117,N_3043,N_3216);
nor U4118 (N_4118,N_2192,N_3103);
nand U4119 (N_4119,N_2410,N_2297);
nor U4120 (N_4120,N_2113,N_3432);
nor U4121 (N_4121,N_3259,N_2764);
nor U4122 (N_4122,N_3338,N_2386);
nand U4123 (N_4123,N_3176,N_2093);
or U4124 (N_4124,N_2565,N_3194);
or U4125 (N_4125,N_2065,N_3044);
xnor U4126 (N_4126,N_3495,N_2165);
or U4127 (N_4127,N_3830,N_2815);
nor U4128 (N_4128,N_2315,N_2550);
and U4129 (N_4129,N_3164,N_2121);
nor U4130 (N_4130,N_3575,N_2645);
nand U4131 (N_4131,N_2886,N_2075);
and U4132 (N_4132,N_2857,N_2170);
and U4133 (N_4133,N_3048,N_3061);
and U4134 (N_4134,N_3745,N_2098);
nor U4135 (N_4135,N_2547,N_3878);
xnor U4136 (N_4136,N_2318,N_3753);
or U4137 (N_4137,N_3635,N_2847);
nand U4138 (N_4138,N_3801,N_3738);
nor U4139 (N_4139,N_2319,N_3847);
nand U4140 (N_4140,N_3691,N_3026);
nor U4141 (N_4141,N_2558,N_2256);
and U4142 (N_4142,N_2001,N_2347);
xnor U4143 (N_4143,N_3579,N_3231);
nor U4144 (N_4144,N_3909,N_2651);
nor U4145 (N_4145,N_3009,N_3714);
and U4146 (N_4146,N_3694,N_3383);
nand U4147 (N_4147,N_2317,N_2311);
nand U4148 (N_4148,N_3240,N_2665);
nor U4149 (N_4149,N_3242,N_3987);
nand U4150 (N_4150,N_3765,N_2367);
nand U4151 (N_4151,N_3892,N_3580);
and U4152 (N_4152,N_2484,N_2264);
xnor U4153 (N_4153,N_2242,N_3425);
and U4154 (N_4154,N_3056,N_2235);
nand U4155 (N_4155,N_2622,N_3182);
or U4156 (N_4156,N_3380,N_3440);
xor U4157 (N_4157,N_2822,N_3199);
or U4158 (N_4158,N_3631,N_2294);
and U4159 (N_4159,N_3392,N_2037);
nor U4160 (N_4160,N_2022,N_3945);
or U4161 (N_4161,N_3113,N_2029);
xnor U4162 (N_4162,N_2801,N_2150);
nand U4163 (N_4163,N_2159,N_2151);
nor U4164 (N_4164,N_2683,N_2255);
nand U4165 (N_4165,N_2322,N_2211);
and U4166 (N_4166,N_2302,N_2798);
xnor U4167 (N_4167,N_2653,N_2304);
nand U4168 (N_4168,N_3196,N_2655);
xor U4169 (N_4169,N_2041,N_2602);
and U4170 (N_4170,N_2031,N_3018);
xor U4171 (N_4171,N_3200,N_2591);
and U4172 (N_4172,N_3799,N_3013);
and U4173 (N_4173,N_2033,N_3864);
nor U4174 (N_4174,N_3818,N_3254);
nand U4175 (N_4175,N_3090,N_2494);
or U4176 (N_4176,N_3632,N_3251);
or U4177 (N_4177,N_3592,N_3703);
nand U4178 (N_4178,N_3910,N_2897);
xnor U4179 (N_4179,N_3419,N_2427);
nand U4180 (N_4180,N_3598,N_2491);
or U4181 (N_4181,N_2850,N_3567);
nand U4182 (N_4182,N_3206,N_2486);
or U4183 (N_4183,N_3036,N_2475);
nor U4184 (N_4184,N_3726,N_3888);
xnor U4185 (N_4185,N_3333,N_3469);
and U4186 (N_4186,N_3900,N_2698);
or U4187 (N_4187,N_2364,N_2989);
and U4188 (N_4188,N_3133,N_2123);
and U4189 (N_4189,N_2955,N_2939);
nand U4190 (N_4190,N_3144,N_3261);
nand U4191 (N_4191,N_3596,N_2556);
xor U4192 (N_4192,N_3709,N_2444);
or U4193 (N_4193,N_2749,N_2933);
nor U4194 (N_4194,N_3188,N_2851);
nor U4195 (N_4195,N_3977,N_2435);
and U4196 (N_4196,N_3907,N_2674);
or U4197 (N_4197,N_3313,N_3503);
nand U4198 (N_4198,N_3610,N_2008);
nor U4199 (N_4199,N_2226,N_2838);
xor U4200 (N_4200,N_3207,N_3919);
and U4201 (N_4201,N_3644,N_3831);
nor U4202 (N_4202,N_2096,N_2928);
and U4203 (N_4203,N_2133,N_3360);
and U4204 (N_4204,N_3494,N_3341);
and U4205 (N_4205,N_3339,N_2398);
or U4206 (N_4206,N_3602,N_3052);
or U4207 (N_4207,N_3542,N_3189);
nor U4208 (N_4208,N_2336,N_2199);
and U4209 (N_4209,N_3344,N_2950);
nand U4210 (N_4210,N_2187,N_2296);
and U4211 (N_4211,N_2868,N_3902);
nor U4212 (N_4212,N_3435,N_2960);
or U4213 (N_4213,N_3011,N_2044);
nor U4214 (N_4214,N_2553,N_3154);
or U4215 (N_4215,N_3371,N_3627);
nor U4216 (N_4216,N_3209,N_3974);
nand U4217 (N_4217,N_3318,N_2848);
nor U4218 (N_4218,N_2377,N_3617);
xor U4219 (N_4219,N_2712,N_3604);
xnor U4220 (N_4220,N_2349,N_3965);
or U4221 (N_4221,N_2035,N_2356);
nor U4222 (N_4222,N_3448,N_2117);
nor U4223 (N_4223,N_2947,N_3787);
and U4224 (N_4224,N_2807,N_2052);
and U4225 (N_4225,N_3306,N_3014);
and U4226 (N_4226,N_2738,N_2202);
and U4227 (N_4227,N_2708,N_3549);
and U4228 (N_4228,N_3424,N_2281);
and U4229 (N_4229,N_3171,N_2659);
xnor U4230 (N_4230,N_2896,N_2275);
nor U4231 (N_4231,N_3405,N_2411);
nand U4232 (N_4232,N_3368,N_2616);
or U4233 (N_4233,N_3953,N_3316);
xor U4234 (N_4234,N_3577,N_2292);
or U4235 (N_4235,N_2293,N_3168);
nor U4236 (N_4236,N_2009,N_3031);
nand U4237 (N_4237,N_3289,N_3678);
nand U4238 (N_4238,N_2740,N_3761);
or U4239 (N_4239,N_2026,N_2510);
and U4240 (N_4240,N_2824,N_3372);
nand U4241 (N_4241,N_3250,N_2603);
xor U4242 (N_4242,N_2340,N_2652);
or U4243 (N_4243,N_2880,N_2495);
and U4244 (N_4244,N_3266,N_3352);
nor U4245 (N_4245,N_2577,N_3197);
xnor U4246 (N_4246,N_2618,N_2463);
nor U4247 (N_4247,N_3719,N_3397);
xnor U4248 (N_4248,N_2039,N_3563);
and U4249 (N_4249,N_3384,N_2178);
nand U4250 (N_4250,N_2077,N_2145);
or U4251 (N_4251,N_3650,N_2114);
nand U4252 (N_4252,N_2105,N_3423);
or U4253 (N_4253,N_3119,N_3106);
or U4254 (N_4254,N_3253,N_3673);
or U4255 (N_4255,N_3589,N_3740);
and U4256 (N_4256,N_3649,N_2504);
nand U4257 (N_4257,N_2051,N_2437);
or U4258 (N_4258,N_2466,N_2775);
nor U4259 (N_4259,N_3433,N_3032);
nand U4260 (N_4260,N_3645,N_2776);
nor U4261 (N_4261,N_2631,N_3326);
and U4262 (N_4262,N_3205,N_2748);
xnor U4263 (N_4263,N_3693,N_3715);
nand U4264 (N_4264,N_2316,N_2985);
or U4265 (N_4265,N_2918,N_2879);
or U4266 (N_4266,N_2094,N_3415);
nand U4267 (N_4267,N_3305,N_2455);
nand U4268 (N_4268,N_2551,N_3226);
or U4269 (N_4269,N_3078,N_3129);
nor U4270 (N_4270,N_3082,N_2018);
nand U4271 (N_4271,N_2308,N_2835);
xor U4272 (N_4272,N_3237,N_3996);
and U4273 (N_4273,N_2662,N_2793);
nand U4274 (N_4274,N_2433,N_2280);
or U4275 (N_4275,N_3790,N_2993);
or U4276 (N_4276,N_3717,N_2759);
nand U4277 (N_4277,N_2607,N_3270);
or U4278 (N_4278,N_3476,N_3852);
or U4279 (N_4279,N_3224,N_2849);
or U4280 (N_4280,N_3844,N_3651);
or U4281 (N_4281,N_3794,N_3532);
xnor U4282 (N_4282,N_2059,N_2991);
nand U4283 (N_4283,N_2532,N_2456);
nand U4284 (N_4284,N_2929,N_3896);
nand U4285 (N_4285,N_3674,N_3152);
nand U4286 (N_4286,N_2111,N_3249);
or U4287 (N_4287,N_2865,N_2770);
or U4288 (N_4288,N_2030,N_2186);
xor U4289 (N_4289,N_3614,N_2704);
xor U4290 (N_4290,N_3590,N_3699);
and U4291 (N_4291,N_3932,N_3742);
and U4292 (N_4292,N_3553,N_3355);
or U4293 (N_4293,N_2025,N_2774);
and U4294 (N_4294,N_2040,N_2753);
nand U4295 (N_4295,N_3361,N_2716);
nor U4296 (N_4296,N_3764,N_3087);
nand U4297 (N_4297,N_2149,N_3963);
and U4298 (N_4298,N_3376,N_2464);
nand U4299 (N_4299,N_3471,N_2062);
nor U4300 (N_4300,N_2952,N_3214);
and U4301 (N_4301,N_3180,N_2705);
xor U4302 (N_4302,N_3422,N_3460);
or U4303 (N_4303,N_2160,N_2417);
nor U4304 (N_4304,N_3335,N_2672);
xnor U4305 (N_4305,N_3130,N_2236);
nand U4306 (N_4306,N_3211,N_2580);
nand U4307 (N_4307,N_2441,N_2782);
nand U4308 (N_4308,N_3885,N_2042);
and U4309 (N_4309,N_2327,N_3697);
nand U4310 (N_4310,N_3603,N_2083);
or U4311 (N_4311,N_2348,N_3121);
xnor U4312 (N_4312,N_2005,N_2461);
and U4313 (N_4313,N_2462,N_2099);
xnor U4314 (N_4314,N_3192,N_2966);
and U4315 (N_4315,N_3116,N_3547);
nand U4316 (N_4316,N_2642,N_3099);
nand U4317 (N_4317,N_3293,N_3245);
nor U4318 (N_4318,N_3796,N_2654);
xnor U4319 (N_4319,N_2617,N_3565);
nand U4320 (N_4320,N_3367,N_3159);
and U4321 (N_4321,N_2266,N_2833);
nor U4322 (N_4322,N_2223,N_2143);
and U4323 (N_4323,N_2596,N_2489);
xnor U4324 (N_4324,N_3141,N_3817);
or U4325 (N_4325,N_2731,N_2036);
and U4326 (N_4326,N_2791,N_3315);
nor U4327 (N_4327,N_2180,N_2924);
or U4328 (N_4328,N_2526,N_3268);
and U4329 (N_4329,N_3109,N_2592);
nand U4330 (N_4330,N_2426,N_3638);
or U4331 (N_4331,N_3486,N_3533);
xnor U4332 (N_4332,N_3859,N_3185);
nor U4333 (N_4333,N_2208,N_3190);
and U4334 (N_4334,N_2423,N_2442);
and U4335 (N_4335,N_2154,N_3721);
and U4336 (N_4336,N_2522,N_2428);
or U4337 (N_4337,N_2195,N_2863);
nand U4338 (N_4338,N_2541,N_3964);
or U4339 (N_4339,N_2309,N_2174);
or U4340 (N_4340,N_3633,N_2946);
and U4341 (N_4341,N_3641,N_2930);
and U4342 (N_4342,N_3791,N_2106);
nor U4343 (N_4343,N_2816,N_3898);
and U4344 (N_4344,N_3126,N_2626);
xor U4345 (N_4345,N_2080,N_3160);
nand U4346 (N_4346,N_3946,N_2888);
nand U4347 (N_4347,N_3498,N_2789);
and U4348 (N_4348,N_2934,N_2300);
or U4349 (N_4349,N_2373,N_3665);
nor U4350 (N_4350,N_3404,N_3004);
or U4351 (N_4351,N_3774,N_3897);
and U4352 (N_4352,N_3223,N_3019);
or U4353 (N_4353,N_2067,N_2011);
xnor U4354 (N_4354,N_3300,N_2074);
and U4355 (N_4355,N_2534,N_2284);
or U4356 (N_4356,N_2061,N_2633);
nor U4357 (N_4357,N_3527,N_2443);
nand U4358 (N_4358,N_3642,N_3978);
or U4359 (N_4359,N_2389,N_3157);
nand U4360 (N_4360,N_2124,N_3822);
xnor U4361 (N_4361,N_3639,N_3669);
nand U4362 (N_4362,N_3507,N_2867);
and U4363 (N_4363,N_3710,N_3795);
and U4364 (N_4364,N_3267,N_3387);
or U4365 (N_4365,N_3983,N_3395);
xor U4366 (N_4366,N_2129,N_2871);
nand U4367 (N_4367,N_3840,N_2097);
nand U4368 (N_4368,N_3329,N_2467);
nor U4369 (N_4369,N_2761,N_3772);
xor U4370 (N_4370,N_2413,N_3287);
xor U4371 (N_4371,N_2076,N_2086);
xnor U4372 (N_4372,N_2746,N_3024);
and U4373 (N_4373,N_3802,N_2525);
or U4374 (N_4374,N_2784,N_3599);
nand U4375 (N_4375,N_2927,N_2161);
nand U4376 (N_4376,N_2954,N_3875);
nor U4377 (N_4377,N_2261,N_2267);
xor U4378 (N_4378,N_3652,N_2222);
nor U4379 (N_4379,N_2120,N_2902);
xor U4380 (N_4380,N_2574,N_2663);
and U4381 (N_4381,N_3447,N_3863);
and U4382 (N_4382,N_3905,N_2917);
or U4383 (N_4383,N_3213,N_2056);
and U4384 (N_4384,N_3518,N_3000);
xor U4385 (N_4385,N_3283,N_2730);
nor U4386 (N_4386,N_3396,N_3028);
xor U4387 (N_4387,N_2689,N_2505);
and U4388 (N_4388,N_3508,N_3952);
nand U4389 (N_4389,N_3280,N_2383);
or U4390 (N_4390,N_3272,N_2515);
and U4391 (N_4391,N_2109,N_2583);
xor U4392 (N_4392,N_3809,N_3008);
and U4393 (N_4393,N_3186,N_3069);
nor U4394 (N_4394,N_3275,N_2420);
nor U4395 (N_4395,N_2248,N_2218);
and U4396 (N_4396,N_2713,N_2387);
nand U4397 (N_4397,N_2352,N_3583);
nor U4398 (N_4398,N_2938,N_2168);
and U4399 (N_4399,N_3893,N_3218);
and U4400 (N_4400,N_2840,N_3944);
nand U4401 (N_4401,N_3016,N_2412);
or U4402 (N_4402,N_3427,N_2263);
xor U4403 (N_4403,N_2682,N_3049);
xnor U4404 (N_4404,N_2201,N_2384);
or U4405 (N_4405,N_2401,N_2245);
nor U4406 (N_4406,N_3228,N_3247);
and U4407 (N_4407,N_3656,N_2543);
xor U4408 (N_4408,N_3672,N_3869);
and U4409 (N_4409,N_3456,N_2247);
xnor U4410 (N_4410,N_3538,N_3463);
and U4411 (N_4411,N_2418,N_3502);
nor U4412 (N_4412,N_3125,N_2003);
nor U4413 (N_4413,N_2872,N_3748);
and U4414 (N_4414,N_3111,N_3991);
nor U4415 (N_4415,N_2756,N_3992);
nand U4416 (N_4416,N_2539,N_2959);
xnor U4417 (N_4417,N_2502,N_2233);
xnor U4418 (N_4418,N_3483,N_2100);
nand U4419 (N_4419,N_3947,N_2996);
nand U4420 (N_4420,N_3516,N_3773);
nand U4421 (N_4421,N_2002,N_2589);
and U4422 (N_4422,N_3350,N_2937);
nand U4423 (N_4423,N_2811,N_2068);
and U4424 (N_4424,N_3092,N_3750);
or U4425 (N_4425,N_2862,N_2881);
nand U4426 (N_4426,N_3920,N_3883);
or U4427 (N_4427,N_2345,N_2610);
nor U4428 (N_4428,N_3478,N_3937);
xor U4429 (N_4429,N_2434,N_2481);
and U4430 (N_4430,N_2940,N_2431);
or U4431 (N_4431,N_2147,N_2176);
or U4432 (N_4432,N_2762,N_3263);
or U4433 (N_4433,N_2588,N_2694);
xnor U4434 (N_4434,N_2079,N_3889);
nand U4435 (N_4435,N_3001,N_3846);
or U4436 (N_4436,N_3870,N_2702);
or U4437 (N_4437,N_2472,N_3936);
nor U4438 (N_4438,N_3551,N_3541);
nor U4439 (N_4439,N_3539,N_2183);
and U4440 (N_4440,N_2122,N_3412);
nor U4441 (N_4441,N_3233,N_3047);
and U4442 (N_4442,N_2611,N_3833);
or U4443 (N_4443,N_3640,N_3767);
nand U4444 (N_4444,N_3346,N_2845);
xnor U4445 (N_4445,N_3766,N_2483);
xor U4446 (N_4446,N_2278,N_3597);
nor U4447 (N_4447,N_3684,N_2800);
xnor U4448 (N_4448,N_2213,N_3094);
xor U4449 (N_4449,N_2823,N_2509);
nand U4450 (N_4450,N_3400,N_2754);
and U4451 (N_4451,N_3501,N_3187);
xor U4452 (N_4452,N_2792,N_3630);
nor U4453 (N_4453,N_3534,N_2070);
or U4454 (N_4454,N_2104,N_3022);
and U4455 (N_4455,N_2189,N_3349);
xnor U4456 (N_4456,N_2678,N_3730);
or U4457 (N_4457,N_2818,N_3509);
xor U4458 (N_4458,N_3628,N_2696);
or U4459 (N_4459,N_2931,N_2891);
nor U4460 (N_4460,N_2637,N_2313);
xor U4461 (N_4461,N_2338,N_2307);
xnor U4462 (N_4462,N_3913,N_3756);
and U4463 (N_4463,N_2019,N_3354);
nand U4464 (N_4464,N_2381,N_3688);
nand U4465 (N_4465,N_2666,N_3813);
xor U4466 (N_4466,N_3059,N_2915);
xnor U4467 (N_4467,N_2579,N_2177);
nand U4468 (N_4468,N_3212,N_2973);
and U4469 (N_4469,N_2141,N_3243);
nand U4470 (N_4470,N_3576,N_2893);
xor U4471 (N_4471,N_3845,N_2414);
or U4472 (N_4472,N_2175,N_3587);
or U4473 (N_4473,N_2204,N_3839);
nand U4474 (N_4474,N_2287,N_3364);
and U4475 (N_4475,N_3975,N_2734);
xnor U4476 (N_4476,N_3124,N_3430);
xnor U4477 (N_4477,N_3015,N_2372);
and U4478 (N_4478,N_3681,N_3148);
xor U4479 (N_4479,N_2511,N_2119);
and U4480 (N_4480,N_2171,N_3276);
nor U4481 (N_4481,N_2291,N_3776);
xor U4482 (N_4482,N_2805,N_2252);
nand U4483 (N_4483,N_3757,N_2469);
and U4484 (N_4484,N_3234,N_2508);
nand U4485 (N_4485,N_3239,N_3374);
nor U4486 (N_4486,N_3788,N_2595);
and U4487 (N_4487,N_3506,N_2540);
nor U4488 (N_4488,N_3411,N_2735);
and U4489 (N_4489,N_3654,N_2354);
or U4490 (N_4490,N_3063,N_3927);
nand U4491 (N_4491,N_2953,N_3948);
xor U4492 (N_4492,N_3406,N_3882);
or U4493 (N_4493,N_2091,N_3320);
nor U4494 (N_4494,N_2992,N_2788);
or U4495 (N_4495,N_2295,N_3439);
nor U4496 (N_4496,N_2214,N_2517);
or U4497 (N_4497,N_2028,N_3564);
nand U4498 (N_4498,N_3225,N_2695);
xor U4499 (N_4499,N_3785,N_2697);
nor U4500 (N_4500,N_2779,N_3464);
and U4501 (N_4501,N_2346,N_3812);
and U4502 (N_4502,N_2399,N_3856);
nand U4503 (N_4503,N_3708,N_3626);
and U4504 (N_4504,N_3561,N_3161);
nor U4505 (N_4505,N_3517,N_3264);
nand U4506 (N_4506,N_3929,N_2623);
xor U4507 (N_4507,N_2209,N_2194);
xor U4508 (N_4508,N_2922,N_3299);
nand U4509 (N_4509,N_3500,N_3449);
and U4510 (N_4510,N_3528,N_3615);
or U4511 (N_4511,N_3066,N_3735);
nand U4512 (N_4512,N_3312,N_2476);
and U4513 (N_4513,N_3664,N_2739);
xor U4514 (N_4514,N_2673,N_3980);
nand U4515 (N_4515,N_2555,N_2419);
nand U4516 (N_4516,N_3807,N_3191);
nand U4517 (N_4517,N_2468,N_3085);
nor U4518 (N_4518,N_2619,N_3173);
and U4519 (N_4519,N_3786,N_3296);
nand U4520 (N_4520,N_2439,N_2344);
xor U4521 (N_4521,N_2394,N_3174);
nand U4522 (N_4522,N_3158,N_3260);
xor U4523 (N_4523,N_2667,N_2135);
nand U4524 (N_4524,N_3737,N_2737);
and U4525 (N_4525,N_2964,N_2380);
and U4526 (N_4526,N_2866,N_3410);
nand U4527 (N_4527,N_3053,N_3611);
nor U4528 (N_4528,N_2911,N_3523);
nand U4529 (N_4529,N_2341,N_3914);
or U4530 (N_4530,N_2956,N_3244);
nor U4531 (N_4531,N_3403,N_2493);
nand U4532 (N_4532,N_2987,N_2385);
nor U4533 (N_4533,N_2570,N_3522);
or U4534 (N_4534,N_2743,N_2262);
or U4535 (N_4535,N_3727,N_3262);
or U4536 (N_4536,N_3918,N_3990);
or U4537 (N_4537,N_3294,N_3749);
nand U4538 (N_4538,N_3662,N_3466);
and U4539 (N_4539,N_2861,N_3378);
nand U4540 (N_4540,N_3866,N_3179);
nand U4541 (N_4541,N_2899,N_2471);
nand U4542 (N_4542,N_2225,N_2599);
and U4543 (N_4543,N_3479,N_2676);
xor U4544 (N_4544,N_3193,N_3823);
xnor U4545 (N_4545,N_3477,N_2478);
or U4546 (N_4546,N_3219,N_3054);
or U4547 (N_4547,N_3930,N_2258);
nand U4548 (N_4548,N_3353,N_3358);
nand U4549 (N_4549,N_3201,N_3408);
and U4550 (N_4550,N_3208,N_2043);
xor U4551 (N_4551,N_2794,N_3770);
and U4552 (N_4552,N_2326,N_3803);
and U4553 (N_4553,N_2339,N_3434);
and U4554 (N_4554,N_3702,N_2943);
xnor U4555 (N_4555,N_3327,N_3972);
or U4556 (N_4556,N_3926,N_2271);
xor U4557 (N_4557,N_2482,N_3544);
nor U4558 (N_4558,N_3690,N_2919);
or U4559 (N_4559,N_3843,N_2628);
xnor U4560 (N_4560,N_3938,N_2717);
xnor U4561 (N_4561,N_3705,N_3997);
nor U4562 (N_4562,N_2545,N_3452);
or U4563 (N_4563,N_2516,N_3002);
xor U4564 (N_4564,N_2169,N_2312);
nand U4565 (N_4565,N_3865,N_3042);
xnor U4566 (N_4566,N_3468,N_3086);
nand U4567 (N_4567,N_2709,N_3304);
or U4568 (N_4568,N_2290,N_2269);
and U4569 (N_4569,N_2131,N_2690);
and U4570 (N_4570,N_3696,N_3083);
or U4571 (N_4571,N_2630,N_3752);
and U4572 (N_4572,N_3815,N_3908);
or U4573 (N_4573,N_2128,N_2563);
nor U4574 (N_4574,N_3971,N_2397);
nor U4575 (N_4575,N_2921,N_2207);
and U4576 (N_4576,N_2392,N_3572);
or U4577 (N_4577,N_3045,N_2436);
xor U4578 (N_4578,N_3838,N_3115);
or U4579 (N_4579,N_3961,N_2368);
xnor U4580 (N_4580,N_2923,N_3499);
xnor U4581 (N_4581,N_3871,N_3685);
nor U4582 (N_4582,N_2627,N_2907);
or U4583 (N_4583,N_2162,N_3711);
or U4584 (N_4584,N_2640,N_2337);
and U4585 (N_4585,N_2283,N_2538);
xnor U4586 (N_4586,N_3958,N_3098);
and U4587 (N_4587,N_3515,N_2721);
nand U4588 (N_4588,N_2671,N_2914);
nor U4589 (N_4589,N_2860,N_3701);
nand U4590 (N_4590,N_3676,N_3235);
nand U4591 (N_4591,N_2615,N_2542);
or U4592 (N_4592,N_2268,N_2365);
or U4593 (N_4593,N_2578,N_2884);
or U4594 (N_4594,N_2328,N_3167);
and U4595 (N_4595,N_2821,N_3282);
xnor U4596 (N_4596,N_3359,N_3600);
nor U4597 (N_4597,N_2968,N_2714);
or U4598 (N_4598,N_2900,N_2806);
nand U4599 (N_4599,N_2841,N_2048);
and U4600 (N_4600,N_2404,N_3149);
nand U4601 (N_4601,N_3618,N_2988);
xnor U4602 (N_4602,N_3379,N_2771);
or U4603 (N_4603,N_3988,N_3917);
and U4604 (N_4604,N_3825,N_2767);
nor U4605 (N_4605,N_3277,N_2537);
nand U4606 (N_4606,N_2826,N_3005);
nor U4607 (N_4607,N_2982,N_2490);
nor U4608 (N_4608,N_3363,N_3916);
xnor U4609 (N_4609,N_2566,N_3431);
or U4610 (N_4610,N_2027,N_2330);
xnor U4611 (N_4611,N_3571,N_2559);
nor U4612 (N_4612,N_2546,N_3556);
or U4613 (N_4613,N_3181,N_2407);
or U4614 (N_4614,N_2710,N_3065);
nand U4615 (N_4615,N_3616,N_2527);
nand U4616 (N_4616,N_3137,N_3894);
xor U4617 (N_4617,N_2306,N_3962);
and U4618 (N_4618,N_2063,N_2751);
nand U4619 (N_4619,N_2084,N_2675);
or U4620 (N_4620,N_3683,N_2701);
nor U4621 (N_4621,N_3145,N_2140);
or U4622 (N_4622,N_3569,N_3490);
or U4623 (N_4623,N_3418,N_3178);
xor U4624 (N_4624,N_2733,N_2681);
or U4625 (N_4625,N_3169,N_2020);
and U4626 (N_4626,N_2163,N_2240);
and U4627 (N_4627,N_3890,N_3873);
nand U4628 (N_4628,N_3529,N_3608);
or U4629 (N_4629,N_2742,N_3511);
xnor U4630 (N_4630,N_2503,N_2474);
nand U4631 (N_4631,N_2488,N_2920);
or U4632 (N_4632,N_2343,N_2625);
nand U4633 (N_4633,N_2408,N_2660);
nand U4634 (N_4634,N_3118,N_3058);
or U4635 (N_4635,N_2685,N_3417);
and U4636 (N_4636,N_3834,N_3887);
nor U4637 (N_4637,N_2182,N_2722);
nand U4638 (N_4638,N_2790,N_2984);
nor U4639 (N_4639,N_2948,N_2379);
nor U4640 (N_4640,N_3728,N_3548);
nor U4641 (N_4641,N_2898,N_2707);
nor U4642 (N_4642,N_3519,N_2817);
and U4643 (N_4643,N_3659,N_2157);
or U4644 (N_4644,N_2299,N_3573);
and U4645 (N_4645,N_3007,N_3744);
and U4646 (N_4646,N_3723,N_3322);
nand U4647 (N_4647,N_2069,N_3646);
and U4648 (N_4648,N_2193,N_2699);
or U4649 (N_4649,N_2834,N_2549);
or U4650 (N_4650,N_3780,N_3110);
and U4651 (N_4651,N_2644,N_2600);
or U4652 (N_4652,N_2768,N_2916);
nand U4653 (N_4653,N_2963,N_2970);
nand U4654 (N_4654,N_3074,N_3401);
or U4655 (N_4655,N_3976,N_2593);
or U4656 (N_4656,N_2554,N_3826);
and U4657 (N_4657,N_2015,N_2055);
nand U4658 (N_4658,N_2718,N_2926);
nand U4659 (N_4659,N_3080,N_3540);
nand U4660 (N_4660,N_3560,N_2972);
xnor U4661 (N_4661,N_3222,N_3369);
nand U4662 (N_4662,N_2137,N_2650);
and U4663 (N_4663,N_2635,N_3775);
xnor U4664 (N_4664,N_3734,N_3020);
xnor U4665 (N_4665,N_3398,N_3718);
xor U4666 (N_4666,N_2197,N_3107);
and U4667 (N_4667,N_2523,N_3956);
nand U4668 (N_4668,N_3342,N_3623);
nor U4669 (N_4669,N_2859,N_2422);
or U4670 (N_4670,N_2719,N_3057);
xor U4671 (N_4671,N_2518,N_3829);
or U4672 (N_4672,N_2760,N_3504);
nor U4673 (N_4673,N_3040,N_2885);
nand U4674 (N_4674,N_3143,N_3810);
xor U4675 (N_4675,N_2852,N_3302);
or U4676 (N_4676,N_3055,N_2590);
or U4677 (N_4677,N_3862,N_3492);
nor U4678 (N_4678,N_3680,N_2536);
or U4679 (N_4679,N_2060,N_2496);
xor U4680 (N_4680,N_2901,N_3290);
nor U4681 (N_4681,N_2249,N_2082);
or U4682 (N_4682,N_3414,N_3402);
nor U4683 (N_4683,N_2839,N_3156);
or U4684 (N_4684,N_3660,N_3970);
xor U4685 (N_4685,N_3150,N_3356);
or U4686 (N_4686,N_2139,N_3345);
or U4687 (N_4687,N_2819,N_3943);
and U4688 (N_4688,N_2711,N_2757);
and U4689 (N_4689,N_3968,N_3695);
or U4690 (N_4690,N_3850,N_2445);
nor U4691 (N_4691,N_3246,N_2032);
nor U4692 (N_4692,N_2006,N_3003);
or U4693 (N_4693,N_3550,N_2303);
nand U4694 (N_4694,N_2842,N_2796);
or U4695 (N_4695,N_2090,N_2331);
nand U4696 (N_4696,N_3428,N_3657);
xor U4697 (N_4697,N_2606,N_2155);
nand U4698 (N_4698,N_2072,N_2827);
and U4699 (N_4699,N_3851,N_3458);
nand U4700 (N_4700,N_2531,N_3781);
xnor U4701 (N_4701,N_3782,N_2250);
nand U4702 (N_4702,N_3798,N_2513);
xnor U4703 (N_4703,N_3891,N_3429);
or U4704 (N_4704,N_3979,N_2146);
xnor U4705 (N_4705,N_2498,N_3487);
xnor U4706 (N_4706,N_3915,N_3899);
nor U4707 (N_4707,N_3381,N_3981);
xor U4708 (N_4708,N_2535,N_3446);
or U4709 (N_4709,N_3619,N_2152);
and U4710 (N_4710,N_2239,N_3806);
xnor U4711 (N_4711,N_3309,N_2126);
nand U4712 (N_4712,N_3140,N_2814);
and U4713 (N_4713,N_2586,N_2575);
xnor U4714 (N_4714,N_3973,N_2470);
nor U4715 (N_4715,N_2323,N_2421);
xor U4716 (N_4716,N_2228,N_2127);
nand U4717 (N_4717,N_3104,N_2230);
and U4718 (N_4718,N_2480,N_2715);
xor U4719 (N_4719,N_2664,N_3819);
xor U4720 (N_4720,N_3072,N_3484);
and U4721 (N_4721,N_2783,N_2726);
nor U4722 (N_4722,N_3279,N_2357);
nor U4723 (N_4723,N_2458,N_2024);
xor U4724 (N_4724,N_3146,N_2856);
and U4725 (N_4725,N_2670,N_2497);
and U4726 (N_4726,N_2894,N_3454);
or U4727 (N_4727,N_2828,N_2895);
nand U4728 (N_4728,N_3443,N_3860);
or U4729 (N_4729,N_2643,N_3088);
xor U4730 (N_4730,N_2986,N_3568);
nand U4731 (N_4731,N_3389,N_2285);
xnor U4732 (N_4732,N_3236,N_3217);
nor U4733 (N_4733,N_2758,N_2878);
xor U4734 (N_4734,N_3624,N_3934);
and U4735 (N_4735,N_3536,N_3347);
nor U4736 (N_4736,N_2962,N_2196);
nor U4737 (N_4737,N_2785,N_2088);
or U4738 (N_4738,N_2215,N_3079);
nor U4739 (N_4739,N_2581,N_3986);
and U4740 (N_4740,N_2567,N_2679);
nor U4741 (N_4741,N_3512,N_3731);
or U4742 (N_4742,N_2983,N_3842);
and U4743 (N_4743,N_3227,N_2803);
and U4744 (N_4744,N_3382,N_2752);
nand U4745 (N_4745,N_3062,N_3297);
nor U4746 (N_4746,N_2144,N_3420);
nand U4747 (N_4747,N_3634,N_2460);
xnor U4748 (N_4748,N_2382,N_2727);
xor U4749 (N_4749,N_2552,N_3027);
nor U4750 (N_4750,N_3827,N_2629);
nor U4751 (N_4751,N_3336,N_2241);
xnor U4752 (N_4752,N_3675,N_2277);
nand U4753 (N_4753,N_2691,N_2706);
or U4754 (N_4754,N_3811,N_2687);
and U4755 (N_4755,N_2447,N_3365);
nand U4756 (N_4756,N_3585,N_2961);
nand U4757 (N_4757,N_2723,N_2621);
nor U4758 (N_4758,N_3901,N_2925);
nor U4759 (N_4759,N_2747,N_3413);
nor U4760 (N_4760,N_3989,N_3096);
nand U4761 (N_4761,N_3091,N_3162);
xor U4762 (N_4762,N_3689,N_3720);
nor U4763 (N_4763,N_2741,N_2276);
nand U4764 (N_4764,N_2501,N_3257);
xor U4765 (N_4765,N_3295,N_3248);
nand U4766 (N_4766,N_3637,N_3800);
nand U4767 (N_4767,N_3636,N_3325);
and U4768 (N_4768,N_3163,N_2778);
nor U4769 (N_4769,N_3758,N_3525);
nand U4770 (N_4770,N_3221,N_3252);
nor U4771 (N_4771,N_2548,N_3629);
or U4772 (N_4772,N_2334,N_3872);
xor U4773 (N_4773,N_2485,N_3643);
or U4774 (N_4774,N_2134,N_2843);
and U4775 (N_4775,N_2813,N_2010);
and U4776 (N_4776,N_3095,N_2661);
and U4777 (N_4777,N_3612,N_2882);
and U4778 (N_4778,N_2057,N_3647);
or U4779 (N_4779,N_2473,N_2990);
xor U4780 (N_4780,N_3814,N_3348);
nand U4781 (N_4781,N_3816,N_2350);
and U4782 (N_4782,N_3102,N_3886);
xor U4783 (N_4783,N_2432,N_2812);
nor U4784 (N_4784,N_2799,N_3729);
nand U4785 (N_4785,N_3747,N_2763);
nand U4786 (N_4786,N_3677,N_2649);
and U4787 (N_4787,N_3394,N_3768);
nand U4788 (N_4788,N_2362,N_2700);
and U4789 (N_4789,N_3172,N_2335);
or U4790 (N_4790,N_3450,N_3609);
nand U4791 (N_4791,N_3220,N_3855);
nor U4792 (N_4792,N_2858,N_2188);
xnor U4793 (N_4793,N_3332,N_2107);
and U4794 (N_4794,N_2224,N_3142);
or U4795 (N_4795,N_3033,N_2594);
xnor U4796 (N_4796,N_3039,N_2320);
nor U4797 (N_4797,N_2451,N_3373);
nor U4798 (N_4798,N_3319,N_2244);
nand U4799 (N_4799,N_2831,N_3754);
nand U4800 (N_4800,N_2978,N_2118);
nor U4801 (N_4801,N_3716,N_2390);
xor U4802 (N_4802,N_2116,N_3725);
nor U4803 (N_4803,N_3281,N_2238);
and U4804 (N_4804,N_3671,N_2243);
nor U4805 (N_4805,N_2585,N_3957);
nand U4806 (N_4806,N_2736,N_2459);
and U4807 (N_4807,N_3969,N_2101);
nand U4808 (N_4808,N_3204,N_2877);
nor U4809 (N_4809,N_2400,N_3837);
nand U4810 (N_4810,N_3505,N_3940);
or U4811 (N_4811,N_2889,N_2363);
and U4812 (N_4812,N_2089,N_2802);
and U4813 (N_4813,N_3531,N_2979);
and U4814 (N_4814,N_2265,N_3258);
nand U4815 (N_4815,N_3998,N_2810);
xnor U4816 (N_4816,N_2598,N_2658);
xor U4817 (N_4817,N_3006,N_2981);
xor U4818 (N_4818,N_2795,N_2429);
or U4819 (N_4819,N_3274,N_3682);
nand U4820 (N_4820,N_3967,N_3377);
xor U4821 (N_4821,N_2974,N_3939);
and U4822 (N_4822,N_3139,N_2179);
or U4823 (N_4823,N_3455,N_2087);
or U4824 (N_4824,N_2732,N_2108);
nor U4825 (N_4825,N_3607,N_2050);
and U4826 (N_4826,N_2669,N_2301);
and U4827 (N_4827,N_2047,N_2409);
or U4828 (N_4828,N_3578,N_3076);
or U4829 (N_4829,N_2234,N_2998);
and U4830 (N_4830,N_3135,N_3491);
and U4831 (N_4831,N_2533,N_2564);
nor U4832 (N_4832,N_2604,N_3117);
nor U4833 (N_4833,N_2825,N_3783);
nand U4834 (N_4834,N_2975,N_3343);
nand U4835 (N_4835,N_3620,N_2251);
or U4836 (N_4836,N_3562,N_2210);
or U4837 (N_4837,N_3698,N_3510);
nor U4838 (N_4838,N_3763,N_3436);
or U4839 (N_4839,N_2584,N_3108);
xnor U4840 (N_4840,N_3789,N_2636);
or U4841 (N_4841,N_3303,N_2544);
and U4842 (N_4842,N_2351,N_2406);
nand U4843 (N_4843,N_2648,N_2403);
nand U4844 (N_4844,N_2457,N_3457);
nand U4845 (N_4845,N_2374,N_2259);
nand U4846 (N_4846,N_2500,N_2680);
xnor U4847 (N_4847,N_2883,N_3481);
nor U4848 (N_4848,N_3880,N_3215);
or U4849 (N_4849,N_2190,N_2935);
nand U4850 (N_4850,N_3853,N_2424);
and U4851 (N_4851,N_2853,N_3399);
or U4852 (N_4852,N_3165,N_2416);
nand U4853 (N_4853,N_3323,N_2609);
or U4854 (N_4854,N_2693,N_2787);
xnor U4855 (N_4855,N_2342,N_3075);
xor U4856 (N_4856,N_3362,N_2568);
and U4857 (N_4857,N_3138,N_2148);
nor U4858 (N_4858,N_3497,N_2904);
nand U4859 (N_4859,N_3238,N_2132);
and U4860 (N_4860,N_3762,N_3393);
and U4861 (N_4861,N_3198,N_3298);
nand U4862 (N_4862,N_3470,N_2809);
nor U4863 (N_4863,N_2360,N_3444);
xor U4864 (N_4864,N_2164,N_2769);
nand U4865 (N_4865,N_2909,N_2632);
or U4866 (N_4866,N_2744,N_2274);
or U4867 (N_4867,N_2560,N_3951);
nand U4868 (N_4868,N_2402,N_3046);
nor U4869 (N_4869,N_3241,N_2772);
xor U4870 (N_4870,N_2053,N_2253);
nor U4871 (N_4871,N_2153,N_2576);
nor U4872 (N_4872,N_3686,N_2965);
nor U4873 (N_4873,N_3475,N_3739);
nand U4874 (N_4874,N_3292,N_3704);
or U4875 (N_4875,N_3175,N_3041);
and U4876 (N_4876,N_2310,N_2524);
xnor U4877 (N_4877,N_2936,N_3658);
xnor U4878 (N_4878,N_3832,N_2971);
or U4879 (N_4879,N_2007,N_2932);
and U4880 (N_4880,N_3570,N_2479);
or U4881 (N_4881,N_2393,N_3895);
or U4882 (N_4882,N_2977,N_2021);
nand U4883 (N_4883,N_3545,N_3526);
or U4884 (N_4884,N_3311,N_3743);
or U4885 (N_4885,N_2530,N_3706);
nor U4886 (N_4886,N_3301,N_3821);
nor U4887 (N_4887,N_3184,N_3385);
nor U4888 (N_4888,N_2728,N_3462);
and U4889 (N_4889,N_2333,N_3195);
nor U4890 (N_4890,N_2808,N_3340);
nand U4891 (N_4891,N_3966,N_3030);
nor U4892 (N_4892,N_3023,N_3736);
xnor U4893 (N_4893,N_3438,N_3351);
or U4894 (N_4894,N_2638,N_3687);
nor U4895 (N_4895,N_3010,N_2016);
or U4896 (N_4896,N_3663,N_3779);
nand U4897 (N_4897,N_2203,N_2045);
and U4898 (N_4898,N_3051,N_3861);
and U4899 (N_4899,N_3064,N_3202);
and U4900 (N_4900,N_3128,N_2282);
or U4901 (N_4901,N_3467,N_2634);
nor U4902 (N_4902,N_3984,N_2361);
nand U4903 (N_4903,N_2876,N_3733);
or U4904 (N_4904,N_3370,N_2448);
or U4905 (N_4905,N_2014,N_3884);
xnor U4906 (N_4906,N_2745,N_2521);
or U4907 (N_4907,N_2514,N_3712);
or U4908 (N_4908,N_2668,N_3613);
or U4909 (N_4909,N_2967,N_3480);
and U4910 (N_4910,N_3848,N_3593);
and U4911 (N_4911,N_2191,N_3820);
nand U4912 (N_4912,N_2359,N_2376);
and U4913 (N_4913,N_2395,N_2854);
xnor U4914 (N_4914,N_3307,N_2452);
nor U4915 (N_4915,N_2260,N_3070);
or U4916 (N_4916,N_2605,N_3655);
or U4917 (N_4917,N_2765,N_2092);
xor U4918 (N_4918,N_3416,N_2477);
and U4919 (N_4919,N_3256,N_2804);
nor U4920 (N_4920,N_2257,N_2836);
xnor U4921 (N_4921,N_3879,N_2198);
nand U4922 (N_4922,N_2601,N_2913);
or U4923 (N_4923,N_2969,N_2391);
nand U4924 (N_4924,N_3284,N_3995);
or U4925 (N_4925,N_3606,N_3391);
or U4926 (N_4926,N_2064,N_2405);
xnor U4927 (N_4927,N_2270,N_2156);
nor U4928 (N_4928,N_2557,N_3670);
nand U4929 (N_4929,N_2465,N_2004);
xnor U4930 (N_4930,N_3445,N_3465);
or U4931 (N_4931,N_3183,N_3921);
and U4932 (N_4932,N_3021,N_2647);
and U4933 (N_4933,N_2624,N_3928);
and U4934 (N_4934,N_2366,N_3037);
nand U4935 (N_4935,N_3286,N_2657);
nor U4936 (N_4936,N_2254,N_2221);
or U4937 (N_4937,N_2321,N_3269);
and U4938 (N_4938,N_2612,N_3101);
xnor U4939 (N_4939,N_2058,N_3123);
and U4940 (N_4940,N_2692,N_2755);
or U4941 (N_4941,N_2071,N_3993);
nand U4942 (N_4942,N_3035,N_3366);
xor U4943 (N_4943,N_2289,N_3574);
and U4944 (N_4944,N_2237,N_2206);
or U4945 (N_4945,N_3808,N_3100);
nand U4946 (N_4946,N_3584,N_2855);
or U4947 (N_4947,N_3050,N_3805);
or U4948 (N_4948,N_3666,N_3012);
nor U4949 (N_4949,N_3621,N_2887);
xor U4950 (N_4950,N_3025,N_2085);
and U4951 (N_4951,N_2499,N_3314);
nor U4952 (N_4952,N_2449,N_2957);
or U4953 (N_4953,N_2905,N_2388);
nor U4954 (N_4954,N_2903,N_3552);
nor U4955 (N_4955,N_3849,N_2450);
nor U4956 (N_4956,N_3120,N_2832);
or U4957 (N_4957,N_2034,N_3931);
or U4958 (N_4958,N_3386,N_2440);
xnor U4959 (N_4959,N_3559,N_2958);
and U4960 (N_4960,N_2273,N_3232);
xnor U4961 (N_4961,N_2724,N_3521);
xnor U4962 (N_4962,N_3959,N_2217);
xor U4963 (N_4963,N_2081,N_2205);
nor U4964 (N_4964,N_3707,N_3955);
nor U4965 (N_4965,N_2378,N_2656);
nand U4966 (N_4966,N_2725,N_3375);
nor U4967 (N_4967,N_3084,N_3265);
nor U4968 (N_4968,N_3857,N_2487);
nand U4969 (N_4969,N_2677,N_3089);
or U4970 (N_4970,N_2573,N_3835);
nand U4971 (N_4971,N_2646,N_3496);
nand U4972 (N_4972,N_3941,N_3824);
xor U4973 (N_4973,N_3854,N_2569);
xnor U4974 (N_4974,N_2115,N_2780);
or U4975 (N_4975,N_3273,N_2184);
and U4976 (N_4976,N_3081,N_3514);
nor U4977 (N_4977,N_2369,N_3134);
xnor U4978 (N_4978,N_3017,N_3942);
or U4979 (N_4979,N_2997,N_2158);
or U4980 (N_4980,N_3472,N_3112);
nand U4981 (N_4981,N_3960,N_3601);
and U4982 (N_4982,N_3537,N_3867);
nand U4983 (N_4983,N_3722,N_3858);
nor U4984 (N_4984,N_3324,N_3451);
or U4985 (N_4985,N_3390,N_3877);
nand U4986 (N_4986,N_3546,N_3127);
and U4987 (N_4987,N_3868,N_3535);
nor U4988 (N_4988,N_3622,N_3473);
or U4989 (N_4989,N_2869,N_3558);
nor U4990 (N_4990,N_3513,N_3255);
or U4991 (N_4991,N_3751,N_2446);
and U4992 (N_4992,N_3077,N_2999);
and U4993 (N_4993,N_2837,N_2941);
xnor U4994 (N_4994,N_2980,N_2013);
xor U4995 (N_4995,N_3034,N_3317);
xor U4996 (N_4996,N_3692,N_2219);
nand U4997 (N_4997,N_3982,N_2375);
or U4998 (N_4998,N_3874,N_3493);
or U4999 (N_4999,N_2370,N_3912);
or U5000 (N_5000,N_3841,N_2909);
nand U5001 (N_5001,N_2192,N_2092);
nor U5002 (N_5002,N_3460,N_2831);
and U5003 (N_5003,N_2574,N_2303);
nor U5004 (N_5004,N_3603,N_2615);
nor U5005 (N_5005,N_3988,N_3939);
and U5006 (N_5006,N_2792,N_3943);
nand U5007 (N_5007,N_3783,N_3452);
and U5008 (N_5008,N_2507,N_2733);
and U5009 (N_5009,N_2236,N_2531);
xnor U5010 (N_5010,N_3680,N_2988);
nand U5011 (N_5011,N_2337,N_2632);
xnor U5012 (N_5012,N_2066,N_2742);
and U5013 (N_5013,N_2500,N_2995);
nor U5014 (N_5014,N_2768,N_2701);
nand U5015 (N_5015,N_2790,N_3620);
nand U5016 (N_5016,N_3069,N_3566);
xnor U5017 (N_5017,N_2031,N_3302);
xor U5018 (N_5018,N_3273,N_2760);
xor U5019 (N_5019,N_3467,N_2987);
or U5020 (N_5020,N_3785,N_2119);
and U5021 (N_5021,N_3247,N_3545);
and U5022 (N_5022,N_2958,N_3706);
nor U5023 (N_5023,N_2303,N_3699);
and U5024 (N_5024,N_2458,N_3216);
nand U5025 (N_5025,N_3528,N_2795);
nand U5026 (N_5026,N_2061,N_3770);
nor U5027 (N_5027,N_2359,N_2466);
or U5028 (N_5028,N_3352,N_3458);
and U5029 (N_5029,N_2575,N_3273);
xor U5030 (N_5030,N_3614,N_3975);
xor U5031 (N_5031,N_2913,N_2277);
nor U5032 (N_5032,N_3085,N_3684);
and U5033 (N_5033,N_3091,N_3134);
xor U5034 (N_5034,N_3529,N_2651);
and U5035 (N_5035,N_2781,N_3712);
nand U5036 (N_5036,N_2494,N_2836);
or U5037 (N_5037,N_2822,N_3299);
xor U5038 (N_5038,N_3487,N_3541);
or U5039 (N_5039,N_3446,N_2026);
or U5040 (N_5040,N_3816,N_2764);
nor U5041 (N_5041,N_3368,N_2809);
nand U5042 (N_5042,N_2490,N_3455);
or U5043 (N_5043,N_2735,N_2451);
nor U5044 (N_5044,N_3906,N_3315);
or U5045 (N_5045,N_3065,N_2999);
and U5046 (N_5046,N_2197,N_2417);
nor U5047 (N_5047,N_2374,N_2761);
and U5048 (N_5048,N_2739,N_3528);
xor U5049 (N_5049,N_3452,N_2617);
nand U5050 (N_5050,N_3938,N_2152);
nand U5051 (N_5051,N_3331,N_3189);
and U5052 (N_5052,N_3327,N_2852);
nor U5053 (N_5053,N_3258,N_3585);
nor U5054 (N_5054,N_2443,N_2301);
or U5055 (N_5055,N_3387,N_2050);
or U5056 (N_5056,N_2242,N_2341);
nor U5057 (N_5057,N_3526,N_2499);
and U5058 (N_5058,N_2572,N_2973);
or U5059 (N_5059,N_3899,N_3906);
and U5060 (N_5060,N_3239,N_2290);
or U5061 (N_5061,N_2230,N_3013);
nor U5062 (N_5062,N_2068,N_3462);
xor U5063 (N_5063,N_3231,N_3613);
xor U5064 (N_5064,N_3229,N_2808);
or U5065 (N_5065,N_2425,N_2094);
and U5066 (N_5066,N_2239,N_3393);
nor U5067 (N_5067,N_3404,N_2552);
xnor U5068 (N_5068,N_3446,N_3898);
nand U5069 (N_5069,N_3713,N_3858);
or U5070 (N_5070,N_2553,N_2601);
or U5071 (N_5071,N_3023,N_2526);
nor U5072 (N_5072,N_3944,N_3219);
and U5073 (N_5073,N_3102,N_2704);
nand U5074 (N_5074,N_2821,N_3409);
nand U5075 (N_5075,N_3476,N_2861);
and U5076 (N_5076,N_2786,N_2898);
or U5077 (N_5077,N_3263,N_3176);
xor U5078 (N_5078,N_2356,N_3805);
and U5079 (N_5079,N_3687,N_3970);
and U5080 (N_5080,N_2790,N_3102);
xnor U5081 (N_5081,N_2342,N_2096);
nor U5082 (N_5082,N_2827,N_2007);
xor U5083 (N_5083,N_2419,N_3116);
nand U5084 (N_5084,N_3519,N_2344);
nand U5085 (N_5085,N_2582,N_2472);
or U5086 (N_5086,N_2383,N_3335);
nor U5087 (N_5087,N_2937,N_2891);
nand U5088 (N_5088,N_3645,N_2557);
or U5089 (N_5089,N_2055,N_2821);
nor U5090 (N_5090,N_3443,N_2943);
or U5091 (N_5091,N_3862,N_2685);
and U5092 (N_5092,N_3657,N_2137);
and U5093 (N_5093,N_3146,N_2045);
or U5094 (N_5094,N_2225,N_3974);
xor U5095 (N_5095,N_3799,N_2004);
nor U5096 (N_5096,N_2167,N_3637);
nand U5097 (N_5097,N_2174,N_3590);
or U5098 (N_5098,N_2359,N_2320);
or U5099 (N_5099,N_2022,N_3897);
nand U5100 (N_5100,N_2748,N_3867);
or U5101 (N_5101,N_2184,N_3003);
xnor U5102 (N_5102,N_3159,N_2169);
xnor U5103 (N_5103,N_2061,N_3830);
and U5104 (N_5104,N_2405,N_3347);
xnor U5105 (N_5105,N_3172,N_3614);
and U5106 (N_5106,N_3927,N_2983);
or U5107 (N_5107,N_2870,N_2766);
nor U5108 (N_5108,N_3705,N_3112);
and U5109 (N_5109,N_2626,N_3001);
or U5110 (N_5110,N_2013,N_2131);
xnor U5111 (N_5111,N_3223,N_2059);
or U5112 (N_5112,N_2859,N_2180);
nor U5113 (N_5113,N_3552,N_3761);
nand U5114 (N_5114,N_2881,N_3904);
nand U5115 (N_5115,N_2386,N_2814);
nor U5116 (N_5116,N_3405,N_2478);
nor U5117 (N_5117,N_3254,N_3109);
nor U5118 (N_5118,N_2280,N_2938);
or U5119 (N_5119,N_2936,N_2696);
nand U5120 (N_5120,N_3727,N_3510);
and U5121 (N_5121,N_3383,N_2354);
nand U5122 (N_5122,N_3044,N_3204);
nand U5123 (N_5123,N_3319,N_2341);
and U5124 (N_5124,N_3695,N_2876);
or U5125 (N_5125,N_2190,N_3887);
nand U5126 (N_5126,N_3063,N_3284);
nor U5127 (N_5127,N_3644,N_2054);
and U5128 (N_5128,N_2126,N_2739);
nand U5129 (N_5129,N_3647,N_2498);
and U5130 (N_5130,N_2690,N_3110);
nand U5131 (N_5131,N_3263,N_2813);
and U5132 (N_5132,N_2822,N_2234);
or U5133 (N_5133,N_3459,N_2345);
nand U5134 (N_5134,N_2734,N_3613);
nand U5135 (N_5135,N_2664,N_3580);
nand U5136 (N_5136,N_2828,N_2778);
nand U5137 (N_5137,N_2091,N_3359);
nor U5138 (N_5138,N_2287,N_3805);
xor U5139 (N_5139,N_3156,N_2988);
nor U5140 (N_5140,N_3287,N_2303);
and U5141 (N_5141,N_3516,N_2519);
xor U5142 (N_5142,N_3308,N_3939);
nand U5143 (N_5143,N_2356,N_2917);
nor U5144 (N_5144,N_3393,N_3768);
or U5145 (N_5145,N_2421,N_2308);
nor U5146 (N_5146,N_2078,N_3323);
xor U5147 (N_5147,N_3032,N_3061);
nor U5148 (N_5148,N_2390,N_2113);
xnor U5149 (N_5149,N_3485,N_2989);
xor U5150 (N_5150,N_2690,N_3316);
xnor U5151 (N_5151,N_2667,N_3565);
xnor U5152 (N_5152,N_2822,N_2478);
or U5153 (N_5153,N_2141,N_2249);
nor U5154 (N_5154,N_3836,N_3700);
xor U5155 (N_5155,N_3097,N_3428);
xor U5156 (N_5156,N_2700,N_2250);
nor U5157 (N_5157,N_2563,N_3974);
nor U5158 (N_5158,N_3223,N_2277);
or U5159 (N_5159,N_2764,N_2850);
nor U5160 (N_5160,N_3886,N_2664);
and U5161 (N_5161,N_3274,N_3226);
or U5162 (N_5162,N_3194,N_2291);
or U5163 (N_5163,N_2882,N_3441);
nand U5164 (N_5164,N_3595,N_3225);
nand U5165 (N_5165,N_2639,N_2789);
xor U5166 (N_5166,N_2248,N_2179);
xnor U5167 (N_5167,N_2326,N_3346);
and U5168 (N_5168,N_2258,N_3517);
nand U5169 (N_5169,N_3893,N_2555);
xor U5170 (N_5170,N_3455,N_2001);
nor U5171 (N_5171,N_3793,N_3581);
nand U5172 (N_5172,N_2898,N_3149);
and U5173 (N_5173,N_2111,N_2540);
nor U5174 (N_5174,N_2544,N_2997);
nor U5175 (N_5175,N_3290,N_3820);
nor U5176 (N_5176,N_2296,N_3533);
nand U5177 (N_5177,N_3859,N_3238);
nor U5178 (N_5178,N_3439,N_3863);
xnor U5179 (N_5179,N_2222,N_3754);
xor U5180 (N_5180,N_2800,N_3566);
nand U5181 (N_5181,N_3700,N_3641);
nand U5182 (N_5182,N_3274,N_3875);
nand U5183 (N_5183,N_2045,N_3728);
nor U5184 (N_5184,N_3491,N_3607);
and U5185 (N_5185,N_2356,N_3463);
and U5186 (N_5186,N_3274,N_3849);
or U5187 (N_5187,N_3116,N_3535);
xor U5188 (N_5188,N_3480,N_2963);
or U5189 (N_5189,N_3543,N_3213);
nand U5190 (N_5190,N_2027,N_3123);
nor U5191 (N_5191,N_2751,N_2646);
or U5192 (N_5192,N_3856,N_3137);
and U5193 (N_5193,N_3198,N_3507);
and U5194 (N_5194,N_2548,N_2319);
nor U5195 (N_5195,N_3479,N_2684);
xor U5196 (N_5196,N_2098,N_3954);
or U5197 (N_5197,N_2312,N_2903);
xor U5198 (N_5198,N_2105,N_2682);
nand U5199 (N_5199,N_3810,N_2870);
xnor U5200 (N_5200,N_3247,N_3034);
or U5201 (N_5201,N_2794,N_3852);
nor U5202 (N_5202,N_2267,N_2425);
nand U5203 (N_5203,N_2965,N_3298);
nand U5204 (N_5204,N_3683,N_2702);
or U5205 (N_5205,N_3556,N_3757);
or U5206 (N_5206,N_3046,N_3709);
nor U5207 (N_5207,N_3844,N_2033);
nand U5208 (N_5208,N_2981,N_3320);
nor U5209 (N_5209,N_3969,N_3650);
or U5210 (N_5210,N_3538,N_3466);
xnor U5211 (N_5211,N_2144,N_3254);
and U5212 (N_5212,N_3158,N_2086);
and U5213 (N_5213,N_3070,N_3878);
xor U5214 (N_5214,N_3152,N_3784);
nand U5215 (N_5215,N_2001,N_2027);
and U5216 (N_5216,N_3177,N_3716);
nand U5217 (N_5217,N_3050,N_3486);
or U5218 (N_5218,N_2859,N_3175);
nor U5219 (N_5219,N_2019,N_3234);
xor U5220 (N_5220,N_3150,N_2376);
and U5221 (N_5221,N_2012,N_3288);
xor U5222 (N_5222,N_3548,N_2218);
or U5223 (N_5223,N_2560,N_3267);
and U5224 (N_5224,N_3007,N_2201);
xnor U5225 (N_5225,N_3290,N_2864);
or U5226 (N_5226,N_2543,N_3902);
xnor U5227 (N_5227,N_3478,N_3116);
xnor U5228 (N_5228,N_2019,N_3459);
or U5229 (N_5229,N_3567,N_3029);
nand U5230 (N_5230,N_3641,N_2138);
nor U5231 (N_5231,N_3349,N_3097);
nor U5232 (N_5232,N_3892,N_3801);
nor U5233 (N_5233,N_3743,N_2062);
nor U5234 (N_5234,N_3211,N_3129);
xor U5235 (N_5235,N_2888,N_2348);
nor U5236 (N_5236,N_2934,N_3185);
nor U5237 (N_5237,N_3762,N_2124);
nand U5238 (N_5238,N_3352,N_3054);
xor U5239 (N_5239,N_2452,N_2999);
nor U5240 (N_5240,N_2524,N_3320);
nand U5241 (N_5241,N_3037,N_3877);
xor U5242 (N_5242,N_3223,N_3512);
nor U5243 (N_5243,N_3703,N_2555);
nor U5244 (N_5244,N_2879,N_3061);
nand U5245 (N_5245,N_3521,N_3016);
nor U5246 (N_5246,N_2832,N_2558);
nor U5247 (N_5247,N_2770,N_2040);
and U5248 (N_5248,N_3971,N_3615);
and U5249 (N_5249,N_3958,N_3500);
xnor U5250 (N_5250,N_3287,N_3339);
or U5251 (N_5251,N_3948,N_3241);
nor U5252 (N_5252,N_3042,N_2928);
and U5253 (N_5253,N_3895,N_2017);
or U5254 (N_5254,N_3888,N_3278);
nor U5255 (N_5255,N_2179,N_3167);
nand U5256 (N_5256,N_2346,N_3704);
xor U5257 (N_5257,N_2299,N_3084);
nand U5258 (N_5258,N_3189,N_2275);
nor U5259 (N_5259,N_2206,N_3685);
and U5260 (N_5260,N_3189,N_2983);
xnor U5261 (N_5261,N_2883,N_2870);
and U5262 (N_5262,N_2690,N_2686);
or U5263 (N_5263,N_3041,N_3805);
nand U5264 (N_5264,N_2879,N_3563);
or U5265 (N_5265,N_3504,N_2799);
xor U5266 (N_5266,N_3242,N_2358);
nand U5267 (N_5267,N_2173,N_3442);
nor U5268 (N_5268,N_2009,N_2645);
nor U5269 (N_5269,N_2158,N_3580);
and U5270 (N_5270,N_3409,N_2442);
nor U5271 (N_5271,N_2434,N_2354);
and U5272 (N_5272,N_3225,N_2751);
and U5273 (N_5273,N_2963,N_3867);
and U5274 (N_5274,N_3215,N_3220);
xnor U5275 (N_5275,N_2466,N_2606);
xnor U5276 (N_5276,N_2107,N_2592);
xnor U5277 (N_5277,N_3455,N_2980);
xnor U5278 (N_5278,N_3652,N_2816);
nor U5279 (N_5279,N_3308,N_3163);
xnor U5280 (N_5280,N_3885,N_3708);
xor U5281 (N_5281,N_2409,N_3370);
and U5282 (N_5282,N_3023,N_3184);
nor U5283 (N_5283,N_3371,N_3058);
nor U5284 (N_5284,N_2872,N_2235);
xnor U5285 (N_5285,N_3694,N_3148);
or U5286 (N_5286,N_3242,N_3537);
xor U5287 (N_5287,N_2272,N_3056);
nand U5288 (N_5288,N_3053,N_3168);
or U5289 (N_5289,N_3910,N_2347);
and U5290 (N_5290,N_2113,N_3258);
nand U5291 (N_5291,N_3965,N_3608);
nand U5292 (N_5292,N_2165,N_3992);
nand U5293 (N_5293,N_2115,N_3114);
and U5294 (N_5294,N_2846,N_2572);
nor U5295 (N_5295,N_3433,N_3885);
nand U5296 (N_5296,N_2447,N_3986);
xor U5297 (N_5297,N_2721,N_2360);
or U5298 (N_5298,N_3282,N_2842);
nand U5299 (N_5299,N_3488,N_3399);
or U5300 (N_5300,N_2127,N_3339);
nand U5301 (N_5301,N_2653,N_3189);
and U5302 (N_5302,N_2751,N_3704);
xor U5303 (N_5303,N_3568,N_3985);
and U5304 (N_5304,N_2265,N_3974);
xor U5305 (N_5305,N_3968,N_3444);
nand U5306 (N_5306,N_3042,N_2184);
and U5307 (N_5307,N_2937,N_3969);
nor U5308 (N_5308,N_3691,N_3206);
or U5309 (N_5309,N_3506,N_2599);
xnor U5310 (N_5310,N_3630,N_2365);
nor U5311 (N_5311,N_2409,N_2157);
and U5312 (N_5312,N_3995,N_2188);
and U5313 (N_5313,N_3391,N_3658);
or U5314 (N_5314,N_2608,N_3382);
nand U5315 (N_5315,N_2353,N_2911);
nor U5316 (N_5316,N_3533,N_3116);
nor U5317 (N_5317,N_2338,N_2156);
nand U5318 (N_5318,N_2627,N_2316);
nor U5319 (N_5319,N_3362,N_2533);
and U5320 (N_5320,N_3735,N_3340);
and U5321 (N_5321,N_3878,N_3377);
or U5322 (N_5322,N_3847,N_2259);
xor U5323 (N_5323,N_2971,N_2824);
or U5324 (N_5324,N_3643,N_2128);
nor U5325 (N_5325,N_3724,N_3398);
nand U5326 (N_5326,N_2559,N_2884);
nor U5327 (N_5327,N_3997,N_3186);
or U5328 (N_5328,N_3303,N_2539);
xor U5329 (N_5329,N_3818,N_2816);
nand U5330 (N_5330,N_2865,N_2449);
nand U5331 (N_5331,N_3463,N_2447);
nand U5332 (N_5332,N_2747,N_2827);
nor U5333 (N_5333,N_2313,N_3895);
nand U5334 (N_5334,N_2062,N_3064);
nor U5335 (N_5335,N_3950,N_2771);
or U5336 (N_5336,N_2753,N_3377);
nor U5337 (N_5337,N_3472,N_2295);
nand U5338 (N_5338,N_3816,N_2675);
or U5339 (N_5339,N_2303,N_2511);
nand U5340 (N_5340,N_2040,N_3592);
nand U5341 (N_5341,N_2770,N_2672);
nor U5342 (N_5342,N_2295,N_2816);
xnor U5343 (N_5343,N_3673,N_2602);
and U5344 (N_5344,N_3446,N_3012);
or U5345 (N_5345,N_2054,N_2484);
or U5346 (N_5346,N_2500,N_2390);
nand U5347 (N_5347,N_3518,N_2964);
nor U5348 (N_5348,N_3729,N_2348);
nor U5349 (N_5349,N_2618,N_2630);
xor U5350 (N_5350,N_3163,N_2200);
nand U5351 (N_5351,N_3037,N_3482);
and U5352 (N_5352,N_2122,N_2924);
and U5353 (N_5353,N_3408,N_2431);
xnor U5354 (N_5354,N_2273,N_2166);
nor U5355 (N_5355,N_2287,N_2493);
nor U5356 (N_5356,N_2308,N_2767);
xnor U5357 (N_5357,N_3305,N_2240);
nand U5358 (N_5358,N_3598,N_2736);
nor U5359 (N_5359,N_2558,N_3113);
nand U5360 (N_5360,N_2746,N_2790);
or U5361 (N_5361,N_2005,N_3072);
or U5362 (N_5362,N_3912,N_2175);
nand U5363 (N_5363,N_2404,N_3524);
and U5364 (N_5364,N_2290,N_3843);
nand U5365 (N_5365,N_3770,N_3484);
and U5366 (N_5366,N_2733,N_2689);
nor U5367 (N_5367,N_3270,N_3850);
and U5368 (N_5368,N_2953,N_2015);
and U5369 (N_5369,N_2820,N_2636);
or U5370 (N_5370,N_3962,N_3072);
or U5371 (N_5371,N_2228,N_2007);
nand U5372 (N_5372,N_2280,N_3496);
nor U5373 (N_5373,N_3873,N_3286);
and U5374 (N_5374,N_2643,N_3789);
nand U5375 (N_5375,N_3540,N_3239);
or U5376 (N_5376,N_3632,N_2033);
nand U5377 (N_5377,N_3762,N_3446);
xnor U5378 (N_5378,N_3729,N_3639);
nor U5379 (N_5379,N_2701,N_2881);
nor U5380 (N_5380,N_3390,N_2902);
nand U5381 (N_5381,N_2064,N_3141);
or U5382 (N_5382,N_2141,N_2064);
nor U5383 (N_5383,N_2995,N_2149);
xnor U5384 (N_5384,N_2818,N_3062);
xor U5385 (N_5385,N_2455,N_3988);
xnor U5386 (N_5386,N_3672,N_2511);
or U5387 (N_5387,N_3107,N_2716);
nand U5388 (N_5388,N_2489,N_3848);
xor U5389 (N_5389,N_2420,N_3155);
nand U5390 (N_5390,N_2124,N_2534);
nand U5391 (N_5391,N_2240,N_3332);
or U5392 (N_5392,N_2105,N_2311);
xor U5393 (N_5393,N_2473,N_3753);
and U5394 (N_5394,N_2484,N_2282);
nand U5395 (N_5395,N_2726,N_2476);
or U5396 (N_5396,N_3949,N_3484);
xnor U5397 (N_5397,N_3978,N_2816);
and U5398 (N_5398,N_2581,N_3070);
xor U5399 (N_5399,N_2183,N_2643);
or U5400 (N_5400,N_2621,N_3161);
nand U5401 (N_5401,N_2375,N_2019);
nor U5402 (N_5402,N_3163,N_3004);
nor U5403 (N_5403,N_3213,N_2773);
xnor U5404 (N_5404,N_3544,N_3331);
or U5405 (N_5405,N_2516,N_2464);
xnor U5406 (N_5406,N_2596,N_3573);
and U5407 (N_5407,N_2534,N_2127);
nand U5408 (N_5408,N_2928,N_2881);
or U5409 (N_5409,N_2997,N_2730);
xor U5410 (N_5410,N_3758,N_3876);
nand U5411 (N_5411,N_2975,N_2391);
xnor U5412 (N_5412,N_3382,N_3672);
xor U5413 (N_5413,N_3177,N_3452);
and U5414 (N_5414,N_2958,N_2722);
nor U5415 (N_5415,N_2524,N_2591);
nand U5416 (N_5416,N_2251,N_2693);
nor U5417 (N_5417,N_3723,N_2623);
and U5418 (N_5418,N_2620,N_2807);
nor U5419 (N_5419,N_2996,N_2726);
or U5420 (N_5420,N_3237,N_2207);
xnor U5421 (N_5421,N_2677,N_2604);
xor U5422 (N_5422,N_2802,N_2975);
nand U5423 (N_5423,N_2767,N_3039);
and U5424 (N_5424,N_2507,N_2460);
nand U5425 (N_5425,N_3704,N_2857);
nor U5426 (N_5426,N_3325,N_2552);
xor U5427 (N_5427,N_3420,N_2897);
xor U5428 (N_5428,N_3746,N_2308);
or U5429 (N_5429,N_3361,N_3642);
or U5430 (N_5430,N_2643,N_2760);
nor U5431 (N_5431,N_2877,N_2392);
or U5432 (N_5432,N_2428,N_2506);
and U5433 (N_5433,N_3572,N_2438);
and U5434 (N_5434,N_3660,N_2209);
nand U5435 (N_5435,N_2232,N_3845);
and U5436 (N_5436,N_2977,N_3134);
or U5437 (N_5437,N_2847,N_3221);
xnor U5438 (N_5438,N_3791,N_3286);
or U5439 (N_5439,N_2198,N_3093);
nor U5440 (N_5440,N_2151,N_2512);
or U5441 (N_5441,N_3001,N_2732);
xor U5442 (N_5442,N_2714,N_3262);
nand U5443 (N_5443,N_2499,N_2945);
nand U5444 (N_5444,N_2782,N_2759);
nand U5445 (N_5445,N_3311,N_3470);
nor U5446 (N_5446,N_3123,N_3263);
nor U5447 (N_5447,N_2406,N_3988);
nand U5448 (N_5448,N_2307,N_2582);
or U5449 (N_5449,N_2183,N_3615);
and U5450 (N_5450,N_2841,N_2668);
xor U5451 (N_5451,N_3807,N_3587);
nor U5452 (N_5452,N_3246,N_3302);
and U5453 (N_5453,N_2059,N_3678);
nor U5454 (N_5454,N_2547,N_3819);
nor U5455 (N_5455,N_2906,N_2173);
nor U5456 (N_5456,N_2083,N_2362);
xor U5457 (N_5457,N_2304,N_3288);
and U5458 (N_5458,N_3935,N_2099);
nor U5459 (N_5459,N_2227,N_3630);
nor U5460 (N_5460,N_3269,N_3378);
and U5461 (N_5461,N_2177,N_3983);
nand U5462 (N_5462,N_2147,N_2059);
or U5463 (N_5463,N_2655,N_2860);
xnor U5464 (N_5464,N_2642,N_3151);
xnor U5465 (N_5465,N_2033,N_3765);
and U5466 (N_5466,N_2722,N_2111);
or U5467 (N_5467,N_2308,N_3980);
nor U5468 (N_5468,N_3077,N_2321);
or U5469 (N_5469,N_3206,N_3936);
nand U5470 (N_5470,N_3238,N_2808);
xor U5471 (N_5471,N_3480,N_2465);
xnor U5472 (N_5472,N_2531,N_3445);
or U5473 (N_5473,N_3332,N_3073);
nand U5474 (N_5474,N_3248,N_3511);
nand U5475 (N_5475,N_3193,N_3485);
nand U5476 (N_5476,N_2805,N_3176);
and U5477 (N_5477,N_2087,N_2280);
nor U5478 (N_5478,N_3967,N_2500);
xnor U5479 (N_5479,N_3729,N_3955);
nor U5480 (N_5480,N_2418,N_2838);
and U5481 (N_5481,N_2502,N_2641);
and U5482 (N_5482,N_3750,N_3412);
or U5483 (N_5483,N_2211,N_3199);
nor U5484 (N_5484,N_2761,N_3223);
xnor U5485 (N_5485,N_2507,N_2042);
nand U5486 (N_5486,N_2678,N_2277);
nor U5487 (N_5487,N_2645,N_3619);
or U5488 (N_5488,N_3243,N_3183);
or U5489 (N_5489,N_2276,N_3419);
nand U5490 (N_5490,N_2286,N_3709);
xnor U5491 (N_5491,N_2942,N_3495);
nor U5492 (N_5492,N_2227,N_3968);
nor U5493 (N_5493,N_2035,N_3131);
nor U5494 (N_5494,N_2965,N_3994);
nor U5495 (N_5495,N_3015,N_2689);
and U5496 (N_5496,N_3468,N_3413);
nand U5497 (N_5497,N_3484,N_2570);
nand U5498 (N_5498,N_2523,N_2222);
xnor U5499 (N_5499,N_3144,N_3719);
or U5500 (N_5500,N_3327,N_3949);
and U5501 (N_5501,N_2219,N_3357);
xor U5502 (N_5502,N_2717,N_3591);
xor U5503 (N_5503,N_2597,N_2047);
nand U5504 (N_5504,N_2392,N_3828);
nor U5505 (N_5505,N_2556,N_3271);
or U5506 (N_5506,N_3239,N_2664);
and U5507 (N_5507,N_3705,N_3379);
nor U5508 (N_5508,N_2300,N_3602);
or U5509 (N_5509,N_3369,N_2816);
nor U5510 (N_5510,N_3444,N_2816);
nor U5511 (N_5511,N_2142,N_3909);
and U5512 (N_5512,N_3479,N_3008);
or U5513 (N_5513,N_3186,N_3311);
and U5514 (N_5514,N_2048,N_3903);
nand U5515 (N_5515,N_3589,N_2127);
nand U5516 (N_5516,N_3017,N_2909);
nor U5517 (N_5517,N_3848,N_2818);
or U5518 (N_5518,N_3864,N_2925);
and U5519 (N_5519,N_2430,N_2802);
nand U5520 (N_5520,N_2485,N_2116);
xor U5521 (N_5521,N_2812,N_3515);
nor U5522 (N_5522,N_3623,N_2350);
and U5523 (N_5523,N_2975,N_2311);
nand U5524 (N_5524,N_2269,N_2855);
nor U5525 (N_5525,N_2937,N_3973);
nor U5526 (N_5526,N_3502,N_2687);
or U5527 (N_5527,N_2865,N_2934);
and U5528 (N_5528,N_3426,N_3096);
nand U5529 (N_5529,N_2221,N_3203);
nor U5530 (N_5530,N_3634,N_2922);
nand U5531 (N_5531,N_2746,N_3947);
or U5532 (N_5532,N_2791,N_2467);
or U5533 (N_5533,N_2861,N_3040);
and U5534 (N_5534,N_3066,N_3537);
nor U5535 (N_5535,N_2116,N_3964);
xnor U5536 (N_5536,N_2441,N_2455);
xor U5537 (N_5537,N_2924,N_2613);
and U5538 (N_5538,N_3035,N_3402);
nor U5539 (N_5539,N_3099,N_3762);
nand U5540 (N_5540,N_3111,N_2020);
nand U5541 (N_5541,N_2412,N_2663);
nand U5542 (N_5542,N_3699,N_3101);
nand U5543 (N_5543,N_2813,N_2246);
and U5544 (N_5544,N_2226,N_2770);
nor U5545 (N_5545,N_2128,N_3855);
xor U5546 (N_5546,N_3524,N_3239);
or U5547 (N_5547,N_2383,N_2404);
and U5548 (N_5548,N_2614,N_3087);
or U5549 (N_5549,N_2714,N_2947);
nand U5550 (N_5550,N_3735,N_3635);
nand U5551 (N_5551,N_3338,N_2633);
nor U5552 (N_5552,N_3021,N_2445);
and U5553 (N_5553,N_2540,N_2885);
or U5554 (N_5554,N_2092,N_3454);
and U5555 (N_5555,N_3671,N_3562);
or U5556 (N_5556,N_3654,N_2721);
or U5557 (N_5557,N_3480,N_2647);
nor U5558 (N_5558,N_2165,N_2812);
nand U5559 (N_5559,N_3887,N_3113);
and U5560 (N_5560,N_2602,N_3153);
nor U5561 (N_5561,N_2473,N_3266);
xor U5562 (N_5562,N_2039,N_3704);
nand U5563 (N_5563,N_3859,N_2839);
nand U5564 (N_5564,N_2317,N_2124);
nor U5565 (N_5565,N_3099,N_2868);
nor U5566 (N_5566,N_2844,N_2092);
nor U5567 (N_5567,N_2033,N_2981);
and U5568 (N_5568,N_3213,N_2165);
nand U5569 (N_5569,N_2435,N_3759);
nand U5570 (N_5570,N_2281,N_3427);
nor U5571 (N_5571,N_2242,N_2972);
nor U5572 (N_5572,N_3240,N_3800);
and U5573 (N_5573,N_3383,N_3421);
or U5574 (N_5574,N_3853,N_2048);
and U5575 (N_5575,N_3516,N_2556);
and U5576 (N_5576,N_2308,N_2759);
and U5577 (N_5577,N_3678,N_2113);
xor U5578 (N_5578,N_3330,N_2056);
and U5579 (N_5579,N_3329,N_2285);
or U5580 (N_5580,N_3326,N_3457);
or U5581 (N_5581,N_2256,N_2084);
xnor U5582 (N_5582,N_2022,N_3039);
xor U5583 (N_5583,N_3862,N_2198);
nand U5584 (N_5584,N_3910,N_2442);
nor U5585 (N_5585,N_2005,N_2752);
or U5586 (N_5586,N_2574,N_2062);
and U5587 (N_5587,N_2121,N_3905);
xor U5588 (N_5588,N_3566,N_3689);
nand U5589 (N_5589,N_2478,N_3154);
nand U5590 (N_5590,N_2450,N_2037);
or U5591 (N_5591,N_3689,N_2892);
or U5592 (N_5592,N_3139,N_3965);
or U5593 (N_5593,N_2486,N_2582);
nor U5594 (N_5594,N_2533,N_2529);
xnor U5595 (N_5595,N_2989,N_3532);
and U5596 (N_5596,N_3051,N_3848);
and U5597 (N_5597,N_2696,N_2087);
or U5598 (N_5598,N_2576,N_2495);
xnor U5599 (N_5599,N_3131,N_3252);
nand U5600 (N_5600,N_3146,N_3691);
or U5601 (N_5601,N_3479,N_3467);
nor U5602 (N_5602,N_3327,N_2548);
nand U5603 (N_5603,N_3601,N_2950);
nand U5604 (N_5604,N_2330,N_3685);
nor U5605 (N_5605,N_3349,N_2116);
and U5606 (N_5606,N_2160,N_3044);
xor U5607 (N_5607,N_3064,N_2005);
nor U5608 (N_5608,N_3242,N_2011);
xor U5609 (N_5609,N_3304,N_2434);
nand U5610 (N_5610,N_2022,N_3561);
nor U5611 (N_5611,N_3833,N_3319);
nor U5612 (N_5612,N_3330,N_2169);
nand U5613 (N_5613,N_3360,N_2870);
nor U5614 (N_5614,N_3369,N_2532);
nand U5615 (N_5615,N_3435,N_2583);
or U5616 (N_5616,N_3248,N_3384);
or U5617 (N_5617,N_3987,N_3710);
nor U5618 (N_5618,N_2409,N_3550);
nand U5619 (N_5619,N_2199,N_3101);
nand U5620 (N_5620,N_2170,N_2775);
nand U5621 (N_5621,N_3645,N_2707);
or U5622 (N_5622,N_3855,N_3528);
and U5623 (N_5623,N_2786,N_3044);
or U5624 (N_5624,N_3802,N_2419);
and U5625 (N_5625,N_3349,N_3262);
nor U5626 (N_5626,N_2451,N_3852);
nand U5627 (N_5627,N_3820,N_3354);
nor U5628 (N_5628,N_2593,N_2956);
and U5629 (N_5629,N_2393,N_3965);
xor U5630 (N_5630,N_3075,N_3448);
nor U5631 (N_5631,N_2100,N_2359);
xnor U5632 (N_5632,N_2791,N_2449);
xnor U5633 (N_5633,N_2469,N_3165);
nor U5634 (N_5634,N_2943,N_3661);
nand U5635 (N_5635,N_2552,N_2347);
nand U5636 (N_5636,N_2230,N_2373);
nor U5637 (N_5637,N_2232,N_3156);
nor U5638 (N_5638,N_2483,N_2304);
nor U5639 (N_5639,N_3181,N_2148);
and U5640 (N_5640,N_2453,N_2760);
nor U5641 (N_5641,N_3105,N_2068);
nor U5642 (N_5642,N_3143,N_3690);
or U5643 (N_5643,N_3841,N_2081);
nor U5644 (N_5644,N_3571,N_2372);
nor U5645 (N_5645,N_2440,N_3179);
and U5646 (N_5646,N_3237,N_2341);
or U5647 (N_5647,N_3474,N_3592);
and U5648 (N_5648,N_2940,N_2519);
nor U5649 (N_5649,N_2972,N_3014);
nand U5650 (N_5650,N_2129,N_3205);
or U5651 (N_5651,N_2264,N_3527);
xor U5652 (N_5652,N_3508,N_2015);
nor U5653 (N_5653,N_2323,N_2682);
xnor U5654 (N_5654,N_2593,N_3623);
nor U5655 (N_5655,N_2143,N_2316);
xor U5656 (N_5656,N_3376,N_2779);
and U5657 (N_5657,N_3337,N_3911);
or U5658 (N_5658,N_2726,N_3830);
nor U5659 (N_5659,N_3856,N_2525);
nand U5660 (N_5660,N_3964,N_2854);
nor U5661 (N_5661,N_2849,N_3496);
xor U5662 (N_5662,N_2086,N_3329);
nor U5663 (N_5663,N_3673,N_2053);
xnor U5664 (N_5664,N_2084,N_3885);
and U5665 (N_5665,N_2409,N_2845);
or U5666 (N_5666,N_3805,N_3947);
nand U5667 (N_5667,N_2467,N_3894);
xor U5668 (N_5668,N_3728,N_2559);
nand U5669 (N_5669,N_3778,N_3701);
xnor U5670 (N_5670,N_3757,N_2274);
nor U5671 (N_5671,N_3451,N_3944);
nand U5672 (N_5672,N_2062,N_3646);
nor U5673 (N_5673,N_3068,N_3322);
nor U5674 (N_5674,N_3347,N_2310);
nor U5675 (N_5675,N_3646,N_3107);
xnor U5676 (N_5676,N_2565,N_3319);
or U5677 (N_5677,N_2698,N_2551);
nand U5678 (N_5678,N_3627,N_3532);
xnor U5679 (N_5679,N_2685,N_2026);
nor U5680 (N_5680,N_2420,N_3962);
nor U5681 (N_5681,N_2695,N_2125);
nor U5682 (N_5682,N_2942,N_3618);
nor U5683 (N_5683,N_2168,N_2237);
and U5684 (N_5684,N_3491,N_2432);
and U5685 (N_5685,N_2696,N_2932);
xor U5686 (N_5686,N_2958,N_2171);
xnor U5687 (N_5687,N_2830,N_3426);
nor U5688 (N_5688,N_2994,N_3427);
and U5689 (N_5689,N_3212,N_3205);
nor U5690 (N_5690,N_3474,N_3745);
nor U5691 (N_5691,N_3236,N_3986);
nand U5692 (N_5692,N_2102,N_3296);
and U5693 (N_5693,N_3418,N_3092);
or U5694 (N_5694,N_2266,N_3621);
or U5695 (N_5695,N_3314,N_2912);
nand U5696 (N_5696,N_2945,N_2052);
xnor U5697 (N_5697,N_2113,N_2314);
and U5698 (N_5698,N_3770,N_2320);
and U5699 (N_5699,N_3264,N_3402);
nand U5700 (N_5700,N_2765,N_2904);
xnor U5701 (N_5701,N_3597,N_3818);
and U5702 (N_5702,N_2946,N_2939);
or U5703 (N_5703,N_2469,N_3474);
or U5704 (N_5704,N_2171,N_3775);
nor U5705 (N_5705,N_3406,N_2267);
xnor U5706 (N_5706,N_2336,N_2998);
and U5707 (N_5707,N_3422,N_3175);
nand U5708 (N_5708,N_3222,N_2841);
or U5709 (N_5709,N_2572,N_2205);
nor U5710 (N_5710,N_2106,N_3217);
nor U5711 (N_5711,N_2217,N_2493);
nor U5712 (N_5712,N_2833,N_2383);
nand U5713 (N_5713,N_3076,N_3741);
or U5714 (N_5714,N_2524,N_2058);
and U5715 (N_5715,N_2365,N_3703);
and U5716 (N_5716,N_2853,N_3277);
xor U5717 (N_5717,N_2914,N_2735);
or U5718 (N_5718,N_2994,N_3816);
nor U5719 (N_5719,N_3074,N_3673);
nand U5720 (N_5720,N_3058,N_3909);
nor U5721 (N_5721,N_3743,N_2958);
nor U5722 (N_5722,N_2750,N_2641);
xor U5723 (N_5723,N_3758,N_3584);
and U5724 (N_5724,N_2310,N_2165);
or U5725 (N_5725,N_2005,N_3195);
or U5726 (N_5726,N_2337,N_3535);
xnor U5727 (N_5727,N_2237,N_3306);
or U5728 (N_5728,N_3526,N_3510);
or U5729 (N_5729,N_2596,N_2348);
nand U5730 (N_5730,N_3686,N_2709);
or U5731 (N_5731,N_3751,N_2682);
xor U5732 (N_5732,N_2799,N_3094);
nand U5733 (N_5733,N_3642,N_2329);
nand U5734 (N_5734,N_2047,N_3939);
xnor U5735 (N_5735,N_2244,N_3844);
nand U5736 (N_5736,N_3407,N_2562);
or U5737 (N_5737,N_3491,N_2335);
and U5738 (N_5738,N_3500,N_3468);
nor U5739 (N_5739,N_2061,N_2943);
and U5740 (N_5740,N_2813,N_3713);
and U5741 (N_5741,N_2042,N_3711);
nor U5742 (N_5742,N_2337,N_2814);
nand U5743 (N_5743,N_2026,N_3714);
and U5744 (N_5744,N_2399,N_3326);
nand U5745 (N_5745,N_3586,N_3509);
nand U5746 (N_5746,N_2848,N_2215);
or U5747 (N_5747,N_3859,N_2402);
xnor U5748 (N_5748,N_2149,N_2537);
and U5749 (N_5749,N_3391,N_3345);
xnor U5750 (N_5750,N_2355,N_2936);
or U5751 (N_5751,N_2493,N_3285);
nand U5752 (N_5752,N_3624,N_3357);
or U5753 (N_5753,N_3152,N_2953);
or U5754 (N_5754,N_2109,N_2151);
nand U5755 (N_5755,N_2638,N_2080);
or U5756 (N_5756,N_2503,N_2537);
xor U5757 (N_5757,N_2802,N_2060);
and U5758 (N_5758,N_2219,N_3718);
nor U5759 (N_5759,N_2137,N_2899);
and U5760 (N_5760,N_3553,N_3281);
nor U5761 (N_5761,N_3831,N_2399);
xor U5762 (N_5762,N_3873,N_2198);
nand U5763 (N_5763,N_2394,N_2648);
nor U5764 (N_5764,N_2938,N_3195);
and U5765 (N_5765,N_3232,N_2918);
and U5766 (N_5766,N_2486,N_2096);
nor U5767 (N_5767,N_2027,N_3340);
nand U5768 (N_5768,N_2117,N_3544);
and U5769 (N_5769,N_2810,N_2561);
nand U5770 (N_5770,N_2831,N_2115);
and U5771 (N_5771,N_2387,N_3303);
nand U5772 (N_5772,N_2106,N_2056);
xnor U5773 (N_5773,N_2458,N_3865);
and U5774 (N_5774,N_3272,N_2633);
xor U5775 (N_5775,N_3241,N_2319);
nand U5776 (N_5776,N_3561,N_3411);
nand U5777 (N_5777,N_2528,N_3428);
or U5778 (N_5778,N_2388,N_3946);
nand U5779 (N_5779,N_2902,N_2978);
nand U5780 (N_5780,N_2804,N_3463);
nand U5781 (N_5781,N_3978,N_3159);
nor U5782 (N_5782,N_3992,N_3236);
or U5783 (N_5783,N_3591,N_2577);
and U5784 (N_5784,N_2067,N_2803);
and U5785 (N_5785,N_3626,N_2757);
xnor U5786 (N_5786,N_3000,N_3329);
or U5787 (N_5787,N_2506,N_3539);
or U5788 (N_5788,N_2589,N_3488);
or U5789 (N_5789,N_2137,N_3343);
nor U5790 (N_5790,N_2138,N_2779);
and U5791 (N_5791,N_3712,N_2121);
xor U5792 (N_5792,N_3901,N_3588);
nor U5793 (N_5793,N_3936,N_3925);
xor U5794 (N_5794,N_2972,N_3577);
nor U5795 (N_5795,N_2209,N_3350);
xnor U5796 (N_5796,N_3383,N_2611);
nor U5797 (N_5797,N_3346,N_2378);
nor U5798 (N_5798,N_2278,N_2198);
xor U5799 (N_5799,N_2683,N_3448);
or U5800 (N_5800,N_2506,N_3116);
or U5801 (N_5801,N_2351,N_3641);
or U5802 (N_5802,N_3728,N_3268);
xnor U5803 (N_5803,N_3822,N_2091);
or U5804 (N_5804,N_2152,N_3627);
nor U5805 (N_5805,N_2620,N_2074);
nor U5806 (N_5806,N_2441,N_2868);
nor U5807 (N_5807,N_2613,N_2797);
and U5808 (N_5808,N_2210,N_3831);
xnor U5809 (N_5809,N_2372,N_3815);
xnor U5810 (N_5810,N_2520,N_3909);
xor U5811 (N_5811,N_2765,N_3685);
xor U5812 (N_5812,N_2120,N_2139);
or U5813 (N_5813,N_3854,N_3680);
nand U5814 (N_5814,N_3783,N_2515);
and U5815 (N_5815,N_2843,N_2767);
and U5816 (N_5816,N_3608,N_3715);
xor U5817 (N_5817,N_3276,N_2458);
and U5818 (N_5818,N_3621,N_2142);
nand U5819 (N_5819,N_3524,N_3004);
or U5820 (N_5820,N_3048,N_3736);
xor U5821 (N_5821,N_2190,N_3584);
or U5822 (N_5822,N_3862,N_2275);
xor U5823 (N_5823,N_3103,N_3573);
or U5824 (N_5824,N_2112,N_3784);
nand U5825 (N_5825,N_3411,N_3545);
nor U5826 (N_5826,N_3354,N_2490);
or U5827 (N_5827,N_3492,N_3863);
xnor U5828 (N_5828,N_3982,N_2145);
nand U5829 (N_5829,N_3543,N_2364);
xnor U5830 (N_5830,N_3815,N_2415);
and U5831 (N_5831,N_3985,N_3527);
nor U5832 (N_5832,N_3868,N_3772);
or U5833 (N_5833,N_2502,N_2036);
nor U5834 (N_5834,N_3414,N_2656);
and U5835 (N_5835,N_3352,N_2114);
nand U5836 (N_5836,N_2788,N_2859);
nor U5837 (N_5837,N_3702,N_2423);
nor U5838 (N_5838,N_3977,N_2414);
and U5839 (N_5839,N_3774,N_3615);
xnor U5840 (N_5840,N_3371,N_2512);
nand U5841 (N_5841,N_2576,N_2788);
and U5842 (N_5842,N_2645,N_3673);
xnor U5843 (N_5843,N_2656,N_3606);
and U5844 (N_5844,N_3778,N_2114);
nand U5845 (N_5845,N_2298,N_2867);
nor U5846 (N_5846,N_3681,N_3978);
or U5847 (N_5847,N_2857,N_3797);
nor U5848 (N_5848,N_2166,N_3672);
xor U5849 (N_5849,N_2465,N_3863);
or U5850 (N_5850,N_3882,N_3530);
nor U5851 (N_5851,N_3594,N_2431);
nand U5852 (N_5852,N_2526,N_3222);
or U5853 (N_5853,N_2405,N_2288);
xnor U5854 (N_5854,N_3456,N_2634);
or U5855 (N_5855,N_3938,N_2218);
nand U5856 (N_5856,N_3232,N_2957);
xor U5857 (N_5857,N_2366,N_2179);
nand U5858 (N_5858,N_2678,N_2254);
xnor U5859 (N_5859,N_3986,N_2486);
or U5860 (N_5860,N_2265,N_2674);
and U5861 (N_5861,N_3057,N_2423);
nor U5862 (N_5862,N_2007,N_2672);
and U5863 (N_5863,N_2863,N_3570);
or U5864 (N_5864,N_3817,N_3333);
nor U5865 (N_5865,N_3161,N_3764);
and U5866 (N_5866,N_3775,N_2817);
nand U5867 (N_5867,N_2704,N_2371);
nor U5868 (N_5868,N_3987,N_2766);
or U5869 (N_5869,N_3531,N_3667);
nor U5870 (N_5870,N_3534,N_2981);
nor U5871 (N_5871,N_2806,N_2363);
or U5872 (N_5872,N_2700,N_3934);
nand U5873 (N_5873,N_3522,N_3758);
xor U5874 (N_5874,N_3410,N_3853);
nand U5875 (N_5875,N_2804,N_2953);
or U5876 (N_5876,N_2605,N_3943);
nand U5877 (N_5877,N_2100,N_3094);
xnor U5878 (N_5878,N_2245,N_2822);
or U5879 (N_5879,N_3443,N_3869);
xor U5880 (N_5880,N_3688,N_2932);
xnor U5881 (N_5881,N_2269,N_2028);
nand U5882 (N_5882,N_2989,N_3656);
nor U5883 (N_5883,N_2605,N_2135);
nor U5884 (N_5884,N_2178,N_3864);
xor U5885 (N_5885,N_3644,N_3867);
nor U5886 (N_5886,N_2643,N_2121);
nand U5887 (N_5887,N_2591,N_3807);
or U5888 (N_5888,N_3550,N_3213);
and U5889 (N_5889,N_3051,N_3548);
or U5890 (N_5890,N_2104,N_3106);
xor U5891 (N_5891,N_3517,N_3629);
nand U5892 (N_5892,N_3299,N_2181);
or U5893 (N_5893,N_2800,N_2514);
and U5894 (N_5894,N_2384,N_3497);
and U5895 (N_5895,N_2432,N_3115);
xor U5896 (N_5896,N_3966,N_3691);
xor U5897 (N_5897,N_3490,N_2651);
or U5898 (N_5898,N_3203,N_3408);
nor U5899 (N_5899,N_3619,N_2132);
nand U5900 (N_5900,N_3382,N_3774);
nor U5901 (N_5901,N_2333,N_2772);
and U5902 (N_5902,N_2681,N_3663);
nand U5903 (N_5903,N_2064,N_2747);
or U5904 (N_5904,N_3298,N_2046);
nand U5905 (N_5905,N_2109,N_2849);
or U5906 (N_5906,N_3619,N_2764);
and U5907 (N_5907,N_3983,N_2502);
or U5908 (N_5908,N_2394,N_3599);
nand U5909 (N_5909,N_3862,N_3111);
and U5910 (N_5910,N_2035,N_2584);
nor U5911 (N_5911,N_3700,N_3086);
nand U5912 (N_5912,N_3274,N_3071);
nor U5913 (N_5913,N_2912,N_3726);
xnor U5914 (N_5914,N_2051,N_2373);
xnor U5915 (N_5915,N_2059,N_2186);
nor U5916 (N_5916,N_2657,N_3991);
and U5917 (N_5917,N_3939,N_3259);
nand U5918 (N_5918,N_3761,N_3095);
and U5919 (N_5919,N_3853,N_2175);
or U5920 (N_5920,N_3688,N_2028);
and U5921 (N_5921,N_2649,N_3190);
nor U5922 (N_5922,N_3660,N_2677);
nand U5923 (N_5923,N_2347,N_2165);
nand U5924 (N_5924,N_3703,N_3284);
and U5925 (N_5925,N_3563,N_2035);
nand U5926 (N_5926,N_2132,N_2779);
nand U5927 (N_5927,N_3614,N_2610);
nand U5928 (N_5928,N_2772,N_2015);
and U5929 (N_5929,N_2448,N_3992);
xnor U5930 (N_5930,N_2231,N_2624);
nand U5931 (N_5931,N_2363,N_2805);
nand U5932 (N_5932,N_2096,N_3886);
xor U5933 (N_5933,N_2407,N_3325);
or U5934 (N_5934,N_3586,N_3468);
and U5935 (N_5935,N_3023,N_3815);
xor U5936 (N_5936,N_3877,N_2919);
xor U5937 (N_5937,N_2857,N_2110);
or U5938 (N_5938,N_2175,N_3820);
nor U5939 (N_5939,N_2103,N_3539);
xor U5940 (N_5940,N_2024,N_2864);
nor U5941 (N_5941,N_3197,N_3688);
xor U5942 (N_5942,N_2070,N_3090);
or U5943 (N_5943,N_3500,N_2720);
nor U5944 (N_5944,N_3104,N_3248);
or U5945 (N_5945,N_3404,N_2652);
or U5946 (N_5946,N_2909,N_3864);
nand U5947 (N_5947,N_3805,N_3468);
nor U5948 (N_5948,N_2076,N_3740);
nand U5949 (N_5949,N_2328,N_3539);
xor U5950 (N_5950,N_3811,N_3308);
or U5951 (N_5951,N_2652,N_3857);
xor U5952 (N_5952,N_2911,N_2828);
nor U5953 (N_5953,N_3511,N_2114);
nor U5954 (N_5954,N_2267,N_3086);
and U5955 (N_5955,N_2069,N_3559);
nor U5956 (N_5956,N_2166,N_3063);
nand U5957 (N_5957,N_3535,N_3065);
nand U5958 (N_5958,N_3111,N_3205);
xor U5959 (N_5959,N_3875,N_2697);
nor U5960 (N_5960,N_2543,N_3781);
nor U5961 (N_5961,N_2997,N_3545);
nor U5962 (N_5962,N_2383,N_3793);
nand U5963 (N_5963,N_2890,N_2999);
nor U5964 (N_5964,N_2298,N_3162);
nand U5965 (N_5965,N_3731,N_2070);
or U5966 (N_5966,N_2418,N_2472);
and U5967 (N_5967,N_2983,N_2796);
and U5968 (N_5968,N_3693,N_2565);
and U5969 (N_5969,N_3982,N_2313);
and U5970 (N_5970,N_3725,N_3262);
or U5971 (N_5971,N_3054,N_3012);
or U5972 (N_5972,N_2021,N_3664);
or U5973 (N_5973,N_3081,N_2177);
and U5974 (N_5974,N_3620,N_3430);
nor U5975 (N_5975,N_3043,N_3780);
nor U5976 (N_5976,N_3075,N_3576);
xnor U5977 (N_5977,N_2844,N_2791);
or U5978 (N_5978,N_3589,N_3461);
or U5979 (N_5979,N_3010,N_2439);
and U5980 (N_5980,N_2552,N_2673);
and U5981 (N_5981,N_2828,N_2026);
and U5982 (N_5982,N_2198,N_2251);
nor U5983 (N_5983,N_3205,N_3667);
nor U5984 (N_5984,N_2958,N_3435);
and U5985 (N_5985,N_3953,N_3171);
nand U5986 (N_5986,N_3660,N_3581);
nand U5987 (N_5987,N_3360,N_2920);
nor U5988 (N_5988,N_3849,N_2668);
nand U5989 (N_5989,N_2447,N_2110);
nor U5990 (N_5990,N_3145,N_2735);
or U5991 (N_5991,N_3972,N_2651);
nand U5992 (N_5992,N_2840,N_3143);
nand U5993 (N_5993,N_3874,N_3868);
or U5994 (N_5994,N_3180,N_3163);
and U5995 (N_5995,N_2235,N_3535);
nand U5996 (N_5996,N_2553,N_2562);
or U5997 (N_5997,N_3232,N_2679);
nor U5998 (N_5998,N_3595,N_3560);
nor U5999 (N_5999,N_2361,N_3373);
or U6000 (N_6000,N_5808,N_5124);
and U6001 (N_6001,N_4217,N_4604);
xor U6002 (N_6002,N_4314,N_5919);
xnor U6003 (N_6003,N_5186,N_4657);
nor U6004 (N_6004,N_4570,N_5282);
or U6005 (N_6005,N_5982,N_4070);
nand U6006 (N_6006,N_4369,N_5498);
nand U6007 (N_6007,N_5351,N_4636);
or U6008 (N_6008,N_5834,N_4237);
nor U6009 (N_6009,N_4871,N_4844);
nor U6010 (N_6010,N_4412,N_5813);
xnor U6011 (N_6011,N_5173,N_4565);
and U6012 (N_6012,N_5913,N_4769);
xor U6013 (N_6013,N_4340,N_4530);
or U6014 (N_6014,N_4977,N_5715);
xor U6015 (N_6015,N_4170,N_4263);
or U6016 (N_6016,N_5859,N_4888);
nor U6017 (N_6017,N_4042,N_5030);
nand U6018 (N_6018,N_5306,N_4824);
nand U6019 (N_6019,N_4509,N_4782);
nor U6020 (N_6020,N_5489,N_5104);
nand U6021 (N_6021,N_5316,N_4551);
and U6022 (N_6022,N_5285,N_5950);
xor U6023 (N_6023,N_5318,N_4862);
xor U6024 (N_6024,N_4525,N_5093);
nand U6025 (N_6025,N_4016,N_4833);
xor U6026 (N_6026,N_5178,N_4726);
and U6027 (N_6027,N_5545,N_5763);
xnor U6028 (N_6028,N_4869,N_4175);
or U6029 (N_6029,N_4994,N_5661);
nand U6030 (N_6030,N_5339,N_5414);
and U6031 (N_6031,N_4278,N_5435);
or U6032 (N_6032,N_4457,N_4533);
xnor U6033 (N_6033,N_4678,N_5029);
and U6034 (N_6034,N_5739,N_5769);
xor U6035 (N_6035,N_5755,N_5829);
and U6036 (N_6036,N_5170,N_5389);
xor U6037 (N_6037,N_4705,N_5821);
or U6038 (N_6038,N_4702,N_4499);
nor U6039 (N_6039,N_4558,N_5594);
and U6040 (N_6040,N_5119,N_4223);
xnor U6041 (N_6041,N_5263,N_4183);
nand U6042 (N_6042,N_5552,N_4789);
and U6043 (N_6043,N_4588,N_4357);
or U6044 (N_6044,N_5957,N_5796);
nand U6045 (N_6045,N_5201,N_5777);
nor U6046 (N_6046,N_4015,N_5698);
nor U6047 (N_6047,N_4718,N_4885);
and U6048 (N_6048,N_5038,N_4786);
and U6049 (N_6049,N_4767,N_5441);
and U6050 (N_6050,N_5592,N_4451);
nand U6051 (N_6051,N_5925,N_5127);
xor U6052 (N_6052,N_4686,N_4436);
or U6053 (N_6053,N_5775,N_4270);
nand U6054 (N_6054,N_4148,N_4923);
or U6055 (N_6055,N_5889,N_4783);
or U6056 (N_6056,N_5874,N_5546);
or U6057 (N_6057,N_4609,N_4747);
or U6058 (N_6058,N_4054,N_4995);
nand U6059 (N_6059,N_5637,N_4130);
or U6060 (N_6060,N_4372,N_5907);
or U6061 (N_6061,N_5336,N_5184);
xnor U6062 (N_6062,N_5118,N_5229);
or U6063 (N_6063,N_5804,N_5419);
xnor U6064 (N_6064,N_4129,N_5144);
xnor U6065 (N_6065,N_5921,N_4075);
xnor U6066 (N_6066,N_4399,N_5892);
or U6067 (N_6067,N_4681,N_4303);
nand U6068 (N_6068,N_5011,N_4300);
nor U6069 (N_6069,N_4689,N_4271);
nand U6070 (N_6070,N_4301,N_5877);
xor U6071 (N_6071,N_4157,N_5936);
nand U6072 (N_6072,N_5729,N_4150);
xor U6073 (N_6073,N_4614,N_5035);
nand U6074 (N_6074,N_5010,N_5811);
nor U6075 (N_6075,N_4543,N_5831);
or U6076 (N_6076,N_5559,N_4750);
or U6077 (N_6077,N_4238,N_4382);
and U6078 (N_6078,N_5644,N_5748);
or U6079 (N_6079,N_5279,N_4302);
nor U6080 (N_6080,N_5329,N_5294);
nor U6081 (N_6081,N_5424,N_5046);
or U6082 (N_6082,N_5601,N_5057);
xnor U6083 (N_6083,N_4002,N_5126);
or U6084 (N_6084,N_4163,N_5550);
or U6085 (N_6085,N_5939,N_5745);
or U6086 (N_6086,N_4470,N_5612);
nor U6087 (N_6087,N_4804,N_4084);
and U6088 (N_6088,N_5416,N_5793);
and U6089 (N_6089,N_4095,N_5569);
nand U6090 (N_6090,N_4280,N_5311);
and U6091 (N_6091,N_5253,N_4641);
or U6092 (N_6092,N_5970,N_4594);
xnor U6093 (N_6093,N_4260,N_5410);
or U6094 (N_6094,N_4608,N_4582);
and U6095 (N_6095,N_4932,N_5437);
xor U6096 (N_6096,N_4692,N_5133);
nand U6097 (N_6097,N_4370,N_4097);
nor U6098 (N_6098,N_5252,N_4896);
xor U6099 (N_6099,N_4899,N_5945);
and U6100 (N_6100,N_5677,N_5560);
or U6101 (N_6101,N_5417,N_5947);
nand U6102 (N_6102,N_5474,N_4355);
xor U6103 (N_6103,N_5959,N_5666);
nand U6104 (N_6104,N_5482,N_4045);
or U6105 (N_6105,N_4631,N_4842);
xnor U6106 (N_6106,N_4714,N_4787);
nand U6107 (N_6107,N_5112,N_4125);
nand U6108 (N_6108,N_5367,N_4388);
nand U6109 (N_6109,N_5841,N_4200);
nand U6110 (N_6110,N_5985,N_5971);
and U6111 (N_6111,N_4746,N_5228);
and U6112 (N_6112,N_4922,N_4014);
and U6113 (N_6113,N_4483,N_4063);
nand U6114 (N_6114,N_4093,N_5565);
xor U6115 (N_6115,N_5708,N_5894);
nand U6116 (N_6116,N_4625,N_5526);
nor U6117 (N_6117,N_4597,N_4521);
and U6118 (N_6118,N_5366,N_4502);
and U6119 (N_6119,N_5703,N_4341);
nand U6120 (N_6120,N_5111,N_4766);
or U6121 (N_6121,N_5182,N_5962);
and U6122 (N_6122,N_5785,N_4098);
xnor U6123 (N_6123,N_4752,N_5451);
nand U6124 (N_6124,N_5700,N_4018);
and U6125 (N_6125,N_5483,N_4936);
nand U6126 (N_6126,N_5710,N_5393);
or U6127 (N_6127,N_5851,N_5617);
or U6128 (N_6128,N_4071,N_5726);
nand U6129 (N_6129,N_5452,N_5232);
or U6130 (N_6130,N_4591,N_5523);
or U6131 (N_6131,N_5534,N_4792);
nand U6132 (N_6132,N_4668,N_4822);
nor U6133 (N_6133,N_5890,N_4527);
xnor U6134 (N_6134,N_5683,N_4571);
and U6135 (N_6135,N_4791,N_5392);
nand U6136 (N_6136,N_5308,N_5885);
xor U6137 (N_6137,N_4665,N_5325);
or U6138 (N_6138,N_4161,N_4317);
nor U6139 (N_6139,N_5760,N_4479);
or U6140 (N_6140,N_5586,N_4354);
xor U6141 (N_6141,N_5384,N_5028);
nand U6142 (N_6142,N_5778,N_4351);
and U6143 (N_6143,N_4957,N_5281);
or U6144 (N_6144,N_4267,N_5718);
xnor U6145 (N_6145,N_5349,N_4032);
xor U6146 (N_6146,N_5828,N_4306);
and U6147 (N_6147,N_4515,N_4443);
or U6148 (N_6148,N_5518,N_4363);
nor U6149 (N_6149,N_4112,N_4915);
nor U6150 (N_6150,N_4773,N_5738);
or U6151 (N_6151,N_5379,N_4383);
and U6152 (N_6152,N_4549,N_5801);
and U6153 (N_6153,N_4394,N_4508);
and U6154 (N_6154,N_5799,N_4975);
nand U6155 (N_6155,N_4319,N_4398);
or U6156 (N_6156,N_4850,N_4122);
and U6157 (N_6157,N_5599,N_4893);
nor U6158 (N_6158,N_4648,N_5634);
nor U6159 (N_6159,N_5802,N_4947);
and U6160 (N_6160,N_5337,N_5116);
xnor U6161 (N_6161,N_4607,N_5762);
nand U6162 (N_6162,N_5260,N_4816);
and U6163 (N_6163,N_5303,N_5444);
and U6164 (N_6164,N_4827,N_5163);
nand U6165 (N_6165,N_4968,N_5205);
nor U6166 (N_6166,N_4198,N_4143);
xnor U6167 (N_6167,N_5678,N_5623);
xnor U6168 (N_6168,N_4496,N_5058);
nand U6169 (N_6169,N_5830,N_5782);
and U6170 (N_6170,N_5231,N_5625);
and U6171 (N_6171,N_4246,N_5912);
xnor U6172 (N_6172,N_5465,N_5973);
nor U6173 (N_6173,N_5324,N_4679);
or U6174 (N_6174,N_5940,N_5624);
nand U6175 (N_6175,N_4992,N_4349);
and U6176 (N_6176,N_5963,N_4040);
or U6177 (N_6177,N_4485,N_5314);
nor U6178 (N_6178,N_5015,N_4442);
xor U6179 (N_6179,N_5531,N_5621);
and U6180 (N_6180,N_5242,N_4945);
nor U6181 (N_6181,N_5404,N_5990);
and U6182 (N_6182,N_5927,N_4249);
or U6183 (N_6183,N_5024,N_5409);
nand U6184 (N_6184,N_4482,N_4779);
or U6185 (N_6185,N_4660,N_4327);
or U6186 (N_6186,N_4078,N_5979);
nor U6187 (N_6187,N_4808,N_4494);
nand U6188 (N_6188,N_4102,N_5132);
or U6189 (N_6189,N_5286,N_5542);
or U6190 (N_6190,N_5911,N_4149);
xnor U6191 (N_6191,N_5338,N_4545);
xnor U6192 (N_6192,N_4963,N_5595);
nand U6193 (N_6193,N_5582,N_5295);
nor U6194 (N_6194,N_5887,N_5169);
nor U6195 (N_6195,N_5615,N_5411);
or U6196 (N_6196,N_5918,N_4446);
or U6197 (N_6197,N_4073,N_5673);
and U6198 (N_6198,N_5044,N_5312);
and U6199 (N_6199,N_5086,N_5245);
xor U6200 (N_6200,N_5378,N_4555);
xor U6201 (N_6201,N_4661,N_5524);
xnor U6202 (N_6202,N_5917,N_5276);
and U6203 (N_6203,N_5564,N_4461);
xnor U6204 (N_6204,N_4642,N_5690);
or U6205 (N_6205,N_5865,N_4882);
nor U6206 (N_6206,N_4420,N_4350);
or U6207 (N_6207,N_5539,N_4931);
or U6208 (N_6208,N_5064,N_4598);
nand U6209 (N_6209,N_5102,N_4364);
nand U6210 (N_6210,N_5167,N_4536);
and U6211 (N_6211,N_5916,N_4449);
nor U6212 (N_6212,N_4511,N_5199);
nand U6213 (N_6213,N_4389,N_4134);
nor U6214 (N_6214,N_4501,N_4210);
or U6215 (N_6215,N_5188,N_5089);
xnor U6216 (N_6216,N_5861,N_5737);
nand U6217 (N_6217,N_5291,N_5369);
nand U6218 (N_6218,N_5398,N_5391);
nor U6219 (N_6219,N_5105,N_5580);
and U6220 (N_6220,N_5005,N_5888);
and U6221 (N_6221,N_4761,N_4219);
and U6222 (N_6222,N_4135,N_5353);
xnor U6223 (N_6223,N_4857,N_4245);
nand U6224 (N_6224,N_5774,N_5767);
and U6225 (N_6225,N_5331,N_4362);
xnor U6226 (N_6226,N_5494,N_5639);
nand U6227 (N_6227,N_4654,N_4425);
and U6228 (N_6228,N_5998,N_5108);
nand U6229 (N_6229,N_5259,N_4074);
or U6230 (N_6230,N_5743,N_5689);
and U6231 (N_6231,N_5098,N_4731);
nand U6232 (N_6232,N_5072,N_4847);
or U6233 (N_6233,N_4182,N_4561);
xor U6234 (N_6234,N_4704,N_4358);
xnor U6235 (N_6235,N_5541,N_5195);
and U6236 (N_6236,N_4321,N_4538);
and U6237 (N_6237,N_5557,N_4682);
and U6238 (N_6238,N_5868,N_5941);
or U6239 (N_6239,N_5380,N_4113);
and U6240 (N_6240,N_4248,N_5997);
nand U6241 (N_6241,N_5744,N_5701);
or U6242 (N_6242,N_4926,N_4178);
nor U6243 (N_6243,N_5114,N_5341);
nand U6244 (N_6244,N_4622,N_4541);
xnor U6245 (N_6245,N_5226,N_4004);
and U6246 (N_6246,N_5532,N_5528);
nand U6247 (N_6247,N_4826,N_5313);
nand U6248 (N_6248,N_4464,N_4956);
and U6249 (N_6249,N_5321,N_4395);
and U6250 (N_6250,N_5334,N_5002);
and U6251 (N_6251,N_4585,N_5930);
nor U6252 (N_6252,N_5400,N_4900);
nand U6253 (N_6253,N_4030,N_5138);
nand U6254 (N_6254,N_5519,N_5884);
nor U6255 (N_6255,N_4308,N_4233);
nand U6256 (N_6256,N_4077,N_5079);
or U6257 (N_6257,N_5672,N_5855);
xor U6258 (N_6258,N_4619,N_5648);
nand U6259 (N_6259,N_4873,N_4277);
xnor U6260 (N_6260,N_5611,N_5593);
nor U6261 (N_6261,N_5045,N_4834);
xor U6262 (N_6262,N_4244,N_5068);
nand U6263 (N_6263,N_4104,N_4522);
and U6264 (N_6264,N_5953,N_5328);
or U6265 (N_6265,N_5641,N_4083);
xor U6266 (N_6266,N_5920,N_5439);
nand U6267 (N_6267,N_4935,N_5469);
and U6268 (N_6268,N_5996,N_4279);
nor U6269 (N_6269,N_5879,N_4514);
and U6270 (N_6270,N_5340,N_4160);
nor U6271 (N_6271,N_5506,N_5515);
nor U6272 (N_6272,N_5923,N_4552);
xor U6273 (N_6273,N_5244,N_5694);
or U6274 (N_6274,N_4544,N_4427);
nor U6275 (N_6275,N_4473,N_4049);
and U6276 (N_6276,N_4402,N_5840);
xor U6277 (N_6277,N_4870,N_4265);
or U6278 (N_6278,N_4700,N_5576);
and U6279 (N_6279,N_5610,N_4730);
nor U6280 (N_6280,N_4950,N_4039);
nor U6281 (N_6281,N_5399,N_4159);
or U6282 (N_6282,N_5589,N_5946);
nand U6283 (N_6283,N_4703,N_4236);
nand U6284 (N_6284,N_4880,N_5951);
and U6285 (N_6285,N_4720,N_4116);
nand U6286 (N_6286,N_5268,N_5810);
nand U6287 (N_6287,N_5000,N_5141);
nor U6288 (N_6288,N_5765,N_4667);
and U6289 (N_6289,N_4964,N_5679);
and U6290 (N_6290,N_5631,N_4339);
or U6291 (N_6291,N_5023,N_4563);
or U6292 (N_6292,N_4003,N_4685);
nand U6293 (N_6293,N_5850,N_5575);
nand U6294 (N_6294,N_4972,N_4484);
and U6295 (N_6295,N_5952,N_5712);
or U6296 (N_6296,N_4179,N_5236);
xnor U6297 (N_6297,N_5554,N_4795);
nand U6298 (N_6298,N_5503,N_4337);
nor U6299 (N_6299,N_5302,N_4624);
xnor U6300 (N_6300,N_5164,N_4912);
nor U6301 (N_6301,N_4874,N_4902);
or U6302 (N_6302,N_4123,N_4456);
nand U6303 (N_6303,N_4020,N_4709);
xnor U6304 (N_6304,N_4408,N_4907);
xnor U6305 (N_6305,N_4776,N_4669);
nand U6306 (N_6306,N_5442,N_4780);
xnor U6307 (N_6307,N_5113,N_4264);
and U6308 (N_6308,N_5548,N_5878);
nand U6309 (N_6309,N_5817,N_4512);
nand U6310 (N_6310,N_5106,N_5402);
nor U6311 (N_6311,N_4276,N_4373);
or U6312 (N_6312,N_5896,N_4173);
nor U6313 (N_6313,N_4414,N_5757);
nand U6314 (N_6314,N_5643,N_4519);
xnor U6315 (N_6315,N_4539,N_4961);
nor U6316 (N_6316,N_5436,N_5561);
and U6317 (N_6317,N_4518,N_4940);
and U6318 (N_6318,N_5794,N_4955);
or U6319 (N_6319,N_5513,N_4055);
nor U6320 (N_6320,N_5750,N_5270);
or U6321 (N_6321,N_5265,N_5434);
nor U6322 (N_6322,N_4859,N_4124);
xor U6323 (N_6323,N_4906,N_5382);
or U6324 (N_6324,N_4232,N_4013);
nand U6325 (N_6325,N_4171,N_5152);
xor U6326 (N_6326,N_5275,N_4380);
or U6327 (N_6327,N_4733,N_4960);
xor U6328 (N_6328,N_4696,N_5994);
and U6329 (N_6329,N_5961,N_4497);
nor U6330 (N_6330,N_5070,N_4294);
or U6331 (N_6331,N_5273,N_5826);
nand U6332 (N_6332,N_5455,N_5875);
nand U6333 (N_6333,N_4487,N_5842);
or U6334 (N_6334,N_4811,N_5177);
xnor U6335 (N_6335,N_5640,N_4021);
xnor U6336 (N_6336,N_5496,N_5633);
xor U6337 (N_6337,N_5572,N_4784);
nand U6338 (N_6338,N_4603,N_5264);
or U6339 (N_6339,N_5838,N_5972);
xor U6340 (N_6340,N_5373,N_4417);
nor U6341 (N_6341,N_4193,N_5854);
nand U6342 (N_6342,N_4556,N_4634);
and U6343 (N_6343,N_5636,N_5759);
or U6344 (N_6344,N_5447,N_5902);
nor U6345 (N_6345,N_4195,N_5733);
nand U6346 (N_6346,N_4728,N_5719);
xor U6347 (N_6347,N_4980,N_4109);
xnor U6348 (N_6348,N_5180,N_4845);
and U6349 (N_6349,N_4821,N_5508);
or U6350 (N_6350,N_4984,N_4225);
or U6351 (N_6351,N_4916,N_4127);
nand U6352 (N_6352,N_4662,N_5059);
xnor U6353 (N_6353,N_5520,N_5571);
or U6354 (N_6354,N_4837,N_5357);
nor U6355 (N_6355,N_5695,N_5618);
nor U6356 (N_6356,N_4537,N_4930);
nor U6357 (N_6357,N_5556,N_4520);
and U6358 (N_6358,N_4928,N_4204);
xnor U6359 (N_6359,N_4510,N_4656);
and U6360 (N_6360,N_4586,N_4831);
nor U6361 (N_6361,N_4296,N_4640);
and U6362 (N_6362,N_4941,N_5342);
and U6363 (N_6363,N_4925,N_4031);
nor U6364 (N_6364,N_4997,N_4413);
nand U6365 (N_6365,N_5898,N_5464);
or U6366 (N_6366,N_5039,N_4567);
and U6367 (N_6367,N_4650,N_4951);
and U6368 (N_6368,N_4197,N_4216);
or U6369 (N_6369,N_5819,N_4424);
and U6370 (N_6370,N_4701,N_5869);
and U6371 (N_6371,N_4818,N_5960);
xnor U6372 (N_6372,N_4905,N_5129);
nand U6373 (N_6373,N_5606,N_5065);
nor U6374 (N_6374,N_4895,N_5751);
and U6375 (N_6375,N_4973,N_4151);
nand U6376 (N_6376,N_5758,N_4111);
xnor U6377 (N_6377,N_5613,N_5022);
nand U6378 (N_6378,N_5607,N_5975);
and U6379 (N_6379,N_5596,N_5728);
and U6380 (N_6380,N_5547,N_4970);
xnor U6381 (N_6381,N_5510,N_5299);
xor U6382 (N_6382,N_5196,N_4981);
and U6383 (N_6383,N_4441,N_5860);
nand U6384 (N_6384,N_4814,N_5446);
nor U6385 (N_6385,N_4005,N_5134);
nand U6386 (N_6386,N_4154,N_4990);
nor U6387 (N_6387,N_4332,N_4763);
xnor U6388 (N_6388,N_4307,N_5208);
nor U6389 (N_6389,N_5401,N_4674);
nand U6390 (N_6390,N_4033,N_4630);
and U6391 (N_6391,N_5307,N_4865);
or U6392 (N_6392,N_4867,N_5063);
and U6393 (N_6393,N_5335,N_4914);
nor U6394 (N_6394,N_4486,N_4954);
and U6395 (N_6395,N_5272,N_4029);
xor U6396 (N_6396,N_4344,N_5194);
and U6397 (N_6397,N_4664,N_4465);
nand U6398 (N_6398,N_5092,N_4145);
nor U6399 (N_6399,N_5988,N_4391);
or U6400 (N_6400,N_5290,N_4721);
nor U6401 (N_6401,N_5047,N_5344);
or U6402 (N_6402,N_4106,N_4100);
and U6403 (N_6403,N_4053,N_5723);
or U6404 (N_6404,N_4708,N_5585);
nand U6405 (N_6405,N_4397,N_5326);
xnor U6406 (N_6406,N_5361,N_4059);
or U6407 (N_6407,N_4167,N_5449);
xnor U6408 (N_6408,N_5013,N_5900);
and U6409 (N_6409,N_5862,N_5317);
or U6410 (N_6410,N_5783,N_5734);
or U6411 (N_6411,N_4258,N_4891);
nand U6412 (N_6412,N_4243,N_5122);
nor U6413 (N_6413,N_4739,N_4794);
nor U6414 (N_6414,N_4697,N_5833);
nor U6415 (N_6415,N_4754,N_5363);
and U6416 (N_6416,N_5460,N_4305);
or U6417 (N_6417,N_5761,N_5543);
nand U6418 (N_6418,N_5685,N_5090);
or U6419 (N_6419,N_5856,N_4387);
and U6420 (N_6420,N_5910,N_4347);
xnor U6421 (N_6421,N_5074,N_4724);
and U6422 (N_6422,N_4601,N_5095);
and U6423 (N_6423,N_5396,N_4866);
nand U6424 (N_6424,N_5073,N_4459);
nand U6425 (N_6425,N_4812,N_5346);
and U6426 (N_6426,N_4432,N_5130);
nand U6427 (N_6427,N_5080,N_4320);
or U6428 (N_6428,N_5635,N_4400);
and U6429 (N_6429,N_5699,N_4220);
or U6430 (N_6430,N_5590,N_5773);
xnor U6431 (N_6431,N_4626,N_5021);
nand U6432 (N_6432,N_5491,N_5372);
nor U6433 (N_6433,N_4165,N_5006);
xnor U6434 (N_6434,N_5210,N_5248);
nor U6435 (N_6435,N_5217,N_5732);
xnor U6436 (N_6436,N_4796,N_5591);
xnor U6437 (N_6437,N_5521,N_4287);
and U6438 (N_6438,N_5725,N_5288);
or U6439 (N_6439,N_5562,N_5720);
and U6440 (N_6440,N_4403,N_4513);
xor U6441 (N_6441,N_4137,N_5240);
and U6442 (N_6442,N_5222,N_5922);
nand U6443 (N_6443,N_4735,N_5175);
nand U6444 (N_6444,N_4168,N_5603);
xor U6445 (N_6445,N_4406,N_4547);
nand U6446 (N_6446,N_4892,N_4490);
or U6447 (N_6447,N_5212,N_4330);
or U6448 (N_6448,N_4807,N_5207);
xnor U6449 (N_6449,N_4851,N_4581);
nand U6450 (N_6450,N_5225,N_5823);
nor U6451 (N_6451,N_5292,N_5667);
xor U6452 (N_6452,N_5747,N_5333);
xor U6453 (N_6453,N_4336,N_4334);
nand U6454 (N_6454,N_5420,N_4114);
nor U6455 (N_6455,N_5781,N_5976);
xor U6456 (N_6456,N_5214,N_4138);
nand U6457 (N_6457,N_5347,N_5405);
and U6458 (N_6458,N_5844,N_5517);
xor U6459 (N_6459,N_5269,N_4829);
xor U6460 (N_6460,N_5493,N_5016);
and U6461 (N_6461,N_5697,N_4901);
or U6462 (N_6462,N_5076,N_5421);
nor U6463 (N_6463,N_5779,N_4452);
nand U6464 (N_6464,N_4176,N_5609);
xnor U6465 (N_6465,N_5485,N_4255);
and U6466 (N_6466,N_5348,N_4006);
or U6467 (N_6467,N_5753,N_4026);
xor U6468 (N_6468,N_5664,N_5852);
nor U6469 (N_6469,N_5407,N_4838);
or U6470 (N_6470,N_4346,N_5165);
nor U6471 (N_6471,N_4352,N_5502);
nor U6472 (N_6472,N_4595,N_5966);
xnor U6473 (N_6473,N_5239,N_4835);
nor U6474 (N_6474,N_5247,N_5262);
nand U6475 (N_6475,N_4745,N_5221);
nand U6476 (N_6476,N_5408,N_4328);
xnor U6477 (N_6477,N_5220,N_5368);
nor U6478 (N_6478,N_5149,N_4396);
nand U6479 (N_6479,N_5671,N_5929);
and U6480 (N_6480,N_5730,N_4934);
xor U6481 (N_6481,N_4861,N_5107);
or U6482 (N_6482,N_5406,N_4559);
xor U6483 (N_6483,N_4201,N_4082);
xnor U6484 (N_6484,N_5551,N_5993);
nor U6485 (N_6485,N_4331,N_5278);
xnor U6486 (N_6486,N_4315,N_5305);
and U6487 (N_6487,N_4800,N_4036);
and U6488 (N_6488,N_4503,N_5620);
nand U6489 (N_6489,N_5218,N_4599);
or U6490 (N_6490,N_5563,N_5103);
nand U6491 (N_6491,N_5786,N_5237);
and U6492 (N_6492,N_5824,N_5162);
xnor U6493 (N_6493,N_4756,N_5764);
nand U6494 (N_6494,N_4325,N_4326);
nand U6495 (N_6495,N_5274,N_4506);
xnor U6496 (N_6496,N_4172,N_4854);
nand U6497 (N_6497,N_5853,N_4072);
or U6498 (N_6498,N_5287,N_4991);
nor U6499 (N_6499,N_4186,N_5145);
or U6500 (N_6500,N_5504,N_4633);
and U6501 (N_6501,N_4230,N_5462);
nor U6502 (N_6502,N_5883,N_5235);
xnor U6503 (N_6503,N_5445,N_4310);
xor U6504 (N_6504,N_5155,N_5684);
or U6505 (N_6505,N_4192,N_5688);
and U6506 (N_6506,N_4738,N_5181);
xnor U6507 (N_6507,N_4471,N_5991);
xor U6508 (N_6508,N_5135,N_4612);
and U6509 (N_6509,N_5096,N_4028);
nor U6510 (N_6510,N_4256,N_5418);
nor U6511 (N_6511,N_4575,N_4024);
nor U6512 (N_6512,N_5301,N_5500);
nand U6513 (N_6513,N_4933,N_4080);
or U6514 (N_6514,N_5867,N_4286);
or U6515 (N_6515,N_4448,N_4121);
nand U6516 (N_6516,N_4898,N_4052);
xor U6517 (N_6517,N_4239,N_4290);
xor U6518 (N_6518,N_4261,N_4146);
nor U6519 (N_6519,N_4468,N_4962);
nand U6520 (N_6520,N_4392,N_4535);
nand U6521 (N_6521,N_5495,N_5481);
nand U6522 (N_6522,N_4534,N_5663);
and U6523 (N_6523,N_5626,N_5646);
or U6524 (N_6524,N_4952,N_4732);
xnor U6525 (N_6525,N_5784,N_4741);
and U6526 (N_6526,N_4578,N_4488);
nand U6527 (N_6527,N_5954,N_5529);
nor U6528 (N_6528,N_4229,N_4115);
nor U6529 (N_6529,N_4643,N_5937);
nand U6530 (N_6530,N_5488,N_4085);
nand U6531 (N_6531,N_4241,N_5300);
nand U6532 (N_6532,N_4979,N_4676);
or U6533 (N_6533,N_5780,N_4989);
and U6534 (N_6534,N_4615,N_4855);
nor U6535 (N_6535,N_4680,N_5835);
xnor U6536 (N_6536,N_5429,N_4670);
nand U6537 (N_6537,N_4046,N_5189);
xnor U6538 (N_6538,N_4592,N_4550);
nor U6539 (N_6539,N_5309,N_5223);
nand U6540 (N_6540,N_4825,N_5527);
and U6541 (N_6541,N_5956,N_5789);
nor U6542 (N_6542,N_5109,N_4740);
nor U6543 (N_6543,N_5176,N_4986);
or U6544 (N_6544,N_5412,N_4785);
and U6545 (N_6545,N_5383,N_4546);
xnor U6546 (N_6546,N_4252,N_4517);
and U6547 (N_6547,N_4273,N_5499);
nand U6548 (N_6548,N_4772,N_5048);
or U6549 (N_6549,N_4155,N_5430);
xnor U6550 (N_6550,N_5662,N_4119);
and U6551 (N_6551,N_5901,N_4128);
xor U6552 (N_6552,N_4268,N_4472);
and U6553 (N_6553,N_4706,N_4462);
or U6554 (N_6554,N_5203,N_4913);
and U6555 (N_6555,N_5581,N_4655);
and U6556 (N_6556,N_4433,N_4879);
and U6557 (N_6557,N_5075,N_5974);
xor U6558 (N_6558,N_4421,N_4429);
xnor U6559 (N_6559,N_5472,N_5087);
and U6560 (N_6560,N_5509,N_4034);
and U6561 (N_6561,N_5914,N_5549);
and U6562 (N_6562,N_4272,N_4969);
nor U6563 (N_6563,N_4639,N_5525);
and U6564 (N_6564,N_5280,N_5036);
xnor U6565 (N_6565,N_5915,N_5986);
nor U6566 (N_6566,N_5656,N_4316);
xnor U6567 (N_6567,N_5933,N_5822);
nor U6568 (N_6568,N_5094,N_4228);
and U6569 (N_6569,N_5752,N_4993);
or U6570 (N_6570,N_4491,N_4426);
and U6571 (N_6571,N_4374,N_5007);
xnor U6572 (N_6572,N_5866,N_4649);
nor U6573 (N_6573,N_5193,N_5955);
and U6574 (N_6574,N_4390,N_5206);
nor U6575 (N_6575,N_5658,N_4493);
nand U6576 (N_6576,N_4507,N_4356);
nand U6577 (N_6577,N_4929,N_4600);
xor U6578 (N_6578,N_4627,N_5362);
nand U6579 (N_6579,N_5807,N_5987);
nor U6580 (N_6580,N_4360,N_4583);
nor U6581 (N_6581,N_4617,N_5501);
nor U6582 (N_6582,N_4068,N_4949);
nor U6583 (N_6583,N_5174,N_4242);
nand U6584 (N_6584,N_5327,N_4207);
and U6585 (N_6585,N_4027,N_5463);
nor U6586 (N_6586,N_5770,N_5190);
xnor U6587 (N_6587,N_4823,N_4638);
nand U6588 (N_6588,N_5457,N_5131);
and U6589 (N_6589,N_5069,N_5864);
nand U6590 (N_6590,N_4579,N_5014);
and U6591 (N_6591,N_4169,N_5578);
and U6592 (N_6592,N_4495,N_4062);
nor U6593 (N_6593,N_5159,N_4047);
or U6594 (N_6594,N_4602,N_5776);
or U6595 (N_6595,N_5791,N_4141);
nor U6596 (N_6596,N_4065,N_5756);
nor U6597 (N_6597,N_4887,N_5980);
xnor U6598 (N_6598,N_4687,N_4205);
and U6599 (N_6599,N_5352,N_4623);
or U6600 (N_6600,N_5450,N_5251);
and U6601 (N_6601,N_5795,N_5084);
nand U6602 (N_6602,N_4903,N_4458);
xnor U6603 (N_6603,N_4943,N_5992);
xor U6604 (N_6604,N_4948,N_4144);
xnor U6605 (N_6605,N_5433,N_4254);
xor U6606 (N_6606,N_4673,N_4474);
nor U6607 (N_6607,N_5627,N_5746);
nand U6608 (N_6608,N_4366,N_5428);
or U6609 (N_6609,N_4177,N_4809);
xnor U6610 (N_6610,N_4688,N_4189);
or U6611 (N_6611,N_5009,N_5574);
nor U6612 (N_6612,N_4645,N_4500);
nor U6613 (N_6613,N_5492,N_5724);
nand U6614 (N_6614,N_4166,N_5091);
xnor U6615 (N_6615,N_5277,N_5150);
nand U6616 (N_6616,N_5657,N_5008);
and U6617 (N_6617,N_4371,N_5516);
and U6618 (N_6618,N_4450,N_5071);
and U6619 (N_6619,N_4889,N_5942);
xnor U6620 (N_6620,N_5387,N_5507);
xnor U6621 (N_6621,N_4467,N_5283);
and U6622 (N_6622,N_5354,N_5903);
nor U6623 (N_6623,N_4295,N_5345);
xor U6624 (N_6624,N_4455,N_4944);
or U6625 (N_6625,N_4755,N_5468);
nand U6626 (N_6626,N_5371,N_4557);
nor U6627 (N_6627,N_4011,N_5544);
and U6628 (N_6628,N_4836,N_4235);
or U6629 (N_6629,N_5995,N_5530);
or U6630 (N_6630,N_5001,N_5928);
nor U6631 (N_6631,N_4710,N_5364);
nand U6632 (N_6632,N_4379,N_4877);
xnor U6633 (N_6633,N_5385,N_4378);
xnor U6634 (N_6634,N_4131,N_5735);
or U6635 (N_6635,N_4529,N_5949);
and U6636 (N_6636,N_4333,N_5969);
and U6637 (N_6637,N_5766,N_5143);
xor U6638 (N_6638,N_4635,N_5296);
or U6639 (N_6639,N_4666,N_5893);
xnor U6640 (N_6640,N_4819,N_5020);
xnor U6641 (N_6641,N_5304,N_4257);
nand U6642 (N_6642,N_5397,N_5660);
or U6643 (N_6643,N_5443,N_5081);
nor U6644 (N_6644,N_4760,N_5148);
nor U6645 (N_6645,N_4532,N_5471);
or U6646 (N_6646,N_4613,N_4606);
or U6647 (N_6647,N_4978,N_4841);
and U6648 (N_6648,N_5470,N_4691);
nand U6649 (N_6649,N_4281,N_4856);
or U6650 (N_6650,N_4203,N_4322);
nor U6651 (N_6651,N_5897,N_4554);
or U6652 (N_6652,N_5238,N_5863);
nor U6653 (N_6653,N_5258,N_4377);
nor U6654 (N_6654,N_5820,N_4088);
and U6655 (N_6655,N_5054,N_5693);
or U6656 (N_6656,N_4904,N_4698);
nor U6657 (N_6657,N_5386,N_4832);
nor U6658 (N_6658,N_4771,N_4911);
nand U6659 (N_6659,N_5692,N_4694);
and U6660 (N_6660,N_4478,N_5376);
nand U6661 (N_6661,N_5727,N_4938);
nand U6662 (N_6662,N_5977,N_4644);
or U6663 (N_6663,N_5358,N_5172);
or U6664 (N_6664,N_4659,N_5659);
xnor U6665 (N_6665,N_5943,N_5948);
or U6666 (N_6666,N_4076,N_5097);
and U6667 (N_6667,N_5025,N_4985);
nor U6668 (N_6668,N_4202,N_5183);
and U6669 (N_6669,N_5847,N_4712);
nor U6670 (N_6670,N_4883,N_4793);
xnor U6671 (N_6671,N_5583,N_5815);
nand U6672 (N_6672,N_4671,N_5123);
nor U6673 (N_6673,N_5706,N_4019);
or U6674 (N_6674,N_4120,N_4231);
or U6675 (N_6675,N_4908,N_5365);
xnor U6676 (N_6676,N_5597,N_5924);
and U6677 (N_6677,N_4191,N_5332);
or U6678 (N_6678,N_4184,N_5459);
xor U6679 (N_6679,N_4743,N_5147);
nor U6680 (N_6680,N_4092,N_4289);
nor U6681 (N_6681,N_4937,N_4725);
nor U6682 (N_6682,N_5213,N_4338);
or U6683 (N_6683,N_5848,N_4878);
or U6684 (N_6684,N_4368,N_4012);
xor U6685 (N_6685,N_4288,N_5803);
or U6686 (N_6686,N_4418,N_5146);
and U6687 (N_6687,N_5876,N_5343);
or U6688 (N_6688,N_5062,N_5832);
nor U6689 (N_6689,N_5191,N_4683);
or U6690 (N_6690,N_4596,N_5839);
xor U6691 (N_6691,N_5082,N_5256);
xnor U6692 (N_6692,N_4096,N_5293);
or U6693 (N_6693,N_5989,N_5536);
nor U6694 (N_6694,N_5423,N_4428);
or U6695 (N_6695,N_4946,N_5736);
and U6696 (N_6696,N_4584,N_5136);
or U6697 (N_6697,N_5846,N_5967);
or U6698 (N_6698,N_5932,N_4215);
xor U6699 (N_6699,N_5771,N_5857);
nand U6700 (N_6700,N_4023,N_4386);
and U6701 (N_6701,N_5604,N_4423);
and U6702 (N_6702,N_4226,N_4348);
and U6703 (N_6703,N_5101,N_5906);
nor U6704 (N_6704,N_4343,N_5137);
or U6705 (N_6705,N_5904,N_4621);
nor U6706 (N_6706,N_4475,N_4974);
or U6707 (N_6707,N_5458,N_5031);
and U6708 (N_6708,N_4684,N_5800);
xor U6709 (N_6709,N_5032,N_5944);
nor U6710 (N_6710,N_4742,N_4007);
nor U6711 (N_6711,N_4610,N_5568);
nor U6712 (N_6712,N_5553,N_4744);
xor U6713 (N_6713,N_5812,N_4573);
nor U6714 (N_6714,N_5768,N_4504);
or U6715 (N_6715,N_4162,N_4010);
nor U6716 (N_6716,N_5818,N_5512);
nor U6717 (N_6717,N_4147,N_5714);
nand U6718 (N_6718,N_5981,N_4437);
and U6719 (N_6719,N_4653,N_5984);
xor U6720 (N_6720,N_4108,N_4342);
nand U6721 (N_6721,N_4778,N_4828);
or U6722 (N_6722,N_4971,N_5602);
and U6723 (N_6723,N_4605,N_5702);
and U6724 (N_6724,N_4367,N_4058);
or U6725 (N_6725,N_5674,N_5787);
nand U6726 (N_6726,N_5187,N_5179);
nand U6727 (N_6727,N_4213,N_4297);
nor U6728 (N_6728,N_4057,N_5845);
and U6729 (N_6729,N_5377,N_5128);
or U6730 (N_6730,N_5968,N_4447);
or U6731 (N_6731,N_5619,N_5573);
xnor U6732 (N_6732,N_4976,N_4959);
or U6733 (N_6733,N_4572,N_4312);
xor U6734 (N_6734,N_4081,N_5638);
nor U6735 (N_6735,N_5600,N_5026);
nand U6736 (N_6736,N_5067,N_5267);
xnor U6737 (N_6737,N_4524,N_5234);
xnor U6738 (N_6738,N_5642,N_4875);
nand U6739 (N_6739,N_5061,N_4410);
nand U6740 (N_6740,N_4777,N_4313);
xnor U6741 (N_6741,N_5478,N_4868);
nand U6742 (N_6742,N_5749,N_4240);
and U6743 (N_6743,N_5157,N_4498);
or U6744 (N_6744,N_5577,N_5166);
nor U6745 (N_6745,N_4920,N_5665);
xnor U6746 (N_6746,N_5540,N_4381);
nand U6747 (N_6747,N_4734,N_4043);
or U6748 (N_6748,N_5983,N_5053);
or U6749 (N_6749,N_5425,N_5881);
and U6750 (N_6750,N_5156,N_5909);
and U6751 (N_6751,N_5843,N_5938);
nor U6752 (N_6752,N_5999,N_5211);
nand U6753 (N_6753,N_5171,N_4553);
nand U6754 (N_6754,N_5707,N_5814);
nand U6755 (N_6755,N_4840,N_4221);
or U6756 (N_6756,N_4206,N_4695);
or U6757 (N_6757,N_4737,N_5533);
nand U6758 (N_6758,N_4758,N_5711);
xor U6759 (N_6759,N_4087,N_5041);
nor U6760 (N_6760,N_4187,N_5033);
nand U6761 (N_6761,N_4376,N_4250);
or U6762 (N_6762,N_4126,N_4110);
or U6763 (N_6763,N_5772,N_5356);
xor U6764 (N_6764,N_4863,N_4419);
and U6765 (N_6765,N_4562,N_4637);
nor U6766 (N_6766,N_5645,N_4987);
xor U6767 (N_6767,N_4345,N_5882);
xnor U6768 (N_6768,N_5448,N_5650);
or U6769 (N_6769,N_5908,N_5200);
and U6770 (N_6770,N_4918,N_4304);
xnor U6771 (N_6771,N_4407,N_5486);
nand U6772 (N_6772,N_5555,N_4560);
nand U6773 (N_6773,N_4768,N_4269);
and U6774 (N_6774,N_4309,N_5243);
xor U6775 (N_6775,N_4860,N_4430);
and U6776 (N_6776,N_4843,N_4318);
xnor U6777 (N_6777,N_4274,N_5040);
xor U6778 (N_6778,N_4651,N_5687);
xor U6779 (N_6779,N_5467,N_5653);
nand U6780 (N_6780,N_5886,N_5390);
or U6781 (N_6781,N_4415,N_5158);
xnor U6782 (N_6782,N_5654,N_4939);
nor U6783 (N_6783,N_5505,N_5395);
nand U6784 (N_6784,N_4748,N_4798);
nor U6785 (N_6785,N_4647,N_4438);
or U6786 (N_6786,N_5049,N_5628);
xor U6787 (N_6787,N_5110,N_5632);
nand U6788 (N_6788,N_5085,N_4646);
xnor U6789 (N_6789,N_5522,N_4086);
nand U6790 (N_6790,N_5934,N_5905);
nand U6791 (N_6791,N_4188,N_5647);
and U6792 (N_6792,N_5899,N_5284);
and U6793 (N_6793,N_4283,N_4133);
or U6794 (N_6794,N_5322,N_5453);
nand U6795 (N_6795,N_4196,N_4199);
xnor U6796 (N_6796,N_5050,N_4262);
nand U6797 (N_6797,N_5558,N_5705);
nor U6798 (N_6798,N_5965,N_5680);
xnor U6799 (N_6799,N_5668,N_5060);
and U6800 (N_6800,N_5440,N_4757);
nor U6801 (N_6801,N_5872,N_5480);
nand U6802 (N_6802,N_4802,N_5320);
or U6803 (N_6803,N_5792,N_5125);
nor U6804 (N_6804,N_5717,N_4444);
and U6805 (N_6805,N_4722,N_5017);
nand U6806 (N_6806,N_4385,N_4048);
xor U6807 (N_6807,N_5323,N_5037);
or U6808 (N_6808,N_4632,N_4409);
nand U6809 (N_6809,N_5806,N_4480);
nor U6810 (N_6810,N_4454,N_4017);
nand U6811 (N_6811,N_4439,N_5652);
nor U6812 (N_6812,N_5043,N_4469);
and U6813 (N_6813,N_4690,N_4251);
nand U6814 (N_6814,N_5375,N_4153);
or U6815 (N_6815,N_4353,N_4365);
and U6816 (N_6816,N_5827,N_4727);
nor U6817 (N_6817,N_4140,N_5538);
or U6818 (N_6818,N_4222,N_4180);
xnor U6819 (N_6819,N_5681,N_5271);
nor U6820 (N_6820,N_4440,N_5359);
xnor U6821 (N_6821,N_4361,N_4061);
nor U6822 (N_6822,N_4707,N_4164);
or U6823 (N_6823,N_4224,N_5721);
or U6824 (N_6824,N_4781,N_4208);
nand U6825 (N_6825,N_4839,N_4953);
xnor U6826 (N_6826,N_4211,N_4996);
and U6827 (N_6827,N_4749,N_4311);
and U6828 (N_6828,N_4815,N_4375);
and U6829 (N_6829,N_4481,N_4716);
nand U6830 (N_6830,N_4967,N_4788);
or U6831 (N_6831,N_4404,N_5066);
nand U6832 (N_6832,N_4035,N_4411);
xor U6833 (N_6833,N_5978,N_5431);
nand U6834 (N_6834,N_4142,N_5216);
or U6835 (N_6835,N_5254,N_4587);
xnor U6836 (N_6836,N_4190,N_4091);
nand U6837 (N_6837,N_4805,N_4463);
nand U6838 (N_6838,N_5027,N_4282);
and U6839 (N_6839,N_4753,N_5535);
xnor U6840 (N_6840,N_5713,N_4405);
and U6841 (N_6841,N_4066,N_4909);
or U6842 (N_6842,N_4105,N_5052);
and U6843 (N_6843,N_4723,N_4060);
and U6844 (N_6844,N_4218,N_4460);
nor U6845 (N_6845,N_5083,N_4897);
nor U6846 (N_6846,N_5588,N_4998);
or U6847 (N_6847,N_4910,N_4616);
nor U6848 (N_6848,N_5142,N_4435);
and U6849 (N_6849,N_5209,N_4069);
nor U6850 (N_6850,N_4001,N_4593);
or U6851 (N_6851,N_4466,N_5608);
nor U6852 (N_6852,N_5466,N_4401);
nand U6853 (N_6853,N_4801,N_4064);
nor U6854 (N_6854,N_4729,N_5497);
xor U6855 (N_6855,N_4416,N_5140);
and U6856 (N_6856,N_5056,N_4580);
xnor U6857 (N_6857,N_4209,N_4813);
nand U6858 (N_6858,N_5350,N_5151);
nor U6859 (N_6859,N_4505,N_4079);
xnor U6860 (N_6860,N_4564,N_5310);
nand U6861 (N_6861,N_5587,N_4008);
and U6862 (N_6862,N_4797,N_5849);
or U6863 (N_6863,N_5388,N_4041);
nand U6864 (N_6864,N_5629,N_4569);
nand U6865 (N_6865,N_4762,N_5670);
xnor U6866 (N_6866,N_5374,N_5880);
nor U6867 (N_6867,N_5475,N_4528);
xor U6868 (N_6868,N_4185,N_4999);
and U6869 (N_6869,N_5675,N_5567);
xnor U6870 (N_6870,N_5935,N_4000);
and U6871 (N_6871,N_4958,N_5651);
nor U6872 (N_6872,N_4574,N_4577);
xnor U6873 (N_6873,N_4253,N_5926);
or U6874 (N_6874,N_5160,N_5704);
nor U6875 (N_6875,N_5413,N_4548);
nand U6876 (N_6876,N_5115,N_5330);
or U6877 (N_6877,N_5614,N_5121);
nor U6878 (N_6878,N_4983,N_5100);
nor U6879 (N_6879,N_5797,N_5381);
nor U6880 (N_6880,N_4067,N_4022);
nor U6881 (N_6881,N_5215,N_4214);
and U6882 (N_6882,N_5426,N_5117);
nor U6883 (N_6883,N_5484,N_5514);
nand U6884 (N_6884,N_4715,N_4774);
nor U6885 (N_6885,N_4453,N_4359);
xnor U6886 (N_6886,N_5185,N_4849);
and U6887 (N_6887,N_5931,N_4830);
nor U6888 (N_6888,N_4736,N_4212);
nand U6889 (N_6889,N_4982,N_5454);
nand U6890 (N_6890,N_4884,N_5479);
and U6891 (N_6891,N_5655,N_4846);
and U6892 (N_6892,N_4589,N_5355);
nor U6893 (N_6893,N_5204,N_4858);
nor U6894 (N_6894,N_5584,N_5241);
nor U6895 (N_6895,N_4677,N_4799);
and U6896 (N_6896,N_5403,N_5360);
nand U6897 (N_6897,N_4770,N_5246);
and U6898 (N_6898,N_5731,N_5537);
nand U6899 (N_6899,N_5394,N_5042);
xnor U6900 (N_6900,N_5230,N_5490);
or U6901 (N_6901,N_4919,N_4259);
nor U6902 (N_6902,N_5266,N_5415);
nand U6903 (N_6903,N_4117,N_5370);
and U6904 (N_6904,N_4099,N_5566);
xnor U6905 (N_6905,N_5077,N_4431);
or U6906 (N_6906,N_4765,N_4759);
nand U6907 (N_6907,N_5261,N_5319);
xnor U6908 (N_6908,N_5836,N_5120);
nand U6909 (N_6909,N_5289,N_5598);
nor U6910 (N_6910,N_4477,N_5964);
and U6911 (N_6911,N_5579,N_5741);
and U6912 (N_6912,N_4526,N_5682);
nor U6913 (N_6913,N_5837,N_4568);
and U6914 (N_6914,N_5858,N_4492);
and U6915 (N_6915,N_4434,N_5895);
nand U6916 (N_6916,N_5161,N_5139);
or U6917 (N_6917,N_4820,N_4921);
and U6918 (N_6918,N_5003,N_4790);
or U6919 (N_6919,N_4942,N_4103);
nand U6920 (N_6920,N_5754,N_5233);
or U6921 (N_6921,N_4628,N_4266);
nor U6922 (N_6922,N_4713,N_4051);
nor U6923 (N_6923,N_4540,N_5873);
or U6924 (N_6924,N_4876,N_5078);
nand U6925 (N_6925,N_4751,N_4089);
nand U6926 (N_6926,N_5297,N_5422);
nand U6927 (N_6927,N_4620,N_5456);
nand U6928 (N_6928,N_4118,N_4881);
xnor U6929 (N_6929,N_5192,N_5691);
or U6930 (N_6930,N_5461,N_5790);
nand U6931 (N_6931,N_5476,N_4817);
nor U6932 (N_6932,N_5088,N_5298);
or U6933 (N_6933,N_5788,N_4542);
xor U6934 (N_6934,N_4853,N_4136);
or U6935 (N_6935,N_4894,N_5798);
or U6936 (N_6936,N_4044,N_5511);
and U6937 (N_6937,N_5257,N_5224);
xnor U6938 (N_6938,N_4094,N_5438);
and U6939 (N_6939,N_4590,N_4886);
or U6940 (N_6940,N_4393,N_4711);
nor U6941 (N_6941,N_5676,N_5805);
xor U6942 (N_6942,N_5709,N_5686);
xnor U6943 (N_6943,N_5153,N_5004);
nor U6944 (N_6944,N_4158,N_5219);
xnor U6945 (N_6945,N_5740,N_4156);
or U6946 (N_6946,N_4658,N_4384);
nor U6947 (N_6947,N_4675,N_5051);
or U6948 (N_6948,N_4476,N_5202);
or U6949 (N_6949,N_4107,N_4652);
xor U6950 (N_6950,N_5825,N_5605);
and U6951 (N_6951,N_4489,N_5249);
nand U6952 (N_6952,N_5154,N_4038);
and U6953 (N_6953,N_5722,N_5034);
or U6954 (N_6954,N_4329,N_5669);
or U6955 (N_6955,N_4247,N_4531);
and U6956 (N_6956,N_4299,N_5630);
nand U6957 (N_6957,N_4152,N_4672);
and U6958 (N_6958,N_4292,N_5227);
xnor U6959 (N_6959,N_4806,N_5168);
xnor U6960 (N_6960,N_4025,N_4324);
xor U6961 (N_6961,N_4775,N_4618);
nand U6962 (N_6962,N_5255,N_5055);
nor U6963 (N_6963,N_5250,N_4275);
and U6964 (N_6964,N_4966,N_4693);
nor U6965 (N_6965,N_4810,N_4291);
and U6966 (N_6966,N_4101,N_4629);
nor U6967 (N_6967,N_4523,N_5019);
nand U6968 (N_6968,N_4445,N_4965);
or U6969 (N_6969,N_4864,N_5473);
nor U6970 (N_6970,N_4917,N_4764);
nor U6971 (N_6971,N_4009,N_5742);
or U6972 (N_6972,N_4227,N_5099);
nor U6973 (N_6973,N_5570,N_5958);
nand U6974 (N_6974,N_5432,N_5696);
nor U6975 (N_6975,N_4848,N_5198);
xnor U6976 (N_6976,N_5427,N_4090);
nand U6977 (N_6977,N_4139,N_5616);
nor U6978 (N_6978,N_5809,N_4803);
nor U6979 (N_6979,N_4293,N_5816);
xnor U6980 (N_6980,N_4566,N_4174);
nor U6981 (N_6981,N_4037,N_4924);
nand U6982 (N_6982,N_4422,N_4717);
or U6983 (N_6983,N_4576,N_4611);
or U6984 (N_6984,N_4516,N_4852);
xnor U6985 (N_6985,N_5871,N_5622);
nand U6986 (N_6986,N_4719,N_4663);
and U6987 (N_6987,N_4181,N_5315);
xnor U6988 (N_6988,N_4234,N_5891);
or U6989 (N_6989,N_5870,N_5012);
or U6990 (N_6990,N_4285,N_4988);
and U6991 (N_6991,N_4335,N_4194);
xor U6992 (N_6992,N_4050,N_4132);
xnor U6993 (N_6993,N_4056,N_5649);
and U6994 (N_6994,N_5477,N_4890);
or U6995 (N_6995,N_5487,N_5716);
xnor U6996 (N_6996,N_5197,N_5018);
nand U6997 (N_6997,N_4699,N_4323);
or U6998 (N_6998,N_4298,N_4284);
nand U6999 (N_6999,N_4927,N_4872);
xnor U7000 (N_7000,N_5202,N_5915);
nor U7001 (N_7001,N_5633,N_5366);
or U7002 (N_7002,N_4320,N_5683);
nand U7003 (N_7003,N_5224,N_4758);
nor U7004 (N_7004,N_4748,N_4662);
xor U7005 (N_7005,N_5490,N_5936);
and U7006 (N_7006,N_4361,N_4229);
xnor U7007 (N_7007,N_5900,N_4379);
nand U7008 (N_7008,N_5907,N_4065);
or U7009 (N_7009,N_5789,N_4540);
nor U7010 (N_7010,N_5709,N_5589);
nor U7011 (N_7011,N_4284,N_4431);
and U7012 (N_7012,N_4500,N_4879);
nand U7013 (N_7013,N_5422,N_5783);
nor U7014 (N_7014,N_5808,N_4103);
and U7015 (N_7015,N_5977,N_5005);
xnor U7016 (N_7016,N_4257,N_5855);
nor U7017 (N_7017,N_4600,N_4676);
nor U7018 (N_7018,N_4593,N_4342);
or U7019 (N_7019,N_5130,N_4155);
nand U7020 (N_7020,N_4444,N_4231);
or U7021 (N_7021,N_5468,N_5232);
nand U7022 (N_7022,N_4800,N_5184);
nor U7023 (N_7023,N_5483,N_5148);
nand U7024 (N_7024,N_5434,N_4282);
nor U7025 (N_7025,N_4988,N_4731);
nor U7026 (N_7026,N_5897,N_5241);
nor U7027 (N_7027,N_5230,N_5426);
and U7028 (N_7028,N_4502,N_4919);
nor U7029 (N_7029,N_4431,N_4125);
and U7030 (N_7030,N_4563,N_4697);
or U7031 (N_7031,N_5501,N_4293);
nand U7032 (N_7032,N_4213,N_4836);
xor U7033 (N_7033,N_5027,N_5104);
and U7034 (N_7034,N_5815,N_4721);
xnor U7035 (N_7035,N_5252,N_5765);
nor U7036 (N_7036,N_5807,N_4163);
nor U7037 (N_7037,N_4501,N_5636);
and U7038 (N_7038,N_4383,N_4385);
and U7039 (N_7039,N_5284,N_4770);
nand U7040 (N_7040,N_4417,N_4084);
xnor U7041 (N_7041,N_4112,N_4373);
nand U7042 (N_7042,N_4779,N_4986);
and U7043 (N_7043,N_5749,N_5254);
nor U7044 (N_7044,N_4102,N_4253);
and U7045 (N_7045,N_4814,N_4033);
nor U7046 (N_7046,N_4769,N_5348);
nand U7047 (N_7047,N_4815,N_5090);
and U7048 (N_7048,N_5462,N_5742);
or U7049 (N_7049,N_4115,N_4109);
nor U7050 (N_7050,N_4638,N_4501);
nand U7051 (N_7051,N_5586,N_4149);
or U7052 (N_7052,N_4795,N_4549);
nand U7053 (N_7053,N_5540,N_5627);
and U7054 (N_7054,N_4506,N_4916);
xnor U7055 (N_7055,N_5262,N_4763);
and U7056 (N_7056,N_4332,N_4543);
or U7057 (N_7057,N_4921,N_4721);
or U7058 (N_7058,N_5910,N_4494);
and U7059 (N_7059,N_5713,N_5579);
nand U7060 (N_7060,N_5271,N_5066);
xor U7061 (N_7061,N_5079,N_5189);
and U7062 (N_7062,N_5833,N_5638);
nor U7063 (N_7063,N_5929,N_5892);
nand U7064 (N_7064,N_4210,N_4355);
nor U7065 (N_7065,N_5750,N_5209);
nand U7066 (N_7066,N_5426,N_4120);
nand U7067 (N_7067,N_4219,N_5416);
and U7068 (N_7068,N_5626,N_4297);
nor U7069 (N_7069,N_5764,N_4879);
nand U7070 (N_7070,N_4280,N_5857);
nand U7071 (N_7071,N_5415,N_4527);
nor U7072 (N_7072,N_4049,N_4944);
and U7073 (N_7073,N_4803,N_4100);
or U7074 (N_7074,N_5034,N_5820);
and U7075 (N_7075,N_5076,N_4903);
or U7076 (N_7076,N_4416,N_5064);
or U7077 (N_7077,N_5744,N_4921);
nor U7078 (N_7078,N_5709,N_4563);
nand U7079 (N_7079,N_4927,N_5325);
xnor U7080 (N_7080,N_5005,N_5850);
nor U7081 (N_7081,N_5938,N_5867);
xnor U7082 (N_7082,N_4404,N_4566);
xnor U7083 (N_7083,N_5091,N_5521);
nor U7084 (N_7084,N_4597,N_5340);
or U7085 (N_7085,N_4693,N_5680);
nor U7086 (N_7086,N_5078,N_4289);
and U7087 (N_7087,N_4958,N_5230);
nand U7088 (N_7088,N_4689,N_4575);
nor U7089 (N_7089,N_5915,N_5096);
nor U7090 (N_7090,N_4467,N_5694);
nand U7091 (N_7091,N_4957,N_5183);
or U7092 (N_7092,N_4014,N_5341);
nand U7093 (N_7093,N_5165,N_4537);
nand U7094 (N_7094,N_4655,N_4947);
or U7095 (N_7095,N_4527,N_5110);
or U7096 (N_7096,N_5818,N_5250);
nor U7097 (N_7097,N_4431,N_5640);
nand U7098 (N_7098,N_5781,N_4511);
nand U7099 (N_7099,N_5478,N_5859);
nand U7100 (N_7100,N_4157,N_4517);
xnor U7101 (N_7101,N_5185,N_4253);
nor U7102 (N_7102,N_5724,N_5123);
or U7103 (N_7103,N_5403,N_5645);
nor U7104 (N_7104,N_5574,N_4523);
and U7105 (N_7105,N_4088,N_5016);
xnor U7106 (N_7106,N_4799,N_4396);
xnor U7107 (N_7107,N_5528,N_4791);
or U7108 (N_7108,N_5238,N_4353);
xnor U7109 (N_7109,N_5448,N_4697);
or U7110 (N_7110,N_4353,N_5342);
nor U7111 (N_7111,N_5219,N_5931);
and U7112 (N_7112,N_4711,N_4410);
and U7113 (N_7113,N_4104,N_4029);
xor U7114 (N_7114,N_5616,N_4497);
or U7115 (N_7115,N_4202,N_4913);
nor U7116 (N_7116,N_4455,N_4616);
nor U7117 (N_7117,N_4175,N_4880);
nand U7118 (N_7118,N_4248,N_5241);
xnor U7119 (N_7119,N_5161,N_4076);
xor U7120 (N_7120,N_4033,N_5132);
or U7121 (N_7121,N_5248,N_5966);
xor U7122 (N_7122,N_5651,N_4759);
and U7123 (N_7123,N_4504,N_4549);
and U7124 (N_7124,N_4775,N_5020);
or U7125 (N_7125,N_4049,N_5265);
xor U7126 (N_7126,N_4599,N_5021);
and U7127 (N_7127,N_4473,N_5717);
and U7128 (N_7128,N_5415,N_4657);
nand U7129 (N_7129,N_5803,N_4597);
and U7130 (N_7130,N_5984,N_5129);
nand U7131 (N_7131,N_5218,N_5733);
nor U7132 (N_7132,N_5066,N_5703);
xnor U7133 (N_7133,N_4829,N_4806);
or U7134 (N_7134,N_5826,N_4121);
nand U7135 (N_7135,N_4288,N_5142);
and U7136 (N_7136,N_5631,N_5633);
and U7137 (N_7137,N_5022,N_4559);
nand U7138 (N_7138,N_4375,N_4114);
nor U7139 (N_7139,N_4365,N_5787);
xor U7140 (N_7140,N_4867,N_5175);
and U7141 (N_7141,N_4964,N_5618);
nand U7142 (N_7142,N_5819,N_5743);
nand U7143 (N_7143,N_5263,N_5772);
nand U7144 (N_7144,N_4436,N_5264);
or U7145 (N_7145,N_5412,N_4176);
or U7146 (N_7146,N_5727,N_5755);
or U7147 (N_7147,N_4243,N_5086);
xnor U7148 (N_7148,N_4692,N_4089);
nor U7149 (N_7149,N_4292,N_4993);
or U7150 (N_7150,N_4556,N_4218);
xnor U7151 (N_7151,N_5258,N_5133);
nand U7152 (N_7152,N_5643,N_4899);
nand U7153 (N_7153,N_4224,N_5146);
or U7154 (N_7154,N_4356,N_4389);
nand U7155 (N_7155,N_4542,N_4662);
nand U7156 (N_7156,N_5373,N_4427);
xor U7157 (N_7157,N_4886,N_5860);
nand U7158 (N_7158,N_5098,N_4313);
or U7159 (N_7159,N_5736,N_4589);
nor U7160 (N_7160,N_4020,N_4705);
or U7161 (N_7161,N_5715,N_5265);
nand U7162 (N_7162,N_4955,N_5082);
xor U7163 (N_7163,N_5696,N_5361);
nand U7164 (N_7164,N_5770,N_4658);
and U7165 (N_7165,N_5645,N_4025);
nand U7166 (N_7166,N_4573,N_4640);
nor U7167 (N_7167,N_5161,N_5912);
nor U7168 (N_7168,N_5370,N_4446);
and U7169 (N_7169,N_5547,N_4325);
and U7170 (N_7170,N_5151,N_5016);
nand U7171 (N_7171,N_5277,N_4121);
nor U7172 (N_7172,N_4818,N_5177);
xnor U7173 (N_7173,N_5307,N_4169);
nor U7174 (N_7174,N_4710,N_4795);
nand U7175 (N_7175,N_4324,N_4014);
xnor U7176 (N_7176,N_4394,N_5967);
and U7177 (N_7177,N_5896,N_4421);
or U7178 (N_7178,N_5223,N_4883);
and U7179 (N_7179,N_4157,N_4398);
and U7180 (N_7180,N_5942,N_5104);
and U7181 (N_7181,N_4050,N_4428);
or U7182 (N_7182,N_4538,N_5139);
or U7183 (N_7183,N_5206,N_4805);
or U7184 (N_7184,N_5509,N_5329);
xor U7185 (N_7185,N_5662,N_4082);
xor U7186 (N_7186,N_4626,N_4405);
nand U7187 (N_7187,N_4989,N_5262);
and U7188 (N_7188,N_4370,N_4528);
nand U7189 (N_7189,N_4257,N_5776);
nand U7190 (N_7190,N_4130,N_4233);
and U7191 (N_7191,N_5811,N_4233);
nand U7192 (N_7192,N_5305,N_4369);
nand U7193 (N_7193,N_5378,N_4870);
xnor U7194 (N_7194,N_4144,N_4881);
nor U7195 (N_7195,N_4930,N_4674);
nand U7196 (N_7196,N_5819,N_5850);
or U7197 (N_7197,N_5107,N_5168);
nand U7198 (N_7198,N_5281,N_4337);
xor U7199 (N_7199,N_4083,N_5567);
nand U7200 (N_7200,N_4939,N_4496);
nor U7201 (N_7201,N_5109,N_4450);
or U7202 (N_7202,N_4582,N_5918);
nor U7203 (N_7203,N_4034,N_4649);
or U7204 (N_7204,N_5417,N_4023);
and U7205 (N_7205,N_5161,N_4081);
nor U7206 (N_7206,N_4640,N_5720);
xnor U7207 (N_7207,N_5612,N_4516);
or U7208 (N_7208,N_4712,N_4723);
nor U7209 (N_7209,N_4079,N_4893);
nand U7210 (N_7210,N_4268,N_4609);
nor U7211 (N_7211,N_4037,N_4715);
xnor U7212 (N_7212,N_5961,N_4562);
or U7213 (N_7213,N_4273,N_5847);
nor U7214 (N_7214,N_4638,N_5414);
and U7215 (N_7215,N_4418,N_4768);
nand U7216 (N_7216,N_5801,N_5424);
nand U7217 (N_7217,N_4009,N_5394);
and U7218 (N_7218,N_5145,N_4975);
xor U7219 (N_7219,N_5630,N_4446);
xnor U7220 (N_7220,N_5024,N_5079);
or U7221 (N_7221,N_4398,N_5666);
nand U7222 (N_7222,N_5217,N_5729);
nand U7223 (N_7223,N_5043,N_5794);
nand U7224 (N_7224,N_4358,N_5615);
nand U7225 (N_7225,N_5870,N_5815);
nand U7226 (N_7226,N_5048,N_5930);
or U7227 (N_7227,N_5960,N_4732);
and U7228 (N_7228,N_4132,N_4484);
xnor U7229 (N_7229,N_5396,N_4145);
and U7230 (N_7230,N_5447,N_5424);
and U7231 (N_7231,N_4319,N_4817);
and U7232 (N_7232,N_4078,N_4735);
nand U7233 (N_7233,N_4650,N_4461);
and U7234 (N_7234,N_5992,N_4444);
and U7235 (N_7235,N_4730,N_5098);
xnor U7236 (N_7236,N_4772,N_4047);
nor U7237 (N_7237,N_4447,N_5407);
or U7238 (N_7238,N_4453,N_5730);
nor U7239 (N_7239,N_4227,N_5523);
nand U7240 (N_7240,N_5643,N_5798);
nor U7241 (N_7241,N_4993,N_5164);
xor U7242 (N_7242,N_5410,N_4650);
nand U7243 (N_7243,N_4585,N_5099);
xor U7244 (N_7244,N_4287,N_4616);
or U7245 (N_7245,N_4880,N_5504);
or U7246 (N_7246,N_4244,N_5243);
and U7247 (N_7247,N_4156,N_5599);
xnor U7248 (N_7248,N_5895,N_4606);
xnor U7249 (N_7249,N_4054,N_5548);
nand U7250 (N_7250,N_4933,N_4742);
or U7251 (N_7251,N_4541,N_5654);
xnor U7252 (N_7252,N_4576,N_4068);
or U7253 (N_7253,N_5327,N_4809);
or U7254 (N_7254,N_4033,N_4551);
xnor U7255 (N_7255,N_5922,N_4152);
and U7256 (N_7256,N_5532,N_4071);
xor U7257 (N_7257,N_4168,N_5196);
nor U7258 (N_7258,N_5277,N_5630);
xnor U7259 (N_7259,N_5593,N_4683);
nand U7260 (N_7260,N_4813,N_5881);
and U7261 (N_7261,N_4492,N_4715);
and U7262 (N_7262,N_5353,N_5023);
or U7263 (N_7263,N_5572,N_4843);
and U7264 (N_7264,N_5129,N_4416);
nand U7265 (N_7265,N_4276,N_5609);
xor U7266 (N_7266,N_5050,N_5394);
xnor U7267 (N_7267,N_5440,N_5088);
and U7268 (N_7268,N_5230,N_4509);
and U7269 (N_7269,N_5918,N_4358);
and U7270 (N_7270,N_4965,N_5146);
and U7271 (N_7271,N_4479,N_5734);
and U7272 (N_7272,N_5314,N_5670);
nand U7273 (N_7273,N_4041,N_5277);
or U7274 (N_7274,N_4289,N_4779);
or U7275 (N_7275,N_5489,N_5472);
or U7276 (N_7276,N_4425,N_4587);
xnor U7277 (N_7277,N_4242,N_5263);
or U7278 (N_7278,N_5741,N_4431);
nor U7279 (N_7279,N_4971,N_4705);
nor U7280 (N_7280,N_5683,N_5448);
or U7281 (N_7281,N_5766,N_5211);
or U7282 (N_7282,N_5738,N_4639);
or U7283 (N_7283,N_5087,N_4093);
and U7284 (N_7284,N_4559,N_4947);
nor U7285 (N_7285,N_5547,N_4524);
or U7286 (N_7286,N_5840,N_4277);
xor U7287 (N_7287,N_4977,N_5439);
nand U7288 (N_7288,N_5787,N_5410);
nor U7289 (N_7289,N_5727,N_5047);
nor U7290 (N_7290,N_5028,N_5369);
nor U7291 (N_7291,N_4812,N_5949);
xor U7292 (N_7292,N_4082,N_5162);
nand U7293 (N_7293,N_4960,N_4237);
xnor U7294 (N_7294,N_4547,N_5354);
nand U7295 (N_7295,N_4513,N_5614);
and U7296 (N_7296,N_5250,N_5124);
xor U7297 (N_7297,N_5380,N_4998);
or U7298 (N_7298,N_5031,N_5578);
xnor U7299 (N_7299,N_5263,N_5324);
and U7300 (N_7300,N_5785,N_4665);
or U7301 (N_7301,N_4540,N_4708);
nand U7302 (N_7302,N_5908,N_5836);
xor U7303 (N_7303,N_5540,N_5082);
nand U7304 (N_7304,N_5396,N_5535);
and U7305 (N_7305,N_4648,N_5405);
nand U7306 (N_7306,N_4972,N_4423);
xnor U7307 (N_7307,N_5200,N_4201);
nand U7308 (N_7308,N_5485,N_5675);
nor U7309 (N_7309,N_4751,N_4964);
xor U7310 (N_7310,N_4211,N_5229);
and U7311 (N_7311,N_5219,N_5061);
and U7312 (N_7312,N_5902,N_5245);
xnor U7313 (N_7313,N_5833,N_5038);
nor U7314 (N_7314,N_4607,N_4480);
xnor U7315 (N_7315,N_5813,N_4860);
xnor U7316 (N_7316,N_4044,N_4970);
nor U7317 (N_7317,N_4946,N_5383);
and U7318 (N_7318,N_5486,N_4431);
or U7319 (N_7319,N_4106,N_4847);
or U7320 (N_7320,N_4415,N_4853);
xnor U7321 (N_7321,N_5114,N_4131);
or U7322 (N_7322,N_4283,N_5567);
xnor U7323 (N_7323,N_4017,N_4751);
nand U7324 (N_7324,N_4239,N_5847);
and U7325 (N_7325,N_4674,N_5077);
xor U7326 (N_7326,N_5591,N_5262);
and U7327 (N_7327,N_4574,N_4171);
and U7328 (N_7328,N_5321,N_5212);
or U7329 (N_7329,N_4977,N_4791);
nand U7330 (N_7330,N_4755,N_5044);
nor U7331 (N_7331,N_4371,N_5078);
or U7332 (N_7332,N_5192,N_5667);
nor U7333 (N_7333,N_4418,N_4214);
nor U7334 (N_7334,N_5236,N_4109);
nand U7335 (N_7335,N_4801,N_4933);
nand U7336 (N_7336,N_5183,N_5870);
or U7337 (N_7337,N_4977,N_5450);
xnor U7338 (N_7338,N_4652,N_5135);
nand U7339 (N_7339,N_4138,N_4413);
or U7340 (N_7340,N_4038,N_5101);
or U7341 (N_7341,N_4179,N_5410);
nor U7342 (N_7342,N_5446,N_4646);
or U7343 (N_7343,N_5836,N_5617);
nand U7344 (N_7344,N_4895,N_5280);
xor U7345 (N_7345,N_5403,N_4732);
nor U7346 (N_7346,N_4107,N_5962);
or U7347 (N_7347,N_5273,N_5866);
nor U7348 (N_7348,N_4917,N_5895);
nor U7349 (N_7349,N_5069,N_5504);
and U7350 (N_7350,N_5043,N_4944);
xor U7351 (N_7351,N_4823,N_5839);
and U7352 (N_7352,N_5988,N_4798);
or U7353 (N_7353,N_5434,N_5205);
nor U7354 (N_7354,N_5702,N_4421);
and U7355 (N_7355,N_4454,N_5293);
xnor U7356 (N_7356,N_5655,N_5923);
or U7357 (N_7357,N_4175,N_4646);
or U7358 (N_7358,N_4244,N_4188);
and U7359 (N_7359,N_4267,N_5429);
or U7360 (N_7360,N_4402,N_5339);
nand U7361 (N_7361,N_4859,N_5305);
and U7362 (N_7362,N_4784,N_5733);
and U7363 (N_7363,N_5833,N_5551);
nor U7364 (N_7364,N_5801,N_5610);
and U7365 (N_7365,N_5411,N_5066);
xor U7366 (N_7366,N_4296,N_5084);
nor U7367 (N_7367,N_5852,N_5842);
and U7368 (N_7368,N_5942,N_4819);
and U7369 (N_7369,N_5838,N_5225);
xnor U7370 (N_7370,N_5371,N_5378);
and U7371 (N_7371,N_5686,N_5103);
xnor U7372 (N_7372,N_4359,N_4125);
xor U7373 (N_7373,N_5245,N_4228);
xor U7374 (N_7374,N_4488,N_4957);
nor U7375 (N_7375,N_5653,N_5927);
nor U7376 (N_7376,N_4500,N_4095);
nor U7377 (N_7377,N_4578,N_4379);
and U7378 (N_7378,N_5116,N_4734);
nand U7379 (N_7379,N_4433,N_4350);
and U7380 (N_7380,N_4432,N_4765);
nor U7381 (N_7381,N_4611,N_4623);
nor U7382 (N_7382,N_4221,N_4824);
or U7383 (N_7383,N_4384,N_4979);
nand U7384 (N_7384,N_4910,N_4956);
xor U7385 (N_7385,N_5053,N_5447);
nor U7386 (N_7386,N_4482,N_5812);
xnor U7387 (N_7387,N_5109,N_4954);
nor U7388 (N_7388,N_5407,N_5726);
nor U7389 (N_7389,N_5148,N_5578);
nand U7390 (N_7390,N_4819,N_5274);
and U7391 (N_7391,N_4249,N_4690);
nand U7392 (N_7392,N_4946,N_5415);
nor U7393 (N_7393,N_4530,N_5417);
nand U7394 (N_7394,N_5331,N_5974);
or U7395 (N_7395,N_5355,N_4105);
or U7396 (N_7396,N_4509,N_5495);
nor U7397 (N_7397,N_4953,N_4748);
or U7398 (N_7398,N_5442,N_4204);
xor U7399 (N_7399,N_5084,N_4175);
nand U7400 (N_7400,N_4610,N_4475);
or U7401 (N_7401,N_5031,N_5165);
nor U7402 (N_7402,N_5087,N_4367);
or U7403 (N_7403,N_4664,N_4452);
xnor U7404 (N_7404,N_5342,N_4138);
nor U7405 (N_7405,N_4909,N_5745);
or U7406 (N_7406,N_4950,N_4811);
nand U7407 (N_7407,N_4927,N_4626);
xor U7408 (N_7408,N_5195,N_5481);
nor U7409 (N_7409,N_4175,N_4804);
xnor U7410 (N_7410,N_4576,N_5283);
or U7411 (N_7411,N_5088,N_5453);
nor U7412 (N_7412,N_4265,N_4623);
xor U7413 (N_7413,N_5896,N_4127);
xor U7414 (N_7414,N_4279,N_5728);
nor U7415 (N_7415,N_4038,N_4308);
xor U7416 (N_7416,N_5061,N_4120);
and U7417 (N_7417,N_5884,N_4448);
xnor U7418 (N_7418,N_5959,N_5183);
nand U7419 (N_7419,N_5911,N_4854);
nand U7420 (N_7420,N_5054,N_4246);
or U7421 (N_7421,N_4581,N_4052);
nor U7422 (N_7422,N_5407,N_5108);
nor U7423 (N_7423,N_5738,N_5452);
or U7424 (N_7424,N_5600,N_4934);
nor U7425 (N_7425,N_5927,N_5644);
or U7426 (N_7426,N_4423,N_4595);
or U7427 (N_7427,N_5608,N_4812);
nor U7428 (N_7428,N_5258,N_5617);
or U7429 (N_7429,N_5877,N_5113);
or U7430 (N_7430,N_5371,N_5665);
and U7431 (N_7431,N_4905,N_4422);
and U7432 (N_7432,N_5496,N_5199);
or U7433 (N_7433,N_5208,N_4403);
nand U7434 (N_7434,N_5819,N_5942);
nand U7435 (N_7435,N_4883,N_4181);
nand U7436 (N_7436,N_5081,N_5118);
nor U7437 (N_7437,N_5918,N_4438);
nand U7438 (N_7438,N_4818,N_5965);
nor U7439 (N_7439,N_5799,N_4403);
nor U7440 (N_7440,N_4233,N_5755);
or U7441 (N_7441,N_5952,N_4168);
and U7442 (N_7442,N_5148,N_5488);
and U7443 (N_7443,N_5249,N_4109);
nand U7444 (N_7444,N_4821,N_5600);
nor U7445 (N_7445,N_5478,N_4397);
xor U7446 (N_7446,N_5448,N_5691);
nor U7447 (N_7447,N_5525,N_4200);
or U7448 (N_7448,N_4007,N_5940);
nor U7449 (N_7449,N_4288,N_4395);
nand U7450 (N_7450,N_5919,N_5815);
xnor U7451 (N_7451,N_4790,N_4403);
xor U7452 (N_7452,N_4021,N_4599);
xnor U7453 (N_7453,N_4384,N_4360);
xor U7454 (N_7454,N_5629,N_5708);
xnor U7455 (N_7455,N_5915,N_4156);
or U7456 (N_7456,N_5583,N_5769);
or U7457 (N_7457,N_4079,N_4261);
or U7458 (N_7458,N_4121,N_5066);
nand U7459 (N_7459,N_5880,N_5284);
and U7460 (N_7460,N_5925,N_5850);
and U7461 (N_7461,N_5896,N_4888);
xnor U7462 (N_7462,N_5306,N_4066);
xor U7463 (N_7463,N_4918,N_4343);
and U7464 (N_7464,N_4317,N_5625);
and U7465 (N_7465,N_5616,N_5168);
or U7466 (N_7466,N_5361,N_4739);
and U7467 (N_7467,N_4312,N_5422);
nor U7468 (N_7468,N_5040,N_5305);
nand U7469 (N_7469,N_4800,N_4218);
nand U7470 (N_7470,N_5419,N_4814);
nand U7471 (N_7471,N_4460,N_4452);
or U7472 (N_7472,N_4429,N_5278);
xnor U7473 (N_7473,N_5086,N_4043);
or U7474 (N_7474,N_5131,N_4103);
xnor U7475 (N_7475,N_4078,N_5787);
and U7476 (N_7476,N_4516,N_4226);
and U7477 (N_7477,N_5108,N_5361);
xnor U7478 (N_7478,N_4026,N_4161);
or U7479 (N_7479,N_5446,N_4861);
nor U7480 (N_7480,N_5131,N_5335);
xor U7481 (N_7481,N_4379,N_4217);
or U7482 (N_7482,N_4684,N_5511);
and U7483 (N_7483,N_4590,N_5184);
or U7484 (N_7484,N_5715,N_4632);
xor U7485 (N_7485,N_5507,N_4922);
xor U7486 (N_7486,N_4395,N_5555);
and U7487 (N_7487,N_4160,N_5240);
xnor U7488 (N_7488,N_5921,N_5237);
xor U7489 (N_7489,N_4725,N_5753);
xnor U7490 (N_7490,N_4445,N_5680);
nand U7491 (N_7491,N_5969,N_5124);
or U7492 (N_7492,N_4191,N_4211);
nor U7493 (N_7493,N_5844,N_4329);
nand U7494 (N_7494,N_5148,N_5353);
nand U7495 (N_7495,N_4500,N_5846);
nand U7496 (N_7496,N_4278,N_4364);
nand U7497 (N_7497,N_4434,N_5381);
nor U7498 (N_7498,N_5759,N_4530);
nor U7499 (N_7499,N_5096,N_5742);
nand U7500 (N_7500,N_4050,N_5948);
nand U7501 (N_7501,N_4400,N_5936);
nor U7502 (N_7502,N_5757,N_5167);
nand U7503 (N_7503,N_5431,N_5312);
xor U7504 (N_7504,N_5182,N_4858);
and U7505 (N_7505,N_5523,N_4318);
and U7506 (N_7506,N_4373,N_4883);
nor U7507 (N_7507,N_5445,N_4007);
nand U7508 (N_7508,N_5879,N_5821);
nand U7509 (N_7509,N_4754,N_5002);
nor U7510 (N_7510,N_5949,N_5935);
and U7511 (N_7511,N_5046,N_4974);
xor U7512 (N_7512,N_4723,N_4530);
and U7513 (N_7513,N_4718,N_5349);
nand U7514 (N_7514,N_5399,N_5423);
nand U7515 (N_7515,N_4676,N_4042);
and U7516 (N_7516,N_5663,N_4661);
nor U7517 (N_7517,N_4621,N_5617);
nand U7518 (N_7518,N_5136,N_5536);
xnor U7519 (N_7519,N_4455,N_5847);
nand U7520 (N_7520,N_5570,N_4811);
xor U7521 (N_7521,N_4273,N_4488);
nand U7522 (N_7522,N_5304,N_5775);
xor U7523 (N_7523,N_5941,N_4036);
or U7524 (N_7524,N_5865,N_5335);
nor U7525 (N_7525,N_4276,N_5120);
or U7526 (N_7526,N_5298,N_5992);
or U7527 (N_7527,N_5749,N_4573);
xor U7528 (N_7528,N_4777,N_4196);
xor U7529 (N_7529,N_4775,N_4342);
or U7530 (N_7530,N_5102,N_5672);
xnor U7531 (N_7531,N_5076,N_4777);
or U7532 (N_7532,N_4196,N_4028);
and U7533 (N_7533,N_4769,N_4494);
nor U7534 (N_7534,N_4775,N_5966);
xor U7535 (N_7535,N_5022,N_5680);
and U7536 (N_7536,N_4205,N_4436);
xnor U7537 (N_7537,N_4203,N_4178);
and U7538 (N_7538,N_5112,N_5812);
xor U7539 (N_7539,N_4189,N_4938);
nor U7540 (N_7540,N_5721,N_5551);
or U7541 (N_7541,N_4715,N_5111);
and U7542 (N_7542,N_5111,N_4127);
nor U7543 (N_7543,N_5048,N_4195);
nor U7544 (N_7544,N_5968,N_4368);
nor U7545 (N_7545,N_5796,N_4945);
nor U7546 (N_7546,N_4273,N_4797);
xnor U7547 (N_7547,N_5817,N_4836);
or U7548 (N_7548,N_5852,N_5167);
xor U7549 (N_7549,N_5292,N_5446);
or U7550 (N_7550,N_5978,N_4214);
or U7551 (N_7551,N_5417,N_4117);
or U7552 (N_7552,N_5197,N_5348);
xor U7553 (N_7553,N_4213,N_5644);
or U7554 (N_7554,N_4687,N_5361);
and U7555 (N_7555,N_5682,N_4110);
or U7556 (N_7556,N_4585,N_4726);
xnor U7557 (N_7557,N_4719,N_5617);
or U7558 (N_7558,N_4680,N_5455);
or U7559 (N_7559,N_5452,N_4300);
nand U7560 (N_7560,N_4654,N_4223);
and U7561 (N_7561,N_5017,N_5925);
nor U7562 (N_7562,N_4900,N_4354);
xnor U7563 (N_7563,N_4712,N_4757);
xor U7564 (N_7564,N_4983,N_4287);
and U7565 (N_7565,N_5322,N_4265);
nor U7566 (N_7566,N_5960,N_4247);
xnor U7567 (N_7567,N_4006,N_4908);
xor U7568 (N_7568,N_5820,N_4555);
and U7569 (N_7569,N_5189,N_4982);
nand U7570 (N_7570,N_4454,N_4474);
nand U7571 (N_7571,N_5809,N_5498);
and U7572 (N_7572,N_5942,N_4142);
nand U7573 (N_7573,N_4421,N_4581);
and U7574 (N_7574,N_5985,N_5911);
nand U7575 (N_7575,N_5883,N_5127);
nand U7576 (N_7576,N_5896,N_5480);
and U7577 (N_7577,N_4833,N_5422);
and U7578 (N_7578,N_5682,N_4589);
or U7579 (N_7579,N_4114,N_4318);
and U7580 (N_7580,N_5673,N_4728);
or U7581 (N_7581,N_4410,N_5558);
xor U7582 (N_7582,N_5413,N_5714);
nor U7583 (N_7583,N_5613,N_4315);
xnor U7584 (N_7584,N_4748,N_5794);
or U7585 (N_7585,N_4276,N_5493);
xnor U7586 (N_7586,N_5591,N_4500);
nand U7587 (N_7587,N_5411,N_5504);
nand U7588 (N_7588,N_4880,N_4191);
xor U7589 (N_7589,N_4946,N_5466);
nor U7590 (N_7590,N_5123,N_4283);
nand U7591 (N_7591,N_4404,N_5884);
xnor U7592 (N_7592,N_4948,N_4347);
and U7593 (N_7593,N_5423,N_4762);
or U7594 (N_7594,N_5710,N_4173);
or U7595 (N_7595,N_4097,N_4835);
xnor U7596 (N_7596,N_4671,N_5749);
and U7597 (N_7597,N_4687,N_4704);
nor U7598 (N_7598,N_4752,N_4858);
and U7599 (N_7599,N_5450,N_4391);
xnor U7600 (N_7600,N_5619,N_5939);
or U7601 (N_7601,N_5810,N_5110);
nand U7602 (N_7602,N_4782,N_4936);
or U7603 (N_7603,N_5195,N_4016);
nand U7604 (N_7604,N_5564,N_5343);
or U7605 (N_7605,N_5499,N_4090);
and U7606 (N_7606,N_4106,N_5351);
nand U7607 (N_7607,N_5893,N_4166);
or U7608 (N_7608,N_4122,N_5874);
or U7609 (N_7609,N_4684,N_4801);
and U7610 (N_7610,N_5597,N_4557);
and U7611 (N_7611,N_4033,N_5273);
nor U7612 (N_7612,N_4568,N_5867);
and U7613 (N_7613,N_5223,N_5170);
or U7614 (N_7614,N_4635,N_4283);
nand U7615 (N_7615,N_5909,N_4607);
and U7616 (N_7616,N_5626,N_5022);
nand U7617 (N_7617,N_5531,N_5119);
xnor U7618 (N_7618,N_5870,N_4349);
and U7619 (N_7619,N_4609,N_5303);
xor U7620 (N_7620,N_4266,N_4320);
and U7621 (N_7621,N_4115,N_5661);
nand U7622 (N_7622,N_5029,N_5108);
or U7623 (N_7623,N_5746,N_5832);
or U7624 (N_7624,N_4391,N_5629);
xnor U7625 (N_7625,N_4264,N_4784);
nor U7626 (N_7626,N_5673,N_4265);
or U7627 (N_7627,N_4779,N_4251);
xnor U7628 (N_7628,N_5582,N_4230);
or U7629 (N_7629,N_4985,N_4216);
xnor U7630 (N_7630,N_4168,N_5602);
and U7631 (N_7631,N_5540,N_4675);
or U7632 (N_7632,N_4887,N_4056);
nor U7633 (N_7633,N_5848,N_5367);
or U7634 (N_7634,N_5848,N_5363);
and U7635 (N_7635,N_4553,N_5857);
or U7636 (N_7636,N_5627,N_4158);
nor U7637 (N_7637,N_4237,N_5207);
nor U7638 (N_7638,N_4419,N_5118);
and U7639 (N_7639,N_5684,N_4728);
nand U7640 (N_7640,N_4798,N_5615);
nor U7641 (N_7641,N_5274,N_4531);
or U7642 (N_7642,N_5856,N_4901);
nor U7643 (N_7643,N_4910,N_4657);
nand U7644 (N_7644,N_4696,N_4798);
xnor U7645 (N_7645,N_4632,N_4127);
nand U7646 (N_7646,N_5209,N_5882);
nor U7647 (N_7647,N_5911,N_4857);
nand U7648 (N_7648,N_5327,N_4340);
xnor U7649 (N_7649,N_5541,N_5340);
and U7650 (N_7650,N_4564,N_5301);
or U7651 (N_7651,N_4272,N_4878);
or U7652 (N_7652,N_5651,N_4575);
xor U7653 (N_7653,N_4947,N_4528);
and U7654 (N_7654,N_4836,N_4130);
xor U7655 (N_7655,N_4365,N_5636);
and U7656 (N_7656,N_4481,N_5469);
and U7657 (N_7657,N_5796,N_4789);
nand U7658 (N_7658,N_4652,N_4934);
xor U7659 (N_7659,N_5365,N_4689);
or U7660 (N_7660,N_5408,N_4000);
nor U7661 (N_7661,N_4149,N_5091);
and U7662 (N_7662,N_5339,N_5023);
and U7663 (N_7663,N_4775,N_5175);
nand U7664 (N_7664,N_5632,N_4622);
nor U7665 (N_7665,N_4195,N_4482);
nand U7666 (N_7666,N_4925,N_5609);
nor U7667 (N_7667,N_5149,N_4609);
nor U7668 (N_7668,N_4687,N_5812);
or U7669 (N_7669,N_4380,N_5922);
or U7670 (N_7670,N_5602,N_5281);
or U7671 (N_7671,N_4871,N_4521);
or U7672 (N_7672,N_4401,N_4298);
or U7673 (N_7673,N_5120,N_4322);
xor U7674 (N_7674,N_4059,N_4158);
and U7675 (N_7675,N_5277,N_5715);
xor U7676 (N_7676,N_5037,N_5198);
nand U7677 (N_7677,N_4948,N_4483);
or U7678 (N_7678,N_5233,N_5364);
nor U7679 (N_7679,N_4155,N_4491);
nand U7680 (N_7680,N_4325,N_4110);
xnor U7681 (N_7681,N_5242,N_4277);
nand U7682 (N_7682,N_5647,N_5417);
nand U7683 (N_7683,N_5514,N_5058);
nand U7684 (N_7684,N_5425,N_4792);
xor U7685 (N_7685,N_4709,N_5625);
nand U7686 (N_7686,N_4590,N_4639);
nor U7687 (N_7687,N_4641,N_4043);
or U7688 (N_7688,N_5861,N_4511);
nand U7689 (N_7689,N_5172,N_4445);
or U7690 (N_7690,N_5210,N_5756);
and U7691 (N_7691,N_5499,N_5264);
or U7692 (N_7692,N_5619,N_5427);
nand U7693 (N_7693,N_4365,N_5096);
nand U7694 (N_7694,N_4973,N_4009);
and U7695 (N_7695,N_4620,N_4259);
and U7696 (N_7696,N_4294,N_5312);
xnor U7697 (N_7697,N_5759,N_4595);
nand U7698 (N_7698,N_5808,N_5293);
or U7699 (N_7699,N_4322,N_4247);
nand U7700 (N_7700,N_5126,N_4421);
and U7701 (N_7701,N_5182,N_5463);
nor U7702 (N_7702,N_5687,N_5974);
xor U7703 (N_7703,N_5415,N_5553);
nand U7704 (N_7704,N_5860,N_5431);
or U7705 (N_7705,N_4722,N_5652);
xor U7706 (N_7706,N_5277,N_5830);
nor U7707 (N_7707,N_5233,N_4348);
nand U7708 (N_7708,N_5519,N_5756);
nor U7709 (N_7709,N_4713,N_5920);
and U7710 (N_7710,N_5556,N_5033);
xnor U7711 (N_7711,N_4697,N_4159);
nand U7712 (N_7712,N_5404,N_5969);
and U7713 (N_7713,N_4875,N_4389);
and U7714 (N_7714,N_5258,N_4487);
and U7715 (N_7715,N_4217,N_5019);
and U7716 (N_7716,N_4131,N_4625);
and U7717 (N_7717,N_5353,N_5158);
nand U7718 (N_7718,N_5962,N_5984);
xor U7719 (N_7719,N_4278,N_4968);
nand U7720 (N_7720,N_4987,N_4244);
nor U7721 (N_7721,N_5267,N_5209);
and U7722 (N_7722,N_4888,N_5373);
or U7723 (N_7723,N_5198,N_5914);
and U7724 (N_7724,N_5079,N_4097);
nand U7725 (N_7725,N_4270,N_5927);
nor U7726 (N_7726,N_5592,N_4342);
or U7727 (N_7727,N_4702,N_4952);
or U7728 (N_7728,N_4434,N_4150);
nor U7729 (N_7729,N_5204,N_4243);
nor U7730 (N_7730,N_4111,N_4240);
or U7731 (N_7731,N_5175,N_5594);
nor U7732 (N_7732,N_5601,N_4615);
or U7733 (N_7733,N_5974,N_4433);
and U7734 (N_7734,N_4407,N_4214);
xnor U7735 (N_7735,N_5140,N_5411);
or U7736 (N_7736,N_4897,N_5578);
nor U7737 (N_7737,N_4869,N_5348);
nor U7738 (N_7738,N_5153,N_5544);
nand U7739 (N_7739,N_5473,N_4985);
and U7740 (N_7740,N_4882,N_4504);
or U7741 (N_7741,N_5061,N_4037);
xor U7742 (N_7742,N_5121,N_5965);
xor U7743 (N_7743,N_5200,N_5941);
nand U7744 (N_7744,N_4706,N_4742);
and U7745 (N_7745,N_4545,N_4995);
nand U7746 (N_7746,N_4421,N_4761);
xnor U7747 (N_7747,N_4845,N_5449);
or U7748 (N_7748,N_5199,N_4547);
xnor U7749 (N_7749,N_4590,N_5770);
and U7750 (N_7750,N_5729,N_4049);
or U7751 (N_7751,N_5076,N_4222);
or U7752 (N_7752,N_4240,N_4134);
nor U7753 (N_7753,N_4426,N_5554);
xor U7754 (N_7754,N_5445,N_5346);
nor U7755 (N_7755,N_5342,N_4700);
xor U7756 (N_7756,N_5284,N_5595);
xor U7757 (N_7757,N_5128,N_4959);
nor U7758 (N_7758,N_4064,N_5718);
xor U7759 (N_7759,N_5128,N_5335);
nand U7760 (N_7760,N_5997,N_5429);
nand U7761 (N_7761,N_5254,N_4726);
and U7762 (N_7762,N_5319,N_4704);
nor U7763 (N_7763,N_4004,N_4035);
nor U7764 (N_7764,N_4522,N_4889);
nand U7765 (N_7765,N_5203,N_4409);
xnor U7766 (N_7766,N_4647,N_4874);
or U7767 (N_7767,N_4491,N_5139);
nand U7768 (N_7768,N_4140,N_4778);
nand U7769 (N_7769,N_4063,N_5022);
nand U7770 (N_7770,N_5639,N_4930);
nand U7771 (N_7771,N_5178,N_5476);
or U7772 (N_7772,N_5763,N_5527);
xnor U7773 (N_7773,N_5928,N_4202);
nor U7774 (N_7774,N_5587,N_5960);
or U7775 (N_7775,N_4009,N_5381);
xnor U7776 (N_7776,N_5967,N_5244);
or U7777 (N_7777,N_4542,N_4541);
nor U7778 (N_7778,N_4716,N_5180);
or U7779 (N_7779,N_4865,N_4528);
and U7780 (N_7780,N_4759,N_4926);
nand U7781 (N_7781,N_4931,N_4006);
or U7782 (N_7782,N_5808,N_4761);
nor U7783 (N_7783,N_4397,N_4394);
xor U7784 (N_7784,N_4087,N_4241);
nand U7785 (N_7785,N_5933,N_4489);
nand U7786 (N_7786,N_5361,N_5334);
nand U7787 (N_7787,N_4587,N_4724);
and U7788 (N_7788,N_4967,N_4432);
or U7789 (N_7789,N_5237,N_4777);
or U7790 (N_7790,N_5593,N_4270);
and U7791 (N_7791,N_5679,N_5398);
nand U7792 (N_7792,N_4239,N_5006);
nand U7793 (N_7793,N_5987,N_5767);
or U7794 (N_7794,N_4202,N_4517);
and U7795 (N_7795,N_5914,N_4305);
and U7796 (N_7796,N_5793,N_5266);
nor U7797 (N_7797,N_5372,N_4328);
xnor U7798 (N_7798,N_5764,N_5523);
or U7799 (N_7799,N_5496,N_5680);
nand U7800 (N_7800,N_4996,N_5117);
or U7801 (N_7801,N_5396,N_5791);
and U7802 (N_7802,N_4226,N_4443);
and U7803 (N_7803,N_5375,N_5092);
nor U7804 (N_7804,N_4870,N_4214);
nor U7805 (N_7805,N_5248,N_4611);
xnor U7806 (N_7806,N_5700,N_4796);
and U7807 (N_7807,N_5421,N_4503);
and U7808 (N_7808,N_5708,N_5915);
or U7809 (N_7809,N_5762,N_4377);
nand U7810 (N_7810,N_4680,N_4197);
nor U7811 (N_7811,N_5382,N_4935);
nand U7812 (N_7812,N_5094,N_4110);
and U7813 (N_7813,N_5088,N_4440);
and U7814 (N_7814,N_4691,N_5728);
or U7815 (N_7815,N_5816,N_4712);
nor U7816 (N_7816,N_5495,N_4730);
and U7817 (N_7817,N_4928,N_5327);
or U7818 (N_7818,N_4083,N_4714);
nand U7819 (N_7819,N_5737,N_4683);
and U7820 (N_7820,N_5789,N_4716);
or U7821 (N_7821,N_5142,N_4478);
nand U7822 (N_7822,N_4344,N_5763);
and U7823 (N_7823,N_4079,N_4643);
nor U7824 (N_7824,N_4052,N_5477);
nand U7825 (N_7825,N_5303,N_4128);
xor U7826 (N_7826,N_5358,N_5956);
and U7827 (N_7827,N_5176,N_5890);
nand U7828 (N_7828,N_5187,N_4634);
and U7829 (N_7829,N_5458,N_4286);
or U7830 (N_7830,N_5628,N_4285);
nand U7831 (N_7831,N_4516,N_5335);
nand U7832 (N_7832,N_5272,N_5626);
nand U7833 (N_7833,N_4209,N_5676);
nor U7834 (N_7834,N_4988,N_5015);
or U7835 (N_7835,N_4496,N_4276);
or U7836 (N_7836,N_4885,N_4606);
and U7837 (N_7837,N_4409,N_4521);
nand U7838 (N_7838,N_4715,N_5918);
and U7839 (N_7839,N_5379,N_4882);
or U7840 (N_7840,N_5747,N_5743);
xnor U7841 (N_7841,N_5467,N_4851);
nand U7842 (N_7842,N_4252,N_5665);
or U7843 (N_7843,N_4389,N_4328);
nand U7844 (N_7844,N_5380,N_4421);
nand U7845 (N_7845,N_5146,N_4816);
or U7846 (N_7846,N_4782,N_4736);
or U7847 (N_7847,N_5184,N_5427);
or U7848 (N_7848,N_4323,N_5293);
nand U7849 (N_7849,N_4877,N_5162);
and U7850 (N_7850,N_4268,N_5302);
or U7851 (N_7851,N_4841,N_5889);
nand U7852 (N_7852,N_5693,N_4372);
and U7853 (N_7853,N_4365,N_5301);
xnor U7854 (N_7854,N_5720,N_4226);
and U7855 (N_7855,N_5367,N_5720);
nand U7856 (N_7856,N_4810,N_5793);
or U7857 (N_7857,N_4966,N_5109);
nor U7858 (N_7858,N_5563,N_4967);
and U7859 (N_7859,N_4423,N_4275);
xnor U7860 (N_7860,N_5274,N_5642);
and U7861 (N_7861,N_5929,N_5392);
nor U7862 (N_7862,N_4647,N_4226);
or U7863 (N_7863,N_4781,N_4764);
nand U7864 (N_7864,N_5112,N_4741);
nor U7865 (N_7865,N_4478,N_5374);
or U7866 (N_7866,N_4884,N_4642);
nor U7867 (N_7867,N_4247,N_5910);
nand U7868 (N_7868,N_5243,N_5465);
nor U7869 (N_7869,N_5880,N_5255);
nor U7870 (N_7870,N_5289,N_5493);
nor U7871 (N_7871,N_4890,N_4122);
nor U7872 (N_7872,N_5528,N_4297);
nand U7873 (N_7873,N_5084,N_4583);
nand U7874 (N_7874,N_5146,N_4863);
or U7875 (N_7875,N_4982,N_4555);
nor U7876 (N_7876,N_5729,N_5924);
xnor U7877 (N_7877,N_5028,N_5057);
nand U7878 (N_7878,N_4927,N_4977);
nand U7879 (N_7879,N_4421,N_5695);
or U7880 (N_7880,N_5480,N_5429);
xnor U7881 (N_7881,N_4137,N_4622);
xnor U7882 (N_7882,N_5376,N_5989);
xor U7883 (N_7883,N_4155,N_4023);
nand U7884 (N_7884,N_5768,N_5363);
and U7885 (N_7885,N_5019,N_4416);
xor U7886 (N_7886,N_5880,N_4249);
or U7887 (N_7887,N_4593,N_4590);
xor U7888 (N_7888,N_4409,N_5111);
and U7889 (N_7889,N_5630,N_4450);
and U7890 (N_7890,N_5562,N_5098);
or U7891 (N_7891,N_4063,N_4985);
or U7892 (N_7892,N_4060,N_4727);
nand U7893 (N_7893,N_4700,N_4818);
and U7894 (N_7894,N_5610,N_4951);
nor U7895 (N_7895,N_5777,N_5952);
nand U7896 (N_7896,N_5999,N_4753);
nor U7897 (N_7897,N_5671,N_4791);
xnor U7898 (N_7898,N_5702,N_4317);
xnor U7899 (N_7899,N_4142,N_5381);
nand U7900 (N_7900,N_4989,N_4525);
nor U7901 (N_7901,N_4853,N_4546);
nor U7902 (N_7902,N_5011,N_4133);
xor U7903 (N_7903,N_5068,N_4435);
nor U7904 (N_7904,N_5739,N_4112);
nor U7905 (N_7905,N_4589,N_4456);
nand U7906 (N_7906,N_4928,N_4196);
or U7907 (N_7907,N_4672,N_5012);
nand U7908 (N_7908,N_4816,N_5246);
xor U7909 (N_7909,N_5582,N_5693);
nand U7910 (N_7910,N_5190,N_4395);
and U7911 (N_7911,N_5684,N_5284);
nor U7912 (N_7912,N_5363,N_5825);
nor U7913 (N_7913,N_5632,N_5787);
nor U7914 (N_7914,N_5728,N_5234);
nor U7915 (N_7915,N_4225,N_4625);
and U7916 (N_7916,N_4118,N_5691);
nor U7917 (N_7917,N_4732,N_4064);
or U7918 (N_7918,N_5632,N_5275);
nand U7919 (N_7919,N_4943,N_4905);
nand U7920 (N_7920,N_4666,N_4768);
and U7921 (N_7921,N_4339,N_5422);
xor U7922 (N_7922,N_5902,N_5612);
nand U7923 (N_7923,N_4089,N_4894);
nor U7924 (N_7924,N_5905,N_5561);
nor U7925 (N_7925,N_4689,N_5627);
nor U7926 (N_7926,N_4826,N_5340);
xnor U7927 (N_7927,N_4363,N_5693);
or U7928 (N_7928,N_5008,N_4703);
nand U7929 (N_7929,N_4418,N_5519);
or U7930 (N_7930,N_5306,N_4802);
xnor U7931 (N_7931,N_4786,N_5378);
or U7932 (N_7932,N_4425,N_5073);
xor U7933 (N_7933,N_4242,N_4879);
and U7934 (N_7934,N_5497,N_4826);
xor U7935 (N_7935,N_4586,N_5795);
and U7936 (N_7936,N_4040,N_5607);
or U7937 (N_7937,N_4813,N_4946);
or U7938 (N_7938,N_4621,N_4006);
nand U7939 (N_7939,N_4488,N_4465);
xor U7940 (N_7940,N_4634,N_5490);
nand U7941 (N_7941,N_5747,N_4392);
nor U7942 (N_7942,N_5540,N_5472);
nand U7943 (N_7943,N_5845,N_5203);
nand U7944 (N_7944,N_4262,N_4116);
or U7945 (N_7945,N_5026,N_4086);
xor U7946 (N_7946,N_4519,N_4562);
nor U7947 (N_7947,N_4424,N_5345);
or U7948 (N_7948,N_5119,N_4698);
nor U7949 (N_7949,N_4078,N_4907);
and U7950 (N_7950,N_4751,N_5103);
nand U7951 (N_7951,N_4437,N_5993);
nand U7952 (N_7952,N_5609,N_5616);
and U7953 (N_7953,N_4713,N_4189);
nor U7954 (N_7954,N_4229,N_5652);
and U7955 (N_7955,N_5093,N_5400);
and U7956 (N_7956,N_5201,N_5819);
and U7957 (N_7957,N_5112,N_4739);
nor U7958 (N_7958,N_4193,N_4502);
and U7959 (N_7959,N_4642,N_4173);
and U7960 (N_7960,N_4564,N_4512);
nor U7961 (N_7961,N_4937,N_5135);
nand U7962 (N_7962,N_4333,N_5175);
and U7963 (N_7963,N_4201,N_5580);
nor U7964 (N_7964,N_5128,N_5801);
nor U7965 (N_7965,N_4163,N_5790);
and U7966 (N_7966,N_4400,N_4661);
nor U7967 (N_7967,N_4124,N_5496);
xor U7968 (N_7968,N_5180,N_4398);
nor U7969 (N_7969,N_5814,N_4462);
nand U7970 (N_7970,N_4451,N_5047);
nand U7971 (N_7971,N_5618,N_4405);
and U7972 (N_7972,N_5850,N_5523);
and U7973 (N_7973,N_4080,N_4646);
nor U7974 (N_7974,N_4118,N_4890);
and U7975 (N_7975,N_5818,N_5085);
nand U7976 (N_7976,N_4206,N_4789);
nand U7977 (N_7977,N_4989,N_5747);
nor U7978 (N_7978,N_5683,N_4205);
nand U7979 (N_7979,N_5153,N_5899);
nand U7980 (N_7980,N_5671,N_5736);
or U7981 (N_7981,N_4637,N_4257);
nor U7982 (N_7982,N_5874,N_5480);
and U7983 (N_7983,N_5025,N_4931);
nand U7984 (N_7984,N_4282,N_4326);
or U7985 (N_7985,N_4113,N_5839);
nand U7986 (N_7986,N_4452,N_4424);
or U7987 (N_7987,N_4549,N_4680);
xnor U7988 (N_7988,N_5279,N_4528);
and U7989 (N_7989,N_5736,N_4603);
or U7990 (N_7990,N_5218,N_4515);
and U7991 (N_7991,N_4648,N_4224);
or U7992 (N_7992,N_4820,N_4409);
xnor U7993 (N_7993,N_4385,N_4624);
nand U7994 (N_7994,N_5193,N_5660);
or U7995 (N_7995,N_5467,N_5056);
xnor U7996 (N_7996,N_5335,N_4222);
xnor U7997 (N_7997,N_5511,N_5885);
nand U7998 (N_7998,N_4167,N_4638);
or U7999 (N_7999,N_4810,N_5517);
nand U8000 (N_8000,N_7463,N_6527);
xor U8001 (N_8001,N_6601,N_6460);
and U8002 (N_8002,N_6818,N_7087);
or U8003 (N_8003,N_6064,N_6716);
xnor U8004 (N_8004,N_7172,N_7183);
nand U8005 (N_8005,N_7438,N_6636);
xor U8006 (N_8006,N_7304,N_7103);
or U8007 (N_8007,N_7575,N_7765);
nand U8008 (N_8008,N_7232,N_6234);
and U8009 (N_8009,N_6967,N_6642);
nor U8010 (N_8010,N_6614,N_6522);
and U8011 (N_8011,N_6715,N_6302);
xnor U8012 (N_8012,N_6795,N_7699);
nor U8013 (N_8013,N_6362,N_6754);
and U8014 (N_8014,N_6127,N_6272);
or U8015 (N_8015,N_7506,N_6609);
nand U8016 (N_8016,N_7863,N_6156);
or U8017 (N_8017,N_7142,N_6870);
nor U8018 (N_8018,N_6359,N_6215);
or U8019 (N_8019,N_7202,N_6864);
and U8020 (N_8020,N_7356,N_6993);
xnor U8021 (N_8021,N_7160,N_6843);
xor U8022 (N_8022,N_7567,N_7195);
nor U8023 (N_8023,N_7889,N_6520);
and U8024 (N_8024,N_7828,N_6361);
or U8025 (N_8025,N_6893,N_7585);
nand U8026 (N_8026,N_7021,N_6277);
nand U8027 (N_8027,N_7564,N_7061);
nor U8028 (N_8028,N_7657,N_7668);
nand U8029 (N_8029,N_7239,N_6348);
and U8030 (N_8030,N_6825,N_7154);
and U8031 (N_8031,N_7445,N_6972);
nor U8032 (N_8032,N_6821,N_7084);
nor U8033 (N_8033,N_6612,N_6856);
and U8034 (N_8034,N_6559,N_6743);
nand U8035 (N_8035,N_7827,N_7462);
or U8036 (N_8036,N_7578,N_7891);
or U8037 (N_8037,N_7342,N_6546);
nand U8038 (N_8038,N_7804,N_7783);
nand U8039 (N_8039,N_7032,N_6652);
xnor U8040 (N_8040,N_6851,N_7034);
nor U8041 (N_8041,N_7182,N_7734);
and U8042 (N_8042,N_7710,N_6790);
nor U8043 (N_8043,N_6845,N_7843);
and U8044 (N_8044,N_7684,N_6093);
nand U8045 (N_8045,N_7265,N_6447);
nand U8046 (N_8046,N_7079,N_6747);
or U8047 (N_8047,N_7313,N_6134);
nor U8048 (N_8048,N_6245,N_6229);
xnor U8049 (N_8049,N_7042,N_7259);
xor U8050 (N_8050,N_6074,N_7784);
xor U8051 (N_8051,N_6943,N_6310);
xor U8052 (N_8052,N_6816,N_7483);
or U8053 (N_8053,N_6668,N_6043);
xnor U8054 (N_8054,N_6321,N_7416);
xnor U8055 (N_8055,N_7256,N_7294);
and U8056 (N_8056,N_7028,N_6633);
nor U8057 (N_8057,N_7701,N_6945);
nor U8058 (N_8058,N_6985,N_7129);
or U8059 (N_8059,N_7543,N_6583);
or U8060 (N_8060,N_6429,N_6305);
or U8061 (N_8061,N_6564,N_6296);
xor U8062 (N_8062,N_7855,N_7215);
or U8063 (N_8063,N_7562,N_6330);
and U8064 (N_8064,N_6751,N_7628);
nor U8065 (N_8065,N_7059,N_6102);
nor U8066 (N_8066,N_7029,N_7662);
nor U8067 (N_8067,N_6646,N_7568);
and U8068 (N_8068,N_6473,N_6530);
nor U8069 (N_8069,N_7083,N_7224);
nand U8070 (N_8070,N_7437,N_6617);
or U8071 (N_8071,N_7381,N_6112);
nor U8072 (N_8072,N_6406,N_6086);
nor U8073 (N_8073,N_6647,N_6107);
nand U8074 (N_8074,N_7524,N_7885);
or U8075 (N_8075,N_6414,N_7989);
nand U8076 (N_8076,N_6045,N_7108);
or U8077 (N_8077,N_7890,N_7687);
and U8078 (N_8078,N_6078,N_7307);
xnor U8079 (N_8079,N_6718,N_7951);
xnor U8080 (N_8080,N_7821,N_7328);
and U8081 (N_8081,N_6929,N_7364);
xor U8082 (N_8082,N_7507,N_7935);
or U8083 (N_8083,N_6641,N_7286);
xnor U8084 (N_8084,N_6576,N_7249);
or U8085 (N_8085,N_6260,N_6920);
or U8086 (N_8086,N_6542,N_7163);
or U8087 (N_8087,N_6944,N_7162);
nor U8088 (N_8088,N_7577,N_6509);
xor U8089 (N_8089,N_7143,N_6243);
xor U8090 (N_8090,N_6360,N_7547);
xnor U8091 (N_8091,N_6340,N_7064);
nor U8092 (N_8092,N_7276,N_7205);
or U8093 (N_8093,N_6145,N_6511);
nand U8094 (N_8094,N_6565,N_6407);
and U8095 (N_8095,N_7428,N_7902);
nand U8096 (N_8096,N_7869,N_6080);
or U8097 (N_8097,N_6274,N_6595);
nor U8098 (N_8098,N_7382,N_7925);
or U8099 (N_8099,N_7988,N_6336);
and U8100 (N_8100,N_6136,N_7361);
and U8101 (N_8101,N_7823,N_7983);
or U8102 (N_8102,N_7515,N_7231);
and U8103 (N_8103,N_7636,N_6173);
nand U8104 (N_8104,N_7112,N_7489);
or U8105 (N_8105,N_7487,N_7597);
nand U8106 (N_8106,N_6817,N_6772);
xnor U8107 (N_8107,N_6143,N_7478);
xor U8108 (N_8108,N_7895,N_7611);
and U8109 (N_8109,N_7803,N_6218);
and U8110 (N_8110,N_6714,N_7786);
and U8111 (N_8111,N_6819,N_7053);
or U8112 (N_8112,N_7810,N_7472);
xor U8113 (N_8113,N_6704,N_6670);
and U8114 (N_8114,N_7390,N_6581);
or U8115 (N_8115,N_7167,N_6717);
or U8116 (N_8116,N_7475,N_7702);
nor U8117 (N_8117,N_7363,N_7082);
or U8118 (N_8118,N_6413,N_6886);
nand U8119 (N_8119,N_6002,N_7229);
nand U8120 (N_8120,N_7090,N_6486);
nand U8121 (N_8121,N_6988,N_6535);
nor U8122 (N_8122,N_7967,N_6536);
nor U8123 (N_8123,N_6664,N_6109);
nor U8124 (N_8124,N_7102,N_7466);
and U8125 (N_8125,N_6774,N_6677);
or U8126 (N_8126,N_6344,N_7186);
nor U8127 (N_8127,N_6586,N_6961);
and U8128 (N_8128,N_7697,N_6177);
or U8129 (N_8129,N_6587,N_6400);
nand U8130 (N_8130,N_6734,N_6651);
nor U8131 (N_8131,N_6608,N_6162);
xor U8132 (N_8132,N_6915,N_7368);
xnor U8133 (N_8133,N_6557,N_7496);
xnor U8134 (N_8134,N_6912,N_7589);
or U8135 (N_8135,N_7455,N_6659);
nor U8136 (N_8136,N_7754,N_7764);
nand U8137 (N_8137,N_6242,N_7576);
xnor U8138 (N_8138,N_6553,N_6802);
and U8139 (N_8139,N_7958,N_6853);
xnor U8140 (N_8140,N_7171,N_6062);
xnor U8141 (N_8141,N_7728,N_7852);
xor U8142 (N_8142,N_6901,N_6213);
xnor U8143 (N_8143,N_7711,N_6973);
or U8144 (N_8144,N_6866,N_6957);
or U8145 (N_8145,N_7759,N_7086);
nand U8146 (N_8146,N_6240,N_7779);
or U8147 (N_8147,N_7196,N_6063);
nand U8148 (N_8148,N_7188,N_7962);
and U8149 (N_8149,N_6026,N_7288);
nor U8150 (N_8150,N_6733,N_7264);
and U8151 (N_8151,N_6159,N_6066);
or U8152 (N_8152,N_6591,N_7114);
xnor U8153 (N_8153,N_6499,N_6932);
and U8154 (N_8154,N_6327,N_6692);
nor U8155 (N_8155,N_7631,N_6847);
nor U8156 (N_8156,N_6322,N_7877);
and U8157 (N_8157,N_6448,N_7647);
xor U8158 (N_8158,N_6709,N_6053);
xor U8159 (N_8159,N_6590,N_7801);
xnor U8160 (N_8160,N_7473,N_7533);
xor U8161 (N_8161,N_6374,N_7400);
or U8162 (N_8162,N_7070,N_7203);
or U8163 (N_8163,N_7847,N_6738);
xor U8164 (N_8164,N_6534,N_7144);
xnor U8165 (N_8165,N_7471,N_7436);
nand U8166 (N_8166,N_6696,N_6404);
nor U8167 (N_8167,N_6169,N_7388);
or U8168 (N_8168,N_7310,N_6742);
nand U8169 (N_8169,N_7035,N_6706);
xnor U8170 (N_8170,N_7905,N_7351);
xnor U8171 (N_8171,N_6098,N_6428);
nand U8172 (N_8172,N_7778,N_6294);
nor U8173 (N_8173,N_6631,N_7777);
xor U8174 (N_8174,N_6637,N_7815);
or U8175 (N_8175,N_7862,N_6962);
nor U8176 (N_8176,N_6380,N_7133);
xnor U8177 (N_8177,N_7594,N_7049);
xnor U8178 (N_8178,N_7817,N_7124);
nand U8179 (N_8179,N_7442,N_6955);
nand U8180 (N_8180,N_7460,N_7494);
nor U8181 (N_8181,N_7329,N_7066);
and U8182 (N_8182,N_7833,N_6172);
nor U8183 (N_8183,N_6402,N_6625);
nor U8184 (N_8184,N_6269,N_6011);
nor U8185 (N_8185,N_7691,N_6487);
xnor U8186 (N_8186,N_7319,N_6057);
or U8187 (N_8187,N_6914,N_6120);
xor U8188 (N_8188,N_6480,N_7528);
xor U8189 (N_8189,N_6088,N_7345);
and U8190 (N_8190,N_7200,N_7639);
nand U8191 (N_8191,N_7943,N_7347);
and U8192 (N_8192,N_7624,N_6390);
and U8193 (N_8193,N_6775,N_7399);
and U8194 (N_8194,N_7263,N_6827);
nand U8195 (N_8195,N_7016,N_7924);
nand U8196 (N_8196,N_6190,N_7735);
and U8197 (N_8197,N_7956,N_7337);
xnor U8198 (N_8198,N_7099,N_6259);
or U8199 (N_8199,N_7403,N_7137);
xor U8200 (N_8200,N_6019,N_7839);
nor U8201 (N_8201,N_6574,N_6090);
nor U8202 (N_8202,N_7175,N_6351);
nor U8203 (N_8203,N_7806,N_6323);
or U8204 (N_8204,N_7616,N_6975);
and U8205 (N_8205,N_7671,N_6698);
xor U8206 (N_8206,N_7015,N_6283);
nand U8207 (N_8207,N_6672,N_7731);
xor U8208 (N_8208,N_7548,N_7014);
and U8209 (N_8209,N_7860,N_7796);
or U8210 (N_8210,N_7527,N_7355);
nor U8211 (N_8211,N_6861,N_6219);
xnor U8212 (N_8212,N_6433,N_6051);
or U8213 (N_8213,N_6965,N_7377);
nor U8214 (N_8214,N_7749,N_6308);
and U8215 (N_8215,N_6452,N_6178);
nor U8216 (N_8216,N_7257,N_6036);
nor U8217 (N_8217,N_6999,N_7703);
nor U8218 (N_8218,N_7914,N_6976);
nand U8219 (N_8219,N_7882,N_6235);
nor U8220 (N_8220,N_7375,N_7880);
nand U8221 (N_8221,N_6504,N_7295);
and U8222 (N_8222,N_7788,N_6158);
xnor U8223 (N_8223,N_7246,N_7170);
xor U8224 (N_8224,N_7676,N_6075);
nand U8225 (N_8225,N_7430,N_6300);
and U8226 (N_8226,N_6376,N_6194);
and U8227 (N_8227,N_7004,N_7707);
nor U8228 (N_8228,N_6065,N_6547);
or U8229 (N_8229,N_6524,N_6179);
nand U8230 (N_8230,N_7739,N_7094);
and U8231 (N_8231,N_6490,N_6092);
xnor U8232 (N_8232,N_6889,N_6757);
and U8233 (N_8233,N_6436,N_6118);
xor U8234 (N_8234,N_6140,N_7227);
and U8235 (N_8235,N_7467,N_6657);
nor U8236 (N_8236,N_7767,N_6822);
or U8237 (N_8237,N_6262,N_6475);
and U8238 (N_8238,N_7682,N_6784);
nor U8239 (N_8239,N_7758,N_6408);
or U8240 (N_8240,N_7516,N_7179);
nand U8241 (N_8241,N_7746,N_6928);
nor U8242 (N_8242,N_6110,N_6027);
xor U8243 (N_8243,N_6111,N_7736);
or U8244 (N_8244,N_7720,N_6862);
or U8245 (N_8245,N_6898,N_6899);
xnor U8246 (N_8246,N_6377,N_7262);
nor U8247 (N_8247,N_7291,N_6076);
xor U8248 (N_8248,N_7787,N_6632);
nor U8249 (N_8249,N_6255,N_7352);
and U8250 (N_8250,N_7406,N_7324);
or U8251 (N_8251,N_7601,N_6220);
nor U8252 (N_8252,N_7492,N_7942);
and U8253 (N_8253,N_7194,N_7448);
nand U8254 (N_8254,N_7374,N_6268);
nor U8255 (N_8255,N_6188,N_7602);
xor U8256 (N_8256,N_7518,N_6001);
and U8257 (N_8257,N_7125,N_6653);
or U8258 (N_8258,N_7113,N_7394);
nor U8259 (N_8259,N_7861,N_7539);
or U8260 (N_8260,N_7561,N_7260);
xor U8261 (N_8261,N_7348,N_6326);
nand U8262 (N_8262,N_7447,N_7148);
or U8263 (N_8263,N_6951,N_6459);
nor U8264 (N_8264,N_7119,N_6554);
nor U8265 (N_8265,N_6378,N_7376);
and U8266 (N_8266,N_7772,N_6033);
nand U8267 (N_8267,N_7479,N_7780);
xor U8268 (N_8268,N_6411,N_6163);
and U8269 (N_8269,N_7680,N_7721);
nand U8270 (N_8270,N_7449,N_7782);
and U8271 (N_8271,N_7752,N_7669);
nand U8272 (N_8272,N_7807,N_7285);
xnor U8273 (N_8273,N_6728,N_7234);
nand U8274 (N_8274,N_6116,N_7809);
nand U8275 (N_8275,N_7012,N_6050);
nand U8276 (N_8276,N_6538,N_7723);
or U8277 (N_8277,N_7106,N_7454);
and U8278 (N_8278,N_7373,N_6598);
nand U8279 (N_8279,N_7921,N_6656);
nor U8280 (N_8280,N_7615,N_7587);
or U8281 (N_8281,N_7916,N_7681);
and U8282 (N_8282,N_6471,N_6798);
nor U8283 (N_8283,N_7730,N_6675);
nor U8284 (N_8284,N_6989,N_6902);
and U8285 (N_8285,N_6338,N_6548);
and U8286 (N_8286,N_6419,N_6839);
nand U8287 (N_8287,N_7440,N_6426);
nor U8288 (N_8288,N_7834,N_6275);
nor U8289 (N_8289,N_6373,N_7679);
nor U8290 (N_8290,N_7063,N_6510);
nand U8291 (N_8291,N_6834,N_6729);
nor U8292 (N_8292,N_6750,N_6479);
xor U8293 (N_8293,N_6732,N_7534);
nor U8294 (N_8294,N_7453,N_6358);
nor U8295 (N_8295,N_6228,N_6895);
xnor U8296 (N_8296,N_6320,N_7490);
nand U8297 (N_8297,N_6405,N_7894);
and U8298 (N_8298,N_6369,N_7424);
xor U8299 (N_8299,N_7903,N_6872);
nand U8300 (N_8300,N_6122,N_7683);
nand U8301 (N_8301,N_7837,N_6777);
nand U8302 (N_8302,N_7936,N_6684);
nor U8303 (N_8303,N_6104,N_6683);
nand U8304 (N_8304,N_6037,N_6152);
xor U8305 (N_8305,N_6392,N_6236);
nor U8306 (N_8306,N_7851,N_7505);
nand U8307 (N_8307,N_6131,N_7140);
or U8308 (N_8308,N_7825,N_7972);
or U8309 (N_8309,N_6410,N_6840);
and U8310 (N_8310,N_6629,N_6495);
nand U8311 (N_8311,N_6648,N_6942);
xor U8312 (N_8312,N_6556,N_7708);
nor U8313 (N_8313,N_7901,N_6804);
nor U8314 (N_8314,N_7098,N_6996);
xor U8315 (N_8315,N_7592,N_6135);
nand U8316 (N_8316,N_7230,N_7135);
xnor U8317 (N_8317,N_7426,N_6301);
xnor U8318 (N_8318,N_7692,N_7411);
and U8319 (N_8319,N_7621,N_6040);
and U8320 (N_8320,N_6254,N_7198);
or U8321 (N_8321,N_6008,N_7514);
nand U8322 (N_8322,N_7405,N_6313);
or U8323 (N_8323,N_7009,N_6755);
nor U8324 (N_8324,N_6599,N_6029);
nor U8325 (N_8325,N_6289,N_6950);
or U8326 (N_8326,N_7044,N_7940);
nor U8327 (N_8327,N_6261,N_7010);
and U8328 (N_8328,N_7159,N_7927);
or U8329 (N_8329,N_6437,N_6981);
or U8330 (N_8330,N_6329,N_6991);
xor U8331 (N_8331,N_6139,N_7820);
and U8332 (N_8332,N_6298,N_6966);
and U8333 (N_8333,N_7068,N_7147);
xnor U8334 (N_8334,N_6690,N_6420);
and U8335 (N_8335,N_7867,N_7946);
nor U8336 (N_8336,N_6334,N_7218);
nand U8337 (N_8337,N_7836,N_6785);
or U8338 (N_8338,N_6153,N_6174);
xnor U8339 (N_8339,N_6431,N_6890);
nor U8340 (N_8340,N_6532,N_6248);
nand U8341 (N_8341,N_6195,N_6384);
nand U8342 (N_8342,N_7495,N_7253);
or U8343 (N_8343,N_6911,N_7209);
nor U8344 (N_8344,N_7718,N_6211);
nor U8345 (N_8345,N_6503,N_6505);
and U8346 (N_8346,N_7091,N_7864);
and U8347 (N_8347,N_7664,N_6891);
xnor U8348 (N_8348,N_6708,N_6610);
or U8349 (N_8349,N_7488,N_7630);
nor U8350 (N_8350,N_6852,N_6666);
and U8351 (N_8351,N_7733,N_6894);
nand U8352 (N_8352,N_6166,N_6282);
xnor U8353 (N_8353,N_7164,N_7663);
xor U8354 (N_8354,N_6842,N_7358);
xnor U8355 (N_8355,N_6563,N_6284);
or U8356 (N_8356,N_6149,N_7856);
xor U8357 (N_8357,N_6725,N_7873);
nand U8358 (N_8358,N_7419,N_6058);
or U8359 (N_8359,N_6416,N_7994);
nand U8360 (N_8360,N_7922,N_7565);
nor U8361 (N_8361,N_7959,N_7075);
xnor U8362 (N_8362,N_6549,N_6031);
or U8363 (N_8363,N_6693,N_7722);
and U8364 (N_8364,N_6626,N_6206);
and U8365 (N_8365,N_6462,N_6316);
or U8366 (N_8366,N_7503,N_6909);
nor U8367 (N_8367,N_6737,N_7579);
or U8368 (N_8368,N_6225,N_6645);
or U8369 (N_8369,N_6982,N_6810);
xnor U8370 (N_8370,N_6567,N_6721);
nor U8371 (N_8371,N_6119,N_7023);
nand U8372 (N_8372,N_6175,N_6458);
and U8373 (N_8373,N_7608,N_7580);
and U8374 (N_8374,N_7391,N_6917);
nand U8375 (N_8375,N_6994,N_7926);
nand U8376 (N_8376,N_6746,N_7333);
nand U8377 (N_8377,N_6465,N_6702);
nand U8378 (N_8378,N_7677,N_7913);
nand U8379 (N_8379,N_7327,N_6669);
nor U8380 (N_8380,N_6874,N_7939);
xnor U8381 (N_8381,N_6766,N_7367);
nand U8382 (N_8382,N_7627,N_6056);
xor U8383 (N_8383,N_6435,N_6309);
nand U8384 (N_8384,N_7790,N_6214);
or U8385 (N_8385,N_7635,N_6028);
xor U8386 (N_8386,N_6468,N_6687);
or U8387 (N_8387,N_7439,N_7963);
nor U8388 (N_8388,N_7210,N_6787);
or U8389 (N_8389,N_7957,N_7665);
and U8390 (N_8390,N_7997,N_7974);
nand U8391 (N_8391,N_7251,N_6180);
xnor U8392 (N_8392,N_6256,N_6295);
nor U8393 (N_8393,N_6061,N_7446);
and U8394 (N_8394,N_7252,N_7293);
or U8395 (N_8395,N_6748,N_6009);
nand U8396 (N_8396,N_6425,N_7541);
and U8397 (N_8397,N_6165,N_6497);
or U8398 (N_8398,N_6386,N_7623);
and U8399 (N_8399,N_7415,N_6793);
nand U8400 (N_8400,N_6528,N_7222);
and U8401 (N_8401,N_6231,N_7769);
nor U8402 (N_8402,N_7225,N_7953);
nor U8403 (N_8403,N_7305,N_7686);
xor U8404 (N_8404,N_7871,N_7629);
nor U8405 (N_8405,N_6032,N_6589);
nor U8406 (N_8406,N_7444,N_6808);
or U8407 (N_8407,N_6394,N_6346);
and U8408 (N_8408,N_6603,N_7551);
xor U8409 (N_8409,N_6201,N_6555);
xor U8410 (N_8410,N_7214,N_7798);
or U8411 (N_8411,N_7158,N_7341);
and U8412 (N_8412,N_6830,N_7584);
nand U8413 (N_8413,N_6811,N_7556);
nand U8414 (N_8414,N_7413,N_7526);
nand U8415 (N_8415,N_6939,N_7174);
nor U8416 (N_8416,N_7987,N_6141);
nand U8417 (N_8417,N_6446,N_7477);
nand U8418 (N_8418,N_7981,N_6125);
nand U8419 (N_8419,N_6807,N_7191);
nor U8420 (N_8420,N_7385,N_6079);
xor U8421 (N_8421,N_7278,N_7641);
and U8422 (N_8422,N_6686,N_6695);
or U8423 (N_8423,N_6541,N_7155);
and U8424 (N_8424,N_6780,N_6740);
xnor U8425 (N_8425,N_7724,N_6919);
nand U8426 (N_8426,N_7985,N_7971);
xnor U8427 (N_8427,N_6726,N_6389);
nand U8428 (N_8428,N_7149,N_7714);
nand U8429 (N_8429,N_7868,N_7052);
and U8430 (N_8430,N_7650,N_6654);
nand U8431 (N_8431,N_7386,N_7993);
and U8432 (N_8432,N_6551,N_7845);
nor U8433 (N_8433,N_6263,N_6154);
nand U8434 (N_8434,N_7306,N_6759);
or U8435 (N_8435,N_6467,N_6638);
xnor U8436 (N_8436,N_7990,N_6117);
or U8437 (N_8437,N_7934,N_7984);
xnor U8438 (N_8438,N_7168,N_6860);
nor U8439 (N_8439,N_6393,N_7673);
or U8440 (N_8440,N_6455,N_7811);
and U8441 (N_8441,N_7693,N_7619);
and U8442 (N_8442,N_7982,N_6339);
xor U8443 (N_8443,N_7027,N_6786);
nand U8444 (N_8444,N_7509,N_6478);
and U8445 (N_8445,N_7950,N_7212);
nor U8446 (N_8446,N_6570,N_7139);
or U8447 (N_8447,N_6496,N_6849);
or U8448 (N_8448,N_7018,N_7713);
and U8449 (N_8449,N_6266,N_6004);
nand U8450 (N_8450,N_7977,N_6935);
xor U8451 (N_8451,N_6771,N_6735);
or U8452 (N_8452,N_7634,N_7604);
and U8453 (N_8453,N_6508,N_7092);
nand U8454 (N_8454,N_6445,N_6903);
or U8455 (N_8455,N_6727,N_6372);
nand U8456 (N_8456,N_6343,N_7331);
and U8457 (N_8457,N_7250,N_6332);
or U8458 (N_8458,N_6068,N_6665);
and U8459 (N_8459,N_7464,N_7300);
and U8460 (N_8460,N_6015,N_6189);
xor U8461 (N_8461,N_6987,N_7241);
and U8462 (N_8462,N_6192,N_6723);
or U8463 (N_8463,N_7076,N_7336);
xnor U8464 (N_8464,N_7132,N_6267);
or U8465 (N_8465,N_7614,N_7161);
xor U8466 (N_8466,N_7540,N_6366);
or U8467 (N_8467,N_7870,N_6789);
and U8468 (N_8468,N_7923,N_6515);
and U8469 (N_8469,N_7056,N_7316);
xor U8470 (N_8470,N_7392,N_7435);
or U8471 (N_8471,N_6409,N_7706);
and U8472 (N_8472,N_7525,N_6682);
xnor U8473 (N_8473,N_6203,N_7109);
and U8474 (N_8474,N_7674,N_6863);
nand U8475 (N_8475,N_7932,N_6841);
nor U8476 (N_8476,N_6325,N_6239);
and U8477 (N_8477,N_6501,N_7409);
nand U8478 (N_8478,N_7789,N_7404);
nand U8479 (N_8479,N_6888,N_6200);
nor U8480 (N_8480,N_7917,N_7334);
and U8481 (N_8481,N_7826,N_7031);
nand U8482 (N_8482,N_6470,N_7685);
xor U8483 (N_8483,N_6087,N_6722);
and U8484 (N_8484,N_7136,N_7121);
nand U8485 (N_8485,N_7704,N_6176);
nor U8486 (N_8486,N_6451,N_6730);
nand U8487 (N_8487,N_6137,N_7211);
nor U8488 (N_8488,N_6673,N_6297);
xor U8489 (N_8489,N_6469,N_6241);
or U8490 (N_8490,N_7732,N_7632);
xnor U8491 (N_8491,N_7899,N_6550);
and U8492 (N_8492,N_7366,N_7970);
and U8493 (N_8493,N_6578,N_6616);
nor U8494 (N_8494,N_6020,N_7011);
and U8495 (N_8495,N_6208,N_7850);
xnor U8496 (N_8496,N_6035,N_7384);
nor U8497 (N_8497,N_6396,N_7221);
xnor U8498 (N_8498,N_6703,N_6788);
and U8499 (N_8499,N_7546,N_6749);
nand U8500 (N_8500,N_7500,N_7039);
nor U8501 (N_8501,N_7431,N_7320);
xnor U8502 (N_8502,N_6237,N_6427);
nor U8503 (N_8503,N_7774,N_7312);
nand U8504 (N_8504,N_6983,N_7365);
nand U8505 (N_8505,N_6797,N_7226);
and U8506 (N_8506,N_7928,N_6199);
nor U8507 (N_8507,N_7085,N_6077);
or U8508 (N_8508,N_7247,N_7583);
or U8509 (N_8509,N_7571,N_6221);
and U8510 (N_8510,N_7491,N_6986);
nand U8511 (N_8511,N_6904,N_7781);
or U8512 (N_8512,N_7793,N_7315);
or U8513 (N_8513,N_7038,N_6744);
nand U8514 (N_8514,N_6472,N_6516);
nand U8515 (N_8515,N_6940,N_7274);
nand U8516 (N_8516,N_6450,N_7881);
or U8517 (N_8517,N_6401,N_6264);
nor U8518 (N_8518,N_6367,N_7192);
nor U8519 (N_8519,N_7768,N_6356);
and U8520 (N_8520,N_7273,N_7559);
and U8521 (N_8521,N_6464,N_6671);
and U8522 (N_8522,N_7645,N_7661);
nor U8523 (N_8523,N_7216,N_6933);
nand U8524 (N_8524,N_7859,N_7240);
and U8525 (N_8525,N_7517,N_6826);
nand U8526 (N_8526,N_7622,N_7452);
or U8527 (N_8527,N_6837,N_6227);
nand U8528 (N_8528,N_6820,N_7357);
nor U8529 (N_8529,N_7818,N_7296);
nor U8530 (N_8530,N_6736,N_6885);
xor U8531 (N_8531,N_7458,N_6946);
nand U8532 (N_8532,N_6623,N_7947);
or U8533 (N_8533,N_7470,N_7794);
or U8534 (N_8534,N_7502,N_6711);
nor U8535 (N_8535,N_7468,N_7248);
xor U8536 (N_8536,N_6941,N_7892);
nand U8537 (N_8537,N_6103,N_7960);
xor U8538 (N_8538,N_6897,N_6526);
or U8539 (N_8539,N_6303,N_6184);
or U8540 (N_8540,N_7968,N_6223);
xor U8541 (N_8541,N_7236,N_7751);
or U8542 (N_8542,N_6443,N_6418);
or U8543 (N_8543,N_7317,N_6291);
nor U8544 (N_8544,N_7020,N_7808);
nor U8545 (N_8545,N_6397,N_6566);
or U8546 (N_8546,N_7207,N_6865);
and U8547 (N_8547,N_6128,N_6921);
xnor U8548 (N_8548,N_7267,N_7887);
nor U8549 (N_8549,N_7741,N_6600);
xnor U8550 (N_8550,N_6907,N_6658);
nand U8551 (N_8551,N_6615,N_6594);
nand U8552 (N_8552,N_6014,N_7271);
and U8553 (N_8553,N_7640,N_6776);
xor U8554 (N_8554,N_6560,N_7417);
xnor U8555 (N_8555,N_6424,N_7969);
nand U8556 (N_8556,N_6403,N_6833);
and U8557 (N_8557,N_6773,N_7838);
or U8558 (N_8558,N_6048,N_6226);
xnor U8559 (N_8559,N_6800,N_7542);
xor U8560 (N_8560,N_7130,N_7067);
and U8561 (N_8561,N_7339,N_7111);
and U8562 (N_8562,N_6923,N_7744);
nand U8563 (N_8563,N_6205,N_6992);
or U8564 (N_8564,N_7637,N_6545);
nor U8565 (N_8565,N_6363,N_7900);
xor U8566 (N_8566,N_7842,N_7675);
and U8567 (N_8567,N_7040,N_7612);
xnor U8568 (N_8568,N_6089,N_7326);
or U8569 (N_8569,N_7323,N_7134);
or U8570 (N_8570,N_7802,N_7805);
nor U8571 (N_8571,N_6936,N_7912);
nand U8572 (N_8572,N_6265,N_7269);
xor U8573 (N_8573,N_6883,N_7308);
and U8574 (N_8574,N_7100,N_6055);
and U8575 (N_8575,N_6824,N_6995);
or U8576 (N_8576,N_7414,N_6521);
xor U8577 (N_8577,N_7266,N_7219);
and U8578 (N_8578,N_7536,N_7513);
nor U8579 (N_8579,N_7760,N_7138);
and U8580 (N_8580,N_6160,N_6382);
xnor U8581 (N_8581,N_6934,N_6335);
nand U8582 (N_8582,N_6537,N_7976);
and U8583 (N_8583,N_6281,N_7625);
and U8584 (N_8584,N_6315,N_7740);
and U8585 (N_8585,N_7653,N_7883);
or U8586 (N_8586,N_6620,N_6271);
nand U8587 (N_8587,N_7688,N_7918);
and U8588 (N_8588,N_6529,N_6354);
nor U8589 (N_8589,N_6859,N_7535);
xor U8590 (N_8590,N_7074,N_7287);
nand U8591 (N_8591,N_7201,N_6222);
nand U8592 (N_8592,N_7407,N_7966);
nor U8593 (N_8593,N_6349,N_6794);
xor U8594 (N_8594,N_6575,N_6954);
and U8595 (N_8595,N_7281,N_6016);
nor U8596 (N_8596,N_7107,N_7799);
xnor U8597 (N_8597,N_6649,N_7213);
nor U8598 (N_8598,N_7949,N_7441);
xnor U8599 (N_8599,N_7771,N_7840);
and U8600 (N_8600,N_6285,N_6258);
nand U8601 (N_8601,N_7907,N_7057);
xor U8602 (N_8602,N_7572,N_7005);
xor U8603 (N_8603,N_7832,N_7127);
nor U8604 (N_8604,N_6970,N_6540);
xor U8605 (N_8605,N_6253,N_6500);
nor U8606 (N_8606,N_7757,N_6288);
xor U8607 (N_8607,N_6984,N_7050);
xor U8608 (N_8608,N_6095,N_7816);
xor U8609 (N_8609,N_7069,N_7931);
or U8610 (N_8610,N_7181,N_6278);
or U8611 (N_8611,N_6927,N_6082);
and U8612 (N_8612,N_7991,N_7055);
or U8613 (N_8613,N_6964,N_6544);
or U8614 (N_8614,N_7242,N_7884);
nor U8615 (N_8615,N_7716,N_6196);
or U8616 (N_8616,N_7146,N_6072);
nor U8617 (N_8617,N_7048,N_7410);
and U8618 (N_8618,N_6232,N_7402);
nand U8619 (N_8619,N_7600,N_6279);
xor U8620 (N_8620,N_7002,N_7829);
or U8621 (N_8621,N_6613,N_6978);
xor U8622 (N_8622,N_6430,N_6129);
nand U8623 (N_8623,N_6124,N_7745);
nor U8624 (N_8624,N_6815,N_7486);
and U8625 (N_8625,N_7325,N_7667);
or U8626 (N_8626,N_7283,N_7062);
or U8627 (N_8627,N_6003,N_6796);
nand U8628 (N_8628,N_6867,N_7228);
xor U8629 (N_8629,N_6597,N_6168);
or U8630 (N_8630,N_7642,N_6918);
and U8631 (N_8631,N_6593,N_6044);
nand U8632 (N_8632,N_6100,N_7220);
nand U8633 (N_8633,N_6434,N_6761);
and U8634 (N_8634,N_6908,N_6352);
nor U8635 (N_8635,N_6650,N_7897);
nand U8636 (N_8636,N_6710,N_6444);
nor U8637 (N_8637,N_6892,N_6034);
nor U8638 (N_8638,N_7770,N_7204);
nand U8639 (N_8639,N_6974,N_7173);
xnor U8640 (N_8640,N_6844,N_7350);
and U8641 (N_8641,N_6365,N_7830);
xor U8642 (N_8642,N_6449,N_7290);
or U8643 (N_8643,N_7036,N_6280);
nand U8644 (N_8644,N_7362,N_7024);
nor U8645 (N_8645,N_6701,N_7145);
xor U8646 (N_8646,N_7141,N_7443);
nand U8647 (N_8647,N_7046,N_6831);
nor U8648 (N_8648,N_7545,N_7700);
and U8649 (N_8649,N_6691,N_7429);
nor U8650 (N_8650,N_7893,N_7177);
nand U8651 (N_8651,N_6767,N_7434);
and U8652 (N_8652,N_6667,N_6519);
and U8653 (N_8653,N_6186,N_7582);
nor U8654 (N_8654,N_6882,N_6155);
and U8655 (N_8655,N_6345,N_7725);
or U8656 (N_8656,N_6769,N_7104);
xor U8657 (N_8657,N_7185,N_6311);
and U8658 (N_8658,N_7785,N_7649);
nand U8659 (N_8659,N_6971,N_6276);
and U8660 (N_8660,N_7910,N_6039);
or U8661 (N_8661,N_6926,N_7844);
xor U8662 (N_8662,N_7217,N_7282);
nor U8663 (N_8663,N_7421,N_7007);
xnor U8664 (N_8664,N_7558,N_7520);
nand U8665 (N_8665,N_7715,N_7763);
nand U8666 (N_8666,N_6568,N_7176);
nor U8667 (N_8667,N_6052,N_6299);
and U8668 (N_8668,N_6251,N_7512);
xnor U8669 (N_8669,N_7353,N_7656);
nand U8670 (N_8670,N_6661,N_7595);
nor U8671 (N_8671,N_7208,N_6182);
xor U8672 (N_8672,N_6552,N_7644);
nand U8673 (N_8673,N_6699,N_6318);
xor U8674 (N_8674,N_7380,N_6307);
xor U8675 (N_8675,N_7690,N_6247);
nand U8676 (N_8676,N_7510,N_6005);
nand U8677 (N_8677,N_7060,N_6132);
and U8678 (N_8678,N_7408,N_6792);
or U8679 (N_8679,N_6069,N_6491);
nand U8680 (N_8680,N_6963,N_7666);
and U8681 (N_8681,N_7022,N_6979);
or U8682 (N_8682,N_6531,N_6949);
xor U8683 (N_8683,N_6572,N_7596);
and U8684 (N_8684,N_6561,N_7255);
nor U8685 (N_8685,N_7279,N_7660);
nand U8686 (N_8686,N_6924,N_6454);
or U8687 (N_8687,N_7180,N_6731);
nand U8688 (N_8688,N_7695,N_7599);
nor U8689 (N_8689,N_6990,N_6762);
nor U8690 (N_8690,N_7848,N_6375);
and U8691 (N_8691,N_6000,N_7919);
or U8692 (N_8692,N_6828,N_7238);
xnor U8693 (N_8693,N_7335,N_6720);
nor U8694 (N_8694,N_7726,N_7378);
nor U8695 (N_8695,N_6115,N_7995);
or U8696 (N_8696,N_6685,N_7762);
or U8697 (N_8697,N_7088,N_6887);
or U8698 (N_8698,N_7717,N_7791);
or U8699 (N_8699,N_7586,N_7719);
and U8700 (N_8700,N_6580,N_7532);
nor U8701 (N_8701,N_7696,N_7116);
xnor U8702 (N_8702,N_6085,N_7909);
xnor U8703 (N_8703,N_6138,N_6607);
nor U8704 (N_8704,N_7309,N_6805);
xor U8705 (N_8705,N_6868,N_6341);
nand U8706 (N_8706,N_6306,N_6876);
xnor U8707 (N_8707,N_6719,N_7054);
and U8708 (N_8708,N_6832,N_6680);
and U8709 (N_8709,N_6342,N_7338);
or U8710 (N_8710,N_7097,N_7193);
xnor U8711 (N_8711,N_6273,N_6611);
xor U8712 (N_8712,N_7944,N_7152);
and U8713 (N_8713,N_7330,N_7422);
nor U8714 (N_8714,N_6579,N_6012);
or U8715 (N_8715,N_7709,N_6046);
or U8716 (N_8716,N_6314,N_6582);
xnor U8717 (N_8717,N_6606,N_6873);
and U8718 (N_8718,N_6482,N_7738);
and U8719 (N_8719,N_7065,N_7866);
nand U8720 (N_8720,N_7555,N_6627);
nand U8721 (N_8721,N_6848,N_7523);
and U8722 (N_8722,N_6287,N_6193);
nand U8723 (N_8723,N_7190,N_6488);
nor U8724 (N_8724,N_6952,N_7560);
xnor U8725 (N_8725,N_7888,N_6113);
and U8726 (N_8726,N_6602,N_6204);
nor U8727 (N_8727,N_6432,N_7272);
nand U8728 (N_8728,N_6770,N_6084);
xnor U8729 (N_8729,N_6006,N_7117);
nor U8730 (N_8730,N_6209,N_6741);
or U8731 (N_8731,N_7030,N_7986);
xnor U8732 (N_8732,N_6038,N_6161);
xnor U8733 (N_8733,N_6838,N_7906);
and U8734 (N_8734,N_7425,N_6502);
nor U8735 (N_8735,N_7254,N_7128);
nor U8736 (N_8736,N_7389,N_6484);
xor U8737 (N_8737,N_6628,N_7813);
and U8738 (N_8738,N_6233,N_6114);
nand U8739 (N_8739,N_7268,N_6130);
nand U8740 (N_8740,N_6621,N_7698);
xor U8741 (N_8741,N_6059,N_7184);
or U8742 (N_8742,N_6622,N_6745);
nor U8743 (N_8743,N_6202,N_7482);
nor U8744 (N_8744,N_7655,N_6512);
and U8745 (N_8745,N_6562,N_7115);
nor U8746 (N_8746,N_7952,N_6823);
nor U8747 (N_8747,N_7071,N_6421);
nand U8748 (N_8748,N_6558,N_7123);
and U8749 (N_8749,N_6042,N_6293);
and U8750 (N_8750,N_7322,N_6525);
or U8751 (N_8751,N_6181,N_7554);
and U8752 (N_8752,N_7387,N_6167);
nor U8753 (N_8753,N_6492,N_7857);
nor U8754 (N_8754,N_7563,N_6758);
nand U8755 (N_8755,N_6023,N_7618);
and U8756 (N_8756,N_6588,N_7878);
and U8757 (N_8757,N_7911,N_7223);
nor U8758 (N_8758,N_6249,N_7033);
and U8759 (N_8759,N_6217,N_6605);
nand U8760 (N_8760,N_6210,N_7165);
and U8761 (N_8761,N_6697,N_7314);
and U8762 (N_8762,N_7609,N_7096);
or U8763 (N_8763,N_7169,N_6415);
or U8764 (N_8764,N_6879,N_6663);
nor U8765 (N_8765,N_7748,N_7156);
nand U8766 (N_8766,N_7080,N_7626);
and U8767 (N_8767,N_6662,N_7131);
or U8768 (N_8768,N_7469,N_6144);
and U8769 (N_8769,N_7978,N_7591);
and U8770 (N_8770,N_6969,N_7465);
xor U8771 (N_8771,N_6958,N_6814);
xnor U8772 (N_8772,N_7996,N_7120);
and U8773 (N_8773,N_7235,N_7646);
and U8774 (N_8774,N_6146,N_6142);
and U8775 (N_8775,N_6513,N_7651);
and U8776 (N_8776,N_6639,N_6147);
nor U8777 (N_8777,N_6968,N_6485);
xnor U8778 (N_8778,N_7544,N_7705);
nor U8779 (N_8779,N_7654,N_6357);
or U8780 (N_8780,N_6099,N_7292);
and U8781 (N_8781,N_6018,N_7360);
nand U8782 (N_8782,N_6543,N_6081);
and U8783 (N_8783,N_7497,N_7206);
xnor U8784 (N_8784,N_6584,N_6655);
nor U8785 (N_8785,N_7041,N_7006);
and U8786 (N_8786,N_7574,N_6712);
and U8787 (N_8787,N_6806,N_6764);
xnor U8788 (N_8788,N_6440,N_6533);
or U8789 (N_8789,N_6368,N_6457);
xnor U8790 (N_8790,N_7670,N_6198);
nand U8791 (N_8791,N_6292,N_6353);
nand U8792 (N_8792,N_6257,N_6238);
nor U8793 (N_8793,N_6461,N_6937);
nor U8794 (N_8794,N_7961,N_7742);
and U8795 (N_8795,N_7590,N_7879);
nand U8796 (N_8796,N_6676,N_7474);
and U8797 (N_8797,N_6304,N_7321);
xnor U8798 (N_8798,N_7643,N_6829);
nand U8799 (N_8799,N_7501,N_6724);
and U8800 (N_8800,N_6185,N_6592);
nand U8801 (N_8801,N_6133,N_7418);
nand U8802 (N_8802,N_6101,N_6877);
and U8803 (N_8803,N_7370,N_6067);
nor U8804 (N_8804,N_6324,N_7303);
xor U8805 (N_8805,N_6573,N_6387);
or U8806 (N_8806,N_7930,N_7233);
nor U8807 (N_8807,N_6596,N_7025);
and U8808 (N_8808,N_6523,N_6489);
and U8809 (N_8809,N_6960,N_6385);
xnor U8810 (N_8810,N_7275,N_6539);
and U8811 (N_8811,N_7737,N_6148);
nand U8812 (N_8812,N_7743,N_6096);
nand U8813 (N_8813,N_7849,N_7853);
or U8814 (N_8814,N_7766,N_6948);
or U8815 (N_8815,N_7393,N_6779);
nor U8816 (N_8816,N_6021,N_7457);
xor U8817 (N_8817,N_6517,N_7875);
or U8818 (N_8818,N_6916,N_6910);
or U8819 (N_8819,N_7245,N_6700);
and U8820 (N_8820,N_7081,N_6604);
xor U8821 (N_8821,N_7531,N_6846);
xor U8822 (N_8822,N_7118,N_7773);
or U8823 (N_8823,N_6871,N_7822);
nand U8824 (N_8824,N_7620,N_6030);
or U8825 (N_8825,N_7831,N_7354);
xor U8826 (N_8826,N_7658,N_6635);
and U8827 (N_8827,N_6395,N_6466);
nand U8828 (N_8828,N_7593,N_7280);
and U8829 (N_8829,N_6010,N_6183);
or U8830 (N_8830,N_7398,N_7261);
nand U8831 (N_8831,N_7566,N_7689);
xnor U8832 (N_8832,N_6422,N_7298);
or U8833 (N_8833,N_7481,N_7197);
and U8834 (N_8834,N_7110,N_6121);
or U8835 (N_8835,N_6835,N_7965);
nand U8836 (N_8836,N_6073,N_7396);
and U8837 (N_8837,N_7051,N_6689);
and U8838 (N_8838,N_6328,N_7898);
xor U8839 (N_8839,N_7607,N_6370);
or U8840 (N_8840,N_6881,N_6688);
and U8841 (N_8841,N_7938,N_6391);
and U8842 (N_8842,N_7151,N_7872);
nand U8843 (N_8843,N_7150,N_6624);
nand U8844 (N_8844,N_7904,N_7729);
xnor U8845 (N_8845,N_6959,N_7199);
and U8846 (N_8846,N_7538,N_6097);
nand U8847 (N_8847,N_6791,N_6931);
xor U8848 (N_8848,N_7073,N_6108);
nor U8849 (N_8849,N_7581,N_6456);
nand U8850 (N_8850,N_7613,N_7297);
nand U8851 (N_8851,N_7058,N_7557);
xnor U8852 (N_8852,N_6956,N_7795);
xor U8853 (N_8853,N_6197,N_7037);
xor U8854 (N_8854,N_6922,N_6399);
nor U8855 (N_8855,N_7908,N_7371);
nand U8856 (N_8856,N_6347,N_6765);
nand U8857 (N_8857,N_6707,N_7712);
nand U8858 (N_8858,N_7750,N_7954);
and U8859 (N_8859,N_7450,N_7284);
nand U8860 (N_8860,N_7941,N_7975);
and U8861 (N_8861,N_6270,N_7610);
and U8862 (N_8862,N_7948,N_6094);
xnor U8863 (N_8863,N_6216,N_7569);
nor U8864 (N_8864,N_6041,N_6713);
nor U8865 (N_8865,N_7797,N_7549);
and U8866 (N_8866,N_7093,N_6763);
nor U8867 (N_8867,N_7876,N_7973);
nor U8868 (N_8868,N_7980,N_6660);
or U8869 (N_8869,N_6739,N_7122);
nor U8870 (N_8870,N_7343,N_6412);
nor U8871 (N_8871,N_6803,N_6333);
xnor U8872 (N_8872,N_7013,N_7423);
and U8873 (N_8873,N_6337,N_7761);
and U8874 (N_8874,N_7570,N_6756);
nand U8875 (N_8875,N_6640,N_7485);
nand U8876 (N_8876,N_7126,N_6423);
or U8877 (N_8877,N_7349,N_7652);
nor U8878 (N_8878,N_6060,N_6049);
xnor U8879 (N_8879,N_7397,N_6007);
or U8880 (N_8880,N_7383,N_6854);
and U8881 (N_8881,N_7017,N_7166);
xor U8882 (N_8882,N_6801,N_7187);
xnor U8883 (N_8883,N_7311,N_7332);
or U8884 (N_8884,N_6809,N_6017);
or U8885 (N_8885,N_6317,N_7237);
nor U8886 (N_8886,N_6679,N_6054);
and U8887 (N_8887,N_7945,N_6507);
xnor U8888 (N_8888,N_7243,N_6474);
nor U8889 (N_8889,N_6783,N_6930);
nor U8890 (N_8890,N_7678,N_6752);
nand U8891 (N_8891,N_7573,N_6678);
nand U8892 (N_8892,N_7747,N_7045);
or U8893 (N_8893,N_7427,N_6047);
nand U8894 (N_8894,N_7937,N_6812);
nand U8895 (N_8895,N_7929,N_6126);
and U8896 (N_8896,N_6705,N_7277);
xor U8897 (N_8897,N_7999,N_6947);
or U8898 (N_8898,N_6481,N_6997);
xor U8899 (N_8899,N_6417,N_6388);
xor U8900 (N_8900,N_7270,N_7189);
xor U8901 (N_8901,N_6760,N_6980);
nand U8902 (N_8902,N_7008,N_6618);
xor U8903 (N_8903,N_7727,N_6643);
or U8904 (N_8904,N_7603,N_6869);
and U8905 (N_8905,N_7379,N_7819);
nand U8906 (N_8906,N_6170,N_7550);
and U8907 (N_8907,N_7499,N_7346);
and U8908 (N_8908,N_6813,N_6938);
nand U8909 (N_8909,N_7101,N_6252);
xor U8910 (N_8910,N_6381,N_6585);
nor U8911 (N_8911,N_7858,N_6884);
nor U8912 (N_8912,N_6850,N_7089);
xor U8913 (N_8913,N_6836,N_6091);
xnor U8914 (N_8914,N_6398,N_7484);
xnor U8915 (N_8915,N_7933,N_7301);
xnor U8916 (N_8916,N_7854,N_7530);
xnor U8917 (N_8917,N_7617,N_7401);
or U8918 (N_8918,N_7289,N_6453);
nand U8919 (N_8919,N_7846,N_6619);
or U8920 (N_8920,N_6371,N_6494);
and U8921 (N_8921,N_6753,N_7498);
or U8922 (N_8922,N_7459,N_7841);
nand U8923 (N_8923,N_7043,N_6083);
nor U8924 (N_8924,N_7800,N_6953);
nand U8925 (N_8925,N_7302,N_7157);
and U8926 (N_8926,N_7299,N_7372);
and U8927 (N_8927,N_7493,N_6906);
xnor U8928 (N_8928,N_6106,N_6925);
and U8929 (N_8929,N_6569,N_6022);
nand U8930 (N_8930,N_6905,N_7915);
nor U8931 (N_8931,N_6998,N_7395);
xnor U8932 (N_8932,N_7998,N_7955);
nor U8933 (N_8933,N_7812,N_6187);
nor U8934 (N_8934,N_6880,N_7672);
nand U8935 (N_8935,N_7776,N_6858);
or U8936 (N_8936,N_7003,N_6364);
xnor U8937 (N_8937,N_6577,N_7886);
nor U8938 (N_8938,N_6071,N_7001);
xor U8939 (N_8939,N_6150,N_7344);
nand U8940 (N_8940,N_6442,N_6476);
and U8941 (N_8941,N_6506,N_7605);
nor U8942 (N_8942,N_7019,N_6694);
nor U8943 (N_8943,N_7369,N_6157);
and U8944 (N_8944,N_6477,N_7178);
and U8945 (N_8945,N_7105,N_7865);
xor U8946 (N_8946,N_7047,N_7420);
nor U8947 (N_8947,N_7476,N_6681);
nand U8948 (N_8948,N_6518,N_6250);
nand U8949 (N_8949,N_6224,N_6514);
and U8950 (N_8950,N_6674,N_6290);
xor U8951 (N_8951,N_6630,N_6634);
nand U8952 (N_8952,N_6331,N_6498);
and U8953 (N_8953,N_6644,N_6286);
xnor U8954 (N_8954,N_7511,N_6230);
and U8955 (N_8955,N_7598,N_6438);
or U8956 (N_8956,N_7456,N_6857);
and U8957 (N_8957,N_7153,N_7432);
xor U8958 (N_8958,N_7835,N_6123);
or U8959 (N_8959,N_7964,N_6350);
and U8960 (N_8960,N_7504,N_7077);
nand U8961 (N_8961,N_6782,N_6781);
and U8962 (N_8962,N_7529,N_6164);
xnor U8963 (N_8963,N_7979,N_7244);
and U8964 (N_8964,N_6070,N_6900);
and U8965 (N_8965,N_7606,N_7026);
and U8966 (N_8966,N_6441,N_6355);
xor U8967 (N_8967,N_7756,N_6778);
or U8968 (N_8968,N_6977,N_6191);
or U8969 (N_8969,N_6319,N_6212);
or U8970 (N_8970,N_6246,N_6244);
nand U8971 (N_8971,N_6913,N_7755);
and U8972 (N_8972,N_7896,N_7522);
or U8973 (N_8973,N_6312,N_7078);
nand U8974 (N_8974,N_7000,N_6875);
xnor U8975 (N_8975,N_6768,N_6105);
nor U8976 (N_8976,N_7433,N_7318);
nand U8977 (N_8977,N_7638,N_7753);
nor U8978 (N_8978,N_7874,N_7412);
and U8979 (N_8979,N_6207,N_6855);
nor U8980 (N_8980,N_6379,N_7552);
and U8981 (N_8981,N_6799,N_7694);
and U8982 (N_8982,N_7992,N_7451);
nor U8983 (N_8983,N_7659,N_6171);
xnor U8984 (N_8984,N_6151,N_6439);
nor U8985 (N_8985,N_6463,N_7521);
nor U8986 (N_8986,N_7480,N_7792);
and U8987 (N_8987,N_6483,N_7095);
and U8988 (N_8988,N_7824,N_6493);
or U8989 (N_8989,N_7633,N_6024);
and U8990 (N_8990,N_7775,N_7461);
or U8991 (N_8991,N_7258,N_7553);
or U8992 (N_8992,N_6896,N_7508);
or U8993 (N_8993,N_7648,N_6571);
xor U8994 (N_8994,N_6013,N_7814);
and U8995 (N_8995,N_7340,N_6383);
xor U8996 (N_8996,N_6878,N_7519);
or U8997 (N_8997,N_7359,N_7588);
nand U8998 (N_8998,N_7920,N_6025);
nand U8999 (N_8999,N_7537,N_7072);
or U9000 (N_9000,N_7698,N_6903);
nor U9001 (N_9001,N_6295,N_7559);
and U9002 (N_9002,N_6649,N_6944);
and U9003 (N_9003,N_7958,N_6694);
and U9004 (N_9004,N_6472,N_7376);
or U9005 (N_9005,N_7818,N_6226);
xor U9006 (N_9006,N_6055,N_7688);
or U9007 (N_9007,N_6265,N_6441);
nor U9008 (N_9008,N_7269,N_6517);
nor U9009 (N_9009,N_7474,N_7662);
nor U9010 (N_9010,N_6205,N_7771);
nor U9011 (N_9011,N_6487,N_6877);
or U9012 (N_9012,N_7530,N_7694);
nor U9013 (N_9013,N_7134,N_7754);
nand U9014 (N_9014,N_7407,N_6160);
nor U9015 (N_9015,N_7185,N_6013);
or U9016 (N_9016,N_6240,N_6841);
and U9017 (N_9017,N_6360,N_7889);
or U9018 (N_9018,N_7305,N_6927);
nand U9019 (N_9019,N_7597,N_6617);
nand U9020 (N_9020,N_7469,N_7950);
and U9021 (N_9021,N_7040,N_6526);
and U9022 (N_9022,N_7999,N_7536);
nor U9023 (N_9023,N_7816,N_7377);
or U9024 (N_9024,N_7230,N_7653);
nand U9025 (N_9025,N_6789,N_7741);
nor U9026 (N_9026,N_7596,N_6475);
xnor U9027 (N_9027,N_6438,N_7914);
xor U9028 (N_9028,N_7287,N_6923);
xor U9029 (N_9029,N_6578,N_6045);
and U9030 (N_9030,N_7826,N_7898);
xnor U9031 (N_9031,N_7179,N_6342);
and U9032 (N_9032,N_7361,N_7109);
nor U9033 (N_9033,N_7918,N_7950);
or U9034 (N_9034,N_6121,N_7488);
nand U9035 (N_9035,N_7668,N_7670);
nand U9036 (N_9036,N_7897,N_6134);
and U9037 (N_9037,N_6180,N_7960);
and U9038 (N_9038,N_6730,N_7500);
nor U9039 (N_9039,N_7767,N_6013);
nor U9040 (N_9040,N_7113,N_7142);
nor U9041 (N_9041,N_6139,N_6267);
and U9042 (N_9042,N_6389,N_6887);
xnor U9043 (N_9043,N_6654,N_7291);
xor U9044 (N_9044,N_7194,N_7684);
nor U9045 (N_9045,N_7341,N_7958);
nor U9046 (N_9046,N_6985,N_6821);
and U9047 (N_9047,N_7792,N_7392);
nand U9048 (N_9048,N_6848,N_6862);
xor U9049 (N_9049,N_7049,N_7125);
or U9050 (N_9050,N_6177,N_7008);
xnor U9051 (N_9051,N_6105,N_6321);
and U9052 (N_9052,N_7331,N_7663);
and U9053 (N_9053,N_7328,N_6911);
nor U9054 (N_9054,N_6822,N_6041);
nand U9055 (N_9055,N_6817,N_6607);
xnor U9056 (N_9056,N_7469,N_7711);
or U9057 (N_9057,N_6132,N_6362);
nand U9058 (N_9058,N_6598,N_7123);
xor U9059 (N_9059,N_6641,N_6903);
nor U9060 (N_9060,N_7527,N_7293);
and U9061 (N_9061,N_6009,N_7861);
or U9062 (N_9062,N_6627,N_6882);
and U9063 (N_9063,N_7624,N_7131);
or U9064 (N_9064,N_6380,N_6974);
nor U9065 (N_9065,N_7234,N_6626);
xor U9066 (N_9066,N_7107,N_6126);
and U9067 (N_9067,N_7709,N_6569);
and U9068 (N_9068,N_6436,N_6834);
or U9069 (N_9069,N_7600,N_7892);
nor U9070 (N_9070,N_6010,N_7515);
nor U9071 (N_9071,N_7176,N_6331);
and U9072 (N_9072,N_7387,N_6644);
nor U9073 (N_9073,N_6645,N_6783);
nand U9074 (N_9074,N_7127,N_6204);
or U9075 (N_9075,N_6601,N_7263);
nor U9076 (N_9076,N_7968,N_7198);
and U9077 (N_9077,N_7908,N_6869);
nand U9078 (N_9078,N_6426,N_7565);
and U9079 (N_9079,N_6001,N_6417);
nor U9080 (N_9080,N_6313,N_7386);
and U9081 (N_9081,N_7094,N_7151);
xor U9082 (N_9082,N_6189,N_6697);
xnor U9083 (N_9083,N_7384,N_6351);
nand U9084 (N_9084,N_6173,N_6977);
xor U9085 (N_9085,N_7835,N_7204);
and U9086 (N_9086,N_6204,N_6808);
xnor U9087 (N_9087,N_6940,N_6859);
xnor U9088 (N_9088,N_6002,N_7584);
nand U9089 (N_9089,N_7685,N_7204);
nand U9090 (N_9090,N_7519,N_6078);
nor U9091 (N_9091,N_7088,N_6960);
nand U9092 (N_9092,N_6377,N_6744);
or U9093 (N_9093,N_6562,N_6925);
or U9094 (N_9094,N_7274,N_7949);
and U9095 (N_9095,N_7710,N_6559);
and U9096 (N_9096,N_7924,N_7603);
nand U9097 (N_9097,N_7581,N_7963);
xnor U9098 (N_9098,N_6226,N_6246);
nand U9099 (N_9099,N_6804,N_6356);
nor U9100 (N_9100,N_7972,N_7475);
and U9101 (N_9101,N_6047,N_6057);
nor U9102 (N_9102,N_6709,N_6276);
nand U9103 (N_9103,N_6565,N_7618);
nor U9104 (N_9104,N_6982,N_6408);
or U9105 (N_9105,N_6125,N_7713);
or U9106 (N_9106,N_7297,N_7350);
xnor U9107 (N_9107,N_6973,N_6148);
xnor U9108 (N_9108,N_7622,N_6995);
xnor U9109 (N_9109,N_7641,N_6466);
or U9110 (N_9110,N_6078,N_7310);
nand U9111 (N_9111,N_6803,N_6787);
nand U9112 (N_9112,N_7144,N_6752);
nand U9113 (N_9113,N_6465,N_7203);
and U9114 (N_9114,N_7492,N_6913);
and U9115 (N_9115,N_6794,N_7916);
or U9116 (N_9116,N_6778,N_6487);
nand U9117 (N_9117,N_7973,N_7315);
or U9118 (N_9118,N_6316,N_6615);
xnor U9119 (N_9119,N_6211,N_6598);
and U9120 (N_9120,N_6017,N_7847);
nor U9121 (N_9121,N_6376,N_6562);
nand U9122 (N_9122,N_7213,N_6560);
or U9123 (N_9123,N_6233,N_7765);
xor U9124 (N_9124,N_6571,N_6078);
nor U9125 (N_9125,N_6334,N_6591);
and U9126 (N_9126,N_7346,N_6679);
or U9127 (N_9127,N_6373,N_7298);
nor U9128 (N_9128,N_7119,N_6914);
xor U9129 (N_9129,N_7433,N_7417);
and U9130 (N_9130,N_7361,N_6457);
nand U9131 (N_9131,N_6619,N_7742);
nor U9132 (N_9132,N_6408,N_7070);
xnor U9133 (N_9133,N_6358,N_7568);
nor U9134 (N_9134,N_7490,N_6947);
and U9135 (N_9135,N_7712,N_7964);
nor U9136 (N_9136,N_6047,N_6186);
nor U9137 (N_9137,N_6601,N_6874);
nor U9138 (N_9138,N_7641,N_6508);
or U9139 (N_9139,N_6781,N_6762);
xor U9140 (N_9140,N_6078,N_6413);
xnor U9141 (N_9141,N_7913,N_6339);
xnor U9142 (N_9142,N_7333,N_7206);
and U9143 (N_9143,N_7009,N_6758);
nor U9144 (N_9144,N_7764,N_6103);
nand U9145 (N_9145,N_7988,N_6624);
or U9146 (N_9146,N_6827,N_6968);
xor U9147 (N_9147,N_7294,N_6571);
nor U9148 (N_9148,N_6936,N_7497);
xnor U9149 (N_9149,N_7548,N_7208);
nor U9150 (N_9150,N_6096,N_7474);
nand U9151 (N_9151,N_6273,N_6980);
xor U9152 (N_9152,N_6785,N_7905);
nor U9153 (N_9153,N_6184,N_6137);
xor U9154 (N_9154,N_7631,N_7079);
and U9155 (N_9155,N_7354,N_6735);
nand U9156 (N_9156,N_6446,N_6469);
nor U9157 (N_9157,N_6895,N_7456);
nand U9158 (N_9158,N_6030,N_7867);
and U9159 (N_9159,N_6849,N_6300);
nand U9160 (N_9160,N_7197,N_6781);
and U9161 (N_9161,N_7920,N_7603);
or U9162 (N_9162,N_6275,N_7973);
xnor U9163 (N_9163,N_7451,N_7733);
and U9164 (N_9164,N_6672,N_6684);
and U9165 (N_9165,N_6162,N_7188);
and U9166 (N_9166,N_6220,N_6021);
or U9167 (N_9167,N_6282,N_6371);
nand U9168 (N_9168,N_6253,N_7003);
or U9169 (N_9169,N_6656,N_7527);
and U9170 (N_9170,N_7538,N_7872);
nand U9171 (N_9171,N_6042,N_6768);
or U9172 (N_9172,N_6089,N_6234);
and U9173 (N_9173,N_7474,N_6688);
nand U9174 (N_9174,N_6605,N_6523);
nand U9175 (N_9175,N_7162,N_7656);
xor U9176 (N_9176,N_6082,N_7496);
or U9177 (N_9177,N_6427,N_7767);
nor U9178 (N_9178,N_6252,N_7363);
and U9179 (N_9179,N_6420,N_6148);
nor U9180 (N_9180,N_6301,N_7927);
nor U9181 (N_9181,N_7110,N_7282);
nand U9182 (N_9182,N_6736,N_7523);
nand U9183 (N_9183,N_7652,N_6440);
xnor U9184 (N_9184,N_6609,N_7273);
xor U9185 (N_9185,N_7718,N_6677);
nand U9186 (N_9186,N_7789,N_6910);
and U9187 (N_9187,N_6139,N_7527);
xnor U9188 (N_9188,N_6254,N_7528);
nor U9189 (N_9189,N_7838,N_7535);
nand U9190 (N_9190,N_7506,N_6367);
xor U9191 (N_9191,N_7809,N_7241);
xnor U9192 (N_9192,N_7113,N_7713);
nand U9193 (N_9193,N_7501,N_6574);
xor U9194 (N_9194,N_6513,N_7201);
or U9195 (N_9195,N_7538,N_6373);
or U9196 (N_9196,N_7076,N_7759);
and U9197 (N_9197,N_7187,N_6643);
or U9198 (N_9198,N_7263,N_7888);
or U9199 (N_9199,N_7793,N_7078);
and U9200 (N_9200,N_6354,N_7965);
or U9201 (N_9201,N_7464,N_6199);
nand U9202 (N_9202,N_7984,N_6142);
xnor U9203 (N_9203,N_6455,N_7315);
or U9204 (N_9204,N_6269,N_7111);
nand U9205 (N_9205,N_7492,N_6605);
xor U9206 (N_9206,N_6110,N_6860);
and U9207 (N_9207,N_6989,N_7932);
and U9208 (N_9208,N_7265,N_7944);
or U9209 (N_9209,N_6450,N_7027);
nand U9210 (N_9210,N_6223,N_6468);
and U9211 (N_9211,N_6332,N_6737);
xnor U9212 (N_9212,N_6977,N_6550);
nor U9213 (N_9213,N_7633,N_6575);
nor U9214 (N_9214,N_7516,N_7622);
and U9215 (N_9215,N_6003,N_6831);
nor U9216 (N_9216,N_6596,N_6617);
xor U9217 (N_9217,N_7816,N_6604);
or U9218 (N_9218,N_6440,N_7812);
nand U9219 (N_9219,N_6556,N_6434);
and U9220 (N_9220,N_6224,N_6325);
and U9221 (N_9221,N_6339,N_6701);
nor U9222 (N_9222,N_7768,N_6785);
and U9223 (N_9223,N_7456,N_6246);
nor U9224 (N_9224,N_6157,N_6144);
or U9225 (N_9225,N_7025,N_7243);
xor U9226 (N_9226,N_6727,N_7545);
xor U9227 (N_9227,N_7675,N_7481);
and U9228 (N_9228,N_6267,N_7485);
nor U9229 (N_9229,N_7986,N_7176);
xor U9230 (N_9230,N_7946,N_7527);
nand U9231 (N_9231,N_6898,N_6203);
and U9232 (N_9232,N_7099,N_7459);
nor U9233 (N_9233,N_6618,N_7868);
nor U9234 (N_9234,N_6043,N_6998);
nand U9235 (N_9235,N_6245,N_6647);
or U9236 (N_9236,N_7921,N_6799);
or U9237 (N_9237,N_6043,N_7271);
or U9238 (N_9238,N_6869,N_6761);
or U9239 (N_9239,N_6400,N_7935);
xnor U9240 (N_9240,N_7253,N_6661);
and U9241 (N_9241,N_6945,N_7937);
nor U9242 (N_9242,N_6830,N_6100);
nor U9243 (N_9243,N_7441,N_7882);
nor U9244 (N_9244,N_7641,N_6032);
xor U9245 (N_9245,N_7302,N_7674);
xnor U9246 (N_9246,N_7487,N_7092);
nand U9247 (N_9247,N_7710,N_7541);
and U9248 (N_9248,N_6553,N_7684);
or U9249 (N_9249,N_6340,N_7824);
xor U9250 (N_9250,N_7208,N_6917);
and U9251 (N_9251,N_6777,N_7909);
or U9252 (N_9252,N_6867,N_7472);
or U9253 (N_9253,N_6011,N_7991);
nor U9254 (N_9254,N_6306,N_6734);
and U9255 (N_9255,N_7816,N_7764);
nand U9256 (N_9256,N_6074,N_6564);
and U9257 (N_9257,N_6018,N_7240);
or U9258 (N_9258,N_6219,N_6634);
and U9259 (N_9259,N_7706,N_7762);
xnor U9260 (N_9260,N_7204,N_7102);
nor U9261 (N_9261,N_7386,N_7303);
and U9262 (N_9262,N_7466,N_6273);
nand U9263 (N_9263,N_7904,N_6905);
xor U9264 (N_9264,N_6282,N_7875);
or U9265 (N_9265,N_7185,N_7968);
and U9266 (N_9266,N_6421,N_6078);
nor U9267 (N_9267,N_6890,N_7621);
or U9268 (N_9268,N_6906,N_7357);
and U9269 (N_9269,N_6376,N_6651);
nor U9270 (N_9270,N_6374,N_6510);
or U9271 (N_9271,N_6271,N_7069);
xor U9272 (N_9272,N_7933,N_6862);
xor U9273 (N_9273,N_7160,N_7962);
nor U9274 (N_9274,N_7313,N_6976);
nand U9275 (N_9275,N_6596,N_7386);
nand U9276 (N_9276,N_6639,N_7615);
nor U9277 (N_9277,N_6482,N_6337);
nand U9278 (N_9278,N_7691,N_7657);
xnor U9279 (N_9279,N_7191,N_6662);
xor U9280 (N_9280,N_7535,N_6391);
nand U9281 (N_9281,N_7043,N_6695);
nand U9282 (N_9282,N_7795,N_6781);
or U9283 (N_9283,N_6133,N_7198);
or U9284 (N_9284,N_6334,N_7705);
or U9285 (N_9285,N_7296,N_6974);
nand U9286 (N_9286,N_6904,N_6993);
nand U9287 (N_9287,N_6399,N_7734);
nand U9288 (N_9288,N_6928,N_6842);
nand U9289 (N_9289,N_7699,N_6424);
xnor U9290 (N_9290,N_6231,N_6397);
xor U9291 (N_9291,N_6309,N_6055);
and U9292 (N_9292,N_6245,N_6440);
and U9293 (N_9293,N_6585,N_6293);
nand U9294 (N_9294,N_6201,N_7295);
nor U9295 (N_9295,N_6073,N_7294);
nor U9296 (N_9296,N_6405,N_6439);
and U9297 (N_9297,N_6779,N_6174);
nand U9298 (N_9298,N_6452,N_6733);
nor U9299 (N_9299,N_6168,N_6623);
nor U9300 (N_9300,N_7149,N_7504);
and U9301 (N_9301,N_7469,N_6919);
and U9302 (N_9302,N_7782,N_6974);
nand U9303 (N_9303,N_6694,N_6299);
xor U9304 (N_9304,N_7492,N_7694);
or U9305 (N_9305,N_6383,N_7406);
xor U9306 (N_9306,N_7226,N_7564);
nand U9307 (N_9307,N_7722,N_7742);
nor U9308 (N_9308,N_6222,N_6486);
or U9309 (N_9309,N_7193,N_6522);
and U9310 (N_9310,N_7270,N_7114);
nor U9311 (N_9311,N_7016,N_7486);
nor U9312 (N_9312,N_6332,N_7441);
nand U9313 (N_9313,N_7121,N_6991);
nand U9314 (N_9314,N_7492,N_7857);
nand U9315 (N_9315,N_6561,N_7580);
nor U9316 (N_9316,N_6604,N_7691);
nand U9317 (N_9317,N_7322,N_7899);
nand U9318 (N_9318,N_6505,N_6858);
nand U9319 (N_9319,N_6340,N_7456);
or U9320 (N_9320,N_7496,N_7168);
nand U9321 (N_9321,N_7845,N_6106);
and U9322 (N_9322,N_6972,N_7240);
xor U9323 (N_9323,N_6232,N_6157);
and U9324 (N_9324,N_6962,N_6380);
nor U9325 (N_9325,N_6027,N_6599);
or U9326 (N_9326,N_7451,N_6750);
or U9327 (N_9327,N_7826,N_6962);
or U9328 (N_9328,N_7358,N_6218);
nand U9329 (N_9329,N_7972,N_7521);
nor U9330 (N_9330,N_6115,N_6395);
or U9331 (N_9331,N_6365,N_7147);
and U9332 (N_9332,N_7144,N_7462);
xor U9333 (N_9333,N_7944,N_7032);
xnor U9334 (N_9334,N_7468,N_7379);
xnor U9335 (N_9335,N_7879,N_7378);
or U9336 (N_9336,N_7932,N_7520);
nand U9337 (N_9337,N_6012,N_6804);
and U9338 (N_9338,N_7259,N_7341);
and U9339 (N_9339,N_6898,N_7918);
xnor U9340 (N_9340,N_6959,N_7918);
nand U9341 (N_9341,N_7046,N_6274);
or U9342 (N_9342,N_6789,N_7688);
nor U9343 (N_9343,N_6124,N_6558);
or U9344 (N_9344,N_7953,N_6156);
or U9345 (N_9345,N_6092,N_6310);
or U9346 (N_9346,N_6148,N_7231);
and U9347 (N_9347,N_7400,N_6764);
nand U9348 (N_9348,N_7770,N_6713);
nand U9349 (N_9349,N_6468,N_6797);
and U9350 (N_9350,N_6348,N_7623);
and U9351 (N_9351,N_7751,N_6454);
or U9352 (N_9352,N_6747,N_7827);
nand U9353 (N_9353,N_6532,N_6655);
nor U9354 (N_9354,N_7267,N_6806);
and U9355 (N_9355,N_6551,N_6143);
nor U9356 (N_9356,N_6123,N_6247);
nand U9357 (N_9357,N_6112,N_7808);
xor U9358 (N_9358,N_7797,N_7002);
nand U9359 (N_9359,N_7214,N_7023);
nand U9360 (N_9360,N_7889,N_6713);
and U9361 (N_9361,N_6965,N_6429);
xor U9362 (N_9362,N_7878,N_7702);
or U9363 (N_9363,N_7877,N_7799);
and U9364 (N_9364,N_7629,N_7110);
or U9365 (N_9365,N_7143,N_7369);
nor U9366 (N_9366,N_6230,N_7293);
xor U9367 (N_9367,N_7924,N_7695);
xor U9368 (N_9368,N_6140,N_6103);
nor U9369 (N_9369,N_7310,N_7117);
nand U9370 (N_9370,N_6273,N_7200);
and U9371 (N_9371,N_6303,N_7179);
and U9372 (N_9372,N_7050,N_6234);
nor U9373 (N_9373,N_6722,N_7034);
or U9374 (N_9374,N_6091,N_6733);
nand U9375 (N_9375,N_6350,N_6339);
nand U9376 (N_9376,N_6730,N_7429);
xor U9377 (N_9377,N_7423,N_6939);
or U9378 (N_9378,N_6208,N_6685);
xnor U9379 (N_9379,N_6657,N_7737);
and U9380 (N_9380,N_6411,N_6945);
xnor U9381 (N_9381,N_6698,N_6367);
and U9382 (N_9382,N_7215,N_6273);
xor U9383 (N_9383,N_6499,N_6906);
and U9384 (N_9384,N_6907,N_6220);
xor U9385 (N_9385,N_6760,N_7358);
nand U9386 (N_9386,N_6890,N_6307);
nand U9387 (N_9387,N_6403,N_6157);
xor U9388 (N_9388,N_7986,N_6069);
or U9389 (N_9389,N_6997,N_7925);
or U9390 (N_9390,N_6521,N_7359);
nor U9391 (N_9391,N_6964,N_6214);
or U9392 (N_9392,N_6653,N_7699);
nand U9393 (N_9393,N_7737,N_7647);
xnor U9394 (N_9394,N_7492,N_6013);
or U9395 (N_9395,N_7686,N_6553);
nor U9396 (N_9396,N_6107,N_6139);
xor U9397 (N_9397,N_7863,N_7070);
or U9398 (N_9398,N_6362,N_6336);
and U9399 (N_9399,N_7682,N_6120);
and U9400 (N_9400,N_6963,N_6342);
and U9401 (N_9401,N_7813,N_7072);
nor U9402 (N_9402,N_7895,N_6210);
and U9403 (N_9403,N_7457,N_6476);
xor U9404 (N_9404,N_7746,N_7910);
nand U9405 (N_9405,N_6523,N_7734);
and U9406 (N_9406,N_7524,N_6979);
or U9407 (N_9407,N_6376,N_7025);
nor U9408 (N_9408,N_7023,N_7364);
and U9409 (N_9409,N_6781,N_6964);
nor U9410 (N_9410,N_6173,N_7717);
xor U9411 (N_9411,N_7504,N_6843);
or U9412 (N_9412,N_6739,N_7335);
xor U9413 (N_9413,N_6158,N_6055);
or U9414 (N_9414,N_6891,N_6011);
nand U9415 (N_9415,N_6784,N_6447);
nand U9416 (N_9416,N_6178,N_7093);
xnor U9417 (N_9417,N_7714,N_7813);
or U9418 (N_9418,N_7684,N_6808);
or U9419 (N_9419,N_6535,N_7683);
xor U9420 (N_9420,N_7957,N_6865);
nor U9421 (N_9421,N_6521,N_7041);
or U9422 (N_9422,N_6677,N_6122);
and U9423 (N_9423,N_6569,N_7434);
or U9424 (N_9424,N_7823,N_6514);
or U9425 (N_9425,N_6051,N_6310);
nor U9426 (N_9426,N_6964,N_6530);
nand U9427 (N_9427,N_6702,N_7587);
xor U9428 (N_9428,N_6837,N_7320);
nand U9429 (N_9429,N_6717,N_6023);
xnor U9430 (N_9430,N_6550,N_7094);
nand U9431 (N_9431,N_6110,N_7451);
and U9432 (N_9432,N_7781,N_6995);
and U9433 (N_9433,N_6523,N_7384);
and U9434 (N_9434,N_7677,N_6252);
nor U9435 (N_9435,N_7230,N_6623);
xnor U9436 (N_9436,N_6646,N_6392);
nand U9437 (N_9437,N_6803,N_7897);
or U9438 (N_9438,N_6241,N_7829);
xor U9439 (N_9439,N_6596,N_6932);
and U9440 (N_9440,N_7687,N_7568);
or U9441 (N_9441,N_7406,N_6763);
nand U9442 (N_9442,N_6914,N_6513);
xor U9443 (N_9443,N_6977,N_7081);
nand U9444 (N_9444,N_7171,N_6055);
nor U9445 (N_9445,N_7215,N_6777);
nand U9446 (N_9446,N_6318,N_6898);
or U9447 (N_9447,N_6977,N_6911);
xnor U9448 (N_9448,N_7344,N_7702);
xnor U9449 (N_9449,N_6726,N_7830);
xor U9450 (N_9450,N_7147,N_6982);
or U9451 (N_9451,N_7397,N_6177);
and U9452 (N_9452,N_7061,N_6109);
nor U9453 (N_9453,N_6668,N_6162);
and U9454 (N_9454,N_6852,N_7555);
or U9455 (N_9455,N_6106,N_7321);
and U9456 (N_9456,N_7931,N_6341);
and U9457 (N_9457,N_6110,N_7611);
nor U9458 (N_9458,N_6172,N_6799);
or U9459 (N_9459,N_7174,N_6060);
nor U9460 (N_9460,N_6067,N_6409);
nor U9461 (N_9461,N_6387,N_7793);
and U9462 (N_9462,N_6007,N_7547);
nand U9463 (N_9463,N_6280,N_6312);
or U9464 (N_9464,N_7070,N_6205);
xnor U9465 (N_9465,N_7311,N_6207);
or U9466 (N_9466,N_7980,N_7371);
and U9467 (N_9467,N_7230,N_6249);
or U9468 (N_9468,N_7457,N_7888);
nand U9469 (N_9469,N_6770,N_6548);
nor U9470 (N_9470,N_6797,N_6169);
or U9471 (N_9471,N_6585,N_6840);
xor U9472 (N_9472,N_6339,N_6364);
or U9473 (N_9473,N_7089,N_6191);
nor U9474 (N_9474,N_7409,N_6226);
and U9475 (N_9475,N_7124,N_6855);
or U9476 (N_9476,N_6125,N_7728);
and U9477 (N_9477,N_7474,N_7736);
xnor U9478 (N_9478,N_6916,N_6575);
nand U9479 (N_9479,N_7534,N_7952);
or U9480 (N_9480,N_7397,N_6367);
or U9481 (N_9481,N_6176,N_6811);
or U9482 (N_9482,N_7072,N_7575);
and U9483 (N_9483,N_7733,N_7170);
and U9484 (N_9484,N_7256,N_6680);
and U9485 (N_9485,N_7755,N_6094);
nand U9486 (N_9486,N_7889,N_6315);
nor U9487 (N_9487,N_6207,N_7315);
nor U9488 (N_9488,N_7955,N_7810);
nor U9489 (N_9489,N_6855,N_6708);
nand U9490 (N_9490,N_7681,N_7182);
xnor U9491 (N_9491,N_6514,N_6934);
or U9492 (N_9492,N_6674,N_6673);
and U9493 (N_9493,N_7789,N_6695);
nor U9494 (N_9494,N_6883,N_6501);
and U9495 (N_9495,N_6864,N_7223);
nand U9496 (N_9496,N_6783,N_6274);
nor U9497 (N_9497,N_7710,N_7988);
nand U9498 (N_9498,N_7610,N_7034);
or U9499 (N_9499,N_6311,N_7480);
nor U9500 (N_9500,N_6180,N_7229);
nand U9501 (N_9501,N_7093,N_6856);
and U9502 (N_9502,N_6371,N_6826);
nor U9503 (N_9503,N_7153,N_6950);
and U9504 (N_9504,N_7195,N_7155);
nor U9505 (N_9505,N_7017,N_6445);
xnor U9506 (N_9506,N_6741,N_6179);
xor U9507 (N_9507,N_6934,N_6012);
or U9508 (N_9508,N_7091,N_6158);
nand U9509 (N_9509,N_6810,N_6578);
and U9510 (N_9510,N_7393,N_7350);
nor U9511 (N_9511,N_7107,N_6204);
nor U9512 (N_9512,N_7745,N_7308);
xnor U9513 (N_9513,N_7069,N_7578);
nor U9514 (N_9514,N_7202,N_7555);
xor U9515 (N_9515,N_6105,N_7793);
nor U9516 (N_9516,N_7991,N_7780);
nand U9517 (N_9517,N_6322,N_7815);
nor U9518 (N_9518,N_6710,N_7083);
or U9519 (N_9519,N_7599,N_7983);
and U9520 (N_9520,N_6073,N_6219);
or U9521 (N_9521,N_6351,N_7028);
nor U9522 (N_9522,N_7776,N_7331);
nor U9523 (N_9523,N_6306,N_6974);
and U9524 (N_9524,N_6559,N_6405);
and U9525 (N_9525,N_6626,N_7458);
nor U9526 (N_9526,N_7634,N_7461);
or U9527 (N_9527,N_7343,N_7604);
or U9528 (N_9528,N_7267,N_7103);
or U9529 (N_9529,N_6545,N_6813);
or U9530 (N_9530,N_7988,N_7838);
nor U9531 (N_9531,N_7022,N_6727);
nor U9532 (N_9532,N_7178,N_6978);
nor U9533 (N_9533,N_7401,N_7605);
nand U9534 (N_9534,N_6012,N_6766);
xnor U9535 (N_9535,N_6793,N_7851);
nand U9536 (N_9536,N_6997,N_7855);
or U9537 (N_9537,N_6802,N_7343);
and U9538 (N_9538,N_7266,N_7581);
or U9539 (N_9539,N_7038,N_7020);
xnor U9540 (N_9540,N_6161,N_6305);
nand U9541 (N_9541,N_6484,N_7863);
xor U9542 (N_9542,N_6625,N_6174);
or U9543 (N_9543,N_6429,N_6336);
nor U9544 (N_9544,N_6477,N_7133);
or U9545 (N_9545,N_7241,N_6889);
nor U9546 (N_9546,N_7623,N_7913);
or U9547 (N_9547,N_7835,N_7335);
xnor U9548 (N_9548,N_6743,N_7606);
nor U9549 (N_9549,N_7916,N_6660);
or U9550 (N_9550,N_7916,N_6622);
or U9551 (N_9551,N_6259,N_6134);
or U9552 (N_9552,N_6760,N_7633);
or U9553 (N_9553,N_6456,N_7325);
nor U9554 (N_9554,N_6613,N_7031);
nand U9555 (N_9555,N_7473,N_6432);
nor U9556 (N_9556,N_7233,N_6976);
and U9557 (N_9557,N_7250,N_7478);
nor U9558 (N_9558,N_6162,N_6083);
or U9559 (N_9559,N_6587,N_7642);
nor U9560 (N_9560,N_6421,N_6210);
nor U9561 (N_9561,N_7010,N_6787);
xnor U9562 (N_9562,N_7941,N_6878);
nor U9563 (N_9563,N_7923,N_6654);
nand U9564 (N_9564,N_6648,N_6797);
xnor U9565 (N_9565,N_7317,N_7343);
and U9566 (N_9566,N_7661,N_6377);
and U9567 (N_9567,N_6800,N_6204);
and U9568 (N_9568,N_7047,N_7276);
nor U9569 (N_9569,N_6170,N_6393);
xnor U9570 (N_9570,N_7250,N_7808);
and U9571 (N_9571,N_6143,N_7518);
and U9572 (N_9572,N_7120,N_7784);
and U9573 (N_9573,N_6243,N_6835);
or U9574 (N_9574,N_7813,N_6225);
nand U9575 (N_9575,N_7515,N_6206);
nand U9576 (N_9576,N_7034,N_7062);
and U9577 (N_9577,N_7011,N_7000);
nor U9578 (N_9578,N_7930,N_6533);
or U9579 (N_9579,N_6010,N_6837);
xor U9580 (N_9580,N_6972,N_6189);
nor U9581 (N_9581,N_6326,N_7011);
nand U9582 (N_9582,N_7084,N_7123);
nand U9583 (N_9583,N_6723,N_7318);
xor U9584 (N_9584,N_6880,N_6586);
xnor U9585 (N_9585,N_7941,N_7865);
nor U9586 (N_9586,N_6222,N_7504);
and U9587 (N_9587,N_7570,N_7806);
xnor U9588 (N_9588,N_6578,N_6710);
and U9589 (N_9589,N_6818,N_7180);
and U9590 (N_9590,N_7896,N_6339);
nand U9591 (N_9591,N_7785,N_6362);
or U9592 (N_9592,N_7451,N_7085);
or U9593 (N_9593,N_7186,N_7594);
nor U9594 (N_9594,N_6998,N_6973);
or U9595 (N_9595,N_7710,N_6226);
nand U9596 (N_9596,N_7880,N_6036);
and U9597 (N_9597,N_6585,N_6275);
nor U9598 (N_9598,N_7905,N_6097);
xnor U9599 (N_9599,N_7552,N_6240);
and U9600 (N_9600,N_7027,N_6203);
nand U9601 (N_9601,N_7313,N_6633);
nor U9602 (N_9602,N_7439,N_6417);
nor U9603 (N_9603,N_6796,N_7635);
nor U9604 (N_9604,N_7871,N_7968);
and U9605 (N_9605,N_7905,N_7953);
nor U9606 (N_9606,N_6083,N_7714);
nor U9607 (N_9607,N_7268,N_7170);
nor U9608 (N_9608,N_7136,N_7302);
nor U9609 (N_9609,N_6494,N_7484);
and U9610 (N_9610,N_6076,N_7367);
nand U9611 (N_9611,N_7797,N_6546);
nor U9612 (N_9612,N_7996,N_7302);
or U9613 (N_9613,N_7128,N_7019);
nor U9614 (N_9614,N_6508,N_7840);
xnor U9615 (N_9615,N_7639,N_7574);
nor U9616 (N_9616,N_6293,N_7037);
and U9617 (N_9617,N_7095,N_6001);
nor U9618 (N_9618,N_6000,N_7154);
and U9619 (N_9619,N_7166,N_7268);
and U9620 (N_9620,N_6232,N_6736);
or U9621 (N_9621,N_7016,N_6588);
and U9622 (N_9622,N_6636,N_6325);
and U9623 (N_9623,N_6765,N_7920);
nor U9624 (N_9624,N_6639,N_7370);
nor U9625 (N_9625,N_7101,N_6996);
nor U9626 (N_9626,N_7240,N_6098);
and U9627 (N_9627,N_6777,N_7972);
xnor U9628 (N_9628,N_7804,N_7271);
xnor U9629 (N_9629,N_6239,N_6642);
and U9630 (N_9630,N_7127,N_7661);
nand U9631 (N_9631,N_6854,N_6986);
and U9632 (N_9632,N_6900,N_7430);
nor U9633 (N_9633,N_7090,N_6065);
or U9634 (N_9634,N_7847,N_6773);
nand U9635 (N_9635,N_7201,N_7780);
nand U9636 (N_9636,N_7032,N_6344);
nand U9637 (N_9637,N_7737,N_6082);
nor U9638 (N_9638,N_7661,N_7833);
nor U9639 (N_9639,N_6287,N_6359);
xor U9640 (N_9640,N_6449,N_7124);
or U9641 (N_9641,N_7671,N_7621);
and U9642 (N_9642,N_6094,N_7677);
xor U9643 (N_9643,N_7517,N_6761);
nor U9644 (N_9644,N_6097,N_6283);
xor U9645 (N_9645,N_7585,N_6636);
nand U9646 (N_9646,N_6208,N_7731);
or U9647 (N_9647,N_7526,N_7716);
and U9648 (N_9648,N_6109,N_7367);
nor U9649 (N_9649,N_7413,N_6408);
nand U9650 (N_9650,N_6729,N_6492);
xnor U9651 (N_9651,N_7455,N_7009);
xor U9652 (N_9652,N_7222,N_7289);
xor U9653 (N_9653,N_7759,N_7047);
xor U9654 (N_9654,N_7581,N_7172);
nand U9655 (N_9655,N_7554,N_6470);
nand U9656 (N_9656,N_6789,N_7839);
nor U9657 (N_9657,N_7267,N_6541);
nor U9658 (N_9658,N_7273,N_6691);
nand U9659 (N_9659,N_7775,N_6454);
xnor U9660 (N_9660,N_6448,N_6357);
nor U9661 (N_9661,N_6748,N_6089);
and U9662 (N_9662,N_7540,N_6127);
or U9663 (N_9663,N_6088,N_6541);
or U9664 (N_9664,N_6010,N_6806);
nand U9665 (N_9665,N_7918,N_6335);
and U9666 (N_9666,N_6315,N_6834);
nand U9667 (N_9667,N_6932,N_7347);
or U9668 (N_9668,N_6689,N_7622);
nor U9669 (N_9669,N_6677,N_7559);
nand U9670 (N_9670,N_7345,N_6060);
or U9671 (N_9671,N_7646,N_7874);
or U9672 (N_9672,N_6831,N_7333);
and U9673 (N_9673,N_7794,N_6792);
or U9674 (N_9674,N_6065,N_7372);
or U9675 (N_9675,N_7381,N_7706);
or U9676 (N_9676,N_6477,N_7614);
nand U9677 (N_9677,N_6510,N_6880);
nand U9678 (N_9678,N_7318,N_7513);
nor U9679 (N_9679,N_7453,N_7698);
and U9680 (N_9680,N_7378,N_7673);
and U9681 (N_9681,N_7664,N_7278);
xnor U9682 (N_9682,N_6470,N_6679);
or U9683 (N_9683,N_7188,N_7256);
and U9684 (N_9684,N_7177,N_6273);
nand U9685 (N_9685,N_7787,N_6714);
xnor U9686 (N_9686,N_7337,N_6079);
and U9687 (N_9687,N_7129,N_6718);
xnor U9688 (N_9688,N_7406,N_7394);
nor U9689 (N_9689,N_6891,N_7551);
xnor U9690 (N_9690,N_6255,N_6632);
or U9691 (N_9691,N_7457,N_7167);
nor U9692 (N_9692,N_7917,N_6780);
or U9693 (N_9693,N_6184,N_6196);
or U9694 (N_9694,N_6524,N_7441);
nor U9695 (N_9695,N_6192,N_6008);
xnor U9696 (N_9696,N_7171,N_6965);
xor U9697 (N_9697,N_7468,N_7149);
xor U9698 (N_9698,N_7992,N_6563);
nand U9699 (N_9699,N_7836,N_7981);
xor U9700 (N_9700,N_6009,N_7640);
nor U9701 (N_9701,N_6941,N_7310);
nand U9702 (N_9702,N_6517,N_7667);
nand U9703 (N_9703,N_7100,N_6701);
xor U9704 (N_9704,N_7139,N_7499);
xor U9705 (N_9705,N_6271,N_6999);
xnor U9706 (N_9706,N_7165,N_6679);
xnor U9707 (N_9707,N_6648,N_7580);
nor U9708 (N_9708,N_6163,N_7523);
or U9709 (N_9709,N_6473,N_7723);
or U9710 (N_9710,N_6763,N_6262);
and U9711 (N_9711,N_7724,N_7227);
and U9712 (N_9712,N_6203,N_6321);
xor U9713 (N_9713,N_6075,N_6997);
xnor U9714 (N_9714,N_7217,N_6849);
and U9715 (N_9715,N_7752,N_6434);
and U9716 (N_9716,N_7294,N_7605);
nor U9717 (N_9717,N_6987,N_7901);
nor U9718 (N_9718,N_6961,N_6159);
nand U9719 (N_9719,N_6179,N_7118);
or U9720 (N_9720,N_7799,N_6556);
or U9721 (N_9721,N_6312,N_6760);
nor U9722 (N_9722,N_6906,N_7596);
xor U9723 (N_9723,N_6967,N_7838);
and U9724 (N_9724,N_6890,N_7542);
nor U9725 (N_9725,N_7845,N_6477);
and U9726 (N_9726,N_6675,N_6363);
nand U9727 (N_9727,N_6154,N_7414);
or U9728 (N_9728,N_6032,N_7114);
nor U9729 (N_9729,N_6374,N_6326);
and U9730 (N_9730,N_6263,N_6158);
nor U9731 (N_9731,N_6888,N_6909);
and U9732 (N_9732,N_7725,N_7819);
or U9733 (N_9733,N_6008,N_6716);
nor U9734 (N_9734,N_6709,N_6820);
nor U9735 (N_9735,N_6796,N_6670);
xnor U9736 (N_9736,N_7357,N_7655);
xnor U9737 (N_9737,N_7473,N_7458);
nand U9738 (N_9738,N_7492,N_7007);
and U9739 (N_9739,N_6762,N_7161);
and U9740 (N_9740,N_6286,N_7931);
and U9741 (N_9741,N_6710,N_7794);
xnor U9742 (N_9742,N_6906,N_7872);
nor U9743 (N_9743,N_6061,N_6317);
nor U9744 (N_9744,N_7948,N_7670);
xor U9745 (N_9745,N_7429,N_7921);
xnor U9746 (N_9746,N_6900,N_7137);
or U9747 (N_9747,N_6436,N_7607);
and U9748 (N_9748,N_6365,N_7017);
xnor U9749 (N_9749,N_6191,N_7568);
nand U9750 (N_9750,N_6760,N_6885);
or U9751 (N_9751,N_7150,N_7961);
or U9752 (N_9752,N_6080,N_7562);
xor U9753 (N_9753,N_6979,N_6052);
or U9754 (N_9754,N_7814,N_6799);
nand U9755 (N_9755,N_7821,N_6334);
nor U9756 (N_9756,N_6103,N_7347);
xnor U9757 (N_9757,N_7329,N_6048);
nor U9758 (N_9758,N_6844,N_7763);
xor U9759 (N_9759,N_6341,N_6627);
and U9760 (N_9760,N_7012,N_7613);
or U9761 (N_9761,N_6008,N_6667);
or U9762 (N_9762,N_7032,N_6156);
nor U9763 (N_9763,N_6478,N_6314);
or U9764 (N_9764,N_7607,N_7258);
nor U9765 (N_9765,N_7339,N_7294);
nand U9766 (N_9766,N_7608,N_6765);
and U9767 (N_9767,N_6412,N_7784);
xor U9768 (N_9768,N_6841,N_6093);
xnor U9769 (N_9769,N_6731,N_7011);
xor U9770 (N_9770,N_7215,N_6969);
and U9771 (N_9771,N_6469,N_7310);
and U9772 (N_9772,N_6989,N_7060);
nor U9773 (N_9773,N_6320,N_7972);
xnor U9774 (N_9774,N_7222,N_6941);
xor U9775 (N_9775,N_7475,N_7538);
and U9776 (N_9776,N_7492,N_6789);
nand U9777 (N_9777,N_6258,N_6586);
xnor U9778 (N_9778,N_7306,N_7402);
xnor U9779 (N_9779,N_6988,N_6688);
or U9780 (N_9780,N_6889,N_7757);
nand U9781 (N_9781,N_6518,N_7070);
xnor U9782 (N_9782,N_6555,N_7161);
or U9783 (N_9783,N_7307,N_7623);
nand U9784 (N_9784,N_7510,N_7063);
or U9785 (N_9785,N_6349,N_6999);
xor U9786 (N_9786,N_7360,N_6021);
and U9787 (N_9787,N_6346,N_7740);
nor U9788 (N_9788,N_7674,N_7292);
or U9789 (N_9789,N_6806,N_7304);
xor U9790 (N_9790,N_7978,N_6516);
xor U9791 (N_9791,N_7706,N_7672);
or U9792 (N_9792,N_7302,N_6910);
nand U9793 (N_9793,N_7957,N_6952);
or U9794 (N_9794,N_6292,N_6977);
nand U9795 (N_9795,N_7837,N_6931);
nand U9796 (N_9796,N_7422,N_7356);
and U9797 (N_9797,N_7253,N_7735);
or U9798 (N_9798,N_6060,N_6262);
xnor U9799 (N_9799,N_6880,N_6902);
xnor U9800 (N_9800,N_6575,N_6962);
xor U9801 (N_9801,N_7577,N_7118);
xnor U9802 (N_9802,N_6641,N_7611);
nor U9803 (N_9803,N_7492,N_7842);
and U9804 (N_9804,N_6322,N_6504);
xnor U9805 (N_9805,N_7154,N_7298);
nor U9806 (N_9806,N_6907,N_6206);
or U9807 (N_9807,N_6717,N_7512);
or U9808 (N_9808,N_7729,N_6897);
nor U9809 (N_9809,N_7209,N_7362);
or U9810 (N_9810,N_7689,N_6243);
xnor U9811 (N_9811,N_6703,N_7338);
and U9812 (N_9812,N_6722,N_6897);
or U9813 (N_9813,N_6550,N_7185);
and U9814 (N_9814,N_6845,N_6205);
xor U9815 (N_9815,N_7655,N_6731);
nand U9816 (N_9816,N_7141,N_6497);
or U9817 (N_9817,N_7523,N_6980);
and U9818 (N_9818,N_6943,N_7177);
and U9819 (N_9819,N_6014,N_7808);
xor U9820 (N_9820,N_6787,N_7951);
xnor U9821 (N_9821,N_6708,N_6558);
or U9822 (N_9822,N_6576,N_6637);
nand U9823 (N_9823,N_6551,N_7560);
nand U9824 (N_9824,N_6577,N_7244);
or U9825 (N_9825,N_6831,N_6707);
nand U9826 (N_9826,N_7107,N_6241);
or U9827 (N_9827,N_7949,N_6673);
nand U9828 (N_9828,N_6769,N_7724);
and U9829 (N_9829,N_6577,N_7081);
nand U9830 (N_9830,N_7600,N_7431);
xnor U9831 (N_9831,N_7320,N_6292);
or U9832 (N_9832,N_7930,N_6893);
and U9833 (N_9833,N_6975,N_6730);
xor U9834 (N_9834,N_6531,N_6773);
nor U9835 (N_9835,N_7912,N_6263);
and U9836 (N_9836,N_6862,N_7147);
xnor U9837 (N_9837,N_6072,N_6294);
nand U9838 (N_9838,N_7530,N_6090);
nand U9839 (N_9839,N_7460,N_7905);
nand U9840 (N_9840,N_7466,N_7148);
or U9841 (N_9841,N_7549,N_6382);
nor U9842 (N_9842,N_7350,N_6787);
nor U9843 (N_9843,N_7920,N_7368);
and U9844 (N_9844,N_6927,N_7098);
nor U9845 (N_9845,N_6403,N_6610);
nand U9846 (N_9846,N_6938,N_6570);
or U9847 (N_9847,N_7536,N_7179);
nand U9848 (N_9848,N_6263,N_6294);
xnor U9849 (N_9849,N_7524,N_6813);
nor U9850 (N_9850,N_7047,N_7316);
xnor U9851 (N_9851,N_7772,N_7364);
and U9852 (N_9852,N_6931,N_7998);
nand U9853 (N_9853,N_7213,N_7896);
nor U9854 (N_9854,N_7918,N_6041);
nand U9855 (N_9855,N_7322,N_6801);
nor U9856 (N_9856,N_6358,N_6429);
xor U9857 (N_9857,N_7953,N_6300);
or U9858 (N_9858,N_7760,N_7804);
or U9859 (N_9859,N_6828,N_6926);
and U9860 (N_9860,N_6373,N_6228);
nand U9861 (N_9861,N_6348,N_6287);
and U9862 (N_9862,N_7942,N_7151);
or U9863 (N_9863,N_7671,N_7576);
or U9864 (N_9864,N_6607,N_7686);
or U9865 (N_9865,N_6657,N_6844);
xor U9866 (N_9866,N_6364,N_6411);
nand U9867 (N_9867,N_6814,N_6588);
and U9868 (N_9868,N_7876,N_6599);
nor U9869 (N_9869,N_6307,N_7613);
nor U9870 (N_9870,N_7650,N_6948);
nand U9871 (N_9871,N_6651,N_7279);
nand U9872 (N_9872,N_7891,N_7980);
xor U9873 (N_9873,N_6202,N_7283);
nor U9874 (N_9874,N_7399,N_7831);
nand U9875 (N_9875,N_6963,N_6147);
nand U9876 (N_9876,N_7003,N_6875);
nor U9877 (N_9877,N_6619,N_7410);
or U9878 (N_9878,N_6522,N_6791);
nand U9879 (N_9879,N_6826,N_6438);
nand U9880 (N_9880,N_7369,N_7434);
and U9881 (N_9881,N_7259,N_7523);
nand U9882 (N_9882,N_6096,N_7646);
nor U9883 (N_9883,N_6110,N_6663);
or U9884 (N_9884,N_7183,N_7777);
or U9885 (N_9885,N_7725,N_7381);
and U9886 (N_9886,N_7099,N_6891);
xor U9887 (N_9887,N_6956,N_7876);
nor U9888 (N_9888,N_6462,N_7963);
nand U9889 (N_9889,N_7320,N_6281);
nor U9890 (N_9890,N_6267,N_7413);
nand U9891 (N_9891,N_6917,N_7275);
xor U9892 (N_9892,N_6565,N_6525);
or U9893 (N_9893,N_6855,N_7283);
nand U9894 (N_9894,N_7297,N_7079);
xnor U9895 (N_9895,N_7661,N_7815);
and U9896 (N_9896,N_6612,N_6734);
nand U9897 (N_9897,N_6427,N_6139);
xor U9898 (N_9898,N_7936,N_6479);
nor U9899 (N_9899,N_7274,N_6558);
and U9900 (N_9900,N_6988,N_6721);
nor U9901 (N_9901,N_7022,N_6600);
nand U9902 (N_9902,N_7572,N_7060);
xor U9903 (N_9903,N_6015,N_6543);
and U9904 (N_9904,N_6342,N_7446);
and U9905 (N_9905,N_7329,N_7778);
xnor U9906 (N_9906,N_6662,N_7475);
xor U9907 (N_9907,N_6967,N_6389);
and U9908 (N_9908,N_7466,N_6813);
nand U9909 (N_9909,N_7462,N_6819);
nor U9910 (N_9910,N_7695,N_7943);
nand U9911 (N_9911,N_7845,N_7101);
and U9912 (N_9912,N_7212,N_6080);
xor U9913 (N_9913,N_6231,N_7491);
nand U9914 (N_9914,N_7677,N_6284);
nand U9915 (N_9915,N_6865,N_7262);
xor U9916 (N_9916,N_7249,N_7179);
nand U9917 (N_9917,N_7239,N_7278);
nor U9918 (N_9918,N_7875,N_6375);
or U9919 (N_9919,N_7114,N_7838);
nor U9920 (N_9920,N_7416,N_6546);
nor U9921 (N_9921,N_6875,N_6359);
nor U9922 (N_9922,N_7143,N_6172);
nor U9923 (N_9923,N_7257,N_7762);
or U9924 (N_9924,N_6844,N_6062);
xnor U9925 (N_9925,N_6979,N_7707);
or U9926 (N_9926,N_6128,N_6997);
and U9927 (N_9927,N_6514,N_7535);
and U9928 (N_9928,N_6879,N_7354);
xor U9929 (N_9929,N_6273,N_6244);
nor U9930 (N_9930,N_6409,N_7976);
and U9931 (N_9931,N_6699,N_6535);
nand U9932 (N_9932,N_6166,N_7491);
xor U9933 (N_9933,N_6693,N_7529);
nand U9934 (N_9934,N_6487,N_6237);
nor U9935 (N_9935,N_7913,N_6935);
xnor U9936 (N_9936,N_7176,N_7687);
and U9937 (N_9937,N_6784,N_7474);
xnor U9938 (N_9938,N_6582,N_7762);
nand U9939 (N_9939,N_7405,N_7941);
or U9940 (N_9940,N_7429,N_7330);
xor U9941 (N_9941,N_7427,N_6626);
xor U9942 (N_9942,N_7771,N_7471);
xor U9943 (N_9943,N_6685,N_6012);
xor U9944 (N_9944,N_6394,N_6375);
or U9945 (N_9945,N_6802,N_7415);
xnor U9946 (N_9946,N_6289,N_6009);
xor U9947 (N_9947,N_6960,N_7065);
nand U9948 (N_9948,N_6512,N_6867);
or U9949 (N_9949,N_6480,N_6890);
and U9950 (N_9950,N_6566,N_6466);
xnor U9951 (N_9951,N_6814,N_7863);
nand U9952 (N_9952,N_7926,N_7482);
nand U9953 (N_9953,N_6595,N_6829);
and U9954 (N_9954,N_6304,N_7268);
and U9955 (N_9955,N_7485,N_7348);
nand U9956 (N_9956,N_6134,N_7755);
and U9957 (N_9957,N_7913,N_7979);
or U9958 (N_9958,N_7214,N_6523);
nor U9959 (N_9959,N_6158,N_7578);
nand U9960 (N_9960,N_6489,N_6771);
nor U9961 (N_9961,N_6498,N_6936);
xor U9962 (N_9962,N_6141,N_6623);
and U9963 (N_9963,N_6728,N_6321);
or U9964 (N_9964,N_7586,N_6985);
and U9965 (N_9965,N_6299,N_7912);
and U9966 (N_9966,N_6119,N_7375);
and U9967 (N_9967,N_6224,N_7921);
nor U9968 (N_9968,N_6798,N_6652);
nand U9969 (N_9969,N_7986,N_7230);
nand U9970 (N_9970,N_7538,N_7217);
nor U9971 (N_9971,N_6806,N_7379);
or U9972 (N_9972,N_6167,N_6037);
nand U9973 (N_9973,N_7506,N_6946);
nor U9974 (N_9974,N_7394,N_7279);
and U9975 (N_9975,N_6156,N_6783);
and U9976 (N_9976,N_6168,N_6086);
xor U9977 (N_9977,N_6369,N_6609);
xnor U9978 (N_9978,N_6708,N_7404);
and U9979 (N_9979,N_6839,N_6911);
or U9980 (N_9980,N_7764,N_6032);
and U9981 (N_9981,N_6492,N_6426);
or U9982 (N_9982,N_6387,N_7719);
xnor U9983 (N_9983,N_7017,N_6076);
xnor U9984 (N_9984,N_6500,N_7317);
nor U9985 (N_9985,N_7986,N_6176);
xnor U9986 (N_9986,N_6528,N_6504);
xnor U9987 (N_9987,N_7168,N_6344);
xnor U9988 (N_9988,N_7280,N_7844);
or U9989 (N_9989,N_6118,N_6764);
and U9990 (N_9990,N_7071,N_7245);
or U9991 (N_9991,N_6927,N_7187);
xnor U9992 (N_9992,N_7306,N_6083);
and U9993 (N_9993,N_7761,N_6072);
and U9994 (N_9994,N_7892,N_6090);
xor U9995 (N_9995,N_6634,N_6232);
or U9996 (N_9996,N_7768,N_7149);
or U9997 (N_9997,N_6573,N_6926);
nor U9998 (N_9998,N_7417,N_7731);
xor U9999 (N_9999,N_7032,N_6807);
nand U10000 (N_10000,N_9529,N_8630);
or U10001 (N_10001,N_8585,N_9210);
nand U10002 (N_10002,N_9813,N_9908);
nor U10003 (N_10003,N_8123,N_9670);
nand U10004 (N_10004,N_9165,N_9414);
xor U10005 (N_10005,N_8328,N_9890);
nor U10006 (N_10006,N_9798,N_9889);
and U10007 (N_10007,N_8834,N_9751);
and U10008 (N_10008,N_9239,N_8467);
or U10009 (N_10009,N_9115,N_9107);
and U10010 (N_10010,N_8959,N_8498);
nor U10011 (N_10011,N_9486,N_8015);
and U10012 (N_10012,N_8295,N_9953);
xnor U10013 (N_10013,N_8455,N_9055);
nor U10014 (N_10014,N_9278,N_9979);
xnor U10015 (N_10015,N_8790,N_8235);
or U10016 (N_10016,N_8872,N_8896);
or U10017 (N_10017,N_8779,N_9647);
nor U10018 (N_10018,N_8196,N_8035);
xor U10019 (N_10019,N_8424,N_8122);
and U10020 (N_10020,N_8603,N_9638);
nand U10021 (N_10021,N_8836,N_8821);
nand U10022 (N_10022,N_8373,N_8485);
or U10023 (N_10023,N_9657,N_8823);
and U10024 (N_10024,N_9745,N_9731);
or U10025 (N_10025,N_9044,N_9807);
nand U10026 (N_10026,N_9926,N_8215);
and U10027 (N_10027,N_9472,N_9284);
nor U10028 (N_10028,N_8162,N_9212);
or U10029 (N_10029,N_9723,N_8155);
and U10030 (N_10030,N_8513,N_9738);
nor U10031 (N_10031,N_9223,N_9185);
nand U10032 (N_10032,N_9648,N_9821);
nor U10033 (N_10033,N_9942,N_9873);
nand U10034 (N_10034,N_9131,N_9976);
and U10035 (N_10035,N_9563,N_9999);
xnor U10036 (N_10036,N_8338,N_8711);
nor U10037 (N_10037,N_8597,N_8897);
and U10038 (N_10038,N_8282,N_9279);
or U10039 (N_10039,N_9915,N_8465);
and U10040 (N_10040,N_9987,N_9154);
and U10041 (N_10041,N_9329,N_9835);
or U10042 (N_10042,N_8783,N_9511);
and U10043 (N_10043,N_8565,N_8631);
xnor U10044 (N_10044,N_9629,N_8146);
and U10045 (N_10045,N_8687,N_8919);
nor U10046 (N_10046,N_9346,N_8780);
and U10047 (N_10047,N_9124,N_8535);
and U10048 (N_10048,N_8331,N_8170);
xor U10049 (N_10049,N_8178,N_8406);
xor U10050 (N_10050,N_8875,N_8322);
and U10051 (N_10051,N_9301,N_8618);
nor U10052 (N_10052,N_8357,N_8566);
xnor U10053 (N_10053,N_8911,N_9056);
and U10054 (N_10054,N_8641,N_9392);
or U10055 (N_10055,N_8871,N_8806);
or U10056 (N_10056,N_9224,N_8494);
nand U10057 (N_10057,N_8008,N_9431);
or U10058 (N_10058,N_9098,N_9747);
nor U10059 (N_10059,N_9378,N_9149);
xor U10060 (N_10060,N_8868,N_9737);
nand U10061 (N_10061,N_8407,N_9029);
nor U10062 (N_10062,N_9537,N_8450);
nand U10063 (N_10063,N_8412,N_9959);
xnor U10064 (N_10064,N_9352,N_8829);
xnor U10065 (N_10065,N_9000,N_8642);
nor U10066 (N_10066,N_8085,N_8231);
nor U10067 (N_10067,N_8564,N_9060);
nor U10068 (N_10068,N_8093,N_9121);
or U10069 (N_10069,N_8058,N_9847);
xor U10070 (N_10070,N_9535,N_9401);
nand U10071 (N_10071,N_8507,N_9887);
nand U10072 (N_10072,N_9317,N_9675);
nand U10073 (N_10073,N_8081,N_9335);
and U10074 (N_10074,N_8908,N_8405);
xnor U10075 (N_10075,N_8510,N_8608);
and U10076 (N_10076,N_8588,N_8761);
nand U10077 (N_10077,N_8057,N_8975);
and U10078 (N_10078,N_9272,N_9138);
xor U10079 (N_10079,N_9885,N_8901);
xnor U10080 (N_10080,N_9422,N_9031);
and U10081 (N_10081,N_8137,N_9856);
xnor U10082 (N_10082,N_9299,N_9480);
and U10083 (N_10083,N_8425,N_9554);
nand U10084 (N_10084,N_8249,N_9771);
xor U10085 (N_10085,N_8429,N_8804);
or U10086 (N_10086,N_8101,N_9664);
xnor U10087 (N_10087,N_8145,N_9226);
nand U10088 (N_10088,N_8402,N_8963);
or U10089 (N_10089,N_9998,N_9957);
xnor U10090 (N_10090,N_8052,N_8175);
and U10091 (N_10091,N_9153,N_9586);
and U10092 (N_10092,N_8973,N_8173);
and U10093 (N_10093,N_8371,N_9386);
nor U10094 (N_10094,N_8278,N_8277);
xnor U10095 (N_10095,N_9892,N_8822);
nor U10096 (N_10096,N_9052,N_8578);
nand U10097 (N_10097,N_8515,N_9155);
and U10098 (N_10098,N_8299,N_9313);
xnor U10099 (N_10099,N_8891,N_9285);
or U10100 (N_10100,N_8443,N_8289);
or U10101 (N_10101,N_8595,N_8300);
xor U10102 (N_10102,N_8064,N_8795);
nor U10103 (N_10103,N_9610,N_9303);
xnor U10104 (N_10104,N_8408,N_8388);
nor U10105 (N_10105,N_8700,N_9420);
or U10106 (N_10106,N_8726,N_8643);
nand U10107 (N_10107,N_9742,N_8359);
nand U10108 (N_10108,N_8898,N_9007);
xor U10109 (N_10109,N_8041,N_9429);
or U10110 (N_10110,N_9250,N_8877);
nor U10111 (N_10111,N_8020,N_9377);
xnor U10112 (N_10112,N_8210,N_9974);
nor U10113 (N_10113,N_9775,N_8153);
or U10114 (N_10114,N_8023,N_9699);
xor U10115 (N_10115,N_8130,N_8718);
nand U10116 (N_10116,N_9577,N_8344);
nand U10117 (N_10117,N_8675,N_9514);
or U10118 (N_10118,N_9050,N_8801);
xnor U10119 (N_10119,N_9641,N_8022);
xor U10120 (N_10120,N_8813,N_8941);
or U10121 (N_10121,N_9411,N_8421);
and U10122 (N_10122,N_9013,N_8342);
nor U10123 (N_10123,N_8204,N_9904);
and U10124 (N_10124,N_8715,N_8915);
or U10125 (N_10125,N_8698,N_9615);
and U10126 (N_10126,N_8870,N_9321);
xnor U10127 (N_10127,N_8648,N_9178);
or U10128 (N_10128,N_8523,N_8923);
or U10129 (N_10129,N_8842,N_8982);
and U10130 (N_10130,N_8548,N_9515);
or U10131 (N_10131,N_8014,N_9839);
nand U10132 (N_10132,N_9366,N_8541);
or U10133 (N_10133,N_9937,N_8593);
nand U10134 (N_10134,N_8308,N_9820);
and U10135 (N_10135,N_9300,N_8283);
or U10136 (N_10136,N_8600,N_8389);
nor U10137 (N_10137,N_8119,N_8841);
xor U10138 (N_10138,N_8094,N_9799);
nor U10139 (N_10139,N_8759,N_9273);
or U10140 (N_10140,N_8219,N_9427);
nor U10141 (N_10141,N_8066,N_8894);
xor U10142 (N_10142,N_9085,N_9071);
nor U10143 (N_10143,N_9528,N_8934);
nor U10144 (N_10144,N_8659,N_9814);
and U10145 (N_10145,N_9965,N_8887);
nor U10146 (N_10146,N_8361,N_9543);
or U10147 (N_10147,N_8457,N_8781);
nand U10148 (N_10148,N_8247,N_9195);
nand U10149 (N_10149,N_9240,N_9614);
nor U10150 (N_10150,N_9795,N_9975);
and U10151 (N_10151,N_9394,N_9968);
or U10152 (N_10152,N_8893,N_9623);
xnor U10153 (N_10153,N_8216,N_9256);
xnor U10154 (N_10154,N_8367,N_8730);
nand U10155 (N_10155,N_9191,N_9171);
nand U10156 (N_10156,N_9069,N_9727);
nor U10157 (N_10157,N_8490,N_9260);
and U10158 (N_10158,N_8892,N_8944);
xor U10159 (N_10159,N_9520,N_8561);
or U10160 (N_10160,N_9588,N_9246);
xor U10161 (N_10161,N_8241,N_8063);
nor U10162 (N_10162,N_8773,N_8569);
and U10163 (N_10163,N_8281,N_8853);
and U10164 (N_10164,N_8310,N_9041);
nor U10165 (N_10165,N_8756,N_8623);
nor U10166 (N_10166,N_8132,N_9184);
nor U10167 (N_10167,N_9880,N_9622);
xnor U10168 (N_10168,N_8148,N_8010);
and U10169 (N_10169,N_8420,N_8859);
or U10170 (N_10170,N_8609,N_9984);
or U10171 (N_10171,N_9454,N_9135);
xor U10172 (N_10172,N_8628,N_8149);
or U10173 (N_10173,N_9596,N_9393);
or U10174 (N_10174,N_9922,N_9749);
or U10175 (N_10175,N_8074,N_9997);
xor U10176 (N_10176,N_9585,N_8360);
xnor U10177 (N_10177,N_9662,N_9833);
and U10178 (N_10178,N_9540,N_8805);
nor U10179 (N_10179,N_8268,N_9557);
or U10180 (N_10180,N_9923,N_8309);
or U10181 (N_10181,N_8599,N_8152);
or U10182 (N_10182,N_9897,N_9921);
xor U10183 (N_10183,N_9983,N_8435);
xor U10184 (N_10184,N_8078,N_9523);
or U10185 (N_10185,N_8418,N_9371);
nand U10186 (N_10186,N_8546,N_9964);
nand U10187 (N_10187,N_9574,N_9952);
or U10188 (N_10188,N_8942,N_9827);
or U10189 (N_10189,N_9591,N_8199);
nor U10190 (N_10190,N_8218,N_9498);
and U10191 (N_10191,N_8994,N_8740);
nand U10192 (N_10192,N_8266,N_8180);
xnor U10193 (N_10193,N_9573,N_8969);
or U10194 (N_10194,N_9989,N_8729);
nor U10195 (N_10195,N_9408,N_8621);
xor U10196 (N_10196,N_8213,N_9914);
or U10197 (N_10197,N_9365,N_8520);
nand U10198 (N_10198,N_8920,N_9842);
xor U10199 (N_10199,N_8778,N_9994);
nor U10200 (N_10200,N_9209,N_9286);
nor U10201 (N_10201,N_8753,N_9175);
or U10202 (N_10202,N_8763,N_9693);
xnor U10203 (N_10203,N_9652,N_8313);
nor U10204 (N_10204,N_9203,N_8258);
and U10205 (N_10205,N_8471,N_9849);
nand U10206 (N_10206,N_8547,N_8723);
or U10207 (N_10207,N_9549,N_8984);
nand U10208 (N_10208,N_8586,N_9562);
xor U10209 (N_10209,N_9973,N_9789);
or U10210 (N_10210,N_8774,N_9846);
or U10211 (N_10211,N_9860,N_9156);
xnor U10212 (N_10212,N_8899,N_9510);
nand U10213 (N_10213,N_8605,N_8990);
xor U10214 (N_10214,N_8741,N_9712);
xnor U10215 (N_10215,N_8895,N_9986);
nand U10216 (N_10216,N_8680,N_8885);
and U10217 (N_10217,N_8886,N_9732);
nor U10218 (N_10218,N_8254,N_9262);
nor U10219 (N_10219,N_9653,N_9811);
nor U10220 (N_10220,N_9206,N_9045);
nor U10221 (N_10221,N_9785,N_9636);
nor U10222 (N_10222,N_9091,N_8632);
and U10223 (N_10223,N_9147,N_9008);
xor U10224 (N_10224,N_9402,N_8193);
xor U10225 (N_10225,N_9101,N_9741);
nand U10226 (N_10226,N_8432,N_9642);
nor U10227 (N_10227,N_9339,N_8952);
xnor U10228 (N_10228,N_9895,N_8906);
nand U10229 (N_10229,N_9395,N_8348);
xnor U10230 (N_10230,N_8707,N_8878);
nand U10231 (N_10231,N_8476,N_9305);
xnor U10232 (N_10232,N_9659,N_8319);
nand U10233 (N_10233,N_9804,N_9981);
and U10234 (N_10234,N_8288,N_9704);
and U10235 (N_10235,N_9691,N_8228);
xnor U10236 (N_10236,N_9656,N_9312);
or U10237 (N_10237,N_8681,N_9536);
xor U10238 (N_10238,N_9764,N_8423);
nand U10239 (N_10239,N_9447,N_9900);
and U10240 (N_10240,N_9748,N_8615);
and U10241 (N_10241,N_8226,N_8748);
or U10242 (N_10242,N_9991,N_8679);
nand U10243 (N_10243,N_9233,N_8927);
nor U10244 (N_10244,N_9319,N_8168);
or U10245 (N_10245,N_9114,N_8368);
or U10246 (N_10246,N_8792,N_8330);
or U10247 (N_10247,N_8109,N_9068);
and U10248 (N_10248,N_9176,N_9719);
nor U10249 (N_10249,N_8921,N_9134);
or U10250 (N_10250,N_9330,N_9913);
or U10251 (N_10251,N_8003,N_9700);
and U10252 (N_10252,N_8928,N_9231);
nor U10253 (N_10253,N_8441,N_9488);
nor U10254 (N_10254,N_8447,N_9449);
nand U10255 (N_10255,N_9370,N_8438);
nor U10256 (N_10256,N_8236,N_8614);
nand U10257 (N_10257,N_9597,N_9126);
nor U10258 (N_10258,N_8932,N_9361);
xor U10259 (N_10259,N_8428,N_9506);
xnor U10260 (N_10260,N_8867,N_9854);
xor U10261 (N_10261,N_9125,N_9465);
nand U10262 (N_10262,N_9826,N_8950);
and U10263 (N_10263,N_8134,N_8011);
nand U10264 (N_10264,N_9197,N_9898);
and U10265 (N_10265,N_8900,N_8579);
nand U10266 (N_10266,N_8694,N_8221);
xor U10267 (N_10267,N_8117,N_9743);
or U10268 (N_10268,N_9452,N_9582);
xnor U10269 (N_10269,N_9426,N_8301);
nor U10270 (N_10270,N_9415,N_8072);
nand U10271 (N_10271,N_8025,N_9479);
or U10272 (N_10272,N_9077,N_9288);
xor U10273 (N_10273,N_9169,N_8954);
or U10274 (N_10274,N_9621,N_8769);
xor U10275 (N_10275,N_9407,N_9220);
xor U10276 (N_10276,N_9302,N_8559);
nand U10277 (N_10277,N_9896,N_9237);
or U10278 (N_10278,N_9949,N_8646);
nor U10279 (N_10279,N_8818,N_9837);
xnor U10280 (N_10280,N_9079,N_8719);
nor U10281 (N_10281,N_9025,N_8888);
nand U10282 (N_10282,N_9461,N_8165);
xnor U10283 (N_10283,N_8883,N_9368);
or U10284 (N_10284,N_9208,N_8169);
nor U10285 (N_10285,N_8206,N_9144);
and U10286 (N_10286,N_8991,N_8720);
nand U10287 (N_10287,N_9482,N_9410);
nand U10288 (N_10288,N_8512,N_8459);
nand U10289 (N_10289,N_9754,N_9266);
nand U10290 (N_10290,N_9531,N_9547);
nor U10291 (N_10291,N_8040,N_9782);
and U10292 (N_10292,N_8069,N_9601);
nand U10293 (N_10293,N_9518,N_9990);
xnor U10294 (N_10294,N_8483,N_8936);
nand U10295 (N_10295,N_9058,N_9172);
nor U10296 (N_10296,N_9513,N_8825);
nand U10297 (N_10297,N_8722,N_9268);
and U10298 (N_10298,N_9589,N_9877);
nor U10299 (N_10299,N_8377,N_8251);
xnor U10300 (N_10300,N_9665,N_8676);
or U10301 (N_10301,N_8107,N_9309);
or U10302 (N_10302,N_9735,N_9823);
xnor U10303 (N_10303,N_9326,N_8250);
nand U10304 (N_10304,N_8957,N_9985);
nand U10305 (N_10305,N_9159,N_8166);
or U10306 (N_10306,N_8924,N_8653);
nor U10307 (N_10307,N_8287,N_8775);
and U10308 (N_10308,N_9522,N_8033);
or U10309 (N_10309,N_8998,N_8222);
nor U10310 (N_10310,N_9720,N_8638);
nor U10311 (N_10311,N_9188,N_9281);
xnor U10312 (N_10312,N_8493,N_8913);
and U10313 (N_10313,N_8261,N_9494);
nand U10314 (N_10314,N_9917,N_9651);
xor U10315 (N_10315,N_9640,N_8242);
or U10316 (N_10316,N_8745,N_8126);
and U10317 (N_10317,N_8849,N_8835);
and U10318 (N_10318,N_8501,N_9910);
nand U10319 (N_10319,N_9687,N_9251);
and U10320 (N_10320,N_9294,N_8550);
nor U10321 (N_10321,N_8404,N_8427);
or U10322 (N_10322,N_9362,N_8750);
or U10323 (N_10323,N_9927,N_9944);
and U10324 (N_10324,N_9831,N_8253);
nor U10325 (N_10325,N_9834,N_9766);
or U10326 (N_10326,N_9800,N_9218);
xor U10327 (N_10327,N_9103,N_8873);
or U10328 (N_10328,N_8336,N_8077);
nor U10329 (N_10329,N_9358,N_9658);
or U10330 (N_10330,N_9342,N_9946);
xnor U10331 (N_10331,N_8186,N_9020);
and U10332 (N_10332,N_9304,N_9808);
nand U10333 (N_10333,N_9087,N_9389);
or U10334 (N_10334,N_8176,N_8038);
and U10335 (N_10335,N_9333,N_9866);
nor U10336 (N_10336,N_9291,N_8912);
nor U10337 (N_10337,N_9066,N_9604);
xor U10338 (N_10338,N_9618,N_8678);
and U10339 (N_10339,N_9059,N_9760);
or U10340 (N_10340,N_8409,N_8470);
nor U10341 (N_10341,N_8082,N_9857);
xnor U10342 (N_10342,N_9812,N_8070);
nor U10343 (N_10343,N_8517,N_9626);
and U10344 (N_10344,N_9503,N_8683);
or U10345 (N_10345,N_9062,N_8831);
or U10346 (N_10346,N_9242,N_9243);
and U10347 (N_10347,N_8863,N_8858);
nor U10348 (N_10348,N_8552,N_8124);
nand U10349 (N_10349,N_8384,N_8154);
and U10350 (N_10350,N_9674,N_9616);
nor U10351 (N_10351,N_9148,N_9469);
nor U10352 (N_10352,N_9779,N_9639);
or U10353 (N_10353,N_8272,N_8815);
nand U10354 (N_10354,N_9061,N_9725);
or U10355 (N_10355,N_9024,N_8393);
or U10356 (N_10356,N_8979,N_8127);
nor U10357 (N_10357,N_8273,N_9097);
and U10358 (N_10358,N_9385,N_9236);
xnor U10359 (N_10359,N_8840,N_8446);
nand U10360 (N_10360,N_8601,N_9718);
and U10361 (N_10361,N_9637,N_9963);
nand U10362 (N_10362,N_9773,N_9609);
or U10363 (N_10363,N_8095,N_8506);
xor U10364 (N_10364,N_8511,N_8482);
xnor U10365 (N_10365,N_9049,N_8100);
or U10366 (N_10366,N_8200,N_9780);
nor U10367 (N_10367,N_9383,N_9355);
or U10368 (N_10368,N_8051,N_8663);
nor U10369 (N_10369,N_9306,N_8852);
xor U10370 (N_10370,N_8061,N_9092);
and U10371 (N_10371,N_9108,N_8545);
and U10372 (N_10372,N_8966,N_9851);
xor U10373 (N_10373,N_8949,N_8037);
nand U10374 (N_10374,N_8211,N_9162);
nand U10375 (N_10375,N_9939,N_8691);
or U10376 (N_10376,N_9878,N_9027);
or U10377 (N_10377,N_9825,N_9701);
or U10378 (N_10378,N_8353,N_9010);
nor U10379 (N_10379,N_8039,N_8198);
nand U10380 (N_10380,N_9275,N_9822);
and U10381 (N_10381,N_8647,N_9364);
nor U10382 (N_10382,N_8262,N_8788);
nand U10383 (N_10383,N_9163,N_9759);
or U10384 (N_10384,N_9527,N_9594);
xnor U10385 (N_10385,N_9711,N_9724);
nand U10386 (N_10386,N_8312,N_8846);
nor U10387 (N_10387,N_9230,N_8233);
or U10388 (N_10388,N_9182,N_9797);
xor U10389 (N_10389,N_9228,N_9861);
nor U10390 (N_10390,N_9222,N_9412);
nor U10391 (N_10391,N_9253,N_9438);
or U10392 (N_10392,N_9507,N_9645);
nor U10393 (N_10393,N_8981,N_8284);
nand U10394 (N_10394,N_9466,N_8819);
or U10395 (N_10395,N_9196,N_8717);
and U10396 (N_10396,N_8797,N_9867);
nand U10397 (N_10397,N_9793,N_9315);
nor U10398 (N_10398,N_9958,N_9595);
nor U10399 (N_10399,N_8065,N_8390);
or U10400 (N_10400,N_8843,N_8789);
or U10401 (N_10401,N_9539,N_8125);
and U10402 (N_10402,N_8861,N_9888);
and U10403 (N_10403,N_8275,N_9471);
xor U10404 (N_10404,N_8060,N_9028);
nor U10405 (N_10405,N_9078,N_9777);
nor U10406 (N_10406,N_9475,N_8724);
xor U10407 (N_10407,N_9853,N_9668);
and U10408 (N_10408,N_8079,N_9519);
and U10409 (N_10409,N_8766,N_9696);
or U10410 (N_10410,N_8531,N_8386);
xnor U10411 (N_10411,N_9967,N_8032);
nor U10412 (N_10412,N_8970,N_8297);
nor U10413 (N_10413,N_8018,N_8824);
nand U10414 (N_10414,N_8129,N_8449);
nor U10415 (N_10415,N_9043,N_8135);
xor U10416 (N_10416,N_8744,N_8291);
nor U10417 (N_10417,N_8862,N_8772);
or U10418 (N_10418,N_9219,N_8433);
and U10419 (N_10419,N_9474,N_8869);
and U10420 (N_10420,N_8150,N_8106);
xnor U10421 (N_10421,N_9509,N_9706);
nor U10422 (N_10422,N_8532,N_9457);
nor U10423 (N_10423,N_9252,N_8478);
or U10424 (N_10424,N_8333,N_8279);
nand U10425 (N_10425,N_9232,N_9063);
or U10426 (N_10426,N_8160,N_8387);
or U10427 (N_10427,N_9102,N_8845);
nor U10428 (N_10428,N_9090,N_8400);
or U10429 (N_10429,N_9015,N_8341);
or U10430 (N_10430,N_8606,N_8854);
nor U10431 (N_10431,N_8487,N_8305);
or U10432 (N_10432,N_8706,N_8009);
or U10433 (N_10433,N_8838,N_8791);
nand U10434 (N_10434,N_9464,N_8240);
or U10435 (N_10435,N_8881,N_8345);
or U10436 (N_10436,N_8537,N_9396);
and U10437 (N_10437,N_9755,N_9140);
xor U10438 (N_10438,N_8484,N_8158);
xor U10439 (N_10439,N_8091,N_9698);
nand U10440 (N_10440,N_8128,N_8110);
nand U10441 (N_10441,N_9037,N_8365);
and U10442 (N_10442,N_9337,N_8334);
nand U10443 (N_10443,N_9158,N_9023);
nor U10444 (N_10444,N_9685,N_9320);
or U10445 (N_10445,N_8047,N_9292);
and U10446 (N_10446,N_9569,N_8464);
or U10447 (N_10447,N_9467,N_9476);
xor U10448 (N_10448,N_8445,N_8195);
nor U10449 (N_10449,N_9139,N_9406);
or U10450 (N_10450,N_9229,N_9611);
or U10451 (N_10451,N_9705,N_9542);
nand U10452 (N_10452,N_9258,N_8839);
nand U10453 (N_10453,N_8255,N_9118);
and U10454 (N_10454,N_9391,N_8903);
and U10455 (N_10455,N_8392,N_9413);
nor U10456 (N_10456,N_8327,N_9109);
and U10457 (N_10457,N_9872,N_8587);
nand U10458 (N_10458,N_9500,N_9568);
and U10459 (N_10459,N_8298,N_9455);
nand U10460 (N_10460,N_8702,N_8640);
nor U10461 (N_10461,N_9132,N_9708);
nor U10462 (N_10462,N_9677,N_8737);
or U10463 (N_10463,N_8933,N_8739);
nand U10464 (N_10464,N_8380,N_8735);
nand U10465 (N_10465,N_9809,N_8097);
or U10466 (N_10466,N_9663,N_8349);
and U10467 (N_10467,N_9739,N_9316);
nor U10468 (N_10468,N_9073,N_9189);
nand U10469 (N_10469,N_8227,N_9274);
and U10470 (N_10470,N_9349,N_8383);
and U10471 (N_10471,N_9094,N_9458);
nor U10472 (N_10472,N_9598,N_9600);
nand U10473 (N_10473,N_9380,N_8762);
and U10474 (N_10474,N_9048,N_8477);
and U10475 (N_10475,N_9492,N_9057);
xnor U10476 (N_10476,N_8024,N_8658);
nor U10477 (N_10477,N_9884,N_8265);
xor U10478 (N_10478,N_8664,N_8049);
and U10479 (N_10479,N_9496,N_9443);
or U10480 (N_10480,N_8879,N_9104);
nand U10481 (N_10481,N_9729,N_8172);
and U10482 (N_10482,N_8381,N_9734);
xnor U10483 (N_10483,N_9409,N_9002);
xor U10484 (N_10484,N_9318,N_9129);
or U10485 (N_10485,N_9980,N_8161);
nor U10486 (N_10486,N_9357,N_8584);
and U10487 (N_10487,N_9756,N_9679);
nor U10488 (N_10488,N_9047,N_9630);
xor U10489 (N_10489,N_9238,N_9669);
and U10490 (N_10490,N_9678,N_9065);
nand U10491 (N_10491,N_9633,N_8050);
or U10492 (N_10492,N_8689,N_9277);
nor U10493 (N_10493,N_9012,N_9681);
and U10494 (N_10494,N_8013,N_8764);
and U10495 (N_10495,N_9116,N_8224);
xnor U10496 (N_10496,N_9961,N_8046);
nand U10497 (N_10497,N_9040,N_9417);
nor U10498 (N_10498,N_9881,N_8940);
nand U10499 (N_10499,N_9830,N_9810);
nand U10500 (N_10500,N_8572,N_8463);
xor U10501 (N_10501,N_9572,N_8865);
xor U10502 (N_10502,N_9201,N_8439);
nor U10503 (N_10503,N_8637,N_8622);
xnor U10504 (N_10504,N_8860,N_9372);
or U10505 (N_10505,N_9310,N_8486);
or U10506 (N_10506,N_9613,N_8133);
xor U10507 (N_10507,N_9022,N_8422);
and U10508 (N_10508,N_9517,N_9907);
nand U10509 (N_10509,N_8461,N_9781);
xnor U10510 (N_10510,N_8257,N_8048);
or U10511 (N_10511,N_9150,N_8649);
xnor U10512 (N_10512,N_9348,N_8067);
nand U10513 (N_10513,N_8332,N_9581);
nor U10514 (N_10514,N_9882,N_8682);
xnor U10515 (N_10515,N_9794,N_8474);
xor U10516 (N_10516,N_8751,N_9841);
nand U10517 (N_10517,N_9966,N_8017);
or U10518 (N_10518,N_8488,N_8121);
or U10519 (N_10519,N_9280,N_8571);
nor U10520 (N_10520,N_9343,N_9200);
or U10521 (N_10521,N_8686,N_8796);
or U10522 (N_10522,N_8182,N_9578);
xor U10523 (N_10523,N_8114,N_8657);
nor U10524 (N_10524,N_8684,N_8356);
and U10525 (N_10525,N_8610,N_8556);
xor U10526 (N_10526,N_9190,N_9398);
xor U10527 (N_10527,N_8746,N_9437);
nand U10528 (N_10528,N_9786,N_8736);
nor U10529 (N_10529,N_8053,N_9521);
nand U10530 (N_10530,N_8713,N_9925);
and U10531 (N_10531,N_9883,N_8996);
and U10532 (N_10532,N_9634,N_8054);
xor U10533 (N_10533,N_8972,N_9332);
or U10534 (N_10534,N_8088,N_8480);
nand U10535 (N_10535,N_8620,N_9533);
and U10536 (N_10536,N_9211,N_9088);
nor U10537 (N_10537,N_9254,N_8542);
and U10538 (N_10538,N_9676,N_8716);
nand U10539 (N_10539,N_8143,N_9912);
nor U10540 (N_10540,N_8355,N_9978);
xor U10541 (N_10541,N_8391,N_8931);
and U10542 (N_10542,N_8787,N_9550);
nand U10543 (N_10543,N_8594,N_8558);
xor U10544 (N_10544,N_9702,N_9970);
xor U10545 (N_10545,N_9607,N_8577);
nor U10546 (N_10546,N_8910,N_9715);
and U10547 (N_10547,N_8758,N_9767);
or U10548 (N_10548,N_8217,N_8001);
nand U10549 (N_10549,N_8670,N_8157);
nand U10550 (N_10550,N_8238,N_8270);
or U10551 (N_10551,N_9039,N_8209);
nand U10552 (N_10552,N_8144,N_8907);
or U10553 (N_10553,N_8084,N_9778);
nand U10554 (N_10554,N_9599,N_8688);
nand U10555 (N_10555,N_9083,N_8530);
or U10556 (N_10556,N_8855,N_8243);
xnor U10557 (N_10557,N_8183,N_9481);
nand U10558 (N_10558,N_9792,N_8174);
and U10559 (N_10559,N_9334,N_9462);
or U10560 (N_10560,N_8378,N_9971);
or U10561 (N_10561,N_8710,N_8514);
or U10562 (N_10562,N_8889,N_8986);
xnor U10563 (N_10563,N_8832,N_9806);
xor U10564 (N_10564,N_8727,N_8504);
nor U10565 (N_10565,N_8645,N_8045);
xnor U10566 (N_10566,N_9893,N_8977);
and U10567 (N_10567,N_8237,N_9502);
or U10568 (N_10568,N_8935,N_9654);
nand U10569 (N_10569,N_8466,N_8318);
and U10570 (N_10570,N_8634,N_9493);
nand U10571 (N_10571,N_9661,N_8473);
and U10572 (N_10572,N_9053,N_8321);
nand U10573 (N_10573,N_9216,N_8904);
and U10574 (N_10574,N_9683,N_8953);
or U10575 (N_10575,N_8800,N_8549);
or U10576 (N_10576,N_8793,N_8598);
or U10577 (N_10577,N_9113,N_8538);
or U10578 (N_10578,N_9784,N_8747);
or U10579 (N_10579,N_9567,N_8246);
nor U10580 (N_10580,N_9388,N_9340);
xnor U10581 (N_10581,N_9345,N_8968);
nand U10582 (N_10582,N_9421,N_8073);
or U10583 (N_10583,N_9730,N_8163);
xnor U10584 (N_10584,N_9198,N_8372);
nor U10585 (N_10585,N_9605,N_9081);
nand U10586 (N_10586,N_9516,N_8416);
nor U10587 (N_10587,N_9864,N_8167);
and U10588 (N_10588,N_8857,N_9419);
nor U10589 (N_10589,N_9095,N_8347);
or U10590 (N_10590,N_9951,N_8343);
and U10591 (N_10591,N_8749,N_8946);
xnor U10592 (N_10592,N_8847,N_8590);
nor U10593 (N_10593,N_9311,N_8499);
xnor U10594 (N_10594,N_8239,N_9560);
xor U10595 (N_10595,N_9244,N_9817);
and U10596 (N_10596,N_9788,N_8662);
nor U10597 (N_10597,N_9328,N_8105);
or U10598 (N_10598,N_9214,N_9671);
or U10599 (N_10599,N_8930,N_8782);
nand U10600 (N_10600,N_8592,N_8993);
or U10601 (N_10601,N_9042,N_9489);
and U10602 (N_10602,N_8444,N_8525);
and U10603 (N_10603,N_9843,N_9992);
xor U10604 (N_10604,N_8448,N_8364);
nand U10605 (N_10605,N_8363,N_9995);
and U10606 (N_10606,N_9941,N_9682);
xnor U10607 (N_10607,N_8118,N_9241);
and U10608 (N_10608,N_9559,N_8043);
and U10609 (N_10609,N_9617,N_9945);
or U10610 (N_10610,N_8714,N_8102);
nor U10611 (N_10611,N_9263,N_8326);
xor U10612 (N_10612,N_8138,N_8808);
nand U10613 (N_10613,N_9463,N_9606);
xnor U10614 (N_10614,N_9017,N_9565);
and U10615 (N_10615,N_8876,N_8087);
xnor U10616 (N_10616,N_8866,N_9526);
xor U10617 (N_10617,N_9005,N_8890);
nand U10618 (N_10618,N_9680,N_8113);
xor U10619 (N_10619,N_8290,N_8755);
and U10620 (N_10620,N_9295,N_8395);
xor U10621 (N_10621,N_8500,N_8902);
or U10622 (N_10622,N_8495,N_9996);
or U10623 (N_10623,N_9894,N_8884);
xor U10624 (N_10624,N_9450,N_9235);
nand U10625 (N_10625,N_9929,N_9845);
xnor U10626 (N_10626,N_8185,N_8794);
xnor U10627 (N_10627,N_8171,N_9379);
and U10628 (N_10628,N_8656,N_9556);
and U10629 (N_10629,N_9545,N_8562);
and U10630 (N_10630,N_9858,N_8677);
xor U10631 (N_10631,N_8528,N_9133);
or U10632 (N_10632,N_8909,N_9227);
xnor U10633 (N_10633,N_8589,N_9202);
and U10634 (N_10634,N_8812,N_8964);
nor U10635 (N_10635,N_8452,N_9298);
nor U10636 (N_10636,N_9325,N_9137);
nor U10637 (N_10637,N_9282,N_8503);
nor U10638 (N_10638,N_8491,N_9602);
xor U10639 (N_10639,N_8140,N_8489);
xnor U10640 (N_10640,N_9733,N_9688);
xnor U10641 (N_10641,N_9082,N_8976);
and U10642 (N_10642,N_8437,N_9631);
nor U10643 (N_10643,N_8864,N_9505);
nand U10644 (N_10644,N_8798,N_9399);
xor U10645 (N_10645,N_9164,N_8985);
nand U10646 (N_10646,N_9276,N_9717);
nand U10647 (N_10647,N_9428,N_8293);
or U10648 (N_10648,N_9004,N_9501);
and U10649 (N_10649,N_9477,N_9369);
nor U10650 (N_10650,N_9360,N_8156);
or U10651 (N_10651,N_8076,N_8536);
nor U10652 (N_10652,N_8752,N_8164);
nand U10653 (N_10653,N_8743,N_9111);
and U10654 (N_10654,N_8693,N_9728);
xor U10655 (N_10655,N_8799,N_9035);
or U10656 (N_10656,N_9351,N_9018);
nor U10657 (N_10657,N_8306,N_9977);
or U10658 (N_10658,N_8362,N_8151);
nor U10659 (N_10659,N_8557,N_8709);
and U10660 (N_10660,N_9403,N_8983);
nand U10661 (N_10661,N_8120,N_8553);
nor U10662 (N_10662,N_9903,N_8229);
nor U10663 (N_10663,N_8264,N_8468);
or U10664 (N_10664,N_9580,N_8099);
nand U10665 (N_10665,N_8434,N_9938);
or U10666 (N_10666,N_9003,N_9405);
nand U10667 (N_10667,N_8551,N_8696);
and U10668 (N_10668,N_9829,N_8816);
or U10669 (N_10669,N_9381,N_9287);
nand U10670 (N_10670,N_8352,N_9962);
or U10671 (N_10671,N_8534,N_8335);
and U10672 (N_10672,N_9323,N_8141);
and U10673 (N_10673,N_9433,N_8828);
nand U10674 (N_10674,N_9544,N_9213);
or U10675 (N_10675,N_9972,N_9532);
or U10676 (N_10676,N_9152,N_9064);
nand U10677 (N_10677,N_9038,N_9001);
nand U10678 (N_10678,N_8650,N_9145);
nand U10679 (N_10679,N_8225,N_9442);
nor U10680 (N_10680,N_8937,N_8325);
and U10681 (N_10681,N_8916,N_8810);
and U10682 (N_10682,N_8627,N_8573);
nor U10683 (N_10683,N_8971,N_8639);
nand U10684 (N_10684,N_9801,N_8591);
xnor U10685 (N_10685,N_8396,N_8667);
or U10686 (N_10686,N_9690,N_9593);
xnor U10687 (N_10687,N_9106,N_8999);
nand U10688 (N_10688,N_8660,N_8784);
or U10689 (N_10689,N_9257,N_9534);
or U10690 (N_10690,N_8654,N_8028);
nor U10691 (N_10691,N_9416,N_9625);
xnor U10692 (N_10692,N_8092,N_9338);
and U10693 (N_10693,N_9508,N_9862);
or U10694 (N_10694,N_9697,N_9512);
xor U10695 (N_10695,N_9470,N_8978);
nand U10696 (N_10696,N_8820,N_8159);
nor U10697 (N_10697,N_9424,N_9649);
or U10698 (N_10698,N_8021,N_8245);
and U10699 (N_10699,N_8701,N_8475);
nand U10700 (N_10700,N_8376,N_8732);
xor U10701 (N_10701,N_8527,N_8624);
xnor U10702 (N_10702,N_9752,N_8703);
and U10703 (N_10703,N_8479,N_8626);
xor U10704 (N_10704,N_8666,N_8337);
nand U10705 (N_10705,N_9935,N_8555);
nand U10706 (N_10706,N_8570,N_8611);
nor U10707 (N_10707,N_9740,N_9173);
nor U10708 (N_10708,N_8296,N_8131);
and U10709 (N_10709,N_9906,N_8181);
or U10710 (N_10710,N_8019,N_8397);
nand U10711 (N_10711,N_9524,N_8286);
nor U10712 (N_10712,N_9954,N_8096);
nand U10713 (N_10713,N_8071,N_9161);
nor U10714 (N_10714,N_9248,N_9293);
nand U10715 (N_10715,N_9123,N_9852);
nand U10716 (N_10716,N_9644,N_9264);
nand U10717 (N_10717,N_9444,N_8770);
nor U10718 (N_10718,N_9956,N_9120);
and U10719 (N_10719,N_8062,N_8139);
nand U10720 (N_10720,N_8472,N_9225);
xnor U10721 (N_10721,N_9863,N_9269);
nand U10722 (N_10722,N_9267,N_8207);
and U10723 (N_10723,N_8192,N_9632);
nand U10724 (N_10724,N_9181,N_8673);
xnor U10725 (N_10725,N_9011,N_8000);
or U10726 (N_10726,N_9643,N_8802);
and U10727 (N_10727,N_9635,N_9689);
and U10728 (N_10728,N_8108,N_8672);
and U10729 (N_10729,N_8302,N_9105);
and U10730 (N_10730,N_9199,N_8765);
nor U10731 (N_10731,N_9112,N_9110);
or U10732 (N_10732,N_9473,N_8103);
nand U10733 (N_10733,N_9548,N_8036);
nand U10734 (N_10734,N_8259,N_9753);
xnor U10735 (N_10735,N_8581,N_9721);
nand U10736 (N_10736,N_8625,N_8992);
or U10737 (N_10737,N_9955,N_8248);
nand U10738 (N_10738,N_8543,N_8956);
and U10739 (N_10739,N_9430,N_9590);
nand U10740 (N_10740,N_8059,N_9046);
or U10741 (N_10741,N_9096,N_8136);
nor U10742 (N_10742,N_9030,N_9871);
and U10743 (N_10743,N_8661,N_9076);
xnor U10744 (N_10744,N_8602,N_9709);
nand U10745 (N_10745,N_8311,N_8469);
or U10746 (N_10746,N_8086,N_9920);
or U10747 (N_10747,N_9307,N_9168);
and U10748 (N_10748,N_8768,N_9460);
nor U10749 (N_10749,N_8314,N_8526);
or U10750 (N_10750,N_9746,N_8055);
nor U10751 (N_10751,N_9271,N_9308);
and U10752 (N_10752,N_8369,N_8005);
nor U10753 (N_10753,N_9790,N_9703);
nor U10754 (N_10754,N_9564,N_8307);
and U10755 (N_10755,N_9816,N_9765);
nor U10756 (N_10756,N_9832,N_9247);
nand U10757 (N_10757,N_9353,N_8274);
and U10758 (N_10758,N_9180,N_9170);
nor U10759 (N_10759,N_8256,N_9818);
and U10760 (N_10760,N_9194,N_9344);
nand U10761 (N_10761,N_8212,N_8083);
or U10762 (N_10762,N_9546,N_9592);
or U10763 (N_10763,N_9612,N_8837);
nand U10764 (N_10764,N_9089,N_9993);
or U10765 (N_10765,N_8415,N_8851);
and U10766 (N_10766,N_9619,N_9255);
or U10767 (N_10767,N_9487,N_9874);
and U10768 (N_10768,N_9136,N_9552);
or U10769 (N_10769,N_8651,N_8016);
nand U10770 (N_10770,N_8202,N_9555);
and U10771 (N_10771,N_8089,N_8522);
or U10772 (N_10772,N_9757,N_9331);
xnor U10773 (N_10773,N_8567,N_8533);
xnor U10774 (N_10774,N_9033,N_9783);
or U10775 (N_10775,N_8733,N_9166);
or U10776 (N_10776,N_8607,N_8636);
and U10777 (N_10777,N_8616,N_9891);
xnor U10778 (N_10778,N_9234,N_9179);
nand U10779 (N_10779,N_8201,N_9988);
nor U10780 (N_10780,N_8191,N_9608);
and U10781 (N_10781,N_8809,N_8034);
xor U10782 (N_10782,N_8426,N_8635);
or U10783 (N_10783,N_9451,N_8563);
or U10784 (N_10784,N_8197,N_8580);
nand U10785 (N_10785,N_8315,N_9776);
and U10786 (N_10786,N_8317,N_9432);
xor U10787 (N_10787,N_8269,N_8929);
or U10788 (N_10788,N_8417,N_9026);
nor U10789 (N_10789,N_9902,N_8002);
xnor U10790 (N_10790,N_8006,N_8738);
and U10791 (N_10791,N_9848,N_8340);
xnor U10792 (N_10792,N_8358,N_9960);
or U10793 (N_10793,N_8285,N_9815);
and U10794 (N_10794,N_8316,N_9722);
or U10795 (N_10795,N_8554,N_8382);
and U10796 (N_10796,N_9924,N_9541);
nor U10797 (N_10797,N_9714,N_9434);
nor U10798 (N_10798,N_8699,N_9650);
nor U10799 (N_10799,N_9446,N_9499);
xnor U10800 (N_10800,N_9051,N_8844);
nand U10801 (N_10801,N_8460,N_8524);
and U10802 (N_10802,N_8583,N_9763);
nand U10803 (N_10803,N_8596,N_8734);
and U10804 (N_10804,N_8712,N_8776);
nand U10805 (N_10805,N_9021,N_8917);
and U10806 (N_10806,N_8029,N_9067);
and U10807 (N_10807,N_9142,N_9576);
and U10808 (N_10808,N_8230,N_8568);
nand U10809 (N_10809,N_8220,N_9850);
and U10810 (N_10810,N_8414,N_8655);
or U10811 (N_10811,N_8962,N_9270);
nor U10812 (N_10812,N_8947,N_9791);
nor U10813 (N_10813,N_9072,N_9418);
nor U10814 (N_10814,N_8177,N_9761);
nand U10815 (N_10815,N_9151,N_8030);
nor U10816 (N_10816,N_8419,N_9006);
and U10817 (N_10817,N_9905,N_9217);
nand U10818 (N_10818,N_8104,N_8430);
and U10819 (N_10819,N_9356,N_9215);
xor U10820 (N_10820,N_9375,N_9387);
or U10821 (N_10821,N_8234,N_9187);
xnor U10822 (N_10822,N_8366,N_8848);
nand U10823 (N_10823,N_8575,N_8492);
and U10824 (N_10824,N_9762,N_8401);
or U10825 (N_10825,N_9672,N_8697);
nand U10826 (N_10826,N_8116,N_8505);
and U10827 (N_10827,N_9770,N_9710);
xor U10828 (N_10828,N_8785,N_9259);
nor U10829 (N_10829,N_8922,N_9367);
nor U10830 (N_10830,N_9167,N_9193);
or U10831 (N_10831,N_9530,N_9192);
and U10832 (N_10832,N_8874,N_9969);
nor U10833 (N_10833,N_8374,N_8850);
nor U10834 (N_10834,N_9441,N_8497);
nor U10835 (N_10835,N_9919,N_8905);
nand U10836 (N_10836,N_9566,N_9768);
and U10837 (N_10837,N_9397,N_9221);
nand U10838 (N_10838,N_9070,N_9459);
xor U10839 (N_10839,N_9436,N_8007);
nand U10840 (N_10840,N_8188,N_8987);
or U10841 (N_10841,N_9204,N_8184);
or U10842 (N_10842,N_9561,N_9296);
xnor U10843 (N_10843,N_9805,N_8974);
or U10844 (N_10844,N_9074,N_8617);
xor U10845 (N_10845,N_9322,N_8945);
nand U10846 (N_10846,N_9869,N_8705);
and U10847 (N_10847,N_8252,N_8292);
xnor U10848 (N_10848,N_9453,N_9859);
xnor U10849 (N_10849,N_8518,N_9283);
or U10850 (N_10850,N_9553,N_8539);
nor U10851 (N_10851,N_8692,N_8652);
and U10852 (N_10852,N_8811,N_8481);
nor U10853 (N_10853,N_9400,N_8370);
nand U10854 (N_10854,N_8708,N_9750);
or U10855 (N_10855,N_8379,N_8685);
nand U10856 (N_10856,N_8516,N_8399);
and U10857 (N_10857,N_9084,N_8760);
and U10858 (N_10858,N_9207,N_9909);
or U10859 (N_10859,N_8560,N_9538);
nor U10860 (N_10860,N_9901,N_8208);
and U10861 (N_10861,N_8704,N_9933);
or U10862 (N_10862,N_8263,N_9290);
nand U10863 (N_10863,N_9289,N_9695);
and U10864 (N_10864,N_8644,N_8451);
nand U10865 (N_10865,N_8232,N_9947);
nor U10866 (N_10866,N_8056,N_9390);
and U10867 (N_10867,N_8436,N_8613);
nand U10868 (N_10868,N_9265,N_9435);
xor U10869 (N_10869,N_9327,N_9157);
and U10870 (N_10870,N_9404,N_9667);
and U10871 (N_10871,N_9796,N_9384);
nor U10872 (N_10872,N_9086,N_9363);
xor U10873 (N_10873,N_8203,N_8456);
or U10874 (N_10874,N_8098,N_9448);
or U10875 (N_10875,N_9928,N_9627);
nand U10876 (N_10876,N_9347,N_9838);
or U10877 (N_10877,N_8267,N_9122);
or U10878 (N_10878,N_9950,N_9844);
or U10879 (N_10879,N_9483,N_8519);
and U10880 (N_10880,N_9943,N_9655);
nand U10881 (N_10881,N_9940,N_9916);
and U10882 (N_10882,N_8988,N_9769);
xnor U10883 (N_10883,N_8398,N_8080);
or U10884 (N_10884,N_8674,N_8731);
or U10885 (N_10885,N_9744,N_8147);
xor U10886 (N_10886,N_8955,N_8012);
nand U10887 (N_10887,N_8410,N_9016);
and U10888 (N_10888,N_8669,N_8394);
or U10889 (N_10889,N_8997,N_9128);
xor U10890 (N_10890,N_9080,N_9787);
or U10891 (N_10891,N_9855,N_8926);
nand U10892 (N_10892,N_9143,N_9819);
or U10893 (N_10893,N_8442,N_9579);
or U10894 (N_10894,N_8540,N_9382);
or U10895 (N_10895,N_9932,N_9141);
nand U10896 (N_10896,N_9802,N_9130);
nor U10897 (N_10897,N_9603,N_8856);
xor U10898 (N_10898,N_9628,N_9686);
or U10899 (N_10899,N_9876,N_9186);
xor U10900 (N_10900,N_9336,N_9666);
or U10901 (N_10901,N_9100,N_8721);
xor U10902 (N_10902,N_8948,N_9774);
and U10903 (N_10903,N_9093,N_9054);
nor U10904 (N_10904,N_8989,N_9982);
or U10905 (N_10905,N_8303,N_8403);
nor U10906 (N_10906,N_8938,N_9865);
nor U10907 (N_10907,N_8833,N_8665);
xnor U10908 (N_10908,N_8742,N_9376);
and U10909 (N_10909,N_8214,N_9445);
or U10910 (N_10910,N_9205,N_9911);
xor U10911 (N_10911,N_8918,N_9439);
nand U10912 (N_10912,N_8943,N_8385);
xor U10913 (N_10913,N_9558,N_9707);
xnor U10914 (N_10914,N_9726,N_8814);
nor U10915 (N_10915,N_9324,N_8454);
or U10916 (N_10916,N_8771,N_8529);
nand U10917 (N_10917,N_8995,N_9836);
nor U10918 (N_10918,N_9034,N_8817);
or U10919 (N_10919,N_9584,N_8767);
and U10920 (N_10920,N_9245,N_8440);
nand U10921 (N_10921,N_9886,N_9099);
or U10922 (N_10922,N_9936,N_8725);
nand U10923 (N_10923,N_9918,N_8803);
or U10924 (N_10924,N_8223,N_9468);
xor U10925 (N_10925,N_9249,N_8502);
nor U10926 (N_10926,N_9374,N_9456);
nor U10927 (N_10927,N_9828,N_8958);
nor U10928 (N_10928,N_8882,N_8453);
and U10929 (N_10929,N_8830,N_9490);
nor U10930 (N_10930,N_9373,N_8914);
or U10931 (N_10931,N_9174,N_9297);
xnor U10932 (N_10932,N_9879,N_8090);
and U10933 (N_10933,N_8354,N_8111);
and U10934 (N_10934,N_8026,N_8194);
xor U10935 (N_10935,N_8115,N_8960);
and U10936 (N_10936,N_9261,N_9177);
nor U10937 (N_10937,N_8458,N_8189);
nor U10938 (N_10938,N_9485,N_9736);
xnor U10939 (N_10939,N_8044,N_8521);
and U10940 (N_10940,N_8280,N_9673);
nand U10941 (N_10941,N_8668,N_8004);
nand U10942 (N_10942,N_9146,N_8276);
or U10943 (N_10943,N_8350,N_8967);
and U10944 (N_10944,N_8329,N_9341);
or U10945 (N_10945,N_9009,N_9875);
xor U10946 (N_10946,N_9314,N_9032);
and U10947 (N_10947,N_8951,N_8346);
and U10948 (N_10948,N_8574,N_8294);
nand U10949 (N_10949,N_8619,N_8582);
and U10950 (N_10950,N_8205,N_8961);
nor U10951 (N_10951,N_9354,N_9620);
xnor U10952 (N_10952,N_9758,N_8757);
xor U10953 (N_10953,N_9716,N_9824);
or U10954 (N_10954,N_8031,N_9868);
or U10955 (N_10955,N_9484,N_9183);
or U10956 (N_10956,N_9350,N_8544);
nor U10957 (N_10957,N_8068,N_9359);
nor U10958 (N_10958,N_8576,N_8320);
nand U10959 (N_10959,N_8431,N_9772);
nor U10960 (N_10960,N_8042,N_8807);
or U10961 (N_10961,N_9571,N_9930);
nand U10962 (N_10962,N_8411,N_9931);
nor U10963 (N_10963,N_9624,N_9504);
nand U10964 (N_10964,N_8187,N_9948);
xor U10965 (N_10965,N_8190,N_9870);
or U10966 (N_10966,N_8980,N_8244);
or U10967 (N_10967,N_9014,N_8604);
nand U10968 (N_10968,N_9425,N_8695);
nor U10969 (N_10969,N_9036,N_8375);
nor U10970 (N_10970,N_8925,N_8271);
nand U10971 (N_10971,N_8413,N_9803);
xnor U10972 (N_10972,N_8671,N_8075);
or U10973 (N_10973,N_8612,N_8633);
nor U10974 (N_10974,N_9575,N_8323);
or U10975 (N_10975,N_9160,N_9440);
xnor U10976 (N_10976,N_8112,N_8496);
nand U10977 (N_10977,N_8690,N_9551);
nor U10978 (N_10978,N_8754,N_8728);
and U10979 (N_10979,N_8260,N_8339);
xnor U10980 (N_10980,N_8827,N_8304);
or U10981 (N_10981,N_9899,N_9423);
or U10982 (N_10982,N_9570,N_9497);
nand U10983 (N_10983,N_8786,N_8351);
nand U10984 (N_10984,N_9117,N_9478);
nand U10985 (N_10985,N_8324,N_8142);
nand U10986 (N_10986,N_8508,N_8826);
nor U10987 (N_10987,N_9934,N_9694);
or U10988 (N_10988,N_8777,N_9119);
and U10989 (N_10989,N_9692,N_9525);
or U10990 (N_10990,N_9495,N_9660);
or U10991 (N_10991,N_8629,N_9840);
nor U10992 (N_10992,N_9583,N_8462);
and U10993 (N_10993,N_8965,N_9075);
nor U10994 (N_10994,N_9019,N_9646);
nor U10995 (N_10995,N_8880,N_8509);
nor U10996 (N_10996,N_9491,N_8939);
or U10997 (N_10997,N_9587,N_9127);
nor U10998 (N_10998,N_8179,N_8027);
xor U10999 (N_10999,N_9713,N_9684);
nand U11000 (N_11000,N_8582,N_9406);
xor U11001 (N_11001,N_9163,N_8873);
and U11002 (N_11002,N_8556,N_9188);
nor U11003 (N_11003,N_9583,N_8974);
or U11004 (N_11004,N_9475,N_9113);
or U11005 (N_11005,N_9009,N_9506);
nand U11006 (N_11006,N_8624,N_9998);
nand U11007 (N_11007,N_8161,N_8224);
and U11008 (N_11008,N_8134,N_9745);
or U11009 (N_11009,N_8036,N_9557);
nand U11010 (N_11010,N_8995,N_8314);
xnor U11011 (N_11011,N_8865,N_9645);
and U11012 (N_11012,N_8647,N_9582);
nand U11013 (N_11013,N_9137,N_8502);
xor U11014 (N_11014,N_8204,N_8786);
and U11015 (N_11015,N_9852,N_9482);
or U11016 (N_11016,N_8548,N_9206);
nand U11017 (N_11017,N_8666,N_9772);
nor U11018 (N_11018,N_9145,N_9522);
and U11019 (N_11019,N_9606,N_8300);
xnor U11020 (N_11020,N_9142,N_8914);
or U11021 (N_11021,N_9662,N_9647);
or U11022 (N_11022,N_8551,N_8987);
and U11023 (N_11023,N_9339,N_9250);
xor U11024 (N_11024,N_8913,N_8626);
or U11025 (N_11025,N_8111,N_8397);
nand U11026 (N_11026,N_9094,N_8945);
or U11027 (N_11027,N_9130,N_9823);
nand U11028 (N_11028,N_9572,N_9331);
or U11029 (N_11029,N_8857,N_8518);
nand U11030 (N_11030,N_9111,N_9388);
nor U11031 (N_11031,N_9946,N_9894);
nor U11032 (N_11032,N_8157,N_9377);
and U11033 (N_11033,N_8011,N_9915);
nand U11034 (N_11034,N_9771,N_9990);
and U11035 (N_11035,N_9647,N_9885);
and U11036 (N_11036,N_9469,N_8217);
nand U11037 (N_11037,N_9874,N_9207);
nand U11038 (N_11038,N_9277,N_8431);
xnor U11039 (N_11039,N_9202,N_8705);
and U11040 (N_11040,N_8993,N_8236);
and U11041 (N_11041,N_9120,N_9284);
nor U11042 (N_11042,N_8436,N_8615);
nor U11043 (N_11043,N_9018,N_9283);
nor U11044 (N_11044,N_8330,N_8211);
nor U11045 (N_11045,N_8160,N_8413);
and U11046 (N_11046,N_8249,N_9984);
xor U11047 (N_11047,N_9943,N_9192);
nand U11048 (N_11048,N_8745,N_8823);
or U11049 (N_11049,N_8687,N_8284);
and U11050 (N_11050,N_8590,N_8151);
or U11051 (N_11051,N_8000,N_9813);
nand U11052 (N_11052,N_8238,N_8638);
xor U11053 (N_11053,N_9165,N_9392);
and U11054 (N_11054,N_9423,N_8100);
xor U11055 (N_11055,N_9246,N_9605);
xnor U11056 (N_11056,N_8333,N_9332);
xnor U11057 (N_11057,N_8480,N_8680);
nor U11058 (N_11058,N_9313,N_9988);
xnor U11059 (N_11059,N_9631,N_8197);
nor U11060 (N_11060,N_8558,N_8689);
nor U11061 (N_11061,N_8398,N_8374);
xnor U11062 (N_11062,N_8229,N_8695);
nand U11063 (N_11063,N_8301,N_9634);
xnor U11064 (N_11064,N_9672,N_9245);
nor U11065 (N_11065,N_8175,N_9707);
xnor U11066 (N_11066,N_8518,N_9342);
nand U11067 (N_11067,N_9252,N_9542);
or U11068 (N_11068,N_9072,N_9716);
and U11069 (N_11069,N_8557,N_9646);
nand U11070 (N_11070,N_8629,N_9044);
xnor U11071 (N_11071,N_8184,N_9305);
xor U11072 (N_11072,N_9468,N_9775);
nor U11073 (N_11073,N_9282,N_8444);
or U11074 (N_11074,N_8137,N_8850);
nor U11075 (N_11075,N_9543,N_9791);
xnor U11076 (N_11076,N_9751,N_9138);
nor U11077 (N_11077,N_8884,N_9160);
and U11078 (N_11078,N_8085,N_9274);
and U11079 (N_11079,N_9240,N_9212);
or U11080 (N_11080,N_8839,N_8453);
and U11081 (N_11081,N_8621,N_8831);
xor U11082 (N_11082,N_8613,N_8011);
nor U11083 (N_11083,N_8772,N_9559);
or U11084 (N_11084,N_8936,N_8138);
xor U11085 (N_11085,N_9867,N_8026);
nor U11086 (N_11086,N_9331,N_9442);
or U11087 (N_11087,N_8591,N_9521);
or U11088 (N_11088,N_9403,N_9915);
or U11089 (N_11089,N_9566,N_9834);
or U11090 (N_11090,N_9563,N_9025);
xor U11091 (N_11091,N_8629,N_9378);
nor U11092 (N_11092,N_8645,N_9752);
or U11093 (N_11093,N_9607,N_8951);
nand U11094 (N_11094,N_9033,N_9647);
or U11095 (N_11095,N_8094,N_8195);
nand U11096 (N_11096,N_8998,N_9877);
or U11097 (N_11097,N_8708,N_8302);
and U11098 (N_11098,N_8687,N_8570);
xnor U11099 (N_11099,N_8378,N_9651);
xnor U11100 (N_11100,N_9951,N_8427);
and U11101 (N_11101,N_9827,N_8581);
xnor U11102 (N_11102,N_9491,N_8984);
xnor U11103 (N_11103,N_8346,N_8582);
nand U11104 (N_11104,N_8621,N_9720);
nand U11105 (N_11105,N_8383,N_8756);
and U11106 (N_11106,N_9746,N_9171);
and U11107 (N_11107,N_9707,N_9731);
nor U11108 (N_11108,N_8608,N_8538);
nand U11109 (N_11109,N_9525,N_8309);
nand U11110 (N_11110,N_9877,N_8170);
xnor U11111 (N_11111,N_8460,N_9545);
or U11112 (N_11112,N_8114,N_9211);
xnor U11113 (N_11113,N_8488,N_8924);
and U11114 (N_11114,N_9547,N_8432);
nor U11115 (N_11115,N_8067,N_8239);
xnor U11116 (N_11116,N_8669,N_9051);
xnor U11117 (N_11117,N_9690,N_8184);
xnor U11118 (N_11118,N_9167,N_8059);
nor U11119 (N_11119,N_9137,N_8598);
xor U11120 (N_11120,N_9374,N_9594);
nand U11121 (N_11121,N_8518,N_8580);
nor U11122 (N_11122,N_8404,N_9595);
xnor U11123 (N_11123,N_8246,N_9993);
or U11124 (N_11124,N_8836,N_9221);
or U11125 (N_11125,N_9604,N_9581);
nand U11126 (N_11126,N_8371,N_9963);
and U11127 (N_11127,N_8006,N_8513);
and U11128 (N_11128,N_9589,N_8893);
xnor U11129 (N_11129,N_8956,N_9857);
nand U11130 (N_11130,N_9168,N_8378);
and U11131 (N_11131,N_8823,N_8166);
xor U11132 (N_11132,N_9404,N_9724);
nor U11133 (N_11133,N_8525,N_9299);
nor U11134 (N_11134,N_8527,N_8248);
nand U11135 (N_11135,N_9084,N_8158);
and U11136 (N_11136,N_8161,N_8921);
nor U11137 (N_11137,N_9382,N_8224);
or U11138 (N_11138,N_8346,N_8822);
and U11139 (N_11139,N_8803,N_9226);
or U11140 (N_11140,N_9425,N_9889);
nand U11141 (N_11141,N_9025,N_9307);
xor U11142 (N_11142,N_8431,N_8361);
nand U11143 (N_11143,N_9467,N_9074);
or U11144 (N_11144,N_8500,N_8331);
or U11145 (N_11145,N_8528,N_9842);
or U11146 (N_11146,N_8672,N_8868);
nor U11147 (N_11147,N_8157,N_9606);
or U11148 (N_11148,N_9326,N_9059);
or U11149 (N_11149,N_8094,N_8450);
or U11150 (N_11150,N_8966,N_8724);
nand U11151 (N_11151,N_8296,N_9962);
xor U11152 (N_11152,N_8862,N_9370);
nand U11153 (N_11153,N_9392,N_8295);
and U11154 (N_11154,N_8157,N_8454);
nand U11155 (N_11155,N_9291,N_8244);
xnor U11156 (N_11156,N_9533,N_8839);
nand U11157 (N_11157,N_9856,N_8270);
nor U11158 (N_11158,N_8123,N_9748);
and U11159 (N_11159,N_9596,N_8627);
and U11160 (N_11160,N_9872,N_9997);
nand U11161 (N_11161,N_8924,N_8781);
nand U11162 (N_11162,N_8297,N_8483);
xor U11163 (N_11163,N_9484,N_8541);
or U11164 (N_11164,N_8740,N_8220);
nor U11165 (N_11165,N_9441,N_8914);
or U11166 (N_11166,N_8827,N_8833);
xor U11167 (N_11167,N_8691,N_9963);
nor U11168 (N_11168,N_9782,N_9129);
xnor U11169 (N_11169,N_8833,N_8848);
xor U11170 (N_11170,N_8125,N_9160);
or U11171 (N_11171,N_9576,N_9481);
and U11172 (N_11172,N_8095,N_8903);
nor U11173 (N_11173,N_8265,N_9464);
xnor U11174 (N_11174,N_8764,N_8248);
nor U11175 (N_11175,N_9489,N_9137);
nor U11176 (N_11176,N_9700,N_9375);
nand U11177 (N_11177,N_9125,N_9398);
and U11178 (N_11178,N_8739,N_9895);
or U11179 (N_11179,N_9269,N_9169);
xnor U11180 (N_11180,N_8010,N_9444);
nor U11181 (N_11181,N_9754,N_8439);
nand U11182 (N_11182,N_9592,N_9049);
nand U11183 (N_11183,N_8051,N_9772);
or U11184 (N_11184,N_8146,N_8060);
or U11185 (N_11185,N_8521,N_9833);
and U11186 (N_11186,N_9239,N_9005);
nor U11187 (N_11187,N_8857,N_8414);
or U11188 (N_11188,N_9199,N_9512);
or U11189 (N_11189,N_9182,N_9355);
nor U11190 (N_11190,N_8803,N_9548);
nor U11191 (N_11191,N_9821,N_9547);
or U11192 (N_11192,N_9036,N_8348);
nor U11193 (N_11193,N_8982,N_8267);
and U11194 (N_11194,N_8516,N_8053);
nand U11195 (N_11195,N_8428,N_9514);
xnor U11196 (N_11196,N_9259,N_8775);
or U11197 (N_11197,N_8884,N_9925);
nor U11198 (N_11198,N_8681,N_9377);
or U11199 (N_11199,N_8584,N_8756);
nor U11200 (N_11200,N_9323,N_9105);
nand U11201 (N_11201,N_9963,N_8995);
xor U11202 (N_11202,N_8571,N_8197);
nand U11203 (N_11203,N_8130,N_8645);
or U11204 (N_11204,N_9718,N_8971);
xor U11205 (N_11205,N_9760,N_8117);
nor U11206 (N_11206,N_9932,N_9163);
and U11207 (N_11207,N_8439,N_9499);
nor U11208 (N_11208,N_9093,N_8652);
and U11209 (N_11209,N_8246,N_9540);
nand U11210 (N_11210,N_8978,N_8796);
nor U11211 (N_11211,N_9159,N_8557);
nand U11212 (N_11212,N_9004,N_8394);
and U11213 (N_11213,N_8538,N_8599);
xor U11214 (N_11214,N_8127,N_8038);
xor U11215 (N_11215,N_8774,N_9087);
nor U11216 (N_11216,N_8008,N_9229);
nor U11217 (N_11217,N_9267,N_8273);
nand U11218 (N_11218,N_8163,N_9458);
nand U11219 (N_11219,N_8125,N_9586);
nor U11220 (N_11220,N_8932,N_8070);
or U11221 (N_11221,N_8945,N_9570);
xnor U11222 (N_11222,N_9754,N_8709);
or U11223 (N_11223,N_8969,N_8247);
nor U11224 (N_11224,N_8684,N_9701);
nand U11225 (N_11225,N_9335,N_9547);
nor U11226 (N_11226,N_8659,N_8469);
nor U11227 (N_11227,N_9503,N_8200);
xnor U11228 (N_11228,N_8016,N_8876);
or U11229 (N_11229,N_9141,N_8303);
or U11230 (N_11230,N_8160,N_8257);
nor U11231 (N_11231,N_8262,N_9279);
and U11232 (N_11232,N_8007,N_8018);
nand U11233 (N_11233,N_9885,N_9792);
nand U11234 (N_11234,N_9013,N_9191);
nand U11235 (N_11235,N_8576,N_8255);
or U11236 (N_11236,N_8385,N_9323);
nor U11237 (N_11237,N_8061,N_9874);
nor U11238 (N_11238,N_8630,N_9367);
or U11239 (N_11239,N_8177,N_8573);
and U11240 (N_11240,N_8030,N_8715);
nor U11241 (N_11241,N_9497,N_9476);
nand U11242 (N_11242,N_9538,N_9436);
xnor U11243 (N_11243,N_9419,N_8067);
xor U11244 (N_11244,N_8071,N_9980);
and U11245 (N_11245,N_8615,N_9095);
nand U11246 (N_11246,N_8238,N_9859);
nor U11247 (N_11247,N_9304,N_9946);
nand U11248 (N_11248,N_8296,N_8140);
or U11249 (N_11249,N_9593,N_9441);
or U11250 (N_11250,N_8775,N_8764);
xnor U11251 (N_11251,N_9494,N_8045);
nand U11252 (N_11252,N_8213,N_8234);
nand U11253 (N_11253,N_9250,N_8057);
xor U11254 (N_11254,N_8008,N_8687);
xnor U11255 (N_11255,N_8139,N_9557);
xor U11256 (N_11256,N_8196,N_9545);
and U11257 (N_11257,N_9784,N_9060);
xor U11258 (N_11258,N_9058,N_9136);
or U11259 (N_11259,N_8896,N_8941);
nand U11260 (N_11260,N_9993,N_9701);
nor U11261 (N_11261,N_9889,N_9138);
and U11262 (N_11262,N_9928,N_8787);
or U11263 (N_11263,N_9878,N_8369);
nor U11264 (N_11264,N_8774,N_9923);
and U11265 (N_11265,N_9570,N_9882);
or U11266 (N_11266,N_9917,N_9489);
nor U11267 (N_11267,N_8379,N_9913);
nand U11268 (N_11268,N_8550,N_8302);
and U11269 (N_11269,N_8452,N_8694);
and U11270 (N_11270,N_8045,N_8546);
or U11271 (N_11271,N_8875,N_9878);
or U11272 (N_11272,N_8188,N_9329);
xor U11273 (N_11273,N_9820,N_8613);
xnor U11274 (N_11274,N_9581,N_9071);
or U11275 (N_11275,N_8369,N_8701);
nand U11276 (N_11276,N_8856,N_8634);
xnor U11277 (N_11277,N_9096,N_8458);
and U11278 (N_11278,N_8237,N_9470);
nand U11279 (N_11279,N_9748,N_9726);
nor U11280 (N_11280,N_9074,N_9815);
nor U11281 (N_11281,N_8419,N_8542);
nand U11282 (N_11282,N_9228,N_9783);
xnor U11283 (N_11283,N_8579,N_9185);
nand U11284 (N_11284,N_8299,N_8509);
and U11285 (N_11285,N_9226,N_8269);
nand U11286 (N_11286,N_8975,N_9163);
nand U11287 (N_11287,N_8752,N_8537);
xnor U11288 (N_11288,N_9355,N_9461);
or U11289 (N_11289,N_8348,N_8084);
nand U11290 (N_11290,N_8562,N_8637);
or U11291 (N_11291,N_9728,N_9172);
nor U11292 (N_11292,N_9936,N_8227);
and U11293 (N_11293,N_9140,N_8186);
nand U11294 (N_11294,N_8407,N_8737);
and U11295 (N_11295,N_8985,N_9859);
nor U11296 (N_11296,N_8488,N_9244);
nand U11297 (N_11297,N_8391,N_8643);
nor U11298 (N_11298,N_8594,N_8314);
and U11299 (N_11299,N_8836,N_9700);
and U11300 (N_11300,N_8507,N_9514);
nand U11301 (N_11301,N_9637,N_9714);
nor U11302 (N_11302,N_8237,N_8140);
or U11303 (N_11303,N_8155,N_9151);
nand U11304 (N_11304,N_9807,N_9006);
nand U11305 (N_11305,N_8952,N_8225);
nand U11306 (N_11306,N_9110,N_8932);
or U11307 (N_11307,N_8700,N_8593);
or U11308 (N_11308,N_8098,N_8891);
nor U11309 (N_11309,N_8883,N_8892);
xor U11310 (N_11310,N_9405,N_8304);
or U11311 (N_11311,N_8257,N_9352);
xor U11312 (N_11312,N_8952,N_9302);
and U11313 (N_11313,N_8784,N_9671);
and U11314 (N_11314,N_8455,N_8490);
or U11315 (N_11315,N_8541,N_8194);
or U11316 (N_11316,N_9916,N_9076);
xnor U11317 (N_11317,N_9413,N_8890);
and U11318 (N_11318,N_8650,N_8173);
xnor U11319 (N_11319,N_8720,N_9271);
xor U11320 (N_11320,N_9550,N_9694);
or U11321 (N_11321,N_8013,N_8674);
nand U11322 (N_11322,N_8134,N_9896);
nand U11323 (N_11323,N_9588,N_9946);
xnor U11324 (N_11324,N_9085,N_8999);
nand U11325 (N_11325,N_9452,N_8982);
or U11326 (N_11326,N_8886,N_8608);
nor U11327 (N_11327,N_8861,N_8330);
nor U11328 (N_11328,N_8353,N_8735);
and U11329 (N_11329,N_9711,N_9988);
and U11330 (N_11330,N_8397,N_8503);
or U11331 (N_11331,N_8624,N_9063);
xor U11332 (N_11332,N_9594,N_8654);
and U11333 (N_11333,N_8616,N_8432);
nand U11334 (N_11334,N_9490,N_9356);
or U11335 (N_11335,N_9888,N_8389);
or U11336 (N_11336,N_8695,N_9967);
nor U11337 (N_11337,N_8023,N_8921);
xnor U11338 (N_11338,N_8358,N_8338);
xor U11339 (N_11339,N_8073,N_9089);
or U11340 (N_11340,N_8268,N_9367);
nor U11341 (N_11341,N_8776,N_9748);
nor U11342 (N_11342,N_9120,N_8418);
xnor U11343 (N_11343,N_8527,N_9047);
xnor U11344 (N_11344,N_8113,N_9883);
and U11345 (N_11345,N_8863,N_9850);
nand U11346 (N_11346,N_9610,N_9468);
and U11347 (N_11347,N_9442,N_8943);
or U11348 (N_11348,N_9576,N_8177);
nor U11349 (N_11349,N_9106,N_9149);
nor U11350 (N_11350,N_8007,N_9370);
nand U11351 (N_11351,N_8230,N_8626);
nand U11352 (N_11352,N_9402,N_9630);
and U11353 (N_11353,N_9647,N_8222);
nor U11354 (N_11354,N_8127,N_8873);
or U11355 (N_11355,N_9601,N_9870);
xnor U11356 (N_11356,N_8587,N_9454);
and U11357 (N_11357,N_8455,N_8939);
nor U11358 (N_11358,N_8794,N_9023);
and U11359 (N_11359,N_9638,N_9274);
xor U11360 (N_11360,N_8015,N_9072);
xnor U11361 (N_11361,N_9307,N_8173);
nand U11362 (N_11362,N_8687,N_8992);
nand U11363 (N_11363,N_9274,N_8962);
xnor U11364 (N_11364,N_9104,N_9963);
xor U11365 (N_11365,N_8797,N_8143);
nor U11366 (N_11366,N_8387,N_8984);
nand U11367 (N_11367,N_8404,N_8657);
nor U11368 (N_11368,N_8998,N_9691);
nor U11369 (N_11369,N_9232,N_9739);
or U11370 (N_11370,N_9246,N_8625);
xnor U11371 (N_11371,N_9558,N_9806);
nand U11372 (N_11372,N_9667,N_9746);
and U11373 (N_11373,N_9545,N_9420);
nor U11374 (N_11374,N_8666,N_9116);
and U11375 (N_11375,N_8064,N_8654);
xnor U11376 (N_11376,N_9017,N_8669);
nand U11377 (N_11377,N_9613,N_9068);
xnor U11378 (N_11378,N_9334,N_9268);
xnor U11379 (N_11379,N_9268,N_8456);
nor U11380 (N_11380,N_8892,N_8005);
nor U11381 (N_11381,N_9815,N_8281);
or U11382 (N_11382,N_8325,N_9827);
nor U11383 (N_11383,N_9247,N_8484);
xor U11384 (N_11384,N_9891,N_9794);
nor U11385 (N_11385,N_8242,N_8045);
nand U11386 (N_11386,N_9615,N_8243);
or U11387 (N_11387,N_8157,N_8663);
xnor U11388 (N_11388,N_8164,N_8271);
nand U11389 (N_11389,N_8578,N_9784);
xor U11390 (N_11390,N_9929,N_9365);
xor U11391 (N_11391,N_8934,N_9866);
nand U11392 (N_11392,N_8428,N_8564);
and U11393 (N_11393,N_9313,N_9806);
nand U11394 (N_11394,N_9308,N_9348);
or U11395 (N_11395,N_9280,N_8541);
nand U11396 (N_11396,N_9583,N_9942);
or U11397 (N_11397,N_8928,N_8150);
nor U11398 (N_11398,N_9313,N_9314);
nor U11399 (N_11399,N_8963,N_8719);
nor U11400 (N_11400,N_8733,N_9040);
nand U11401 (N_11401,N_8514,N_9229);
or U11402 (N_11402,N_9465,N_8206);
and U11403 (N_11403,N_9628,N_9279);
and U11404 (N_11404,N_9402,N_9997);
and U11405 (N_11405,N_8449,N_9737);
nor U11406 (N_11406,N_9861,N_9179);
xnor U11407 (N_11407,N_9706,N_9928);
and U11408 (N_11408,N_8894,N_8855);
nor U11409 (N_11409,N_9767,N_8247);
and U11410 (N_11410,N_9392,N_9428);
nand U11411 (N_11411,N_9068,N_9502);
nor U11412 (N_11412,N_9823,N_8290);
and U11413 (N_11413,N_8522,N_9374);
nor U11414 (N_11414,N_9596,N_9591);
nor U11415 (N_11415,N_8775,N_9123);
nor U11416 (N_11416,N_9764,N_9114);
and U11417 (N_11417,N_8904,N_9608);
xor U11418 (N_11418,N_9847,N_9060);
nand U11419 (N_11419,N_8324,N_9134);
nand U11420 (N_11420,N_8815,N_8206);
and U11421 (N_11421,N_9370,N_8475);
nor U11422 (N_11422,N_9801,N_9270);
or U11423 (N_11423,N_9738,N_9781);
and U11424 (N_11424,N_9427,N_9347);
and U11425 (N_11425,N_8845,N_9585);
and U11426 (N_11426,N_8389,N_9024);
and U11427 (N_11427,N_9373,N_8345);
and U11428 (N_11428,N_9359,N_8553);
or U11429 (N_11429,N_8492,N_8652);
nand U11430 (N_11430,N_8931,N_8790);
nor U11431 (N_11431,N_9256,N_9133);
and U11432 (N_11432,N_8658,N_9059);
and U11433 (N_11433,N_8834,N_9287);
nand U11434 (N_11434,N_8766,N_8850);
nor U11435 (N_11435,N_8402,N_8368);
or U11436 (N_11436,N_8872,N_9201);
or U11437 (N_11437,N_9189,N_9637);
xnor U11438 (N_11438,N_9682,N_9890);
nand U11439 (N_11439,N_8765,N_9908);
nand U11440 (N_11440,N_8317,N_9501);
or U11441 (N_11441,N_9159,N_9453);
and U11442 (N_11442,N_9729,N_8320);
xor U11443 (N_11443,N_8965,N_9990);
nor U11444 (N_11444,N_9523,N_9440);
nor U11445 (N_11445,N_8009,N_8895);
and U11446 (N_11446,N_8898,N_9261);
nor U11447 (N_11447,N_9671,N_9463);
and U11448 (N_11448,N_8169,N_8311);
nand U11449 (N_11449,N_8579,N_9598);
or U11450 (N_11450,N_8828,N_8303);
or U11451 (N_11451,N_8201,N_8052);
xnor U11452 (N_11452,N_9834,N_9486);
and U11453 (N_11453,N_9293,N_8206);
and U11454 (N_11454,N_9212,N_9432);
nand U11455 (N_11455,N_8591,N_8638);
or U11456 (N_11456,N_9706,N_9101);
xor U11457 (N_11457,N_8607,N_8263);
or U11458 (N_11458,N_9063,N_9393);
nor U11459 (N_11459,N_9540,N_9801);
xnor U11460 (N_11460,N_9451,N_8074);
or U11461 (N_11461,N_9442,N_9628);
nor U11462 (N_11462,N_8065,N_9810);
nor U11463 (N_11463,N_8701,N_8239);
nand U11464 (N_11464,N_8538,N_9660);
and U11465 (N_11465,N_9181,N_8933);
nor U11466 (N_11466,N_8896,N_9517);
or U11467 (N_11467,N_8785,N_8744);
nand U11468 (N_11468,N_9742,N_8011);
nor U11469 (N_11469,N_9896,N_9196);
nand U11470 (N_11470,N_8512,N_9826);
or U11471 (N_11471,N_9317,N_9475);
nand U11472 (N_11472,N_9836,N_8886);
nor U11473 (N_11473,N_9037,N_9492);
nor U11474 (N_11474,N_8444,N_8226);
nor U11475 (N_11475,N_8876,N_8864);
or U11476 (N_11476,N_9965,N_9959);
nand U11477 (N_11477,N_9356,N_9622);
or U11478 (N_11478,N_9136,N_8824);
nor U11479 (N_11479,N_9004,N_8209);
nand U11480 (N_11480,N_9888,N_8530);
nor U11481 (N_11481,N_8219,N_9805);
or U11482 (N_11482,N_9340,N_9559);
and U11483 (N_11483,N_8141,N_8190);
xor U11484 (N_11484,N_8886,N_9148);
and U11485 (N_11485,N_8413,N_9774);
xor U11486 (N_11486,N_9551,N_8730);
and U11487 (N_11487,N_8252,N_8221);
nor U11488 (N_11488,N_9702,N_9542);
and U11489 (N_11489,N_9415,N_8267);
nor U11490 (N_11490,N_8893,N_9271);
nor U11491 (N_11491,N_9634,N_8478);
xnor U11492 (N_11492,N_9760,N_9524);
or U11493 (N_11493,N_9702,N_8581);
nand U11494 (N_11494,N_9838,N_8004);
xor U11495 (N_11495,N_9654,N_9933);
nor U11496 (N_11496,N_8488,N_9234);
and U11497 (N_11497,N_9829,N_8862);
xnor U11498 (N_11498,N_9931,N_8430);
or U11499 (N_11499,N_9022,N_8159);
and U11500 (N_11500,N_9047,N_9481);
xor U11501 (N_11501,N_8808,N_8877);
or U11502 (N_11502,N_9051,N_9021);
nor U11503 (N_11503,N_8239,N_8179);
nor U11504 (N_11504,N_8144,N_9586);
or U11505 (N_11505,N_8845,N_9765);
nor U11506 (N_11506,N_9143,N_8532);
nand U11507 (N_11507,N_9920,N_9604);
xnor U11508 (N_11508,N_8180,N_9140);
and U11509 (N_11509,N_8538,N_9154);
or U11510 (N_11510,N_8639,N_8834);
nor U11511 (N_11511,N_8954,N_9424);
and U11512 (N_11512,N_8790,N_8483);
nor U11513 (N_11513,N_8444,N_9390);
or U11514 (N_11514,N_9528,N_9425);
or U11515 (N_11515,N_8574,N_9781);
nor U11516 (N_11516,N_8745,N_9737);
nand U11517 (N_11517,N_8355,N_8356);
nor U11518 (N_11518,N_8536,N_9147);
and U11519 (N_11519,N_9133,N_8081);
and U11520 (N_11520,N_8727,N_9972);
nor U11521 (N_11521,N_9164,N_8604);
nand U11522 (N_11522,N_9494,N_8399);
or U11523 (N_11523,N_9423,N_8634);
nor U11524 (N_11524,N_9335,N_8953);
or U11525 (N_11525,N_9546,N_8075);
and U11526 (N_11526,N_9801,N_8845);
and U11527 (N_11527,N_8787,N_9118);
and U11528 (N_11528,N_8881,N_8112);
or U11529 (N_11529,N_8743,N_8104);
xor U11530 (N_11530,N_8343,N_9778);
nand U11531 (N_11531,N_9394,N_8481);
nor U11532 (N_11532,N_9152,N_8652);
nor U11533 (N_11533,N_9978,N_9844);
or U11534 (N_11534,N_9122,N_9956);
xor U11535 (N_11535,N_8330,N_8015);
nand U11536 (N_11536,N_8562,N_9557);
and U11537 (N_11537,N_8904,N_9156);
nand U11538 (N_11538,N_8985,N_8503);
or U11539 (N_11539,N_8735,N_8820);
xor U11540 (N_11540,N_9871,N_8472);
or U11541 (N_11541,N_9202,N_8230);
and U11542 (N_11542,N_9388,N_9395);
and U11543 (N_11543,N_9851,N_8961);
nand U11544 (N_11544,N_9386,N_9178);
nor U11545 (N_11545,N_9100,N_8775);
nor U11546 (N_11546,N_8803,N_9038);
and U11547 (N_11547,N_8183,N_9581);
xnor U11548 (N_11548,N_8751,N_8174);
nand U11549 (N_11549,N_8689,N_8031);
xnor U11550 (N_11550,N_8799,N_9274);
and U11551 (N_11551,N_9963,N_8801);
or U11552 (N_11552,N_9725,N_9024);
or U11553 (N_11553,N_9178,N_9890);
xnor U11554 (N_11554,N_9981,N_8667);
or U11555 (N_11555,N_9658,N_8163);
or U11556 (N_11556,N_9759,N_9691);
or U11557 (N_11557,N_9450,N_8567);
nand U11558 (N_11558,N_8600,N_8388);
and U11559 (N_11559,N_8492,N_9209);
and U11560 (N_11560,N_9570,N_9491);
nor U11561 (N_11561,N_9706,N_8404);
or U11562 (N_11562,N_9532,N_9959);
nand U11563 (N_11563,N_9469,N_9478);
and U11564 (N_11564,N_9390,N_8826);
or U11565 (N_11565,N_9510,N_9015);
xor U11566 (N_11566,N_8595,N_9928);
nand U11567 (N_11567,N_9814,N_8909);
or U11568 (N_11568,N_8095,N_8119);
nand U11569 (N_11569,N_9004,N_8954);
nand U11570 (N_11570,N_9515,N_9914);
and U11571 (N_11571,N_9910,N_8605);
or U11572 (N_11572,N_8667,N_9736);
xnor U11573 (N_11573,N_9957,N_9971);
nand U11574 (N_11574,N_8095,N_8252);
nor U11575 (N_11575,N_9250,N_9971);
or U11576 (N_11576,N_9270,N_9648);
xor U11577 (N_11577,N_9789,N_9049);
or U11578 (N_11578,N_9072,N_8473);
or U11579 (N_11579,N_8294,N_8291);
xnor U11580 (N_11580,N_9726,N_9384);
nand U11581 (N_11581,N_8256,N_9950);
nand U11582 (N_11582,N_9516,N_9757);
nand U11583 (N_11583,N_9038,N_9186);
and U11584 (N_11584,N_8530,N_8586);
or U11585 (N_11585,N_8314,N_9736);
xor U11586 (N_11586,N_9973,N_9991);
nand U11587 (N_11587,N_8984,N_8440);
and U11588 (N_11588,N_8120,N_8431);
or U11589 (N_11589,N_9779,N_9830);
and U11590 (N_11590,N_9400,N_9354);
nand U11591 (N_11591,N_9867,N_9094);
nor U11592 (N_11592,N_9447,N_8385);
nor U11593 (N_11593,N_9406,N_8441);
nand U11594 (N_11594,N_9351,N_8234);
nor U11595 (N_11595,N_8583,N_9986);
nor U11596 (N_11596,N_9002,N_8481);
nor U11597 (N_11597,N_9528,N_8042);
or U11598 (N_11598,N_8740,N_9046);
nor U11599 (N_11599,N_9922,N_8707);
and U11600 (N_11600,N_9132,N_8843);
nor U11601 (N_11601,N_9310,N_9044);
nor U11602 (N_11602,N_8081,N_9816);
or U11603 (N_11603,N_9293,N_8693);
or U11604 (N_11604,N_8747,N_9486);
nand U11605 (N_11605,N_9952,N_8682);
nand U11606 (N_11606,N_8567,N_9977);
or U11607 (N_11607,N_8487,N_8050);
nand U11608 (N_11608,N_9235,N_8398);
nor U11609 (N_11609,N_9712,N_8103);
and U11610 (N_11610,N_9512,N_8345);
xor U11611 (N_11611,N_8671,N_8012);
nor U11612 (N_11612,N_9749,N_9949);
nor U11613 (N_11613,N_9669,N_9880);
nand U11614 (N_11614,N_9433,N_9518);
xnor U11615 (N_11615,N_9658,N_8539);
and U11616 (N_11616,N_9131,N_9238);
xnor U11617 (N_11617,N_8063,N_8555);
and U11618 (N_11618,N_9526,N_8983);
xnor U11619 (N_11619,N_9164,N_9778);
and U11620 (N_11620,N_9573,N_9753);
nor U11621 (N_11621,N_9311,N_8817);
and U11622 (N_11622,N_8760,N_8776);
nand U11623 (N_11623,N_8332,N_8213);
nand U11624 (N_11624,N_8127,N_8064);
xnor U11625 (N_11625,N_9681,N_8603);
nor U11626 (N_11626,N_9229,N_8869);
nor U11627 (N_11627,N_9900,N_9038);
nor U11628 (N_11628,N_9549,N_9671);
and U11629 (N_11629,N_8492,N_8665);
and U11630 (N_11630,N_8922,N_8554);
and U11631 (N_11631,N_8576,N_9764);
or U11632 (N_11632,N_9576,N_8037);
nor U11633 (N_11633,N_8899,N_8550);
nand U11634 (N_11634,N_9835,N_8851);
and U11635 (N_11635,N_9160,N_8742);
or U11636 (N_11636,N_8375,N_8380);
and U11637 (N_11637,N_9467,N_9707);
and U11638 (N_11638,N_8345,N_9075);
or U11639 (N_11639,N_8720,N_9545);
xor U11640 (N_11640,N_8829,N_8943);
or U11641 (N_11641,N_8460,N_9661);
or U11642 (N_11642,N_9590,N_9515);
nor U11643 (N_11643,N_8060,N_8382);
or U11644 (N_11644,N_9965,N_9075);
xnor U11645 (N_11645,N_8116,N_9360);
and U11646 (N_11646,N_9059,N_8122);
or U11647 (N_11647,N_9671,N_8275);
or U11648 (N_11648,N_8051,N_8306);
xnor U11649 (N_11649,N_8747,N_9407);
or U11650 (N_11650,N_8088,N_9648);
and U11651 (N_11651,N_8494,N_8082);
nand U11652 (N_11652,N_8489,N_9686);
xnor U11653 (N_11653,N_8139,N_8604);
nand U11654 (N_11654,N_9150,N_8086);
xor U11655 (N_11655,N_9372,N_8959);
and U11656 (N_11656,N_9554,N_8321);
and U11657 (N_11657,N_8910,N_8550);
nand U11658 (N_11658,N_9903,N_9569);
or U11659 (N_11659,N_9172,N_8216);
nand U11660 (N_11660,N_9441,N_9320);
nand U11661 (N_11661,N_8076,N_9534);
xnor U11662 (N_11662,N_8034,N_9812);
xor U11663 (N_11663,N_9598,N_9929);
nor U11664 (N_11664,N_9532,N_9053);
nand U11665 (N_11665,N_8711,N_8713);
and U11666 (N_11666,N_9629,N_8099);
nand U11667 (N_11667,N_8760,N_8991);
xor U11668 (N_11668,N_9016,N_8585);
and U11669 (N_11669,N_8503,N_8430);
xor U11670 (N_11670,N_8364,N_8760);
xnor U11671 (N_11671,N_9439,N_8718);
nor U11672 (N_11672,N_8750,N_8472);
nor U11673 (N_11673,N_8163,N_8845);
and U11674 (N_11674,N_8997,N_9789);
nor U11675 (N_11675,N_8482,N_9021);
nor U11676 (N_11676,N_9034,N_9152);
xor U11677 (N_11677,N_9017,N_8261);
nor U11678 (N_11678,N_9005,N_9193);
nand U11679 (N_11679,N_8480,N_9808);
or U11680 (N_11680,N_8563,N_9421);
nand U11681 (N_11681,N_9492,N_8814);
nor U11682 (N_11682,N_8633,N_8725);
nand U11683 (N_11683,N_8132,N_8361);
nor U11684 (N_11684,N_8419,N_9409);
nor U11685 (N_11685,N_9261,N_8454);
nor U11686 (N_11686,N_8302,N_8280);
xnor U11687 (N_11687,N_8890,N_9408);
xor U11688 (N_11688,N_9931,N_9035);
or U11689 (N_11689,N_9697,N_9021);
nand U11690 (N_11690,N_9375,N_9302);
xor U11691 (N_11691,N_9402,N_8595);
or U11692 (N_11692,N_9696,N_8613);
nand U11693 (N_11693,N_9235,N_9963);
xnor U11694 (N_11694,N_9646,N_8886);
and U11695 (N_11695,N_9718,N_8823);
nand U11696 (N_11696,N_9654,N_9750);
nand U11697 (N_11697,N_8642,N_9156);
or U11698 (N_11698,N_8539,N_9087);
and U11699 (N_11699,N_9525,N_8416);
nand U11700 (N_11700,N_8404,N_9154);
or U11701 (N_11701,N_8976,N_8114);
xor U11702 (N_11702,N_9272,N_9642);
and U11703 (N_11703,N_8309,N_8889);
nand U11704 (N_11704,N_9702,N_9410);
and U11705 (N_11705,N_8150,N_8101);
nor U11706 (N_11706,N_9307,N_8976);
or U11707 (N_11707,N_8764,N_8407);
nand U11708 (N_11708,N_8733,N_8065);
and U11709 (N_11709,N_9626,N_8899);
nand U11710 (N_11710,N_8253,N_8922);
xnor U11711 (N_11711,N_8866,N_9666);
xnor U11712 (N_11712,N_8129,N_8038);
and U11713 (N_11713,N_9421,N_9759);
xnor U11714 (N_11714,N_9454,N_8840);
nand U11715 (N_11715,N_8651,N_8208);
xor U11716 (N_11716,N_8261,N_9399);
xnor U11717 (N_11717,N_9707,N_8602);
nand U11718 (N_11718,N_8067,N_8463);
xnor U11719 (N_11719,N_8185,N_9661);
xnor U11720 (N_11720,N_9330,N_9632);
xor U11721 (N_11721,N_8524,N_9208);
nor U11722 (N_11722,N_8570,N_8668);
or U11723 (N_11723,N_9607,N_9627);
nand U11724 (N_11724,N_9793,N_8499);
and U11725 (N_11725,N_8283,N_8896);
or U11726 (N_11726,N_9212,N_8220);
nand U11727 (N_11727,N_9942,N_8800);
nand U11728 (N_11728,N_8588,N_8882);
or U11729 (N_11729,N_9370,N_9049);
nand U11730 (N_11730,N_8566,N_8713);
or U11731 (N_11731,N_8349,N_9305);
nand U11732 (N_11732,N_9053,N_9038);
nor U11733 (N_11733,N_8366,N_9677);
nor U11734 (N_11734,N_8221,N_8995);
nand U11735 (N_11735,N_8930,N_9285);
nand U11736 (N_11736,N_8674,N_9852);
nand U11737 (N_11737,N_9231,N_8957);
or U11738 (N_11738,N_8574,N_8591);
xnor U11739 (N_11739,N_9439,N_8148);
nand U11740 (N_11740,N_9815,N_9793);
nand U11741 (N_11741,N_9250,N_8607);
and U11742 (N_11742,N_8200,N_9855);
nand U11743 (N_11743,N_8941,N_9883);
or U11744 (N_11744,N_8557,N_9276);
nand U11745 (N_11745,N_9888,N_9500);
nor U11746 (N_11746,N_9972,N_9010);
nand U11747 (N_11747,N_8978,N_8708);
nor U11748 (N_11748,N_8792,N_9570);
or U11749 (N_11749,N_9680,N_9559);
or U11750 (N_11750,N_9662,N_9568);
or U11751 (N_11751,N_9800,N_8479);
nand U11752 (N_11752,N_9279,N_8769);
nor U11753 (N_11753,N_8134,N_8600);
nand U11754 (N_11754,N_8284,N_8985);
nor U11755 (N_11755,N_9515,N_8298);
and U11756 (N_11756,N_9273,N_8694);
nand U11757 (N_11757,N_9187,N_8192);
xor U11758 (N_11758,N_8343,N_8313);
nand U11759 (N_11759,N_9339,N_9901);
nor U11760 (N_11760,N_8816,N_9858);
nand U11761 (N_11761,N_9595,N_8852);
xnor U11762 (N_11762,N_8895,N_8301);
nand U11763 (N_11763,N_9770,N_8818);
and U11764 (N_11764,N_9791,N_8428);
or U11765 (N_11765,N_9039,N_8908);
and U11766 (N_11766,N_8879,N_8355);
xnor U11767 (N_11767,N_9963,N_8285);
or U11768 (N_11768,N_8416,N_9918);
nor U11769 (N_11769,N_8006,N_9460);
or U11770 (N_11770,N_9939,N_8479);
nand U11771 (N_11771,N_9944,N_9362);
nor U11772 (N_11772,N_9425,N_8312);
xor U11773 (N_11773,N_8273,N_8696);
or U11774 (N_11774,N_9546,N_8415);
nor U11775 (N_11775,N_8428,N_8211);
xnor U11776 (N_11776,N_8883,N_8353);
or U11777 (N_11777,N_8377,N_8950);
or U11778 (N_11778,N_8163,N_9820);
xnor U11779 (N_11779,N_9179,N_8324);
nor U11780 (N_11780,N_8145,N_8635);
nor U11781 (N_11781,N_9793,N_9675);
nor U11782 (N_11782,N_8792,N_8504);
nand U11783 (N_11783,N_8988,N_9828);
xnor U11784 (N_11784,N_8067,N_9616);
and U11785 (N_11785,N_8289,N_8245);
and U11786 (N_11786,N_9913,N_8223);
nor U11787 (N_11787,N_8352,N_8454);
and U11788 (N_11788,N_9358,N_9959);
or U11789 (N_11789,N_8146,N_9547);
xnor U11790 (N_11790,N_9039,N_9407);
nand U11791 (N_11791,N_9702,N_9439);
nand U11792 (N_11792,N_8330,N_8365);
nand U11793 (N_11793,N_9623,N_8523);
nor U11794 (N_11794,N_9138,N_8811);
and U11795 (N_11795,N_9274,N_9612);
xor U11796 (N_11796,N_8962,N_8039);
nand U11797 (N_11797,N_8225,N_8072);
or U11798 (N_11798,N_9895,N_8514);
and U11799 (N_11799,N_9109,N_8558);
xnor U11800 (N_11800,N_8197,N_8151);
or U11801 (N_11801,N_8871,N_9115);
nand U11802 (N_11802,N_9816,N_9341);
or U11803 (N_11803,N_8935,N_8172);
xnor U11804 (N_11804,N_8682,N_9759);
xor U11805 (N_11805,N_9505,N_9653);
xor U11806 (N_11806,N_9223,N_9081);
nand U11807 (N_11807,N_9140,N_9498);
nor U11808 (N_11808,N_9451,N_8906);
xor U11809 (N_11809,N_8176,N_8988);
or U11810 (N_11810,N_9125,N_8490);
nand U11811 (N_11811,N_8835,N_9146);
nor U11812 (N_11812,N_8957,N_9422);
or U11813 (N_11813,N_8676,N_9702);
nand U11814 (N_11814,N_8183,N_8697);
and U11815 (N_11815,N_8314,N_9405);
or U11816 (N_11816,N_9415,N_9267);
or U11817 (N_11817,N_8045,N_8019);
xor U11818 (N_11818,N_8171,N_9023);
xor U11819 (N_11819,N_9710,N_8601);
nand U11820 (N_11820,N_8774,N_9339);
nor U11821 (N_11821,N_9340,N_8310);
nor U11822 (N_11822,N_8175,N_8513);
and U11823 (N_11823,N_8114,N_9855);
xnor U11824 (N_11824,N_8197,N_8131);
nand U11825 (N_11825,N_9204,N_9150);
nor U11826 (N_11826,N_9959,N_9538);
nand U11827 (N_11827,N_8925,N_9325);
and U11828 (N_11828,N_9042,N_9276);
and U11829 (N_11829,N_8985,N_9197);
and U11830 (N_11830,N_8120,N_9322);
xor U11831 (N_11831,N_8283,N_9452);
or U11832 (N_11832,N_9088,N_9862);
nor U11833 (N_11833,N_8226,N_8090);
nand U11834 (N_11834,N_8086,N_9016);
nand U11835 (N_11835,N_9267,N_8084);
xnor U11836 (N_11836,N_9568,N_9802);
and U11837 (N_11837,N_8757,N_8020);
and U11838 (N_11838,N_9884,N_9997);
xnor U11839 (N_11839,N_8299,N_8366);
nor U11840 (N_11840,N_8967,N_9440);
nand U11841 (N_11841,N_8044,N_8397);
and U11842 (N_11842,N_9221,N_9475);
xor U11843 (N_11843,N_8372,N_8743);
xor U11844 (N_11844,N_8768,N_8460);
and U11845 (N_11845,N_8437,N_8644);
or U11846 (N_11846,N_8127,N_9757);
nor U11847 (N_11847,N_9894,N_8778);
and U11848 (N_11848,N_9593,N_9024);
nor U11849 (N_11849,N_9715,N_9376);
xnor U11850 (N_11850,N_9848,N_9120);
nand U11851 (N_11851,N_8113,N_9615);
nor U11852 (N_11852,N_9604,N_8151);
and U11853 (N_11853,N_8162,N_9296);
and U11854 (N_11854,N_9870,N_9742);
nand U11855 (N_11855,N_9719,N_9055);
nor U11856 (N_11856,N_8284,N_8735);
xnor U11857 (N_11857,N_9559,N_9770);
or U11858 (N_11858,N_8974,N_9027);
nand U11859 (N_11859,N_8314,N_8547);
nand U11860 (N_11860,N_9529,N_9349);
nor U11861 (N_11861,N_8084,N_9373);
and U11862 (N_11862,N_8478,N_8831);
or U11863 (N_11863,N_9638,N_8924);
xor U11864 (N_11864,N_8462,N_9599);
xor U11865 (N_11865,N_9928,N_9115);
xor U11866 (N_11866,N_8081,N_9337);
nand U11867 (N_11867,N_8151,N_9235);
nand U11868 (N_11868,N_9328,N_9740);
xnor U11869 (N_11869,N_8049,N_9049);
and U11870 (N_11870,N_9574,N_8701);
xnor U11871 (N_11871,N_8239,N_8193);
or U11872 (N_11872,N_8313,N_8786);
or U11873 (N_11873,N_8277,N_8373);
xnor U11874 (N_11874,N_9315,N_9056);
xnor U11875 (N_11875,N_9406,N_9268);
xnor U11876 (N_11876,N_9576,N_8639);
xor U11877 (N_11877,N_9232,N_9879);
and U11878 (N_11878,N_9014,N_8073);
nand U11879 (N_11879,N_9291,N_8925);
or U11880 (N_11880,N_8942,N_9896);
nand U11881 (N_11881,N_9156,N_8963);
and U11882 (N_11882,N_9422,N_9373);
nand U11883 (N_11883,N_8909,N_9033);
xnor U11884 (N_11884,N_9405,N_9897);
or U11885 (N_11885,N_9608,N_9175);
and U11886 (N_11886,N_9038,N_8313);
and U11887 (N_11887,N_9243,N_8790);
or U11888 (N_11888,N_8153,N_8204);
and U11889 (N_11889,N_8156,N_9464);
or U11890 (N_11890,N_8478,N_8447);
and U11891 (N_11891,N_9505,N_8665);
xor U11892 (N_11892,N_9067,N_9812);
nor U11893 (N_11893,N_9327,N_9637);
nand U11894 (N_11894,N_8285,N_8742);
and U11895 (N_11895,N_8119,N_9950);
xnor U11896 (N_11896,N_9663,N_8060);
or U11897 (N_11897,N_9407,N_9055);
and U11898 (N_11898,N_8121,N_8890);
xor U11899 (N_11899,N_8527,N_9967);
xor U11900 (N_11900,N_9397,N_9046);
xnor U11901 (N_11901,N_8389,N_8679);
nand U11902 (N_11902,N_9673,N_9762);
and U11903 (N_11903,N_8868,N_8443);
or U11904 (N_11904,N_9606,N_9127);
or U11905 (N_11905,N_8172,N_9109);
or U11906 (N_11906,N_9915,N_8520);
or U11907 (N_11907,N_8950,N_9925);
xnor U11908 (N_11908,N_9283,N_8021);
xnor U11909 (N_11909,N_9717,N_9465);
nand U11910 (N_11910,N_8115,N_9978);
or U11911 (N_11911,N_8644,N_9216);
xnor U11912 (N_11912,N_8675,N_8731);
xnor U11913 (N_11913,N_9069,N_9580);
nand U11914 (N_11914,N_8833,N_8786);
xor U11915 (N_11915,N_8060,N_9469);
and U11916 (N_11916,N_9818,N_9440);
xor U11917 (N_11917,N_8648,N_9524);
and U11918 (N_11918,N_8332,N_9059);
xor U11919 (N_11919,N_8718,N_9038);
xnor U11920 (N_11920,N_9746,N_8826);
nand U11921 (N_11921,N_8569,N_9595);
or U11922 (N_11922,N_8001,N_8902);
xnor U11923 (N_11923,N_8975,N_9792);
xnor U11924 (N_11924,N_9342,N_8969);
nor U11925 (N_11925,N_8486,N_8957);
and U11926 (N_11926,N_8538,N_8341);
or U11927 (N_11927,N_8107,N_8870);
or U11928 (N_11928,N_8133,N_8769);
nand U11929 (N_11929,N_8849,N_8583);
or U11930 (N_11930,N_8946,N_8073);
and U11931 (N_11931,N_9000,N_9045);
and U11932 (N_11932,N_8373,N_9816);
nor U11933 (N_11933,N_9841,N_8625);
nor U11934 (N_11934,N_9032,N_9436);
nor U11935 (N_11935,N_9812,N_9429);
xor U11936 (N_11936,N_9808,N_9342);
and U11937 (N_11937,N_8706,N_8389);
and U11938 (N_11938,N_8454,N_9228);
and U11939 (N_11939,N_8983,N_9967);
nand U11940 (N_11940,N_8392,N_9872);
nor U11941 (N_11941,N_9059,N_8473);
nand U11942 (N_11942,N_9751,N_9814);
nand U11943 (N_11943,N_8847,N_8168);
xnor U11944 (N_11944,N_8375,N_8249);
nand U11945 (N_11945,N_8708,N_9922);
xor U11946 (N_11946,N_9995,N_9901);
or U11947 (N_11947,N_8815,N_9194);
and U11948 (N_11948,N_8978,N_8743);
or U11949 (N_11949,N_9207,N_9663);
or U11950 (N_11950,N_9341,N_8412);
nand U11951 (N_11951,N_9579,N_9517);
and U11952 (N_11952,N_9996,N_8268);
or U11953 (N_11953,N_9046,N_8034);
or U11954 (N_11954,N_9960,N_9839);
nor U11955 (N_11955,N_9045,N_9112);
and U11956 (N_11956,N_8654,N_8770);
or U11957 (N_11957,N_9039,N_9377);
nor U11958 (N_11958,N_8624,N_8696);
and U11959 (N_11959,N_9596,N_8874);
or U11960 (N_11960,N_8425,N_9855);
xor U11961 (N_11961,N_9080,N_9558);
and U11962 (N_11962,N_9631,N_8914);
nor U11963 (N_11963,N_8823,N_8688);
or U11964 (N_11964,N_8231,N_9691);
or U11965 (N_11965,N_8884,N_8054);
or U11966 (N_11966,N_9544,N_8099);
and U11967 (N_11967,N_8210,N_8647);
nor U11968 (N_11968,N_9162,N_8759);
nor U11969 (N_11969,N_8831,N_8532);
nor U11970 (N_11970,N_9946,N_8873);
xor U11971 (N_11971,N_9399,N_9802);
or U11972 (N_11972,N_9566,N_9797);
xor U11973 (N_11973,N_9751,N_8441);
nor U11974 (N_11974,N_9515,N_8150);
nor U11975 (N_11975,N_9035,N_8264);
xor U11976 (N_11976,N_8410,N_9796);
xor U11977 (N_11977,N_8833,N_9143);
nand U11978 (N_11978,N_8414,N_9909);
nand U11979 (N_11979,N_8858,N_8924);
nand U11980 (N_11980,N_9096,N_8875);
or U11981 (N_11981,N_9161,N_9719);
xnor U11982 (N_11982,N_9178,N_8469);
or U11983 (N_11983,N_9011,N_8442);
and U11984 (N_11984,N_8629,N_8418);
nand U11985 (N_11985,N_8871,N_8128);
nand U11986 (N_11986,N_9227,N_8216);
nand U11987 (N_11987,N_8701,N_9730);
nand U11988 (N_11988,N_9930,N_8514);
or U11989 (N_11989,N_9868,N_8086);
xor U11990 (N_11990,N_9320,N_9863);
nand U11991 (N_11991,N_8107,N_8938);
and U11992 (N_11992,N_8394,N_9347);
xnor U11993 (N_11993,N_8502,N_8550);
and U11994 (N_11994,N_9470,N_8820);
nor U11995 (N_11995,N_8941,N_8963);
and U11996 (N_11996,N_8972,N_9156);
nand U11997 (N_11997,N_8572,N_9083);
or U11998 (N_11998,N_9678,N_9193);
nor U11999 (N_11999,N_8485,N_8023);
nand U12000 (N_12000,N_10217,N_10521);
xor U12001 (N_12001,N_10032,N_11595);
nor U12002 (N_12002,N_11237,N_10092);
and U12003 (N_12003,N_10837,N_11824);
xor U12004 (N_12004,N_11800,N_10757);
and U12005 (N_12005,N_10879,N_11869);
and U12006 (N_12006,N_10011,N_10216);
nand U12007 (N_12007,N_11296,N_11113);
nand U12008 (N_12008,N_11329,N_10138);
xor U12009 (N_12009,N_10730,N_10401);
xnor U12010 (N_12010,N_10386,N_11611);
nor U12011 (N_12011,N_11600,N_11517);
or U12012 (N_12012,N_10589,N_11487);
and U12013 (N_12013,N_11854,N_10617);
or U12014 (N_12014,N_10137,N_10173);
or U12015 (N_12015,N_10736,N_10029);
nand U12016 (N_12016,N_11432,N_11683);
xnor U12017 (N_12017,N_10647,N_10670);
or U12018 (N_12018,N_11986,N_11837);
xor U12019 (N_12019,N_10315,N_11176);
xor U12020 (N_12020,N_10447,N_11424);
and U12021 (N_12021,N_11377,N_11759);
or U12022 (N_12022,N_11575,N_11499);
or U12023 (N_12023,N_10362,N_10595);
and U12024 (N_12024,N_11642,N_10165);
nand U12025 (N_12025,N_10363,N_11395);
nand U12026 (N_12026,N_11425,N_10506);
or U12027 (N_12027,N_11646,N_11262);
nor U12028 (N_12028,N_11875,N_11579);
xnor U12029 (N_12029,N_10466,N_11334);
and U12030 (N_12030,N_10831,N_10596);
nand U12031 (N_12031,N_10820,N_10365);
xnor U12032 (N_12032,N_11051,N_11735);
nor U12033 (N_12033,N_10225,N_11355);
xor U12034 (N_12034,N_10327,N_10373);
and U12035 (N_12035,N_10944,N_11239);
nand U12036 (N_12036,N_11586,N_11682);
nand U12037 (N_12037,N_10220,N_10110);
xnor U12038 (N_12038,N_11242,N_10369);
xor U12039 (N_12039,N_11382,N_11036);
or U12040 (N_12040,N_11139,N_10146);
nand U12041 (N_12041,N_11401,N_11736);
and U12042 (N_12042,N_10525,N_10295);
nand U12043 (N_12043,N_10324,N_11946);
and U12044 (N_12044,N_11005,N_11535);
and U12045 (N_12045,N_10231,N_11099);
xnor U12046 (N_12046,N_10815,N_11598);
xnor U12047 (N_12047,N_10697,N_11229);
nor U12048 (N_12048,N_11378,N_10250);
xor U12049 (N_12049,N_11158,N_11720);
xor U12050 (N_12050,N_10177,N_11591);
and U12051 (N_12051,N_11650,N_11443);
or U12052 (N_12052,N_10323,N_11997);
xnor U12053 (N_12053,N_10667,N_10824);
nor U12054 (N_12054,N_10080,N_11070);
xnor U12055 (N_12055,N_11008,N_11449);
or U12056 (N_12056,N_10314,N_11033);
or U12057 (N_12057,N_11776,N_11961);
and U12058 (N_12058,N_10618,N_11657);
and U12059 (N_12059,N_11190,N_11474);
nor U12060 (N_12060,N_11612,N_11659);
or U12061 (N_12061,N_10724,N_11688);
and U12062 (N_12062,N_11536,N_11872);
or U12063 (N_12063,N_10266,N_11325);
nand U12064 (N_12064,N_10756,N_11696);
and U12065 (N_12065,N_11290,N_10611);
nor U12066 (N_12066,N_10883,N_10119);
nand U12067 (N_12067,N_11321,N_11938);
or U12068 (N_12068,N_10869,N_11057);
or U12069 (N_12069,N_11301,N_11669);
or U12070 (N_12070,N_11898,N_11153);
or U12071 (N_12071,N_10790,N_10579);
and U12072 (N_12072,N_10406,N_10052);
nor U12073 (N_12073,N_10583,N_11966);
and U12074 (N_12074,N_11471,N_10574);
nor U12075 (N_12075,N_11857,N_10448);
or U12076 (N_12076,N_11253,N_10560);
or U12077 (N_12077,N_11364,N_11353);
and U12078 (N_12078,N_11210,N_11677);
nand U12079 (N_12079,N_11891,N_11529);
nor U12080 (N_12080,N_11760,N_11721);
nand U12081 (N_12081,N_11170,N_10278);
xor U12082 (N_12082,N_11465,N_10361);
and U12083 (N_12083,N_11254,N_10294);
nor U12084 (N_12084,N_10038,N_11808);
nor U12085 (N_12085,N_10704,N_11422);
xor U12086 (N_12086,N_10115,N_11665);
nand U12087 (N_12087,N_10750,N_11151);
xor U12088 (N_12088,N_10874,N_10972);
xor U12089 (N_12089,N_10843,N_10908);
and U12090 (N_12090,N_10580,N_11435);
nand U12091 (N_12091,N_10097,N_10631);
and U12092 (N_12092,N_10603,N_10546);
nor U12093 (N_12093,N_11624,N_11480);
xnor U12094 (N_12094,N_10798,N_11410);
and U12095 (N_12095,N_10243,N_10805);
nor U12096 (N_12096,N_10239,N_11715);
nand U12097 (N_12097,N_10850,N_11848);
nand U12098 (N_12098,N_10348,N_10274);
or U12099 (N_12099,N_10460,N_10399);
or U12100 (N_12100,N_11813,N_10985);
nor U12101 (N_12101,N_10811,N_11178);
nand U12102 (N_12102,N_11928,N_11116);
nand U12103 (N_12103,N_11668,N_10427);
and U12104 (N_12104,N_11658,N_10979);
or U12105 (N_12105,N_10069,N_10451);
and U12106 (N_12106,N_11980,N_11552);
xnor U12107 (N_12107,N_10718,N_11032);
and U12108 (N_12108,N_10727,N_11020);
and U12109 (N_12109,N_11128,N_10488);
xor U12110 (N_12110,N_11147,N_10566);
xor U12111 (N_12111,N_10584,N_11880);
or U12112 (N_12112,N_11939,N_10997);
or U12113 (N_12113,N_11630,N_10691);
nand U12114 (N_12114,N_10233,N_11693);
and U12115 (N_12115,N_10792,N_10818);
or U12116 (N_12116,N_11098,N_10986);
nor U12117 (N_12117,N_10331,N_11007);
and U12118 (N_12118,N_11962,N_11701);
xnor U12119 (N_12119,N_11492,N_11916);
nand U12120 (N_12120,N_11930,N_10206);
nand U12121 (N_12121,N_11900,N_10089);
and U12122 (N_12122,N_10397,N_10507);
nor U12123 (N_12123,N_11732,N_11040);
xnor U12124 (N_12124,N_11285,N_10433);
xor U12125 (N_12125,N_10517,N_10957);
and U12126 (N_12126,N_11617,N_10126);
and U12127 (N_12127,N_10135,N_11590);
and U12128 (N_12128,N_10129,N_11063);
and U12129 (N_12129,N_11416,N_10413);
xor U12130 (N_12130,N_11100,N_10454);
xnor U12131 (N_12131,N_11649,N_11507);
nand U12132 (N_12132,N_11518,N_11015);
and U12133 (N_12133,N_10856,N_10846);
xnor U12134 (N_12134,N_10533,N_10068);
xor U12135 (N_12135,N_10558,N_10376);
or U12136 (N_12136,N_11025,N_10844);
and U12137 (N_12137,N_10588,N_11264);
and U12138 (N_12138,N_11896,N_11951);
and U12139 (N_12139,N_11358,N_10563);
xor U12140 (N_12140,N_10190,N_11613);
xnor U12141 (N_12141,N_11685,N_10031);
nor U12142 (N_12142,N_11684,N_10728);
or U12143 (N_12143,N_10495,N_10019);
nor U12144 (N_12144,N_11194,N_10561);
and U12145 (N_12145,N_11046,N_11545);
and U12146 (N_12146,N_10802,N_10240);
and U12147 (N_12147,N_10259,N_10938);
nand U12148 (N_12148,N_11494,N_10030);
and U12149 (N_12149,N_10419,N_11910);
xnor U12150 (N_12150,N_11431,N_10576);
nand U12151 (N_12151,N_11868,N_11490);
or U12152 (N_12152,N_10567,N_11862);
or U12153 (N_12153,N_11690,N_10484);
or U12154 (N_12154,N_10270,N_11454);
xnor U12155 (N_12155,N_11220,N_10304);
and U12156 (N_12156,N_11905,N_11346);
or U12157 (N_12157,N_10439,N_10519);
and U12158 (N_12158,N_10890,N_11212);
nor U12159 (N_12159,N_11469,N_10594);
nand U12160 (N_12160,N_11300,N_11433);
or U12161 (N_12161,N_10998,N_10022);
and U12162 (N_12162,N_10570,N_10077);
nand U12163 (N_12163,N_10035,N_11619);
nor U12164 (N_12164,N_11095,N_10497);
nand U12165 (N_12165,N_11281,N_11949);
nor U12166 (N_12166,N_11342,N_11618);
and U12167 (N_12167,N_10087,N_11144);
xor U12168 (N_12168,N_11884,N_10208);
xor U12169 (N_12169,N_11127,N_10659);
nor U12170 (N_12170,N_11064,N_11430);
xnor U12171 (N_12171,N_11833,N_11394);
or U12172 (N_12172,N_11597,N_10255);
nand U12173 (N_12173,N_11805,N_11204);
xnor U12174 (N_12174,N_10573,N_10139);
xor U12175 (N_12175,N_10449,N_11687);
or U12176 (N_12176,N_11981,N_10426);
xnor U12177 (N_12177,N_10131,N_11525);
and U12178 (N_12178,N_10272,N_11909);
nand U12179 (N_12179,N_11562,N_11198);
or U12180 (N_12180,N_10234,N_10287);
nor U12181 (N_12181,N_11581,N_11014);
and U12182 (N_12182,N_11234,N_11415);
xnor U12183 (N_12183,N_10298,N_11041);
and U12184 (N_12184,N_11052,N_10403);
or U12185 (N_12185,N_11976,N_10857);
xnor U12186 (N_12186,N_10422,N_11527);
or U12187 (N_12187,N_11705,N_10641);
and U12188 (N_12188,N_10524,N_10425);
xnor U12189 (N_12189,N_11027,N_11344);
nor U12190 (N_12190,N_11149,N_10123);
and U12191 (N_12191,N_10329,N_11692);
nor U12192 (N_12192,N_11573,N_10776);
xnor U12193 (N_12193,N_10926,N_11266);
or U12194 (N_12194,N_10710,N_10302);
xor U12195 (N_12195,N_10917,N_10597);
nor U12196 (N_12196,N_10630,N_11973);
or U12197 (N_12197,N_11140,N_11870);
nor U12198 (N_12198,N_11944,N_11023);
nor U12199 (N_12199,N_10352,N_11024);
nor U12200 (N_12200,N_11460,N_11162);
nand U12201 (N_12201,N_11123,N_11785);
nor U12202 (N_12202,N_11817,N_10181);
or U12203 (N_12203,N_11643,N_10411);
xnor U12204 (N_12204,N_11273,N_10207);
and U12205 (N_12205,N_11967,N_11689);
and U12206 (N_12206,N_10404,N_10799);
and U12207 (N_12207,N_10714,N_10845);
nand U12208 (N_12208,N_11164,N_10292);
or U12209 (N_12209,N_10531,N_10388);
xnor U12210 (N_12210,N_10765,N_11505);
or U12211 (N_12211,N_11935,N_10340);
nand U12212 (N_12212,N_11495,N_11724);
xnor U12213 (N_12213,N_10334,N_10513);
xnor U12214 (N_12214,N_11082,N_11085);
nand U12215 (N_12215,N_11769,N_10347);
nor U12216 (N_12216,N_10078,N_10158);
nor U12217 (N_12217,N_10389,N_10796);
nand U12218 (N_12218,N_11777,N_11216);
and U12219 (N_12219,N_11340,N_11404);
and U12220 (N_12220,N_10410,N_11578);
xnor U12221 (N_12221,N_10627,N_11634);
or U12222 (N_12222,N_11514,N_11902);
xor U12223 (N_12223,N_10241,N_11468);
nand U12224 (N_12224,N_10509,N_10142);
nor U12225 (N_12225,N_11592,N_10854);
nor U12226 (N_12226,N_11791,N_11241);
and U12227 (N_12227,N_10434,N_11637);
nor U12228 (N_12228,N_11335,N_11115);
nor U12229 (N_12229,N_10505,N_10203);
nor U12230 (N_12230,N_11661,N_11933);
nor U12231 (N_12231,N_10620,N_11803);
xnor U12232 (N_12232,N_11067,N_11625);
nor U12233 (N_12233,N_10305,N_11411);
and U12234 (N_12234,N_10248,N_11038);
and U12235 (N_12235,N_11680,N_11143);
or U12236 (N_12236,N_11319,N_10600);
nand U12237 (N_12237,N_10933,N_10858);
nor U12238 (N_12238,N_10064,N_10366);
nor U12239 (N_12239,N_11062,N_10187);
nor U12240 (N_12240,N_10868,N_10375);
and U12241 (N_12241,N_10694,N_11493);
nand U12242 (N_12242,N_11899,N_11440);
xnor U12243 (N_12243,N_11927,N_10923);
xnor U12244 (N_12244,N_10554,N_10830);
xnor U12245 (N_12245,N_10984,N_11801);
nand U12246 (N_12246,N_10742,N_10380);
xnor U12247 (N_12247,N_10499,N_10585);
and U12248 (N_12248,N_11137,N_10812);
xor U12249 (N_12249,N_10920,N_11858);
and U12250 (N_12250,N_11974,N_11093);
or U12251 (N_12251,N_11631,N_10456);
nor U12252 (N_12252,N_11039,N_10127);
or U12253 (N_12253,N_10477,N_10381);
nand U12254 (N_12254,N_11950,N_10819);
or U12255 (N_12255,N_11538,N_10117);
xor U12256 (N_12256,N_11714,N_10669);
or U12257 (N_12257,N_10145,N_11742);
nor U12258 (N_12258,N_11171,N_11125);
nor U12259 (N_12259,N_11716,N_10023);
and U12260 (N_12260,N_11348,N_10632);
nor U12261 (N_12261,N_11269,N_10467);
and U12262 (N_12262,N_11350,N_11882);
or U12263 (N_12263,N_10515,N_10464);
or U12264 (N_12264,N_10424,N_10940);
or U12265 (N_12265,N_11345,N_11810);
xnor U12266 (N_12266,N_10085,N_11305);
or U12267 (N_12267,N_10120,N_11585);
or U12268 (N_12268,N_11488,N_10510);
xnor U12269 (N_12269,N_11712,N_10800);
nor U12270 (N_12270,N_10128,N_10476);
and U12271 (N_12271,N_11989,N_10823);
xnor U12272 (N_12272,N_10599,N_11531);
nor U12273 (N_12273,N_11840,N_10921);
nor U12274 (N_12274,N_11897,N_10125);
xor U12275 (N_12275,N_11456,N_10354);
nand U12276 (N_12276,N_11504,N_10981);
xnor U12277 (N_12277,N_11632,N_10260);
nand U12278 (N_12278,N_10209,N_10096);
xnor U12279 (N_12279,N_10257,N_10319);
nor U12280 (N_12280,N_11926,N_10478);
or U12281 (N_12281,N_11744,N_11920);
or U12282 (N_12282,N_10199,N_10429);
and U12283 (N_12283,N_10547,N_10614);
xnor U12284 (N_12284,N_10849,N_10452);
or U12285 (N_12285,N_10283,N_11663);
and U12286 (N_12286,N_10414,N_11112);
or U12287 (N_12287,N_10288,N_10212);
nand U12288 (N_12288,N_10913,N_11741);
nor U12289 (N_12289,N_11486,N_10191);
and U12290 (N_12290,N_10291,N_11011);
xnor U12291 (N_12291,N_10744,N_10832);
xnor U12292 (N_12292,N_11703,N_10677);
xnor U12293 (N_12293,N_11574,N_11271);
nor U12294 (N_12294,N_10925,N_11277);
and U12295 (N_12295,N_11357,N_10176);
and U12296 (N_12296,N_11207,N_11437);
xor U12297 (N_12297,N_10383,N_10061);
xnor U12298 (N_12298,N_10320,N_10624);
nand U12299 (N_12299,N_11850,N_11044);
nand U12300 (N_12300,N_10564,N_10775);
nor U12301 (N_12301,N_11075,N_10277);
xor U12302 (N_12302,N_11396,N_10312);
nand U12303 (N_12303,N_11569,N_11626);
xor U12304 (N_12304,N_11349,N_11594);
or U12305 (N_12305,N_11111,N_11268);
xor U12306 (N_12306,N_10643,N_10771);
and U12307 (N_12307,N_11155,N_11955);
nand U12308 (N_12308,N_10947,N_10688);
or U12309 (N_12309,N_10695,N_11278);
and U12310 (N_12310,N_10934,N_11936);
and U12311 (N_12311,N_11104,N_10379);
or U12312 (N_12312,N_11026,N_10167);
or U12313 (N_12313,N_10322,N_11609);
or U12314 (N_12314,N_10218,N_11699);
xor U12315 (N_12315,N_11423,N_11713);
and U12316 (N_12316,N_10057,N_11148);
nand U12317 (N_12317,N_11169,N_11876);
nand U12318 (N_12318,N_11530,N_10578);
or U12319 (N_12319,N_10793,N_10109);
xor U12320 (N_12320,N_10747,N_10680);
and U12321 (N_12321,N_10102,N_11879);
nand U12322 (N_12322,N_10058,N_10968);
or U12323 (N_12323,N_10651,N_10678);
xnor U12324 (N_12324,N_10027,N_11131);
and U12325 (N_12325,N_11292,N_10893);
nand U12326 (N_12326,N_10945,N_10723);
nand U12327 (N_12327,N_10044,N_10784);
xnor U12328 (N_12328,N_11390,N_11546);
xor U12329 (N_12329,N_10939,N_11621);
xnor U12330 (N_12330,N_10619,N_11445);
nand U12331 (N_12331,N_10518,N_10071);
nand U12332 (N_12332,N_11751,N_10999);
or U12333 (N_12333,N_10418,N_10350);
nor U12334 (N_12334,N_10671,N_11819);
nor U12335 (N_12335,N_11218,N_10219);
and U12336 (N_12336,N_11351,N_11758);
xnor U12337 (N_12337,N_11385,N_10457);
and U12338 (N_12338,N_10821,N_10729);
nor U12339 (N_12339,N_10280,N_10178);
nor U12340 (N_12340,N_10663,N_10001);
nand U12341 (N_12341,N_11602,N_10221);
nand U12342 (N_12342,N_11477,N_11794);
xor U12343 (N_12343,N_10084,N_11219);
or U12344 (N_12344,N_10244,N_10014);
or U12345 (N_12345,N_10400,N_10367);
nand U12346 (N_12346,N_11931,N_10701);
nor U12347 (N_12347,N_10215,N_10889);
or U12348 (N_12348,N_11640,N_11745);
nand U12349 (N_12349,N_11167,N_11419);
xnor U12350 (N_12350,N_11109,N_10358);
and U12351 (N_12351,N_11089,N_10196);
nand U12352 (N_12352,N_10059,N_11359);
or U12353 (N_12353,N_10861,N_11746);
or U12354 (N_12354,N_11244,N_11584);
nor U12355 (N_12355,N_10664,N_11077);
nor U12356 (N_12356,N_10872,N_10734);
xor U12357 (N_12357,N_10970,N_10770);
nor U12358 (N_12358,N_11387,N_11072);
or U12359 (N_12359,N_11403,N_11076);
nand U12360 (N_12360,N_10516,N_11734);
or U12361 (N_12361,N_10755,N_11436);
and U12362 (N_12362,N_11034,N_10786);
xnor U12363 (N_12363,N_10955,N_11230);
nor U12364 (N_12364,N_11448,N_11883);
or U12365 (N_12365,N_10708,N_10807);
and U12366 (N_12366,N_11783,N_10762);
or U12367 (N_12367,N_11172,N_10605);
and U12368 (N_12368,N_10496,N_11547);
or U12369 (N_12369,N_10346,N_11959);
nand U12370 (N_12370,N_11402,N_11126);
or U12371 (N_12371,N_11280,N_10238);
and U12372 (N_12372,N_10500,N_11577);
nand U12373 (N_12373,N_10699,N_11583);
nor U12374 (N_12374,N_10592,N_11199);
or U12375 (N_12375,N_11161,N_10245);
xor U12376 (N_12376,N_10928,N_11347);
and U12377 (N_12377,N_10896,N_11283);
or U12378 (N_12378,N_10289,N_10942);
and U12379 (N_12379,N_11629,N_11059);
nand U12380 (N_12380,N_10436,N_10247);
nand U12381 (N_12381,N_10835,N_11270);
and U12382 (N_12382,N_10417,N_11568);
nand U12383 (N_12383,N_11965,N_10772);
nand U12384 (N_12384,N_11922,N_11481);
nand U12385 (N_12385,N_10106,N_10349);
nor U12386 (N_12386,N_10549,N_10094);
or U12387 (N_12387,N_11320,N_11146);
xor U12388 (N_12388,N_11091,N_11773);
and U12389 (N_12389,N_11987,N_10335);
xor U12390 (N_12390,N_11509,N_10613);
or U12391 (N_12391,N_11561,N_10189);
and U12392 (N_12392,N_10444,N_11937);
and U12393 (N_12393,N_10310,N_11168);
or U12394 (N_12394,N_10638,N_11826);
nand U12395 (N_12395,N_11604,N_11695);
and U12396 (N_12396,N_10543,N_10055);
and U12397 (N_12397,N_11614,N_11616);
nor U12398 (N_12398,N_10956,N_10825);
xor U12399 (N_12399,N_11878,N_10306);
and U12400 (N_12400,N_11316,N_10179);
and U12401 (N_12401,N_10881,N_11388);
nand U12402 (N_12402,N_10152,N_11915);
nand U12403 (N_12403,N_11917,N_10491);
xor U12404 (N_12404,N_10650,N_11255);
and U12405 (N_12405,N_10194,N_10474);
or U12406 (N_12406,N_11214,N_11257);
and U12407 (N_12407,N_10606,N_10387);
and U12408 (N_12408,N_10490,N_10164);
nor U12409 (N_12409,N_10950,N_10261);
nand U12410 (N_12410,N_10885,N_10285);
xor U12411 (N_12411,N_11798,N_11589);
xnor U12412 (N_12412,N_11587,N_11710);
xnor U12413 (N_12413,N_10508,N_11940);
nor U12414 (N_12414,N_10931,N_10286);
or U12415 (N_12415,N_10256,N_10787);
and U12416 (N_12416,N_11467,N_11990);
or U12417 (N_12417,N_11846,N_10017);
and U12418 (N_12418,N_10502,N_10141);
nor U12419 (N_12419,N_10943,N_10646);
or U12420 (N_12420,N_10205,N_10912);
nor U12421 (N_12421,N_11893,N_11543);
nand U12422 (N_12422,N_11781,N_11224);
nor U12423 (N_12423,N_10333,N_10735);
and U12424 (N_12424,N_10649,N_11331);
and U12425 (N_12425,N_11588,N_10204);
xnor U12426 (N_12426,N_10405,N_10591);
or U12427 (N_12427,N_10122,N_11209);
xor U12428 (N_12428,N_11097,N_11670);
nand U12429 (N_12429,N_10859,N_10937);
or U12430 (N_12430,N_11279,N_10160);
and U12431 (N_12431,N_11282,N_10246);
nand U12432 (N_12432,N_11635,N_11017);
nand U12433 (N_12433,N_11698,N_11322);
nand U12434 (N_12434,N_11318,N_11603);
and U12435 (N_12435,N_11941,N_11638);
nand U12436 (N_12436,N_10767,N_10674);
nor U12437 (N_12437,N_10668,N_11370);
nand U12438 (N_12438,N_11737,N_11233);
xor U12439 (N_12439,N_10842,N_11016);
nor U12440 (N_12440,N_11472,N_11399);
nand U12441 (N_12441,N_10267,N_11768);
and U12442 (N_12442,N_11775,N_11828);
or U12443 (N_12443,N_10853,N_10415);
and U12444 (N_12444,N_11903,N_11238);
nor U12445 (N_12445,N_10154,N_10781);
or U12446 (N_12446,N_10300,N_11983);
nand U12447 (N_12447,N_11311,N_11145);
and U12448 (N_12448,N_11809,N_10157);
nor U12449 (N_12449,N_10351,N_10276);
nor U12450 (N_12450,N_11165,N_10398);
nand U12451 (N_12451,N_10919,N_11464);
or U12452 (N_12452,N_11553,N_10722);
nor U12453 (N_12453,N_10015,N_10769);
or U12454 (N_12454,N_11524,N_11303);
nor U12455 (N_12455,N_10833,N_10623);
xnor U12456 (N_12456,N_10441,N_11885);
and U12457 (N_12457,N_11376,N_10693);
nor U12458 (N_12458,N_11755,N_11451);
nor U12459 (N_12459,N_11332,N_10150);
xnor U12460 (N_12460,N_10982,N_10758);
nor U12461 (N_12461,N_11380,N_10635);
or U12462 (N_12462,N_11954,N_11496);
or U12463 (N_12463,N_11455,N_11183);
and U12464 (N_12464,N_10236,N_10275);
nand U12465 (N_12465,N_11202,N_10282);
and U12466 (N_12466,N_10337,N_11205);
nand U12467 (N_12467,N_10301,N_11134);
xnor U12468 (N_12468,N_11799,N_11867);
nand U12469 (N_12469,N_11188,N_11037);
nor U12470 (N_12470,N_10065,N_10235);
and U12471 (N_12471,N_10904,N_10607);
nand U12472 (N_12472,N_11708,N_10661);
and U12473 (N_12473,N_10384,N_11782);
nor U12474 (N_12474,N_10076,N_11406);
xnor U12475 (N_12475,N_11019,N_11929);
nor U12476 (N_12476,N_10099,N_11888);
xor U12477 (N_12477,N_11836,N_11117);
and U12478 (N_12478,N_11726,N_10169);
nand U12479 (N_12479,N_10124,N_10809);
or U12480 (N_12480,N_11101,N_10910);
xnor U12481 (N_12481,N_10171,N_10273);
nor U12482 (N_12482,N_11313,N_10759);
and U12483 (N_12483,N_10797,N_10535);
nor U12484 (N_12484,N_10892,N_11010);
nand U12485 (N_12485,N_11259,N_11786);
or U12486 (N_12486,N_11361,N_10332);
nor U12487 (N_12487,N_10504,N_11778);
or U12488 (N_12488,N_11838,N_10922);
xor U12489 (N_12489,N_11136,N_10132);
and U12490 (N_12490,N_10598,N_11152);
nor U12491 (N_12491,N_11906,N_10480);
xnor U12492 (N_12492,N_11943,N_11606);
nor U12493 (N_12493,N_10430,N_10341);
nand U12494 (N_12494,N_10924,N_10801);
or U12495 (N_12495,N_11434,N_11717);
nor U12496 (N_12496,N_10378,N_10785);
and U12497 (N_12497,N_10000,N_10214);
nand U12498 (N_12498,N_11919,N_10705);
or U12499 (N_12499,N_11654,N_10990);
or U12500 (N_12500,N_10170,N_11256);
nand U12501 (N_12501,N_10745,N_10703);
xnor U12502 (N_12502,N_11853,N_10309);
or U12503 (N_12503,N_10959,N_11516);
or U12504 (N_12504,N_11338,N_11029);
nand U12505 (N_12505,N_11293,N_11834);
nor U12506 (N_12506,N_10840,N_11009);
and U12507 (N_12507,N_11520,N_10980);
nor U12508 (N_12508,N_10039,N_10371);
nand U12509 (N_12509,N_10902,N_10104);
or U12510 (N_12510,N_11083,N_11180);
nor U12511 (N_12511,N_10752,N_11565);
nand U12512 (N_12512,N_10100,N_10666);
or U12513 (N_12513,N_11774,N_10852);
xor U12514 (N_12514,N_11130,N_11772);
nor U12515 (N_12515,N_11790,N_10459);
nor U12516 (N_12516,N_10726,N_11118);
or U12517 (N_12517,N_10465,N_11132);
or U12518 (N_12518,N_10967,N_10882);
nor U12519 (N_12519,N_10114,N_11557);
nand U12520 (N_12520,N_10550,N_10918);
or U12521 (N_12521,N_11375,N_10538);
nor U12522 (N_12522,N_10174,N_11213);
xnor U12523 (N_12523,N_10895,N_10200);
nor U12524 (N_12524,N_11473,N_10472);
nor U12525 (N_12525,N_11337,N_11223);
or U12526 (N_12526,N_10296,N_10034);
xnor U12527 (N_12527,N_10473,N_10746);
nand U12528 (N_12528,N_10829,N_10530);
nor U12529 (N_12529,N_11821,N_11500);
or U12530 (N_12530,N_11362,N_10148);
or U12531 (N_12531,N_10992,N_10359);
xor U12532 (N_12532,N_11418,N_11442);
nand U12533 (N_12533,N_10090,N_11250);
or U12534 (N_12534,N_10356,N_11551);
xor U12535 (N_12535,N_10900,N_11166);
nor U12536 (N_12536,N_10860,N_10702);
and U12537 (N_12537,N_10370,N_10079);
nand U12538 (N_12538,N_11645,N_10754);
and U12539 (N_12539,N_11275,N_10739);
and U12540 (N_12540,N_11295,N_11142);
nor U12541 (N_12541,N_10264,N_11633);
xnor U12542 (N_12542,N_10681,N_10687);
or U12543 (N_12543,N_10626,N_10783);
and U12544 (N_12544,N_10374,N_11912);
or U12545 (N_12545,N_11088,N_10760);
or U12546 (N_12546,N_11907,N_11263);
nand U12547 (N_12547,N_10886,N_10808);
and U12548 (N_12548,N_10093,N_10440);
and U12549 (N_12549,N_11558,N_10232);
or U12550 (N_12550,N_11429,N_11749);
or U12551 (N_12551,N_11327,N_10432);
nand U12552 (N_12552,N_11078,N_11796);
or U12553 (N_12553,N_11763,N_10060);
and U12554 (N_12554,N_11236,N_10684);
and U12555 (N_12555,N_10344,N_11003);
nand U12556 (N_12556,N_10720,N_10230);
nor U12557 (N_12557,N_11135,N_11728);
nor U12558 (N_12558,N_11042,N_11065);
and U12559 (N_12559,N_11648,N_10328);
nor U12560 (N_12560,N_11022,N_11489);
and U12561 (N_12561,N_11555,N_10013);
xor U12562 (N_12562,N_11855,N_11963);
xnor U12563 (N_12563,N_10213,N_10763);
nand U12564 (N_12564,N_10222,N_10006);
nor U12565 (N_12565,N_11608,N_10541);
xor U12566 (N_12566,N_10501,N_10806);
nor U12567 (N_12567,N_10622,N_11969);
nor U12568 (N_12568,N_11823,N_10468);
nand U12569 (N_12569,N_11122,N_10455);
xor U12570 (N_12570,N_10713,N_10053);
xnor U12571 (N_12571,N_11818,N_10905);
nand U12572 (N_12572,N_11780,N_11971);
or U12573 (N_12573,N_10977,N_10268);
and U12574 (N_12574,N_10050,N_11339);
xnor U12575 (N_12575,N_11047,N_11925);
and U12576 (N_12576,N_11049,N_10529);
xnor U12577 (N_12577,N_10828,N_11087);
xor U12578 (N_12578,N_11757,N_10482);
xor U12579 (N_12579,N_10548,N_10048);
xor U12580 (N_12580,N_11719,N_10339);
nand U12581 (N_12581,N_11739,N_10091);
and U12582 (N_12582,N_10458,N_10717);
nand U12583 (N_12583,N_10625,N_11240);
or U12584 (N_12584,N_11383,N_10721);
xor U12585 (N_12585,N_11767,N_11408);
nand U12586 (N_12586,N_11765,N_10527);
or U12587 (N_12587,N_11119,N_11924);
nand U12588 (N_12588,N_11420,N_11956);
or U12589 (N_12589,N_11193,N_10644);
nand U12590 (N_12590,N_11409,N_11452);
xnor U12591 (N_12591,N_10601,N_11484);
or U12592 (N_12592,N_11615,N_11560);
xnor U12593 (N_12593,N_11326,N_10162);
and U12594 (N_12594,N_11675,N_10046);
or U12595 (N_12595,N_10450,N_10003);
xor U12596 (N_12596,N_10198,N_11567);
xor U12597 (N_12597,N_11074,N_11391);
nand U12598 (N_12598,N_10753,N_10195);
xor U12599 (N_12599,N_11540,N_11222);
nor U12600 (N_12600,N_10966,N_10211);
or U12601 (N_12601,N_11852,N_10151);
nand U12602 (N_12602,N_10539,N_11324);
and U12603 (N_12603,N_11221,N_11312);
xnor U12604 (N_12604,N_10498,N_11822);
xnor U12605 (N_12605,N_10159,N_10738);
and U12606 (N_12606,N_11328,N_11729);
xor U12607 (N_12607,N_10112,N_10976);
nand U12608 (N_12608,N_10066,N_11672);
nor U12609 (N_12609,N_11333,N_10437);
and U12610 (N_12610,N_11753,N_11028);
nand U12611 (N_12611,N_11877,N_11972);
nor U12612 (N_12612,N_11860,N_11203);
xor U12613 (N_12613,N_10862,N_10503);
and U12614 (N_12614,N_10407,N_11627);
nand U12615 (N_12615,N_10265,N_10153);
nor U12616 (N_12616,N_11886,N_10402);
nor U12617 (N_12617,N_11173,N_10847);
xor U12618 (N_12618,N_11502,N_10149);
nand U12619 (N_12619,N_11686,N_10989);
and U12620 (N_12620,N_10952,N_10009);
or U12621 (N_12621,N_11539,N_10675);
and U12622 (N_12622,N_10486,N_11094);
and U12623 (N_12623,N_11841,N_11506);
nand U12624 (N_12624,N_10062,N_11461);
nor U12625 (N_12625,N_10897,N_11666);
and U12626 (N_12626,N_10621,N_10838);
nand U12627 (N_12627,N_11181,N_11352);
nand U12628 (N_12628,N_10743,N_10423);
nand U12629 (N_12629,N_11793,N_11641);
nor U12630 (N_12630,N_10224,N_11610);
and U12631 (N_12631,N_11895,N_11738);
nand U12632 (N_12632,N_11012,N_10116);
nor U12633 (N_12633,N_10445,N_10876);
xor U12634 (N_12634,N_11462,N_10706);
nand U12635 (N_12635,N_11660,N_10994);
nand U12636 (N_12636,N_11678,N_11770);
xnor U12637 (N_12637,N_11482,N_10047);
or U12638 (N_12638,N_10442,N_10113);
nand U12639 (N_12639,N_11952,N_11157);
nor U12640 (N_12640,N_11288,N_11994);
xor U12641 (N_12641,N_10193,N_11050);
and U12642 (N_12642,N_10075,N_11563);
nand U12643 (N_12643,N_11752,N_10018);
or U12644 (N_12644,N_11302,N_10263);
xnor U12645 (N_12645,N_11185,N_11227);
and U12646 (N_12646,N_10685,N_11232);
nand U12647 (N_12647,N_10227,N_11991);
nand U12648 (N_12648,N_10741,N_11056);
or U12649 (N_12649,N_11526,N_10562);
and U12650 (N_12650,N_10867,N_10056);
nand U12651 (N_12651,N_11289,N_10740);
nand U12652 (N_12652,N_11881,N_10875);
or U12653 (N_12653,N_11532,N_10969);
nor U12654 (N_12654,N_10487,N_10827);
xor U12655 (N_12655,N_10817,N_10732);
nor U12656 (N_12656,N_10719,N_11623);
or U12657 (N_12657,N_10353,N_11412);
and U12658 (N_12658,N_10907,N_10682);
and U12659 (N_12659,N_11294,N_10184);
or U12660 (N_12660,N_11845,N_11195);
or U12661 (N_12661,N_10610,N_11559);
nor U12662 (N_12662,N_11541,N_10012);
or U12663 (N_12663,N_11667,N_11628);
and U12664 (N_12664,N_11141,N_11802);
xnor U12665 (N_12665,N_11960,N_11084);
nor U12666 (N_12666,N_11384,N_11369);
or U12667 (N_12667,N_11733,N_10834);
and U12668 (N_12668,N_10098,N_10545);
nand U12669 (N_12669,N_11674,N_10587);
or U12670 (N_12670,N_10636,N_11873);
and U12671 (N_12671,N_11114,N_11197);
nand U12672 (N_12672,N_10629,N_10155);
nand U12673 (N_12673,N_10511,N_10903);
xnor U12674 (N_12674,N_11398,N_11979);
nand U12675 (N_12675,N_10658,N_11215);
nor U12676 (N_12676,N_11175,N_10642);
and U12677 (N_12677,N_10338,N_11570);
nor U12678 (N_12678,N_10036,N_10202);
and U12679 (N_12679,N_11620,N_11446);
and U12680 (N_12680,N_11341,N_11154);
xor U12681 (N_12681,N_10672,N_11371);
and U12682 (N_12682,N_11513,N_11368);
nor U12683 (N_12683,N_10299,N_11671);
nand U12684 (N_12684,N_11655,N_10147);
or U12685 (N_12685,N_11291,N_10608);
and U12686 (N_12686,N_10095,N_11847);
nor U12687 (N_12687,N_11365,N_11835);
nor U12688 (N_12688,N_10008,N_10791);
and U12689 (N_12689,N_11918,N_10462);
nor U12690 (N_12690,N_11908,N_11308);
nor U12691 (N_12691,N_10780,N_11814);
xor U12692 (N_12692,N_11914,N_11523);
nand U12693 (N_12693,N_11556,N_11276);
nand U12694 (N_12694,N_10991,N_10586);
nor U12695 (N_12695,N_10711,N_10313);
xnor U12696 (N_12696,N_10010,N_10254);
nand U12697 (N_12697,N_10841,N_11725);
nor U12698 (N_12698,N_11815,N_11664);
nor U12699 (N_12699,N_10172,N_11438);
xor U12700 (N_12700,N_10737,N_10183);
nand U12701 (N_12701,N_11762,N_11191);
and U12702 (N_12702,N_11287,N_11691);
or U12703 (N_12703,N_11159,N_10185);
nand U12704 (N_12704,N_11911,N_11913);
or U12705 (N_12705,N_10870,N_11400);
and U12706 (N_12706,N_11787,N_11286);
or U12707 (N_12707,N_10391,N_11681);
or U12708 (N_12708,N_10866,N_10166);
nand U12709 (N_12709,N_11747,N_11607);
nand U12710 (N_12710,N_11392,N_11599);
nand U12711 (N_12711,N_11748,N_10996);
and U12712 (N_12712,N_10271,N_11977);
and U12713 (N_12713,N_11761,N_10226);
xnor U12714 (N_12714,N_11110,N_10707);
nor U12715 (N_12715,N_10025,N_10914);
nand U12716 (N_12716,N_11004,N_10385);
xnor U12717 (N_12717,N_10074,N_11727);
xor U12718 (N_12718,N_10602,N_10878);
xor U12719 (N_12719,N_11208,N_10253);
or U12720 (N_12720,N_10565,N_11512);
and U12721 (N_12721,N_11309,N_10637);
or U12722 (N_12722,N_11073,N_11812);
and U12723 (N_12723,N_10690,N_10953);
nand U12724 (N_12724,N_10408,N_11478);
or U12725 (N_12725,N_11582,N_11475);
xnor U12726 (N_12726,N_10660,N_10026);
or U12727 (N_12727,N_11414,N_10612);
or U12728 (N_12728,N_11831,N_10073);
nor U12729 (N_12729,N_11550,N_11196);
nand U12730 (N_12730,N_11673,N_10049);
or U12731 (N_12731,N_11508,N_11466);
nand U12732 (N_12732,N_10935,N_11576);
nor U12733 (N_12733,N_10394,N_10540);
or U12734 (N_12734,N_10929,N_11228);
or U12735 (N_12735,N_10005,N_11298);
or U12736 (N_12736,N_10930,N_10766);
and U12737 (N_12737,N_10435,N_10665);
xor U12738 (N_12738,N_11080,N_10143);
xnor U12739 (N_12739,N_11718,N_11124);
xor U12740 (N_12740,N_11035,N_11999);
xnor U12741 (N_12741,N_11483,N_10884);
nor U12742 (N_12742,N_11779,N_10279);
nand U12743 (N_12743,N_10993,N_10083);
and U12744 (N_12744,N_11086,N_10804);
nand U12745 (N_12745,N_11103,N_11225);
xnor U12746 (N_12746,N_10461,N_11031);
and U12747 (N_12747,N_11457,N_10186);
xnor U12748 (N_12748,N_10995,N_11510);
or U12749 (N_12749,N_10639,N_10471);
nor U12750 (N_12750,N_10901,N_10575);
nor U12751 (N_12751,N_11427,N_10067);
and U12752 (N_12752,N_10242,N_10372);
nand U12753 (N_12753,N_11957,N_11866);
and U12754 (N_12754,N_11580,N_11068);
and U12755 (N_12755,N_10443,N_10698);
nand U12756 (N_12756,N_10512,N_11515);
or U12757 (N_12757,N_11373,N_11497);
xor U12758 (N_12758,N_11001,N_11307);
nand U12759 (N_12759,N_10709,N_10489);
nor U12760 (N_12760,N_10107,N_10168);
nor U12761 (N_12761,N_10891,N_10716);
xnor U12762 (N_12762,N_11189,N_11844);
nand U12763 (N_12763,N_10470,N_10485);
or U12764 (N_12764,N_10042,N_11970);
and U12765 (N_12765,N_10020,N_11367);
and U12766 (N_12766,N_10182,N_11636);
nor U12767 (N_12767,N_11820,N_10816);
xor U12768 (N_12768,N_10392,N_10520);
or U12769 (N_12769,N_10686,N_11647);
and U12770 (N_12770,N_11639,N_11996);
nor U12771 (N_12771,N_11246,N_11096);
or U12772 (N_12772,N_11788,N_11447);
nand U12773 (N_12773,N_11184,N_10021);
or U12774 (N_12774,N_10420,N_11121);
or U12775 (N_12775,N_10409,N_10761);
nand U12776 (N_12776,N_10428,N_10101);
nand U12777 (N_12777,N_11921,N_10864);
nor U12778 (N_12778,N_11192,N_11887);
and U12779 (N_12779,N_11656,N_11066);
nand U12780 (N_12780,N_10318,N_10308);
nand U12781 (N_12781,N_10555,N_11120);
xor U12782 (N_12782,N_11843,N_10712);
or U12783 (N_12783,N_10103,N_11043);
nand U12784 (N_12784,N_10559,N_10577);
xnor U12785 (N_12785,N_10814,N_10475);
nor U12786 (N_12786,N_11439,N_10640);
nor U12787 (N_12787,N_10088,N_10469);
xnor U12788 (N_12788,N_11784,N_11771);
nand U12789 (N_12789,N_11958,N_11055);
nor U12790 (N_12790,N_11544,N_11138);
nor U12791 (N_12791,N_11243,N_10016);
xor U12792 (N_12792,N_11849,N_10258);
nor U12793 (N_12793,N_10961,N_11730);
nor U12794 (N_12794,N_10063,N_10004);
nand U12795 (N_12795,N_11542,N_11795);
nor U12796 (N_12796,N_10865,N_10140);
xnor U12797 (N_12797,N_11314,N_10700);
and U12798 (N_12798,N_10311,N_11330);
and U12799 (N_12799,N_11274,N_11479);
xor U12800 (N_12800,N_10648,N_11002);
and U12801 (N_12801,N_11754,N_10974);
xor U12802 (N_12802,N_10360,N_10794);
nor U12803 (N_12803,N_11235,N_11393);
or U12804 (N_12804,N_11984,N_10782);
nor U12805 (N_12805,N_10528,N_10813);
nor U12806 (N_12806,N_10954,N_10948);
xor U12807 (N_12807,N_10163,N_11258);
and U12808 (N_12808,N_11789,N_11842);
nand U12809 (N_12809,N_10863,N_11564);
xor U12810 (N_12810,N_11596,N_10514);
and U12811 (N_12811,N_11968,N_11503);
or U12812 (N_12812,N_10051,N_10326);
nor U12813 (N_12813,N_10748,N_10316);
and U12814 (N_12814,N_10393,N_11090);
and U12815 (N_12815,N_11694,N_10108);
nand U12816 (N_12816,N_10251,N_10290);
nand U12817 (N_12817,N_10175,N_11397);
nor U12818 (N_12818,N_10572,N_10645);
nand U12819 (N_12819,N_10281,N_10581);
or U12820 (N_12820,N_10887,N_10396);
nand U12821 (N_12821,N_11304,N_11622);
xnor U12822 (N_12822,N_11261,N_11133);
nor U12823 (N_12823,N_10342,N_11386);
and U12824 (N_12824,N_11998,N_10916);
nand U12825 (N_12825,N_10725,N_10615);
nor U12826 (N_12826,N_10542,N_11000);
xnor U12827 (N_12827,N_11252,N_10118);
nand U12828 (N_12828,N_11245,N_11519);
nor U12829 (N_12829,N_10357,N_11679);
and U12830 (N_12830,N_10569,N_11537);
and U12831 (N_12831,N_10652,N_11060);
nor U12832 (N_12832,N_10906,N_11816);
nor U12833 (N_12833,N_10773,N_11743);
nand U12834 (N_12834,N_11081,N_10894);
and U12835 (N_12835,N_10551,N_11179);
xnor U12836 (N_12836,N_10653,N_10523);
nand U12837 (N_12837,N_11548,N_10960);
nor U12838 (N_12838,N_10037,N_10544);
and U12839 (N_12839,N_11992,N_10774);
nor U12840 (N_12840,N_10040,N_10964);
or U12841 (N_12841,N_11336,N_11945);
nor U12842 (N_12842,N_11106,N_11160);
xor U12843 (N_12843,N_11706,N_10136);
nor U12844 (N_12844,N_10851,N_10715);
and U12845 (N_12845,N_11459,N_11343);
nand U12846 (N_12846,N_11150,N_11711);
nand U12847 (N_12847,N_10364,N_10228);
or U12848 (N_12848,N_10552,N_10877);
nand U12849 (N_12849,N_10826,N_10336);
nand U12850 (N_12850,N_10571,N_11187);
nand U12851 (N_12851,N_10683,N_10144);
xnor U12852 (N_12852,N_11934,N_11722);
xor U12853 (N_12853,N_11444,N_10958);
or U12854 (N_12854,N_11297,N_10557);
or U12855 (N_12855,N_11260,N_11653);
and U12856 (N_12856,N_10043,N_11174);
nand U12857 (N_12857,N_11374,N_10237);
or U12858 (N_12858,N_11018,N_10962);
xor U12859 (N_12859,N_11206,N_11904);
nand U12860 (N_12860,N_10463,N_10438);
and U12861 (N_12861,N_10262,N_10284);
nor U12862 (N_12862,N_11108,N_10789);
nand U12863 (N_12863,N_10777,N_11200);
nor U12864 (N_12864,N_11964,N_10909);
xnor U12865 (N_12865,N_11177,N_10161);
xnor U12866 (N_12866,N_11476,N_10307);
or U12867 (N_12867,N_11360,N_10733);
xnor U12868 (N_12868,N_11163,N_10822);
nand U12869 (N_12869,N_11766,N_11901);
and U12870 (N_12870,N_11756,N_11859);
xnor U12871 (N_12871,N_11306,N_11470);
nor U12872 (N_12872,N_11450,N_10616);
nand U12873 (N_12873,N_10963,N_10483);
xor U12874 (N_12874,N_11707,N_10446);
nor U12875 (N_12875,N_10382,N_11792);
nor U12876 (N_12876,N_10479,N_10007);
and U12877 (N_12877,N_11750,N_11839);
and U12878 (N_12878,N_11323,N_11379);
nand U12879 (N_12879,N_10526,N_11804);
or U12880 (N_12880,N_10628,N_10532);
xor U12881 (N_12881,N_11806,N_10041);
and U12882 (N_12882,N_10971,N_11942);
nand U12883 (N_12883,N_11249,N_11549);
nor U12884 (N_12884,N_11491,N_11021);
and U12885 (N_12885,N_10788,N_11463);
nand U12886 (N_12886,N_10634,N_10553);
and U12887 (N_12887,N_11299,N_10676);
nand U12888 (N_12888,N_11995,N_11453);
nand U12889 (N_12889,N_11417,N_11315);
nand U12890 (N_12890,N_10941,N_10033);
xnor U12891 (N_12891,N_11988,N_10568);
nand U12892 (N_12892,N_11006,N_10946);
or U12893 (N_12893,N_11601,N_10325);
and U12894 (N_12894,N_11284,N_10390);
nor U12895 (N_12895,N_11201,N_11593);
xor U12896 (N_12896,N_11889,N_11265);
xor U12897 (N_12897,N_11413,N_11811);
nand U12898 (N_12898,N_10303,N_11829);
nand U12899 (N_12899,N_10028,N_11985);
xnor U12900 (N_12900,N_10368,N_11702);
xnor U12901 (N_12901,N_10082,N_10249);
nand U12902 (N_12902,N_11013,N_11948);
xnor U12903 (N_12903,N_11030,N_10188);
xnor U12904 (N_12904,N_10192,N_11947);
xnor U12905 (N_12905,N_11061,N_11923);
or U12906 (N_12906,N_11156,N_10810);
nor U12907 (N_12907,N_10293,N_10002);
nand U12908 (N_12908,N_10839,N_11389);
and U12909 (N_12909,N_11102,N_10377);
nor U12910 (N_12910,N_10045,N_11372);
xnor U12911 (N_12911,N_11054,N_11105);
xnor U12912 (N_12912,N_10795,N_11676);
and U12913 (N_12913,N_11662,N_10534);
and U12914 (N_12914,N_11807,N_10252);
or U12915 (N_12915,N_10911,N_10975);
or U12916 (N_12916,N_10899,N_11217);
nand U12917 (N_12917,N_11533,N_10330);
or U12918 (N_12918,N_11356,N_11993);
or U12919 (N_12919,N_10416,N_11458);
or U12920 (N_12920,N_10927,N_11731);
xor U12921 (N_12921,N_11069,N_11485);
nor U12922 (N_12922,N_10072,N_10556);
xor U12923 (N_12923,N_11226,N_10848);
xnor U12924 (N_12924,N_11107,N_11366);
or U12925 (N_12925,N_11231,N_11851);
nand U12926 (N_12926,N_11182,N_11498);
nor U12927 (N_12927,N_10493,N_11709);
or U12928 (N_12928,N_11571,N_10105);
or U12929 (N_12929,N_11501,N_10764);
or U12930 (N_12930,N_10803,N_11894);
nand U12931 (N_12931,N_10778,N_10421);
and U12932 (N_12932,N_11251,N_11053);
nand U12933 (N_12933,N_10888,N_11522);
xnor U12934 (N_12934,N_10321,N_11048);
nand U12935 (N_12935,N_11871,N_11832);
nor U12936 (N_12936,N_10431,N_11421);
nor U12937 (N_12937,N_11186,N_11310);
or U12938 (N_12938,N_10779,N_11317);
nor U12939 (N_12939,N_11652,N_11566);
and U12940 (N_12940,N_11932,N_11863);
nand U12941 (N_12941,N_10983,N_10494);
or U12942 (N_12942,N_11651,N_11953);
or U12943 (N_12943,N_10536,N_10156);
and U12944 (N_12944,N_10915,N_11441);
and U12945 (N_12945,N_10988,N_11129);
nor U12946 (N_12946,N_10978,N_10871);
nand U12947 (N_12947,N_10836,N_11354);
or U12948 (N_12948,N_11874,N_10656);
or U12949 (N_12949,N_10965,N_11071);
nand U12950 (N_12950,N_10936,N_10673);
nand U12951 (N_12951,N_10932,N_11528);
or U12952 (N_12952,N_10197,N_10604);
and U12953 (N_12953,N_11045,N_11825);
xor U12954 (N_12954,N_10134,N_11092);
xnor U12955 (N_12955,N_10582,N_10898);
or U12956 (N_12956,N_10269,N_11521);
and U12957 (N_12957,N_10689,N_10537);
xor U12958 (N_12958,N_10949,N_10751);
or U12959 (N_12959,N_10655,N_10111);
nor U12960 (N_12960,N_10522,N_10130);
and U12961 (N_12961,N_10355,N_10180);
nor U12962 (N_12962,N_11267,N_10873);
or U12963 (N_12963,N_10086,N_10054);
nor U12964 (N_12964,N_10696,N_10343);
or U12965 (N_12965,N_10654,N_10223);
or U12966 (N_12966,N_10609,N_11975);
and U12967 (N_12967,N_11978,N_11740);
nand U12968 (N_12968,N_11856,N_10880);
nand U12969 (N_12969,N_11058,N_11827);
nand U12970 (N_12970,N_11892,N_10492);
nor U12971 (N_12971,N_10855,N_11764);
nand U12972 (N_12972,N_11700,N_11890);
nand U12973 (N_12973,N_11644,N_11861);
nor U12974 (N_12974,N_11511,N_10229);
nand U12975 (N_12975,N_11211,N_11405);
or U12976 (N_12976,N_10987,N_10692);
and U12977 (N_12977,N_11248,N_10412);
nand U12978 (N_12978,N_10657,N_10395);
xor U12979 (N_12979,N_10453,N_10133);
or U12980 (N_12980,N_10749,N_10768);
xor U12981 (N_12981,N_11723,N_10633);
nand U12982 (N_12982,N_10317,N_11407);
nor U12983 (N_12983,N_11426,N_11554);
nand U12984 (N_12984,N_10951,N_10731);
nand U12985 (N_12985,N_11428,N_10679);
nand U12986 (N_12986,N_10662,N_11982);
nand U12987 (N_12987,N_11247,N_11381);
and U12988 (N_12988,N_10210,N_10481);
nand U12989 (N_12989,N_11272,N_11797);
xor U12990 (N_12990,N_11534,N_11605);
and U12991 (N_12991,N_11704,N_10345);
xor U12992 (N_12992,N_10593,N_11864);
nor U12993 (N_12993,N_10201,N_11079);
nand U12994 (N_12994,N_10081,N_10973);
and U12995 (N_12995,N_10024,N_11572);
or U12996 (N_12996,N_11865,N_11363);
and U12997 (N_12997,N_10070,N_10121);
or U12998 (N_12998,N_10590,N_11697);
xnor U12999 (N_12999,N_10297,N_11830);
nor U13000 (N_13000,N_11196,N_10709);
nor U13001 (N_13001,N_10418,N_11985);
nand U13002 (N_13002,N_10389,N_10062);
and U13003 (N_13003,N_10624,N_10164);
or U13004 (N_13004,N_10304,N_10506);
or U13005 (N_13005,N_11591,N_11974);
or U13006 (N_13006,N_10698,N_11588);
xnor U13007 (N_13007,N_10503,N_11464);
nand U13008 (N_13008,N_11687,N_11645);
nor U13009 (N_13009,N_11744,N_10371);
nand U13010 (N_13010,N_10996,N_11577);
nand U13011 (N_13011,N_11587,N_10735);
nor U13012 (N_13012,N_10348,N_10655);
and U13013 (N_13013,N_11592,N_10542);
nor U13014 (N_13014,N_10599,N_10347);
nand U13015 (N_13015,N_10072,N_11791);
or U13016 (N_13016,N_11038,N_10780);
and U13017 (N_13017,N_11545,N_10167);
nor U13018 (N_13018,N_10286,N_10199);
or U13019 (N_13019,N_10878,N_11360);
xor U13020 (N_13020,N_10461,N_10789);
nand U13021 (N_13021,N_11667,N_10873);
and U13022 (N_13022,N_11022,N_11886);
xnor U13023 (N_13023,N_11358,N_11619);
and U13024 (N_13024,N_10257,N_11133);
nor U13025 (N_13025,N_10703,N_11569);
and U13026 (N_13026,N_10378,N_10456);
nor U13027 (N_13027,N_11721,N_10388);
or U13028 (N_13028,N_10731,N_11961);
nand U13029 (N_13029,N_11962,N_11892);
or U13030 (N_13030,N_11913,N_11297);
nand U13031 (N_13031,N_10753,N_11812);
nand U13032 (N_13032,N_11171,N_10348);
or U13033 (N_13033,N_11999,N_10164);
and U13034 (N_13034,N_11885,N_10845);
or U13035 (N_13035,N_11567,N_10791);
nor U13036 (N_13036,N_10479,N_11975);
nand U13037 (N_13037,N_10039,N_10642);
or U13038 (N_13038,N_10745,N_11575);
nand U13039 (N_13039,N_11026,N_10220);
nor U13040 (N_13040,N_10486,N_11277);
or U13041 (N_13041,N_11964,N_10099);
or U13042 (N_13042,N_10193,N_10484);
and U13043 (N_13043,N_11948,N_10548);
nor U13044 (N_13044,N_11937,N_10332);
xnor U13045 (N_13045,N_11365,N_11014);
or U13046 (N_13046,N_11617,N_11652);
xnor U13047 (N_13047,N_11770,N_10357);
and U13048 (N_13048,N_11006,N_11700);
xor U13049 (N_13049,N_11590,N_11360);
nor U13050 (N_13050,N_11211,N_10152);
xor U13051 (N_13051,N_11541,N_11949);
nor U13052 (N_13052,N_10328,N_10512);
nor U13053 (N_13053,N_11188,N_11819);
nand U13054 (N_13054,N_10775,N_10976);
xor U13055 (N_13055,N_11108,N_11552);
nor U13056 (N_13056,N_11897,N_11476);
nor U13057 (N_13057,N_11694,N_11735);
nand U13058 (N_13058,N_10014,N_10757);
and U13059 (N_13059,N_10258,N_10882);
nor U13060 (N_13060,N_10180,N_11718);
or U13061 (N_13061,N_11004,N_11373);
nand U13062 (N_13062,N_10768,N_10138);
xnor U13063 (N_13063,N_10199,N_10476);
or U13064 (N_13064,N_11668,N_10628);
nor U13065 (N_13065,N_10564,N_11964);
xnor U13066 (N_13066,N_11135,N_11667);
nand U13067 (N_13067,N_11635,N_11563);
xnor U13068 (N_13068,N_10401,N_11441);
nor U13069 (N_13069,N_11603,N_11534);
xnor U13070 (N_13070,N_11952,N_11882);
nand U13071 (N_13071,N_10338,N_11217);
and U13072 (N_13072,N_10520,N_11846);
nor U13073 (N_13073,N_11354,N_11915);
or U13074 (N_13074,N_10944,N_10734);
nand U13075 (N_13075,N_11298,N_10152);
or U13076 (N_13076,N_10779,N_11880);
nor U13077 (N_13077,N_10606,N_11663);
nor U13078 (N_13078,N_11586,N_11409);
or U13079 (N_13079,N_11571,N_10384);
xor U13080 (N_13080,N_10193,N_11948);
xor U13081 (N_13081,N_10941,N_11858);
nor U13082 (N_13082,N_10152,N_10081);
nor U13083 (N_13083,N_11608,N_10070);
and U13084 (N_13084,N_10752,N_10811);
xor U13085 (N_13085,N_10530,N_11921);
nand U13086 (N_13086,N_11328,N_11630);
nand U13087 (N_13087,N_10822,N_10290);
xor U13088 (N_13088,N_10082,N_11851);
nand U13089 (N_13089,N_11316,N_10249);
or U13090 (N_13090,N_10822,N_11962);
nor U13091 (N_13091,N_10345,N_10175);
xnor U13092 (N_13092,N_11208,N_10720);
or U13093 (N_13093,N_11689,N_10070);
and U13094 (N_13094,N_10200,N_11226);
and U13095 (N_13095,N_11616,N_11968);
and U13096 (N_13096,N_11521,N_10055);
and U13097 (N_13097,N_10856,N_10296);
nor U13098 (N_13098,N_11628,N_11849);
nor U13099 (N_13099,N_11898,N_10938);
and U13100 (N_13100,N_10011,N_11141);
or U13101 (N_13101,N_10027,N_10899);
and U13102 (N_13102,N_10929,N_11890);
nand U13103 (N_13103,N_10733,N_10402);
or U13104 (N_13104,N_11162,N_11401);
xnor U13105 (N_13105,N_11893,N_11652);
nor U13106 (N_13106,N_10888,N_10452);
nand U13107 (N_13107,N_10290,N_11646);
or U13108 (N_13108,N_11114,N_11036);
xor U13109 (N_13109,N_11857,N_11823);
nor U13110 (N_13110,N_10554,N_11320);
xor U13111 (N_13111,N_10008,N_10297);
nand U13112 (N_13112,N_10787,N_11087);
xnor U13113 (N_13113,N_11175,N_10962);
xnor U13114 (N_13114,N_11397,N_10961);
or U13115 (N_13115,N_10397,N_11598);
and U13116 (N_13116,N_10530,N_11899);
xor U13117 (N_13117,N_11600,N_11425);
and U13118 (N_13118,N_10308,N_11431);
and U13119 (N_13119,N_10010,N_11174);
nor U13120 (N_13120,N_11549,N_11460);
xnor U13121 (N_13121,N_11388,N_11652);
and U13122 (N_13122,N_11080,N_10262);
or U13123 (N_13123,N_10431,N_11870);
and U13124 (N_13124,N_11521,N_11994);
nand U13125 (N_13125,N_10414,N_10493);
xor U13126 (N_13126,N_11264,N_10617);
nor U13127 (N_13127,N_11871,N_11314);
xnor U13128 (N_13128,N_11882,N_11997);
or U13129 (N_13129,N_11082,N_10240);
nand U13130 (N_13130,N_10834,N_10220);
or U13131 (N_13131,N_10773,N_10083);
and U13132 (N_13132,N_10934,N_11093);
or U13133 (N_13133,N_10043,N_10383);
nor U13134 (N_13134,N_10189,N_11976);
xor U13135 (N_13135,N_11275,N_11222);
or U13136 (N_13136,N_10230,N_10122);
nand U13137 (N_13137,N_11644,N_11956);
or U13138 (N_13138,N_11234,N_11245);
or U13139 (N_13139,N_10865,N_11737);
nand U13140 (N_13140,N_10491,N_10801);
and U13141 (N_13141,N_11769,N_10142);
and U13142 (N_13142,N_11039,N_11304);
and U13143 (N_13143,N_10493,N_11948);
xor U13144 (N_13144,N_10959,N_10226);
xor U13145 (N_13145,N_10610,N_10408);
and U13146 (N_13146,N_11639,N_10167);
or U13147 (N_13147,N_10705,N_10733);
or U13148 (N_13148,N_11204,N_11167);
xor U13149 (N_13149,N_11722,N_10529);
and U13150 (N_13150,N_11869,N_11582);
or U13151 (N_13151,N_10023,N_11198);
nor U13152 (N_13152,N_10661,N_11767);
nor U13153 (N_13153,N_11997,N_11485);
nand U13154 (N_13154,N_10154,N_10751);
and U13155 (N_13155,N_11300,N_11692);
and U13156 (N_13156,N_11796,N_10098);
xnor U13157 (N_13157,N_10431,N_11566);
nand U13158 (N_13158,N_11068,N_11143);
nor U13159 (N_13159,N_11087,N_11198);
nor U13160 (N_13160,N_10360,N_11733);
nand U13161 (N_13161,N_10162,N_11799);
xnor U13162 (N_13162,N_11375,N_11339);
xor U13163 (N_13163,N_10136,N_11769);
and U13164 (N_13164,N_11407,N_10111);
nand U13165 (N_13165,N_10533,N_11190);
nand U13166 (N_13166,N_10425,N_10231);
nor U13167 (N_13167,N_10328,N_10023);
nand U13168 (N_13168,N_10162,N_11731);
nand U13169 (N_13169,N_10320,N_10777);
nand U13170 (N_13170,N_10340,N_11709);
nand U13171 (N_13171,N_11128,N_10623);
and U13172 (N_13172,N_10412,N_11684);
nand U13173 (N_13173,N_11463,N_11792);
nand U13174 (N_13174,N_11684,N_10860);
xor U13175 (N_13175,N_11062,N_10472);
nor U13176 (N_13176,N_11525,N_10510);
nand U13177 (N_13177,N_11446,N_11281);
and U13178 (N_13178,N_10175,N_11183);
xor U13179 (N_13179,N_11024,N_11017);
nor U13180 (N_13180,N_11173,N_10185);
or U13181 (N_13181,N_10700,N_11853);
xor U13182 (N_13182,N_10287,N_11266);
nor U13183 (N_13183,N_10856,N_11749);
nor U13184 (N_13184,N_10009,N_10222);
xor U13185 (N_13185,N_10507,N_11058);
nor U13186 (N_13186,N_10837,N_10021);
nand U13187 (N_13187,N_11582,N_10766);
and U13188 (N_13188,N_11742,N_11980);
and U13189 (N_13189,N_10967,N_11654);
nor U13190 (N_13190,N_10961,N_10768);
nor U13191 (N_13191,N_10107,N_10817);
or U13192 (N_13192,N_10692,N_10750);
nor U13193 (N_13193,N_11029,N_10595);
xor U13194 (N_13194,N_10128,N_10607);
nor U13195 (N_13195,N_11551,N_11627);
xnor U13196 (N_13196,N_10602,N_10395);
nand U13197 (N_13197,N_10964,N_11241);
and U13198 (N_13198,N_11852,N_10319);
nor U13199 (N_13199,N_10898,N_11498);
xor U13200 (N_13200,N_10048,N_11675);
nand U13201 (N_13201,N_10812,N_11467);
or U13202 (N_13202,N_10644,N_10189);
or U13203 (N_13203,N_10526,N_10572);
nor U13204 (N_13204,N_11606,N_11795);
xor U13205 (N_13205,N_11142,N_11382);
xor U13206 (N_13206,N_11366,N_11651);
nor U13207 (N_13207,N_11139,N_10183);
nor U13208 (N_13208,N_10855,N_10152);
nand U13209 (N_13209,N_11000,N_10203);
or U13210 (N_13210,N_10495,N_10087);
nor U13211 (N_13211,N_11071,N_10358);
nor U13212 (N_13212,N_11579,N_10606);
xnor U13213 (N_13213,N_11526,N_11749);
nor U13214 (N_13214,N_11394,N_11006);
and U13215 (N_13215,N_10588,N_10313);
xnor U13216 (N_13216,N_11659,N_10560);
nand U13217 (N_13217,N_11989,N_11853);
nand U13218 (N_13218,N_11307,N_10681);
or U13219 (N_13219,N_11576,N_10098);
nor U13220 (N_13220,N_10840,N_10141);
and U13221 (N_13221,N_10862,N_11417);
nand U13222 (N_13222,N_10019,N_11481);
xor U13223 (N_13223,N_11647,N_11075);
and U13224 (N_13224,N_10839,N_10939);
and U13225 (N_13225,N_10970,N_11448);
xnor U13226 (N_13226,N_10967,N_10585);
or U13227 (N_13227,N_11693,N_11446);
nor U13228 (N_13228,N_11113,N_11017);
or U13229 (N_13229,N_10578,N_11430);
or U13230 (N_13230,N_11594,N_10570);
or U13231 (N_13231,N_10453,N_10730);
nor U13232 (N_13232,N_10553,N_10387);
nor U13233 (N_13233,N_11224,N_11593);
nor U13234 (N_13234,N_10325,N_10643);
or U13235 (N_13235,N_10861,N_10131);
xnor U13236 (N_13236,N_11740,N_11165);
and U13237 (N_13237,N_11035,N_11284);
or U13238 (N_13238,N_10071,N_11040);
and U13239 (N_13239,N_11399,N_11526);
nand U13240 (N_13240,N_10551,N_11036);
and U13241 (N_13241,N_10983,N_11243);
and U13242 (N_13242,N_10088,N_11971);
xnor U13243 (N_13243,N_10324,N_10461);
nand U13244 (N_13244,N_11690,N_10438);
and U13245 (N_13245,N_11221,N_10641);
nand U13246 (N_13246,N_11905,N_11786);
nor U13247 (N_13247,N_10259,N_11128);
xnor U13248 (N_13248,N_10389,N_10668);
nand U13249 (N_13249,N_11951,N_10627);
xnor U13250 (N_13250,N_10032,N_10470);
nor U13251 (N_13251,N_10474,N_10648);
xnor U13252 (N_13252,N_10639,N_10036);
xor U13253 (N_13253,N_11195,N_10809);
or U13254 (N_13254,N_10929,N_10423);
nand U13255 (N_13255,N_10789,N_11636);
or U13256 (N_13256,N_11435,N_10780);
nand U13257 (N_13257,N_10179,N_10481);
or U13258 (N_13258,N_10088,N_11278);
nor U13259 (N_13259,N_11791,N_11069);
nor U13260 (N_13260,N_11822,N_10427);
nor U13261 (N_13261,N_10337,N_10084);
and U13262 (N_13262,N_11825,N_11684);
nor U13263 (N_13263,N_11650,N_11131);
nor U13264 (N_13264,N_11122,N_11522);
or U13265 (N_13265,N_10020,N_11857);
nand U13266 (N_13266,N_10618,N_11171);
or U13267 (N_13267,N_11696,N_10026);
xor U13268 (N_13268,N_11058,N_10446);
nand U13269 (N_13269,N_11937,N_10140);
xor U13270 (N_13270,N_10866,N_11312);
and U13271 (N_13271,N_10892,N_10197);
and U13272 (N_13272,N_11565,N_10526);
nor U13273 (N_13273,N_11805,N_10781);
xor U13274 (N_13274,N_10874,N_10865);
nor U13275 (N_13275,N_11514,N_10838);
or U13276 (N_13276,N_10401,N_10777);
xnor U13277 (N_13277,N_11561,N_10300);
nor U13278 (N_13278,N_10651,N_11409);
and U13279 (N_13279,N_10428,N_10190);
and U13280 (N_13280,N_11193,N_10004);
nand U13281 (N_13281,N_10965,N_11035);
nor U13282 (N_13282,N_11008,N_11850);
nand U13283 (N_13283,N_11508,N_10601);
or U13284 (N_13284,N_11575,N_11979);
and U13285 (N_13285,N_11754,N_11525);
nor U13286 (N_13286,N_11327,N_11094);
and U13287 (N_13287,N_11600,N_10777);
nor U13288 (N_13288,N_11229,N_11974);
xnor U13289 (N_13289,N_11387,N_11124);
nor U13290 (N_13290,N_10276,N_10914);
and U13291 (N_13291,N_11613,N_11292);
and U13292 (N_13292,N_10817,N_11145);
xor U13293 (N_13293,N_11456,N_11283);
and U13294 (N_13294,N_10546,N_10288);
nand U13295 (N_13295,N_11831,N_11445);
nor U13296 (N_13296,N_11420,N_11712);
xnor U13297 (N_13297,N_11866,N_10631);
xnor U13298 (N_13298,N_11278,N_10390);
or U13299 (N_13299,N_10354,N_11524);
or U13300 (N_13300,N_10909,N_10518);
nand U13301 (N_13301,N_10264,N_10922);
and U13302 (N_13302,N_11626,N_10990);
and U13303 (N_13303,N_10431,N_10685);
and U13304 (N_13304,N_10715,N_11408);
xor U13305 (N_13305,N_11960,N_11471);
or U13306 (N_13306,N_10425,N_11280);
xor U13307 (N_13307,N_10820,N_11841);
xnor U13308 (N_13308,N_10425,N_11226);
or U13309 (N_13309,N_11079,N_10679);
xor U13310 (N_13310,N_10736,N_11569);
nand U13311 (N_13311,N_10227,N_11469);
nor U13312 (N_13312,N_11825,N_11654);
and U13313 (N_13313,N_11962,N_10194);
nand U13314 (N_13314,N_10031,N_10515);
nand U13315 (N_13315,N_10812,N_10839);
xor U13316 (N_13316,N_11367,N_11852);
nor U13317 (N_13317,N_11842,N_10887);
nor U13318 (N_13318,N_11268,N_10185);
nor U13319 (N_13319,N_11326,N_10660);
or U13320 (N_13320,N_10752,N_10517);
nor U13321 (N_13321,N_11666,N_11028);
and U13322 (N_13322,N_11002,N_11162);
nor U13323 (N_13323,N_11125,N_11781);
nor U13324 (N_13324,N_11597,N_11936);
xnor U13325 (N_13325,N_11357,N_10356);
or U13326 (N_13326,N_10244,N_11927);
nor U13327 (N_13327,N_11438,N_10014);
nor U13328 (N_13328,N_11297,N_10315);
or U13329 (N_13329,N_10568,N_11404);
nand U13330 (N_13330,N_10173,N_11046);
or U13331 (N_13331,N_10425,N_10760);
and U13332 (N_13332,N_11251,N_11703);
nand U13333 (N_13333,N_10440,N_11986);
xnor U13334 (N_13334,N_10941,N_11494);
xor U13335 (N_13335,N_10228,N_10573);
xor U13336 (N_13336,N_10066,N_10285);
xor U13337 (N_13337,N_11687,N_10559);
and U13338 (N_13338,N_11307,N_11432);
or U13339 (N_13339,N_11750,N_10007);
nor U13340 (N_13340,N_10645,N_11308);
nand U13341 (N_13341,N_10858,N_10008);
xnor U13342 (N_13342,N_11523,N_11260);
nor U13343 (N_13343,N_11687,N_10172);
or U13344 (N_13344,N_11684,N_10311);
nand U13345 (N_13345,N_11886,N_10160);
xor U13346 (N_13346,N_10374,N_10560);
nor U13347 (N_13347,N_11699,N_10023);
xor U13348 (N_13348,N_11034,N_11795);
nand U13349 (N_13349,N_10147,N_10660);
xor U13350 (N_13350,N_10410,N_11263);
xnor U13351 (N_13351,N_11307,N_11460);
and U13352 (N_13352,N_10965,N_11428);
and U13353 (N_13353,N_11851,N_10613);
xnor U13354 (N_13354,N_10119,N_10075);
nor U13355 (N_13355,N_10131,N_10021);
xor U13356 (N_13356,N_10450,N_10805);
xor U13357 (N_13357,N_11315,N_10839);
nand U13358 (N_13358,N_10244,N_10240);
and U13359 (N_13359,N_11336,N_10555);
and U13360 (N_13360,N_11810,N_11688);
nand U13361 (N_13361,N_11874,N_10634);
nand U13362 (N_13362,N_11479,N_10105);
nand U13363 (N_13363,N_11068,N_11764);
nand U13364 (N_13364,N_10822,N_11428);
nand U13365 (N_13365,N_11738,N_10514);
nand U13366 (N_13366,N_10021,N_11609);
xor U13367 (N_13367,N_11364,N_11246);
xnor U13368 (N_13368,N_10537,N_11684);
nand U13369 (N_13369,N_11678,N_11743);
or U13370 (N_13370,N_11812,N_10826);
and U13371 (N_13371,N_11054,N_11228);
nand U13372 (N_13372,N_11825,N_10330);
nand U13373 (N_13373,N_11868,N_10904);
nor U13374 (N_13374,N_10651,N_11752);
nor U13375 (N_13375,N_11775,N_11413);
nor U13376 (N_13376,N_10140,N_10498);
or U13377 (N_13377,N_11126,N_10662);
nand U13378 (N_13378,N_10625,N_10520);
or U13379 (N_13379,N_11179,N_11932);
nor U13380 (N_13380,N_10453,N_11596);
and U13381 (N_13381,N_10533,N_10364);
nand U13382 (N_13382,N_10504,N_10515);
xnor U13383 (N_13383,N_10752,N_10423);
or U13384 (N_13384,N_11429,N_10736);
nand U13385 (N_13385,N_10717,N_11954);
xnor U13386 (N_13386,N_10521,N_10627);
nand U13387 (N_13387,N_10365,N_11856);
and U13388 (N_13388,N_11551,N_11731);
and U13389 (N_13389,N_11737,N_10302);
or U13390 (N_13390,N_11429,N_10856);
and U13391 (N_13391,N_10893,N_10337);
xor U13392 (N_13392,N_11732,N_10470);
nor U13393 (N_13393,N_10189,N_10074);
or U13394 (N_13394,N_10534,N_10731);
and U13395 (N_13395,N_11716,N_10174);
and U13396 (N_13396,N_10080,N_11576);
and U13397 (N_13397,N_10280,N_11490);
nand U13398 (N_13398,N_11617,N_11057);
nor U13399 (N_13399,N_11582,N_11605);
and U13400 (N_13400,N_10181,N_10879);
and U13401 (N_13401,N_10497,N_10244);
xor U13402 (N_13402,N_10839,N_10079);
nor U13403 (N_13403,N_11207,N_10972);
xor U13404 (N_13404,N_11154,N_10993);
and U13405 (N_13405,N_11485,N_11171);
nor U13406 (N_13406,N_10294,N_10802);
nor U13407 (N_13407,N_11946,N_10491);
and U13408 (N_13408,N_11355,N_10898);
nand U13409 (N_13409,N_11708,N_10520);
or U13410 (N_13410,N_10543,N_11875);
and U13411 (N_13411,N_11831,N_11687);
nand U13412 (N_13412,N_11522,N_10253);
nand U13413 (N_13413,N_11137,N_11982);
nor U13414 (N_13414,N_11766,N_10676);
nor U13415 (N_13415,N_10776,N_11511);
xnor U13416 (N_13416,N_11073,N_10375);
or U13417 (N_13417,N_11534,N_10492);
and U13418 (N_13418,N_11988,N_11263);
nand U13419 (N_13419,N_10564,N_10137);
nand U13420 (N_13420,N_10180,N_11131);
xnor U13421 (N_13421,N_11607,N_10476);
or U13422 (N_13422,N_11894,N_10575);
or U13423 (N_13423,N_11308,N_11653);
nor U13424 (N_13424,N_10787,N_11442);
xor U13425 (N_13425,N_10734,N_10977);
or U13426 (N_13426,N_11840,N_10928);
nor U13427 (N_13427,N_11111,N_11647);
nand U13428 (N_13428,N_10642,N_10701);
nand U13429 (N_13429,N_11912,N_11511);
and U13430 (N_13430,N_10946,N_11410);
xnor U13431 (N_13431,N_11884,N_11168);
nor U13432 (N_13432,N_10923,N_11082);
nand U13433 (N_13433,N_10948,N_11709);
and U13434 (N_13434,N_11762,N_11453);
nand U13435 (N_13435,N_10414,N_10060);
xnor U13436 (N_13436,N_10111,N_10184);
nand U13437 (N_13437,N_10110,N_11790);
xnor U13438 (N_13438,N_11711,N_10487);
and U13439 (N_13439,N_11899,N_11020);
nor U13440 (N_13440,N_11560,N_11315);
or U13441 (N_13441,N_10757,N_11650);
nand U13442 (N_13442,N_11622,N_11916);
nand U13443 (N_13443,N_10825,N_11702);
or U13444 (N_13444,N_11408,N_11464);
or U13445 (N_13445,N_11572,N_11592);
or U13446 (N_13446,N_11048,N_11285);
and U13447 (N_13447,N_11779,N_10528);
xor U13448 (N_13448,N_11726,N_11252);
or U13449 (N_13449,N_10596,N_10411);
nand U13450 (N_13450,N_10307,N_11192);
and U13451 (N_13451,N_11577,N_10044);
xor U13452 (N_13452,N_10701,N_11996);
xor U13453 (N_13453,N_11550,N_10622);
nor U13454 (N_13454,N_11010,N_11348);
xnor U13455 (N_13455,N_11684,N_10400);
nor U13456 (N_13456,N_11721,N_11187);
xor U13457 (N_13457,N_11408,N_11642);
and U13458 (N_13458,N_10336,N_10303);
nor U13459 (N_13459,N_10823,N_11184);
or U13460 (N_13460,N_10462,N_11603);
nor U13461 (N_13461,N_11584,N_10375);
or U13462 (N_13462,N_11665,N_10821);
or U13463 (N_13463,N_10308,N_11708);
nand U13464 (N_13464,N_11241,N_11690);
nor U13465 (N_13465,N_10134,N_10078);
xor U13466 (N_13466,N_10460,N_11697);
and U13467 (N_13467,N_10106,N_10059);
nand U13468 (N_13468,N_11158,N_11848);
nand U13469 (N_13469,N_10896,N_10558);
and U13470 (N_13470,N_11835,N_10477);
and U13471 (N_13471,N_11229,N_10696);
xnor U13472 (N_13472,N_11887,N_10449);
xor U13473 (N_13473,N_11355,N_11763);
nand U13474 (N_13474,N_10287,N_11009);
and U13475 (N_13475,N_10093,N_11652);
nor U13476 (N_13476,N_10621,N_11894);
and U13477 (N_13477,N_11768,N_11893);
nand U13478 (N_13478,N_10670,N_11643);
or U13479 (N_13479,N_11325,N_11050);
nor U13480 (N_13480,N_10232,N_11858);
xnor U13481 (N_13481,N_10055,N_10558);
and U13482 (N_13482,N_11589,N_10968);
xor U13483 (N_13483,N_11035,N_10950);
and U13484 (N_13484,N_10319,N_11712);
nand U13485 (N_13485,N_11923,N_10309);
nand U13486 (N_13486,N_10568,N_10335);
xnor U13487 (N_13487,N_11188,N_10376);
and U13488 (N_13488,N_11743,N_10637);
or U13489 (N_13489,N_10293,N_11706);
nor U13490 (N_13490,N_11713,N_10851);
nor U13491 (N_13491,N_10044,N_10750);
and U13492 (N_13492,N_11707,N_11514);
nand U13493 (N_13493,N_11905,N_10119);
xor U13494 (N_13494,N_10252,N_10027);
nor U13495 (N_13495,N_11229,N_11725);
and U13496 (N_13496,N_10633,N_10449);
xor U13497 (N_13497,N_11542,N_10567);
or U13498 (N_13498,N_11830,N_10605);
nand U13499 (N_13499,N_11557,N_11529);
nor U13500 (N_13500,N_11698,N_10976);
nor U13501 (N_13501,N_10973,N_10063);
nor U13502 (N_13502,N_11018,N_11024);
nor U13503 (N_13503,N_10036,N_11750);
or U13504 (N_13504,N_10631,N_10123);
or U13505 (N_13505,N_11906,N_11852);
and U13506 (N_13506,N_11748,N_10885);
nand U13507 (N_13507,N_11696,N_10937);
and U13508 (N_13508,N_10806,N_10066);
nor U13509 (N_13509,N_11974,N_10225);
or U13510 (N_13510,N_11652,N_11502);
nand U13511 (N_13511,N_10499,N_11049);
and U13512 (N_13512,N_10232,N_11487);
nand U13513 (N_13513,N_11372,N_11601);
and U13514 (N_13514,N_11887,N_11769);
nand U13515 (N_13515,N_11915,N_10437);
nand U13516 (N_13516,N_10290,N_10670);
or U13517 (N_13517,N_11898,N_10048);
nor U13518 (N_13518,N_10846,N_10885);
and U13519 (N_13519,N_10022,N_11961);
nor U13520 (N_13520,N_10822,N_11067);
or U13521 (N_13521,N_10352,N_11870);
nor U13522 (N_13522,N_11082,N_11382);
or U13523 (N_13523,N_11481,N_10048);
or U13524 (N_13524,N_10776,N_10117);
nor U13525 (N_13525,N_10046,N_10329);
nor U13526 (N_13526,N_10212,N_11571);
or U13527 (N_13527,N_11697,N_11182);
nand U13528 (N_13528,N_10920,N_11074);
nand U13529 (N_13529,N_10098,N_10143);
or U13530 (N_13530,N_11385,N_10116);
nor U13531 (N_13531,N_10237,N_10943);
nand U13532 (N_13532,N_11204,N_10066);
nor U13533 (N_13533,N_10208,N_11688);
and U13534 (N_13534,N_10128,N_10634);
xnor U13535 (N_13535,N_11152,N_10742);
nor U13536 (N_13536,N_10219,N_11248);
and U13537 (N_13537,N_11466,N_10288);
or U13538 (N_13538,N_11783,N_11252);
or U13539 (N_13539,N_10087,N_10195);
or U13540 (N_13540,N_10071,N_10015);
nor U13541 (N_13541,N_10621,N_11480);
nand U13542 (N_13542,N_11338,N_10035);
or U13543 (N_13543,N_10003,N_10044);
nand U13544 (N_13544,N_11390,N_11293);
or U13545 (N_13545,N_11890,N_10543);
xnor U13546 (N_13546,N_10471,N_10952);
or U13547 (N_13547,N_11436,N_10253);
or U13548 (N_13548,N_11210,N_10995);
or U13549 (N_13549,N_10274,N_11678);
nor U13550 (N_13550,N_11252,N_10379);
and U13551 (N_13551,N_10350,N_11247);
xnor U13552 (N_13552,N_11000,N_10074);
and U13553 (N_13553,N_11685,N_11743);
nor U13554 (N_13554,N_10877,N_11813);
and U13555 (N_13555,N_10213,N_11152);
xnor U13556 (N_13556,N_11806,N_11004);
nand U13557 (N_13557,N_11110,N_11645);
or U13558 (N_13558,N_10617,N_11435);
nor U13559 (N_13559,N_10572,N_10496);
and U13560 (N_13560,N_11272,N_11059);
xor U13561 (N_13561,N_11405,N_11610);
nand U13562 (N_13562,N_11442,N_11612);
nand U13563 (N_13563,N_11614,N_11851);
nand U13564 (N_13564,N_10345,N_11306);
nor U13565 (N_13565,N_10727,N_11827);
nand U13566 (N_13566,N_10420,N_10393);
or U13567 (N_13567,N_10141,N_11950);
or U13568 (N_13568,N_11088,N_10748);
or U13569 (N_13569,N_11347,N_10545);
nor U13570 (N_13570,N_11841,N_10054);
and U13571 (N_13571,N_10166,N_11882);
and U13572 (N_13572,N_11418,N_10985);
and U13573 (N_13573,N_11281,N_10354);
and U13574 (N_13574,N_11637,N_10121);
or U13575 (N_13575,N_11688,N_10281);
nand U13576 (N_13576,N_10095,N_11605);
xnor U13577 (N_13577,N_11163,N_11455);
xor U13578 (N_13578,N_11322,N_10039);
nor U13579 (N_13579,N_10075,N_11130);
and U13580 (N_13580,N_11227,N_10899);
nand U13581 (N_13581,N_11140,N_10340);
or U13582 (N_13582,N_10363,N_11668);
or U13583 (N_13583,N_11768,N_11169);
and U13584 (N_13584,N_10061,N_10200);
xor U13585 (N_13585,N_10208,N_11560);
nor U13586 (N_13586,N_10298,N_11623);
nand U13587 (N_13587,N_10479,N_10545);
nand U13588 (N_13588,N_10341,N_10745);
or U13589 (N_13589,N_11987,N_11900);
nor U13590 (N_13590,N_11696,N_10203);
xnor U13591 (N_13591,N_11313,N_11155);
and U13592 (N_13592,N_11469,N_10608);
and U13593 (N_13593,N_10727,N_11246);
xnor U13594 (N_13594,N_10278,N_10625);
nor U13595 (N_13595,N_11159,N_11083);
or U13596 (N_13596,N_10476,N_10426);
and U13597 (N_13597,N_10523,N_10454);
nand U13598 (N_13598,N_10193,N_11658);
or U13599 (N_13599,N_10034,N_11938);
and U13600 (N_13600,N_10544,N_11556);
or U13601 (N_13601,N_11185,N_11589);
and U13602 (N_13602,N_10860,N_11114);
xnor U13603 (N_13603,N_11107,N_11101);
or U13604 (N_13604,N_11159,N_11024);
nor U13605 (N_13605,N_11386,N_10157);
or U13606 (N_13606,N_10952,N_11025);
nand U13607 (N_13607,N_10055,N_10514);
nand U13608 (N_13608,N_11289,N_11137);
nor U13609 (N_13609,N_10870,N_10233);
xnor U13610 (N_13610,N_11302,N_11344);
nor U13611 (N_13611,N_10268,N_11111);
or U13612 (N_13612,N_11044,N_11924);
and U13613 (N_13613,N_11918,N_11720);
nand U13614 (N_13614,N_11021,N_11323);
or U13615 (N_13615,N_11216,N_10697);
and U13616 (N_13616,N_10849,N_11926);
xor U13617 (N_13617,N_11944,N_11569);
xnor U13618 (N_13618,N_11832,N_10041);
nand U13619 (N_13619,N_11471,N_10573);
or U13620 (N_13620,N_10575,N_11381);
nor U13621 (N_13621,N_10363,N_10775);
nor U13622 (N_13622,N_10307,N_11263);
xor U13623 (N_13623,N_10575,N_10410);
xor U13624 (N_13624,N_10869,N_11577);
and U13625 (N_13625,N_10635,N_11869);
and U13626 (N_13626,N_10261,N_10910);
and U13627 (N_13627,N_11443,N_11095);
xor U13628 (N_13628,N_11073,N_11971);
and U13629 (N_13629,N_10824,N_11231);
and U13630 (N_13630,N_11592,N_10467);
nand U13631 (N_13631,N_11733,N_10522);
nor U13632 (N_13632,N_10840,N_10194);
nor U13633 (N_13633,N_10777,N_10222);
and U13634 (N_13634,N_10490,N_11601);
xnor U13635 (N_13635,N_10489,N_10411);
nand U13636 (N_13636,N_10170,N_10103);
and U13637 (N_13637,N_10221,N_11772);
nand U13638 (N_13638,N_11655,N_10514);
xnor U13639 (N_13639,N_11485,N_11317);
nand U13640 (N_13640,N_10218,N_10533);
xor U13641 (N_13641,N_10779,N_10633);
or U13642 (N_13642,N_11864,N_10344);
nor U13643 (N_13643,N_10119,N_10624);
xor U13644 (N_13644,N_10771,N_11923);
and U13645 (N_13645,N_11510,N_10831);
nor U13646 (N_13646,N_10218,N_10485);
or U13647 (N_13647,N_10385,N_10959);
and U13648 (N_13648,N_10093,N_11373);
or U13649 (N_13649,N_11777,N_10002);
nor U13650 (N_13650,N_11654,N_10892);
nand U13651 (N_13651,N_10199,N_10928);
or U13652 (N_13652,N_10122,N_11413);
xnor U13653 (N_13653,N_11863,N_11504);
or U13654 (N_13654,N_10816,N_10558);
nor U13655 (N_13655,N_11613,N_10027);
nand U13656 (N_13656,N_10424,N_10354);
xor U13657 (N_13657,N_10912,N_11119);
and U13658 (N_13658,N_11881,N_11907);
and U13659 (N_13659,N_11259,N_10768);
nand U13660 (N_13660,N_10369,N_10216);
or U13661 (N_13661,N_11216,N_10016);
or U13662 (N_13662,N_11316,N_10888);
xor U13663 (N_13663,N_10392,N_10117);
or U13664 (N_13664,N_11811,N_10699);
xor U13665 (N_13665,N_10381,N_10872);
nand U13666 (N_13666,N_10300,N_10965);
xnor U13667 (N_13667,N_11067,N_11056);
or U13668 (N_13668,N_11935,N_10599);
nor U13669 (N_13669,N_11718,N_11175);
and U13670 (N_13670,N_10369,N_10513);
xnor U13671 (N_13671,N_10924,N_11106);
or U13672 (N_13672,N_11134,N_10264);
nand U13673 (N_13673,N_10236,N_11624);
and U13674 (N_13674,N_11025,N_10960);
or U13675 (N_13675,N_11624,N_10486);
nor U13676 (N_13676,N_10113,N_11194);
or U13677 (N_13677,N_11423,N_10891);
and U13678 (N_13678,N_11270,N_10467);
xor U13679 (N_13679,N_10491,N_11651);
nor U13680 (N_13680,N_11693,N_11746);
xor U13681 (N_13681,N_11321,N_11920);
or U13682 (N_13682,N_11291,N_11990);
nand U13683 (N_13683,N_10191,N_11698);
xor U13684 (N_13684,N_10424,N_10136);
nand U13685 (N_13685,N_11077,N_10563);
nand U13686 (N_13686,N_11175,N_11999);
nand U13687 (N_13687,N_10924,N_10469);
and U13688 (N_13688,N_10922,N_10678);
nor U13689 (N_13689,N_10783,N_10181);
nand U13690 (N_13690,N_11262,N_11272);
and U13691 (N_13691,N_10593,N_10311);
or U13692 (N_13692,N_10103,N_10835);
nor U13693 (N_13693,N_11703,N_10429);
xor U13694 (N_13694,N_11540,N_10293);
nand U13695 (N_13695,N_11901,N_11893);
or U13696 (N_13696,N_11676,N_10756);
and U13697 (N_13697,N_10269,N_11823);
or U13698 (N_13698,N_10527,N_10415);
nand U13699 (N_13699,N_11769,N_10352);
and U13700 (N_13700,N_10009,N_11206);
or U13701 (N_13701,N_10879,N_11824);
or U13702 (N_13702,N_10863,N_11833);
nand U13703 (N_13703,N_11851,N_10771);
nand U13704 (N_13704,N_10385,N_11708);
and U13705 (N_13705,N_11059,N_10126);
and U13706 (N_13706,N_10113,N_10135);
and U13707 (N_13707,N_11005,N_11143);
or U13708 (N_13708,N_10935,N_11066);
nor U13709 (N_13709,N_10698,N_11501);
xnor U13710 (N_13710,N_10249,N_10396);
nor U13711 (N_13711,N_10762,N_11513);
nand U13712 (N_13712,N_11189,N_11969);
nor U13713 (N_13713,N_11520,N_10162);
or U13714 (N_13714,N_11004,N_11324);
nor U13715 (N_13715,N_11097,N_11121);
nor U13716 (N_13716,N_10180,N_10783);
or U13717 (N_13717,N_11315,N_11840);
and U13718 (N_13718,N_11586,N_11551);
xnor U13719 (N_13719,N_10390,N_11404);
and U13720 (N_13720,N_11063,N_11592);
xnor U13721 (N_13721,N_11446,N_10628);
xor U13722 (N_13722,N_10635,N_11926);
or U13723 (N_13723,N_11535,N_11898);
nor U13724 (N_13724,N_11009,N_11287);
or U13725 (N_13725,N_11292,N_10981);
and U13726 (N_13726,N_10898,N_10960);
xor U13727 (N_13727,N_10041,N_10943);
nor U13728 (N_13728,N_10546,N_11667);
nor U13729 (N_13729,N_11802,N_10100);
nand U13730 (N_13730,N_11414,N_11018);
xnor U13731 (N_13731,N_11544,N_10843);
and U13732 (N_13732,N_10100,N_11116);
nand U13733 (N_13733,N_10534,N_11981);
or U13734 (N_13734,N_11332,N_10732);
nand U13735 (N_13735,N_10136,N_10323);
nand U13736 (N_13736,N_10290,N_11154);
or U13737 (N_13737,N_11529,N_10414);
xor U13738 (N_13738,N_10454,N_10308);
xnor U13739 (N_13739,N_10784,N_10291);
nor U13740 (N_13740,N_11687,N_11326);
and U13741 (N_13741,N_11204,N_11289);
xor U13742 (N_13742,N_11609,N_10052);
nor U13743 (N_13743,N_11737,N_10615);
xor U13744 (N_13744,N_11322,N_10773);
xor U13745 (N_13745,N_11034,N_10676);
xor U13746 (N_13746,N_11053,N_11766);
or U13747 (N_13747,N_10869,N_10879);
nand U13748 (N_13748,N_11616,N_10280);
nor U13749 (N_13749,N_10252,N_10455);
or U13750 (N_13750,N_11044,N_11042);
xor U13751 (N_13751,N_11839,N_11580);
nor U13752 (N_13752,N_11405,N_11922);
nor U13753 (N_13753,N_10160,N_11920);
xnor U13754 (N_13754,N_11791,N_10554);
or U13755 (N_13755,N_10957,N_10576);
and U13756 (N_13756,N_11803,N_10341);
nor U13757 (N_13757,N_11177,N_11575);
nand U13758 (N_13758,N_10010,N_10291);
nor U13759 (N_13759,N_11306,N_10920);
or U13760 (N_13760,N_11892,N_11203);
and U13761 (N_13761,N_11150,N_10917);
or U13762 (N_13762,N_11289,N_10538);
nor U13763 (N_13763,N_11618,N_11427);
nor U13764 (N_13764,N_11542,N_10679);
nand U13765 (N_13765,N_11047,N_11531);
and U13766 (N_13766,N_10064,N_11126);
xnor U13767 (N_13767,N_10519,N_10200);
and U13768 (N_13768,N_11876,N_11907);
xnor U13769 (N_13769,N_10052,N_10558);
nand U13770 (N_13770,N_10840,N_11366);
xor U13771 (N_13771,N_10326,N_11876);
nand U13772 (N_13772,N_11507,N_10917);
and U13773 (N_13773,N_10455,N_10154);
nor U13774 (N_13774,N_11677,N_11801);
xor U13775 (N_13775,N_11469,N_10954);
nor U13776 (N_13776,N_11624,N_11459);
xnor U13777 (N_13777,N_11801,N_11017);
nand U13778 (N_13778,N_11314,N_10660);
or U13779 (N_13779,N_11418,N_11482);
nand U13780 (N_13780,N_11093,N_11104);
or U13781 (N_13781,N_10459,N_11043);
or U13782 (N_13782,N_10678,N_10734);
or U13783 (N_13783,N_10812,N_10014);
nand U13784 (N_13784,N_10265,N_11721);
or U13785 (N_13785,N_11983,N_11180);
or U13786 (N_13786,N_11553,N_11108);
nor U13787 (N_13787,N_11638,N_11589);
and U13788 (N_13788,N_10949,N_10938);
and U13789 (N_13789,N_10022,N_11088);
nand U13790 (N_13790,N_10770,N_10213);
nand U13791 (N_13791,N_11041,N_11213);
xnor U13792 (N_13792,N_10889,N_11998);
and U13793 (N_13793,N_10554,N_10056);
or U13794 (N_13794,N_11625,N_11194);
nor U13795 (N_13795,N_10618,N_11886);
nor U13796 (N_13796,N_11990,N_11164);
nand U13797 (N_13797,N_11425,N_11226);
nand U13798 (N_13798,N_10358,N_10186);
or U13799 (N_13799,N_10894,N_11929);
nand U13800 (N_13800,N_11021,N_11865);
or U13801 (N_13801,N_11076,N_11616);
or U13802 (N_13802,N_10440,N_10007);
or U13803 (N_13803,N_10555,N_11641);
nand U13804 (N_13804,N_10539,N_11672);
xor U13805 (N_13805,N_10721,N_10060);
nor U13806 (N_13806,N_11712,N_11643);
nand U13807 (N_13807,N_11918,N_10750);
or U13808 (N_13808,N_10155,N_11690);
or U13809 (N_13809,N_11384,N_10131);
nand U13810 (N_13810,N_11639,N_11746);
nor U13811 (N_13811,N_10172,N_10334);
and U13812 (N_13812,N_10846,N_10748);
xor U13813 (N_13813,N_10673,N_10966);
xor U13814 (N_13814,N_11756,N_10915);
and U13815 (N_13815,N_11207,N_10908);
and U13816 (N_13816,N_11076,N_10535);
and U13817 (N_13817,N_11766,N_11918);
xnor U13818 (N_13818,N_11839,N_11742);
or U13819 (N_13819,N_10029,N_10935);
nand U13820 (N_13820,N_11075,N_11747);
or U13821 (N_13821,N_10905,N_11945);
or U13822 (N_13822,N_10497,N_10799);
nor U13823 (N_13823,N_10925,N_10418);
or U13824 (N_13824,N_11209,N_11488);
and U13825 (N_13825,N_10317,N_11031);
or U13826 (N_13826,N_11868,N_11032);
or U13827 (N_13827,N_10878,N_10994);
xnor U13828 (N_13828,N_10760,N_11518);
nand U13829 (N_13829,N_11385,N_11771);
nand U13830 (N_13830,N_11449,N_11536);
nor U13831 (N_13831,N_10688,N_10771);
nor U13832 (N_13832,N_11644,N_11653);
and U13833 (N_13833,N_10167,N_11231);
or U13834 (N_13834,N_11846,N_10739);
nand U13835 (N_13835,N_10530,N_10342);
nor U13836 (N_13836,N_11984,N_11766);
xor U13837 (N_13837,N_11911,N_11365);
nor U13838 (N_13838,N_10826,N_11636);
nor U13839 (N_13839,N_11059,N_10121);
and U13840 (N_13840,N_11269,N_10940);
xor U13841 (N_13841,N_10857,N_11339);
and U13842 (N_13842,N_10274,N_11522);
or U13843 (N_13843,N_10480,N_11392);
nor U13844 (N_13844,N_11376,N_11184);
and U13845 (N_13845,N_11163,N_10099);
nand U13846 (N_13846,N_11886,N_10817);
and U13847 (N_13847,N_11615,N_11519);
or U13848 (N_13848,N_10168,N_10495);
or U13849 (N_13849,N_10940,N_11914);
and U13850 (N_13850,N_11630,N_11954);
nor U13851 (N_13851,N_10387,N_10040);
nor U13852 (N_13852,N_10304,N_11610);
nand U13853 (N_13853,N_11122,N_10306);
xor U13854 (N_13854,N_10435,N_11223);
nor U13855 (N_13855,N_10001,N_11973);
nor U13856 (N_13856,N_10433,N_10216);
nand U13857 (N_13857,N_11027,N_10892);
and U13858 (N_13858,N_11853,N_11656);
nand U13859 (N_13859,N_11104,N_11833);
xnor U13860 (N_13860,N_11838,N_11701);
nor U13861 (N_13861,N_10737,N_10678);
or U13862 (N_13862,N_10203,N_10209);
or U13863 (N_13863,N_10989,N_10254);
nor U13864 (N_13864,N_10752,N_10906);
nor U13865 (N_13865,N_11234,N_11216);
nand U13866 (N_13866,N_11538,N_10618);
xnor U13867 (N_13867,N_10112,N_10570);
xnor U13868 (N_13868,N_10333,N_11352);
and U13869 (N_13869,N_10065,N_11485);
xnor U13870 (N_13870,N_10149,N_10211);
nor U13871 (N_13871,N_10112,N_10660);
nor U13872 (N_13872,N_10119,N_10566);
nor U13873 (N_13873,N_10307,N_11174);
xor U13874 (N_13874,N_10662,N_11540);
nor U13875 (N_13875,N_11542,N_11459);
nor U13876 (N_13876,N_11400,N_10393);
and U13877 (N_13877,N_11776,N_11770);
xor U13878 (N_13878,N_11367,N_11311);
nand U13879 (N_13879,N_10842,N_10067);
xnor U13880 (N_13880,N_11874,N_10122);
and U13881 (N_13881,N_10791,N_10122);
nand U13882 (N_13882,N_10322,N_10864);
xor U13883 (N_13883,N_10978,N_11242);
or U13884 (N_13884,N_10464,N_11538);
or U13885 (N_13885,N_11694,N_10827);
nand U13886 (N_13886,N_11798,N_10285);
and U13887 (N_13887,N_11168,N_11431);
nor U13888 (N_13888,N_11981,N_10286);
nor U13889 (N_13889,N_10367,N_11787);
xnor U13890 (N_13890,N_11173,N_11752);
and U13891 (N_13891,N_11717,N_11360);
nor U13892 (N_13892,N_11878,N_10412);
or U13893 (N_13893,N_11875,N_11685);
and U13894 (N_13894,N_11347,N_10171);
nand U13895 (N_13895,N_10903,N_10522);
or U13896 (N_13896,N_10136,N_11131);
nand U13897 (N_13897,N_11490,N_11900);
nand U13898 (N_13898,N_10704,N_11201);
xor U13899 (N_13899,N_10320,N_11221);
nand U13900 (N_13900,N_10941,N_10866);
nor U13901 (N_13901,N_11444,N_11091);
and U13902 (N_13902,N_11105,N_10885);
or U13903 (N_13903,N_10272,N_10126);
nor U13904 (N_13904,N_11984,N_10295);
or U13905 (N_13905,N_10401,N_11560);
or U13906 (N_13906,N_11872,N_11548);
or U13907 (N_13907,N_11955,N_11132);
xnor U13908 (N_13908,N_11905,N_11174);
or U13909 (N_13909,N_11518,N_11464);
xnor U13910 (N_13910,N_11899,N_11161);
xor U13911 (N_13911,N_11917,N_11694);
and U13912 (N_13912,N_10903,N_11883);
nor U13913 (N_13913,N_11830,N_10043);
or U13914 (N_13914,N_11078,N_11732);
xor U13915 (N_13915,N_10235,N_11243);
nor U13916 (N_13916,N_11944,N_10696);
nor U13917 (N_13917,N_11172,N_10049);
nor U13918 (N_13918,N_10916,N_11535);
xnor U13919 (N_13919,N_10974,N_11790);
and U13920 (N_13920,N_10526,N_10985);
nand U13921 (N_13921,N_11085,N_11826);
nand U13922 (N_13922,N_11038,N_11398);
and U13923 (N_13923,N_10591,N_10277);
or U13924 (N_13924,N_11903,N_11799);
and U13925 (N_13925,N_11691,N_10632);
xnor U13926 (N_13926,N_10371,N_10972);
nor U13927 (N_13927,N_10569,N_10326);
or U13928 (N_13928,N_10946,N_11118);
and U13929 (N_13929,N_11670,N_11372);
nand U13930 (N_13930,N_11066,N_11690);
and U13931 (N_13931,N_11934,N_10710);
xnor U13932 (N_13932,N_11316,N_10629);
nand U13933 (N_13933,N_11194,N_11777);
and U13934 (N_13934,N_11806,N_10778);
nor U13935 (N_13935,N_10072,N_11352);
or U13936 (N_13936,N_10765,N_10556);
or U13937 (N_13937,N_11315,N_11519);
or U13938 (N_13938,N_10468,N_10386);
nand U13939 (N_13939,N_11587,N_11716);
and U13940 (N_13940,N_11294,N_10152);
or U13941 (N_13941,N_11784,N_11411);
nand U13942 (N_13942,N_11134,N_10182);
nand U13943 (N_13943,N_10318,N_11306);
and U13944 (N_13944,N_11897,N_10506);
nand U13945 (N_13945,N_10541,N_10574);
and U13946 (N_13946,N_11588,N_11225);
or U13947 (N_13947,N_11000,N_11662);
xor U13948 (N_13948,N_10981,N_10684);
or U13949 (N_13949,N_11765,N_11245);
or U13950 (N_13950,N_11873,N_11269);
nor U13951 (N_13951,N_11223,N_11244);
nand U13952 (N_13952,N_10091,N_11581);
nor U13953 (N_13953,N_11928,N_10968);
nor U13954 (N_13954,N_11988,N_10076);
xnor U13955 (N_13955,N_10967,N_11317);
nor U13956 (N_13956,N_11216,N_11920);
xor U13957 (N_13957,N_11593,N_11630);
nor U13958 (N_13958,N_10630,N_11563);
nor U13959 (N_13959,N_11385,N_10155);
nor U13960 (N_13960,N_10835,N_10514);
nand U13961 (N_13961,N_11388,N_10259);
and U13962 (N_13962,N_11249,N_11860);
xnor U13963 (N_13963,N_11798,N_10129);
nor U13964 (N_13964,N_10611,N_10876);
nor U13965 (N_13965,N_11188,N_10721);
nand U13966 (N_13966,N_10915,N_10108);
nor U13967 (N_13967,N_11041,N_10613);
nor U13968 (N_13968,N_10599,N_10643);
or U13969 (N_13969,N_10627,N_11231);
xnor U13970 (N_13970,N_11635,N_10635);
xnor U13971 (N_13971,N_10677,N_10887);
nor U13972 (N_13972,N_10398,N_10977);
and U13973 (N_13973,N_10855,N_11545);
nand U13974 (N_13974,N_10834,N_11471);
and U13975 (N_13975,N_10524,N_10334);
nor U13976 (N_13976,N_10879,N_11277);
nor U13977 (N_13977,N_10667,N_10154);
xnor U13978 (N_13978,N_11444,N_10586);
and U13979 (N_13979,N_10976,N_11477);
nor U13980 (N_13980,N_11429,N_11784);
or U13981 (N_13981,N_11431,N_10870);
nand U13982 (N_13982,N_11450,N_10014);
nor U13983 (N_13983,N_10561,N_10000);
and U13984 (N_13984,N_10104,N_10460);
and U13985 (N_13985,N_10596,N_11194);
nand U13986 (N_13986,N_10791,N_10844);
nand U13987 (N_13987,N_10556,N_10191);
or U13988 (N_13988,N_11126,N_11556);
nor U13989 (N_13989,N_11836,N_11214);
and U13990 (N_13990,N_11921,N_11995);
xnor U13991 (N_13991,N_10586,N_11017);
nor U13992 (N_13992,N_11899,N_11516);
nor U13993 (N_13993,N_11603,N_11162);
nand U13994 (N_13994,N_10157,N_10313);
nor U13995 (N_13995,N_11975,N_11700);
nor U13996 (N_13996,N_11771,N_10973);
and U13997 (N_13997,N_10211,N_10558);
and U13998 (N_13998,N_11201,N_10748);
nand U13999 (N_13999,N_10286,N_11994);
nor U14000 (N_14000,N_12678,N_12745);
or U14001 (N_14001,N_12279,N_12626);
xnor U14002 (N_14002,N_12668,N_13584);
nor U14003 (N_14003,N_13705,N_12784);
xor U14004 (N_14004,N_12005,N_13582);
xor U14005 (N_14005,N_13749,N_13733);
and U14006 (N_14006,N_13998,N_13549);
xor U14007 (N_14007,N_12473,N_12887);
and U14008 (N_14008,N_13277,N_13695);
nand U14009 (N_14009,N_12184,N_12709);
xor U14010 (N_14010,N_13264,N_12409);
and U14011 (N_14011,N_13445,N_12810);
nor U14012 (N_14012,N_13250,N_13873);
nor U14013 (N_14013,N_12416,N_13910);
or U14014 (N_14014,N_12286,N_12221);
xor U14015 (N_14015,N_12646,N_13139);
xnor U14016 (N_14016,N_12202,N_13049);
and U14017 (N_14017,N_12232,N_13259);
and U14018 (N_14018,N_13073,N_13739);
or U14019 (N_14019,N_13794,N_13260);
xnor U14020 (N_14020,N_13058,N_12431);
xor U14021 (N_14021,N_12971,N_13334);
nor U14022 (N_14022,N_12871,N_12213);
xor U14023 (N_14023,N_12450,N_12345);
xnor U14024 (N_14024,N_12151,N_13692);
nand U14025 (N_14025,N_12837,N_13123);
nand U14026 (N_14026,N_12956,N_12672);
nor U14027 (N_14027,N_12856,N_12911);
or U14028 (N_14028,N_13978,N_13149);
xnor U14029 (N_14029,N_12316,N_13649);
xor U14030 (N_14030,N_12739,N_12460);
xnor U14031 (N_14031,N_12650,N_12240);
xnor U14032 (N_14032,N_13187,N_13542);
or U14033 (N_14033,N_13252,N_12660);
and U14034 (N_14034,N_13031,N_13848);
or U14035 (N_14035,N_13239,N_12259);
xor U14036 (N_14036,N_12265,N_13107);
and U14037 (N_14037,N_12950,N_13147);
nand U14038 (N_14038,N_13788,N_13092);
nor U14039 (N_14039,N_12793,N_12860);
or U14040 (N_14040,N_12169,N_12145);
nor U14041 (N_14041,N_13625,N_13764);
nor U14042 (N_14042,N_12116,N_12456);
nor U14043 (N_14043,N_12329,N_12731);
or U14044 (N_14044,N_12719,N_12025);
and U14045 (N_14045,N_13547,N_13833);
nor U14046 (N_14046,N_12912,N_13245);
nand U14047 (N_14047,N_12146,N_12339);
nand U14048 (N_14048,N_12968,N_13561);
nand U14049 (N_14049,N_13660,N_13479);
nor U14050 (N_14050,N_13249,N_13784);
nand U14051 (N_14051,N_12225,N_12595);
and U14052 (N_14052,N_13867,N_13986);
nor U14053 (N_14053,N_13436,N_12804);
nand U14054 (N_14054,N_13514,N_12308);
or U14055 (N_14055,N_13106,N_13229);
or U14056 (N_14056,N_13418,N_12640);
xnor U14057 (N_14057,N_12051,N_12104);
xor U14058 (N_14058,N_12742,N_13127);
nand U14059 (N_14059,N_12740,N_13129);
and U14060 (N_14060,N_12323,N_12870);
and U14061 (N_14061,N_13940,N_12497);
nor U14062 (N_14062,N_12771,N_12774);
or U14063 (N_14063,N_12762,N_12717);
xnor U14064 (N_14064,N_12189,N_12706);
nand U14065 (N_14065,N_13911,N_12182);
and U14066 (N_14066,N_13120,N_13521);
xnor U14067 (N_14067,N_13415,N_13932);
nor U14068 (N_14068,N_13390,N_13208);
nand U14069 (N_14069,N_12724,N_13172);
nand U14070 (N_14070,N_13146,N_12609);
nor U14071 (N_14071,N_12734,N_12920);
xnor U14072 (N_14072,N_12233,N_13484);
nand U14073 (N_14073,N_13079,N_13237);
nand U14074 (N_14074,N_12608,N_13019);
xnor U14075 (N_14075,N_12055,N_12273);
or U14076 (N_14076,N_13592,N_13642);
xor U14077 (N_14077,N_13078,N_12236);
nand U14078 (N_14078,N_12092,N_13340);
nand U14079 (N_14079,N_12970,N_13011);
xor U14080 (N_14080,N_13095,N_13556);
and U14081 (N_14081,N_13723,N_12004);
and U14082 (N_14082,N_13992,N_13879);
xor U14083 (N_14083,N_13022,N_13295);
or U14084 (N_14084,N_12661,N_13615);
or U14085 (N_14085,N_13718,N_12079);
nand U14086 (N_14086,N_13033,N_13708);
nand U14087 (N_14087,N_13535,N_13388);
nand U14088 (N_14088,N_12113,N_12297);
xor U14089 (N_14089,N_12832,N_13770);
and U14090 (N_14090,N_12399,N_12099);
and U14091 (N_14091,N_13319,N_13168);
and U14092 (N_14092,N_13653,N_12040);
nor U14093 (N_14093,N_12061,N_13412);
and U14094 (N_14094,N_12546,N_13359);
nand U14095 (N_14095,N_12635,N_13533);
nor U14096 (N_14096,N_13899,N_13368);
xnor U14097 (N_14097,N_13894,N_12893);
nor U14098 (N_14098,N_13071,N_12611);
xor U14099 (N_14099,N_13581,N_12052);
xnor U14100 (N_14100,N_13552,N_13416);
or U14101 (N_14101,N_12408,N_13793);
and U14102 (N_14102,N_12375,N_13905);
xnor U14103 (N_14103,N_13975,N_12226);
or U14104 (N_14104,N_12934,N_13750);
nand U14105 (N_14105,N_12868,N_12366);
nand U14106 (N_14106,N_13673,N_13009);
nand U14107 (N_14107,N_12000,N_12536);
nand U14108 (N_14108,N_13765,N_13385);
or U14109 (N_14109,N_12918,N_12899);
nand U14110 (N_14110,N_12303,N_13926);
nand U14111 (N_14111,N_13667,N_12384);
and U14112 (N_14112,N_13101,N_13357);
nor U14113 (N_14113,N_13468,N_13288);
nor U14114 (N_14114,N_13613,N_12886);
xnor U14115 (N_14115,N_12892,N_13029);
and U14116 (N_14116,N_13039,N_13866);
and U14117 (N_14117,N_13456,N_13119);
or U14118 (N_14118,N_13504,N_12154);
nand U14119 (N_14119,N_12959,N_13994);
and U14120 (N_14120,N_12948,N_12614);
nand U14121 (N_14121,N_12435,N_12618);
and U14122 (N_14122,N_12074,N_12861);
and U14123 (N_14123,N_12160,N_13666);
nor U14124 (N_14124,N_13499,N_13554);
xnor U14125 (N_14125,N_13353,N_13137);
nor U14126 (N_14126,N_13644,N_12035);
nand U14127 (N_14127,N_13217,N_13448);
or U14128 (N_14128,N_13602,N_12754);
xnor U14129 (N_14129,N_13763,N_13989);
nand U14130 (N_14130,N_13186,N_12991);
nor U14131 (N_14131,N_13382,N_12597);
nand U14132 (N_14132,N_13800,N_12628);
nand U14133 (N_14133,N_13324,N_13293);
xnor U14134 (N_14134,N_12556,N_13111);
nand U14135 (N_14135,N_12028,N_12364);
nor U14136 (N_14136,N_13704,N_12328);
xnor U14137 (N_14137,N_13219,N_12951);
nor U14138 (N_14138,N_12667,N_13849);
or U14139 (N_14139,N_12508,N_13462);
nand U14140 (N_14140,N_12965,N_13795);
and U14141 (N_14141,N_13636,N_13258);
nor U14142 (N_14142,N_12819,N_12922);
nand U14143 (N_14143,N_12442,N_13893);
and U14144 (N_14144,N_12823,N_13752);
xor U14145 (N_14145,N_12209,N_12685);
or U14146 (N_14146,N_12673,N_13426);
and U14147 (N_14147,N_13256,N_13929);
nand U14148 (N_14148,N_12797,N_13224);
xor U14149 (N_14149,N_12084,N_12507);
or U14150 (N_14150,N_12141,N_12166);
or U14151 (N_14151,N_12007,N_12142);
or U14152 (N_14152,N_12386,N_12287);
xor U14153 (N_14153,N_12923,N_13278);
or U14154 (N_14154,N_13045,N_12326);
nand U14155 (N_14155,N_12398,N_13375);
xnor U14156 (N_14156,N_13883,N_13126);
or U14157 (N_14157,N_12479,N_13493);
xor U14158 (N_14158,N_12124,N_13344);
nand U14159 (N_14159,N_13452,N_12088);
xor U14160 (N_14160,N_13842,N_13774);
or U14161 (N_14161,N_13315,N_12363);
nand U14162 (N_14162,N_12835,N_12484);
nor U14163 (N_14163,N_12163,N_12809);
nor U14164 (N_14164,N_13656,N_12670);
xor U14165 (N_14165,N_12468,N_13672);
nor U14166 (N_14166,N_13616,N_12231);
nor U14167 (N_14167,N_13059,N_13401);
xor U14168 (N_14168,N_12952,N_12068);
nor U14169 (N_14169,N_12540,N_12926);
nor U14170 (N_14170,N_12177,N_13691);
nand U14171 (N_14171,N_13302,N_13373);
nor U14172 (N_14172,N_12583,N_13520);
and U14173 (N_14173,N_13417,N_12302);
xor U14174 (N_14174,N_12347,N_13182);
or U14175 (N_14175,N_13906,N_13051);
nor U14176 (N_14176,N_12982,N_13527);
nor U14177 (N_14177,N_12106,N_12176);
nand U14178 (N_14178,N_12657,N_12137);
nor U14179 (N_14179,N_12346,N_12524);
xor U14180 (N_14180,N_13920,N_12790);
nor U14181 (N_14181,N_12187,N_13222);
nor U14182 (N_14182,N_12758,N_12291);
xor U14183 (N_14183,N_13701,N_13632);
xnor U14184 (N_14184,N_13036,N_12907);
and U14185 (N_14185,N_13394,N_12331);
nand U14186 (N_14186,N_13367,N_13458);
or U14187 (N_14187,N_12630,N_12437);
nor U14188 (N_14188,N_12144,N_13060);
nor U14189 (N_14189,N_13698,N_13934);
xnor U14190 (N_14190,N_12714,N_12586);
nor U14191 (N_14191,N_13536,N_12889);
and U14192 (N_14192,N_12420,N_12716);
xor U14193 (N_14193,N_13709,N_13944);
nand U14194 (N_14194,N_13973,N_13604);
nand U14195 (N_14195,N_12275,N_13610);
nand U14196 (N_14196,N_13122,N_13922);
xnor U14197 (N_14197,N_13886,N_12876);
nor U14198 (N_14198,N_12200,N_12537);
xor U14199 (N_14199,N_13465,N_13786);
nor U14200 (N_14200,N_13726,N_12281);
nand U14201 (N_14201,N_12374,N_12400);
and U14202 (N_14202,N_12593,N_12503);
nor U14203 (N_14203,N_12422,N_13745);
and U14204 (N_14204,N_12909,N_12094);
nor U14205 (N_14205,N_13803,N_12805);
nor U14206 (N_14206,N_13568,N_12263);
nor U14207 (N_14207,N_13635,N_12875);
and U14208 (N_14208,N_12150,N_13952);
or U14209 (N_14209,N_13303,N_13880);
nor U14210 (N_14210,N_12481,N_12551);
nor U14211 (N_14211,N_13606,N_12833);
or U14212 (N_14212,N_12188,N_13280);
or U14213 (N_14213,N_12368,N_12550);
nor U14214 (N_14214,N_12625,N_13938);
nand U14215 (N_14215,N_13969,N_13690);
nor U14216 (N_14216,N_12278,N_13299);
xnor U14217 (N_14217,N_13243,N_12012);
xor U14218 (N_14218,N_13735,N_12223);
and U14219 (N_14219,N_13518,N_12489);
or U14220 (N_14220,N_13835,N_12836);
nand U14221 (N_14221,N_12394,N_12987);
nor U14222 (N_14222,N_12679,N_13016);
xor U14223 (N_14223,N_13464,N_12781);
nand U14224 (N_14224,N_12598,N_12652);
and U14225 (N_14225,N_13025,N_12649);
nor U14226 (N_14226,N_12973,N_13083);
or U14227 (N_14227,N_12541,N_13943);
xnor U14228 (N_14228,N_13050,N_12534);
or U14229 (N_14229,N_12268,N_13525);
xor U14230 (N_14230,N_12908,N_12057);
nand U14231 (N_14231,N_13289,N_12696);
and U14232 (N_14232,N_13196,N_12186);
or U14233 (N_14233,N_13169,N_13034);
and U14234 (N_14234,N_13366,N_13273);
nor U14235 (N_14235,N_12885,N_13870);
and U14236 (N_14236,N_13771,N_13790);
nand U14237 (N_14237,N_13242,N_13980);
or U14238 (N_14238,N_13055,N_13189);
nand U14239 (N_14239,N_12462,N_12319);
nor U14240 (N_14240,N_12372,N_12874);
xor U14241 (N_14241,N_12568,N_13837);
or U14242 (N_14242,N_13395,N_13824);
or U14243 (N_14243,N_12882,N_13223);
or U14244 (N_14244,N_12750,N_12834);
xnor U14245 (N_14245,N_13074,N_13724);
nand U14246 (N_14246,N_13204,N_13634);
xor U14247 (N_14247,N_12822,N_13668);
or U14248 (N_14248,N_13159,N_13348);
xor U14249 (N_14249,N_12808,N_13676);
nand U14250 (N_14250,N_13915,N_13335);
nor U14251 (N_14251,N_13455,N_13453);
xnor U14252 (N_14252,N_13342,N_12691);
nand U14253 (N_14253,N_13398,N_12463);
nor U14254 (N_14254,N_13290,N_12410);
or U14255 (N_14255,N_12975,N_13825);
nor U14256 (N_14256,N_12490,N_13816);
and U14257 (N_14257,N_12304,N_13160);
xor U14258 (N_14258,N_12299,N_12501);
nor U14259 (N_14259,N_13102,N_13865);
and U14260 (N_14260,N_12054,N_13946);
nor U14261 (N_14261,N_12554,N_12341);
nor U14262 (N_14262,N_13923,N_13609);
xnor U14263 (N_14263,N_12872,N_12839);
nor U14264 (N_14264,N_13438,N_13630);
and U14265 (N_14265,N_13826,N_13598);
nor U14266 (N_14266,N_13832,N_13467);
xor U14267 (N_14267,N_13881,N_13971);
nor U14268 (N_14268,N_13386,N_12457);
nor U14269 (N_14269,N_12185,N_13796);
or U14270 (N_14270,N_12152,N_12561);
or U14271 (N_14271,N_13772,N_12354);
and U14272 (N_14272,N_12794,N_13492);
xnor U14273 (N_14273,N_13560,N_13163);
xnor U14274 (N_14274,N_12049,N_12174);
or U14275 (N_14275,N_12582,N_12205);
nand U14276 (N_14276,N_12320,N_12990);
nand U14277 (N_14277,N_12905,N_12132);
nor U14278 (N_14278,N_13347,N_13015);
xnor U14279 (N_14279,N_13231,N_13785);
xor U14280 (N_14280,N_12827,N_13731);
and U14281 (N_14281,N_13097,N_13988);
and U14282 (N_14282,N_12727,N_13206);
or U14283 (N_14283,N_12476,N_12208);
and U14284 (N_14284,N_12746,N_13017);
xnor U14285 (N_14285,N_13140,N_12356);
nand U14286 (N_14286,N_12445,N_13587);
nor U14287 (N_14287,N_13311,N_13333);
xor U14288 (N_14288,N_13753,N_13109);
and U14289 (N_14289,N_13885,N_13874);
and U14290 (N_14290,N_13935,N_13850);
xor U14291 (N_14291,N_12545,N_13283);
nand U14292 (N_14292,N_12690,N_12623);
xnor U14293 (N_14293,N_12171,N_13688);
and U14294 (N_14294,N_13046,N_13914);
or U14295 (N_14295,N_13639,N_13638);
or U14296 (N_14296,N_12418,N_13352);
nand U14297 (N_14297,N_13450,N_12643);
xor U14298 (N_14298,N_13012,N_13593);
and U14299 (N_14299,N_12728,N_12429);
xor U14300 (N_14300,N_12441,N_13516);
or U14301 (N_14301,N_13312,N_12558);
or U14302 (N_14302,N_12337,N_13823);
xor U14303 (N_14303,N_12680,N_13852);
and U14304 (N_14304,N_13791,N_13207);
nand U14305 (N_14305,N_12769,N_13558);
nand U14306 (N_14306,N_13047,N_12659);
xnor U14307 (N_14307,N_13967,N_12335);
nand U14308 (N_14308,N_12482,N_13736);
xor U14309 (N_14309,N_13836,N_13681);
xnor U14310 (N_14310,N_13236,N_12111);
nor U14311 (N_14311,N_12961,N_12238);
nor U14312 (N_14312,N_13430,N_13135);
or U14313 (N_14313,N_13631,N_12962);
or U14314 (N_14314,N_12107,N_13809);
or U14315 (N_14315,N_13351,N_13563);
and U14316 (N_14316,N_13364,N_12523);
and U14317 (N_14317,N_13979,N_13872);
xnor U14318 (N_14318,N_12483,N_13117);
and U14319 (N_14319,N_13010,N_13362);
and U14320 (N_14320,N_13907,N_13799);
and U14321 (N_14321,N_12036,N_12569);
and U14322 (N_14322,N_12309,N_13118);
or U14323 (N_14323,N_13629,N_13662);
nand U14324 (N_14324,N_13645,N_12034);
nand U14325 (N_14325,N_13044,N_12677);
xnor U14326 (N_14326,N_13459,N_12857);
nor U14327 (N_14327,N_13072,N_12653);
or U14328 (N_14328,N_13839,N_13573);
and U14329 (N_14329,N_13624,N_13580);
xnor U14330 (N_14330,N_12447,N_12413);
and U14331 (N_14331,N_13328,N_13575);
and U14332 (N_14332,N_12066,N_12715);
nor U14333 (N_14333,N_13683,N_13337);
or U14334 (N_14334,N_13588,N_12566);
or U14335 (N_14335,N_12675,N_13743);
nand U14336 (N_14336,N_12840,N_13761);
xor U14337 (N_14337,N_13528,N_12131);
and U14338 (N_14338,N_13310,N_13970);
nor U14339 (N_14339,N_13797,N_12465);
nor U14340 (N_14340,N_13781,N_12984);
nor U14341 (N_14341,N_12378,N_13847);
and U14342 (N_14342,N_12665,N_12513);
and U14343 (N_14343,N_13145,N_13498);
nand U14344 (N_14344,N_13605,N_12547);
and U14345 (N_14345,N_12996,N_13089);
nor U14346 (N_14346,N_12071,N_13953);
nand U14347 (N_14347,N_13226,N_13255);
nor U14348 (N_14348,N_13776,N_13096);
and U14349 (N_14349,N_12925,N_12325);
xnor U14350 (N_14350,N_12194,N_13287);
xor U14351 (N_14351,N_13308,N_13005);
xnor U14352 (N_14352,N_12604,N_13913);
nand U14353 (N_14353,N_12427,N_13699);
nand U14354 (N_14354,N_13860,N_13900);
xnor U14355 (N_14355,N_13951,N_12367);
or U14356 (N_14356,N_13671,N_12557);
and U14357 (N_14357,N_13266,N_12500);
nor U14358 (N_14358,N_12162,N_13004);
nand U14359 (N_14359,N_13291,N_12041);
nand U14360 (N_14360,N_12786,N_12852);
or U14361 (N_14361,N_12748,N_13959);
nor U14362 (N_14362,N_12032,N_13003);
or U14363 (N_14363,N_13454,N_13263);
or U14364 (N_14364,N_13829,N_13028);
nor U14365 (N_14365,N_12656,N_13247);
or U14366 (N_14366,N_12383,N_12651);
and U14367 (N_14367,N_13661,N_12078);
nand U14368 (N_14368,N_12571,N_12620);
xnor U14369 (N_14369,N_12343,N_12744);
and U14370 (N_14370,N_12009,N_12914);
and U14371 (N_14371,N_13136,N_12601);
nand U14372 (N_14372,N_13460,N_13802);
nor U14373 (N_14373,N_13779,N_13719);
nor U14374 (N_14374,N_13345,N_12768);
nand U14375 (N_14375,N_12488,N_13360);
or U14376 (N_14376,N_12538,N_13611);
and U14377 (N_14377,N_13654,N_13817);
nor U14378 (N_14378,N_13548,N_12283);
nand U14379 (N_14379,N_13155,N_12747);
xnor U14380 (N_14380,N_12527,N_13727);
and U14381 (N_14381,N_13318,N_12756);
nand U14382 (N_14382,N_13405,N_13294);
nand U14383 (N_14383,N_13669,N_13828);
xnor U14384 (N_14384,N_12778,N_12376);
and U14385 (N_14385,N_13532,N_12307);
and U14386 (N_14386,N_13819,N_12594);
nor U14387 (N_14387,N_12432,N_12033);
or U14388 (N_14388,N_13052,N_12493);
nor U14389 (N_14389,N_13307,N_13658);
or U14390 (N_14390,N_12743,N_13399);
xor U14391 (N_14391,N_13216,N_12924);
or U14392 (N_14392,N_13144,N_12671);
or U14393 (N_14393,N_13884,N_12779);
or U14394 (N_14394,N_13449,N_13361);
xnor U14395 (N_14395,N_13421,N_13152);
nand U14396 (N_14396,N_13777,N_13070);
or U14397 (N_14397,N_13553,N_12097);
nand U14398 (N_14398,N_12548,N_12070);
and U14399 (N_14399,N_12644,N_13463);
nor U14400 (N_14400,N_12689,N_12241);
nor U14401 (N_14401,N_12845,N_12890);
and U14402 (N_14402,N_13132,N_12058);
or U14403 (N_14403,N_13768,N_12075);
nand U14404 (N_14404,N_12932,N_13868);
or U14405 (N_14405,N_13643,N_12247);
xnor U14406 (N_14406,N_12164,N_12864);
xor U14407 (N_14407,N_12411,N_12387);
xnor U14408 (N_14408,N_12935,N_12867);
nor U14409 (N_14409,N_13203,N_12179);
and U14410 (N_14410,N_13178,N_12694);
nand U14411 (N_14411,N_12738,N_13475);
nor U14412 (N_14412,N_13921,N_13627);
nor U14413 (N_14413,N_12532,N_12831);
and U14414 (N_14414,N_13389,N_12544);
xnor U14415 (N_14415,N_12392,N_13420);
xor U14416 (N_14416,N_13728,N_12552);
xor U14417 (N_14417,N_13936,N_13756);
and U14418 (N_14418,N_13087,N_13018);
or U14419 (N_14419,N_12921,N_13928);
or U14420 (N_14420,N_12397,N_12947);
and U14421 (N_14421,N_13517,N_13040);
nand U14422 (N_14422,N_13717,N_13268);
nand U14423 (N_14423,N_12796,N_13325);
nor U14424 (N_14424,N_12414,N_12621);
nand U14425 (N_14425,N_13177,N_13156);
and U14426 (N_14426,N_12167,N_13843);
and U14427 (N_14427,N_13043,N_13383);
and U14428 (N_14428,N_13001,N_13148);
nand U14429 (N_14429,N_13762,N_12469);
nand U14430 (N_14430,N_13747,N_12780);
xor U14431 (N_14431,N_13541,N_12043);
and U14432 (N_14432,N_13141,N_13088);
xnor U14433 (N_14433,N_13945,N_13714);
xnor U14434 (N_14434,N_13339,N_12130);
or U14435 (N_14435,N_12828,N_13664);
xnor U14436 (N_14436,N_13716,N_13876);
nand U14437 (N_14437,N_13737,N_13190);
nand U14438 (N_14438,N_13869,N_12382);
nand U14439 (N_14439,N_13422,N_12114);
and U14440 (N_14440,N_13586,N_13767);
nor U14441 (N_14441,N_12849,N_12253);
nand U14442 (N_14442,N_12138,N_12274);
or U14443 (N_14443,N_13164,N_13937);
or U14444 (N_14444,N_13100,N_13298);
or U14445 (N_14445,N_12988,N_12322);
and U14446 (N_14446,N_13758,N_12385);
and U14447 (N_14447,N_13410,N_13725);
nand U14448 (N_14448,N_13966,N_12393);
or U14449 (N_14449,N_13509,N_13210);
nor U14450 (N_14450,N_12492,N_13194);
and U14451 (N_14451,N_13218,N_12127);
and U14452 (N_14452,N_12310,N_12622);
nor U14453 (N_14453,N_13578,N_13569);
nor U14454 (N_14454,N_12153,N_12093);
nand U14455 (N_14455,N_12317,N_12178);
nand U14456 (N_14456,N_12726,N_13076);
nand U14457 (N_14457,N_13822,N_12332);
nor U14458 (N_14458,N_12110,N_12504);
nor U14459 (N_14459,N_12528,N_13623);
and U14460 (N_14460,N_13529,N_13614);
xnor U14461 (N_14461,N_13371,N_13917);
nor U14462 (N_14462,N_13748,N_13999);
and U14463 (N_14463,N_12444,N_12321);
nor U14464 (N_14464,N_13775,N_12301);
nor U14465 (N_14465,N_13284,N_12261);
or U14466 (N_14466,N_12664,N_12076);
nand U14467 (N_14467,N_13470,N_12841);
nand U14468 (N_14468,N_12772,N_13081);
xnor U14469 (N_14469,N_12686,N_13806);
or U14470 (N_14470,N_12428,N_12446);
nor U14471 (N_14471,N_12883,N_12461);
nand U14472 (N_14472,N_13659,N_13128);
xor U14473 (N_14473,N_12904,N_12412);
nor U14474 (N_14474,N_12008,N_12511);
nand U14475 (N_14475,N_12073,N_12901);
and U14476 (N_14476,N_12135,N_13732);
xor U14477 (N_14477,N_12139,N_12369);
nand U14478 (N_14478,N_12436,N_12239);
xnor U14479 (N_14479,N_12014,N_13235);
nand U14480 (N_14480,N_12843,N_12931);
and U14481 (N_14481,N_12105,N_12521);
and U14482 (N_14482,N_13875,N_13840);
nor U14483 (N_14483,N_12405,N_12958);
xnor U14484 (N_14484,N_12474,N_12525);
and U14485 (N_14485,N_12192,N_12451);
or U14486 (N_14486,N_12616,N_13007);
nor U14487 (N_14487,N_12877,N_12001);
nand U14488 (N_14488,N_13392,N_13502);
and U14489 (N_14489,N_13595,N_13985);
xor U14490 (N_14490,N_13038,N_12276);
and U14491 (N_14491,N_12605,N_12285);
or U14492 (N_14492,N_13094,N_13265);
and U14493 (N_14493,N_12030,N_12421);
and U14494 (N_14494,N_13056,N_12198);
nand U14495 (N_14495,N_12516,N_13505);
or U14496 (N_14496,N_12264,N_13209);
xnor U14497 (N_14497,N_12564,N_12662);
nor U14498 (N_14498,N_12117,N_13507);
nor U14499 (N_14499,N_13991,N_12477);
or U14500 (N_14500,N_13179,N_12292);
nand U14501 (N_14501,N_13804,N_13675);
or U14502 (N_14502,N_12266,N_12807);
and U14503 (N_14503,N_12520,N_12969);
or U14504 (N_14504,N_13949,N_13896);
nand U14505 (N_14505,N_12898,N_13530);
xor U14506 (N_14506,N_12318,N_13711);
xor U14507 (N_14507,N_12989,N_12949);
or U14508 (N_14508,N_13491,N_12063);
or U14509 (N_14509,N_12280,N_12210);
and U14510 (N_14510,N_12560,N_13406);
nand U14511 (N_14511,N_13327,N_12338);
or U14512 (N_14512,N_12183,N_12161);
nor U14513 (N_14513,N_13621,N_12606);
nor U14514 (N_14514,N_13429,N_12195);
nor U14515 (N_14515,N_12933,N_12895);
nand U14516 (N_14516,N_13300,N_12122);
xnor U14517 (N_14517,N_13130,N_13689);
and U14518 (N_14518,N_13651,N_13811);
xor U14519 (N_14519,N_12475,N_12976);
xnor U14520 (N_14520,N_12994,N_13077);
nor U14521 (N_14521,N_13407,N_12838);
nor U14522 (N_14522,N_13027,N_13570);
nand U14523 (N_14523,N_13175,N_13846);
and U14524 (N_14524,N_12083,N_12723);
and U14525 (N_14525,N_13244,N_12342);
nor U14526 (N_14526,N_12349,N_12284);
or U14527 (N_14527,N_12175,N_12584);
xnor U14528 (N_14528,N_13808,N_12944);
and U14529 (N_14529,N_12718,N_12173);
nand U14530 (N_14530,N_13261,N_13165);
or U14531 (N_14531,N_13956,N_13687);
nand U14532 (N_14532,N_13431,N_13411);
xnor U14533 (N_14533,N_12494,N_12943);
or U14534 (N_14534,N_12509,N_12518);
and U14535 (N_14535,N_13908,N_12954);
xor U14536 (N_14536,N_13272,N_13314);
nand U14537 (N_14537,N_12902,N_13646);
or U14538 (N_14538,N_13707,N_13597);
xnor U14539 (N_14539,N_12641,N_13798);
nand U14540 (N_14540,N_12228,N_13983);
and U14541 (N_14541,N_12082,N_12234);
and U14542 (N_14542,N_12355,N_12067);
and U14543 (N_14543,N_13984,N_13024);
xor U14544 (N_14544,N_12531,N_12787);
and U14545 (N_14545,N_13608,N_13890);
nor U14546 (N_14546,N_13856,N_13506);
nor U14547 (N_14547,N_13564,N_13600);
xor U14548 (N_14548,N_13650,N_13655);
xnor U14549 (N_14549,N_13489,N_13968);
xnor U14550 (N_14550,N_12207,N_13254);
nor U14551 (N_14551,N_13330,N_12777);
or U14552 (N_14552,N_12978,N_12749);
nand U14553 (N_14553,N_13982,N_12352);
xnor U14554 (N_14554,N_12995,N_12458);
nor U14555 (N_14555,N_13354,N_12257);
xor U14556 (N_14556,N_13153,N_13301);
and U14557 (N_14557,N_12765,N_12655);
nand U14558 (N_14558,N_12633,N_12681);
xnor U14559 (N_14559,N_13590,N_13710);
nor U14560 (N_14560,N_13065,N_13281);
or U14561 (N_14561,N_13116,N_13897);
xor U14562 (N_14562,N_12866,N_12454);
or U14563 (N_14563,N_13901,N_12751);
and U14564 (N_14564,N_12080,N_13086);
nor U14565 (N_14565,N_12024,N_12964);
nand U14566 (N_14566,N_13579,N_12023);
or U14567 (N_14567,N_13482,N_12425);
nand U14568 (N_14568,N_12224,N_12391);
or U14569 (N_14569,N_13519,N_12941);
nand U14570 (N_14570,N_13841,N_12775);
nand U14571 (N_14571,N_13167,N_12567);
and U14572 (N_14572,N_12599,N_12002);
or U14573 (N_14573,N_13336,N_12939);
xor U14574 (N_14574,N_13706,N_12021);
and U14575 (N_14575,N_13686,N_13855);
or U14576 (N_14576,N_12917,N_12294);
nand U14577 (N_14577,N_13037,N_12697);
xor U14578 (N_14578,N_12816,N_12589);
nand U14579 (N_14579,N_13863,N_13497);
nand U14580 (N_14580,N_13341,N_12072);
or U14581 (N_14581,N_12235,N_12219);
nor U14582 (N_14582,N_13020,N_12443);
or U14583 (N_14583,N_12015,N_13693);
or U14584 (N_14584,N_12855,N_12782);
nand U14585 (N_14585,N_13104,N_13323);
and U14586 (N_14586,N_13241,N_12340);
nor U14587 (N_14587,N_13807,N_12448);
and U14588 (N_14588,N_12499,N_13955);
or U14589 (N_14589,N_13197,N_12380);
or U14590 (N_14590,N_12426,N_13657);
xnor U14591 (N_14591,N_12913,N_12467);
nand U14592 (N_14592,N_12217,N_12757);
and U14593 (N_14593,N_13909,N_12613);
and U14594 (N_14594,N_12098,N_12631);
and U14595 (N_14595,N_12053,N_13562);
nor U14596 (N_14596,N_13927,N_12663);
nor U14597 (N_14597,N_13730,N_12577);
xor U14598 (N_14598,N_13198,N_13538);
or U14599 (N_14599,N_12103,N_13143);
xor U14600 (N_14600,N_12156,N_12801);
xor U14601 (N_14601,N_13787,N_12216);
nand U14602 (N_14602,N_13939,N_12199);
xnor U14603 (N_14603,N_12842,N_13296);
and U14604 (N_14604,N_13678,N_13480);
xnor U14605 (N_14605,N_13942,N_12647);
or U14606 (N_14606,N_12576,N_13282);
nor U14607 (N_14607,N_13363,N_13262);
and U14608 (N_14608,N_13895,N_13996);
or U14609 (N_14609,N_12741,N_13276);
or U14610 (N_14610,N_12529,N_12218);
nand U14611 (N_14611,N_13757,N_12419);
nor U14612 (N_14612,N_13545,N_12133);
xor U14613 (N_14613,N_12048,N_12878);
xnor U14614 (N_14614,N_12282,N_13684);
xor U14615 (N_14615,N_12118,N_13814);
xor U14616 (N_14616,N_12830,N_13534);
and U14617 (N_14617,N_12243,N_12829);
nand U14618 (N_14618,N_13919,N_13601);
and U14619 (N_14619,N_13964,N_12602);
or U14620 (N_14620,N_12395,N_13490);
nor U14621 (N_14621,N_12916,N_12172);
or U14622 (N_14622,N_13510,N_12977);
nand U14623 (N_14623,N_12371,N_12776);
and U14624 (N_14624,N_12543,N_12042);
nand U14625 (N_14625,N_13376,N_12936);
xor U14626 (N_14626,N_13769,N_13474);
xor U14627 (N_14627,N_13782,N_13061);
xor U14628 (N_14628,N_12256,N_13925);
or U14629 (N_14629,N_13378,N_12624);
nand U14630 (N_14630,N_13557,N_13062);
nor U14631 (N_14631,N_12588,N_13286);
nor U14632 (N_14632,N_12654,N_12848);
xor U14633 (N_14633,N_13652,N_12795);
and U14634 (N_14634,N_12288,N_13522);
xnor U14635 (N_14635,N_12825,N_13121);
nand U14636 (N_14636,N_13715,N_12574);
or U14637 (N_14637,N_12423,N_12896);
xor U14638 (N_14638,N_12682,N_13511);
and U14639 (N_14639,N_12884,N_13574);
xnor U14640 (N_14640,N_12579,N_12370);
xor U14641 (N_14641,N_12634,N_13439);
nor U14642 (N_14642,N_12453,N_12290);
xor U14643 (N_14643,N_12565,N_12981);
xor U14644 (N_14644,N_13306,N_13640);
nand U14645 (N_14645,N_12963,N_12115);
nand U14646 (N_14646,N_12535,N_13075);
xnor U14647 (N_14647,N_13485,N_12244);
nand U14648 (N_14648,N_12222,N_13858);
or U14649 (N_14649,N_13435,N_13212);
or U14650 (N_14650,N_13150,N_13161);
or U14651 (N_14651,N_12305,N_12632);
nand U14652 (N_14652,N_12676,N_13054);
or U14653 (N_14653,N_13703,N_12732);
xnor U14654 (N_14654,N_13002,N_12617);
nor U14655 (N_14655,N_13903,N_13882);
nor U14656 (N_14656,N_13171,N_13697);
or U14657 (N_14657,N_13384,N_13338);
and U14658 (N_14658,N_13789,N_13396);
nor U14659 (N_14659,N_12039,N_13346);
and U14660 (N_14660,N_12191,N_12271);
and U14661 (N_14661,N_12707,N_13734);
nand U14662 (N_14662,N_13215,N_13403);
or U14663 (N_14663,N_13269,N_12206);
nand U14664 (N_14664,N_12246,N_12311);
xor U14665 (N_14665,N_12854,N_13487);
xnor U14666 (N_14666,N_13713,N_12245);
xnor U14667 (N_14667,N_12143,N_12900);
or U14668 (N_14668,N_13851,N_12077);
or U14669 (N_14669,N_13205,N_13068);
xor U14670 (N_14670,N_13812,N_13526);
and U14671 (N_14671,N_13032,N_13871);
nor U14672 (N_14672,N_12940,N_12495);
nand U14673 (N_14673,N_12126,N_12851);
or U14674 (N_14674,N_12700,N_12250);
xor U14675 (N_14675,N_12381,N_12357);
xor U14676 (N_14676,N_13067,N_12480);
nand U14677 (N_14677,N_12487,N_13057);
nand U14678 (N_14678,N_12251,N_13437);
nor U14679 (N_14679,N_13887,N_13577);
and U14680 (N_14680,N_13486,N_13965);
or U14681 (N_14681,N_12575,N_12197);
and U14682 (N_14682,N_12974,N_13200);
xor U14683 (N_14683,N_13138,N_12229);
or U14684 (N_14684,N_12424,N_13234);
and U14685 (N_14685,N_12360,N_13993);
nor U14686 (N_14686,N_12915,N_13700);
and U14687 (N_14687,N_12315,N_12459);
and U14688 (N_14688,N_12514,N_13603);
xor U14689 (N_14689,N_13960,N_12314);
xnor U14690 (N_14690,N_13838,N_13477);
nand U14691 (N_14691,N_13110,N_13014);
xor U14692 (N_14692,N_13898,N_13862);
nor U14693 (N_14693,N_12619,N_13270);
nor U14694 (N_14694,N_13594,N_13783);
or U14695 (N_14695,N_12695,N_13576);
and U14696 (N_14696,N_12903,N_13166);
nand U14697 (N_14697,N_12471,N_13742);
nand U14698 (N_14698,N_12581,N_13350);
nor U14699 (N_14699,N_12764,N_13091);
xnor U14700 (N_14700,N_13744,N_12464);
nand U14701 (N_14701,N_13021,N_12180);
or U14702 (N_14702,N_13930,N_12125);
and U14703 (N_14703,N_12800,N_12767);
or U14704 (N_14704,N_13674,N_12711);
or U14705 (N_14705,N_12708,N_12615);
nor U14706 (N_14706,N_13864,N_12018);
or U14707 (N_14707,N_13679,N_13108);
or U14708 (N_14708,N_12955,N_13954);
nand U14709 (N_14709,N_12237,N_13612);
xor U14710 (N_14710,N_13877,N_12888);
nor U14711 (N_14711,N_12573,N_12788);
xor U14712 (N_14712,N_12945,N_12894);
nor U14713 (N_14713,N_12702,N_13257);
xnor U14714 (N_14714,N_13188,N_13457);
nor U14715 (N_14715,N_13637,N_13326);
nand U14716 (N_14716,N_12262,N_12003);
and U14717 (N_14717,N_12439,N_13820);
nor U14718 (N_14718,N_12373,N_13064);
and U14719 (N_14719,N_13211,N_12496);
nand U14720 (N_14720,N_13647,N_12992);
nor U14721 (N_14721,N_12300,N_12249);
nand U14722 (N_14722,N_13267,N_12610);
nand U14723 (N_14723,N_13317,N_13854);
and U14724 (N_14724,N_13377,N_12260);
xor U14725 (N_14725,N_13622,N_12906);
nor U14726 (N_14726,N_12612,N_13124);
nor U14727 (N_14727,N_13444,N_13232);
xor U14728 (N_14728,N_12095,N_13183);
nor U14729 (N_14729,N_13997,N_12362);
or U14730 (N_14730,N_13663,N_12629);
xor U14731 (N_14731,N_12636,N_12648);
or U14732 (N_14732,N_13501,N_12879);
or U14733 (N_14733,N_12553,N_13888);
nand U14734 (N_14734,N_12220,N_12255);
xor U14735 (N_14735,N_12798,N_13090);
and U14736 (N_14736,N_12815,N_13746);
and U14737 (N_14737,N_12853,N_12324);
nand U14738 (N_14738,N_13013,N_12639);
xor U14739 (N_14739,N_12937,N_12938);
or U14740 (N_14740,N_13821,N_12683);
xor U14741 (N_14741,N_12563,N_12733);
and U14742 (N_14742,N_13042,N_13981);
nand U14743 (N_14743,N_12056,N_13961);
or U14744 (N_14744,N_13026,N_12064);
nand U14745 (N_14745,N_12522,N_12865);
xnor U14746 (N_14746,N_13759,N_13066);
or U14747 (N_14747,N_13950,N_13274);
or U14748 (N_14748,N_12519,N_13495);
nand U14749 (N_14749,N_12763,N_13181);
nor U14750 (N_14750,N_12844,N_13192);
xor U14751 (N_14751,N_13738,N_12204);
nand U14752 (N_14752,N_12472,N_12967);
and U14753 (N_14753,N_13413,N_12272);
nand U14754 (N_14754,N_12334,N_12510);
nand U14755 (N_14755,N_13633,N_12590);
nor U14756 (N_14756,N_13425,N_13332);
nand U14757 (N_14757,N_12269,N_12379);
or U14758 (N_14758,N_13424,N_12060);
and U14759 (N_14759,N_12134,N_13115);
nor U14760 (N_14760,N_12736,N_13729);
and U14761 (N_14761,N_12821,N_12351);
or U14762 (N_14762,N_12669,N_13133);
xnor U14763 (N_14763,N_12986,N_13356);
nor U14764 (N_14764,N_12637,N_12402);
and U14765 (N_14765,N_13585,N_13933);
nor U14766 (N_14766,N_12159,N_12157);
xnor U14767 (N_14767,N_13619,N_13830);
nor U14768 (N_14768,N_13185,N_12147);
or U14769 (N_14769,N_12037,N_13404);
or U14770 (N_14770,N_13488,N_12930);
nor U14771 (N_14771,N_13543,N_13316);
or U14772 (N_14772,N_13006,N_13599);
and U14773 (N_14773,N_13931,N_12946);
nor U14774 (N_14774,N_13349,N_13099);
nand U14775 (N_14775,N_12242,N_12713);
nor U14776 (N_14776,N_12390,N_12919);
or U14777 (N_14777,N_13792,N_13414);
nand U14778 (N_14778,N_12491,N_13891);
nor U14779 (N_14779,N_12957,N_12817);
nor U14780 (N_14780,N_12312,N_13571);
or U14781 (N_14781,N_13685,N_12802);
or U14782 (N_14782,N_12396,N_12555);
xor U14783 (N_14783,N_13381,N_13008);
nor U14784 (N_14784,N_12858,N_12148);
or U14785 (N_14785,N_12020,N_12897);
and U14786 (N_14786,N_12814,N_13271);
xnor U14787 (N_14787,N_13483,N_13285);
nand U14788 (N_14788,N_12596,N_13370);
xnor U14789 (N_14789,N_12306,N_13125);
nand U14790 (N_14790,N_13972,N_13473);
nor U14791 (N_14791,N_13827,N_12592);
and U14792 (N_14792,N_13478,N_13041);
xor U14793 (N_14793,N_12168,N_13741);
nand U14794 (N_14794,N_13322,N_13995);
nand U14795 (N_14795,N_13515,N_12267);
and U14796 (N_14796,N_12712,N_13080);
nor U14797 (N_14797,N_13607,N_12783);
nand U14798 (N_14798,N_12773,N_12022);
nor U14799 (N_14799,N_13801,N_13114);
or U14800 (N_14800,N_12087,N_13628);
nand U14801 (N_14801,N_13540,N_12019);
and U14802 (N_14802,N_13225,N_13496);
nor U14803 (N_14803,N_13844,N_13947);
or U14804 (N_14804,N_12031,N_12038);
nor U14805 (N_14805,N_13904,N_13400);
nand U14806 (N_14806,N_13329,N_13112);
and U14807 (N_14807,N_12722,N_13191);
and U14808 (N_14808,N_13754,N_12293);
xnor U14809 (N_14809,N_13892,N_13551);
nor U14810 (N_14810,N_13958,N_13313);
nand U14811 (N_14811,N_12140,N_13641);
nor U14812 (N_14812,N_12701,N_13990);
nand U14813 (N_14813,N_13924,N_12415);
nor U14814 (N_14814,N_12017,N_12972);
nor U14815 (N_14815,N_12090,N_13780);
nand U14816 (N_14816,N_13379,N_13358);
or U14817 (N_14817,N_12953,N_13369);
and U14818 (N_14818,N_13246,N_13184);
nor U14819 (N_14819,N_13402,N_13162);
nand U14820 (N_14820,N_12693,N_12006);
and U14821 (N_14821,N_12998,N_13583);
nand U14822 (N_14822,N_12081,N_12455);
nor U14823 (N_14823,N_12515,N_12666);
nand U14824 (N_14824,N_12406,N_13193);
and U14825 (N_14825,N_13591,N_12928);
nor U14826 (N_14826,N_13157,N_12109);
xor U14827 (N_14827,N_13248,N_12699);
and U14828 (N_14828,N_13461,N_12600);
and U14829 (N_14829,N_13443,N_12155);
nor U14830 (N_14830,N_12365,N_12862);
nor U14831 (N_14831,N_12258,N_13648);
xnor U14832 (N_14832,N_13253,N_12136);
nand U14833 (N_14833,N_12983,N_12703);
xnor U14834 (N_14834,N_12013,N_13912);
xnor U14835 (N_14835,N_13423,N_12539);
or U14836 (N_14836,N_13199,N_13760);
and U14837 (N_14837,N_12214,N_12086);
nand U14838 (N_14838,N_12587,N_12108);
nand U14839 (N_14839,N_12120,N_12730);
and U14840 (N_14840,N_13620,N_12820);
or U14841 (N_14841,N_13805,N_12658);
nand U14842 (N_14842,N_12766,N_13134);
nand U14843 (N_14843,N_13251,N_13539);
xor U14844 (N_14844,N_12170,N_13053);
and U14845 (N_14845,N_12591,N_13694);
nor U14846 (N_14846,N_12478,N_13845);
or U14847 (N_14847,N_13589,N_13331);
nor U14848 (N_14848,N_12761,N_13297);
nor U14849 (N_14849,N_13665,N_13503);
and U14850 (N_14850,N_13500,N_12486);
or U14851 (N_14851,N_13712,N_12704);
nor U14852 (N_14852,N_13813,N_13962);
and U14853 (N_14853,N_13158,N_12880);
or U14854 (N_14854,N_12401,N_12485);
and U14855 (N_14855,N_13918,N_12403);
or U14856 (N_14856,N_12069,N_12254);
nor U14857 (N_14857,N_13227,N_12050);
xor U14858 (N_14858,N_12859,N_12526);
nor U14859 (N_14859,N_13214,N_12230);
nand U14860 (N_14860,N_12470,N_13546);
and U14861 (N_14861,N_13702,N_12698);
nand U14862 (N_14862,N_13292,N_13213);
nor U14863 (N_14863,N_13063,N_12129);
and U14864 (N_14864,N_13471,N_13093);
xor U14865 (N_14865,N_13085,N_13974);
nor U14866 (N_14866,N_13567,N_12201);
nor U14867 (N_14867,N_12846,N_12752);
nor U14868 (N_14868,N_13550,N_12102);
and U14869 (N_14869,N_13720,N_13105);
or U14870 (N_14870,N_13466,N_13508);
and U14871 (N_14871,N_12826,N_13030);
or U14872 (N_14872,N_12215,N_12128);
xnor U14873 (N_14873,N_13113,N_13170);
nor U14874 (N_14874,N_13472,N_13987);
and U14875 (N_14875,N_12193,N_13393);
xnor U14876 (N_14876,N_13523,N_12252);
and U14877 (N_14877,N_13446,N_12211);
nand U14878 (N_14878,N_13889,N_13372);
nor U14879 (N_14879,N_13220,N_13559);
nor U14880 (N_14880,N_12811,N_13084);
and U14881 (N_14881,N_12929,N_12863);
nor U14882 (N_14882,N_13572,N_13677);
or U14883 (N_14883,N_13566,N_13151);
and U14884 (N_14884,N_13154,N_12313);
nand U14885 (N_14885,N_12333,N_13048);
or U14886 (N_14886,N_12813,N_12101);
nor U14887 (N_14887,N_12687,N_12542);
xnor U14888 (N_14888,N_12710,N_13082);
and U14889 (N_14889,N_12533,N_12059);
nand U14890 (N_14890,N_12585,N_13976);
or U14891 (N_14891,N_12089,N_12123);
or U14892 (N_14892,N_12792,N_12642);
or U14893 (N_14893,N_13941,N_12549);
nor U14894 (N_14894,N_13778,N_12026);
and U14895 (N_14895,N_13343,N_13419);
nor U14896 (N_14896,N_13304,N_13451);
nand U14897 (N_14897,N_13230,N_13834);
or U14898 (N_14898,N_12607,N_12085);
nand U14899 (N_14899,N_13279,N_12735);
nor U14900 (N_14900,N_13494,N_13512);
or U14901 (N_14901,N_12824,N_12270);
xnor U14902 (N_14902,N_12638,N_13555);
nor U14903 (N_14903,N_12806,N_13722);
nand U14904 (N_14904,N_12721,N_13831);
and U14905 (N_14905,N_12559,N_13818);
xor U14906 (N_14906,N_13174,N_12891);
and U14907 (N_14907,N_12196,N_12359);
xnor U14908 (N_14908,N_12227,N_12869);
nand U14909 (N_14909,N_12119,N_12505);
nand U14910 (N_14910,N_12096,N_12578);
nor U14911 (N_14911,N_12498,N_12100);
xor U14912 (N_14912,N_12433,N_12980);
nor U14913 (N_14913,N_13861,N_13513);
or U14914 (N_14914,N_12407,N_12881);
and U14915 (N_14915,N_12873,N_13440);
nor U14916 (N_14916,N_12298,N_13201);
nand U14917 (N_14917,N_13309,N_13537);
nor U14918 (N_14918,N_13320,N_12044);
and U14919 (N_14919,N_12512,N_13374);
and U14920 (N_14920,N_13240,N_13408);
nor U14921 (N_14921,N_13098,N_12010);
xor U14922 (N_14922,N_12942,N_13131);
nor U14923 (N_14923,N_12530,N_13469);
xor U14924 (N_14924,N_12791,N_12212);
or U14925 (N_14925,N_12580,N_12737);
nand U14926 (N_14926,N_12506,N_12112);
or U14927 (N_14927,N_13103,N_13853);
xor U14928 (N_14928,N_13023,N_12016);
nand U14929 (N_14929,N_12336,N_12165);
or U14930 (N_14930,N_13857,N_12960);
nor U14931 (N_14931,N_13957,N_13355);
and U14932 (N_14932,N_13069,N_13442);
xnor U14933 (N_14933,N_12645,N_12753);
nand U14934 (N_14934,N_13321,N_13815);
nor U14935 (N_14935,N_12350,N_13476);
nor U14936 (N_14936,N_12047,N_13626);
nor U14937 (N_14937,N_13617,N_13434);
nor U14938 (N_14938,N_13696,N_12388);
or U14939 (N_14939,N_13773,N_13380);
nor U14940 (N_14940,N_13524,N_12562);
or U14941 (N_14941,N_12692,N_12759);
and U14942 (N_14942,N_12296,N_12295);
nor U14943 (N_14943,N_12330,N_13233);
or U14944 (N_14944,N_13810,N_13721);
nor U14945 (N_14945,N_12570,N_12979);
and U14946 (N_14946,N_13176,N_12674);
and U14947 (N_14947,N_12572,N_13000);
or U14948 (N_14948,N_13751,N_12029);
xor U14949 (N_14949,N_12818,N_12203);
xor U14950 (N_14950,N_12729,N_13766);
nand U14951 (N_14951,N_13755,N_12725);
nor U14952 (N_14952,N_12502,N_13397);
or U14953 (N_14953,N_12720,N_12770);
nor U14954 (N_14954,N_13428,N_12158);
or U14955 (N_14955,N_12190,N_13916);
or U14956 (N_14956,N_12627,N_13275);
nor U14957 (N_14957,N_13565,N_13544);
and U14958 (N_14958,N_12062,N_12993);
nand U14959 (N_14959,N_13618,N_12755);
nor U14960 (N_14960,N_12248,N_12149);
nor U14961 (N_14961,N_12434,N_12417);
nand U14962 (N_14962,N_12785,N_13859);
nor U14963 (N_14963,N_13670,N_12404);
xnor U14964 (N_14964,N_12927,N_12799);
or U14965 (N_14965,N_12985,N_12850);
or U14966 (N_14966,N_12027,N_13195);
nand U14967 (N_14967,N_12517,N_13963);
and U14968 (N_14968,N_12688,N_12046);
or U14969 (N_14969,N_12344,N_13447);
nor U14970 (N_14970,N_12438,N_12389);
or U14971 (N_14971,N_13481,N_12440);
or U14972 (N_14972,N_13387,N_12121);
nand U14973 (N_14973,N_13596,N_12847);
and U14974 (N_14974,N_12999,N_12789);
xor U14975 (N_14975,N_13391,N_12684);
xor U14976 (N_14976,N_12966,N_12466);
xnor U14977 (N_14977,N_13238,N_12327);
nor U14978 (N_14978,N_12181,N_13682);
nor U14979 (N_14979,N_13432,N_12277);
nor U14980 (N_14980,N_13531,N_12091);
nor U14981 (N_14981,N_13433,N_12377);
nand U14982 (N_14982,N_12045,N_13173);
xor U14983 (N_14983,N_13878,N_12348);
and U14984 (N_14984,N_13409,N_13427);
nand U14985 (N_14985,N_13228,N_13977);
or U14986 (N_14986,N_13680,N_13441);
xnor U14987 (N_14987,N_13305,N_13180);
nor U14988 (N_14988,N_13902,N_12011);
and U14989 (N_14989,N_12803,N_13202);
nor U14990 (N_14990,N_12065,N_12452);
or U14991 (N_14991,N_13740,N_12603);
and U14992 (N_14992,N_13365,N_13142);
nand U14993 (N_14993,N_13035,N_12289);
nand U14994 (N_14994,N_12760,N_13948);
nand U14995 (N_14995,N_12910,N_12705);
or U14996 (N_14996,N_12449,N_12997);
nor U14997 (N_14997,N_12358,N_12361);
nand U14998 (N_14998,N_12430,N_12353);
nand U14999 (N_14999,N_13221,N_12812);
nand U15000 (N_15000,N_12742,N_12015);
or U15001 (N_15001,N_12103,N_12183);
or U15002 (N_15002,N_12651,N_12634);
nand U15003 (N_15003,N_13146,N_12242);
nor U15004 (N_15004,N_13061,N_13525);
xnor U15005 (N_15005,N_13559,N_12546);
or U15006 (N_15006,N_13655,N_12155);
xor U15007 (N_15007,N_12087,N_12231);
or U15008 (N_15008,N_12684,N_13774);
nand U15009 (N_15009,N_13322,N_12989);
nand U15010 (N_15010,N_13512,N_12836);
nand U15011 (N_15011,N_12980,N_13955);
or U15012 (N_15012,N_13506,N_13901);
nor U15013 (N_15013,N_13314,N_13800);
nor U15014 (N_15014,N_13024,N_13019);
nand U15015 (N_15015,N_12274,N_13858);
or U15016 (N_15016,N_12236,N_12705);
or U15017 (N_15017,N_12633,N_12746);
xor U15018 (N_15018,N_13367,N_12361);
nor U15019 (N_15019,N_12259,N_13222);
or U15020 (N_15020,N_12933,N_13118);
xor U15021 (N_15021,N_12655,N_12411);
or U15022 (N_15022,N_12345,N_13088);
or U15023 (N_15023,N_13277,N_13239);
nand U15024 (N_15024,N_12784,N_13309);
nand U15025 (N_15025,N_13289,N_12874);
nand U15026 (N_15026,N_13918,N_13126);
or U15027 (N_15027,N_13787,N_13332);
nand U15028 (N_15028,N_12754,N_12382);
nand U15029 (N_15029,N_13999,N_13523);
xnor U15030 (N_15030,N_12332,N_13005);
nor U15031 (N_15031,N_12361,N_13765);
nor U15032 (N_15032,N_12697,N_13907);
nand U15033 (N_15033,N_12396,N_12535);
and U15034 (N_15034,N_12360,N_12781);
or U15035 (N_15035,N_12523,N_13167);
or U15036 (N_15036,N_13579,N_13003);
and U15037 (N_15037,N_12734,N_13924);
nor U15038 (N_15038,N_12794,N_13157);
nor U15039 (N_15039,N_13436,N_12815);
or U15040 (N_15040,N_13715,N_12767);
and U15041 (N_15041,N_13713,N_13028);
nor U15042 (N_15042,N_13308,N_13597);
nand U15043 (N_15043,N_12523,N_13404);
xor U15044 (N_15044,N_12202,N_13335);
or U15045 (N_15045,N_13163,N_13062);
xnor U15046 (N_15046,N_12108,N_12073);
and U15047 (N_15047,N_13008,N_13660);
or U15048 (N_15048,N_12847,N_12145);
or U15049 (N_15049,N_13099,N_13055);
nand U15050 (N_15050,N_12552,N_13021);
xnor U15051 (N_15051,N_13307,N_13362);
xnor U15052 (N_15052,N_12498,N_13265);
xnor U15053 (N_15053,N_13241,N_12920);
or U15054 (N_15054,N_13897,N_12264);
or U15055 (N_15055,N_12624,N_13974);
xor U15056 (N_15056,N_12555,N_12266);
and U15057 (N_15057,N_13901,N_12191);
xnor U15058 (N_15058,N_13323,N_12201);
or U15059 (N_15059,N_12446,N_12226);
and U15060 (N_15060,N_13823,N_13205);
and U15061 (N_15061,N_12939,N_12553);
nor U15062 (N_15062,N_12339,N_13081);
xor U15063 (N_15063,N_13190,N_12492);
xnor U15064 (N_15064,N_12129,N_12683);
or U15065 (N_15065,N_13157,N_13440);
and U15066 (N_15066,N_13449,N_12381);
and U15067 (N_15067,N_12119,N_13471);
or U15068 (N_15068,N_13534,N_12417);
nand U15069 (N_15069,N_13297,N_12232);
xnor U15070 (N_15070,N_13143,N_13648);
or U15071 (N_15071,N_13505,N_13229);
xnor U15072 (N_15072,N_12948,N_12435);
nor U15073 (N_15073,N_13816,N_13472);
or U15074 (N_15074,N_12369,N_12017);
or U15075 (N_15075,N_13483,N_12786);
nand U15076 (N_15076,N_13925,N_12281);
or U15077 (N_15077,N_12338,N_13079);
or U15078 (N_15078,N_13563,N_12279);
nand U15079 (N_15079,N_12086,N_13538);
or U15080 (N_15080,N_12231,N_13778);
and U15081 (N_15081,N_13689,N_13174);
xnor U15082 (N_15082,N_12884,N_12686);
xor U15083 (N_15083,N_12069,N_12628);
xnor U15084 (N_15084,N_13144,N_13849);
nand U15085 (N_15085,N_13280,N_13152);
xor U15086 (N_15086,N_13166,N_13861);
nor U15087 (N_15087,N_12539,N_12222);
or U15088 (N_15088,N_13708,N_13729);
xor U15089 (N_15089,N_12054,N_12983);
nand U15090 (N_15090,N_12934,N_12324);
nand U15091 (N_15091,N_13129,N_12108);
nor U15092 (N_15092,N_12276,N_12022);
nor U15093 (N_15093,N_12431,N_13681);
nand U15094 (N_15094,N_13122,N_12364);
nor U15095 (N_15095,N_12060,N_12917);
and U15096 (N_15096,N_12631,N_13428);
nand U15097 (N_15097,N_13983,N_12590);
xnor U15098 (N_15098,N_13735,N_13637);
and U15099 (N_15099,N_12404,N_12495);
or U15100 (N_15100,N_12087,N_13028);
or U15101 (N_15101,N_12328,N_12982);
xnor U15102 (N_15102,N_12183,N_13080);
nor U15103 (N_15103,N_13185,N_13615);
xor U15104 (N_15104,N_12839,N_12514);
or U15105 (N_15105,N_13050,N_13428);
xnor U15106 (N_15106,N_13024,N_12742);
xor U15107 (N_15107,N_13440,N_13529);
nand U15108 (N_15108,N_12049,N_13747);
or U15109 (N_15109,N_12807,N_13838);
xnor U15110 (N_15110,N_13519,N_13364);
nor U15111 (N_15111,N_12836,N_12984);
nand U15112 (N_15112,N_13043,N_13197);
nand U15113 (N_15113,N_13758,N_12698);
or U15114 (N_15114,N_13619,N_13467);
nand U15115 (N_15115,N_12555,N_13396);
nor U15116 (N_15116,N_12559,N_13058);
or U15117 (N_15117,N_13212,N_13104);
and U15118 (N_15118,N_12498,N_13099);
nor U15119 (N_15119,N_13698,N_12905);
xor U15120 (N_15120,N_13835,N_12204);
xor U15121 (N_15121,N_12035,N_12539);
nand U15122 (N_15122,N_12712,N_13472);
nor U15123 (N_15123,N_12425,N_12953);
and U15124 (N_15124,N_13957,N_12419);
or U15125 (N_15125,N_13955,N_13595);
or U15126 (N_15126,N_12478,N_13716);
nor U15127 (N_15127,N_13969,N_13950);
xnor U15128 (N_15128,N_12655,N_12246);
nand U15129 (N_15129,N_12915,N_13109);
xnor U15130 (N_15130,N_12781,N_13826);
nor U15131 (N_15131,N_12421,N_12914);
nor U15132 (N_15132,N_13601,N_13638);
xnor U15133 (N_15133,N_13391,N_13859);
nand U15134 (N_15134,N_13020,N_12558);
and U15135 (N_15135,N_13872,N_12017);
or U15136 (N_15136,N_13849,N_13435);
or U15137 (N_15137,N_13596,N_12971);
and U15138 (N_15138,N_12046,N_13086);
and U15139 (N_15139,N_13233,N_12637);
and U15140 (N_15140,N_13413,N_13696);
xnor U15141 (N_15141,N_13178,N_13482);
xor U15142 (N_15142,N_12066,N_12254);
nand U15143 (N_15143,N_12320,N_12647);
nor U15144 (N_15144,N_12739,N_13291);
or U15145 (N_15145,N_13218,N_13917);
or U15146 (N_15146,N_13161,N_13012);
nor U15147 (N_15147,N_13191,N_12788);
and U15148 (N_15148,N_13055,N_13291);
and U15149 (N_15149,N_12060,N_12063);
or U15150 (N_15150,N_12405,N_13586);
nor U15151 (N_15151,N_13219,N_13197);
xnor U15152 (N_15152,N_13456,N_13656);
xor U15153 (N_15153,N_12819,N_13982);
nand U15154 (N_15154,N_12900,N_13490);
nor U15155 (N_15155,N_12907,N_13968);
xor U15156 (N_15156,N_13113,N_12123);
or U15157 (N_15157,N_13386,N_12508);
nand U15158 (N_15158,N_12634,N_13795);
nor U15159 (N_15159,N_13345,N_12742);
and U15160 (N_15160,N_13852,N_12464);
or U15161 (N_15161,N_13836,N_13864);
nand U15162 (N_15162,N_13876,N_12420);
or U15163 (N_15163,N_13786,N_12863);
xnor U15164 (N_15164,N_12086,N_12030);
nor U15165 (N_15165,N_12261,N_13762);
or U15166 (N_15166,N_13845,N_12776);
xnor U15167 (N_15167,N_12391,N_13864);
nand U15168 (N_15168,N_13767,N_12067);
and U15169 (N_15169,N_13793,N_13896);
xnor U15170 (N_15170,N_12846,N_13703);
or U15171 (N_15171,N_12382,N_12951);
or U15172 (N_15172,N_13122,N_13632);
nand U15173 (N_15173,N_13594,N_12139);
nor U15174 (N_15174,N_12418,N_13716);
nor U15175 (N_15175,N_13910,N_13751);
nand U15176 (N_15176,N_12676,N_12888);
and U15177 (N_15177,N_12505,N_12456);
and U15178 (N_15178,N_13874,N_13099);
and U15179 (N_15179,N_13688,N_12084);
xnor U15180 (N_15180,N_12589,N_12962);
or U15181 (N_15181,N_12512,N_13207);
or U15182 (N_15182,N_13036,N_12953);
or U15183 (N_15183,N_12212,N_13609);
or U15184 (N_15184,N_13452,N_12057);
or U15185 (N_15185,N_12977,N_12376);
or U15186 (N_15186,N_13857,N_13451);
xnor U15187 (N_15187,N_12123,N_13557);
and U15188 (N_15188,N_13784,N_13981);
xnor U15189 (N_15189,N_13030,N_12508);
xnor U15190 (N_15190,N_12330,N_13589);
nor U15191 (N_15191,N_13121,N_13378);
or U15192 (N_15192,N_13548,N_13274);
nand U15193 (N_15193,N_12691,N_12777);
nand U15194 (N_15194,N_13195,N_12726);
or U15195 (N_15195,N_13444,N_12424);
xor U15196 (N_15196,N_13007,N_12162);
nand U15197 (N_15197,N_12382,N_13474);
and U15198 (N_15198,N_12147,N_12676);
xor U15199 (N_15199,N_12327,N_13608);
nor U15200 (N_15200,N_13858,N_13101);
xnor U15201 (N_15201,N_12038,N_13299);
or U15202 (N_15202,N_12844,N_12996);
and U15203 (N_15203,N_13612,N_13794);
nor U15204 (N_15204,N_13930,N_12996);
or U15205 (N_15205,N_12606,N_13354);
and U15206 (N_15206,N_13262,N_12636);
and U15207 (N_15207,N_12712,N_13714);
nor U15208 (N_15208,N_13350,N_12103);
xnor U15209 (N_15209,N_12345,N_12605);
xnor U15210 (N_15210,N_13113,N_13154);
nand U15211 (N_15211,N_12982,N_13344);
nor U15212 (N_15212,N_12086,N_12534);
nor U15213 (N_15213,N_12916,N_13588);
nand U15214 (N_15214,N_12047,N_13322);
nand U15215 (N_15215,N_12685,N_13248);
nor U15216 (N_15216,N_13446,N_13071);
nor U15217 (N_15217,N_12140,N_12751);
nand U15218 (N_15218,N_13668,N_12842);
nand U15219 (N_15219,N_13156,N_13561);
xor U15220 (N_15220,N_13249,N_13105);
and U15221 (N_15221,N_13944,N_13921);
nand U15222 (N_15222,N_12452,N_12441);
xnor U15223 (N_15223,N_13374,N_12761);
and U15224 (N_15224,N_13467,N_12450);
nand U15225 (N_15225,N_13588,N_13490);
and U15226 (N_15226,N_12063,N_13074);
xnor U15227 (N_15227,N_13039,N_13115);
nor U15228 (N_15228,N_13709,N_13730);
xor U15229 (N_15229,N_12173,N_13670);
and U15230 (N_15230,N_13584,N_13157);
nor U15231 (N_15231,N_13697,N_12178);
nand U15232 (N_15232,N_12054,N_13465);
nand U15233 (N_15233,N_12977,N_13289);
nand U15234 (N_15234,N_13631,N_13126);
xnor U15235 (N_15235,N_13120,N_13604);
or U15236 (N_15236,N_12287,N_12113);
or U15237 (N_15237,N_13062,N_12809);
xor U15238 (N_15238,N_13161,N_12319);
or U15239 (N_15239,N_13497,N_13070);
or U15240 (N_15240,N_13524,N_13875);
nand U15241 (N_15241,N_13069,N_12067);
nor U15242 (N_15242,N_12686,N_12294);
nor U15243 (N_15243,N_13718,N_12521);
nor U15244 (N_15244,N_12037,N_13786);
nor U15245 (N_15245,N_13215,N_12402);
xnor U15246 (N_15246,N_12449,N_13366);
nand U15247 (N_15247,N_13684,N_13053);
nor U15248 (N_15248,N_12902,N_13504);
or U15249 (N_15249,N_12717,N_12009);
nor U15250 (N_15250,N_13814,N_13419);
xor U15251 (N_15251,N_13583,N_12207);
and U15252 (N_15252,N_13018,N_13427);
or U15253 (N_15253,N_12315,N_13917);
nor U15254 (N_15254,N_12070,N_13306);
and U15255 (N_15255,N_13414,N_13647);
xnor U15256 (N_15256,N_13042,N_12146);
xor U15257 (N_15257,N_13407,N_12781);
xor U15258 (N_15258,N_12238,N_12166);
nor U15259 (N_15259,N_12159,N_12464);
and U15260 (N_15260,N_13395,N_12035);
or U15261 (N_15261,N_12503,N_12471);
or U15262 (N_15262,N_13091,N_12575);
or U15263 (N_15263,N_12825,N_13486);
and U15264 (N_15264,N_12936,N_12120);
or U15265 (N_15265,N_12900,N_13869);
nor U15266 (N_15266,N_12589,N_12623);
nor U15267 (N_15267,N_12526,N_12424);
or U15268 (N_15268,N_12888,N_12447);
nor U15269 (N_15269,N_12970,N_13340);
xnor U15270 (N_15270,N_13174,N_12397);
nand U15271 (N_15271,N_12905,N_13220);
and U15272 (N_15272,N_13044,N_12387);
or U15273 (N_15273,N_13814,N_12342);
or U15274 (N_15274,N_13217,N_12981);
or U15275 (N_15275,N_13616,N_13666);
and U15276 (N_15276,N_13629,N_13452);
nand U15277 (N_15277,N_13054,N_12568);
and U15278 (N_15278,N_12402,N_12821);
nand U15279 (N_15279,N_12782,N_12128);
and U15280 (N_15280,N_13505,N_12821);
xnor U15281 (N_15281,N_13904,N_12585);
nand U15282 (N_15282,N_12653,N_12242);
and U15283 (N_15283,N_13306,N_12031);
xor U15284 (N_15284,N_13630,N_13388);
nand U15285 (N_15285,N_12586,N_13586);
nor U15286 (N_15286,N_13231,N_12024);
xor U15287 (N_15287,N_13529,N_12609);
nand U15288 (N_15288,N_12051,N_13951);
nor U15289 (N_15289,N_12251,N_13735);
nand U15290 (N_15290,N_12330,N_12509);
or U15291 (N_15291,N_12780,N_13677);
xnor U15292 (N_15292,N_12329,N_13320);
xor U15293 (N_15293,N_13582,N_12478);
nor U15294 (N_15294,N_13553,N_13049);
nor U15295 (N_15295,N_12817,N_12009);
xnor U15296 (N_15296,N_12584,N_12156);
nor U15297 (N_15297,N_12088,N_13698);
xor U15298 (N_15298,N_12050,N_13012);
and U15299 (N_15299,N_12969,N_12085);
and U15300 (N_15300,N_12977,N_12742);
xnor U15301 (N_15301,N_13574,N_12784);
and U15302 (N_15302,N_13791,N_12094);
nand U15303 (N_15303,N_12273,N_12699);
xnor U15304 (N_15304,N_13867,N_12738);
xor U15305 (N_15305,N_12231,N_12456);
nand U15306 (N_15306,N_13299,N_13199);
nor U15307 (N_15307,N_13767,N_13869);
xor U15308 (N_15308,N_12549,N_12968);
and U15309 (N_15309,N_13328,N_13955);
xor U15310 (N_15310,N_13771,N_13370);
or U15311 (N_15311,N_12948,N_12059);
nand U15312 (N_15312,N_12095,N_12051);
and U15313 (N_15313,N_12785,N_12925);
or U15314 (N_15314,N_13796,N_13497);
and U15315 (N_15315,N_12194,N_13686);
or U15316 (N_15316,N_13791,N_12895);
xor U15317 (N_15317,N_13293,N_13255);
or U15318 (N_15318,N_12217,N_12793);
and U15319 (N_15319,N_13655,N_12739);
and U15320 (N_15320,N_12841,N_12776);
or U15321 (N_15321,N_13300,N_12182);
xor U15322 (N_15322,N_13361,N_12096);
nor U15323 (N_15323,N_13404,N_12046);
and U15324 (N_15324,N_12612,N_13157);
and U15325 (N_15325,N_12732,N_12600);
or U15326 (N_15326,N_13429,N_12714);
xnor U15327 (N_15327,N_12530,N_13411);
nand U15328 (N_15328,N_13060,N_12298);
and U15329 (N_15329,N_13019,N_13281);
and U15330 (N_15330,N_12523,N_12383);
nor U15331 (N_15331,N_12973,N_12473);
nor U15332 (N_15332,N_13588,N_13693);
nand U15333 (N_15333,N_13355,N_13479);
and U15334 (N_15334,N_13893,N_12603);
or U15335 (N_15335,N_12633,N_12381);
nand U15336 (N_15336,N_13226,N_13436);
nor U15337 (N_15337,N_12695,N_13770);
and U15338 (N_15338,N_12058,N_12434);
nor U15339 (N_15339,N_13262,N_13977);
and U15340 (N_15340,N_12394,N_12636);
nor U15341 (N_15341,N_13669,N_13772);
xnor U15342 (N_15342,N_13447,N_12197);
nand U15343 (N_15343,N_12735,N_12683);
and U15344 (N_15344,N_13495,N_13395);
nor U15345 (N_15345,N_13439,N_12402);
or U15346 (N_15346,N_13690,N_12376);
or U15347 (N_15347,N_12475,N_13155);
xnor U15348 (N_15348,N_12276,N_12207);
or U15349 (N_15349,N_13829,N_12565);
nor U15350 (N_15350,N_13882,N_13188);
nand U15351 (N_15351,N_12453,N_13783);
xnor U15352 (N_15352,N_12281,N_13803);
nor U15353 (N_15353,N_13878,N_13461);
xnor U15354 (N_15354,N_12003,N_13761);
or U15355 (N_15355,N_12605,N_13536);
nor U15356 (N_15356,N_13037,N_12890);
and U15357 (N_15357,N_13346,N_13949);
and U15358 (N_15358,N_12075,N_12574);
or U15359 (N_15359,N_13514,N_12094);
xor U15360 (N_15360,N_13661,N_13563);
nand U15361 (N_15361,N_13733,N_13809);
nor U15362 (N_15362,N_13186,N_12213);
nand U15363 (N_15363,N_12648,N_13992);
nand U15364 (N_15364,N_12987,N_12495);
nor U15365 (N_15365,N_12989,N_12962);
nand U15366 (N_15366,N_12962,N_12749);
and U15367 (N_15367,N_12122,N_13285);
xnor U15368 (N_15368,N_13398,N_12070);
or U15369 (N_15369,N_13932,N_13253);
or U15370 (N_15370,N_13226,N_12173);
or U15371 (N_15371,N_13128,N_13369);
xor U15372 (N_15372,N_12268,N_12180);
and U15373 (N_15373,N_13287,N_12266);
nand U15374 (N_15374,N_12333,N_13332);
and U15375 (N_15375,N_13433,N_12322);
or U15376 (N_15376,N_13383,N_13747);
nor U15377 (N_15377,N_13385,N_13326);
or U15378 (N_15378,N_12281,N_12946);
nand U15379 (N_15379,N_13394,N_13727);
and U15380 (N_15380,N_13183,N_13656);
or U15381 (N_15381,N_12428,N_12615);
nand U15382 (N_15382,N_13863,N_12306);
nand U15383 (N_15383,N_13788,N_13696);
nor U15384 (N_15384,N_12946,N_12586);
nand U15385 (N_15385,N_12083,N_13887);
and U15386 (N_15386,N_12777,N_13992);
or U15387 (N_15387,N_13359,N_12338);
xnor U15388 (N_15388,N_13249,N_12273);
or U15389 (N_15389,N_12833,N_13893);
and U15390 (N_15390,N_13407,N_12989);
and U15391 (N_15391,N_13138,N_12070);
and U15392 (N_15392,N_12112,N_13525);
or U15393 (N_15393,N_13379,N_13436);
nand U15394 (N_15394,N_12196,N_12689);
xor U15395 (N_15395,N_13149,N_13122);
and U15396 (N_15396,N_12903,N_12081);
nand U15397 (N_15397,N_12772,N_12664);
or U15398 (N_15398,N_13329,N_13498);
and U15399 (N_15399,N_12373,N_13383);
or U15400 (N_15400,N_13535,N_12174);
and U15401 (N_15401,N_13148,N_13575);
nor U15402 (N_15402,N_12540,N_12061);
nand U15403 (N_15403,N_12834,N_13288);
and U15404 (N_15404,N_13063,N_13561);
nor U15405 (N_15405,N_12010,N_12388);
nor U15406 (N_15406,N_13362,N_12089);
and U15407 (N_15407,N_13067,N_13393);
nor U15408 (N_15408,N_12586,N_12797);
and U15409 (N_15409,N_12659,N_12048);
and U15410 (N_15410,N_13529,N_13372);
or U15411 (N_15411,N_13941,N_13438);
nand U15412 (N_15412,N_12763,N_12654);
and U15413 (N_15413,N_13747,N_12519);
xor U15414 (N_15414,N_12082,N_12026);
and U15415 (N_15415,N_13675,N_12454);
xor U15416 (N_15416,N_12543,N_13513);
xor U15417 (N_15417,N_13744,N_12766);
or U15418 (N_15418,N_13108,N_13189);
or U15419 (N_15419,N_12291,N_12080);
or U15420 (N_15420,N_12763,N_12432);
nor U15421 (N_15421,N_12892,N_13462);
nor U15422 (N_15422,N_12886,N_12878);
and U15423 (N_15423,N_12135,N_13625);
and U15424 (N_15424,N_12276,N_13123);
or U15425 (N_15425,N_12170,N_12083);
and U15426 (N_15426,N_13109,N_12140);
and U15427 (N_15427,N_13108,N_13899);
and U15428 (N_15428,N_12530,N_12481);
or U15429 (N_15429,N_13798,N_13000);
or U15430 (N_15430,N_13052,N_12003);
or U15431 (N_15431,N_12373,N_13225);
nand U15432 (N_15432,N_12426,N_12170);
and U15433 (N_15433,N_12808,N_12851);
nand U15434 (N_15434,N_12159,N_13714);
nor U15435 (N_15435,N_12450,N_12720);
nor U15436 (N_15436,N_13323,N_13547);
nand U15437 (N_15437,N_12410,N_12405);
or U15438 (N_15438,N_12731,N_12090);
nand U15439 (N_15439,N_13457,N_13219);
or U15440 (N_15440,N_12079,N_12862);
or U15441 (N_15441,N_13111,N_12927);
or U15442 (N_15442,N_12549,N_12874);
and U15443 (N_15443,N_13130,N_12936);
or U15444 (N_15444,N_13234,N_12355);
nor U15445 (N_15445,N_13775,N_13405);
or U15446 (N_15446,N_13681,N_12633);
and U15447 (N_15447,N_12555,N_13440);
nand U15448 (N_15448,N_12618,N_12293);
nand U15449 (N_15449,N_12549,N_12524);
xor U15450 (N_15450,N_13232,N_12323);
or U15451 (N_15451,N_13835,N_13307);
nor U15452 (N_15452,N_13959,N_12545);
xnor U15453 (N_15453,N_12680,N_13714);
and U15454 (N_15454,N_12184,N_13263);
xor U15455 (N_15455,N_12106,N_13590);
and U15456 (N_15456,N_13219,N_12899);
or U15457 (N_15457,N_13915,N_13555);
and U15458 (N_15458,N_13021,N_12534);
and U15459 (N_15459,N_13362,N_13395);
and U15460 (N_15460,N_13296,N_12022);
nand U15461 (N_15461,N_12581,N_12420);
and U15462 (N_15462,N_13946,N_13790);
nor U15463 (N_15463,N_12049,N_12422);
or U15464 (N_15464,N_12900,N_12189);
xor U15465 (N_15465,N_13657,N_12460);
xor U15466 (N_15466,N_13054,N_13833);
nand U15467 (N_15467,N_12453,N_13400);
or U15468 (N_15468,N_13430,N_12612);
xor U15469 (N_15469,N_13939,N_13607);
nor U15470 (N_15470,N_12867,N_12394);
nor U15471 (N_15471,N_12385,N_12530);
nor U15472 (N_15472,N_12574,N_12488);
nand U15473 (N_15473,N_13470,N_12205);
and U15474 (N_15474,N_13068,N_13146);
and U15475 (N_15475,N_12949,N_13137);
nand U15476 (N_15476,N_13589,N_13987);
or U15477 (N_15477,N_13137,N_12781);
or U15478 (N_15478,N_13769,N_12421);
nor U15479 (N_15479,N_12500,N_13810);
and U15480 (N_15480,N_13464,N_13132);
nor U15481 (N_15481,N_13053,N_12325);
nor U15482 (N_15482,N_12086,N_12439);
nand U15483 (N_15483,N_13501,N_12768);
and U15484 (N_15484,N_12448,N_13198);
nand U15485 (N_15485,N_13613,N_13383);
or U15486 (N_15486,N_13025,N_12454);
nand U15487 (N_15487,N_13759,N_13756);
xnor U15488 (N_15488,N_12635,N_13477);
or U15489 (N_15489,N_12512,N_13726);
and U15490 (N_15490,N_12949,N_13512);
nand U15491 (N_15491,N_12348,N_13520);
or U15492 (N_15492,N_12666,N_12089);
nand U15493 (N_15493,N_13612,N_12716);
or U15494 (N_15494,N_12094,N_13082);
or U15495 (N_15495,N_12934,N_12095);
or U15496 (N_15496,N_13938,N_12212);
nand U15497 (N_15497,N_12704,N_13189);
and U15498 (N_15498,N_13783,N_12861);
nand U15499 (N_15499,N_13812,N_12406);
xor U15500 (N_15500,N_12464,N_12535);
xnor U15501 (N_15501,N_13151,N_12734);
nor U15502 (N_15502,N_13695,N_12388);
nor U15503 (N_15503,N_12301,N_12744);
or U15504 (N_15504,N_12777,N_13486);
or U15505 (N_15505,N_13571,N_13580);
and U15506 (N_15506,N_13809,N_12761);
xor U15507 (N_15507,N_13226,N_12601);
xnor U15508 (N_15508,N_13904,N_13886);
nand U15509 (N_15509,N_12093,N_12842);
or U15510 (N_15510,N_13083,N_12548);
nand U15511 (N_15511,N_13528,N_13336);
xnor U15512 (N_15512,N_13956,N_12429);
and U15513 (N_15513,N_13806,N_13327);
and U15514 (N_15514,N_13213,N_12001);
xor U15515 (N_15515,N_12406,N_13526);
xor U15516 (N_15516,N_13764,N_12196);
nor U15517 (N_15517,N_13651,N_13345);
nand U15518 (N_15518,N_13495,N_13103);
nor U15519 (N_15519,N_13734,N_13789);
xnor U15520 (N_15520,N_13800,N_12624);
xnor U15521 (N_15521,N_12095,N_13395);
nand U15522 (N_15522,N_13672,N_12712);
nand U15523 (N_15523,N_12934,N_12875);
nand U15524 (N_15524,N_13321,N_13039);
nor U15525 (N_15525,N_12548,N_12165);
or U15526 (N_15526,N_12381,N_12950);
xor U15527 (N_15527,N_12039,N_12860);
or U15528 (N_15528,N_12001,N_13523);
nand U15529 (N_15529,N_12529,N_13684);
nand U15530 (N_15530,N_13006,N_13044);
or U15531 (N_15531,N_13914,N_13720);
nand U15532 (N_15532,N_12674,N_13487);
or U15533 (N_15533,N_12591,N_12213);
nand U15534 (N_15534,N_13537,N_13482);
xnor U15535 (N_15535,N_12136,N_12398);
and U15536 (N_15536,N_13521,N_13286);
or U15537 (N_15537,N_12878,N_13561);
xor U15538 (N_15538,N_13256,N_12946);
and U15539 (N_15539,N_12176,N_13394);
or U15540 (N_15540,N_12440,N_12608);
and U15541 (N_15541,N_12179,N_12479);
and U15542 (N_15542,N_13319,N_13412);
xor U15543 (N_15543,N_12351,N_12297);
nand U15544 (N_15544,N_12468,N_13469);
and U15545 (N_15545,N_12486,N_12978);
and U15546 (N_15546,N_13089,N_13056);
nor U15547 (N_15547,N_13319,N_12958);
nor U15548 (N_15548,N_13015,N_12879);
nand U15549 (N_15549,N_13496,N_12377);
or U15550 (N_15550,N_12549,N_13960);
nand U15551 (N_15551,N_12569,N_13271);
and U15552 (N_15552,N_12468,N_13719);
xnor U15553 (N_15553,N_13597,N_12155);
xor U15554 (N_15554,N_13119,N_13806);
nor U15555 (N_15555,N_12456,N_13968);
or U15556 (N_15556,N_12545,N_12577);
xnor U15557 (N_15557,N_13490,N_12666);
and U15558 (N_15558,N_13964,N_13273);
or U15559 (N_15559,N_13469,N_12902);
nand U15560 (N_15560,N_12716,N_13786);
or U15561 (N_15561,N_13025,N_12303);
nor U15562 (N_15562,N_12876,N_12204);
xor U15563 (N_15563,N_12923,N_12804);
nand U15564 (N_15564,N_12961,N_12499);
xor U15565 (N_15565,N_12587,N_12382);
and U15566 (N_15566,N_13203,N_12658);
nor U15567 (N_15567,N_12118,N_13667);
or U15568 (N_15568,N_12837,N_13266);
or U15569 (N_15569,N_12146,N_13120);
or U15570 (N_15570,N_13032,N_13407);
and U15571 (N_15571,N_12536,N_12638);
nand U15572 (N_15572,N_13754,N_13054);
and U15573 (N_15573,N_13019,N_12222);
nor U15574 (N_15574,N_12559,N_12689);
nand U15575 (N_15575,N_13678,N_12063);
xor U15576 (N_15576,N_12779,N_13431);
nor U15577 (N_15577,N_12808,N_13609);
xor U15578 (N_15578,N_12731,N_12702);
nor U15579 (N_15579,N_13206,N_13138);
or U15580 (N_15580,N_13502,N_13482);
nand U15581 (N_15581,N_12860,N_12657);
nor U15582 (N_15582,N_12368,N_12042);
and U15583 (N_15583,N_12791,N_12182);
nand U15584 (N_15584,N_12066,N_12721);
nor U15585 (N_15585,N_12110,N_12556);
nor U15586 (N_15586,N_12559,N_13772);
nand U15587 (N_15587,N_12618,N_13503);
and U15588 (N_15588,N_12640,N_13710);
xor U15589 (N_15589,N_12769,N_13551);
nor U15590 (N_15590,N_13182,N_13162);
nand U15591 (N_15591,N_13571,N_13822);
xor U15592 (N_15592,N_13362,N_12662);
xnor U15593 (N_15593,N_13901,N_12018);
and U15594 (N_15594,N_13395,N_13842);
nand U15595 (N_15595,N_13547,N_12529);
nor U15596 (N_15596,N_12075,N_13223);
and U15597 (N_15597,N_13304,N_13921);
nand U15598 (N_15598,N_12287,N_13023);
or U15599 (N_15599,N_12249,N_13902);
and U15600 (N_15600,N_13931,N_12142);
or U15601 (N_15601,N_12171,N_12175);
xnor U15602 (N_15602,N_12463,N_12556);
nor U15603 (N_15603,N_13169,N_13913);
nand U15604 (N_15604,N_13482,N_13335);
and U15605 (N_15605,N_12713,N_12515);
or U15606 (N_15606,N_12943,N_12807);
or U15607 (N_15607,N_13491,N_13044);
or U15608 (N_15608,N_13299,N_12151);
nor U15609 (N_15609,N_12358,N_13519);
xor U15610 (N_15610,N_12144,N_12406);
and U15611 (N_15611,N_13986,N_12995);
and U15612 (N_15612,N_12058,N_13739);
and U15613 (N_15613,N_12113,N_12087);
nand U15614 (N_15614,N_13720,N_12792);
nor U15615 (N_15615,N_12161,N_12188);
and U15616 (N_15616,N_12153,N_13715);
or U15617 (N_15617,N_13450,N_12274);
or U15618 (N_15618,N_12022,N_13157);
and U15619 (N_15619,N_12893,N_13073);
nand U15620 (N_15620,N_13587,N_12940);
nor U15621 (N_15621,N_13555,N_13541);
xor U15622 (N_15622,N_12634,N_12295);
and U15623 (N_15623,N_12823,N_13743);
nor U15624 (N_15624,N_13649,N_12670);
nor U15625 (N_15625,N_13602,N_13573);
nand U15626 (N_15626,N_12920,N_12477);
or U15627 (N_15627,N_12906,N_12734);
and U15628 (N_15628,N_12815,N_13082);
xnor U15629 (N_15629,N_13894,N_12362);
or U15630 (N_15630,N_12578,N_12550);
nand U15631 (N_15631,N_12364,N_13377);
nand U15632 (N_15632,N_12197,N_12026);
nand U15633 (N_15633,N_12262,N_12375);
xnor U15634 (N_15634,N_13630,N_13407);
nor U15635 (N_15635,N_12247,N_13319);
or U15636 (N_15636,N_13378,N_13575);
or U15637 (N_15637,N_12607,N_12398);
nor U15638 (N_15638,N_13559,N_13320);
xnor U15639 (N_15639,N_12916,N_13124);
nor U15640 (N_15640,N_13432,N_12606);
nor U15641 (N_15641,N_12420,N_13580);
and U15642 (N_15642,N_12566,N_13777);
xnor U15643 (N_15643,N_13826,N_13377);
or U15644 (N_15644,N_13508,N_12259);
xnor U15645 (N_15645,N_12317,N_13291);
xnor U15646 (N_15646,N_13222,N_12377);
and U15647 (N_15647,N_12008,N_12801);
and U15648 (N_15648,N_12084,N_13099);
nor U15649 (N_15649,N_13196,N_13379);
nand U15650 (N_15650,N_13008,N_12362);
nand U15651 (N_15651,N_12867,N_13537);
or U15652 (N_15652,N_13630,N_12538);
or U15653 (N_15653,N_12772,N_13023);
and U15654 (N_15654,N_13747,N_13835);
or U15655 (N_15655,N_12009,N_12180);
or U15656 (N_15656,N_12532,N_13079);
or U15657 (N_15657,N_12140,N_12503);
and U15658 (N_15658,N_13559,N_12450);
or U15659 (N_15659,N_13104,N_13797);
and U15660 (N_15660,N_12969,N_13986);
xor U15661 (N_15661,N_12592,N_13915);
and U15662 (N_15662,N_12900,N_12417);
nor U15663 (N_15663,N_12164,N_12748);
xor U15664 (N_15664,N_12996,N_13918);
and U15665 (N_15665,N_13448,N_13932);
xnor U15666 (N_15666,N_13372,N_12789);
nand U15667 (N_15667,N_13963,N_13186);
xnor U15668 (N_15668,N_12495,N_13067);
nor U15669 (N_15669,N_13273,N_13643);
or U15670 (N_15670,N_12538,N_12423);
or U15671 (N_15671,N_13223,N_12317);
nand U15672 (N_15672,N_13371,N_13458);
xor U15673 (N_15673,N_12455,N_12726);
xor U15674 (N_15674,N_13286,N_12631);
nand U15675 (N_15675,N_13396,N_13084);
and U15676 (N_15676,N_12610,N_13287);
nor U15677 (N_15677,N_12876,N_12437);
xor U15678 (N_15678,N_13078,N_13908);
nor U15679 (N_15679,N_12742,N_12979);
and U15680 (N_15680,N_12022,N_13074);
xor U15681 (N_15681,N_12278,N_12561);
and U15682 (N_15682,N_13712,N_13360);
xor U15683 (N_15683,N_12369,N_13421);
and U15684 (N_15684,N_12426,N_13079);
or U15685 (N_15685,N_13103,N_13092);
and U15686 (N_15686,N_12229,N_13808);
nor U15687 (N_15687,N_12716,N_13146);
nor U15688 (N_15688,N_12127,N_13142);
and U15689 (N_15689,N_12337,N_12373);
xor U15690 (N_15690,N_13587,N_12599);
nor U15691 (N_15691,N_13613,N_12496);
nand U15692 (N_15692,N_13397,N_12293);
and U15693 (N_15693,N_12039,N_13469);
or U15694 (N_15694,N_12369,N_13585);
nand U15695 (N_15695,N_13843,N_12915);
or U15696 (N_15696,N_12139,N_13334);
or U15697 (N_15697,N_12376,N_12864);
nand U15698 (N_15698,N_12021,N_13764);
or U15699 (N_15699,N_13104,N_12861);
xor U15700 (N_15700,N_13109,N_12936);
or U15701 (N_15701,N_13260,N_13342);
nor U15702 (N_15702,N_13891,N_12544);
or U15703 (N_15703,N_12777,N_12074);
nand U15704 (N_15704,N_13239,N_13920);
xor U15705 (N_15705,N_12060,N_12630);
xnor U15706 (N_15706,N_12431,N_12007);
nand U15707 (N_15707,N_12892,N_13429);
and U15708 (N_15708,N_12886,N_12188);
nor U15709 (N_15709,N_13340,N_13148);
nand U15710 (N_15710,N_12897,N_13325);
nor U15711 (N_15711,N_12648,N_13467);
nand U15712 (N_15712,N_13454,N_12967);
nand U15713 (N_15713,N_12328,N_12643);
xor U15714 (N_15714,N_12275,N_12210);
or U15715 (N_15715,N_13554,N_12425);
nand U15716 (N_15716,N_13257,N_12371);
or U15717 (N_15717,N_13430,N_13652);
nor U15718 (N_15718,N_12831,N_13922);
nand U15719 (N_15719,N_13163,N_12657);
and U15720 (N_15720,N_12198,N_12673);
or U15721 (N_15721,N_13214,N_12497);
nand U15722 (N_15722,N_13733,N_13094);
and U15723 (N_15723,N_13833,N_12905);
xnor U15724 (N_15724,N_12771,N_13230);
xor U15725 (N_15725,N_13211,N_12117);
or U15726 (N_15726,N_12610,N_12486);
nor U15727 (N_15727,N_13365,N_12140);
and U15728 (N_15728,N_13510,N_12079);
and U15729 (N_15729,N_12945,N_13252);
nor U15730 (N_15730,N_12772,N_13723);
or U15731 (N_15731,N_13948,N_12302);
xor U15732 (N_15732,N_12506,N_12664);
or U15733 (N_15733,N_13132,N_12275);
nor U15734 (N_15734,N_13142,N_13564);
xor U15735 (N_15735,N_12014,N_12203);
or U15736 (N_15736,N_12768,N_12440);
nor U15737 (N_15737,N_12361,N_12871);
nand U15738 (N_15738,N_13545,N_12713);
or U15739 (N_15739,N_13486,N_13980);
or U15740 (N_15740,N_12861,N_12335);
nand U15741 (N_15741,N_12633,N_12166);
and U15742 (N_15742,N_13657,N_12374);
and U15743 (N_15743,N_13396,N_12198);
nand U15744 (N_15744,N_13584,N_13786);
nor U15745 (N_15745,N_12098,N_12418);
nor U15746 (N_15746,N_12747,N_12205);
nor U15747 (N_15747,N_13623,N_12030);
nand U15748 (N_15748,N_13033,N_12387);
nor U15749 (N_15749,N_13642,N_12039);
nor U15750 (N_15750,N_12963,N_12238);
and U15751 (N_15751,N_12300,N_13537);
and U15752 (N_15752,N_13001,N_12699);
and U15753 (N_15753,N_12011,N_13012);
nor U15754 (N_15754,N_12228,N_12053);
nand U15755 (N_15755,N_13462,N_13173);
nand U15756 (N_15756,N_12007,N_12401);
or U15757 (N_15757,N_12992,N_13218);
xor U15758 (N_15758,N_12587,N_13824);
and U15759 (N_15759,N_13018,N_13212);
nand U15760 (N_15760,N_12679,N_12398);
nor U15761 (N_15761,N_12114,N_13966);
nand U15762 (N_15762,N_13365,N_12307);
nor U15763 (N_15763,N_13711,N_12196);
xor U15764 (N_15764,N_12191,N_13438);
or U15765 (N_15765,N_12546,N_13260);
and U15766 (N_15766,N_13668,N_13852);
nand U15767 (N_15767,N_13094,N_13994);
nor U15768 (N_15768,N_13987,N_13110);
nand U15769 (N_15769,N_13961,N_12138);
and U15770 (N_15770,N_13244,N_13983);
nor U15771 (N_15771,N_12925,N_13236);
and U15772 (N_15772,N_12616,N_12714);
nand U15773 (N_15773,N_13898,N_13101);
or U15774 (N_15774,N_13299,N_12339);
nor U15775 (N_15775,N_12003,N_12139);
xnor U15776 (N_15776,N_13087,N_13628);
xor U15777 (N_15777,N_13264,N_13987);
and U15778 (N_15778,N_13023,N_13313);
nor U15779 (N_15779,N_12622,N_13859);
or U15780 (N_15780,N_13525,N_12604);
xnor U15781 (N_15781,N_13610,N_12440);
nand U15782 (N_15782,N_12677,N_12827);
xor U15783 (N_15783,N_12257,N_13248);
nand U15784 (N_15784,N_13513,N_12004);
and U15785 (N_15785,N_12226,N_12096);
or U15786 (N_15786,N_12153,N_12173);
and U15787 (N_15787,N_12182,N_13838);
or U15788 (N_15788,N_13860,N_12032);
nand U15789 (N_15789,N_13320,N_13536);
nor U15790 (N_15790,N_13266,N_12200);
xnor U15791 (N_15791,N_12906,N_12325);
nand U15792 (N_15792,N_13136,N_13974);
and U15793 (N_15793,N_12160,N_13923);
and U15794 (N_15794,N_12386,N_12255);
nor U15795 (N_15795,N_13633,N_12301);
nor U15796 (N_15796,N_12440,N_13891);
or U15797 (N_15797,N_12059,N_13914);
nand U15798 (N_15798,N_13175,N_12728);
xor U15799 (N_15799,N_13047,N_12750);
nor U15800 (N_15800,N_13154,N_12189);
and U15801 (N_15801,N_13466,N_12766);
xor U15802 (N_15802,N_12936,N_13384);
or U15803 (N_15803,N_12713,N_13230);
or U15804 (N_15804,N_13305,N_13651);
xnor U15805 (N_15805,N_12569,N_12145);
xnor U15806 (N_15806,N_13865,N_12153);
nand U15807 (N_15807,N_13476,N_12133);
and U15808 (N_15808,N_12652,N_13831);
xor U15809 (N_15809,N_13689,N_13638);
xnor U15810 (N_15810,N_12017,N_13207);
and U15811 (N_15811,N_13593,N_12519);
nor U15812 (N_15812,N_13797,N_12072);
or U15813 (N_15813,N_13680,N_13364);
nor U15814 (N_15814,N_13147,N_12778);
or U15815 (N_15815,N_12973,N_12799);
xnor U15816 (N_15816,N_13802,N_12951);
nand U15817 (N_15817,N_13952,N_12807);
and U15818 (N_15818,N_13761,N_12712);
xnor U15819 (N_15819,N_13001,N_12515);
xor U15820 (N_15820,N_13009,N_13884);
or U15821 (N_15821,N_12861,N_13566);
or U15822 (N_15822,N_13918,N_12107);
and U15823 (N_15823,N_12519,N_12819);
nor U15824 (N_15824,N_12072,N_13586);
xor U15825 (N_15825,N_13823,N_13474);
nor U15826 (N_15826,N_13463,N_13514);
xnor U15827 (N_15827,N_12877,N_12726);
xnor U15828 (N_15828,N_12841,N_13246);
or U15829 (N_15829,N_13415,N_12686);
xnor U15830 (N_15830,N_12947,N_13669);
nor U15831 (N_15831,N_12967,N_12685);
xnor U15832 (N_15832,N_13655,N_13680);
nand U15833 (N_15833,N_12428,N_12502);
and U15834 (N_15834,N_13590,N_13200);
nand U15835 (N_15835,N_13596,N_13236);
and U15836 (N_15836,N_12718,N_13316);
or U15837 (N_15837,N_12852,N_12847);
and U15838 (N_15838,N_12709,N_12724);
xnor U15839 (N_15839,N_13527,N_12078);
nor U15840 (N_15840,N_13691,N_12842);
nor U15841 (N_15841,N_13357,N_13617);
or U15842 (N_15842,N_12827,N_12624);
or U15843 (N_15843,N_12183,N_13245);
nand U15844 (N_15844,N_13662,N_13628);
nor U15845 (N_15845,N_13473,N_12443);
or U15846 (N_15846,N_13465,N_12442);
and U15847 (N_15847,N_13473,N_13840);
or U15848 (N_15848,N_12313,N_12144);
nand U15849 (N_15849,N_13359,N_12312);
xor U15850 (N_15850,N_13487,N_12838);
and U15851 (N_15851,N_13566,N_12087);
or U15852 (N_15852,N_12983,N_12736);
and U15853 (N_15853,N_12975,N_13203);
nor U15854 (N_15854,N_12207,N_13186);
nor U15855 (N_15855,N_13460,N_12225);
and U15856 (N_15856,N_12397,N_12247);
xnor U15857 (N_15857,N_13515,N_13819);
or U15858 (N_15858,N_12947,N_13718);
nor U15859 (N_15859,N_12096,N_13790);
xor U15860 (N_15860,N_13497,N_13567);
and U15861 (N_15861,N_12622,N_12199);
xor U15862 (N_15862,N_12024,N_13692);
or U15863 (N_15863,N_13769,N_12019);
nor U15864 (N_15864,N_13353,N_13197);
and U15865 (N_15865,N_13415,N_12766);
nand U15866 (N_15866,N_12602,N_12880);
and U15867 (N_15867,N_12966,N_13637);
nand U15868 (N_15868,N_12848,N_12317);
xor U15869 (N_15869,N_12918,N_12425);
or U15870 (N_15870,N_12572,N_13700);
xnor U15871 (N_15871,N_12244,N_12159);
and U15872 (N_15872,N_12312,N_13703);
and U15873 (N_15873,N_12376,N_13608);
xor U15874 (N_15874,N_12332,N_12569);
nor U15875 (N_15875,N_13115,N_12629);
nor U15876 (N_15876,N_12163,N_12451);
and U15877 (N_15877,N_12009,N_12470);
nor U15878 (N_15878,N_13935,N_13043);
nor U15879 (N_15879,N_12160,N_13851);
xor U15880 (N_15880,N_12757,N_13096);
or U15881 (N_15881,N_13356,N_13514);
nor U15882 (N_15882,N_12631,N_13715);
and U15883 (N_15883,N_13511,N_13727);
xnor U15884 (N_15884,N_12072,N_13133);
nand U15885 (N_15885,N_13806,N_12297);
nand U15886 (N_15886,N_13126,N_13991);
and U15887 (N_15887,N_12509,N_13205);
nand U15888 (N_15888,N_12445,N_12229);
or U15889 (N_15889,N_12130,N_12735);
xor U15890 (N_15890,N_12089,N_13067);
or U15891 (N_15891,N_13074,N_13054);
nand U15892 (N_15892,N_12635,N_12910);
or U15893 (N_15893,N_13091,N_12885);
nand U15894 (N_15894,N_12488,N_13406);
nand U15895 (N_15895,N_12177,N_12091);
and U15896 (N_15896,N_13593,N_12787);
xnor U15897 (N_15897,N_13196,N_12294);
and U15898 (N_15898,N_13582,N_12434);
or U15899 (N_15899,N_13187,N_12591);
or U15900 (N_15900,N_12455,N_12494);
or U15901 (N_15901,N_12394,N_13288);
nor U15902 (N_15902,N_12267,N_13362);
nor U15903 (N_15903,N_12772,N_13902);
and U15904 (N_15904,N_13662,N_12555);
or U15905 (N_15905,N_12072,N_12687);
and U15906 (N_15906,N_12661,N_12334);
xnor U15907 (N_15907,N_13657,N_13917);
xnor U15908 (N_15908,N_12008,N_12260);
xnor U15909 (N_15909,N_13987,N_12410);
and U15910 (N_15910,N_12573,N_12990);
and U15911 (N_15911,N_13248,N_13164);
or U15912 (N_15912,N_13538,N_12189);
and U15913 (N_15913,N_12411,N_13230);
and U15914 (N_15914,N_13249,N_12550);
and U15915 (N_15915,N_13057,N_13693);
or U15916 (N_15916,N_13614,N_12623);
or U15917 (N_15917,N_13725,N_13106);
nand U15918 (N_15918,N_12703,N_12511);
xnor U15919 (N_15919,N_12843,N_13932);
or U15920 (N_15920,N_13198,N_12397);
and U15921 (N_15921,N_12823,N_13708);
nor U15922 (N_15922,N_13406,N_13052);
nor U15923 (N_15923,N_12204,N_12626);
or U15924 (N_15924,N_12167,N_13026);
xor U15925 (N_15925,N_12825,N_12962);
nand U15926 (N_15926,N_13813,N_13456);
or U15927 (N_15927,N_13215,N_12267);
or U15928 (N_15928,N_13548,N_12383);
nand U15929 (N_15929,N_13132,N_12609);
or U15930 (N_15930,N_13792,N_12914);
or U15931 (N_15931,N_12446,N_12838);
or U15932 (N_15932,N_12354,N_12990);
nor U15933 (N_15933,N_13925,N_12963);
and U15934 (N_15934,N_12428,N_13165);
nand U15935 (N_15935,N_13868,N_13391);
nand U15936 (N_15936,N_12546,N_13920);
and U15937 (N_15937,N_13126,N_13578);
nor U15938 (N_15938,N_12057,N_13173);
nor U15939 (N_15939,N_12291,N_13267);
nand U15940 (N_15940,N_13412,N_12920);
and U15941 (N_15941,N_12612,N_12916);
or U15942 (N_15942,N_13834,N_12392);
xnor U15943 (N_15943,N_12149,N_12903);
nand U15944 (N_15944,N_13943,N_12204);
nand U15945 (N_15945,N_13278,N_12600);
nor U15946 (N_15946,N_13282,N_12182);
and U15947 (N_15947,N_12476,N_13365);
xnor U15948 (N_15948,N_13100,N_13372);
nor U15949 (N_15949,N_12461,N_12342);
and U15950 (N_15950,N_12185,N_13500);
and U15951 (N_15951,N_12701,N_12258);
nor U15952 (N_15952,N_13762,N_13031);
nor U15953 (N_15953,N_13455,N_12942);
or U15954 (N_15954,N_12877,N_12760);
nor U15955 (N_15955,N_12595,N_12927);
or U15956 (N_15956,N_12704,N_13949);
and U15957 (N_15957,N_13371,N_13769);
and U15958 (N_15958,N_13617,N_13996);
nand U15959 (N_15959,N_12244,N_13508);
nand U15960 (N_15960,N_12868,N_12341);
or U15961 (N_15961,N_12420,N_13687);
nand U15962 (N_15962,N_12166,N_12618);
or U15963 (N_15963,N_12615,N_13609);
xnor U15964 (N_15964,N_13335,N_13530);
nand U15965 (N_15965,N_12229,N_13340);
nor U15966 (N_15966,N_13986,N_12353);
nor U15967 (N_15967,N_12867,N_13148);
nand U15968 (N_15968,N_12891,N_13749);
xnor U15969 (N_15969,N_13715,N_13005);
nor U15970 (N_15970,N_12932,N_12396);
nor U15971 (N_15971,N_13583,N_12153);
xor U15972 (N_15972,N_12547,N_12690);
nand U15973 (N_15973,N_13007,N_13296);
nor U15974 (N_15974,N_12702,N_12499);
nand U15975 (N_15975,N_13200,N_12518);
or U15976 (N_15976,N_12049,N_12684);
nand U15977 (N_15977,N_13553,N_13646);
nand U15978 (N_15978,N_12777,N_13171);
nand U15979 (N_15979,N_12965,N_13635);
nand U15980 (N_15980,N_12405,N_12284);
or U15981 (N_15981,N_13915,N_13480);
and U15982 (N_15982,N_13500,N_13682);
and U15983 (N_15983,N_13389,N_12739);
xor U15984 (N_15984,N_13273,N_13268);
or U15985 (N_15985,N_12026,N_12586);
and U15986 (N_15986,N_13700,N_12021);
nor U15987 (N_15987,N_13056,N_12727);
or U15988 (N_15988,N_12228,N_13195);
nor U15989 (N_15989,N_12311,N_12641);
nor U15990 (N_15990,N_13708,N_13039);
or U15991 (N_15991,N_13417,N_13653);
or U15992 (N_15992,N_12360,N_12269);
or U15993 (N_15993,N_13429,N_12149);
xnor U15994 (N_15994,N_13558,N_12836);
nor U15995 (N_15995,N_13996,N_12237);
xor U15996 (N_15996,N_12442,N_12268);
and U15997 (N_15997,N_13706,N_12774);
nor U15998 (N_15998,N_13573,N_12266);
and U15999 (N_15999,N_13330,N_13557);
xnor U16000 (N_16000,N_14051,N_14310);
or U16001 (N_16001,N_14294,N_15636);
xor U16002 (N_16002,N_14233,N_15772);
nand U16003 (N_16003,N_14222,N_14651);
nand U16004 (N_16004,N_14205,N_15907);
and U16005 (N_16005,N_14068,N_15961);
nor U16006 (N_16006,N_14836,N_15930);
xnor U16007 (N_16007,N_15076,N_14073);
or U16008 (N_16008,N_15047,N_14638);
and U16009 (N_16009,N_14047,N_15672);
nor U16010 (N_16010,N_15426,N_15006);
nand U16011 (N_16011,N_15832,N_14612);
nor U16012 (N_16012,N_15881,N_14594);
or U16013 (N_16013,N_15761,N_14963);
nand U16014 (N_16014,N_15387,N_14718);
or U16015 (N_16015,N_14693,N_15141);
nor U16016 (N_16016,N_15021,N_15521);
or U16017 (N_16017,N_14914,N_15234);
and U16018 (N_16018,N_14758,N_15785);
nor U16019 (N_16019,N_14636,N_14216);
xnor U16020 (N_16020,N_15773,N_14690);
xor U16021 (N_16021,N_15688,N_15026);
nor U16022 (N_16022,N_15470,N_14146);
or U16023 (N_16023,N_15032,N_14588);
or U16024 (N_16024,N_14004,N_15992);
nor U16025 (N_16025,N_15462,N_15430);
nand U16026 (N_16026,N_15108,N_14341);
nand U16027 (N_16027,N_14140,N_15712);
xor U16028 (N_16028,N_15856,N_15455);
nor U16029 (N_16029,N_15633,N_14145);
nand U16030 (N_16030,N_14811,N_15257);
or U16031 (N_16031,N_14157,N_14895);
nor U16032 (N_16032,N_14135,N_15517);
xor U16033 (N_16033,N_14962,N_14517);
nor U16034 (N_16034,N_14491,N_15184);
nand U16035 (N_16035,N_15869,N_15478);
or U16036 (N_16036,N_14655,N_15438);
or U16037 (N_16037,N_14451,N_15227);
nor U16038 (N_16038,N_15694,N_15115);
nand U16039 (N_16039,N_15147,N_14650);
and U16040 (N_16040,N_14452,N_15955);
nand U16041 (N_16041,N_14494,N_15499);
nand U16042 (N_16042,N_15632,N_14030);
or U16043 (N_16043,N_15657,N_14862);
nor U16044 (N_16044,N_15619,N_14761);
nor U16045 (N_16045,N_15029,N_14695);
nor U16046 (N_16046,N_15651,N_15630);
xor U16047 (N_16047,N_15638,N_15028);
nor U16048 (N_16048,N_15725,N_15213);
nand U16049 (N_16049,N_15963,N_15642);
or U16050 (N_16050,N_14187,N_15728);
or U16051 (N_16051,N_15755,N_14337);
or U16052 (N_16052,N_14119,N_15970);
nand U16053 (N_16053,N_14617,N_14580);
and U16054 (N_16054,N_14344,N_15854);
nor U16055 (N_16055,N_14391,N_15165);
and U16056 (N_16056,N_15464,N_14592);
xor U16057 (N_16057,N_14720,N_14256);
and U16058 (N_16058,N_15899,N_14887);
and U16059 (N_16059,N_15673,N_14502);
nor U16060 (N_16060,N_14953,N_14029);
nand U16061 (N_16061,N_15779,N_14893);
and U16062 (N_16062,N_14958,N_14738);
nand U16063 (N_16063,N_14375,N_14192);
or U16064 (N_16064,N_14826,N_14669);
nand U16065 (N_16065,N_14453,N_15824);
or U16066 (N_16066,N_14608,N_15127);
or U16067 (N_16067,N_14522,N_15682);
and U16068 (N_16068,N_15681,N_14759);
xor U16069 (N_16069,N_14353,N_15668);
and U16070 (N_16070,N_15142,N_14412);
nor U16071 (N_16071,N_14202,N_15511);
and U16072 (N_16072,N_15372,N_15847);
xnor U16073 (N_16073,N_14463,N_14723);
or U16074 (N_16074,N_15014,N_14242);
xnor U16075 (N_16075,N_15878,N_14629);
nand U16076 (N_16076,N_15046,N_15347);
nor U16077 (N_16077,N_14010,N_14214);
xor U16078 (N_16078,N_15523,N_14854);
nor U16079 (N_16079,N_14539,N_15676);
nand U16080 (N_16080,N_14628,N_14886);
nor U16081 (N_16081,N_14911,N_14957);
xor U16082 (N_16082,N_14841,N_14827);
or U16083 (N_16083,N_15034,N_14998);
nor U16084 (N_16084,N_15648,N_14550);
nor U16085 (N_16085,N_14076,N_14942);
nand U16086 (N_16086,N_14467,N_15095);
and U16087 (N_16087,N_15553,N_15435);
nor U16088 (N_16088,N_15312,N_14392);
or U16089 (N_16089,N_15828,N_15411);
xor U16090 (N_16090,N_14368,N_14888);
nor U16091 (N_16091,N_15285,N_14874);
nor U16092 (N_16092,N_14171,N_15802);
or U16093 (N_16093,N_15889,N_14034);
or U16094 (N_16094,N_14218,N_15966);
nor U16095 (N_16095,N_14945,N_15259);
xnor U16096 (N_16096,N_15666,N_15857);
nor U16097 (N_16097,N_15538,N_14177);
or U16098 (N_16098,N_15621,N_14969);
and U16099 (N_16099,N_15152,N_14543);
xor U16100 (N_16100,N_15224,N_15090);
xnor U16101 (N_16101,N_15405,N_15965);
or U16102 (N_16102,N_14829,N_15422);
and U16103 (N_16103,N_14993,N_15902);
or U16104 (N_16104,N_15071,N_14511);
or U16105 (N_16105,N_14288,N_15010);
nor U16106 (N_16106,N_14990,N_14148);
xnor U16107 (N_16107,N_14560,N_15222);
nor U16108 (N_16108,N_14763,N_15585);
xnor U16109 (N_16109,N_15567,N_15606);
nand U16110 (N_16110,N_15448,N_15377);
or U16111 (N_16111,N_14744,N_14696);
nor U16112 (N_16112,N_15256,N_15116);
or U16113 (N_16113,N_14038,N_15101);
nand U16114 (N_16114,N_14673,N_15043);
nand U16115 (N_16115,N_14386,N_14694);
xnor U16116 (N_16116,N_14885,N_15846);
nor U16117 (N_16117,N_14845,N_15089);
nand U16118 (N_16118,N_14363,N_14587);
or U16119 (N_16119,N_14684,N_14204);
and U16120 (N_16120,N_14141,N_15231);
and U16121 (N_16121,N_14406,N_15226);
and U16122 (N_16122,N_15744,N_15137);
and U16123 (N_16123,N_14975,N_14479);
or U16124 (N_16124,N_15397,N_15172);
xor U16125 (N_16125,N_15486,N_14301);
nand U16126 (N_16126,N_14848,N_15806);
or U16127 (N_16127,N_15713,N_14727);
nor U16128 (N_16128,N_14852,N_15178);
nand U16129 (N_16129,N_14474,N_14999);
xor U16130 (N_16130,N_15102,N_15583);
and U16131 (N_16131,N_14324,N_15436);
and U16132 (N_16132,N_15807,N_15526);
and U16133 (N_16133,N_14524,N_14314);
and U16134 (N_16134,N_15106,N_14036);
or U16135 (N_16135,N_15193,N_15879);
or U16136 (N_16136,N_15974,N_14797);
nor U16137 (N_16137,N_14287,N_14509);
or U16138 (N_16138,N_15004,N_14615);
xor U16139 (N_16139,N_14475,N_15876);
and U16140 (N_16140,N_14871,N_15508);
and U16141 (N_16141,N_14211,N_15041);
nand U16142 (N_16142,N_15243,N_14109);
or U16143 (N_16143,N_14173,N_15914);
nand U16144 (N_16144,N_14482,N_15645);
and U16145 (N_16145,N_15975,N_14290);
and U16146 (N_16146,N_14947,N_14316);
or U16147 (N_16147,N_14994,N_15817);
nand U16148 (N_16148,N_15297,N_15431);
and U16149 (N_16149,N_14203,N_15888);
or U16150 (N_16150,N_14997,N_14924);
and U16151 (N_16151,N_15404,N_15597);
xor U16152 (N_16152,N_14544,N_15505);
nand U16153 (N_16153,N_14199,N_15190);
or U16154 (N_16154,N_14825,N_14666);
nor U16155 (N_16155,N_14901,N_14422);
and U16156 (N_16156,N_14151,N_15057);
and U16157 (N_16157,N_14163,N_14193);
nor U16158 (N_16158,N_14159,N_15983);
nand U16159 (N_16159,N_15420,N_14915);
xor U16160 (N_16160,N_15502,N_15515);
nor U16161 (N_16161,N_14261,N_14627);
nand U16162 (N_16162,N_14737,N_15616);
or U16163 (N_16163,N_15530,N_14367);
xnor U16164 (N_16164,N_14323,N_15734);
or U16165 (N_16165,N_15920,N_14147);
xor U16166 (N_16166,N_15622,N_14069);
xor U16167 (N_16167,N_14860,N_15180);
or U16168 (N_16168,N_15308,N_14382);
nor U16169 (N_16169,N_15640,N_14668);
or U16170 (N_16170,N_14979,N_14383);
and U16171 (N_16171,N_14454,N_14625);
nand U16172 (N_16172,N_15836,N_15546);
and U16173 (N_16173,N_15305,N_14951);
xnor U16174 (N_16174,N_15726,N_14918);
nor U16175 (N_16175,N_14447,N_15995);
nand U16176 (N_16176,N_14961,N_14044);
nand U16177 (N_16177,N_15939,N_14390);
and U16178 (N_16178,N_14074,N_15829);
and U16179 (N_16179,N_15037,N_15366);
xnor U16180 (N_16180,N_14439,N_14903);
xor U16181 (N_16181,N_15655,N_15985);
or U16182 (N_16182,N_14342,N_15803);
nand U16183 (N_16183,N_15381,N_15592);
and U16184 (N_16184,N_14019,N_15011);
nor U16185 (N_16185,N_15368,N_14505);
nor U16186 (N_16186,N_15494,N_15456);
nor U16187 (N_16187,N_14849,N_14906);
xor U16188 (N_16188,N_14514,N_15501);
nand U16189 (N_16189,N_14596,N_14264);
and U16190 (N_16190,N_14967,N_14042);
nor U16191 (N_16191,N_14156,N_14465);
nor U16192 (N_16192,N_14527,N_15428);
nand U16193 (N_16193,N_14080,N_14013);
and U16194 (N_16194,N_15631,N_14533);
or U16195 (N_16195,N_14081,N_15774);
xnor U16196 (N_16196,N_15450,N_14118);
nand U16197 (N_16197,N_15649,N_14691);
nand U16198 (N_16198,N_14520,N_15241);
nor U16199 (N_16199,N_14736,N_14433);
nor U16200 (N_16200,N_14676,N_15738);
nor U16201 (N_16201,N_15793,N_14351);
or U16202 (N_16202,N_14660,N_14236);
nor U16203 (N_16203,N_14403,N_14111);
and U16204 (N_16204,N_15194,N_15341);
nor U16205 (N_16205,N_14456,N_14714);
xor U16206 (N_16206,N_14682,N_15084);
nand U16207 (N_16207,N_14165,N_15540);
xnor U16208 (N_16208,N_14062,N_15625);
xnor U16209 (N_16209,N_14959,N_15702);
or U16210 (N_16210,N_14415,N_14806);
and U16211 (N_16211,N_14133,N_14486);
and U16212 (N_16212,N_15359,N_15268);
nor U16213 (N_16213,N_14282,N_15276);
xor U16214 (N_16214,N_15841,N_14851);
nor U16215 (N_16215,N_15598,N_15075);
and U16216 (N_16216,N_15659,N_14426);
xor U16217 (N_16217,N_15446,N_15618);
nand U16218 (N_16218,N_14096,N_15573);
and U16219 (N_16219,N_14106,N_14754);
xor U16220 (N_16220,N_14518,N_15595);
nor U16221 (N_16221,N_14674,N_14102);
xnor U16222 (N_16222,N_14313,N_14757);
and U16223 (N_16223,N_14899,N_14480);
nand U16224 (N_16224,N_15483,N_15394);
or U16225 (N_16225,N_14364,N_15557);
nand U16226 (N_16226,N_15253,N_14462);
and U16227 (N_16227,N_14869,N_14298);
nand U16228 (N_16228,N_15972,N_15944);
or U16229 (N_16229,N_14457,N_14755);
nor U16230 (N_16230,N_15809,N_14956);
nand U16231 (N_16231,N_14750,N_15692);
xnor U16232 (N_16232,N_15842,N_14379);
and U16233 (N_16233,N_14226,N_14050);
nor U16234 (N_16234,N_14430,N_15848);
or U16235 (N_16235,N_15936,N_14941);
or U16236 (N_16236,N_15261,N_15155);
nand U16237 (N_16237,N_15286,N_15263);
nor U16238 (N_16238,N_15782,N_15236);
or U16239 (N_16239,N_14002,N_15689);
nand U16240 (N_16240,N_14041,N_14440);
and U16241 (N_16241,N_14333,N_15861);
or U16242 (N_16242,N_14803,N_14984);
xnor U16243 (N_16243,N_15294,N_14438);
nand U16244 (N_16244,N_14624,N_14598);
nand U16245 (N_16245,N_14965,N_15249);
and U16246 (N_16246,N_15434,N_15062);
nand U16247 (N_16247,N_14410,N_14824);
nand U16248 (N_16248,N_14978,N_14441);
nand U16249 (N_16249,N_15128,N_15821);
and U16250 (N_16250,N_14014,N_14488);
and U16251 (N_16251,N_14976,N_15851);
xnor U16252 (N_16252,N_14605,N_15904);
nor U16253 (N_16253,N_15707,N_15467);
nor U16254 (N_16254,N_14729,N_15087);
nand U16255 (N_16255,N_14540,N_14458);
nand U16256 (N_16256,N_14427,N_15392);
or U16257 (N_16257,N_14882,N_15278);
nand U16258 (N_16258,N_14122,N_15602);
xnor U16259 (N_16259,N_15476,N_14890);
or U16260 (N_16260,N_15956,N_14212);
nand U16261 (N_16261,N_14566,N_14986);
xor U16262 (N_16262,N_15018,N_15912);
or U16263 (N_16263,N_14989,N_15903);
nand U16264 (N_16264,N_14362,N_15999);
nor U16265 (N_16265,N_15801,N_14709);
nor U16266 (N_16266,N_15416,N_15739);
or U16267 (N_16267,N_14556,N_14328);
nand U16268 (N_16268,N_15069,N_15429);
nor U16269 (N_16269,N_14970,N_14920);
xnor U16270 (N_16270,N_15852,N_14253);
xor U16271 (N_16271,N_15072,N_15160);
nor U16272 (N_16272,N_14220,N_14123);
nand U16273 (N_16273,N_15709,N_14131);
xnor U16274 (N_16274,N_15711,N_14648);
nand U16275 (N_16275,N_15157,N_15035);
xor U16276 (N_16276,N_15036,N_15110);
nand U16277 (N_16277,N_14232,N_14278);
xnor U16278 (N_16278,N_15423,N_15780);
or U16279 (N_16279,N_14358,N_15161);
and U16280 (N_16280,N_15230,N_14935);
or U16281 (N_16281,N_14190,N_14529);
xor U16282 (N_16282,N_14468,N_14400);
xnor U16283 (N_16283,N_15153,N_14435);
nor U16284 (N_16284,N_15729,N_15537);
or U16285 (N_16285,N_15192,N_15547);
or U16286 (N_16286,N_14273,N_15866);
or U16287 (N_16287,N_14219,N_15503);
nand U16288 (N_16288,N_15144,N_14670);
nand U16289 (N_16289,N_15229,N_14700);
or U16290 (N_16290,N_14745,N_15960);
and U16291 (N_16291,N_15695,N_14807);
xor U16292 (N_16292,N_14856,N_14420);
nor U16293 (N_16293,N_14103,N_15317);
nor U16294 (N_16294,N_14545,N_15096);
or U16295 (N_16295,N_14161,N_14774);
nand U16296 (N_16296,N_15635,N_14315);
or U16297 (N_16297,N_14040,N_14105);
or U16298 (N_16298,N_15045,N_15056);
or U16299 (N_16299,N_15252,N_15882);
and U16300 (N_16300,N_14089,N_15383);
xor U16301 (N_16301,N_14320,N_15427);
xnor U16302 (N_16302,N_15384,N_14922);
nand U16303 (N_16303,N_15559,N_15701);
or U16304 (N_16304,N_15174,N_14814);
and U16305 (N_16305,N_15292,N_15457);
nor U16306 (N_16306,N_15741,N_14707);
and U16307 (N_16307,N_15313,N_15958);
or U16308 (N_16308,N_14181,N_14092);
and U16309 (N_16309,N_14237,N_14176);
nor U16310 (N_16310,N_15528,N_15590);
or U16311 (N_16311,N_15525,N_15825);
and U16312 (N_16312,N_15111,N_14292);
nand U16313 (N_16313,N_15009,N_15560);
xnor U16314 (N_16314,N_14577,N_15444);
or U16315 (N_16315,N_15977,N_15652);
or U16316 (N_16316,N_15507,N_15207);
xor U16317 (N_16317,N_15837,N_15319);
nor U16318 (N_16318,N_15524,N_14722);
nor U16319 (N_16319,N_14571,N_14780);
xor U16320 (N_16320,N_15813,N_15419);
or U16321 (N_16321,N_15209,N_15896);
nor U16322 (N_16322,N_14552,N_14561);
nand U16323 (N_16323,N_15445,N_15534);
and U16324 (N_16324,N_14506,N_14779);
and U16325 (N_16325,N_14078,N_15346);
or U16326 (N_16326,N_15973,N_15277);
or U16327 (N_16327,N_14859,N_15040);
xnor U16328 (N_16328,N_14568,N_15300);
or U16329 (N_16329,N_14338,N_15104);
xor U16330 (N_16330,N_14641,N_14416);
or U16331 (N_16331,N_15548,N_14618);
and U16332 (N_16332,N_14706,N_14542);
xor U16333 (N_16333,N_14916,N_15345);
xnor U16334 (N_16334,N_15599,N_15048);
and U16335 (N_16335,N_14209,N_14373);
or U16336 (N_16336,N_14756,N_15629);
or U16337 (N_16337,N_14272,N_15910);
nor U16338 (N_16338,N_14631,N_15238);
xnor U16339 (N_16339,N_15460,N_15219);
or U16340 (N_16340,N_15786,N_14322);
nand U16341 (N_16341,N_15050,N_14576);
and U16342 (N_16342,N_15760,N_14857);
and U16343 (N_16343,N_14546,N_14083);
nand U16344 (N_16344,N_14645,N_15182);
or U16345 (N_16345,N_14549,N_14419);
and U16346 (N_16346,N_15703,N_15061);
xor U16347 (N_16347,N_14469,N_14389);
or U16348 (N_16348,N_15171,N_14183);
nand U16349 (N_16349,N_15059,N_14789);
nand U16350 (N_16350,N_15715,N_15031);
and U16351 (N_16351,N_14252,N_15593);
or U16352 (N_16352,N_14000,N_14084);
nor U16353 (N_16353,N_14200,N_14032);
nor U16354 (N_16354,N_15280,N_15686);
and U16355 (N_16355,N_14622,N_15731);
nand U16356 (N_16356,N_14091,N_14595);
nor U16357 (N_16357,N_14126,N_15073);
or U16358 (N_16358,N_14153,N_15990);
nor U16359 (N_16359,N_14178,N_14490);
nor U16360 (N_16360,N_14235,N_14633);
or U16361 (N_16361,N_15271,N_15151);
and U16362 (N_16362,N_15762,N_15477);
or U16363 (N_16363,N_15099,N_14217);
xnor U16364 (N_16364,N_15927,N_14286);
and U16365 (N_16365,N_15862,N_15091);
nand U16366 (N_16366,N_15791,N_14910);
or U16367 (N_16367,N_14124,N_15466);
nor U16368 (N_16368,N_15044,N_15940);
and U16369 (N_16369,N_14285,N_14508);
and U16370 (N_16370,N_14088,N_15781);
or U16371 (N_16371,N_15225,N_14837);
nor U16372 (N_16372,N_14354,N_14726);
xor U16373 (N_16373,N_14553,N_15380);
or U16374 (N_16374,N_15399,N_15342);
or U16375 (N_16375,N_14346,N_15566);
and U16376 (N_16376,N_15361,N_14672);
or U16377 (N_16377,N_14481,N_14158);
xnor U16378 (N_16378,N_15131,N_15808);
nand U16379 (N_16379,N_15125,N_15982);
nor U16380 (N_16380,N_14634,N_14066);
xnor U16381 (N_16381,N_15175,N_14705);
or U16382 (N_16382,N_14277,N_14329);
xor U16383 (N_16383,N_14713,N_15938);
or U16384 (N_16384,N_15202,N_15260);
and U16385 (N_16385,N_15812,N_15900);
nand U16386 (N_16386,N_14664,N_14503);
nor U16387 (N_16387,N_15699,N_15105);
xnor U16388 (N_16388,N_14283,N_14746);
xnor U16389 (N_16389,N_15693,N_14461);
and U16390 (N_16390,N_15201,N_15665);
nand U16391 (N_16391,N_15232,N_15932);
or U16392 (N_16392,N_15107,N_15552);
or U16393 (N_16393,N_15946,N_14775);
nand U16394 (N_16394,N_14995,N_14818);
and U16395 (N_16395,N_14024,N_15212);
and U16396 (N_16396,N_15465,N_15403);
and U16397 (N_16397,N_15203,N_15242);
nor U16398 (N_16398,N_15382,N_15169);
and U16399 (N_16399,N_15647,N_14265);
xnor U16400 (N_16400,N_14581,N_15223);
and U16401 (N_16401,N_14493,N_15962);
xor U16402 (N_16402,N_14782,N_15082);
xor U16403 (N_16403,N_14611,N_14471);
or U16404 (N_16404,N_14449,N_14489);
nand U16405 (N_16405,N_15255,N_15964);
or U16406 (N_16406,N_15675,N_15957);
or U16407 (N_16407,N_14330,N_14369);
nand U16408 (N_16408,N_15533,N_15060);
nor U16409 (N_16409,N_14712,N_14431);
or U16410 (N_16410,N_14271,N_15270);
nand U16411 (N_16411,N_14610,N_14308);
and U16412 (N_16412,N_15459,N_15826);
or U16413 (N_16413,N_14239,N_15066);
nand U16414 (N_16414,N_14413,N_15287);
nor U16415 (N_16415,N_15757,N_14099);
nor U16416 (N_16416,N_14331,N_15704);
or U16417 (N_16417,N_15442,N_14340);
nor U16418 (N_16418,N_14831,N_15838);
and U16419 (N_16419,N_15240,N_15674);
nor U16420 (N_16420,N_14783,N_14699);
xnor U16421 (N_16421,N_14855,N_14304);
nor U16422 (N_16422,N_14478,N_15835);
xnor U16423 (N_16423,N_15777,N_15098);
or U16424 (N_16424,N_15579,N_15819);
and U16425 (N_16425,N_15281,N_14548);
or U16426 (N_16426,N_15208,N_15475);
nor U16427 (N_16427,N_15378,N_14525);
or U16428 (N_16428,N_15950,N_14725);
or U16429 (N_16429,N_14866,N_15706);
nand U16430 (N_16430,N_15070,N_14653);
xor U16431 (N_16431,N_14930,N_15764);
nor U16432 (N_16432,N_15425,N_14864);
nor U16433 (N_16433,N_14484,N_14819);
or U16434 (N_16434,N_15318,N_14195);
nand U16435 (N_16435,N_14828,N_14681);
nor U16436 (N_16436,N_14234,N_14477);
nor U16437 (N_16437,N_14685,N_14143);
nor U16438 (N_16438,N_14637,N_14460);
nor U16439 (N_16439,N_14663,N_15811);
nand U16440 (N_16440,N_15605,N_14094);
xor U16441 (N_16441,N_15463,N_15554);
xnor U16442 (N_16442,N_14917,N_14455);
nand U16443 (N_16443,N_15316,N_15544);
or U16444 (N_16444,N_15587,N_15604);
nand U16445 (N_16445,N_15293,N_14473);
and U16446 (N_16446,N_15615,N_14541);
and U16447 (N_16447,N_15749,N_15008);
nor U16448 (N_16448,N_14626,N_15471);
xor U16449 (N_16449,N_14025,N_15564);
xor U16450 (N_16450,N_14747,N_15140);
and U16451 (N_16451,N_15574,N_15441);
and U16452 (N_16452,N_15221,N_14035);
and U16453 (N_16453,N_14777,N_15054);
xnor U16454 (N_16454,N_14408,N_15085);
or U16455 (N_16455,N_14948,N_14361);
or U16456 (N_16456,N_14059,N_14950);
and U16457 (N_16457,N_14334,N_14215);
or U16458 (N_16458,N_15437,N_15181);
and U16459 (N_16459,N_15913,N_15197);
nand U16460 (N_16460,N_14428,N_15690);
and U16461 (N_16461,N_15798,N_14349);
and U16462 (N_16462,N_15732,N_14343);
and U16463 (N_16463,N_15258,N_15562);
nand U16464 (N_16464,N_15469,N_14380);
or U16465 (N_16465,N_14671,N_14760);
nand U16466 (N_16466,N_14110,N_15816);
and U16467 (N_16467,N_14302,N_14245);
nor U16468 (N_16468,N_14735,N_15109);
xnor U16469 (N_16469,N_14259,N_14832);
and U16470 (N_16470,N_14227,N_14138);
or U16471 (N_16471,N_15133,N_15484);
xnor U16472 (N_16472,N_15576,N_14968);
nor U16473 (N_16473,N_15325,N_15696);
nand U16474 (N_16474,N_15291,N_15078);
xor U16475 (N_16475,N_14701,N_15833);
xor U16476 (N_16476,N_15228,N_15730);
nor U16477 (N_16477,N_15756,N_14377);
xnor U16478 (N_16478,N_14197,N_15354);
and U16479 (N_16479,N_14790,N_15284);
nor U16480 (N_16480,N_15401,N_15132);
xor U16481 (N_16481,N_15988,N_14052);
nor U16482 (N_16482,N_14805,N_14100);
and U16483 (N_16483,N_15506,N_15997);
nand U16484 (N_16484,N_15733,N_15189);
and U16485 (N_16485,N_14532,N_15612);
xnor U16486 (N_16486,N_14731,N_14393);
nand U16487 (N_16487,N_14255,N_14309);
nand U16488 (N_16488,N_14823,N_14892);
nand U16489 (N_16489,N_15183,N_15660);
nor U16490 (N_16490,N_14009,N_15969);
and U16491 (N_16491,N_14872,N_14800);
nor U16492 (N_16492,N_15885,N_15915);
and U16493 (N_16493,N_15700,N_14778);
nor U16494 (N_16494,N_15186,N_15052);
nand U16495 (N_16495,N_14813,N_14840);
xnor U16496 (N_16496,N_14675,N_14130);
and U16497 (N_16497,N_15370,N_14987);
nor U16498 (N_16498,N_15330,N_14752);
nand U16499 (N_16499,N_14240,N_14597);
or U16500 (N_16500,N_14698,N_14804);
or U16501 (N_16501,N_15295,N_15385);
or U16502 (N_16502,N_14894,N_14749);
and U16503 (N_16503,N_14276,N_15767);
nor U16504 (N_16504,N_14401,N_15871);
xor U16505 (N_16505,N_14563,N_14307);
or U16506 (N_16506,N_14168,N_15563);
or U16507 (N_16507,N_15299,N_15518);
and U16508 (N_16508,N_15017,N_15120);
nor U16509 (N_16509,N_15978,N_14244);
nor U16510 (N_16510,N_14977,N_15875);
xor U16511 (N_16511,N_14873,N_14710);
xnor U16512 (N_16512,N_15943,N_14360);
nand U16513 (N_16513,N_14652,N_15565);
xor U16514 (N_16514,N_14248,N_14768);
xor U16515 (N_16515,N_15698,N_14937);
and U16516 (N_16516,N_14053,N_15398);
and U16517 (N_16517,N_15020,N_15919);
xor U16518 (N_16518,N_14319,N_14144);
nor U16519 (N_16519,N_15549,N_14932);
nor U16520 (N_16520,N_15898,N_15283);
and U16521 (N_16521,N_14904,N_15641);
nand U16522 (N_16522,N_15513,N_15480);
or U16523 (N_16523,N_14085,N_15763);
and U16524 (N_16524,N_15577,N_14281);
and U16525 (N_16525,N_14347,N_15472);
nor U16526 (N_16526,N_14792,N_15931);
nand U16527 (N_16527,N_14877,N_14258);
xnor U16528 (N_16528,N_15892,N_15247);
nor U16529 (N_16529,N_15296,N_15748);
xnor U16530 (N_16530,N_14528,N_15374);
nand U16531 (N_16531,N_15134,N_15123);
xnor U16532 (N_16532,N_15391,N_15770);
nor U16533 (N_16533,N_14500,N_15923);
and U16534 (N_16534,N_14799,N_15080);
xnor U16535 (N_16535,N_14210,N_15077);
xor U16536 (N_16536,N_14724,N_15307);
nand U16537 (N_16537,N_14424,N_14927);
nor U16538 (N_16538,N_15164,N_14575);
nand U16539 (N_16539,N_15705,N_14679);
nand U16540 (N_16540,N_15130,N_14359);
nand U16541 (N_16541,N_14274,N_15979);
xnor U16542 (N_16542,N_15769,N_15188);
and U16543 (N_16543,N_14381,N_14604);
or U16544 (N_16544,N_14291,N_14064);
nor U16545 (N_16545,N_15531,N_15558);
or U16546 (N_16546,N_14983,N_14101);
nand U16547 (N_16547,N_15492,N_15288);
nand U16548 (N_16548,N_15139,N_14981);
and U16549 (N_16549,N_14001,N_14125);
nor U16550 (N_16550,N_15408,N_14398);
and U16551 (N_16551,N_15512,N_14250);
nand U16552 (N_16552,N_14027,N_14046);
nor U16553 (N_16553,N_15794,N_15584);
or U16554 (N_16554,N_14483,N_14097);
or U16555 (N_16555,N_15400,N_14345);
and U16556 (N_16556,N_14936,N_14788);
or U16557 (N_16557,N_15339,N_15063);
xor U16558 (N_16558,N_14833,N_15343);
or U16559 (N_16559,N_15129,N_14365);
xnor U16560 (N_16560,N_14371,N_15245);
xor U16561 (N_16561,N_14912,N_15872);
and U16562 (N_16562,N_14198,N_14357);
and U16563 (N_16563,N_15822,N_15929);
nand U16564 (N_16564,N_14880,N_15362);
nand U16565 (N_16565,N_14898,N_15344);
and U16566 (N_16566,N_15895,N_15685);
nand U16567 (N_16567,N_14223,N_14771);
and U16568 (N_16568,N_14764,N_14058);
nand U16569 (N_16569,N_14485,N_15264);
xor U16570 (N_16570,N_15326,N_14697);
nor U16571 (N_16571,N_14213,N_15306);
nor U16572 (N_16572,N_15218,N_14399);
xnor U16573 (N_16573,N_14142,N_14661);
xor U16574 (N_16574,N_15971,N_15664);
and U16575 (N_16575,N_14554,N_14169);
xnor U16576 (N_16576,N_14817,N_14402);
xnor U16577 (N_16577,N_14603,N_15628);
and U16578 (N_16578,N_14573,N_15357);
nor U16579 (N_16579,N_14786,N_14376);
nand U16580 (N_16580,N_14031,N_14822);
nor U16581 (N_16581,N_15473,N_14425);
or U16582 (N_16582,N_14026,N_14472);
nor U16583 (N_16583,N_15662,N_15984);
xor U16584 (N_16584,N_14955,N_14878);
or U16585 (N_16585,N_14311,N_15414);
or U16586 (N_16586,N_15170,N_15007);
xnor U16587 (N_16587,N_15928,N_14012);
or U16588 (N_16588,N_14136,N_14414);
and U16589 (N_16589,N_14523,N_14908);
nor U16590 (N_16590,N_14842,N_14971);
or U16591 (N_16591,N_14196,N_14678);
or U16592 (N_16592,N_15933,N_14926);
or U16593 (N_16593,N_15830,N_14154);
nand U16594 (N_16594,N_14996,N_15839);
nor U16595 (N_16595,N_14112,N_14839);
nand U16596 (N_16596,N_14350,N_14246);
nor U16597 (N_16597,N_14228,N_14429);
or U16598 (N_16598,N_14268,N_15827);
xor U16599 (N_16599,N_15388,N_14476);
nor U16600 (N_16600,N_14923,N_15086);
nand U16601 (N_16601,N_14409,N_15254);
nor U16602 (N_16602,N_14991,N_14870);
nand U16603 (N_16603,N_15449,N_14972);
and U16604 (N_16604,N_14662,N_15451);
nand U16605 (N_16605,N_14513,N_14623);
nor U16606 (N_16606,N_14728,N_14879);
nor U16607 (N_16607,N_15156,N_15329);
nor U16608 (N_16608,N_15766,N_15849);
nor U16609 (N_16609,N_14295,N_15868);
xnor U16610 (N_16610,N_15027,N_15415);
or U16611 (N_16611,N_15015,N_14781);
xnor U16612 (N_16612,N_14045,N_15677);
nand U16613 (N_16613,N_14352,N_15336);
nor U16614 (N_16614,N_14221,N_14421);
or U16615 (N_16615,N_15796,N_15667);
or U16616 (N_16616,N_14619,N_15925);
xor U16617 (N_16617,N_15937,N_15055);
or U16618 (N_16618,N_15083,N_15421);
and U16619 (N_16619,N_14405,N_14843);
nor U16620 (N_16620,N_15723,N_14115);
or U16621 (N_16621,N_15177,N_14443);
or U16622 (N_16622,N_14562,N_14861);
nand U16623 (N_16623,N_15393,N_15214);
or U16624 (N_16624,N_14665,N_15614);
nor U16625 (N_16625,N_15987,N_14583);
nor U16626 (N_16626,N_14796,N_15146);
nor U16627 (N_16627,N_14584,N_14207);
nand U16628 (N_16628,N_14654,N_15775);
or U16629 (N_16629,N_15262,N_14275);
or U16630 (N_16630,N_15002,N_14086);
nand U16631 (N_16631,N_15350,N_14189);
or U16632 (N_16632,N_14858,N_15887);
nor U16633 (N_16633,N_15543,N_15924);
xnor U16634 (N_16634,N_15601,N_15859);
or U16635 (N_16635,N_15539,N_15353);
and U16636 (N_16636,N_14466,N_14057);
and U16637 (N_16637,N_15409,N_15850);
xnor U16638 (N_16638,N_15068,N_15805);
xor U16639 (N_16639,N_14586,N_14838);
xor U16640 (N_16640,N_14411,N_15025);
and U16641 (N_16641,N_14075,N_14022);
xnor U16642 (N_16642,N_14289,N_15092);
nor U16643 (N_16643,N_15149,N_14018);
nand U16644 (N_16644,N_14884,N_14098);
nand U16645 (N_16645,N_14335,N_15038);
or U16646 (N_16646,N_14853,N_14769);
and U16647 (N_16647,N_15064,N_15112);
nand U16648 (N_16648,N_15216,N_15784);
and U16649 (N_16649,N_14120,N_14751);
xor U16650 (N_16650,N_14164,N_15949);
nor U16651 (N_16651,N_15575,N_15752);
nand U16652 (N_16652,N_14572,N_15787);
nand U16653 (N_16653,N_14905,N_14964);
or U16654 (N_16654,N_14614,N_14966);
or U16655 (N_16655,N_14740,N_14687);
and U16656 (N_16656,N_15000,N_15759);
nor U16657 (N_16657,N_14384,N_15024);
nand U16658 (N_16658,N_15371,N_14254);
nor U16659 (N_16659,N_15389,N_14262);
nand U16660 (N_16660,N_14267,N_15671);
nor U16661 (N_16661,N_14060,N_15561);
xnor U16662 (N_16662,N_14704,N_15893);
or U16663 (N_16663,N_14011,N_15654);
and U16664 (N_16664,N_14230,N_15498);
or U16665 (N_16665,N_15154,N_15863);
nor U16666 (N_16666,N_14224,N_14711);
nand U16667 (N_16667,N_14450,N_14512);
and U16668 (N_16668,N_15315,N_15282);
or U16669 (N_16669,N_15582,N_14793);
or U16670 (N_16670,N_15148,N_15670);
and U16671 (N_16671,N_15637,N_14909);
nor U16672 (N_16672,N_15721,N_15220);
xor U16673 (N_16673,N_15179,N_14184);
xor U16674 (N_16674,N_14632,N_15323);
nor U16675 (N_16675,N_15555,N_14815);
nor U16676 (N_16676,N_15765,N_15406);
nor U16677 (N_16677,N_15352,N_15375);
or U16678 (N_16678,N_14809,N_15504);
nor U16679 (N_16679,N_14802,N_15921);
and U16680 (N_16680,N_14061,N_15745);
xnor U16681 (N_16681,N_15373,N_14980);
nand U16682 (N_16682,N_15743,N_15333);
and U16683 (N_16683,N_15418,N_14152);
and U16684 (N_16684,N_15079,N_15980);
and U16685 (N_16685,N_15883,N_15855);
or U16686 (N_16686,N_14515,N_14497);
nand U16687 (N_16687,N_15551,N_15858);
nand U16688 (N_16688,N_14021,N_15658);
or U16689 (N_16689,N_14943,N_14721);
nor U16690 (N_16690,N_14748,N_15627);
and U16691 (N_16691,N_14688,N_14812);
or U16692 (N_16692,N_15122,N_14470);
or U16693 (N_16693,N_15239,N_15039);
nor U16694 (N_16694,N_15407,N_14640);
and U16695 (N_16695,N_14913,N_15669);
nand U16696 (N_16696,N_15905,N_14850);
nand U16697 (N_16697,N_14356,N_15447);
or U16698 (N_16698,N_14875,N_14992);
or U16699 (N_16699,N_14784,N_14023);
xnor U16700 (N_16700,N_14835,N_15714);
nor U16701 (N_16701,N_15051,N_14593);
xnor U16702 (N_16702,N_15163,N_15269);
nand U16703 (N_16703,N_14929,N_15314);
and U16704 (N_16704,N_14260,N_15158);
xor U16705 (N_16705,N_15493,N_15049);
xnor U16706 (N_16706,N_15251,N_14891);
xor U16707 (N_16707,N_14113,N_14116);
or U16708 (N_16708,N_15211,N_14266);
nor U16709 (N_16709,N_15541,N_14332);
xor U16710 (N_16710,N_15363,N_14791);
nand U16711 (N_16711,N_14743,N_14715);
nor U16712 (N_16712,N_15653,N_15206);
or U16713 (N_16713,N_15804,N_14149);
nand U16714 (N_16714,N_15623,N_15114);
nor U16715 (N_16715,N_15369,N_14039);
nand U16716 (N_16716,N_15510,N_14876);
xor U16717 (N_16717,N_15981,N_15716);
nand U16718 (N_16718,N_14974,N_15103);
and U16719 (N_16719,N_15679,N_15634);
nor U16720 (N_16720,N_15886,N_14559);
or U16721 (N_16721,N_15536,N_14536);
nor U16722 (N_16722,N_14569,N_14229);
and U16723 (N_16723,N_15440,N_14609);
or U16724 (N_16724,N_15996,N_15113);
or U16725 (N_16725,N_14821,N_15093);
and U16726 (N_16726,N_14336,N_14263);
xnor U16727 (N_16727,N_14206,N_14072);
or U16728 (N_16728,N_15783,N_15355);
nand U16729 (N_16729,N_15289,N_15663);
xor U16730 (N_16730,N_15136,N_15119);
nor U16731 (N_16731,N_14733,N_15650);
nor U16732 (N_16732,N_15529,N_15198);
nand U16733 (N_16733,N_15081,N_14397);
and U16734 (N_16734,N_14208,N_15452);
or U16735 (N_16735,N_15022,N_15267);
nor U16736 (N_16736,N_15708,N_15489);
xor U16737 (N_16737,N_15867,N_15348);
nor U16738 (N_16738,N_14507,N_14499);
nor U16739 (N_16739,N_14647,N_14296);
or U16740 (N_16740,N_15916,N_15834);
and U16741 (N_16741,N_15624,N_15591);
and U16742 (N_16742,N_15611,N_15166);
xnor U16743 (N_16743,N_15482,N_15067);
xor U16744 (N_16744,N_15844,N_14243);
or U16745 (N_16745,N_14973,N_14739);
xnor U16746 (N_16746,N_14847,N_14241);
xnor U16747 (N_16747,N_15795,N_14117);
nand U16748 (N_16748,N_15952,N_15568);
nor U16749 (N_16749,N_15845,N_15479);
or U16750 (N_16750,N_14547,N_15874);
nor U16751 (N_16751,N_14621,N_15074);
and U16752 (N_16752,N_14504,N_15758);
or U16753 (N_16753,N_15168,N_14534);
nor U16754 (N_16754,N_14188,N_14327);
nor U16755 (N_16755,N_14558,N_14762);
or U16756 (N_16756,N_15556,N_15840);
and U16757 (N_16757,N_14982,N_14578);
nand U16758 (N_16758,N_15274,N_14137);
xnor U16759 (N_16759,N_14093,N_15788);
or U16760 (N_16760,N_14201,N_14616);
or U16761 (N_16761,N_14938,N_15792);
or U16762 (N_16762,N_15747,N_14988);
or U16763 (N_16763,N_14734,N_15126);
nor U16764 (N_16764,N_15327,N_15490);
and U16765 (N_16765,N_14172,N_15908);
or U16766 (N_16766,N_14538,N_15735);
xor U16767 (N_16767,N_14785,N_15453);
nand U16768 (N_16768,N_14599,N_14630);
nand U16769 (N_16769,N_15986,N_15402);
and U16770 (N_16770,N_15310,N_15290);
nand U16771 (N_16771,N_14388,N_14551);
xnor U16772 (N_16772,N_15509,N_15516);
xor U16773 (N_16773,N_15273,N_14606);
xor U16774 (N_16774,N_14742,N_14303);
xor U16775 (N_16775,N_14940,N_15870);
or U16776 (N_16776,N_14703,N_14155);
nand U16777 (N_16777,N_14590,N_15578);
and U16778 (N_16778,N_15753,N_15818);
nand U16779 (N_16779,N_14132,N_14418);
and U16780 (N_16780,N_15364,N_15609);
xor U16781 (N_16781,N_15487,N_15322);
and U16782 (N_16782,N_15331,N_15030);
nor U16783 (N_16783,N_15613,N_14326);
xnor U16784 (N_16784,N_15880,N_14048);
or U16785 (N_16785,N_14020,N_14741);
nand U16786 (N_16786,N_14056,N_14087);
or U16787 (N_16787,N_15410,N_15443);
nand U16788 (N_16788,N_15522,N_14444);
nand U16789 (N_16789,N_15412,N_15320);
and U16790 (N_16790,N_14166,N_14643);
xnor U16791 (N_16791,N_15620,N_15736);
and U16792 (N_16792,N_15603,N_14321);
and U16793 (N_16793,N_14985,N_15349);
nand U16794 (N_16794,N_15481,N_14535);
and U16795 (N_16795,N_15909,N_15013);
nand U16796 (N_16796,N_14667,N_15724);
or U16797 (N_16797,N_15167,N_15691);
and U16798 (N_16798,N_14355,N_14325);
and U16799 (N_16799,N_15687,N_15303);
nor U16800 (N_16800,N_15717,N_14531);
and U16801 (N_16801,N_14407,N_15432);
or U16802 (N_16802,N_14366,N_14753);
nor U16803 (N_16803,N_15520,N_15433);
xor U16804 (N_16804,N_14776,N_15185);
nor U16805 (N_16805,N_15740,N_15719);
or U16806 (N_16806,N_14432,N_15005);
and U16807 (N_16807,N_15461,N_14417);
and U16808 (N_16808,N_15265,N_15358);
or U16809 (N_16809,N_14300,N_15118);
nor U16810 (N_16810,N_14613,N_15088);
and U16811 (N_16811,N_14006,N_14279);
or U16812 (N_16812,N_15321,N_15396);
or U16813 (N_16813,N_14716,N_15023);
or U16814 (N_16814,N_15572,N_15911);
nor U16815 (N_16815,N_15058,N_15589);
xor U16816 (N_16816,N_14708,N_15191);
or U16817 (N_16817,N_15379,N_14766);
nor U16818 (N_16818,N_15491,N_14090);
nand U16819 (N_16819,N_14251,N_14635);
nor U16820 (N_16820,N_14767,N_15012);
nand U16821 (N_16821,N_14820,N_15935);
xor U16822 (N_16822,N_14495,N_14387);
xnor U16823 (N_16823,N_14043,N_15332);
xor U16824 (N_16824,N_15210,N_14656);
nor U16825 (N_16825,N_14049,N_14591);
and U16826 (N_16826,N_14339,N_15065);
nor U16827 (N_16827,N_15610,N_15947);
and U16828 (N_16828,N_14555,N_15600);
or U16829 (N_16829,N_15121,N_15897);
and U16830 (N_16830,N_15356,N_14732);
or U16831 (N_16831,N_15094,N_15683);
nor U16832 (N_16832,N_15159,N_14772);
xor U16833 (N_16833,N_14510,N_15532);
xnor U16834 (N_16834,N_14934,N_14249);
xnor U16835 (N_16835,N_14644,N_15884);
and U16836 (N_16836,N_15823,N_15337);
nand U16837 (N_16837,N_15942,N_14492);
nand U16838 (N_16838,N_15360,N_15820);
xnor U16839 (N_16839,N_14487,N_15810);
nand U16840 (N_16840,N_15789,N_15646);
and U16841 (N_16841,N_14657,N_15100);
and U16842 (N_16842,N_14037,N_15338);
and U16843 (N_16843,N_14003,N_15413);
xor U16844 (N_16844,N_15586,N_14659);
and U16845 (N_16845,N_14810,N_15495);
xor U16846 (N_16846,N_14808,N_14702);
or U16847 (N_16847,N_15968,N_14602);
xnor U16848 (N_16848,N_14689,N_14564);
and U16849 (N_16849,N_15488,N_15003);
nor U16850 (N_16850,N_14526,N_15244);
and U16851 (N_16851,N_14600,N_15439);
xnor U16852 (N_16852,N_14928,N_15710);
nor U16853 (N_16853,N_14231,N_14816);
and U16854 (N_16854,N_15535,N_15275);
and U16855 (N_16855,N_14284,N_14293);
and U16856 (N_16856,N_15279,N_14305);
xor U16857 (N_16857,N_15814,N_14830);
or U16858 (N_16858,N_14692,N_15815);
nor U16859 (N_16859,N_15527,N_15588);
and U16860 (N_16860,N_14017,N_15643);
nor U16861 (N_16861,N_14658,N_14082);
xor U16862 (N_16862,N_14773,N_15235);
xnor U16863 (N_16863,N_14108,N_14642);
or U16864 (N_16864,N_15831,N_14306);
xnor U16865 (N_16865,N_14180,N_15594);
nand U16866 (N_16866,N_14128,N_14374);
nand U16867 (N_16867,N_15922,N_15891);
nor U16868 (N_16868,N_14070,N_15199);
and U16869 (N_16869,N_15746,N_15334);
xor U16870 (N_16870,N_14238,N_14516);
or U16871 (N_16871,N_14445,N_14501);
nand U16872 (N_16872,N_15309,N_15860);
or U16873 (N_16873,N_14434,N_14834);
nand U16874 (N_16874,N_14299,N_15250);
nor U16875 (N_16875,N_14016,N_14378);
and U16876 (N_16876,N_15843,N_15145);
nand U16877 (N_16877,N_14194,N_15376);
and U16878 (N_16878,N_14280,N_14071);
nor U16879 (N_16879,N_14395,N_14719);
nand U16880 (N_16880,N_14385,N_15335);
xnor U16881 (N_16881,N_15644,N_14921);
nand U16882 (N_16882,N_14129,N_15967);
nand U16883 (N_16883,N_14175,N_14919);
and U16884 (N_16884,N_15926,N_14005);
or U16885 (N_16885,N_14787,N_14370);
nor U16886 (N_16886,N_14537,N_14312);
or U16887 (N_16887,N_15143,N_14114);
nor U16888 (N_16888,N_15607,N_15545);
or U16889 (N_16889,N_14496,N_14801);
xnor U16890 (N_16890,N_15124,N_15751);
nand U16891 (N_16891,N_15237,N_15205);
xor U16892 (N_16892,N_15542,N_15873);
xnor U16893 (N_16893,N_15053,N_15162);
or U16894 (N_16894,N_15117,N_14318);
or U16895 (N_16895,N_15768,N_15424);
nand U16896 (N_16896,N_15998,N_14521);
and U16897 (N_16897,N_15718,N_14191);
and U16898 (N_16898,N_15608,N_15135);
nor U16899 (N_16899,N_15042,N_14055);
and U16900 (N_16900,N_14270,N_15266);
or U16901 (N_16901,N_14939,N_14139);
xnor U16902 (N_16902,N_15865,N_14944);
nand U16903 (N_16903,N_15945,N_15639);
nor U16904 (N_16904,N_15722,N_15195);
or U16905 (N_16905,N_15951,N_15991);
and U16906 (N_16906,N_14107,N_15215);
xnor U16907 (N_16907,N_14054,N_14436);
and U16908 (N_16908,N_14730,N_15941);
xnor U16909 (N_16909,N_15019,N_14437);
and U16910 (N_16910,N_14954,N_15304);
or U16911 (N_16911,N_15496,N_15853);
nand U16912 (N_16912,N_15680,N_14297);
nor U16913 (N_16913,N_14127,N_15720);
nand U16914 (N_16914,N_15138,N_15727);
nand U16915 (N_16915,N_14686,N_15626);
xor U16916 (N_16916,N_15298,N_15656);
nor U16917 (N_16917,N_14907,N_15906);
nand U16918 (N_16918,N_15771,N_14607);
xor U16919 (N_16919,N_14717,N_15187);
xnor U16920 (N_16920,N_14863,N_14579);
xnor U16921 (N_16921,N_15569,N_14015);
and U16922 (N_16922,N_14931,N_15581);
or U16923 (N_16923,N_14174,N_14646);
and U16924 (N_16924,N_15328,N_14897);
nor U16925 (N_16925,N_14868,N_15351);
xnor U16926 (N_16926,N_15954,N_15468);
nand U16927 (N_16927,N_15797,N_15800);
xor U16928 (N_16928,N_14846,N_15390);
nand U16929 (N_16929,N_14095,N_14889);
or U16930 (N_16930,N_15340,N_15580);
nor U16931 (N_16931,N_14396,N_14649);
xor U16932 (N_16932,N_14557,N_15894);
and U16933 (N_16933,N_15200,N_15799);
and U16934 (N_16934,N_15877,N_14317);
nor U16935 (N_16935,N_15953,N_14798);
and U16936 (N_16936,N_15367,N_15737);
nand U16937 (N_16937,N_15989,N_14162);
and U16938 (N_16938,N_14372,N_14185);
and U16939 (N_16939,N_15790,N_14946);
and U16940 (N_16940,N_14134,N_14065);
nor U16941 (N_16941,N_15500,N_15454);
nor U16942 (N_16942,N_14170,N_15173);
xor U16943 (N_16943,N_15776,N_15661);
nand U16944 (N_16944,N_14269,N_15001);
nand U16945 (N_16945,N_14423,N_15697);
xnor U16946 (N_16946,N_15514,N_15959);
nand U16947 (N_16947,N_15890,N_15684);
nor U16948 (N_16948,N_14900,N_14952);
nand U16949 (N_16949,N_14150,N_15474);
and U16950 (N_16950,N_14464,N_14007);
nor U16951 (N_16951,N_15596,N_15754);
and U16952 (N_16952,N_15750,N_14902);
nor U16953 (N_16953,N_14179,N_15176);
nor U16954 (N_16954,N_14519,N_14589);
or U16955 (N_16955,N_15617,N_15571);
xnor U16956 (N_16956,N_14867,N_14844);
nor U16957 (N_16957,N_14077,N_14639);
xnor U16958 (N_16958,N_15864,N_14565);
or U16959 (N_16959,N_14459,N_14765);
and U16960 (N_16960,N_15994,N_14770);
nor U16961 (N_16961,N_14620,N_14121);
or U16962 (N_16962,N_15272,N_14933);
or U16963 (N_16963,N_15901,N_14104);
or U16964 (N_16964,N_15365,N_15386);
and U16965 (N_16965,N_14348,N_14257);
or U16966 (N_16966,N_14677,N_14448);
nor U16967 (N_16967,N_14585,N_14033);
and U16968 (N_16968,N_15395,N_14446);
nand U16969 (N_16969,N_15233,N_14683);
xor U16970 (N_16970,N_15918,N_15976);
nand U16971 (N_16971,N_14028,N_14881);
or U16972 (N_16972,N_15519,N_14160);
nor U16973 (N_16973,N_15246,N_15150);
nor U16974 (N_16974,N_15204,N_14680);
nand U16975 (N_16975,N_15678,N_15934);
and U16976 (N_16976,N_14498,N_15097);
xnor U16977 (N_16977,N_14925,N_15248);
and U16978 (N_16978,N_15917,N_15196);
xor U16979 (N_16979,N_14795,N_14794);
and U16980 (N_16980,N_15570,N_14601);
nand U16981 (N_16981,N_14567,N_15497);
or U16982 (N_16982,N_14570,N_14530);
nor U16983 (N_16983,N_14404,N_15311);
nor U16984 (N_16984,N_14008,N_15948);
nor U16985 (N_16985,N_14063,N_14079);
xor U16986 (N_16986,N_15016,N_14225);
or U16987 (N_16987,N_14883,N_14186);
or U16988 (N_16988,N_14442,N_14960);
and U16989 (N_16989,N_15302,N_15033);
and U16990 (N_16990,N_15993,N_14182);
and U16991 (N_16991,N_14865,N_15417);
nand U16992 (N_16992,N_14394,N_15217);
xor U16993 (N_16993,N_14067,N_14896);
or U16994 (N_16994,N_15485,N_15458);
or U16995 (N_16995,N_14167,N_15301);
nor U16996 (N_16996,N_15324,N_15742);
nand U16997 (N_16997,N_14574,N_15778);
nor U16998 (N_16998,N_14949,N_14247);
nand U16999 (N_16999,N_14582,N_15550);
and U17000 (N_17000,N_14329,N_15300);
nor U17001 (N_17001,N_15075,N_14018);
xnor U17002 (N_17002,N_15273,N_14159);
nand U17003 (N_17003,N_14449,N_15893);
nand U17004 (N_17004,N_14088,N_15192);
or U17005 (N_17005,N_14147,N_14345);
xnor U17006 (N_17006,N_15070,N_15911);
xor U17007 (N_17007,N_15098,N_14051);
and U17008 (N_17008,N_14379,N_14684);
or U17009 (N_17009,N_14498,N_15949);
nand U17010 (N_17010,N_15856,N_15548);
xor U17011 (N_17011,N_14698,N_15760);
nor U17012 (N_17012,N_15462,N_15102);
and U17013 (N_17013,N_14631,N_14124);
xor U17014 (N_17014,N_14074,N_14851);
and U17015 (N_17015,N_14066,N_15738);
xnor U17016 (N_17016,N_14114,N_14107);
nand U17017 (N_17017,N_15448,N_14602);
or U17018 (N_17018,N_15847,N_15884);
nand U17019 (N_17019,N_15354,N_14328);
nand U17020 (N_17020,N_14057,N_15761);
or U17021 (N_17021,N_14781,N_15287);
xor U17022 (N_17022,N_15709,N_15486);
nor U17023 (N_17023,N_15870,N_14059);
nor U17024 (N_17024,N_14135,N_15721);
nand U17025 (N_17025,N_15886,N_15306);
nor U17026 (N_17026,N_15894,N_15752);
nor U17027 (N_17027,N_15681,N_14630);
and U17028 (N_17028,N_15630,N_14788);
and U17029 (N_17029,N_15691,N_15266);
nor U17030 (N_17030,N_15703,N_15834);
nor U17031 (N_17031,N_15247,N_14914);
xor U17032 (N_17032,N_15382,N_15110);
and U17033 (N_17033,N_15786,N_15217);
nand U17034 (N_17034,N_14813,N_15141);
or U17035 (N_17035,N_15651,N_14446);
or U17036 (N_17036,N_14625,N_15947);
xnor U17037 (N_17037,N_14257,N_14835);
nor U17038 (N_17038,N_15168,N_15007);
or U17039 (N_17039,N_14254,N_14577);
nor U17040 (N_17040,N_15305,N_14145);
and U17041 (N_17041,N_15658,N_14856);
nor U17042 (N_17042,N_15093,N_14136);
xnor U17043 (N_17043,N_14265,N_14300);
or U17044 (N_17044,N_15390,N_15575);
and U17045 (N_17045,N_14100,N_14284);
nor U17046 (N_17046,N_15745,N_14841);
or U17047 (N_17047,N_14111,N_15752);
and U17048 (N_17048,N_14347,N_15228);
nor U17049 (N_17049,N_15196,N_15979);
or U17050 (N_17050,N_14134,N_15428);
nand U17051 (N_17051,N_15257,N_15481);
and U17052 (N_17052,N_15274,N_15437);
xor U17053 (N_17053,N_14305,N_14586);
and U17054 (N_17054,N_14513,N_14953);
nand U17055 (N_17055,N_15809,N_15539);
nor U17056 (N_17056,N_14616,N_14497);
xor U17057 (N_17057,N_15461,N_15650);
and U17058 (N_17058,N_15282,N_15343);
or U17059 (N_17059,N_15886,N_15447);
or U17060 (N_17060,N_15297,N_14966);
or U17061 (N_17061,N_15655,N_14014);
or U17062 (N_17062,N_14277,N_15400);
xnor U17063 (N_17063,N_15219,N_15221);
nor U17064 (N_17064,N_14365,N_14499);
nor U17065 (N_17065,N_15487,N_14984);
nand U17066 (N_17066,N_15822,N_15268);
xnor U17067 (N_17067,N_14840,N_15432);
and U17068 (N_17068,N_15656,N_15508);
nor U17069 (N_17069,N_14447,N_15510);
and U17070 (N_17070,N_15408,N_15494);
and U17071 (N_17071,N_14683,N_15467);
nor U17072 (N_17072,N_15222,N_15826);
xor U17073 (N_17073,N_15018,N_15236);
or U17074 (N_17074,N_14548,N_14164);
or U17075 (N_17075,N_14964,N_14401);
nor U17076 (N_17076,N_14285,N_15172);
nor U17077 (N_17077,N_14114,N_14984);
or U17078 (N_17078,N_15696,N_14779);
and U17079 (N_17079,N_14886,N_14340);
nand U17080 (N_17080,N_15290,N_14067);
nor U17081 (N_17081,N_15984,N_15061);
nand U17082 (N_17082,N_15562,N_14633);
nor U17083 (N_17083,N_14223,N_15587);
and U17084 (N_17084,N_14952,N_14820);
nor U17085 (N_17085,N_14318,N_14440);
xor U17086 (N_17086,N_14233,N_14419);
xor U17087 (N_17087,N_15627,N_14970);
or U17088 (N_17088,N_14807,N_15082);
xnor U17089 (N_17089,N_15569,N_15962);
nor U17090 (N_17090,N_15027,N_14461);
or U17091 (N_17091,N_15589,N_15700);
or U17092 (N_17092,N_14105,N_14186);
nand U17093 (N_17093,N_15306,N_15911);
and U17094 (N_17094,N_14296,N_14248);
and U17095 (N_17095,N_14932,N_14486);
nor U17096 (N_17096,N_15165,N_14646);
or U17097 (N_17097,N_14130,N_15718);
nand U17098 (N_17098,N_14842,N_14834);
and U17099 (N_17099,N_14920,N_14230);
and U17100 (N_17100,N_15240,N_14020);
xnor U17101 (N_17101,N_15826,N_15580);
and U17102 (N_17102,N_15497,N_14968);
or U17103 (N_17103,N_14907,N_14654);
xnor U17104 (N_17104,N_14231,N_15166);
and U17105 (N_17105,N_14508,N_15580);
or U17106 (N_17106,N_15620,N_15819);
and U17107 (N_17107,N_14389,N_15428);
or U17108 (N_17108,N_15276,N_14994);
xnor U17109 (N_17109,N_14938,N_15530);
or U17110 (N_17110,N_14713,N_15628);
nand U17111 (N_17111,N_14862,N_14657);
and U17112 (N_17112,N_14223,N_14135);
or U17113 (N_17113,N_15221,N_15563);
and U17114 (N_17114,N_14048,N_15038);
nor U17115 (N_17115,N_15418,N_15176);
nand U17116 (N_17116,N_15195,N_15827);
nand U17117 (N_17117,N_15963,N_15351);
xnor U17118 (N_17118,N_14609,N_15510);
nand U17119 (N_17119,N_14950,N_14021);
nor U17120 (N_17120,N_15143,N_15716);
nand U17121 (N_17121,N_14997,N_15375);
xnor U17122 (N_17122,N_15765,N_15092);
or U17123 (N_17123,N_14329,N_15371);
or U17124 (N_17124,N_14819,N_14329);
and U17125 (N_17125,N_14532,N_14167);
nor U17126 (N_17126,N_14748,N_14572);
and U17127 (N_17127,N_15914,N_15806);
nand U17128 (N_17128,N_14488,N_15699);
nand U17129 (N_17129,N_14366,N_15217);
nand U17130 (N_17130,N_14723,N_15905);
and U17131 (N_17131,N_15275,N_15169);
or U17132 (N_17132,N_14903,N_15957);
and U17133 (N_17133,N_15401,N_14350);
or U17134 (N_17134,N_15284,N_14904);
nand U17135 (N_17135,N_15609,N_15150);
nand U17136 (N_17136,N_15652,N_15342);
nand U17137 (N_17137,N_14793,N_15687);
and U17138 (N_17138,N_14496,N_14189);
and U17139 (N_17139,N_15569,N_15922);
nor U17140 (N_17140,N_14341,N_15989);
and U17141 (N_17141,N_15799,N_15817);
nand U17142 (N_17142,N_15099,N_15899);
and U17143 (N_17143,N_14351,N_14932);
and U17144 (N_17144,N_15743,N_15240);
nor U17145 (N_17145,N_14595,N_14880);
or U17146 (N_17146,N_14684,N_15389);
nor U17147 (N_17147,N_14760,N_14023);
nor U17148 (N_17148,N_14972,N_14721);
or U17149 (N_17149,N_15869,N_14151);
nand U17150 (N_17150,N_15960,N_15767);
nand U17151 (N_17151,N_14479,N_15611);
nand U17152 (N_17152,N_14131,N_14837);
nor U17153 (N_17153,N_14929,N_14690);
nor U17154 (N_17154,N_14082,N_14911);
xnor U17155 (N_17155,N_15184,N_14447);
nor U17156 (N_17156,N_15750,N_15444);
nor U17157 (N_17157,N_15403,N_14732);
or U17158 (N_17158,N_15481,N_15041);
nor U17159 (N_17159,N_14016,N_14222);
xnor U17160 (N_17160,N_14373,N_15180);
nor U17161 (N_17161,N_15484,N_15636);
nor U17162 (N_17162,N_14785,N_15397);
or U17163 (N_17163,N_14867,N_14000);
or U17164 (N_17164,N_14468,N_15564);
nor U17165 (N_17165,N_14899,N_15069);
or U17166 (N_17166,N_14147,N_15634);
or U17167 (N_17167,N_15699,N_14469);
and U17168 (N_17168,N_15741,N_14313);
nand U17169 (N_17169,N_14107,N_15388);
and U17170 (N_17170,N_15563,N_14197);
nand U17171 (N_17171,N_15073,N_14512);
or U17172 (N_17172,N_14458,N_15091);
or U17173 (N_17173,N_15074,N_15473);
and U17174 (N_17174,N_15590,N_14593);
xor U17175 (N_17175,N_14546,N_14424);
nor U17176 (N_17176,N_14659,N_14144);
and U17177 (N_17177,N_14276,N_15884);
or U17178 (N_17178,N_15828,N_14367);
nand U17179 (N_17179,N_15167,N_14380);
nand U17180 (N_17180,N_15255,N_15920);
or U17181 (N_17181,N_15287,N_15750);
xnor U17182 (N_17182,N_14128,N_15905);
and U17183 (N_17183,N_14336,N_14406);
xor U17184 (N_17184,N_14902,N_15628);
xor U17185 (N_17185,N_14538,N_14492);
and U17186 (N_17186,N_14670,N_15977);
and U17187 (N_17187,N_14010,N_15317);
nand U17188 (N_17188,N_15323,N_15477);
and U17189 (N_17189,N_14832,N_15651);
xor U17190 (N_17190,N_15640,N_14860);
and U17191 (N_17191,N_15958,N_14333);
nand U17192 (N_17192,N_15058,N_15478);
nand U17193 (N_17193,N_14022,N_14802);
xor U17194 (N_17194,N_14370,N_14055);
and U17195 (N_17195,N_14225,N_14550);
nand U17196 (N_17196,N_14515,N_15987);
xor U17197 (N_17197,N_14707,N_15239);
and U17198 (N_17198,N_14835,N_14356);
or U17199 (N_17199,N_15164,N_15749);
and U17200 (N_17200,N_15481,N_14706);
nor U17201 (N_17201,N_14086,N_15892);
and U17202 (N_17202,N_14119,N_14087);
xnor U17203 (N_17203,N_14998,N_15357);
xnor U17204 (N_17204,N_15418,N_15843);
nor U17205 (N_17205,N_14481,N_14220);
and U17206 (N_17206,N_15704,N_14341);
nand U17207 (N_17207,N_15023,N_14730);
or U17208 (N_17208,N_15402,N_14191);
or U17209 (N_17209,N_15595,N_15652);
nor U17210 (N_17210,N_15086,N_15963);
or U17211 (N_17211,N_14490,N_15159);
or U17212 (N_17212,N_14387,N_14932);
xor U17213 (N_17213,N_14001,N_15140);
and U17214 (N_17214,N_14628,N_15647);
nand U17215 (N_17215,N_15158,N_15187);
xor U17216 (N_17216,N_14781,N_14580);
and U17217 (N_17217,N_15957,N_15954);
nor U17218 (N_17218,N_15501,N_14648);
nand U17219 (N_17219,N_15656,N_15170);
nor U17220 (N_17220,N_15589,N_14555);
nand U17221 (N_17221,N_14098,N_15963);
or U17222 (N_17222,N_15538,N_14994);
nand U17223 (N_17223,N_15455,N_15797);
or U17224 (N_17224,N_15728,N_15032);
nor U17225 (N_17225,N_14868,N_15561);
and U17226 (N_17226,N_14970,N_15347);
or U17227 (N_17227,N_15353,N_15617);
and U17228 (N_17228,N_14005,N_14418);
or U17229 (N_17229,N_14042,N_15619);
xor U17230 (N_17230,N_14501,N_15940);
nor U17231 (N_17231,N_14903,N_14962);
xor U17232 (N_17232,N_15738,N_15008);
and U17233 (N_17233,N_15996,N_14081);
or U17234 (N_17234,N_15853,N_15743);
or U17235 (N_17235,N_15148,N_15966);
nor U17236 (N_17236,N_14305,N_14913);
xor U17237 (N_17237,N_15824,N_15816);
or U17238 (N_17238,N_15787,N_14481);
xnor U17239 (N_17239,N_15767,N_14153);
or U17240 (N_17240,N_14289,N_14275);
xnor U17241 (N_17241,N_14624,N_15680);
and U17242 (N_17242,N_15231,N_14768);
nor U17243 (N_17243,N_14291,N_15944);
and U17244 (N_17244,N_14228,N_14765);
nand U17245 (N_17245,N_15160,N_15163);
nand U17246 (N_17246,N_14502,N_15036);
nor U17247 (N_17247,N_14860,N_15614);
nor U17248 (N_17248,N_14937,N_15141);
xor U17249 (N_17249,N_15978,N_15931);
or U17250 (N_17250,N_15661,N_15277);
and U17251 (N_17251,N_15866,N_14115);
xor U17252 (N_17252,N_14086,N_14640);
and U17253 (N_17253,N_15087,N_14636);
or U17254 (N_17254,N_14823,N_14104);
and U17255 (N_17255,N_14488,N_14177);
or U17256 (N_17256,N_15948,N_14676);
xor U17257 (N_17257,N_14217,N_15264);
nand U17258 (N_17258,N_15721,N_15490);
nand U17259 (N_17259,N_14760,N_14124);
nand U17260 (N_17260,N_14988,N_14009);
nand U17261 (N_17261,N_15571,N_14082);
or U17262 (N_17262,N_15756,N_15925);
nand U17263 (N_17263,N_14570,N_14248);
nor U17264 (N_17264,N_15044,N_15838);
nand U17265 (N_17265,N_14918,N_15890);
nor U17266 (N_17266,N_15851,N_14443);
xnor U17267 (N_17267,N_15915,N_15353);
nand U17268 (N_17268,N_15890,N_15446);
nor U17269 (N_17269,N_15664,N_14604);
xor U17270 (N_17270,N_15880,N_14932);
xnor U17271 (N_17271,N_14286,N_15133);
xnor U17272 (N_17272,N_15951,N_14136);
xor U17273 (N_17273,N_15835,N_14842);
xor U17274 (N_17274,N_14618,N_15685);
xor U17275 (N_17275,N_14828,N_14619);
nand U17276 (N_17276,N_15883,N_15616);
nor U17277 (N_17277,N_15947,N_14291);
or U17278 (N_17278,N_15715,N_15128);
xnor U17279 (N_17279,N_15812,N_15119);
nor U17280 (N_17280,N_14134,N_15240);
and U17281 (N_17281,N_15427,N_14361);
or U17282 (N_17282,N_14206,N_15987);
nand U17283 (N_17283,N_14157,N_15186);
nor U17284 (N_17284,N_14364,N_14656);
xor U17285 (N_17285,N_15237,N_14099);
and U17286 (N_17286,N_14844,N_15350);
or U17287 (N_17287,N_14156,N_15095);
or U17288 (N_17288,N_14908,N_15381);
or U17289 (N_17289,N_15970,N_14474);
nand U17290 (N_17290,N_14467,N_14527);
nand U17291 (N_17291,N_14859,N_14805);
nor U17292 (N_17292,N_15529,N_14207);
or U17293 (N_17293,N_14696,N_14582);
nand U17294 (N_17294,N_14583,N_14069);
nand U17295 (N_17295,N_15780,N_15074);
and U17296 (N_17296,N_14913,N_15560);
or U17297 (N_17297,N_14864,N_14726);
nor U17298 (N_17298,N_15579,N_15696);
nor U17299 (N_17299,N_14079,N_15596);
or U17300 (N_17300,N_15820,N_15603);
or U17301 (N_17301,N_15606,N_15485);
nor U17302 (N_17302,N_14551,N_15029);
nand U17303 (N_17303,N_14910,N_14152);
or U17304 (N_17304,N_15412,N_15364);
nor U17305 (N_17305,N_14076,N_15428);
nor U17306 (N_17306,N_15318,N_14842);
or U17307 (N_17307,N_14529,N_15132);
nand U17308 (N_17308,N_14207,N_14461);
or U17309 (N_17309,N_14954,N_14630);
xor U17310 (N_17310,N_14194,N_14162);
xnor U17311 (N_17311,N_14832,N_15134);
xor U17312 (N_17312,N_15493,N_14185);
xnor U17313 (N_17313,N_14367,N_15065);
nor U17314 (N_17314,N_15089,N_14014);
and U17315 (N_17315,N_14287,N_15820);
nor U17316 (N_17316,N_14963,N_15089);
nand U17317 (N_17317,N_15834,N_14520);
nand U17318 (N_17318,N_14329,N_14234);
or U17319 (N_17319,N_14839,N_15540);
nand U17320 (N_17320,N_15820,N_15186);
nand U17321 (N_17321,N_14115,N_15360);
nor U17322 (N_17322,N_14571,N_14897);
nor U17323 (N_17323,N_14179,N_14981);
nor U17324 (N_17324,N_14789,N_14133);
nor U17325 (N_17325,N_15257,N_15226);
nor U17326 (N_17326,N_14455,N_15267);
xor U17327 (N_17327,N_15620,N_15550);
nand U17328 (N_17328,N_14155,N_15563);
nand U17329 (N_17329,N_14469,N_14587);
nor U17330 (N_17330,N_15241,N_15440);
or U17331 (N_17331,N_15693,N_14416);
nor U17332 (N_17332,N_14269,N_14783);
xnor U17333 (N_17333,N_14738,N_15490);
nand U17334 (N_17334,N_15327,N_15181);
and U17335 (N_17335,N_14895,N_15047);
nor U17336 (N_17336,N_14821,N_15264);
nand U17337 (N_17337,N_14172,N_15698);
or U17338 (N_17338,N_14359,N_14783);
or U17339 (N_17339,N_15707,N_14612);
or U17340 (N_17340,N_15189,N_15975);
nor U17341 (N_17341,N_15071,N_15653);
xor U17342 (N_17342,N_14378,N_15811);
xor U17343 (N_17343,N_14859,N_15524);
nand U17344 (N_17344,N_15806,N_14494);
xnor U17345 (N_17345,N_14450,N_15290);
or U17346 (N_17346,N_14822,N_14657);
or U17347 (N_17347,N_14976,N_14041);
xnor U17348 (N_17348,N_14038,N_14828);
or U17349 (N_17349,N_14470,N_14639);
nor U17350 (N_17350,N_15568,N_15263);
nand U17351 (N_17351,N_15212,N_15914);
nor U17352 (N_17352,N_14755,N_14485);
nor U17353 (N_17353,N_14609,N_15025);
xor U17354 (N_17354,N_14000,N_15687);
and U17355 (N_17355,N_15495,N_14620);
xor U17356 (N_17356,N_14173,N_15960);
nand U17357 (N_17357,N_14122,N_14403);
and U17358 (N_17358,N_14724,N_14397);
nor U17359 (N_17359,N_14885,N_14507);
xnor U17360 (N_17360,N_14721,N_15104);
xor U17361 (N_17361,N_15356,N_15037);
xnor U17362 (N_17362,N_14186,N_14880);
xor U17363 (N_17363,N_15239,N_15691);
nand U17364 (N_17364,N_14618,N_15345);
or U17365 (N_17365,N_14837,N_14868);
nor U17366 (N_17366,N_14373,N_14039);
nor U17367 (N_17367,N_14040,N_14265);
nor U17368 (N_17368,N_15899,N_14455);
nor U17369 (N_17369,N_14297,N_15403);
or U17370 (N_17370,N_15264,N_15921);
and U17371 (N_17371,N_14697,N_14465);
xnor U17372 (N_17372,N_14953,N_14010);
and U17373 (N_17373,N_14843,N_14771);
nand U17374 (N_17374,N_15668,N_14110);
nor U17375 (N_17375,N_15836,N_15187);
xnor U17376 (N_17376,N_15886,N_15483);
xnor U17377 (N_17377,N_15433,N_15130);
and U17378 (N_17378,N_15198,N_15448);
or U17379 (N_17379,N_14880,N_15118);
xnor U17380 (N_17380,N_14884,N_15132);
nor U17381 (N_17381,N_15443,N_15478);
nand U17382 (N_17382,N_14616,N_14963);
and U17383 (N_17383,N_15150,N_15863);
xor U17384 (N_17384,N_15646,N_15766);
nor U17385 (N_17385,N_14206,N_15502);
nand U17386 (N_17386,N_14394,N_15169);
nand U17387 (N_17387,N_15799,N_15471);
and U17388 (N_17388,N_15418,N_14926);
xnor U17389 (N_17389,N_15759,N_15507);
nor U17390 (N_17390,N_14766,N_14953);
xnor U17391 (N_17391,N_14258,N_15772);
xor U17392 (N_17392,N_14054,N_14018);
nand U17393 (N_17393,N_15271,N_15434);
and U17394 (N_17394,N_15969,N_15036);
xnor U17395 (N_17395,N_15231,N_14003);
nand U17396 (N_17396,N_15771,N_15258);
nor U17397 (N_17397,N_14614,N_15341);
or U17398 (N_17398,N_15301,N_15169);
nor U17399 (N_17399,N_15920,N_15589);
and U17400 (N_17400,N_15929,N_14764);
nand U17401 (N_17401,N_14236,N_15753);
nand U17402 (N_17402,N_15037,N_14041);
or U17403 (N_17403,N_15115,N_15081);
nand U17404 (N_17404,N_15255,N_14098);
nor U17405 (N_17405,N_15384,N_15502);
or U17406 (N_17406,N_15537,N_14095);
nor U17407 (N_17407,N_14815,N_14619);
xor U17408 (N_17408,N_15768,N_15851);
nor U17409 (N_17409,N_15287,N_15542);
nand U17410 (N_17410,N_14408,N_14246);
nand U17411 (N_17411,N_14909,N_15531);
nor U17412 (N_17412,N_14223,N_15221);
or U17413 (N_17413,N_14561,N_14527);
xnor U17414 (N_17414,N_14082,N_14034);
and U17415 (N_17415,N_14063,N_14105);
nor U17416 (N_17416,N_14896,N_15094);
and U17417 (N_17417,N_14175,N_14546);
xnor U17418 (N_17418,N_14320,N_14295);
nand U17419 (N_17419,N_14085,N_14303);
and U17420 (N_17420,N_14426,N_15706);
nand U17421 (N_17421,N_15095,N_15278);
xor U17422 (N_17422,N_15893,N_14317);
or U17423 (N_17423,N_15865,N_14400);
xor U17424 (N_17424,N_15443,N_15305);
and U17425 (N_17425,N_14259,N_15356);
xnor U17426 (N_17426,N_14780,N_14015);
nand U17427 (N_17427,N_15627,N_14545);
xor U17428 (N_17428,N_15680,N_14257);
nor U17429 (N_17429,N_14299,N_15261);
and U17430 (N_17430,N_14527,N_15414);
nor U17431 (N_17431,N_14956,N_15126);
or U17432 (N_17432,N_15099,N_15159);
and U17433 (N_17433,N_15269,N_14180);
nand U17434 (N_17434,N_15776,N_15257);
or U17435 (N_17435,N_15147,N_14943);
nor U17436 (N_17436,N_14288,N_15095);
xnor U17437 (N_17437,N_14971,N_15003);
and U17438 (N_17438,N_14282,N_14254);
nand U17439 (N_17439,N_14203,N_14364);
nand U17440 (N_17440,N_15898,N_14110);
nand U17441 (N_17441,N_14454,N_15167);
and U17442 (N_17442,N_15603,N_14136);
or U17443 (N_17443,N_15656,N_15857);
xor U17444 (N_17444,N_14433,N_15858);
and U17445 (N_17445,N_14011,N_14090);
nor U17446 (N_17446,N_14562,N_14615);
nor U17447 (N_17447,N_14557,N_14781);
xor U17448 (N_17448,N_15258,N_14608);
xor U17449 (N_17449,N_15355,N_15116);
nor U17450 (N_17450,N_15009,N_14193);
or U17451 (N_17451,N_14584,N_14755);
and U17452 (N_17452,N_14742,N_15312);
nor U17453 (N_17453,N_14726,N_15288);
or U17454 (N_17454,N_15472,N_15804);
and U17455 (N_17455,N_15095,N_15339);
and U17456 (N_17456,N_14692,N_15758);
nand U17457 (N_17457,N_14167,N_14583);
xnor U17458 (N_17458,N_15443,N_14588);
or U17459 (N_17459,N_15791,N_15546);
xnor U17460 (N_17460,N_14697,N_15216);
nor U17461 (N_17461,N_14539,N_15741);
xnor U17462 (N_17462,N_14282,N_15915);
or U17463 (N_17463,N_15157,N_15947);
or U17464 (N_17464,N_15728,N_14103);
or U17465 (N_17465,N_15851,N_15820);
or U17466 (N_17466,N_14307,N_14874);
nor U17467 (N_17467,N_15189,N_15659);
xor U17468 (N_17468,N_14446,N_14127);
xnor U17469 (N_17469,N_14578,N_14589);
nand U17470 (N_17470,N_14136,N_14946);
nand U17471 (N_17471,N_15132,N_14249);
or U17472 (N_17472,N_14438,N_14794);
nand U17473 (N_17473,N_14482,N_15781);
nor U17474 (N_17474,N_15392,N_15118);
xor U17475 (N_17475,N_15956,N_15571);
and U17476 (N_17476,N_14681,N_14139);
xor U17477 (N_17477,N_15113,N_14172);
or U17478 (N_17478,N_15957,N_15968);
xor U17479 (N_17479,N_14533,N_15422);
or U17480 (N_17480,N_14916,N_15422);
or U17481 (N_17481,N_15795,N_15468);
or U17482 (N_17482,N_15099,N_15557);
and U17483 (N_17483,N_15039,N_15643);
nand U17484 (N_17484,N_15389,N_15088);
nand U17485 (N_17485,N_14238,N_14668);
nor U17486 (N_17486,N_15345,N_14940);
and U17487 (N_17487,N_15510,N_15404);
or U17488 (N_17488,N_15591,N_14162);
xor U17489 (N_17489,N_14863,N_15690);
nor U17490 (N_17490,N_15815,N_15910);
xnor U17491 (N_17491,N_14098,N_15102);
or U17492 (N_17492,N_14223,N_15665);
or U17493 (N_17493,N_14722,N_15947);
and U17494 (N_17494,N_15183,N_15637);
nand U17495 (N_17495,N_14105,N_15327);
nor U17496 (N_17496,N_14530,N_14817);
nand U17497 (N_17497,N_15259,N_14410);
nand U17498 (N_17498,N_15434,N_14682);
xnor U17499 (N_17499,N_15705,N_15529);
or U17500 (N_17500,N_14495,N_14667);
and U17501 (N_17501,N_15537,N_14874);
and U17502 (N_17502,N_15668,N_15942);
nor U17503 (N_17503,N_15380,N_14593);
nor U17504 (N_17504,N_15883,N_15913);
xnor U17505 (N_17505,N_14793,N_15183);
nand U17506 (N_17506,N_15980,N_14714);
nand U17507 (N_17507,N_15381,N_15730);
xnor U17508 (N_17508,N_15195,N_15959);
or U17509 (N_17509,N_15211,N_15893);
xnor U17510 (N_17510,N_15474,N_15140);
or U17511 (N_17511,N_14992,N_14951);
and U17512 (N_17512,N_14685,N_15462);
xnor U17513 (N_17513,N_14557,N_15569);
and U17514 (N_17514,N_14196,N_15635);
and U17515 (N_17515,N_14232,N_15353);
xor U17516 (N_17516,N_15364,N_15999);
and U17517 (N_17517,N_14679,N_15169);
nand U17518 (N_17518,N_15274,N_14734);
or U17519 (N_17519,N_15715,N_15603);
nor U17520 (N_17520,N_15880,N_15917);
nand U17521 (N_17521,N_14776,N_14471);
xor U17522 (N_17522,N_14495,N_15175);
nor U17523 (N_17523,N_15180,N_14015);
or U17524 (N_17524,N_15094,N_14132);
or U17525 (N_17525,N_15658,N_14746);
and U17526 (N_17526,N_15136,N_14226);
or U17527 (N_17527,N_14793,N_15031);
xor U17528 (N_17528,N_14253,N_14130);
or U17529 (N_17529,N_14260,N_15098);
nand U17530 (N_17530,N_15312,N_14597);
and U17531 (N_17531,N_14637,N_15060);
and U17532 (N_17532,N_14891,N_15630);
nor U17533 (N_17533,N_15460,N_15681);
and U17534 (N_17534,N_14014,N_15509);
or U17535 (N_17535,N_14002,N_15551);
xor U17536 (N_17536,N_14759,N_15742);
and U17537 (N_17537,N_15042,N_15272);
nand U17538 (N_17538,N_14070,N_15647);
xnor U17539 (N_17539,N_15102,N_14073);
or U17540 (N_17540,N_14923,N_15483);
nor U17541 (N_17541,N_15926,N_15772);
or U17542 (N_17542,N_15482,N_15641);
nand U17543 (N_17543,N_14196,N_15339);
and U17544 (N_17544,N_14039,N_14253);
xor U17545 (N_17545,N_15921,N_15170);
nor U17546 (N_17546,N_14983,N_15669);
nor U17547 (N_17547,N_14166,N_14460);
xnor U17548 (N_17548,N_14867,N_14769);
nor U17549 (N_17549,N_15548,N_15513);
nor U17550 (N_17550,N_15079,N_15226);
nand U17551 (N_17551,N_15406,N_14218);
nand U17552 (N_17552,N_14513,N_15655);
and U17553 (N_17553,N_14738,N_14891);
or U17554 (N_17554,N_14971,N_15030);
or U17555 (N_17555,N_15660,N_14923);
and U17556 (N_17556,N_15401,N_15000);
nand U17557 (N_17557,N_15129,N_14226);
or U17558 (N_17558,N_15452,N_15041);
or U17559 (N_17559,N_14469,N_14161);
nand U17560 (N_17560,N_14036,N_15277);
or U17561 (N_17561,N_14453,N_15230);
or U17562 (N_17562,N_15242,N_15412);
and U17563 (N_17563,N_14888,N_14475);
nand U17564 (N_17564,N_15515,N_15161);
xnor U17565 (N_17565,N_15662,N_15177);
nand U17566 (N_17566,N_15560,N_14163);
nand U17567 (N_17567,N_14489,N_14691);
xor U17568 (N_17568,N_15338,N_15607);
nand U17569 (N_17569,N_14567,N_14696);
nor U17570 (N_17570,N_15261,N_14995);
nand U17571 (N_17571,N_14366,N_14386);
or U17572 (N_17572,N_14878,N_15046);
and U17573 (N_17573,N_14214,N_14958);
or U17574 (N_17574,N_14689,N_14968);
xor U17575 (N_17575,N_14615,N_14097);
nor U17576 (N_17576,N_14862,N_15140);
and U17577 (N_17577,N_15867,N_15953);
nor U17578 (N_17578,N_14619,N_14212);
nand U17579 (N_17579,N_15405,N_14512);
or U17580 (N_17580,N_15320,N_14328);
nand U17581 (N_17581,N_14626,N_14843);
or U17582 (N_17582,N_15116,N_14953);
nand U17583 (N_17583,N_14071,N_15728);
or U17584 (N_17584,N_14449,N_14363);
and U17585 (N_17585,N_15068,N_15703);
nand U17586 (N_17586,N_15487,N_15096);
or U17587 (N_17587,N_14840,N_14762);
and U17588 (N_17588,N_15607,N_14635);
xnor U17589 (N_17589,N_15520,N_14836);
and U17590 (N_17590,N_15004,N_15526);
and U17591 (N_17591,N_14589,N_15989);
and U17592 (N_17592,N_14767,N_14020);
nand U17593 (N_17593,N_14318,N_15193);
xnor U17594 (N_17594,N_14990,N_14184);
or U17595 (N_17595,N_15248,N_14405);
or U17596 (N_17596,N_14336,N_15266);
nand U17597 (N_17597,N_14656,N_15209);
xnor U17598 (N_17598,N_14728,N_14291);
xnor U17599 (N_17599,N_14889,N_15031);
and U17600 (N_17600,N_15906,N_14584);
or U17601 (N_17601,N_14948,N_14463);
xnor U17602 (N_17602,N_15850,N_14067);
and U17603 (N_17603,N_15790,N_15723);
nand U17604 (N_17604,N_15913,N_15233);
nand U17605 (N_17605,N_15541,N_14522);
xnor U17606 (N_17606,N_15109,N_14320);
and U17607 (N_17607,N_15416,N_14869);
xnor U17608 (N_17608,N_15202,N_14080);
and U17609 (N_17609,N_15644,N_15276);
nor U17610 (N_17610,N_15073,N_15722);
and U17611 (N_17611,N_14862,N_15246);
and U17612 (N_17612,N_14333,N_14799);
or U17613 (N_17613,N_15010,N_15793);
nor U17614 (N_17614,N_14507,N_14486);
or U17615 (N_17615,N_15907,N_14457);
and U17616 (N_17616,N_14575,N_15021);
nor U17617 (N_17617,N_14265,N_14443);
nand U17618 (N_17618,N_15236,N_14662);
or U17619 (N_17619,N_14723,N_14389);
or U17620 (N_17620,N_15291,N_15706);
nand U17621 (N_17621,N_15558,N_14260);
and U17622 (N_17622,N_15658,N_14325);
or U17623 (N_17623,N_15455,N_15126);
or U17624 (N_17624,N_15287,N_15746);
or U17625 (N_17625,N_15085,N_15906);
nor U17626 (N_17626,N_14041,N_15310);
xor U17627 (N_17627,N_14058,N_14457);
and U17628 (N_17628,N_14779,N_15860);
and U17629 (N_17629,N_15766,N_15275);
and U17630 (N_17630,N_14681,N_14263);
nand U17631 (N_17631,N_15061,N_15847);
or U17632 (N_17632,N_15845,N_14645);
xor U17633 (N_17633,N_15870,N_14307);
or U17634 (N_17634,N_15853,N_15190);
and U17635 (N_17635,N_15784,N_14878);
xnor U17636 (N_17636,N_15009,N_14447);
and U17637 (N_17637,N_15938,N_15446);
and U17638 (N_17638,N_15725,N_15338);
xnor U17639 (N_17639,N_14995,N_15391);
xnor U17640 (N_17640,N_15844,N_14421);
and U17641 (N_17641,N_15815,N_15432);
nand U17642 (N_17642,N_15898,N_14154);
nand U17643 (N_17643,N_14495,N_15289);
xor U17644 (N_17644,N_14546,N_14817);
and U17645 (N_17645,N_14380,N_15970);
and U17646 (N_17646,N_14963,N_15562);
xnor U17647 (N_17647,N_14989,N_15676);
xor U17648 (N_17648,N_15634,N_15403);
xor U17649 (N_17649,N_14670,N_14324);
nand U17650 (N_17650,N_15527,N_15006);
nand U17651 (N_17651,N_14875,N_14794);
nor U17652 (N_17652,N_15409,N_14351);
nand U17653 (N_17653,N_14930,N_14407);
nor U17654 (N_17654,N_14900,N_15178);
nor U17655 (N_17655,N_14689,N_14247);
and U17656 (N_17656,N_14368,N_15947);
nand U17657 (N_17657,N_14292,N_15127);
and U17658 (N_17658,N_14880,N_14962);
nand U17659 (N_17659,N_14789,N_14815);
and U17660 (N_17660,N_14489,N_15959);
nor U17661 (N_17661,N_14563,N_14914);
or U17662 (N_17662,N_15696,N_15828);
nor U17663 (N_17663,N_15578,N_14600);
xnor U17664 (N_17664,N_15025,N_15601);
nand U17665 (N_17665,N_15303,N_14160);
or U17666 (N_17666,N_14283,N_14960);
nand U17667 (N_17667,N_15868,N_14302);
nor U17668 (N_17668,N_14075,N_15956);
nor U17669 (N_17669,N_14461,N_14687);
xnor U17670 (N_17670,N_14593,N_14196);
nand U17671 (N_17671,N_15356,N_14311);
nand U17672 (N_17672,N_15588,N_15638);
nor U17673 (N_17673,N_15047,N_14426);
nor U17674 (N_17674,N_15181,N_14743);
nand U17675 (N_17675,N_15429,N_14715);
nand U17676 (N_17676,N_15463,N_15720);
nand U17677 (N_17677,N_14177,N_15770);
nand U17678 (N_17678,N_14241,N_14935);
nor U17679 (N_17679,N_14398,N_14588);
and U17680 (N_17680,N_14764,N_14387);
or U17681 (N_17681,N_15899,N_14693);
nor U17682 (N_17682,N_14437,N_14684);
nand U17683 (N_17683,N_14399,N_15465);
nand U17684 (N_17684,N_14939,N_15473);
and U17685 (N_17685,N_15264,N_14543);
nor U17686 (N_17686,N_14948,N_15659);
nand U17687 (N_17687,N_15259,N_14879);
and U17688 (N_17688,N_14038,N_15097);
and U17689 (N_17689,N_15656,N_14539);
xor U17690 (N_17690,N_14629,N_15204);
xnor U17691 (N_17691,N_15001,N_15195);
nor U17692 (N_17692,N_14978,N_15002);
or U17693 (N_17693,N_15859,N_15998);
nand U17694 (N_17694,N_15169,N_15913);
and U17695 (N_17695,N_14166,N_14900);
and U17696 (N_17696,N_15413,N_15820);
and U17697 (N_17697,N_15145,N_14125);
or U17698 (N_17698,N_15352,N_15033);
or U17699 (N_17699,N_14462,N_14601);
nand U17700 (N_17700,N_14989,N_15288);
nand U17701 (N_17701,N_14170,N_15830);
nor U17702 (N_17702,N_15196,N_14005);
nand U17703 (N_17703,N_14095,N_15480);
nand U17704 (N_17704,N_14307,N_15086);
and U17705 (N_17705,N_14224,N_14289);
xnor U17706 (N_17706,N_14670,N_14509);
nand U17707 (N_17707,N_15847,N_14060);
and U17708 (N_17708,N_14363,N_15153);
nand U17709 (N_17709,N_15578,N_14532);
nand U17710 (N_17710,N_14570,N_15513);
xnor U17711 (N_17711,N_15904,N_15617);
and U17712 (N_17712,N_14817,N_15540);
nand U17713 (N_17713,N_14572,N_15446);
xnor U17714 (N_17714,N_14938,N_14450);
nand U17715 (N_17715,N_15916,N_14428);
or U17716 (N_17716,N_15533,N_15983);
xnor U17717 (N_17717,N_14470,N_15967);
nand U17718 (N_17718,N_14811,N_14898);
and U17719 (N_17719,N_15457,N_14779);
and U17720 (N_17720,N_14214,N_14026);
nor U17721 (N_17721,N_15484,N_14728);
and U17722 (N_17722,N_14138,N_14681);
nand U17723 (N_17723,N_14461,N_14808);
xnor U17724 (N_17724,N_15937,N_14504);
nand U17725 (N_17725,N_15424,N_15560);
or U17726 (N_17726,N_15006,N_15923);
and U17727 (N_17727,N_15367,N_14822);
nor U17728 (N_17728,N_14428,N_15238);
xor U17729 (N_17729,N_15204,N_14753);
nand U17730 (N_17730,N_14959,N_14666);
nand U17731 (N_17731,N_14305,N_14512);
nand U17732 (N_17732,N_14674,N_14672);
xor U17733 (N_17733,N_15662,N_14626);
xor U17734 (N_17734,N_14524,N_15403);
and U17735 (N_17735,N_15084,N_14900);
or U17736 (N_17736,N_15973,N_14513);
nor U17737 (N_17737,N_15270,N_14339);
nor U17738 (N_17738,N_14226,N_14748);
xnor U17739 (N_17739,N_15156,N_14065);
or U17740 (N_17740,N_15562,N_15176);
nor U17741 (N_17741,N_14415,N_15422);
nor U17742 (N_17742,N_15553,N_14618);
and U17743 (N_17743,N_14375,N_15431);
nand U17744 (N_17744,N_15316,N_14784);
and U17745 (N_17745,N_14700,N_15911);
or U17746 (N_17746,N_14820,N_15498);
and U17747 (N_17747,N_14497,N_15374);
nor U17748 (N_17748,N_14276,N_15530);
xor U17749 (N_17749,N_14322,N_14979);
and U17750 (N_17750,N_14953,N_14161);
xor U17751 (N_17751,N_15318,N_14190);
nor U17752 (N_17752,N_15089,N_15697);
and U17753 (N_17753,N_14524,N_14782);
and U17754 (N_17754,N_14308,N_14957);
nand U17755 (N_17755,N_15453,N_14750);
xnor U17756 (N_17756,N_14877,N_14254);
nor U17757 (N_17757,N_14331,N_14539);
xor U17758 (N_17758,N_14665,N_14413);
or U17759 (N_17759,N_15824,N_15384);
nand U17760 (N_17760,N_14169,N_14408);
or U17761 (N_17761,N_14235,N_14870);
xor U17762 (N_17762,N_15469,N_14425);
xor U17763 (N_17763,N_14226,N_14293);
nor U17764 (N_17764,N_14235,N_15587);
xnor U17765 (N_17765,N_15534,N_14014);
nand U17766 (N_17766,N_14750,N_15214);
nor U17767 (N_17767,N_15616,N_15350);
xor U17768 (N_17768,N_15974,N_14282);
nand U17769 (N_17769,N_14484,N_15120);
and U17770 (N_17770,N_14310,N_15638);
nor U17771 (N_17771,N_14772,N_14749);
xnor U17772 (N_17772,N_14741,N_15157);
and U17773 (N_17773,N_14099,N_15911);
or U17774 (N_17774,N_15620,N_15877);
nor U17775 (N_17775,N_14104,N_14946);
and U17776 (N_17776,N_14755,N_15462);
xor U17777 (N_17777,N_15771,N_15352);
or U17778 (N_17778,N_14179,N_14369);
and U17779 (N_17779,N_15272,N_15783);
nor U17780 (N_17780,N_14217,N_15802);
and U17781 (N_17781,N_15342,N_14871);
or U17782 (N_17782,N_15571,N_14518);
or U17783 (N_17783,N_15428,N_14976);
or U17784 (N_17784,N_14622,N_15013);
xnor U17785 (N_17785,N_15729,N_14973);
or U17786 (N_17786,N_14505,N_15672);
xor U17787 (N_17787,N_15682,N_15076);
nor U17788 (N_17788,N_15076,N_14308);
or U17789 (N_17789,N_14384,N_14489);
xor U17790 (N_17790,N_15602,N_14977);
nand U17791 (N_17791,N_14418,N_15163);
nor U17792 (N_17792,N_15478,N_14195);
xor U17793 (N_17793,N_15154,N_15911);
and U17794 (N_17794,N_15753,N_14595);
or U17795 (N_17795,N_14830,N_15803);
nand U17796 (N_17796,N_15965,N_14858);
xor U17797 (N_17797,N_14726,N_14928);
and U17798 (N_17798,N_15088,N_15365);
and U17799 (N_17799,N_15402,N_14427);
or U17800 (N_17800,N_14448,N_15177);
nand U17801 (N_17801,N_14920,N_15202);
nand U17802 (N_17802,N_15075,N_15662);
nor U17803 (N_17803,N_14646,N_15337);
nor U17804 (N_17804,N_14175,N_14083);
xnor U17805 (N_17805,N_14511,N_15083);
nor U17806 (N_17806,N_15530,N_15370);
xnor U17807 (N_17807,N_15350,N_15745);
nor U17808 (N_17808,N_15019,N_14923);
xnor U17809 (N_17809,N_15567,N_14021);
nor U17810 (N_17810,N_14579,N_14225);
or U17811 (N_17811,N_15117,N_15735);
xnor U17812 (N_17812,N_14309,N_14433);
nor U17813 (N_17813,N_14674,N_15056);
nor U17814 (N_17814,N_15160,N_14474);
and U17815 (N_17815,N_14864,N_15989);
nor U17816 (N_17816,N_14039,N_15093);
xnor U17817 (N_17817,N_14132,N_14151);
xor U17818 (N_17818,N_15380,N_15829);
or U17819 (N_17819,N_14698,N_15465);
nor U17820 (N_17820,N_14753,N_14882);
xnor U17821 (N_17821,N_14679,N_15339);
nor U17822 (N_17822,N_15496,N_15394);
nor U17823 (N_17823,N_14996,N_14938);
and U17824 (N_17824,N_14616,N_14804);
and U17825 (N_17825,N_15116,N_15356);
xnor U17826 (N_17826,N_14760,N_15298);
or U17827 (N_17827,N_14801,N_15302);
xnor U17828 (N_17828,N_15197,N_15989);
xor U17829 (N_17829,N_15117,N_15045);
or U17830 (N_17830,N_14693,N_14643);
xnor U17831 (N_17831,N_15169,N_14918);
and U17832 (N_17832,N_15617,N_15270);
nand U17833 (N_17833,N_14344,N_15666);
nor U17834 (N_17834,N_15425,N_15104);
nor U17835 (N_17835,N_15560,N_14342);
nor U17836 (N_17836,N_14627,N_14994);
xnor U17837 (N_17837,N_14420,N_14291);
nand U17838 (N_17838,N_15647,N_14414);
or U17839 (N_17839,N_14894,N_15714);
nand U17840 (N_17840,N_14064,N_15334);
nand U17841 (N_17841,N_14692,N_14499);
and U17842 (N_17842,N_15002,N_15513);
and U17843 (N_17843,N_14736,N_15249);
nor U17844 (N_17844,N_14839,N_15268);
nor U17845 (N_17845,N_14496,N_15378);
and U17846 (N_17846,N_14786,N_14215);
nand U17847 (N_17847,N_15260,N_15833);
nand U17848 (N_17848,N_14287,N_14431);
or U17849 (N_17849,N_15878,N_14631);
nor U17850 (N_17850,N_14372,N_14611);
nand U17851 (N_17851,N_14295,N_14228);
or U17852 (N_17852,N_15977,N_14078);
and U17853 (N_17853,N_14500,N_15816);
and U17854 (N_17854,N_14978,N_15790);
and U17855 (N_17855,N_15808,N_15921);
nor U17856 (N_17856,N_15224,N_14247);
and U17857 (N_17857,N_15149,N_14411);
xnor U17858 (N_17858,N_14682,N_14482);
nand U17859 (N_17859,N_14809,N_14400);
xnor U17860 (N_17860,N_14472,N_15234);
nand U17861 (N_17861,N_14808,N_15521);
and U17862 (N_17862,N_14773,N_14504);
and U17863 (N_17863,N_14172,N_14502);
and U17864 (N_17864,N_15833,N_15479);
and U17865 (N_17865,N_15310,N_14092);
nand U17866 (N_17866,N_14452,N_15601);
or U17867 (N_17867,N_14824,N_14435);
nand U17868 (N_17868,N_14511,N_15530);
nand U17869 (N_17869,N_15864,N_15417);
xor U17870 (N_17870,N_15432,N_15813);
and U17871 (N_17871,N_14341,N_14386);
and U17872 (N_17872,N_14026,N_15385);
xor U17873 (N_17873,N_15637,N_14251);
or U17874 (N_17874,N_14778,N_15784);
and U17875 (N_17875,N_14174,N_15313);
and U17876 (N_17876,N_14507,N_15112);
and U17877 (N_17877,N_14566,N_15117);
or U17878 (N_17878,N_15958,N_15263);
or U17879 (N_17879,N_14414,N_14939);
and U17880 (N_17880,N_14190,N_14552);
nand U17881 (N_17881,N_14667,N_15358);
nand U17882 (N_17882,N_15231,N_15909);
nor U17883 (N_17883,N_15104,N_14414);
nor U17884 (N_17884,N_15989,N_15201);
nand U17885 (N_17885,N_14793,N_14688);
or U17886 (N_17886,N_14740,N_14213);
nand U17887 (N_17887,N_14066,N_15869);
or U17888 (N_17888,N_15178,N_14811);
nand U17889 (N_17889,N_14156,N_15860);
or U17890 (N_17890,N_14911,N_14422);
nor U17891 (N_17891,N_14915,N_14864);
nand U17892 (N_17892,N_14019,N_14684);
and U17893 (N_17893,N_15059,N_14270);
or U17894 (N_17894,N_15515,N_15891);
or U17895 (N_17895,N_15306,N_14047);
nand U17896 (N_17896,N_15649,N_14970);
nor U17897 (N_17897,N_14148,N_14715);
nor U17898 (N_17898,N_15935,N_15488);
xor U17899 (N_17899,N_15600,N_14944);
and U17900 (N_17900,N_15573,N_14902);
nor U17901 (N_17901,N_14212,N_14218);
xnor U17902 (N_17902,N_15354,N_14555);
and U17903 (N_17903,N_14385,N_14432);
nand U17904 (N_17904,N_15497,N_14831);
or U17905 (N_17905,N_15027,N_14899);
xnor U17906 (N_17906,N_14527,N_14125);
nand U17907 (N_17907,N_14099,N_15976);
and U17908 (N_17908,N_15829,N_15242);
or U17909 (N_17909,N_15084,N_14904);
nand U17910 (N_17910,N_14693,N_14753);
or U17911 (N_17911,N_14879,N_14895);
nand U17912 (N_17912,N_14033,N_15559);
nor U17913 (N_17913,N_15677,N_15098);
and U17914 (N_17914,N_15467,N_15232);
xor U17915 (N_17915,N_15149,N_14902);
nand U17916 (N_17916,N_15492,N_14775);
or U17917 (N_17917,N_15759,N_14598);
nor U17918 (N_17918,N_14523,N_15797);
or U17919 (N_17919,N_15246,N_15629);
nand U17920 (N_17920,N_14525,N_15459);
or U17921 (N_17921,N_14894,N_14082);
xnor U17922 (N_17922,N_15908,N_15974);
nor U17923 (N_17923,N_15564,N_15968);
nor U17924 (N_17924,N_14901,N_15792);
xnor U17925 (N_17925,N_14470,N_14144);
nor U17926 (N_17926,N_14503,N_15675);
or U17927 (N_17927,N_15416,N_15058);
nand U17928 (N_17928,N_14786,N_14225);
or U17929 (N_17929,N_14743,N_15121);
nor U17930 (N_17930,N_15918,N_14815);
or U17931 (N_17931,N_14577,N_15371);
xnor U17932 (N_17932,N_15987,N_15762);
xor U17933 (N_17933,N_14167,N_14335);
and U17934 (N_17934,N_14889,N_14329);
nor U17935 (N_17935,N_14220,N_15039);
nor U17936 (N_17936,N_15392,N_15611);
or U17937 (N_17937,N_15261,N_15958);
and U17938 (N_17938,N_14002,N_14283);
and U17939 (N_17939,N_14479,N_14051);
xnor U17940 (N_17940,N_14337,N_14689);
xor U17941 (N_17941,N_15661,N_15280);
or U17942 (N_17942,N_15006,N_14674);
nor U17943 (N_17943,N_15795,N_14741);
or U17944 (N_17944,N_15167,N_14902);
xnor U17945 (N_17945,N_15525,N_14467);
nor U17946 (N_17946,N_14858,N_15028);
nand U17947 (N_17947,N_15283,N_14719);
or U17948 (N_17948,N_14154,N_14510);
and U17949 (N_17949,N_14900,N_14610);
nor U17950 (N_17950,N_15783,N_14325);
and U17951 (N_17951,N_15884,N_15330);
nor U17952 (N_17952,N_14582,N_14536);
xnor U17953 (N_17953,N_15570,N_14020);
nor U17954 (N_17954,N_15158,N_14424);
xor U17955 (N_17955,N_15786,N_14134);
nor U17956 (N_17956,N_14674,N_14737);
nor U17957 (N_17957,N_14391,N_15720);
xor U17958 (N_17958,N_15692,N_14184);
nor U17959 (N_17959,N_15548,N_15499);
nand U17960 (N_17960,N_15750,N_15689);
and U17961 (N_17961,N_14794,N_14537);
xnor U17962 (N_17962,N_15698,N_14533);
nand U17963 (N_17963,N_15746,N_15473);
xnor U17964 (N_17964,N_15449,N_15749);
nor U17965 (N_17965,N_14206,N_14917);
nor U17966 (N_17966,N_15089,N_14655);
nand U17967 (N_17967,N_15395,N_15712);
nor U17968 (N_17968,N_14405,N_15062);
xor U17969 (N_17969,N_15551,N_14671);
and U17970 (N_17970,N_14767,N_14670);
or U17971 (N_17971,N_15736,N_15242);
or U17972 (N_17972,N_14487,N_15752);
nor U17973 (N_17973,N_15257,N_15187);
and U17974 (N_17974,N_14168,N_14801);
nor U17975 (N_17975,N_15439,N_14009);
and U17976 (N_17976,N_15124,N_15133);
xnor U17977 (N_17977,N_15922,N_15621);
nor U17978 (N_17978,N_15942,N_14575);
xnor U17979 (N_17979,N_15626,N_14383);
nor U17980 (N_17980,N_15111,N_14798);
and U17981 (N_17981,N_14238,N_14991);
or U17982 (N_17982,N_14173,N_14411);
xor U17983 (N_17983,N_14850,N_15638);
or U17984 (N_17984,N_15905,N_15792);
nand U17985 (N_17985,N_14000,N_15717);
and U17986 (N_17986,N_14340,N_14977);
xor U17987 (N_17987,N_15319,N_14616);
nand U17988 (N_17988,N_15205,N_15827);
xnor U17989 (N_17989,N_14063,N_14715);
and U17990 (N_17990,N_15991,N_14701);
nand U17991 (N_17991,N_14871,N_15777);
xor U17992 (N_17992,N_14284,N_15158);
nor U17993 (N_17993,N_14580,N_15296);
or U17994 (N_17994,N_14931,N_15060);
and U17995 (N_17995,N_14494,N_14305);
nand U17996 (N_17996,N_14426,N_15574);
nor U17997 (N_17997,N_14888,N_15523);
or U17998 (N_17998,N_15320,N_15292);
nor U17999 (N_17999,N_14474,N_15885);
nor U18000 (N_18000,N_17299,N_17016);
xnor U18001 (N_18001,N_17807,N_16199);
nand U18002 (N_18002,N_17477,N_17968);
xor U18003 (N_18003,N_16736,N_17028);
and U18004 (N_18004,N_17543,N_16061);
and U18005 (N_18005,N_17263,N_16322);
xor U18006 (N_18006,N_16975,N_16896);
nand U18007 (N_18007,N_16688,N_16841);
nor U18008 (N_18008,N_16514,N_16050);
and U18009 (N_18009,N_16887,N_16918);
xnor U18010 (N_18010,N_17893,N_17230);
nand U18011 (N_18011,N_17170,N_17873);
nand U18012 (N_18012,N_16861,N_16686);
and U18013 (N_18013,N_17582,N_16234);
nor U18014 (N_18014,N_16992,N_17800);
xor U18015 (N_18015,N_17554,N_17812);
and U18016 (N_18016,N_17720,N_16373);
or U18017 (N_18017,N_17247,N_17441);
nor U18018 (N_18018,N_16340,N_17465);
nor U18019 (N_18019,N_16266,N_17594);
and U18020 (N_18020,N_17446,N_17516);
xnor U18021 (N_18021,N_16761,N_17671);
nor U18022 (N_18022,N_17866,N_16518);
nor U18023 (N_18023,N_16549,N_17875);
and U18024 (N_18024,N_17082,N_16201);
and U18025 (N_18025,N_16587,N_17957);
nand U18026 (N_18026,N_16353,N_16468);
xnor U18027 (N_18027,N_16030,N_16315);
and U18028 (N_18028,N_16123,N_17488);
nand U18029 (N_18029,N_16959,N_17047);
xnor U18030 (N_18030,N_16693,N_16342);
and U18031 (N_18031,N_16239,N_17117);
and U18032 (N_18032,N_17819,N_17851);
nor U18033 (N_18033,N_17629,N_16140);
nor U18034 (N_18034,N_16594,N_16306);
or U18035 (N_18035,N_17002,N_16742);
or U18036 (N_18036,N_17176,N_16296);
or U18037 (N_18037,N_17288,N_17559);
xnor U18038 (N_18038,N_16665,N_16560);
and U18039 (N_18039,N_17236,N_16211);
and U18040 (N_18040,N_17502,N_17788);
nand U18041 (N_18041,N_16557,N_16161);
nand U18042 (N_18042,N_16247,N_16104);
nor U18043 (N_18043,N_17798,N_16631);
nand U18044 (N_18044,N_17626,N_17769);
xnor U18045 (N_18045,N_16949,N_16605);
and U18046 (N_18046,N_17311,N_16085);
and U18047 (N_18047,N_17303,N_16544);
xor U18048 (N_18048,N_17237,N_17436);
xnor U18049 (N_18049,N_16596,N_16777);
nand U18050 (N_18050,N_17621,N_16607);
nor U18051 (N_18051,N_16370,N_17438);
xnor U18052 (N_18052,N_16972,N_17512);
nand U18053 (N_18053,N_16856,N_16358);
xnor U18054 (N_18054,N_16153,N_17696);
nor U18055 (N_18055,N_17903,N_16931);
or U18056 (N_18056,N_16522,N_17505);
and U18057 (N_18057,N_17432,N_16822);
and U18058 (N_18058,N_16895,N_16794);
xnor U18059 (N_18059,N_16126,N_16844);
and U18060 (N_18060,N_17442,N_17617);
nand U18061 (N_18061,N_17847,N_17894);
nor U18062 (N_18062,N_16619,N_17802);
xnor U18063 (N_18063,N_17300,N_17031);
nor U18064 (N_18064,N_16878,N_16568);
nor U18065 (N_18065,N_16954,N_16465);
nor U18066 (N_18066,N_17659,N_16865);
or U18067 (N_18067,N_17849,N_17168);
and U18068 (N_18068,N_17540,N_16305);
and U18069 (N_18069,N_16369,N_16337);
xor U18070 (N_18070,N_17218,N_16415);
nand U18071 (N_18071,N_16538,N_16964);
nand U18072 (N_18072,N_16450,N_16175);
or U18073 (N_18073,N_16111,N_17015);
or U18074 (N_18074,N_16097,N_16849);
nor U18075 (N_18075,N_16067,N_17402);
nor U18076 (N_18076,N_16937,N_16205);
and U18077 (N_18077,N_16355,N_16851);
nor U18078 (N_18078,N_16825,N_17040);
xor U18079 (N_18079,N_16729,N_16824);
or U18080 (N_18080,N_16716,N_17634);
and U18081 (N_18081,N_16169,N_16018);
and U18082 (N_18082,N_17585,N_16419);
or U18083 (N_18083,N_17815,N_17244);
and U18084 (N_18084,N_17508,N_16669);
or U18085 (N_18085,N_16252,N_16545);
and U18086 (N_18086,N_16692,N_16476);
and U18087 (N_18087,N_16280,N_17640);
xor U18088 (N_18088,N_17904,N_16267);
and U18089 (N_18089,N_16333,N_16304);
and U18090 (N_18090,N_16082,N_16566);
nand U18091 (N_18091,N_17426,N_16399);
nor U18092 (N_18092,N_16592,N_17538);
and U18093 (N_18093,N_16130,N_16830);
xor U18094 (N_18094,N_16412,N_16057);
and U18095 (N_18095,N_17937,N_16614);
and U18096 (N_18096,N_17909,N_17324);
and U18097 (N_18097,N_16022,N_16866);
xnor U18098 (N_18098,N_17868,N_17273);
nor U18099 (N_18099,N_16170,N_16970);
or U18100 (N_18100,N_17497,N_16311);
xnor U18101 (N_18101,N_16236,N_16223);
xnor U18102 (N_18102,N_17166,N_17231);
nor U18103 (N_18103,N_17032,N_16204);
or U18104 (N_18104,N_17586,N_17058);
xor U18105 (N_18105,N_17984,N_16277);
xor U18106 (N_18106,N_17569,N_17858);
or U18107 (N_18107,N_17575,N_17074);
xnor U18108 (N_18108,N_16255,N_17454);
xor U18109 (N_18109,N_16935,N_17378);
and U18110 (N_18110,N_17274,N_16441);
xor U18111 (N_18111,N_17533,N_17949);
or U18112 (N_18112,N_16681,N_17056);
or U18113 (N_18113,N_16109,N_17207);
and U18114 (N_18114,N_17782,N_17654);
or U18115 (N_18115,N_17691,N_17356);
or U18116 (N_18116,N_16754,N_17899);
and U18117 (N_18117,N_17422,N_17383);
and U18118 (N_18118,N_17752,N_16184);
xnor U18119 (N_18119,N_17456,N_16455);
and U18120 (N_18120,N_16318,N_16656);
or U18121 (N_18121,N_16100,N_17639);
xor U18122 (N_18122,N_17185,N_17776);
and U18123 (N_18123,N_16941,N_17154);
or U18124 (N_18124,N_17066,N_17081);
or U18125 (N_18125,N_16770,N_17307);
xor U18126 (N_18126,N_16135,N_16682);
nand U18127 (N_18127,N_16554,N_17805);
and U18128 (N_18128,N_16758,N_17353);
nand U18129 (N_18129,N_17572,N_16447);
nand U18130 (N_18130,N_16013,N_17319);
nor U18131 (N_18131,N_17503,N_17126);
nor U18132 (N_18132,N_16046,N_17843);
nand U18133 (N_18133,N_16214,N_16915);
xor U18134 (N_18134,N_16445,N_17820);
and U18135 (N_18135,N_16227,N_16750);
or U18136 (N_18136,N_17960,N_16490);
nand U18137 (N_18137,N_16747,N_16723);
nor U18138 (N_18138,N_17914,N_17862);
xor U18139 (N_18139,N_16558,N_16722);
nor U18140 (N_18140,N_17388,N_17605);
and U18141 (N_18141,N_17315,N_17260);
or U18142 (N_18142,N_16038,N_16217);
nand U18143 (N_18143,N_16299,N_17774);
nor U18144 (N_18144,N_17528,N_16833);
or U18145 (N_18145,N_17008,N_17039);
xnor U18146 (N_18146,N_16623,N_17114);
or U18147 (N_18147,N_16696,N_17712);
or U18148 (N_18148,N_16584,N_17200);
or U18149 (N_18149,N_17033,N_16483);
nor U18150 (N_18150,N_17547,N_17293);
nor U18151 (N_18151,N_17487,N_17272);
and U18152 (N_18152,N_17332,N_16933);
nand U18153 (N_18153,N_17208,N_16843);
xor U18154 (N_18154,N_16049,N_16238);
or U18155 (N_18155,N_16570,N_17053);
xnor U18156 (N_18156,N_16690,N_17881);
nand U18157 (N_18157,N_16640,N_16601);
xnor U18158 (N_18158,N_16071,N_17956);
and U18159 (N_18159,N_16287,N_16102);
nand U18160 (N_18160,N_16341,N_17989);
nor U18161 (N_18161,N_16927,N_16569);
or U18162 (N_18162,N_17616,N_17418);
and U18163 (N_18163,N_16683,N_16814);
xnor U18164 (N_18164,N_16995,N_16733);
nand U18165 (N_18165,N_17146,N_16962);
xnor U18166 (N_18166,N_16114,N_17281);
nor U18167 (N_18167,N_17202,N_17558);
nand U18168 (N_18168,N_17062,N_16948);
xnor U18169 (N_18169,N_16352,N_17323);
and U18170 (N_18170,N_16826,N_16783);
nand U18171 (N_18171,N_16414,N_17832);
xnor U18172 (N_18172,N_17337,N_16892);
xnor U18173 (N_18173,N_16345,N_17211);
and U18174 (N_18174,N_17308,N_17745);
or U18175 (N_18175,N_17024,N_16986);
nand U18176 (N_18176,N_17048,N_17700);
xor U18177 (N_18177,N_17362,N_17596);
and U18178 (N_18178,N_17334,N_16324);
nand U18179 (N_18179,N_17717,N_17125);
and U18180 (N_18180,N_17359,N_17997);
or U18181 (N_18181,N_17287,N_17987);
and U18182 (N_18182,N_17797,N_17859);
xnor U18183 (N_18183,N_16746,N_17922);
xnor U18184 (N_18184,N_16885,N_17553);
or U18185 (N_18185,N_16137,N_17913);
and U18186 (N_18186,N_17496,N_16491);
xnor U18187 (N_18187,N_16606,N_17493);
xnor U18188 (N_18188,N_16612,N_16743);
or U18189 (N_18189,N_17076,N_16738);
and U18190 (N_18190,N_16982,N_16916);
nand U18191 (N_18191,N_17612,N_17112);
nand U18192 (N_18192,N_16556,N_17761);
or U18193 (N_18193,N_17719,N_16157);
xnor U18194 (N_18194,N_17004,N_17734);
and U18195 (N_18195,N_16543,N_16804);
xor U18196 (N_18196,N_17233,N_17980);
or U18197 (N_18197,N_16293,N_17063);
xor U18198 (N_18198,N_16854,N_16620);
nand U18199 (N_18199,N_17365,N_17938);
xor U18200 (N_18200,N_16232,N_17119);
or U18201 (N_18201,N_16479,N_17374);
nor U18202 (N_18202,N_16245,N_17361);
nand U18203 (N_18203,N_16151,N_17035);
nand U18204 (N_18204,N_16260,N_16210);
or U18205 (N_18205,N_17628,N_16537);
nand U18206 (N_18206,N_16624,N_16098);
and U18207 (N_18207,N_16703,N_16166);
xnor U18208 (N_18208,N_17204,N_17759);
or U18209 (N_18209,N_16812,N_16350);
nor U18210 (N_18210,N_17565,N_17291);
or U18211 (N_18211,N_17013,N_17742);
nor U18212 (N_18212,N_17445,N_16721);
and U18213 (N_18213,N_17216,N_16590);
nor U18214 (N_18214,N_17789,N_16903);
nand U18215 (N_18215,N_17919,N_16105);
nor U18216 (N_18216,N_16025,N_17182);
and U18217 (N_18217,N_16857,N_16752);
or U18218 (N_18218,N_16712,N_17138);
nor U18219 (N_18219,N_17557,N_16346);
nand U18220 (N_18220,N_17526,N_17672);
nor U18221 (N_18221,N_16519,N_17305);
or U18222 (N_18222,N_17682,N_17998);
or U18223 (N_18223,N_17986,N_16430);
nor U18224 (N_18224,N_16081,N_16165);
and U18225 (N_18225,N_16993,N_16460);
or U18226 (N_18226,N_16636,N_16316);
xor U18227 (N_18227,N_16778,N_16384);
nor U18228 (N_18228,N_16110,N_16326);
nand U18229 (N_18229,N_17132,N_17971);
xor U18230 (N_18230,N_16446,N_16036);
or U18231 (N_18231,N_17129,N_17725);
nand U18232 (N_18232,N_16372,N_16839);
nor U18233 (N_18233,N_16477,N_17990);
or U18234 (N_18234,N_17923,N_16871);
or U18235 (N_18235,N_16862,N_17666);
or U18236 (N_18236,N_16835,N_17088);
nor U18237 (N_18237,N_16732,N_17049);
xor U18238 (N_18238,N_17107,N_16595);
nor U18239 (N_18239,N_17799,N_17555);
xor U18240 (N_18240,N_17243,N_17195);
and U18241 (N_18241,N_17282,N_16883);
nor U18242 (N_18242,N_16443,N_17622);
nand U18243 (N_18243,N_17214,N_17384);
and U18244 (N_18244,N_17609,N_17579);
or U18245 (N_18245,N_16968,N_17395);
nor U18246 (N_18246,N_17372,N_17886);
xor U18247 (N_18247,N_16759,N_16695);
xnor U18248 (N_18248,N_16344,N_17698);
nor U18249 (N_18249,N_17552,N_17642);
and U18250 (N_18250,N_17366,N_17743);
and U18251 (N_18251,N_16760,N_16630);
nand U18252 (N_18252,N_17163,N_17994);
and U18253 (N_18253,N_17226,N_16409);
and U18254 (N_18254,N_17522,N_16449);
xnor U18255 (N_18255,N_16128,N_17905);
nor U18256 (N_18256,N_17780,N_17452);
nand U18257 (N_18257,N_17958,N_17327);
and U18258 (N_18258,N_16043,N_17775);
nor U18259 (N_18259,N_16437,N_16579);
xor U18260 (N_18260,N_16610,N_16901);
nor U18261 (N_18261,N_17785,N_17674);
or U18262 (N_18262,N_16718,N_16107);
or U18263 (N_18263,N_16454,N_17751);
nand U18264 (N_18264,N_17570,N_17965);
or U18265 (N_18265,N_17412,N_17706);
xor U18266 (N_18266,N_17294,N_16063);
nand U18267 (N_18267,N_16108,N_17153);
nor U18268 (N_18268,N_16652,N_16991);
or U18269 (N_18269,N_17094,N_16699);
or U18270 (N_18270,N_16406,N_16094);
and U18271 (N_18271,N_16662,N_17246);
nor U18272 (N_18272,N_16563,N_16495);
or U18273 (N_18273,N_16088,N_17702);
and U18274 (N_18274,N_16797,N_16325);
or U18275 (N_18275,N_17673,N_17003);
and U18276 (N_18276,N_17993,N_17590);
nor U18277 (N_18277,N_17173,N_17373);
and U18278 (N_18278,N_17045,N_16354);
or U18279 (N_18279,N_16789,N_16782);
and U18280 (N_18280,N_17637,N_17977);
nor U18281 (N_18281,N_17150,N_16235);
or U18282 (N_18282,N_16766,N_16578);
and U18283 (N_18283,N_16946,N_16881);
nand U18284 (N_18284,N_17517,N_17038);
nor U18285 (N_18285,N_17005,N_17145);
nand U18286 (N_18286,N_16654,N_16188);
and U18287 (N_18287,N_16378,N_16575);
xnor U18288 (N_18288,N_16251,N_16075);
xor U18289 (N_18289,N_16428,N_17128);
nand U18290 (N_18290,N_17541,N_16600);
nand U18291 (N_18291,N_17917,N_16942);
nand U18292 (N_18292,N_16668,N_16106);
nand U18293 (N_18293,N_17001,N_17969);
or U18294 (N_18294,N_16648,N_17205);
or U18295 (N_18295,N_17277,N_17421);
nand U18296 (N_18296,N_17576,N_17695);
nor U18297 (N_18297,N_16228,N_16643);
xnor U18298 (N_18298,N_16134,N_17587);
nor U18299 (N_18299,N_17492,N_16509);
or U18300 (N_18300,N_17275,N_17343);
nor U18301 (N_18301,N_17762,N_17827);
or U18302 (N_18302,N_16837,N_16178);
nor U18303 (N_18303,N_17222,N_17865);
or U18304 (N_18304,N_16285,N_17018);
xnor U18305 (N_18305,N_16499,N_17321);
or U18306 (N_18306,N_17861,N_17228);
xor U18307 (N_18307,N_16086,N_17724);
xnor U18308 (N_18308,N_17408,N_16216);
xor U18309 (N_18309,N_17611,N_17618);
or U18310 (N_18310,N_17765,N_16513);
and U18311 (N_18311,N_17556,N_16504);
nor U18312 (N_18312,N_16850,N_17283);
xnor U18313 (N_18313,N_16027,N_17741);
and U18314 (N_18314,N_16259,N_16039);
and U18315 (N_18315,N_17346,N_16016);
nand U18316 (N_18316,N_16551,N_17597);
or U18317 (N_18317,N_16290,N_16113);
or U18318 (N_18318,N_16374,N_16250);
nand U18319 (N_18319,N_17511,N_16142);
nor U18320 (N_18320,N_16967,N_17813);
nand U18321 (N_18321,N_16221,N_16158);
nand U18322 (N_18322,N_17479,N_17007);
and U18323 (N_18323,N_16307,N_17602);
nand U18324 (N_18324,N_17021,N_17921);
nand U18325 (N_18325,N_17836,N_16055);
xnor U18326 (N_18326,N_16459,N_17783);
and U18327 (N_18327,N_17846,N_16160);
nand U18328 (N_18328,N_17889,N_17407);
nor U18329 (N_18329,N_17793,N_16740);
or U18330 (N_18330,N_17073,N_17023);
or U18331 (N_18331,N_17221,N_17855);
nand U18332 (N_18332,N_17437,N_16427);
nor U18333 (N_18333,N_16001,N_16112);
or U18334 (N_18334,N_17701,N_17000);
and U18335 (N_18335,N_16131,N_17506);
nand U18336 (N_18336,N_17747,N_16559);
nor U18337 (N_18337,N_17241,N_16377);
and U18338 (N_18338,N_17703,N_17382);
nor U18339 (N_18339,N_16505,N_16198);
nor U18340 (N_18340,N_16727,N_16263);
nand U18341 (N_18341,N_16541,N_16371);
or U18342 (N_18342,N_16626,N_16283);
xor U18343 (N_18343,N_16803,N_17856);
nor U18344 (N_18344,N_17514,N_17726);
and U18345 (N_18345,N_16502,N_16405);
xnor U18346 (N_18346,N_16663,N_16254);
and U18347 (N_18347,N_16133,N_17947);
or U18348 (N_18348,N_16737,N_17255);
xnor U18349 (N_18349,N_17190,N_16748);
nand U18350 (N_18350,N_16339,N_17995);
xnor U18351 (N_18351,N_16674,N_16385);
nand U18352 (N_18352,N_17106,N_17464);
xor U18353 (N_18353,N_16336,N_16842);
nand U18354 (N_18354,N_17790,N_17310);
nand U18355 (N_18355,N_17380,N_17883);
xnor U18356 (N_18356,N_17268,N_16388);
or U18357 (N_18357,N_17369,N_17261);
and U18358 (N_18358,N_17444,N_17439);
nor U18359 (N_18359,N_16950,N_16434);
xnor U18360 (N_18360,N_17649,N_16567);
and U18361 (N_18361,N_16909,N_17959);
nand U18362 (N_18362,N_17093,N_17684);
or U18363 (N_18363,N_17071,N_16642);
nand U18364 (N_18364,N_17735,N_16660);
and U18365 (N_18365,N_17070,N_16395);
or U18366 (N_18366,N_17091,N_17580);
nor U18367 (N_18367,N_16202,N_16284);
or U18368 (N_18368,N_17826,N_17060);
and U18369 (N_18369,N_16691,N_16646);
or U18370 (N_18370,N_17838,N_16951);
or U18371 (N_18371,N_17962,N_17095);
nand U18372 (N_18372,N_16528,N_16319);
xor U18373 (N_18373,N_16571,N_17668);
xnor U18374 (N_18374,N_17396,N_16297);
nor U18375 (N_18375,N_16422,N_17416);
xnor U18376 (N_18376,N_17518,N_17571);
and U18377 (N_18377,N_16507,N_16368);
xnor U18378 (N_18378,N_16772,N_17970);
nor U18379 (N_18379,N_16029,N_16226);
or U18380 (N_18380,N_16091,N_17227);
nand U18381 (N_18381,N_16832,N_17925);
or U18382 (N_18382,N_17803,N_17086);
or U18383 (N_18383,N_16291,N_16886);
xnor U18384 (N_18384,N_17413,N_17607);
and U18385 (N_18385,N_16731,N_17489);
nand U18386 (N_18386,N_16220,N_16320);
or U18387 (N_18387,N_16979,N_16180);
or U18388 (N_18388,N_17860,N_16125);
or U18389 (N_18389,N_17924,N_16819);
or U18390 (N_18390,N_16894,N_17055);
or U18391 (N_18391,N_16185,N_17447);
and U18392 (N_18392,N_17911,N_16553);
or U18393 (N_18393,N_16080,N_16420);
or U18394 (N_18394,N_16791,N_16511);
xor U18395 (N_18395,N_16257,N_16521);
nor U18396 (N_18396,N_16990,N_16079);
or U18397 (N_18397,N_16035,N_17061);
nor U18398 (N_18398,N_16644,N_16302);
nand U18399 (N_18399,N_16998,N_16795);
xor U18400 (N_18400,N_16884,N_17850);
and U18401 (N_18401,N_17581,N_16829);
nand U18402 (N_18402,N_17306,N_17219);
xnor U18403 (N_18403,N_16321,N_16963);
xnor U18404 (N_18404,N_16853,N_17072);
xor U18405 (N_18405,N_16241,N_17834);
or U18406 (N_18406,N_17895,N_16928);
or U18407 (N_18407,N_16664,N_16390);
xor U18408 (N_18408,N_17186,N_17157);
and U18409 (N_18409,N_17907,N_17583);
nand U18410 (N_18410,N_16003,N_17728);
nor U18411 (N_18411,N_17852,N_16520);
nand U18412 (N_18412,N_17767,N_17665);
xor U18413 (N_18413,N_16658,N_17317);
and U18414 (N_18414,N_16516,N_16313);
nor U18415 (N_18415,N_16880,N_16429);
xor U18416 (N_18416,N_17561,N_17951);
nand U18417 (N_18417,N_16059,N_16197);
and U18418 (N_18418,N_16855,N_17213);
and U18419 (N_18419,N_17364,N_17390);
or U18420 (N_18420,N_16966,N_17501);
and U18421 (N_18421,N_16264,N_17954);
or U18422 (N_18422,N_16739,N_17030);
and U18423 (N_18423,N_17297,N_16168);
nand U18424 (N_18424,N_16670,N_17768);
nor U18425 (N_18425,N_16701,N_16467);
nor U18426 (N_18426,N_16816,N_17285);
nor U18427 (N_18427,N_17292,N_17089);
and U18428 (N_18428,N_17469,N_16510);
nor U18429 (N_18429,N_17485,N_17593);
nor U18430 (N_18430,N_17839,N_17036);
and U18431 (N_18431,N_17972,N_17286);
or U18432 (N_18432,N_17351,N_17521);
nor U18433 (N_18433,N_17338,N_17270);
and U18434 (N_18434,N_16529,N_17451);
nor U18435 (N_18435,N_17916,N_16805);
nand U18436 (N_18436,N_16763,N_17652);
nor U18437 (N_18437,N_17874,N_17758);
and U18438 (N_18438,N_17491,N_17052);
or U18439 (N_18439,N_16181,N_17624);
and U18440 (N_18440,N_16162,N_17795);
nor U18441 (N_18441,N_17127,N_17755);
nand U18442 (N_18442,N_16700,N_16191);
xor U18443 (N_18443,N_17116,N_16464);
or U18444 (N_18444,N_17159,N_16172);
and U18445 (N_18445,N_17635,N_17314);
and U18446 (N_18446,N_17817,N_17738);
nand U18447 (N_18447,N_17209,N_16536);
or U18448 (N_18448,N_17316,N_16119);
or U18449 (N_18449,N_17867,N_17131);
nand U18450 (N_18450,N_16484,N_17080);
and U18451 (N_18451,N_17906,N_16776);
and U18452 (N_18452,N_16376,N_16045);
and U18453 (N_18453,N_16099,N_16195);
nor U18454 (N_18454,N_17011,N_16327);
nor U18455 (N_18455,N_17375,N_17620);
and U18456 (N_18456,N_17651,N_16637);
nand U18457 (N_18457,N_16093,N_17474);
nand U18458 (N_18458,N_16847,N_16332);
xnor U18459 (N_18459,N_16070,N_16042);
or U18460 (N_18460,N_17676,N_16194);
xnor U18461 (N_18461,N_17660,N_17896);
nor U18462 (N_18462,N_16249,N_16303);
or U18463 (N_18463,N_17462,N_17941);
nor U18464 (N_18464,N_16011,N_17425);
xor U18465 (N_18465,N_17796,N_17471);
nor U18466 (N_18466,N_16064,N_16143);
nor U18467 (N_18467,N_17863,N_16244);
nor U18468 (N_18468,N_17713,N_17589);
nor U18469 (N_18469,N_17428,N_17026);
nor U18470 (N_18470,N_16478,N_16715);
nand U18471 (N_18471,N_16628,N_17619);
nand U18472 (N_18472,N_16934,N_16010);
xor U18473 (N_18473,N_16347,N_16047);
xnor U18474 (N_18474,N_17876,N_16889);
xnor U18475 (N_18475,N_17433,N_17169);
nor U18476 (N_18476,N_17870,N_16209);
nand U18477 (N_18477,N_17885,N_16989);
or U18478 (N_18478,N_16281,N_17367);
or U18479 (N_18479,N_16497,N_16083);
nand U18480 (N_18480,N_16383,N_16831);
xor U18481 (N_18481,N_17625,N_16481);
nor U18482 (N_18482,N_17239,N_16330);
nand U18483 (N_18483,N_17644,N_17358);
nand U18484 (N_18484,N_17973,N_17705);
and U18485 (N_18485,N_17662,N_16159);
or U18486 (N_18486,N_16980,N_17225);
and U18487 (N_18487,N_16547,N_16391);
nand U18488 (N_18488,N_17804,N_16815);
nor U18489 (N_18489,N_17101,N_16604);
nand U18490 (N_18490,N_17449,N_17406);
and U18491 (N_18491,N_17431,N_16418);
nor U18492 (N_18492,N_17584,N_16279);
nor U18493 (N_18493,N_17171,N_17523);
and U18494 (N_18494,N_16356,N_17256);
nand U18495 (N_18495,N_17423,N_16393);
nand U18496 (N_18496,N_17398,N_17453);
nand U18497 (N_18497,N_17068,N_17099);
or U18498 (N_18498,N_16425,N_16867);
nand U18499 (N_18499,N_16882,N_16359);
nand U18500 (N_18500,N_16734,N_17155);
nand U18501 (N_18501,N_17842,N_17857);
nor U18502 (N_18502,N_17535,N_16751);
or U18503 (N_18503,N_17187,N_17296);
nor U18504 (N_18504,N_17473,N_17403);
nor U18505 (N_18505,N_16037,N_16486);
nand U18506 (N_18506,N_16271,N_16394);
nor U18507 (N_18507,N_16863,N_16349);
or U18508 (N_18508,N_16403,N_16453);
or U18509 (N_18509,N_17120,N_16720);
xor U18510 (N_18510,N_17687,N_16961);
and U18511 (N_18511,N_17495,N_17429);
xnor U18512 (N_18512,N_16456,N_17961);
nand U18513 (N_18513,N_16506,N_16402);
and U18514 (N_18514,N_16936,N_16877);
xor U18515 (N_18515,N_16820,N_17050);
or U18516 (N_18516,N_16807,N_16404);
nor U18517 (N_18517,N_17996,N_17830);
nor U18518 (N_18518,N_16526,N_17900);
xor U18519 (N_18519,N_17191,N_16233);
xor U18520 (N_18520,N_17242,N_16410);
nor U18521 (N_18521,N_16956,N_16955);
nor U18522 (N_18522,N_17918,N_17808);
or U18523 (N_18523,N_17313,N_17257);
xor U18524 (N_18524,N_17262,N_16586);
xnor U18525 (N_18525,N_17302,N_17065);
xor U18526 (N_18526,N_16762,N_16196);
xnor U18527 (N_18527,N_16019,N_17198);
xnor U18528 (N_18528,N_17766,N_17588);
and U18529 (N_18529,N_17633,N_16470);
xnor U18530 (N_18530,N_16078,N_17463);
xor U18531 (N_18531,N_16176,N_16472);
nor U18532 (N_18532,N_17295,N_17678);
or U18533 (N_18533,N_17494,N_16496);
nand U18534 (N_18534,N_17560,N_16627);
and U18535 (N_18535,N_16957,N_17711);
or U18536 (N_18536,N_16407,N_16103);
nand U18537 (N_18537,N_17848,N_16095);
or U18538 (N_18538,N_16845,N_16069);
nor U18539 (N_18539,N_16120,N_17475);
nand U18540 (N_18540,N_16523,N_16163);
and U18541 (N_18541,N_16367,N_17017);
and U18542 (N_18542,N_16002,N_16489);
nor U18543 (N_18543,N_17199,N_16268);
nand U18544 (N_18544,N_17733,N_17212);
and U18545 (N_18545,N_16294,N_16146);
nand U18546 (N_18546,N_17680,N_17232);
nor U18547 (N_18547,N_17536,N_17670);
nor U18548 (N_18548,N_17709,N_17598);
and U18549 (N_18549,N_17342,N_16308);
nand U18550 (N_18550,N_16629,N_16508);
nor U18551 (N_18551,N_16246,N_16334);
xor U18552 (N_18552,N_17884,N_16911);
xor U18553 (N_18553,N_16741,N_17087);
xor U18554 (N_18554,N_17051,N_16440);
nand U18555 (N_18555,N_17340,N_17936);
nor U18556 (N_18556,N_17841,N_16634);
or U18557 (N_18557,N_17215,N_17203);
or U18558 (N_18558,N_16331,N_17147);
nor U18559 (N_18559,N_16953,N_16338);
or U18560 (N_18560,N_17266,N_17304);
and U18561 (N_18561,N_16532,N_17410);
and U18562 (N_18562,N_17764,N_17392);
nand U18563 (N_18563,N_17542,N_17109);
nand U18564 (N_18564,N_16540,N_17641);
xnor U18565 (N_18565,N_17771,N_17650);
and U18566 (N_18566,N_17606,N_17945);
nand U18567 (N_18567,N_17891,N_17164);
nand U18568 (N_18568,N_16984,N_17520);
nor U18569 (N_18569,N_17991,N_16300);
xnor U18570 (N_18570,N_16288,N_16651);
and U18571 (N_18571,N_16597,N_17483);
nand U18572 (N_18572,N_16432,N_17638);
and U18573 (N_18573,N_16122,N_16698);
nor U18574 (N_18574,N_16190,N_16398);
or U18575 (N_18575,N_17245,N_17686);
xor U18576 (N_18576,N_17054,N_16118);
and U18577 (N_18577,N_16744,N_16771);
nand U18578 (N_18578,N_16893,N_16997);
nand U18579 (N_18579,N_16272,N_16421);
nor U18580 (N_18580,N_16392,N_17537);
nand U18581 (N_18581,N_16348,N_16977);
nand U18582 (N_18582,N_17910,N_17545);
and U18583 (N_18583,N_17577,N_16375);
nand U18584 (N_18584,N_17006,N_17509);
nand U18585 (N_18585,N_16177,N_17335);
or U18586 (N_18586,N_16564,N_17175);
nor U18587 (N_18587,N_16756,N_17835);
or U18588 (N_18588,N_16117,N_17544);
xnor U18589 (N_18589,N_17902,N_16387);
nor U18590 (N_18590,N_17044,N_17331);
xor U18591 (N_18591,N_16562,N_17604);
nor U18592 (N_18592,N_17196,N_16360);
xnor U18593 (N_18593,N_16275,N_17427);
xor U18594 (N_18594,N_17248,N_16174);
xor U18595 (N_18595,N_16243,N_17756);
and U18596 (N_18596,N_16021,N_17411);
and U18597 (N_18597,N_17118,N_16574);
xor U18598 (N_18598,N_16719,N_17124);
nand U18599 (N_18599,N_16138,N_17329);
or U18600 (N_18600,N_17144,N_16952);
nor U18601 (N_18601,N_17946,N_16786);
or U18602 (N_18602,N_16416,N_16498);
or U18603 (N_18603,N_17882,N_16056);
nor U18604 (N_18604,N_16999,N_16048);
or U18605 (N_18605,N_16906,N_17754);
or U18606 (N_18606,N_17880,N_16973);
and U18607 (N_18607,N_16785,N_16276);
or U18608 (N_18608,N_17376,N_17539);
nor U18609 (N_18609,N_16436,N_17908);
nor U18610 (N_18610,N_16066,N_17928);
xnor U18611 (N_18611,N_17854,N_17699);
or U18612 (N_18612,N_16473,N_17950);
nor U18613 (N_18613,N_17172,N_16458);
xnor U18614 (N_18614,N_16074,N_16366);
or U18615 (N_18615,N_16488,N_16269);
or U18616 (N_18616,N_17963,N_16524);
and U18617 (N_18617,N_16902,N_16397);
nand U18618 (N_18618,N_17077,N_16565);
or U18619 (N_18619,N_16981,N_17265);
and U18620 (N_18620,N_17763,N_16728);
and U18621 (N_18621,N_16400,N_17352);
xor U18622 (N_18622,N_16004,N_17507);
nand U18623 (N_18623,N_16647,N_16714);
xnor U18624 (N_18624,N_17822,N_16167);
nor U18625 (N_18625,N_17692,N_17357);
nor U18626 (N_18626,N_17791,N_17948);
nor U18627 (N_18627,N_17809,N_16846);
nor U18628 (N_18628,N_16020,N_16539);
nor U18629 (N_18629,N_16357,N_17193);
or U18630 (N_18630,N_17974,N_16753);
or U18631 (N_18631,N_17363,N_17929);
nand U18632 (N_18632,N_16875,N_17632);
and U18633 (N_18633,N_17550,N_17636);
xnor U18634 (N_18634,N_16677,N_16608);
or U18635 (N_18635,N_16225,N_16485);
and U18636 (N_18636,N_17148,N_16230);
nand U18637 (N_18637,N_17685,N_17325);
nand U18638 (N_18638,N_17600,N_16312);
or U18639 (N_18639,N_16278,N_16919);
or U18640 (N_18640,N_17529,N_16828);
and U18641 (N_18641,N_16917,N_17610);
nand U18642 (N_18642,N_16840,N_17664);
or U18643 (N_18643,N_17389,N_16796);
or U18644 (N_18644,N_16218,N_16983);
xnor U18645 (N_18645,N_16033,N_16775);
or U18646 (N_18646,N_17057,N_17669);
or U18647 (N_18647,N_16779,N_17794);
nand U18648 (N_18648,N_17476,N_16207);
or U18649 (N_18649,N_16248,N_17940);
and U18650 (N_18650,N_16438,N_17689);
and U18651 (N_18651,N_17723,N_17320);
or U18652 (N_18652,N_17810,N_17490);
and U18653 (N_18653,N_17746,N_16411);
nor U18654 (N_18654,N_16905,N_16148);
or U18655 (N_18655,N_17714,N_16672);
xor U18656 (N_18656,N_16589,N_16920);
xor U18657 (N_18657,N_16452,N_16193);
xor U18658 (N_18658,N_16041,N_16707);
nand U18659 (N_18659,N_17524,N_17141);
nand U18660 (N_18660,N_16351,N_17111);
and U18661 (N_18661,N_17981,N_16869);
and U18662 (N_18662,N_16076,N_16155);
nand U18663 (N_18663,N_17130,N_16965);
nand U18664 (N_18664,N_17748,N_16784);
nand U18665 (N_18665,N_17934,N_16710);
nand U18666 (N_18666,N_17663,N_16859);
or U18667 (N_18667,N_16694,N_17530);
and U18668 (N_18668,N_16073,N_17419);
xnor U18669 (N_18669,N_17892,N_16958);
and U18670 (N_18670,N_17760,N_16602);
nand U18671 (N_18671,N_17653,N_16611);
nor U18672 (N_18672,N_17280,N_17400);
or U18673 (N_18673,N_16213,N_16527);
xnor U18674 (N_18674,N_16792,N_17098);
xnor U18675 (N_18675,N_16676,N_17103);
nor U18676 (N_18676,N_16380,N_17704);
nand U18677 (N_18677,N_17818,N_17440);
and U18678 (N_18678,N_16317,N_16872);
and U18679 (N_18679,N_17786,N_16147);
or U18680 (N_18680,N_16386,N_16132);
or U18681 (N_18681,N_16960,N_17531);
and U18682 (N_18682,N_17677,N_16127);
nand U18683 (N_18683,N_16426,N_16899);
xnor U18684 (N_18684,N_17391,N_17096);
or U18685 (N_18685,N_17059,N_16687);
or U18686 (N_18686,N_16706,N_16994);
xnor U18687 (N_18687,N_16650,N_16530);
nand U18688 (N_18688,N_16577,N_16768);
nor U18689 (N_18689,N_17234,N_16381);
xnor U18690 (N_18690,N_17468,N_17189);
xor U18691 (N_18691,N_16800,N_16335);
or U18692 (N_18692,N_17935,N_16408);
nor U18693 (N_18693,N_16591,N_16799);
xor U18694 (N_18694,N_17979,N_17551);
and U18695 (N_18695,N_16187,N_16939);
nor U18696 (N_18696,N_16535,N_17301);
and U18697 (N_18697,N_16183,N_16724);
and U18698 (N_18698,N_17646,N_16769);
nand U18699 (N_18699,N_16765,N_17694);
and U18700 (N_18700,N_16976,N_17042);
or U18701 (N_18701,N_17271,N_17944);
nor U18702 (N_18702,N_17546,N_16077);
nand U18703 (N_18703,N_16542,N_16811);
xnor U18704 (N_18704,N_17566,N_16996);
xor U18705 (N_18705,N_17484,N_16874);
or U18706 (N_18706,N_16343,N_16115);
or U18707 (N_18707,N_17716,N_17955);
and U18708 (N_18708,N_17259,N_17890);
nand U18709 (N_18709,N_17603,N_16907);
nor U18710 (N_18710,N_16657,N_16735);
or U18711 (N_18711,N_16396,N_17184);
nor U18712 (N_18712,N_17739,N_16534);
xor U18713 (N_18713,N_17010,N_17278);
and U18714 (N_18714,N_17252,N_17344);
nor U18715 (N_18715,N_16179,N_17753);
and U18716 (N_18716,N_17201,N_17727);
xor U18717 (N_18717,N_16781,N_17814);
nor U18718 (N_18718,N_17253,N_16617);
or U18719 (N_18719,N_16680,N_16615);
nor U18720 (N_18720,N_17210,N_17083);
xor U18721 (N_18721,N_16200,N_17014);
or U18722 (N_18722,N_16908,N_16689);
nand U18723 (N_18723,N_17869,N_16625);
xnor U18724 (N_18724,N_16898,N_16500);
nand U18725 (N_18725,N_17085,N_17887);
nand U18726 (N_18726,N_17975,N_17988);
nand U18727 (N_18727,N_17450,N_17041);
nor U18728 (N_18728,N_16090,N_17330);
or U18729 (N_18729,N_17710,N_16834);
and U18730 (N_18730,N_16622,N_17688);
xor U18731 (N_18731,N_17417,N_17177);
and U18732 (N_18732,N_16224,N_17149);
or U18733 (N_18733,N_17415,N_16868);
nand U18734 (N_18734,N_17414,N_16032);
nor U18735 (N_18735,N_16978,N_17568);
xor U18736 (N_18736,N_17387,N_17264);
nand U18737 (N_18737,N_16988,N_17467);
nor U18738 (N_18738,N_16024,N_16860);
xor U18739 (N_18739,N_17901,N_16129);
xor U18740 (N_18740,N_16666,N_16969);
xor U18741 (N_18741,N_16708,N_16145);
and U18742 (N_18742,N_16362,N_16633);
or U18743 (N_18743,N_16154,N_17912);
and U18744 (N_18744,N_16096,N_17837);
nand U18745 (N_18745,N_17615,N_16469);
nand U18746 (N_18746,N_17133,N_16023);
or U18747 (N_18747,N_17188,N_16040);
or U18748 (N_18748,N_17595,N_17844);
and U18749 (N_18749,N_16793,N_16890);
or U18750 (N_18750,N_17985,N_16767);
nor U18751 (N_18751,N_16203,N_17355);
and U18752 (N_18752,N_17864,N_16044);
xnor U18753 (N_18753,N_17368,N_16286);
nor U18754 (N_18754,N_17573,N_17269);
nor U18755 (N_18755,N_17658,N_16679);
xor U18756 (N_18756,N_16548,N_17290);
nor U18757 (N_18757,N_16661,N_17915);
nor U18758 (N_18758,N_17397,N_17339);
or U18759 (N_18759,N_16910,N_17933);
xnor U18760 (N_18760,N_16533,N_17105);
xnor U18761 (N_18761,N_16141,N_17075);
nand U18762 (N_18762,N_16301,N_17736);
nand U18763 (N_18763,N_16725,N_16121);
and U18764 (N_18764,N_17043,N_16925);
xnor U18765 (N_18765,N_17840,N_16552);
xnor U18766 (N_18766,N_17122,N_17707);
nand U18767 (N_18767,N_16987,N_16932);
and U18768 (N_18768,N_17527,N_17498);
xor U18769 (N_18769,N_16827,N_16231);
nand U18770 (N_18770,N_17137,N_17174);
and U18771 (N_18771,N_17420,N_17657);
nand U18772 (N_18772,N_16144,N_16655);
nand U18773 (N_18773,N_16572,N_17434);
nor U18774 (N_18774,N_17326,N_16219);
nand U18775 (N_18775,N_16433,N_16621);
or U18776 (N_18776,N_17435,N_17160);
and U18777 (N_18777,N_16442,N_16616);
nor U18778 (N_18778,N_16054,N_16940);
nand U18779 (N_18779,N_17647,N_17347);
and U18780 (N_18780,N_17284,N_16139);
nor U18781 (N_18781,N_16943,N_16705);
and U18782 (N_18782,N_16186,N_17757);
nand U18783 (N_18783,N_16517,N_16823);
nor U18784 (N_18784,N_16821,N_16208);
xor U18785 (N_18785,N_17009,N_17348);
and U18786 (N_18786,N_17729,N_17027);
or U18787 (N_18787,N_16053,N_17481);
xor U18788 (N_18788,N_16515,N_17627);
nor U18789 (N_18789,N_16052,N_17104);
xor U18790 (N_18790,N_17599,N_16439);
or U18791 (N_18791,N_16487,N_16424);
xnor U18792 (N_18792,N_16328,N_17386);
nand U18793 (N_18793,N_17515,N_16864);
and U18794 (N_18794,N_16282,N_16755);
xnor U18795 (N_18795,N_17878,N_17161);
and U18796 (N_18796,N_16212,N_17722);
nand U18797 (N_18797,N_17370,N_16944);
or U18798 (N_18798,N_17328,N_16482);
or U18799 (N_18799,N_16365,N_17816);
xnor U18800 (N_18800,N_17478,N_17178);
or U18801 (N_18801,N_17360,N_17480);
nor U18802 (N_18802,N_16603,N_16466);
and U18803 (N_18803,N_16101,N_17194);
or U18804 (N_18804,N_17482,N_17371);
and U18805 (N_18805,N_16493,N_16985);
xor U18806 (N_18806,N_16256,N_17667);
or U18807 (N_18807,N_16364,N_16717);
nand U18808 (N_18808,N_16164,N_17192);
nand U18809 (N_18809,N_16007,N_17549);
xor U18810 (N_18810,N_16475,N_17350);
nand U18811 (N_18811,N_16034,N_16242);
xnor U18812 (N_18812,N_16389,N_17322);
or U18813 (N_18813,N_16525,N_16704);
xor U18814 (N_18814,N_17249,N_17224);
and U18815 (N_18815,N_16582,N_16014);
xor U18816 (N_18816,N_16382,N_17134);
xnor U18817 (N_18817,N_17770,N_16323);
nor U18818 (N_18818,N_16838,N_17472);
xor U18819 (N_18819,N_16492,N_17777);
and U18820 (N_18820,N_17457,N_17534);
xnor U18821 (N_18821,N_17179,N_17254);
or U18822 (N_18822,N_16417,N_16087);
nand U18823 (N_18823,N_16599,N_17853);
nand U18824 (N_18824,N_16583,N_16790);
nor U18825 (N_18825,N_17470,N_17409);
nand U18826 (N_18826,N_16156,N_16062);
and U18827 (N_18827,N_16060,N_16031);
nor U18828 (N_18828,N_16361,N_17064);
nor U18829 (N_18829,N_17165,N_17821);
nor U18830 (N_18830,N_17336,N_17811);
nand U18831 (N_18831,N_16274,N_16089);
nand U18832 (N_18832,N_17592,N_17393);
xnor U18833 (N_18833,N_16580,N_17183);
xor U18834 (N_18834,N_16229,N_17162);
or U18835 (N_18835,N_16008,N_17926);
xor U18836 (N_18836,N_17121,N_16237);
nor U18837 (N_18837,N_16471,N_16573);
and U18838 (N_18838,N_16000,N_16474);
and U18839 (N_18839,N_17999,N_17983);
and U18840 (N_18840,N_16363,N_16808);
xnor U18841 (N_18841,N_16806,N_17732);
nor U18842 (N_18842,N_17258,N_17136);
nor U18843 (N_18843,N_17504,N_17721);
nor U18844 (N_18844,N_16051,N_16463);
nor U18845 (N_18845,N_16945,N_16295);
nor U18846 (N_18846,N_16757,N_17877);
xnor U18847 (N_18847,N_16974,N_17992);
xor U18848 (N_18848,N_17078,N_17158);
xor U18849 (N_18849,N_16206,N_16923);
nand U18850 (N_18850,N_16189,N_17379);
or U18851 (N_18851,N_17394,N_17110);
xnor U18852 (N_18852,N_16645,N_17466);
and U18853 (N_18853,N_17067,N_16684);
nand U18854 (N_18854,N_17443,N_16451);
or U18855 (N_18855,N_16938,N_16801);
xnor U18856 (N_18856,N_16270,N_16265);
nor U18857 (N_18857,N_16818,N_16310);
and U18858 (N_18858,N_16561,N_17354);
or U18859 (N_18859,N_17718,N_16836);
nand U18860 (N_18860,N_17267,N_17737);
and U18861 (N_18861,N_16912,N_16598);
xnor U18862 (N_18862,N_17888,N_16550);
nor U18863 (N_18863,N_16711,N_17567);
and U18864 (N_18864,N_17574,N_16192);
nor U18865 (N_18865,N_16653,N_17648);
and U18866 (N_18866,N_16462,N_17385);
nand U18867 (N_18867,N_17381,N_17289);
nor U18868 (N_18868,N_16124,N_17250);
nand U18869 (N_18869,N_17879,N_16667);
xor U18870 (N_18870,N_16273,N_16065);
and U18871 (N_18871,N_16017,N_16581);
nor U18872 (N_18872,N_17113,N_17298);
or U18873 (N_18873,N_16531,N_17792);
nor U18874 (N_18874,N_17715,N_17978);
or U18875 (N_18875,N_16149,N_16635);
nor U18876 (N_18876,N_16494,N_17206);
nand U18877 (N_18877,N_16173,N_17424);
xor U18878 (N_18878,N_17140,N_16084);
or U18879 (N_18879,N_16897,N_16262);
nand U18880 (N_18880,N_16150,N_17333);
or U18881 (N_18881,N_16593,N_17079);
xnor U18882 (N_18882,N_17656,N_17781);
or U18883 (N_18883,N_16924,N_16904);
or U18884 (N_18884,N_17223,N_16730);
or U18885 (N_18885,N_17037,N_17519);
nand U18886 (N_18886,N_16005,N_17180);
or U18887 (N_18887,N_17115,N_17020);
nor U18888 (N_18888,N_16298,N_17749);
and U18889 (N_18889,N_17708,N_17276);
nand U18890 (N_18890,N_17601,N_17608);
and U18891 (N_18891,N_16798,N_17591);
xnor U18892 (N_18892,N_16678,N_17845);
xnor U18893 (N_18893,N_16028,N_16749);
and U18894 (N_18894,N_16809,N_17661);
nand U18895 (N_18895,N_16618,N_16152);
and U18896 (N_18896,N_17486,N_17097);
xnor U18897 (N_18897,N_17090,N_16006);
and U18898 (N_18898,N_17029,N_16261);
and U18899 (N_18899,N_16588,N_16136);
nand U18900 (N_18900,N_17318,N_17151);
and U18901 (N_18901,N_16379,N_16713);
nand U18902 (N_18902,N_17461,N_17525);
or U18903 (N_18903,N_16503,N_17499);
nand U18904 (N_18904,N_17309,N_16930);
or U18905 (N_18905,N_17772,N_17645);
or U18906 (N_18906,N_16292,N_16921);
and U18907 (N_18907,N_16813,N_16314);
nand U18908 (N_18908,N_16116,N_16182);
and U18909 (N_18909,N_16309,N_17787);
or U18910 (N_18910,N_16764,N_17069);
nand U18911 (N_18911,N_17806,N_17240);
or U18912 (N_18912,N_16222,N_16891);
nor U18913 (N_18913,N_16171,N_17345);
nor U18914 (N_18914,N_16448,N_17779);
xor U18915 (N_18915,N_17613,N_16641);
or U18916 (N_18916,N_17927,N_17932);
and U18917 (N_18917,N_17679,N_16012);
nand U18918 (N_18918,N_17025,N_17084);
nand U18919 (N_18919,N_16092,N_16709);
nor U18920 (N_18920,N_16659,N_17238);
and U18921 (N_18921,N_17349,N_17197);
and U18922 (N_18922,N_16649,N_16745);
or U18923 (N_18923,N_16673,N_17801);
nor U18924 (N_18924,N_16922,N_17939);
nand U18925 (N_18925,N_17102,N_16848);
or U18926 (N_18926,N_16914,N_17405);
nor U18927 (N_18927,N_16858,N_17181);
or U18928 (N_18928,N_16780,N_17217);
and U18929 (N_18929,N_17744,N_17156);
nor U18930 (N_18930,N_17898,N_17341);
nor U18931 (N_18931,N_17828,N_16258);
and U18932 (N_18932,N_17510,N_17377);
and U18933 (N_18933,N_16009,N_16638);
nor U18934 (N_18934,N_16774,N_17404);
and U18935 (N_18935,N_16461,N_16702);
or U18936 (N_18936,N_16639,N_17976);
or U18937 (N_18937,N_16852,N_16685);
nor U18938 (N_18938,N_17135,N_16788);
or U18939 (N_18939,N_16971,N_16888);
xor U18940 (N_18940,N_17578,N_17831);
xor U18941 (N_18941,N_17825,N_17046);
nand U18942 (N_18942,N_17139,N_17943);
nor U18943 (N_18943,N_17614,N_16457);
nor U18944 (N_18944,N_16913,N_17931);
nor U18945 (N_18945,N_17623,N_17683);
nor U18946 (N_18946,N_16253,N_17548);
xor U18947 (N_18947,N_17823,N_16873);
and U18948 (N_18948,N_16423,N_17022);
nor U18949 (N_18949,N_16613,N_16555);
xnor U18950 (N_18950,N_16609,N_17235);
or U18951 (N_18951,N_16026,N_16671);
or U18952 (N_18952,N_16675,N_17631);
nand U18953 (N_18953,N_17953,N_16585);
or U18954 (N_18954,N_17279,N_17312);
nor U18955 (N_18955,N_17143,N_17920);
nor U18956 (N_18956,N_17630,N_17460);
nand U18957 (N_18957,N_17829,N_17532);
nand U18958 (N_18958,N_17778,N_17563);
xnor U18959 (N_18959,N_16726,N_17152);
xor U18960 (N_18960,N_17964,N_16413);
and U18961 (N_18961,N_17123,N_16802);
nand U18962 (N_18962,N_17100,N_17942);
or U18963 (N_18963,N_16435,N_17681);
xor U18964 (N_18964,N_17229,N_17399);
or U18965 (N_18965,N_17872,N_16926);
nand U18966 (N_18966,N_17401,N_16015);
and U18967 (N_18967,N_16215,N_16501);
nor U18968 (N_18968,N_17967,N_17142);
and U18969 (N_18969,N_16072,N_17643);
nor U18970 (N_18970,N_17982,N_16289);
nand U18971 (N_18971,N_17966,N_16947);
and U18972 (N_18972,N_17564,N_17430);
and U18973 (N_18973,N_17897,N_17824);
nor U18974 (N_18974,N_17655,N_16444);
or U18975 (N_18975,N_16576,N_16787);
xnor U18976 (N_18976,N_16773,N_16546);
or U18977 (N_18977,N_16879,N_16876);
xnor U18978 (N_18978,N_17012,N_17448);
nand U18979 (N_18979,N_17693,N_16632);
and U18980 (N_18980,N_16480,N_17455);
nor U18981 (N_18981,N_16929,N_17092);
and U18982 (N_18982,N_17513,N_16870);
nand U18983 (N_18983,N_17034,N_17773);
nand U18984 (N_18984,N_17730,N_17952);
nor U18985 (N_18985,N_16058,N_17167);
and U18986 (N_18986,N_16810,N_17220);
nor U18987 (N_18987,N_16817,N_17251);
and U18988 (N_18988,N_17833,N_17108);
and U18989 (N_18989,N_17750,N_17562);
nand U18990 (N_18990,N_16900,N_17930);
or U18991 (N_18991,N_16329,N_17697);
nand U18992 (N_18992,N_17740,N_17731);
xor U18993 (N_18993,N_17458,N_16240);
xnor U18994 (N_18994,N_17019,N_17871);
or U18995 (N_18995,N_16401,N_16431);
and U18996 (N_18996,N_17500,N_16068);
and U18997 (N_18997,N_17784,N_17459);
xnor U18998 (N_18998,N_17690,N_17675);
or U18999 (N_18999,N_16697,N_16512);
nand U19000 (N_19000,N_17221,N_17038);
and U19001 (N_19001,N_16721,N_16470);
and U19002 (N_19002,N_16809,N_17001);
nor U19003 (N_19003,N_17104,N_17059);
and U19004 (N_19004,N_17252,N_16432);
and U19005 (N_19005,N_16677,N_16479);
xor U19006 (N_19006,N_16222,N_17964);
nor U19007 (N_19007,N_16310,N_16350);
nand U19008 (N_19008,N_17399,N_17845);
nand U19009 (N_19009,N_17638,N_17452);
nand U19010 (N_19010,N_17058,N_16257);
and U19011 (N_19011,N_17364,N_16452);
nor U19012 (N_19012,N_17645,N_16309);
nand U19013 (N_19013,N_17773,N_16277);
nand U19014 (N_19014,N_17101,N_17968);
nand U19015 (N_19015,N_16656,N_16920);
xor U19016 (N_19016,N_16238,N_16902);
or U19017 (N_19017,N_16039,N_16591);
nand U19018 (N_19018,N_16844,N_16074);
nand U19019 (N_19019,N_17986,N_17712);
nor U19020 (N_19020,N_16214,N_17906);
nor U19021 (N_19021,N_17497,N_16176);
nand U19022 (N_19022,N_16075,N_17292);
nor U19023 (N_19023,N_16390,N_17269);
nand U19024 (N_19024,N_16759,N_17373);
nor U19025 (N_19025,N_17676,N_16728);
nor U19026 (N_19026,N_16866,N_16335);
xnor U19027 (N_19027,N_17054,N_16797);
nand U19028 (N_19028,N_17563,N_16683);
nor U19029 (N_19029,N_16001,N_16266);
and U19030 (N_19030,N_16769,N_17009);
or U19031 (N_19031,N_16498,N_16752);
nand U19032 (N_19032,N_16552,N_17558);
or U19033 (N_19033,N_16404,N_16846);
nand U19034 (N_19034,N_16334,N_16555);
nand U19035 (N_19035,N_16915,N_17552);
and U19036 (N_19036,N_16867,N_17427);
or U19037 (N_19037,N_16086,N_16140);
nand U19038 (N_19038,N_17062,N_16551);
nor U19039 (N_19039,N_16982,N_17453);
nor U19040 (N_19040,N_17592,N_17860);
nand U19041 (N_19041,N_16954,N_16092);
nor U19042 (N_19042,N_17415,N_17931);
nand U19043 (N_19043,N_17719,N_16181);
or U19044 (N_19044,N_17177,N_17072);
xor U19045 (N_19045,N_17567,N_16854);
and U19046 (N_19046,N_16615,N_16900);
or U19047 (N_19047,N_16397,N_17142);
xnor U19048 (N_19048,N_16143,N_16748);
nand U19049 (N_19049,N_16648,N_16597);
nand U19050 (N_19050,N_16699,N_17844);
nor U19051 (N_19051,N_16255,N_16500);
or U19052 (N_19052,N_17796,N_16327);
nand U19053 (N_19053,N_17793,N_16592);
nor U19054 (N_19054,N_17091,N_16261);
xnor U19055 (N_19055,N_16772,N_17485);
nand U19056 (N_19056,N_16856,N_16535);
or U19057 (N_19057,N_17029,N_17794);
nand U19058 (N_19058,N_17490,N_17255);
or U19059 (N_19059,N_17725,N_16663);
nand U19060 (N_19060,N_17384,N_16268);
xnor U19061 (N_19061,N_17501,N_16722);
or U19062 (N_19062,N_17224,N_16437);
xnor U19063 (N_19063,N_17605,N_16653);
and U19064 (N_19064,N_17344,N_16640);
nor U19065 (N_19065,N_16685,N_17535);
nor U19066 (N_19066,N_17680,N_17611);
and U19067 (N_19067,N_16852,N_16252);
or U19068 (N_19068,N_17549,N_16473);
or U19069 (N_19069,N_16137,N_17180);
or U19070 (N_19070,N_16607,N_17965);
or U19071 (N_19071,N_17745,N_16475);
nor U19072 (N_19072,N_16724,N_17368);
nor U19073 (N_19073,N_17456,N_17679);
and U19074 (N_19074,N_16853,N_17043);
nand U19075 (N_19075,N_16294,N_16625);
nor U19076 (N_19076,N_16104,N_17150);
and U19077 (N_19077,N_16790,N_16578);
and U19078 (N_19078,N_16785,N_16469);
nor U19079 (N_19079,N_16655,N_16106);
or U19080 (N_19080,N_16376,N_16068);
or U19081 (N_19081,N_16636,N_17532);
and U19082 (N_19082,N_16140,N_17547);
nor U19083 (N_19083,N_16496,N_16377);
or U19084 (N_19084,N_17121,N_17827);
nand U19085 (N_19085,N_17408,N_16145);
nand U19086 (N_19086,N_17684,N_16582);
and U19087 (N_19087,N_17285,N_16643);
xnor U19088 (N_19088,N_16242,N_16048);
nand U19089 (N_19089,N_17485,N_16398);
or U19090 (N_19090,N_17305,N_17812);
nand U19091 (N_19091,N_16882,N_17700);
or U19092 (N_19092,N_17157,N_16487);
nor U19093 (N_19093,N_16763,N_17168);
nand U19094 (N_19094,N_17153,N_17459);
nor U19095 (N_19095,N_17133,N_17819);
nor U19096 (N_19096,N_17693,N_17688);
xor U19097 (N_19097,N_17895,N_16342);
xnor U19098 (N_19098,N_16651,N_16268);
nand U19099 (N_19099,N_17279,N_16055);
or U19100 (N_19100,N_16243,N_17093);
nor U19101 (N_19101,N_17097,N_17031);
and U19102 (N_19102,N_17746,N_17994);
xor U19103 (N_19103,N_17898,N_17208);
and U19104 (N_19104,N_16356,N_17442);
xor U19105 (N_19105,N_17545,N_16142);
or U19106 (N_19106,N_17962,N_16247);
and U19107 (N_19107,N_17866,N_17725);
nand U19108 (N_19108,N_17946,N_16859);
and U19109 (N_19109,N_16827,N_16681);
nand U19110 (N_19110,N_17416,N_17838);
xnor U19111 (N_19111,N_17802,N_16571);
xor U19112 (N_19112,N_16857,N_16513);
nand U19113 (N_19113,N_16025,N_16550);
and U19114 (N_19114,N_17497,N_17916);
nand U19115 (N_19115,N_17891,N_17999);
and U19116 (N_19116,N_17389,N_17031);
or U19117 (N_19117,N_17702,N_17529);
and U19118 (N_19118,N_17139,N_17391);
xor U19119 (N_19119,N_17369,N_17408);
nand U19120 (N_19120,N_17087,N_17708);
nor U19121 (N_19121,N_16764,N_16869);
or U19122 (N_19122,N_16415,N_16669);
and U19123 (N_19123,N_17518,N_16490);
and U19124 (N_19124,N_16503,N_16846);
xnor U19125 (N_19125,N_17465,N_17724);
xor U19126 (N_19126,N_17483,N_16559);
and U19127 (N_19127,N_17660,N_16086);
nor U19128 (N_19128,N_17096,N_16952);
nor U19129 (N_19129,N_16446,N_17900);
nand U19130 (N_19130,N_16324,N_16297);
nor U19131 (N_19131,N_17881,N_16839);
nand U19132 (N_19132,N_17015,N_17987);
nand U19133 (N_19133,N_16534,N_17563);
nand U19134 (N_19134,N_17702,N_16512);
or U19135 (N_19135,N_16818,N_17795);
or U19136 (N_19136,N_16902,N_17211);
xnor U19137 (N_19137,N_17457,N_16239);
or U19138 (N_19138,N_16463,N_17809);
nand U19139 (N_19139,N_17703,N_16805);
nand U19140 (N_19140,N_17225,N_17791);
and U19141 (N_19141,N_17932,N_16332);
nor U19142 (N_19142,N_17492,N_16584);
and U19143 (N_19143,N_17657,N_16352);
and U19144 (N_19144,N_17459,N_17554);
nor U19145 (N_19145,N_17892,N_16358);
nor U19146 (N_19146,N_16208,N_17883);
and U19147 (N_19147,N_17559,N_17937);
nor U19148 (N_19148,N_17629,N_16256);
xor U19149 (N_19149,N_16623,N_17701);
nand U19150 (N_19150,N_16359,N_17837);
or U19151 (N_19151,N_16610,N_17426);
and U19152 (N_19152,N_17701,N_17330);
nand U19153 (N_19153,N_16759,N_17633);
nor U19154 (N_19154,N_17509,N_17155);
nor U19155 (N_19155,N_16436,N_17971);
xnor U19156 (N_19156,N_17230,N_17106);
nand U19157 (N_19157,N_17420,N_17706);
nor U19158 (N_19158,N_16762,N_16770);
nor U19159 (N_19159,N_17739,N_17867);
nand U19160 (N_19160,N_17699,N_17479);
nand U19161 (N_19161,N_17182,N_16803);
nor U19162 (N_19162,N_16737,N_17809);
nand U19163 (N_19163,N_16581,N_16992);
or U19164 (N_19164,N_17076,N_17818);
xnor U19165 (N_19165,N_16311,N_17414);
xnor U19166 (N_19166,N_16527,N_17474);
xor U19167 (N_19167,N_17699,N_17588);
and U19168 (N_19168,N_16628,N_17746);
nand U19169 (N_19169,N_16367,N_16923);
or U19170 (N_19170,N_17264,N_16400);
nor U19171 (N_19171,N_17248,N_16915);
or U19172 (N_19172,N_16125,N_16208);
or U19173 (N_19173,N_17669,N_17434);
xnor U19174 (N_19174,N_17301,N_16996);
nand U19175 (N_19175,N_16970,N_16748);
nand U19176 (N_19176,N_17312,N_17053);
nand U19177 (N_19177,N_17567,N_16264);
or U19178 (N_19178,N_16367,N_17642);
and U19179 (N_19179,N_17488,N_16912);
nand U19180 (N_19180,N_16672,N_17461);
and U19181 (N_19181,N_17449,N_16498);
xor U19182 (N_19182,N_17229,N_17392);
and U19183 (N_19183,N_17791,N_16326);
nand U19184 (N_19184,N_17324,N_17247);
nor U19185 (N_19185,N_16251,N_16376);
or U19186 (N_19186,N_16184,N_16516);
and U19187 (N_19187,N_16520,N_16925);
xnor U19188 (N_19188,N_16561,N_16043);
or U19189 (N_19189,N_16146,N_17135);
or U19190 (N_19190,N_16580,N_16453);
xor U19191 (N_19191,N_17056,N_17228);
xnor U19192 (N_19192,N_17960,N_17885);
or U19193 (N_19193,N_17449,N_16494);
or U19194 (N_19194,N_17804,N_17896);
or U19195 (N_19195,N_16056,N_16571);
xor U19196 (N_19196,N_17730,N_17851);
xnor U19197 (N_19197,N_17838,N_16865);
nor U19198 (N_19198,N_16014,N_17963);
nand U19199 (N_19199,N_16934,N_16787);
nor U19200 (N_19200,N_17129,N_16423);
or U19201 (N_19201,N_17346,N_17088);
xor U19202 (N_19202,N_16031,N_17573);
nor U19203 (N_19203,N_17071,N_17156);
and U19204 (N_19204,N_16695,N_17123);
nand U19205 (N_19205,N_16805,N_17517);
nand U19206 (N_19206,N_17877,N_16008);
or U19207 (N_19207,N_17613,N_16847);
xor U19208 (N_19208,N_16437,N_16165);
nor U19209 (N_19209,N_16768,N_17855);
nor U19210 (N_19210,N_17635,N_17880);
nor U19211 (N_19211,N_16539,N_16201);
nor U19212 (N_19212,N_17521,N_17528);
nand U19213 (N_19213,N_17727,N_17211);
or U19214 (N_19214,N_17617,N_16648);
xor U19215 (N_19215,N_17683,N_16651);
and U19216 (N_19216,N_17146,N_16656);
nor U19217 (N_19217,N_17531,N_16411);
and U19218 (N_19218,N_16297,N_17141);
nor U19219 (N_19219,N_17169,N_17392);
nand U19220 (N_19220,N_17803,N_17508);
nand U19221 (N_19221,N_16318,N_17785);
nor U19222 (N_19222,N_16318,N_17675);
or U19223 (N_19223,N_17540,N_16443);
nand U19224 (N_19224,N_17111,N_17013);
and U19225 (N_19225,N_17425,N_16268);
and U19226 (N_19226,N_17246,N_17576);
and U19227 (N_19227,N_17863,N_16441);
xnor U19228 (N_19228,N_17709,N_16400);
xnor U19229 (N_19229,N_17418,N_16137);
and U19230 (N_19230,N_16318,N_17591);
nand U19231 (N_19231,N_17314,N_16454);
or U19232 (N_19232,N_17610,N_17828);
and U19233 (N_19233,N_16351,N_17657);
or U19234 (N_19234,N_17929,N_17993);
xor U19235 (N_19235,N_16393,N_17732);
nand U19236 (N_19236,N_16004,N_17196);
or U19237 (N_19237,N_16016,N_16136);
xor U19238 (N_19238,N_17586,N_16361);
xnor U19239 (N_19239,N_17273,N_17208);
and U19240 (N_19240,N_16910,N_17842);
and U19241 (N_19241,N_17528,N_17518);
nand U19242 (N_19242,N_16932,N_16513);
or U19243 (N_19243,N_17418,N_16365);
nand U19244 (N_19244,N_17996,N_17226);
xnor U19245 (N_19245,N_16809,N_17356);
and U19246 (N_19246,N_16765,N_16119);
or U19247 (N_19247,N_17576,N_17288);
and U19248 (N_19248,N_17469,N_17622);
and U19249 (N_19249,N_17294,N_16162);
and U19250 (N_19250,N_17634,N_16490);
nor U19251 (N_19251,N_17193,N_16315);
nand U19252 (N_19252,N_16268,N_17717);
xnor U19253 (N_19253,N_17332,N_17754);
xnor U19254 (N_19254,N_17275,N_17510);
nor U19255 (N_19255,N_16818,N_16405);
nand U19256 (N_19256,N_17182,N_17984);
or U19257 (N_19257,N_17500,N_16900);
and U19258 (N_19258,N_17698,N_17430);
nor U19259 (N_19259,N_17663,N_16196);
nor U19260 (N_19260,N_16997,N_16782);
or U19261 (N_19261,N_16664,N_17626);
nand U19262 (N_19262,N_17749,N_16954);
or U19263 (N_19263,N_16888,N_17540);
or U19264 (N_19264,N_17049,N_17547);
nand U19265 (N_19265,N_17393,N_17474);
or U19266 (N_19266,N_17537,N_16497);
and U19267 (N_19267,N_17722,N_16166);
and U19268 (N_19268,N_16641,N_17763);
or U19269 (N_19269,N_16724,N_16387);
xor U19270 (N_19270,N_17050,N_16056);
or U19271 (N_19271,N_16315,N_17404);
or U19272 (N_19272,N_17735,N_16551);
or U19273 (N_19273,N_16579,N_16743);
nor U19274 (N_19274,N_16616,N_16035);
xnor U19275 (N_19275,N_16609,N_16911);
nor U19276 (N_19276,N_17460,N_16371);
or U19277 (N_19277,N_16010,N_16421);
nor U19278 (N_19278,N_16952,N_16371);
nor U19279 (N_19279,N_16697,N_16850);
nand U19280 (N_19280,N_16731,N_16952);
xor U19281 (N_19281,N_17373,N_17269);
nor U19282 (N_19282,N_16922,N_17854);
nand U19283 (N_19283,N_17234,N_16475);
xor U19284 (N_19284,N_17157,N_16898);
nor U19285 (N_19285,N_16739,N_17622);
or U19286 (N_19286,N_17311,N_16782);
nor U19287 (N_19287,N_17227,N_16429);
nand U19288 (N_19288,N_17225,N_17946);
xnor U19289 (N_19289,N_17077,N_17206);
and U19290 (N_19290,N_17790,N_16574);
and U19291 (N_19291,N_16550,N_16640);
and U19292 (N_19292,N_16168,N_16753);
nor U19293 (N_19293,N_17441,N_16510);
and U19294 (N_19294,N_17575,N_16864);
nand U19295 (N_19295,N_17728,N_17925);
or U19296 (N_19296,N_16267,N_16934);
nand U19297 (N_19297,N_17273,N_16285);
xnor U19298 (N_19298,N_17916,N_17152);
and U19299 (N_19299,N_17169,N_16210);
nor U19300 (N_19300,N_17865,N_17408);
nand U19301 (N_19301,N_17558,N_16081);
and U19302 (N_19302,N_17105,N_16692);
or U19303 (N_19303,N_17529,N_16812);
xnor U19304 (N_19304,N_16056,N_16208);
or U19305 (N_19305,N_16519,N_17076);
nor U19306 (N_19306,N_17311,N_16270);
nor U19307 (N_19307,N_17967,N_16353);
nor U19308 (N_19308,N_16592,N_17972);
or U19309 (N_19309,N_16685,N_16025);
or U19310 (N_19310,N_17046,N_17509);
xnor U19311 (N_19311,N_17503,N_16683);
and U19312 (N_19312,N_16118,N_17518);
and U19313 (N_19313,N_16850,N_16038);
nand U19314 (N_19314,N_17741,N_17903);
xnor U19315 (N_19315,N_17035,N_16805);
xor U19316 (N_19316,N_17706,N_17797);
or U19317 (N_19317,N_17826,N_17056);
xnor U19318 (N_19318,N_16932,N_16788);
xnor U19319 (N_19319,N_17064,N_16585);
nor U19320 (N_19320,N_16392,N_16099);
or U19321 (N_19321,N_16289,N_16147);
nand U19322 (N_19322,N_16499,N_16476);
nor U19323 (N_19323,N_16536,N_16999);
and U19324 (N_19324,N_17663,N_16655);
xor U19325 (N_19325,N_17504,N_16222);
xnor U19326 (N_19326,N_16421,N_17204);
nor U19327 (N_19327,N_16747,N_16251);
nor U19328 (N_19328,N_16243,N_17364);
or U19329 (N_19329,N_17251,N_17810);
or U19330 (N_19330,N_16915,N_17573);
xnor U19331 (N_19331,N_17888,N_17167);
or U19332 (N_19332,N_16893,N_17569);
nand U19333 (N_19333,N_16158,N_17433);
nand U19334 (N_19334,N_17984,N_16067);
or U19335 (N_19335,N_17848,N_17518);
and U19336 (N_19336,N_17225,N_16533);
nor U19337 (N_19337,N_17015,N_17061);
xor U19338 (N_19338,N_17656,N_16712);
and U19339 (N_19339,N_17092,N_17571);
nand U19340 (N_19340,N_16622,N_16540);
xnor U19341 (N_19341,N_16391,N_17012);
and U19342 (N_19342,N_16558,N_16119);
or U19343 (N_19343,N_17421,N_16880);
and U19344 (N_19344,N_17244,N_16919);
or U19345 (N_19345,N_16801,N_17484);
xor U19346 (N_19346,N_17124,N_16673);
nand U19347 (N_19347,N_17476,N_17467);
nor U19348 (N_19348,N_16996,N_16313);
and U19349 (N_19349,N_17591,N_17127);
and U19350 (N_19350,N_17422,N_17518);
and U19351 (N_19351,N_17987,N_17234);
nor U19352 (N_19352,N_17830,N_16878);
nor U19353 (N_19353,N_17916,N_17605);
nand U19354 (N_19354,N_16225,N_16687);
xnor U19355 (N_19355,N_17895,N_17605);
or U19356 (N_19356,N_16422,N_17401);
and U19357 (N_19357,N_17186,N_17544);
nand U19358 (N_19358,N_16131,N_17580);
or U19359 (N_19359,N_17567,N_16644);
and U19360 (N_19360,N_17264,N_17963);
nor U19361 (N_19361,N_16074,N_17887);
or U19362 (N_19362,N_17648,N_16418);
and U19363 (N_19363,N_17944,N_17332);
nor U19364 (N_19364,N_16942,N_17863);
xnor U19365 (N_19365,N_16550,N_16022);
and U19366 (N_19366,N_17948,N_17734);
nand U19367 (N_19367,N_17722,N_16989);
nor U19368 (N_19368,N_17467,N_16879);
xnor U19369 (N_19369,N_17832,N_16877);
nor U19370 (N_19370,N_16684,N_16732);
xor U19371 (N_19371,N_16423,N_16635);
or U19372 (N_19372,N_16420,N_17819);
nand U19373 (N_19373,N_16793,N_16640);
xor U19374 (N_19374,N_16883,N_16742);
nand U19375 (N_19375,N_16829,N_16796);
nor U19376 (N_19376,N_17706,N_17578);
nor U19377 (N_19377,N_17795,N_16965);
nand U19378 (N_19378,N_17410,N_17061);
xnor U19379 (N_19379,N_17610,N_16974);
xnor U19380 (N_19380,N_16725,N_16649);
xnor U19381 (N_19381,N_17570,N_17736);
xor U19382 (N_19382,N_16915,N_17721);
nand U19383 (N_19383,N_16488,N_16736);
xnor U19384 (N_19384,N_16245,N_17580);
or U19385 (N_19385,N_16695,N_17057);
nand U19386 (N_19386,N_17853,N_17986);
xnor U19387 (N_19387,N_16822,N_16214);
or U19388 (N_19388,N_16104,N_16578);
xor U19389 (N_19389,N_17945,N_17007);
xnor U19390 (N_19390,N_17683,N_17868);
xnor U19391 (N_19391,N_17745,N_17230);
xor U19392 (N_19392,N_17311,N_17019);
xor U19393 (N_19393,N_16269,N_16047);
and U19394 (N_19394,N_16578,N_16175);
and U19395 (N_19395,N_16784,N_17191);
or U19396 (N_19396,N_17757,N_16103);
xor U19397 (N_19397,N_17005,N_16328);
nand U19398 (N_19398,N_17097,N_17801);
nor U19399 (N_19399,N_16315,N_17335);
nand U19400 (N_19400,N_16917,N_17028);
or U19401 (N_19401,N_17186,N_16772);
or U19402 (N_19402,N_17912,N_16626);
or U19403 (N_19403,N_17337,N_16743);
and U19404 (N_19404,N_17990,N_17124);
nor U19405 (N_19405,N_16798,N_16069);
xnor U19406 (N_19406,N_17433,N_16447);
or U19407 (N_19407,N_17082,N_16890);
nor U19408 (N_19408,N_17045,N_17297);
nand U19409 (N_19409,N_17556,N_16970);
nor U19410 (N_19410,N_17245,N_16758);
nand U19411 (N_19411,N_16527,N_16424);
nor U19412 (N_19412,N_16738,N_17541);
nor U19413 (N_19413,N_17330,N_16718);
and U19414 (N_19414,N_17945,N_16836);
nor U19415 (N_19415,N_17337,N_16787);
and U19416 (N_19416,N_17589,N_16211);
xnor U19417 (N_19417,N_17748,N_17480);
nand U19418 (N_19418,N_16753,N_16127);
or U19419 (N_19419,N_17731,N_16865);
xnor U19420 (N_19420,N_16446,N_17726);
nor U19421 (N_19421,N_16708,N_16610);
nor U19422 (N_19422,N_16902,N_17943);
nand U19423 (N_19423,N_16139,N_16947);
xor U19424 (N_19424,N_16387,N_16397);
xor U19425 (N_19425,N_17348,N_17420);
and U19426 (N_19426,N_16800,N_17492);
xnor U19427 (N_19427,N_16737,N_16010);
or U19428 (N_19428,N_16315,N_17956);
and U19429 (N_19429,N_16169,N_17037);
nor U19430 (N_19430,N_16941,N_16837);
or U19431 (N_19431,N_16323,N_16228);
nand U19432 (N_19432,N_16678,N_17079);
and U19433 (N_19433,N_16568,N_17726);
nor U19434 (N_19434,N_17851,N_16572);
xnor U19435 (N_19435,N_16791,N_17280);
xor U19436 (N_19436,N_16423,N_16503);
and U19437 (N_19437,N_16498,N_17473);
and U19438 (N_19438,N_16878,N_16921);
and U19439 (N_19439,N_16257,N_16799);
xor U19440 (N_19440,N_17105,N_17438);
and U19441 (N_19441,N_17676,N_17886);
xnor U19442 (N_19442,N_16553,N_16645);
nor U19443 (N_19443,N_17600,N_17558);
nand U19444 (N_19444,N_17373,N_16735);
xnor U19445 (N_19445,N_17230,N_16784);
xor U19446 (N_19446,N_16689,N_16117);
nand U19447 (N_19447,N_17145,N_17746);
nand U19448 (N_19448,N_16016,N_17375);
nor U19449 (N_19449,N_17920,N_16842);
and U19450 (N_19450,N_16517,N_16205);
nand U19451 (N_19451,N_16544,N_17890);
nor U19452 (N_19452,N_16054,N_17669);
and U19453 (N_19453,N_17805,N_16797);
or U19454 (N_19454,N_17674,N_16128);
nand U19455 (N_19455,N_16744,N_17907);
or U19456 (N_19456,N_16849,N_16334);
or U19457 (N_19457,N_17187,N_16079);
and U19458 (N_19458,N_16970,N_17620);
and U19459 (N_19459,N_16987,N_17091);
and U19460 (N_19460,N_17666,N_16539);
and U19461 (N_19461,N_17915,N_17124);
nand U19462 (N_19462,N_16339,N_16067);
or U19463 (N_19463,N_16042,N_17245);
and U19464 (N_19464,N_16658,N_16577);
nand U19465 (N_19465,N_17728,N_17748);
nand U19466 (N_19466,N_17053,N_17088);
and U19467 (N_19467,N_17791,N_17262);
nand U19468 (N_19468,N_17638,N_16930);
or U19469 (N_19469,N_16981,N_17994);
nor U19470 (N_19470,N_16523,N_16097);
nand U19471 (N_19471,N_16615,N_17914);
and U19472 (N_19472,N_16783,N_16022);
nor U19473 (N_19473,N_17215,N_16933);
and U19474 (N_19474,N_16133,N_16551);
and U19475 (N_19475,N_17310,N_17907);
xor U19476 (N_19476,N_17838,N_17576);
nand U19477 (N_19477,N_16847,N_17906);
or U19478 (N_19478,N_16116,N_17114);
xor U19479 (N_19479,N_17978,N_16273);
nand U19480 (N_19480,N_17738,N_16256);
or U19481 (N_19481,N_17104,N_16959);
and U19482 (N_19482,N_17204,N_16627);
xor U19483 (N_19483,N_16143,N_17444);
nand U19484 (N_19484,N_17275,N_17732);
nand U19485 (N_19485,N_16255,N_17224);
nand U19486 (N_19486,N_17542,N_16646);
and U19487 (N_19487,N_16419,N_16501);
or U19488 (N_19488,N_16283,N_17007);
xnor U19489 (N_19489,N_16494,N_16615);
or U19490 (N_19490,N_17562,N_16666);
xor U19491 (N_19491,N_17733,N_16086);
nand U19492 (N_19492,N_17193,N_17691);
xnor U19493 (N_19493,N_17757,N_17544);
or U19494 (N_19494,N_16762,N_16174);
xnor U19495 (N_19495,N_16324,N_17892);
nand U19496 (N_19496,N_16156,N_17834);
nor U19497 (N_19497,N_16800,N_17576);
xnor U19498 (N_19498,N_16689,N_16241);
nand U19499 (N_19499,N_16685,N_16862);
xor U19500 (N_19500,N_17615,N_17623);
nor U19501 (N_19501,N_17492,N_17017);
or U19502 (N_19502,N_17785,N_16795);
nor U19503 (N_19503,N_17311,N_16319);
nand U19504 (N_19504,N_17400,N_16553);
nor U19505 (N_19505,N_16730,N_17628);
nor U19506 (N_19506,N_17774,N_17605);
or U19507 (N_19507,N_16237,N_17510);
and U19508 (N_19508,N_16579,N_16684);
nor U19509 (N_19509,N_16666,N_17488);
nor U19510 (N_19510,N_16048,N_16042);
and U19511 (N_19511,N_17460,N_16954);
and U19512 (N_19512,N_17604,N_17134);
xnor U19513 (N_19513,N_16215,N_16076);
nor U19514 (N_19514,N_16997,N_16630);
or U19515 (N_19515,N_17818,N_16193);
nand U19516 (N_19516,N_17314,N_17056);
or U19517 (N_19517,N_16133,N_16201);
or U19518 (N_19518,N_16888,N_17770);
xor U19519 (N_19519,N_17680,N_17713);
xnor U19520 (N_19520,N_17786,N_16798);
xnor U19521 (N_19521,N_17117,N_17707);
or U19522 (N_19522,N_17287,N_16268);
and U19523 (N_19523,N_16346,N_16219);
nand U19524 (N_19524,N_16612,N_17153);
or U19525 (N_19525,N_17516,N_17529);
xnor U19526 (N_19526,N_17440,N_17870);
and U19527 (N_19527,N_17794,N_16831);
xnor U19528 (N_19528,N_16902,N_16175);
or U19529 (N_19529,N_17626,N_17481);
or U19530 (N_19530,N_16019,N_17471);
nor U19531 (N_19531,N_17901,N_16620);
xor U19532 (N_19532,N_17205,N_17321);
xnor U19533 (N_19533,N_16032,N_16473);
or U19534 (N_19534,N_16883,N_17861);
nand U19535 (N_19535,N_16785,N_17376);
xor U19536 (N_19536,N_16497,N_16932);
or U19537 (N_19537,N_16835,N_16186);
and U19538 (N_19538,N_16994,N_16900);
or U19539 (N_19539,N_16693,N_17335);
and U19540 (N_19540,N_16599,N_17631);
nand U19541 (N_19541,N_17135,N_17070);
and U19542 (N_19542,N_16916,N_16282);
nor U19543 (N_19543,N_16179,N_16895);
or U19544 (N_19544,N_17208,N_16125);
nor U19545 (N_19545,N_16884,N_17472);
nor U19546 (N_19546,N_16833,N_16988);
nand U19547 (N_19547,N_17408,N_16963);
nand U19548 (N_19548,N_16614,N_16559);
nand U19549 (N_19549,N_17534,N_16698);
or U19550 (N_19550,N_16526,N_17075);
nand U19551 (N_19551,N_17374,N_16907);
nand U19552 (N_19552,N_17469,N_17870);
xnor U19553 (N_19553,N_17892,N_17816);
or U19554 (N_19554,N_17277,N_16478);
and U19555 (N_19555,N_17899,N_17181);
and U19556 (N_19556,N_17094,N_16117);
and U19557 (N_19557,N_16579,N_16966);
nor U19558 (N_19558,N_17099,N_16796);
and U19559 (N_19559,N_16932,N_16174);
and U19560 (N_19560,N_16738,N_17294);
or U19561 (N_19561,N_17123,N_16084);
nand U19562 (N_19562,N_16512,N_16996);
nor U19563 (N_19563,N_17942,N_16825);
or U19564 (N_19564,N_16745,N_16601);
and U19565 (N_19565,N_16761,N_16050);
nand U19566 (N_19566,N_16856,N_17273);
and U19567 (N_19567,N_17253,N_16241);
or U19568 (N_19568,N_17010,N_16703);
nor U19569 (N_19569,N_17064,N_16349);
nor U19570 (N_19570,N_16164,N_16293);
or U19571 (N_19571,N_16586,N_17040);
xor U19572 (N_19572,N_16789,N_17687);
xor U19573 (N_19573,N_16007,N_17148);
and U19574 (N_19574,N_17508,N_17778);
nand U19575 (N_19575,N_17892,N_17289);
and U19576 (N_19576,N_17518,N_17059);
nor U19577 (N_19577,N_17040,N_17196);
or U19578 (N_19578,N_17621,N_16790);
xor U19579 (N_19579,N_17996,N_17252);
nor U19580 (N_19580,N_17933,N_17622);
nor U19581 (N_19581,N_16005,N_16436);
nand U19582 (N_19582,N_17470,N_17094);
nor U19583 (N_19583,N_17295,N_16387);
xnor U19584 (N_19584,N_16529,N_17728);
or U19585 (N_19585,N_17267,N_16301);
xor U19586 (N_19586,N_17293,N_16412);
nand U19587 (N_19587,N_16178,N_17060);
nand U19588 (N_19588,N_16720,N_17502);
nor U19589 (N_19589,N_17979,N_16315);
nand U19590 (N_19590,N_17977,N_17396);
and U19591 (N_19591,N_17355,N_16738);
and U19592 (N_19592,N_16632,N_16866);
nor U19593 (N_19593,N_16310,N_17580);
and U19594 (N_19594,N_16590,N_17008);
and U19595 (N_19595,N_17496,N_16359);
nand U19596 (N_19596,N_16902,N_17670);
xor U19597 (N_19597,N_16799,N_16452);
nor U19598 (N_19598,N_16527,N_16782);
nor U19599 (N_19599,N_16307,N_16367);
and U19600 (N_19600,N_16330,N_16037);
nor U19601 (N_19601,N_16941,N_17022);
nor U19602 (N_19602,N_17296,N_16994);
or U19603 (N_19603,N_17210,N_17246);
nor U19604 (N_19604,N_17121,N_16826);
nor U19605 (N_19605,N_17822,N_16695);
nand U19606 (N_19606,N_17614,N_16421);
or U19607 (N_19607,N_17027,N_16564);
nand U19608 (N_19608,N_17221,N_17475);
xor U19609 (N_19609,N_17901,N_17234);
nand U19610 (N_19610,N_17192,N_17342);
xnor U19611 (N_19611,N_17717,N_16075);
nor U19612 (N_19612,N_16086,N_16816);
nor U19613 (N_19613,N_16047,N_16465);
nor U19614 (N_19614,N_17324,N_17846);
and U19615 (N_19615,N_17045,N_17602);
nor U19616 (N_19616,N_17684,N_17821);
nor U19617 (N_19617,N_16448,N_16591);
nor U19618 (N_19618,N_16949,N_16261);
or U19619 (N_19619,N_16718,N_16699);
or U19620 (N_19620,N_16179,N_16153);
and U19621 (N_19621,N_16304,N_17785);
nand U19622 (N_19622,N_17216,N_17953);
and U19623 (N_19623,N_16074,N_16735);
xor U19624 (N_19624,N_17537,N_16103);
or U19625 (N_19625,N_16491,N_16571);
or U19626 (N_19626,N_17293,N_16989);
nor U19627 (N_19627,N_16915,N_16089);
nor U19628 (N_19628,N_16169,N_16167);
and U19629 (N_19629,N_17676,N_16144);
nor U19630 (N_19630,N_17142,N_17791);
nor U19631 (N_19631,N_17627,N_17648);
nor U19632 (N_19632,N_16512,N_17279);
xor U19633 (N_19633,N_16976,N_16090);
and U19634 (N_19634,N_16821,N_16211);
and U19635 (N_19635,N_17746,N_16482);
nand U19636 (N_19636,N_16965,N_17331);
or U19637 (N_19637,N_16297,N_16557);
and U19638 (N_19638,N_16348,N_17968);
and U19639 (N_19639,N_16099,N_16095);
nor U19640 (N_19640,N_17012,N_16642);
and U19641 (N_19641,N_17114,N_16269);
or U19642 (N_19642,N_16208,N_17232);
and U19643 (N_19643,N_17734,N_17285);
nand U19644 (N_19644,N_17412,N_16628);
nand U19645 (N_19645,N_16367,N_16882);
nand U19646 (N_19646,N_17019,N_16145);
xnor U19647 (N_19647,N_17186,N_17516);
xor U19648 (N_19648,N_16693,N_16326);
nand U19649 (N_19649,N_17080,N_16520);
xor U19650 (N_19650,N_16612,N_16663);
nor U19651 (N_19651,N_16833,N_16432);
xnor U19652 (N_19652,N_16432,N_17140);
and U19653 (N_19653,N_17250,N_16448);
or U19654 (N_19654,N_16960,N_16225);
nor U19655 (N_19655,N_17847,N_17002);
xor U19656 (N_19656,N_17152,N_17809);
xor U19657 (N_19657,N_16549,N_16615);
or U19658 (N_19658,N_17500,N_17142);
nand U19659 (N_19659,N_16673,N_17572);
nor U19660 (N_19660,N_17085,N_16351);
nor U19661 (N_19661,N_17202,N_16603);
and U19662 (N_19662,N_17469,N_16587);
nor U19663 (N_19663,N_17656,N_17384);
or U19664 (N_19664,N_17646,N_16560);
nor U19665 (N_19665,N_16235,N_17147);
nor U19666 (N_19666,N_16247,N_17619);
nor U19667 (N_19667,N_17593,N_16498);
nor U19668 (N_19668,N_17119,N_16638);
nor U19669 (N_19669,N_17329,N_16365);
or U19670 (N_19670,N_17465,N_16736);
and U19671 (N_19671,N_16586,N_16785);
and U19672 (N_19672,N_16013,N_16841);
nor U19673 (N_19673,N_17852,N_17575);
xnor U19674 (N_19674,N_17029,N_17693);
or U19675 (N_19675,N_16808,N_17364);
xor U19676 (N_19676,N_17097,N_16117);
nand U19677 (N_19677,N_16388,N_16455);
or U19678 (N_19678,N_16570,N_16919);
nor U19679 (N_19679,N_16424,N_16664);
nand U19680 (N_19680,N_16836,N_17813);
nor U19681 (N_19681,N_17827,N_17733);
and U19682 (N_19682,N_16209,N_16463);
nand U19683 (N_19683,N_17163,N_16486);
or U19684 (N_19684,N_16055,N_16113);
nand U19685 (N_19685,N_17522,N_16669);
and U19686 (N_19686,N_17230,N_16419);
or U19687 (N_19687,N_16280,N_16192);
nor U19688 (N_19688,N_17369,N_16373);
nor U19689 (N_19689,N_16965,N_16907);
or U19690 (N_19690,N_16353,N_17201);
or U19691 (N_19691,N_16714,N_17772);
nand U19692 (N_19692,N_17039,N_16570);
nor U19693 (N_19693,N_17797,N_17258);
nand U19694 (N_19694,N_16731,N_16997);
nand U19695 (N_19695,N_16029,N_17631);
xnor U19696 (N_19696,N_16519,N_17985);
xor U19697 (N_19697,N_16774,N_16927);
nor U19698 (N_19698,N_17973,N_17145);
xor U19699 (N_19699,N_16184,N_16888);
nand U19700 (N_19700,N_16599,N_17597);
xnor U19701 (N_19701,N_16675,N_16765);
nand U19702 (N_19702,N_16860,N_17773);
nor U19703 (N_19703,N_17148,N_17621);
xnor U19704 (N_19704,N_16141,N_17527);
and U19705 (N_19705,N_17749,N_16028);
nor U19706 (N_19706,N_16451,N_16435);
xor U19707 (N_19707,N_16452,N_17377);
or U19708 (N_19708,N_16579,N_17090);
and U19709 (N_19709,N_16005,N_17300);
nand U19710 (N_19710,N_17253,N_17642);
nand U19711 (N_19711,N_17949,N_17559);
nand U19712 (N_19712,N_16969,N_17061);
nor U19713 (N_19713,N_17430,N_16305);
and U19714 (N_19714,N_17091,N_17037);
and U19715 (N_19715,N_17512,N_17790);
nor U19716 (N_19716,N_16737,N_16607);
nand U19717 (N_19717,N_16998,N_17679);
and U19718 (N_19718,N_17531,N_16213);
nor U19719 (N_19719,N_16344,N_16398);
xor U19720 (N_19720,N_16640,N_16183);
or U19721 (N_19721,N_16703,N_17970);
nand U19722 (N_19722,N_17854,N_17663);
or U19723 (N_19723,N_16938,N_17755);
nor U19724 (N_19724,N_17212,N_16535);
xor U19725 (N_19725,N_16366,N_17676);
or U19726 (N_19726,N_16322,N_17999);
nor U19727 (N_19727,N_16094,N_16452);
xnor U19728 (N_19728,N_17425,N_17107);
nand U19729 (N_19729,N_17063,N_17373);
xnor U19730 (N_19730,N_17616,N_17225);
xnor U19731 (N_19731,N_17306,N_17915);
and U19732 (N_19732,N_16849,N_17862);
nor U19733 (N_19733,N_16814,N_17357);
or U19734 (N_19734,N_17551,N_17139);
nor U19735 (N_19735,N_16749,N_16640);
nor U19736 (N_19736,N_16828,N_16855);
nand U19737 (N_19737,N_16586,N_16635);
xnor U19738 (N_19738,N_16796,N_16507);
nand U19739 (N_19739,N_16194,N_16556);
and U19740 (N_19740,N_16951,N_16685);
xor U19741 (N_19741,N_16654,N_16291);
and U19742 (N_19742,N_17391,N_17528);
nor U19743 (N_19743,N_16115,N_17441);
nor U19744 (N_19744,N_17033,N_17105);
xnor U19745 (N_19745,N_17103,N_17372);
xnor U19746 (N_19746,N_17830,N_17513);
nand U19747 (N_19747,N_16725,N_17503);
and U19748 (N_19748,N_17951,N_16215);
nand U19749 (N_19749,N_16483,N_16013);
xor U19750 (N_19750,N_17362,N_16217);
nand U19751 (N_19751,N_17867,N_16432);
nor U19752 (N_19752,N_17566,N_16830);
nor U19753 (N_19753,N_16756,N_17846);
xnor U19754 (N_19754,N_16044,N_16346);
nor U19755 (N_19755,N_16095,N_16100);
or U19756 (N_19756,N_16156,N_16784);
or U19757 (N_19757,N_16916,N_16021);
or U19758 (N_19758,N_17303,N_16541);
xor U19759 (N_19759,N_17424,N_17081);
xnor U19760 (N_19760,N_17547,N_17121);
xnor U19761 (N_19761,N_16724,N_16346);
nand U19762 (N_19762,N_16621,N_17599);
xnor U19763 (N_19763,N_16494,N_16239);
nor U19764 (N_19764,N_17674,N_16896);
or U19765 (N_19765,N_16538,N_16341);
nor U19766 (N_19766,N_16743,N_16815);
nor U19767 (N_19767,N_17149,N_17522);
xnor U19768 (N_19768,N_16239,N_16759);
and U19769 (N_19769,N_16675,N_17313);
nor U19770 (N_19770,N_16000,N_16959);
and U19771 (N_19771,N_16559,N_17787);
nand U19772 (N_19772,N_16770,N_17832);
nor U19773 (N_19773,N_16758,N_17933);
nor U19774 (N_19774,N_17136,N_17052);
and U19775 (N_19775,N_17640,N_17624);
xnor U19776 (N_19776,N_16561,N_17965);
nand U19777 (N_19777,N_17507,N_16155);
nand U19778 (N_19778,N_16081,N_17154);
xnor U19779 (N_19779,N_16318,N_17151);
xnor U19780 (N_19780,N_17197,N_17458);
or U19781 (N_19781,N_16952,N_17787);
nor U19782 (N_19782,N_17135,N_16124);
nand U19783 (N_19783,N_17742,N_17727);
xnor U19784 (N_19784,N_17684,N_16836);
and U19785 (N_19785,N_17354,N_16191);
nor U19786 (N_19786,N_17082,N_17875);
xnor U19787 (N_19787,N_17110,N_17458);
nor U19788 (N_19788,N_16869,N_16046);
and U19789 (N_19789,N_17411,N_16295);
and U19790 (N_19790,N_16638,N_16349);
nand U19791 (N_19791,N_17040,N_17785);
or U19792 (N_19792,N_16572,N_17960);
or U19793 (N_19793,N_16228,N_17097);
nor U19794 (N_19794,N_16039,N_16398);
nand U19795 (N_19795,N_17716,N_16080);
xor U19796 (N_19796,N_17228,N_17877);
nor U19797 (N_19797,N_16284,N_17948);
xor U19798 (N_19798,N_17877,N_17762);
and U19799 (N_19799,N_17333,N_16711);
nor U19800 (N_19800,N_16226,N_17554);
or U19801 (N_19801,N_16870,N_17616);
or U19802 (N_19802,N_17378,N_16003);
nand U19803 (N_19803,N_17631,N_16601);
nor U19804 (N_19804,N_17054,N_17811);
xor U19805 (N_19805,N_16517,N_16603);
or U19806 (N_19806,N_17837,N_17159);
and U19807 (N_19807,N_16740,N_16040);
nand U19808 (N_19808,N_17233,N_16115);
nor U19809 (N_19809,N_16206,N_16554);
or U19810 (N_19810,N_16436,N_17061);
nand U19811 (N_19811,N_16737,N_17930);
and U19812 (N_19812,N_17484,N_17531);
and U19813 (N_19813,N_16139,N_17745);
nor U19814 (N_19814,N_16659,N_16777);
or U19815 (N_19815,N_17616,N_16487);
nor U19816 (N_19816,N_17372,N_16874);
xnor U19817 (N_19817,N_16594,N_16054);
nand U19818 (N_19818,N_16668,N_17833);
and U19819 (N_19819,N_16207,N_17543);
or U19820 (N_19820,N_16868,N_17624);
nor U19821 (N_19821,N_16864,N_17446);
nand U19822 (N_19822,N_17860,N_17390);
and U19823 (N_19823,N_17022,N_17209);
xor U19824 (N_19824,N_17990,N_16765);
nand U19825 (N_19825,N_16693,N_16509);
and U19826 (N_19826,N_17059,N_17994);
or U19827 (N_19827,N_16695,N_16631);
xor U19828 (N_19828,N_17970,N_16918);
and U19829 (N_19829,N_16541,N_16555);
or U19830 (N_19830,N_16117,N_17399);
nor U19831 (N_19831,N_17587,N_16152);
nand U19832 (N_19832,N_16616,N_17812);
or U19833 (N_19833,N_16423,N_16114);
nor U19834 (N_19834,N_16675,N_17409);
and U19835 (N_19835,N_17594,N_16644);
or U19836 (N_19836,N_16809,N_17431);
xor U19837 (N_19837,N_17676,N_16840);
and U19838 (N_19838,N_17510,N_16960);
xnor U19839 (N_19839,N_17428,N_17400);
or U19840 (N_19840,N_17338,N_17036);
nor U19841 (N_19841,N_16292,N_17848);
nand U19842 (N_19842,N_16546,N_17745);
and U19843 (N_19843,N_17346,N_17928);
xor U19844 (N_19844,N_16063,N_17186);
or U19845 (N_19845,N_16553,N_16954);
nor U19846 (N_19846,N_16125,N_16583);
nand U19847 (N_19847,N_17381,N_16975);
nand U19848 (N_19848,N_17504,N_17791);
xnor U19849 (N_19849,N_16787,N_17281);
nor U19850 (N_19850,N_17453,N_17295);
and U19851 (N_19851,N_16600,N_16863);
and U19852 (N_19852,N_17428,N_17569);
and U19853 (N_19853,N_17282,N_16206);
nor U19854 (N_19854,N_16601,N_16643);
and U19855 (N_19855,N_16212,N_17843);
nor U19856 (N_19856,N_16988,N_17627);
and U19857 (N_19857,N_16315,N_16809);
and U19858 (N_19858,N_17862,N_17484);
xnor U19859 (N_19859,N_16710,N_16481);
nor U19860 (N_19860,N_17787,N_17070);
and U19861 (N_19861,N_17242,N_17517);
nor U19862 (N_19862,N_16221,N_17633);
nor U19863 (N_19863,N_16822,N_17666);
and U19864 (N_19864,N_16332,N_17886);
nand U19865 (N_19865,N_17727,N_17509);
nand U19866 (N_19866,N_17703,N_16177);
nand U19867 (N_19867,N_17503,N_17773);
or U19868 (N_19868,N_16575,N_17007);
and U19869 (N_19869,N_16891,N_16963);
nor U19870 (N_19870,N_16310,N_16171);
or U19871 (N_19871,N_16035,N_16462);
and U19872 (N_19872,N_16080,N_17277);
nor U19873 (N_19873,N_16329,N_16057);
nor U19874 (N_19874,N_17226,N_17684);
nor U19875 (N_19875,N_17747,N_17039);
nand U19876 (N_19876,N_16482,N_17967);
nor U19877 (N_19877,N_16954,N_17675);
xor U19878 (N_19878,N_16473,N_17904);
nand U19879 (N_19879,N_16226,N_16905);
xnor U19880 (N_19880,N_16091,N_16000);
xnor U19881 (N_19881,N_17961,N_17906);
xor U19882 (N_19882,N_17069,N_17822);
and U19883 (N_19883,N_16457,N_17576);
xor U19884 (N_19884,N_17672,N_16631);
nand U19885 (N_19885,N_17036,N_16529);
or U19886 (N_19886,N_17117,N_17069);
and U19887 (N_19887,N_16041,N_16636);
and U19888 (N_19888,N_17281,N_16192);
nand U19889 (N_19889,N_16404,N_17278);
and U19890 (N_19890,N_17554,N_17305);
xnor U19891 (N_19891,N_16223,N_16575);
nor U19892 (N_19892,N_16171,N_17814);
nand U19893 (N_19893,N_17787,N_17158);
nor U19894 (N_19894,N_17839,N_16978);
nand U19895 (N_19895,N_17570,N_16840);
and U19896 (N_19896,N_16608,N_16985);
nand U19897 (N_19897,N_16156,N_16437);
nor U19898 (N_19898,N_17421,N_16318);
xor U19899 (N_19899,N_16499,N_17895);
and U19900 (N_19900,N_17894,N_16027);
nor U19901 (N_19901,N_17432,N_16853);
nor U19902 (N_19902,N_17936,N_16218);
nor U19903 (N_19903,N_17389,N_17499);
nand U19904 (N_19904,N_17989,N_16675);
xnor U19905 (N_19905,N_16833,N_16064);
nor U19906 (N_19906,N_17330,N_17076);
xnor U19907 (N_19907,N_16396,N_16914);
or U19908 (N_19908,N_17489,N_16592);
and U19909 (N_19909,N_16872,N_16713);
and U19910 (N_19910,N_17961,N_17942);
nand U19911 (N_19911,N_16102,N_16031);
nand U19912 (N_19912,N_16914,N_17912);
or U19913 (N_19913,N_16745,N_16277);
nor U19914 (N_19914,N_17867,N_17630);
nor U19915 (N_19915,N_17654,N_17817);
xnor U19916 (N_19916,N_17685,N_17558);
nand U19917 (N_19917,N_16902,N_17145);
or U19918 (N_19918,N_16609,N_16710);
nor U19919 (N_19919,N_17459,N_17152);
or U19920 (N_19920,N_16565,N_16244);
and U19921 (N_19921,N_16714,N_16104);
nand U19922 (N_19922,N_17590,N_16798);
nor U19923 (N_19923,N_17459,N_16777);
and U19924 (N_19924,N_16047,N_17699);
xor U19925 (N_19925,N_16305,N_17331);
nand U19926 (N_19926,N_16097,N_17866);
nor U19927 (N_19927,N_16902,N_16486);
nand U19928 (N_19928,N_17299,N_16462);
nand U19929 (N_19929,N_17893,N_16194);
and U19930 (N_19930,N_17408,N_16878);
nand U19931 (N_19931,N_17706,N_16412);
xor U19932 (N_19932,N_16635,N_16110);
nor U19933 (N_19933,N_16498,N_16572);
xor U19934 (N_19934,N_16469,N_16963);
nor U19935 (N_19935,N_16563,N_16488);
xnor U19936 (N_19936,N_17824,N_16690);
or U19937 (N_19937,N_16717,N_16532);
xor U19938 (N_19938,N_16187,N_17103);
nor U19939 (N_19939,N_16232,N_16217);
nand U19940 (N_19940,N_16804,N_16188);
or U19941 (N_19941,N_16737,N_17710);
or U19942 (N_19942,N_17815,N_17348);
and U19943 (N_19943,N_17045,N_17076);
and U19944 (N_19944,N_17645,N_17785);
nand U19945 (N_19945,N_17406,N_17596);
and U19946 (N_19946,N_17179,N_17950);
nor U19947 (N_19947,N_16625,N_17942);
and U19948 (N_19948,N_17346,N_16456);
and U19949 (N_19949,N_16370,N_16010);
nand U19950 (N_19950,N_17055,N_17940);
and U19951 (N_19951,N_17946,N_16638);
or U19952 (N_19952,N_17021,N_16737);
and U19953 (N_19953,N_17423,N_16324);
xor U19954 (N_19954,N_17088,N_17280);
or U19955 (N_19955,N_16020,N_17641);
xor U19956 (N_19956,N_17716,N_17987);
nor U19957 (N_19957,N_16924,N_17090);
or U19958 (N_19958,N_17569,N_16184);
nand U19959 (N_19959,N_17737,N_16925);
and U19960 (N_19960,N_17893,N_17339);
nand U19961 (N_19961,N_17706,N_17052);
nand U19962 (N_19962,N_17153,N_16037);
xor U19963 (N_19963,N_16521,N_17245);
xor U19964 (N_19964,N_16296,N_17065);
nand U19965 (N_19965,N_16833,N_16422);
nand U19966 (N_19966,N_17400,N_17144);
or U19967 (N_19967,N_17370,N_16331);
nand U19968 (N_19968,N_17472,N_17663);
nor U19969 (N_19969,N_16121,N_17600);
nor U19970 (N_19970,N_16602,N_16352);
nor U19971 (N_19971,N_16826,N_16319);
and U19972 (N_19972,N_17366,N_17559);
and U19973 (N_19973,N_17331,N_17636);
nand U19974 (N_19974,N_17775,N_16334);
nand U19975 (N_19975,N_16530,N_16762);
or U19976 (N_19976,N_16818,N_17637);
or U19977 (N_19977,N_17710,N_17766);
xor U19978 (N_19978,N_17012,N_16011);
and U19979 (N_19979,N_17324,N_16940);
or U19980 (N_19980,N_17449,N_17789);
nand U19981 (N_19981,N_17352,N_17518);
or U19982 (N_19982,N_16630,N_17919);
and U19983 (N_19983,N_16930,N_17878);
nand U19984 (N_19984,N_16844,N_16387);
and U19985 (N_19985,N_16115,N_17299);
nand U19986 (N_19986,N_16460,N_16501);
or U19987 (N_19987,N_16046,N_17946);
xor U19988 (N_19988,N_17062,N_16747);
nand U19989 (N_19989,N_17646,N_17977);
nor U19990 (N_19990,N_16708,N_16623);
and U19991 (N_19991,N_16252,N_16102);
nand U19992 (N_19992,N_17791,N_17336);
and U19993 (N_19993,N_17277,N_17892);
or U19994 (N_19994,N_17291,N_16597);
and U19995 (N_19995,N_17160,N_16802);
nand U19996 (N_19996,N_16075,N_17941);
and U19997 (N_19997,N_17700,N_17724);
xnor U19998 (N_19998,N_17673,N_16171);
nor U19999 (N_19999,N_17077,N_17407);
and U20000 (N_20000,N_19191,N_19330);
or U20001 (N_20001,N_18182,N_19393);
or U20002 (N_20002,N_18514,N_19140);
or U20003 (N_20003,N_18490,N_19049);
nand U20004 (N_20004,N_19283,N_18866);
nand U20005 (N_20005,N_19300,N_18336);
and U20006 (N_20006,N_19204,N_18334);
and U20007 (N_20007,N_19489,N_19856);
nor U20008 (N_20008,N_19170,N_18066);
and U20009 (N_20009,N_19534,N_19697);
xnor U20010 (N_20010,N_19171,N_19174);
xor U20011 (N_20011,N_19553,N_18238);
xnor U20012 (N_20012,N_18725,N_19360);
nor U20013 (N_20013,N_19863,N_18338);
and U20014 (N_20014,N_19507,N_18147);
or U20015 (N_20015,N_19168,N_18222);
xor U20016 (N_20016,N_18511,N_18790);
or U20017 (N_20017,N_19898,N_18635);
nand U20018 (N_20018,N_18747,N_18224);
nand U20019 (N_20019,N_19816,N_18285);
nor U20020 (N_20020,N_18632,N_18452);
or U20021 (N_20021,N_19595,N_19304);
or U20022 (N_20022,N_18375,N_19135);
and U20023 (N_20023,N_19799,N_19707);
and U20024 (N_20024,N_19095,N_18071);
nor U20025 (N_20025,N_19109,N_19787);
nor U20026 (N_20026,N_18557,N_19552);
nand U20027 (N_20027,N_19518,N_18534);
nor U20028 (N_20028,N_18077,N_19568);
nor U20029 (N_20029,N_19163,N_19169);
or U20030 (N_20030,N_18296,N_18259);
or U20031 (N_20031,N_18035,N_18096);
nor U20032 (N_20032,N_19546,N_18012);
and U20033 (N_20033,N_19399,N_18703);
or U20034 (N_20034,N_18158,N_18543);
and U20035 (N_20035,N_19466,N_19993);
nor U20036 (N_20036,N_19597,N_18544);
nand U20037 (N_20037,N_18308,N_19090);
xnor U20038 (N_20038,N_19992,N_19366);
and U20039 (N_20039,N_18652,N_19797);
nor U20040 (N_20040,N_18559,N_19849);
or U20041 (N_20041,N_18713,N_18762);
xor U20042 (N_20042,N_19016,N_18636);
or U20043 (N_20043,N_18440,N_19275);
nand U20044 (N_20044,N_19352,N_18433);
nor U20045 (N_20045,N_19130,N_18893);
and U20046 (N_20046,N_18168,N_19529);
nand U20047 (N_20047,N_18914,N_19886);
nor U20048 (N_20048,N_18954,N_19487);
nor U20049 (N_20049,N_19019,N_18247);
nand U20050 (N_20050,N_19225,N_18665);
nor U20051 (N_20051,N_19535,N_19616);
nor U20052 (N_20052,N_18860,N_19820);
and U20053 (N_20053,N_19607,N_18844);
nand U20054 (N_20054,N_18122,N_19394);
or U20055 (N_20055,N_18955,N_19005);
or U20056 (N_20056,N_18664,N_19955);
nand U20057 (N_20057,N_19277,N_19326);
nor U20058 (N_20058,N_18272,N_18851);
nand U20059 (N_20059,N_18102,N_18822);
or U20060 (N_20060,N_18563,N_18082);
or U20061 (N_20061,N_18803,N_19630);
xor U20062 (N_20062,N_18701,N_19721);
nor U20063 (N_20063,N_18568,N_18030);
or U20064 (N_20064,N_18633,N_19289);
xor U20065 (N_20065,N_18760,N_19162);
nor U20066 (N_20066,N_19857,N_18005);
xor U20067 (N_20067,N_19754,N_19122);
or U20068 (N_20068,N_18835,N_18289);
nor U20069 (N_20069,N_18029,N_19753);
xnor U20070 (N_20070,N_19691,N_19236);
xor U20071 (N_20071,N_19295,N_19824);
or U20072 (N_20072,N_18867,N_18039);
xnor U20073 (N_20073,N_19773,N_18898);
xor U20074 (N_20074,N_18146,N_18373);
nand U20075 (N_20075,N_18998,N_19108);
or U20076 (N_20076,N_18832,N_19664);
and U20077 (N_20077,N_18442,N_19063);
nor U20078 (N_20078,N_19615,N_18078);
xnor U20079 (N_20079,N_19195,N_18004);
nor U20080 (N_20080,N_18143,N_18922);
xnor U20081 (N_20081,N_18989,N_19506);
or U20082 (N_20082,N_19087,N_18817);
and U20083 (N_20083,N_19240,N_19980);
nand U20084 (N_20084,N_18582,N_19491);
xnor U20085 (N_20085,N_19934,N_19390);
and U20086 (N_20086,N_18706,N_18971);
xnor U20087 (N_20087,N_19207,N_18885);
nor U20088 (N_20088,N_19759,N_19335);
and U20089 (N_20089,N_19059,N_19986);
nand U20090 (N_20090,N_18927,N_19965);
or U20091 (N_20091,N_18092,N_19316);
nand U20092 (N_20092,N_19792,N_18780);
and U20093 (N_20093,N_19337,N_18074);
or U20094 (N_20094,N_18681,N_18435);
nand U20095 (N_20095,N_19788,N_18230);
nand U20096 (N_20096,N_18977,N_18492);
nor U20097 (N_20097,N_18166,N_19806);
or U20098 (N_20098,N_19011,N_19643);
xnor U20099 (N_20099,N_19895,N_19502);
nor U20100 (N_20100,N_18424,N_19091);
nand U20101 (N_20101,N_18972,N_18983);
xor U20102 (N_20102,N_19488,N_18729);
nor U20103 (N_20103,N_18060,N_19678);
or U20104 (N_20104,N_18990,N_18397);
nand U20105 (N_20105,N_18763,N_19235);
xor U20106 (N_20106,N_18402,N_18600);
nor U20107 (N_20107,N_18572,N_18391);
nor U20108 (N_20108,N_18930,N_18431);
xor U20109 (N_20109,N_19966,N_19409);
nand U20110 (N_20110,N_19132,N_18831);
and U20111 (N_20111,N_18303,N_19948);
and U20112 (N_20112,N_18597,N_18819);
or U20113 (N_20113,N_19186,N_18718);
or U20114 (N_20114,N_18390,N_19967);
xnor U20115 (N_20115,N_19351,N_18133);
xnor U20116 (N_20116,N_19810,N_19877);
nor U20117 (N_20117,N_18484,N_18687);
nand U20118 (N_20118,N_19447,N_18352);
nor U20119 (N_20119,N_19575,N_19157);
nand U20120 (N_20120,N_18364,N_19252);
nor U20121 (N_20121,N_18468,N_18073);
nand U20122 (N_20122,N_18907,N_19148);
xor U20123 (N_20123,N_19545,N_19264);
nor U20124 (N_20124,N_18612,N_18340);
xor U20125 (N_20125,N_18804,N_19740);
or U20126 (N_20126,N_18466,N_18294);
nor U20127 (N_20127,N_19724,N_19377);
nand U20128 (N_20128,N_18761,N_19920);
xnor U20129 (N_20129,N_18674,N_19818);
and U20130 (N_20130,N_18770,N_19407);
nand U20131 (N_20131,N_18061,N_18801);
and U20132 (N_20132,N_18996,N_19854);
and U20133 (N_20133,N_18883,N_19349);
nand U20134 (N_20134,N_19048,N_19017);
xnor U20135 (N_20135,N_18510,N_19670);
or U20136 (N_20136,N_18614,N_18946);
xnor U20137 (N_20137,N_18538,N_18891);
xnor U20138 (N_20138,N_19836,N_18644);
xor U20139 (N_20139,N_18174,N_18639);
xor U20140 (N_20140,N_18889,N_18536);
or U20141 (N_20141,N_19514,N_18067);
nand U20142 (N_20142,N_19183,N_18054);
nand U20143 (N_20143,N_19242,N_19246);
and U20144 (N_20144,N_18877,N_19528);
or U20145 (N_20145,N_18624,N_19778);
or U20146 (N_20146,N_19975,N_19257);
nand U20147 (N_20147,N_19729,N_19714);
and U20148 (N_20148,N_19805,N_18669);
nor U20149 (N_20149,N_19984,N_18052);
nor U20150 (N_20150,N_19782,N_18697);
or U20151 (N_20151,N_19583,N_18820);
or U20152 (N_20152,N_19560,N_19100);
nor U20153 (N_20153,N_18087,N_19141);
nor U20154 (N_20154,N_18556,N_19471);
nor U20155 (N_20155,N_19710,N_18611);
xnor U20156 (N_20156,N_19635,N_18615);
and U20157 (N_20157,N_18566,N_19228);
xnor U20158 (N_20158,N_18290,N_19777);
or U20159 (N_20159,N_19290,N_19718);
xor U20160 (N_20160,N_19562,N_18522);
or U20161 (N_20161,N_18252,N_18156);
and U20162 (N_20162,N_19230,N_19780);
nor U20163 (N_20163,N_19403,N_18164);
nand U20164 (N_20164,N_18455,N_19903);
xnor U20165 (N_20165,N_18117,N_19524);
nor U20166 (N_20166,N_18311,N_19313);
or U20167 (N_20167,N_18199,N_19702);
nor U20168 (N_20168,N_18666,N_18362);
nor U20169 (N_20169,N_18281,N_18553);
and U20170 (N_20170,N_19896,N_18127);
nand U20171 (N_20171,N_18917,N_18273);
or U20172 (N_20172,N_19189,N_19279);
xnor U20173 (N_20173,N_19159,N_18836);
xor U20174 (N_20174,N_18549,N_19860);
and U20175 (N_20175,N_19268,N_18830);
and U20176 (N_20176,N_18346,N_19259);
nor U20177 (N_20177,N_19943,N_18858);
nand U20178 (N_20178,N_19770,N_18190);
xor U20179 (N_20179,N_18018,N_18302);
nand U20180 (N_20180,N_18261,N_18848);
or U20181 (N_20181,N_18354,N_19968);
xor U20182 (N_20182,N_19266,N_19124);
or U20183 (N_20183,N_19716,N_18620);
xnor U20184 (N_20184,N_18111,N_18266);
or U20185 (N_20185,N_18098,N_18523);
xor U20186 (N_20186,N_18943,N_18220);
nand U20187 (N_20187,N_18084,N_19558);
or U20188 (N_20188,N_19699,N_18382);
or U20189 (N_20189,N_19004,N_18807);
and U20190 (N_20190,N_18815,N_19591);
xor U20191 (N_20191,N_18876,N_18861);
or U20192 (N_20192,N_19609,N_18828);
and U20193 (N_20193,N_18276,N_19062);
nand U20194 (N_20194,N_18240,N_19176);
nor U20195 (N_20195,N_18886,N_19241);
xor U20196 (N_20196,N_19387,N_18865);
nand U20197 (N_20197,N_19334,N_19873);
nand U20198 (N_20198,N_19646,N_19097);
nor U20199 (N_20199,N_19610,N_19054);
nand U20200 (N_20200,N_19869,N_18331);
nand U20201 (N_20201,N_18297,N_19404);
nand U20202 (N_20202,N_18902,N_19400);
xnor U20203 (N_20203,N_19160,N_18504);
or U20204 (N_20204,N_18888,N_18229);
nor U20205 (N_20205,N_18890,N_18715);
or U20206 (N_20206,N_18135,N_18080);
nor U20207 (N_20207,N_18618,N_19258);
and U20208 (N_20208,N_18043,N_18376);
xnor U20209 (N_20209,N_18862,N_19478);
or U20210 (N_20210,N_18319,N_18952);
nand U20211 (N_20211,N_18965,N_19315);
nand U20212 (N_20212,N_19009,N_18217);
or U20213 (N_20213,N_19479,N_19434);
nor U20214 (N_20214,N_18313,N_18027);
xor U20215 (N_20215,N_18816,N_18975);
xor U20216 (N_20216,N_18179,N_18593);
or U20217 (N_20217,N_19842,N_18467);
or U20218 (N_20218,N_19789,N_19752);
and U20219 (N_20219,N_18347,N_18598);
xor U20220 (N_20220,N_19309,N_18200);
and U20221 (N_20221,N_19324,N_18839);
nand U20222 (N_20222,N_19733,N_18274);
xnor U20223 (N_20223,N_18337,N_19775);
nand U20224 (N_20224,N_19861,N_19631);
nor U20225 (N_20225,N_18516,N_19379);
and U20226 (N_20226,N_19372,N_19867);
xnor U20227 (N_20227,N_18163,N_19288);
nor U20228 (N_20228,N_19310,N_18743);
and U20229 (N_20229,N_18314,N_19604);
or U20230 (N_20230,N_18567,N_18962);
xnor U20231 (N_20231,N_19276,N_19526);
nor U20232 (N_20232,N_19500,N_18932);
and U20233 (N_20233,N_18683,N_18947);
or U20234 (N_20234,N_19515,N_18833);
and U20235 (N_20235,N_18970,N_18020);
and U20236 (N_20236,N_18837,N_19203);
nor U20237 (N_20237,N_19651,N_18976);
and U20238 (N_20238,N_18642,N_19738);
nor U20239 (N_20239,N_18404,N_19131);
and U20240 (N_20240,N_19929,N_18180);
xor U20241 (N_20241,N_19462,N_18233);
or U20242 (N_20242,N_19231,N_19041);
xor U20243 (N_20243,N_18900,N_19667);
xor U20244 (N_20244,N_18416,N_19022);
nand U20245 (N_20245,N_18806,N_19779);
nor U20246 (N_20246,N_18728,N_18245);
nand U20247 (N_20247,N_18695,N_19850);
nor U20248 (N_20248,N_18478,N_19215);
nand U20249 (N_20249,N_19501,N_19505);
or U20250 (N_20250,N_18894,N_19858);
or U20251 (N_20251,N_18570,N_18388);
and U20252 (N_20252,N_19255,N_18509);
xnor U20253 (N_20253,N_18505,N_19701);
nand U20254 (N_20254,N_19812,N_18063);
xnor U20255 (N_20255,N_18854,N_18776);
nand U20256 (N_20256,N_18257,N_18076);
nor U20257 (N_20257,N_19641,N_19089);
nor U20258 (N_20258,N_18793,N_18772);
nor U20259 (N_20259,N_19866,N_18961);
or U20260 (N_20260,N_19226,N_19119);
or U20261 (N_20261,N_19184,N_18269);
and U20262 (N_20262,N_19987,N_19638);
and U20263 (N_20263,N_19033,N_18749);
nor U20264 (N_20264,N_19765,N_19074);
or U20265 (N_20265,N_19563,N_18344);
and U20266 (N_20266,N_18110,N_19991);
and U20267 (N_20267,N_19293,N_18533);
xnor U20268 (N_20268,N_19477,N_19239);
nand U20269 (N_20269,N_18797,N_19767);
nand U20270 (N_20270,N_18560,N_18320);
nand U20271 (N_20271,N_18441,N_19549);
nand U20272 (N_20272,N_18381,N_19743);
or U20273 (N_20273,N_19603,N_18910);
xor U20274 (N_20274,N_18204,N_18722);
xnor U20275 (N_20275,N_18656,N_19154);
or U20276 (N_20276,N_19726,N_18342);
or U20277 (N_20277,N_19695,N_18757);
nand U20278 (N_20278,N_18141,N_19247);
or U20279 (N_20279,N_19414,N_19446);
nor U20280 (N_20280,N_18155,N_19431);
nand U20281 (N_20281,N_19668,N_19213);
or U20282 (N_20282,N_18449,N_19134);
xnor U20283 (N_20283,N_18472,N_19730);
nand U20284 (N_20284,N_19055,N_18583);
xnor U20285 (N_20285,N_18434,N_18169);
xor U20286 (N_20286,N_18811,N_18855);
nand U20287 (N_20287,N_18978,N_18950);
and U20288 (N_20288,N_19322,N_18649);
nor U20289 (N_20289,N_18814,N_18630);
nor U20290 (N_20290,N_19598,N_18032);
and U20291 (N_20291,N_18445,N_19893);
nor U20292 (N_20292,N_19318,N_19385);
xnor U20293 (N_20293,N_18775,N_19067);
and U20294 (N_20294,N_19273,N_19922);
nand U20295 (N_20295,N_19755,N_18643);
and U20296 (N_20296,N_19210,N_18070);
xor U20297 (N_20297,N_18069,N_19852);
nor U20298 (N_20298,N_19373,N_19143);
nand U20299 (N_20299,N_19574,N_18106);
or U20300 (N_20300,N_19803,N_19722);
nand U20301 (N_20301,N_18226,N_18904);
and U20302 (N_20302,N_18145,N_19959);
or U20303 (N_20303,N_19826,N_19227);
or U20304 (N_20304,N_19748,N_18335);
or U20305 (N_20305,N_19149,N_18916);
nand U20306 (N_20306,N_19569,N_18227);
nor U20307 (N_20307,N_19152,N_18678);
nor U20308 (N_20308,N_18209,N_18963);
xor U20309 (N_20309,N_18040,N_18037);
nand U20310 (N_20310,N_18878,N_18931);
nand U20311 (N_20311,N_18654,N_19881);
xor U20312 (N_20312,N_19249,N_18564);
or U20313 (N_20313,N_18154,N_18842);
or U20314 (N_20314,N_18979,N_18144);
or U20315 (N_20315,N_18909,N_18545);
xnor U20316 (N_20316,N_19694,N_19460);
and U20317 (N_20317,N_19296,N_19619);
xor U20318 (N_20318,N_18824,N_18000);
nor U20319 (N_20319,N_19899,N_19985);
or U20320 (N_20320,N_19870,N_19329);
and U20321 (N_20321,N_19926,N_18095);
or U20322 (N_20322,N_19072,N_18808);
xnor U20323 (N_20323,N_18960,N_18994);
nand U20324 (N_20324,N_18244,N_18400);
nand U20325 (N_20325,N_19713,N_18707);
nor U20326 (N_20326,N_18263,N_19650);
or U20327 (N_20327,N_18634,N_18873);
nand U20328 (N_20328,N_19673,N_18184);
xor U20329 (N_20329,N_19761,N_19188);
or U20330 (N_20330,N_18912,N_19923);
xor U20331 (N_20331,N_18350,N_18631);
xor U20332 (N_20332,N_18050,N_18906);
and U20333 (N_20333,N_18512,N_19177);
xnor U20334 (N_20334,N_18495,N_18363);
nor U20335 (N_20335,N_19199,N_19118);
nand U20336 (N_20336,N_19212,N_18231);
nand U20337 (N_20337,N_18462,N_18389);
nor U20338 (N_20338,N_18892,N_18126);
nor U20339 (N_20339,N_19843,N_18675);
xnor U20340 (N_20340,N_18726,N_19282);
nor U20341 (N_20341,N_18409,N_18689);
nor U20342 (N_20342,N_18958,N_19474);
and U20343 (N_20343,N_19064,N_19876);
or U20344 (N_20344,N_18679,N_18500);
or U20345 (N_20345,N_19617,N_18953);
nand U20346 (N_20346,N_18599,N_18370);
xnor U20347 (N_20347,N_18021,N_18491);
nand U20348 (N_20348,N_19470,N_18714);
or U20349 (N_20349,N_19859,N_18371);
or U20350 (N_20350,N_18766,N_19823);
or U20351 (N_20351,N_19564,N_19561);
or U20352 (N_20352,N_18268,N_19871);
nor U20353 (N_20353,N_19925,N_18913);
nor U20354 (N_20354,N_19439,N_19080);
or U20355 (N_20355,N_18939,N_19681);
xor U20356 (N_20356,N_18298,N_19178);
nand U20357 (N_20357,N_18361,N_18571);
or U20358 (N_20358,N_19175,N_19437);
nor U20359 (N_20359,N_19442,N_19164);
xor U20360 (N_20360,N_19565,N_18090);
nand U20361 (N_20361,N_19874,N_18015);
nand U20362 (N_20362,N_19051,N_18194);
nor U20363 (N_20363,N_19031,N_19034);
xnor U20364 (N_20364,N_19342,N_19126);
nor U20365 (N_20365,N_18368,N_18677);
nand U20366 (N_20366,N_19793,N_18595);
nor U20367 (N_20367,N_19301,N_18136);
nor U20368 (N_20368,N_18422,N_19682);
nand U20369 (N_20369,N_18993,N_19750);
and U20370 (N_20370,N_19653,N_19116);
or U20371 (N_20371,N_18781,N_19592);
nand U20372 (N_20372,N_19086,N_19205);
xor U20373 (N_20373,N_19909,N_18365);
or U20374 (N_20374,N_19092,N_18315);
nor U20375 (N_20375,N_19465,N_18104);
nand U20376 (N_20376,N_19760,N_18055);
nor U20377 (N_20377,N_18283,N_19737);
and U20378 (N_20378,N_19504,N_19815);
xnor U20379 (N_20379,N_19368,N_18938);
or U20380 (N_20380,N_19637,N_18869);
nor U20381 (N_20381,N_18602,N_18805);
nor U20382 (N_20382,N_19361,N_18506);
xnor U20383 (N_20383,N_19795,N_19953);
and U20384 (N_20384,N_18942,N_19093);
xnor U20385 (N_20385,N_19411,N_19305);
nor U20386 (N_20386,N_18609,N_19885);
nand U20387 (N_20387,N_18300,N_18195);
nor U20388 (N_20388,N_18755,N_18264);
and U20389 (N_20389,N_19219,N_18525);
nand U20390 (N_20390,N_18629,N_18554);
nand U20391 (N_20391,N_19359,N_19888);
xnor U20392 (N_20392,N_19901,N_19657);
and U20393 (N_20393,N_18202,N_19884);
nand U20394 (N_20394,N_18119,N_19261);
nand U20395 (N_20395,N_18608,N_19350);
and U20396 (N_20396,N_19516,N_18800);
and U20397 (N_20397,N_19634,N_19050);
nor U20398 (N_20398,N_18459,N_18278);
and U20399 (N_20399,N_19445,N_18019);
xor U20400 (N_20400,N_19040,N_19254);
and U20401 (N_20401,N_18871,N_18610);
nor U20402 (N_20402,N_18705,N_19998);
nor U20403 (N_20403,N_19686,N_18577);
or U20404 (N_20404,N_18765,N_19757);
nor U20405 (N_20405,N_19066,N_19596);
nor U20406 (N_20406,N_18648,N_19832);
nor U20407 (N_20407,N_19081,N_18053);
or U20408 (N_20408,N_18905,N_18437);
nor U20409 (N_20409,N_19454,N_19693);
and U20410 (N_20410,N_19455,N_18246);
nand U20411 (N_20411,N_19606,N_18210);
nand U20412 (N_20412,N_18162,N_18650);
xor U20413 (N_20413,N_19397,N_18358);
nor U20414 (N_20414,N_19408,N_19547);
nor U20415 (N_20415,N_19913,N_18540);
nor U20416 (N_20416,N_19994,N_18345);
and U20417 (N_20417,N_18688,N_19572);
nand U20418 (N_20418,N_19539,N_18109);
and U20419 (N_20419,N_19232,N_18575);
nand U20420 (N_20420,N_19223,N_19660);
or U20421 (N_20421,N_19928,N_19015);
or U20422 (N_20422,N_18089,N_18480);
and U20423 (N_20423,N_18139,N_18286);
nor U20424 (N_20424,N_18051,N_18251);
and U20425 (N_20425,N_19807,N_19023);
nand U20426 (N_20426,N_18895,N_18647);
xor U20427 (N_20427,N_18881,N_18925);
xnor U20428 (N_20428,N_18017,N_19811);
nand U20429 (N_20429,N_18426,N_18232);
and U20430 (N_20430,N_18756,N_18698);
and U20431 (N_20431,N_19035,N_19425);
and U20432 (N_20432,N_18573,N_19949);
xnor U20433 (N_20433,N_19763,N_19971);
or U20434 (N_20434,N_19639,N_19421);
xnor U20435 (N_20435,N_18105,N_18011);
xnor U20436 (N_20436,N_19785,N_18619);
xor U20437 (N_20437,N_19665,N_19344);
nand U20438 (N_20438,N_18456,N_18640);
or U20439 (N_20439,N_18542,N_19648);
and U20440 (N_20440,N_19263,N_19626);
nor U20441 (N_20441,N_18115,N_19083);
and U20442 (N_20442,N_19530,N_19099);
nor U20443 (N_20443,N_19957,N_18348);
nand U20444 (N_20444,N_18548,N_18079);
or U20445 (N_20445,N_18696,N_18524);
nand U20446 (N_20446,N_18987,N_18395);
nor U20447 (N_20447,N_19999,N_19892);
xor U20448 (N_20448,N_19735,N_19703);
or U20449 (N_20449,N_18530,N_18153);
and U20450 (N_20450,N_19527,N_18493);
nor U20451 (N_20451,N_18288,N_19057);
nor U20452 (N_20452,N_18585,N_19593);
xnor U20453 (N_20453,N_19520,N_19156);
xnor U20454 (N_20454,N_19768,N_19769);
or U20455 (N_20455,N_18686,N_19731);
or U20456 (N_20456,N_18262,N_19997);
xor U20457 (N_20457,N_18929,N_19416);
nand U20458 (N_20458,N_18517,N_19060);
nand U20459 (N_20459,N_18584,N_19822);
nor U20460 (N_20460,N_18001,N_18008);
nor U20461 (N_20461,N_19904,N_19623);
or U20462 (N_20462,N_18737,N_18586);
or U20463 (N_20463,N_19555,N_19840);
xor U20464 (N_20464,N_18857,N_18736);
xor U20465 (N_20465,N_18042,N_18207);
nand U20466 (N_20466,N_19221,N_19036);
nand U20467 (N_20467,N_18408,N_18684);
xor U20468 (N_20468,N_19580,N_18081);
xor U20469 (N_20469,N_18420,N_19137);
and U20470 (N_20470,N_19587,N_19981);
nand U20471 (N_20471,N_18377,N_19484);
and U20472 (N_20472,N_19312,N_18520);
nand U20473 (N_20473,N_18065,N_19386);
xor U20474 (N_20474,N_18185,N_19392);
nor U20475 (N_20475,N_19389,N_19030);
and U20476 (N_20476,N_18138,N_18667);
nor U20477 (N_20477,N_19883,N_19941);
nor U20478 (N_20478,N_19192,N_18915);
or U20479 (N_20479,N_19675,N_19197);
nand U20480 (N_20480,N_18058,N_19383);
and U20481 (N_20481,N_18752,N_19503);
or U20482 (N_20482,N_18708,N_18537);
and U20483 (N_20483,N_19078,N_19307);
nor U20484 (N_20484,N_19222,N_19417);
nand U20485 (N_20485,N_19911,N_18821);
or U20486 (N_20486,N_18576,N_19625);
nand U20487 (N_20487,N_18956,N_19864);
nor U20488 (N_20488,N_19094,N_19636);
xor U20489 (N_20489,N_18280,N_19155);
or U20490 (N_20490,N_19936,N_18009);
nor U20491 (N_20491,N_19391,N_18007);
nor U20492 (N_20492,N_18321,N_19586);
nor U20493 (N_20493,N_19085,N_18845);
nor U20494 (N_20494,N_19308,N_18360);
and U20495 (N_20495,N_18118,N_19581);
xor U20496 (N_20496,N_19910,N_18341);
or U20497 (N_20497,N_19728,N_19771);
nor U20498 (N_20498,N_19029,N_19962);
nand U20499 (N_20499,N_18739,N_19677);
nand U20500 (N_20500,N_19989,N_18253);
nand U20501 (N_20501,N_18601,N_18613);
nor U20502 (N_20502,N_19136,N_19996);
or U20503 (N_20503,N_18405,N_18868);
or U20504 (N_20504,N_18234,N_19828);
and U20505 (N_20505,N_19432,N_19193);
nand U20506 (N_20506,N_19946,N_19600);
and U20507 (N_20507,N_19358,N_19972);
xnor U20508 (N_20508,N_19894,N_19747);
and U20509 (N_20509,N_19374,N_19933);
xnor U20510 (N_20510,N_19053,N_19882);
and U20511 (N_20511,N_18489,N_19878);
nor U20512 (N_20512,N_18398,N_19448);
or U20513 (N_20513,N_19357,N_18394);
nor U20514 (N_20514,N_19459,N_18161);
nor U20515 (N_20515,N_18176,N_19521);
or U20516 (N_20516,N_18148,N_18849);
xnor U20517 (N_20517,N_18870,N_19237);
and U20518 (N_20518,N_18062,N_19690);
nand U20519 (N_20519,N_18788,N_18719);
or U20520 (N_20520,N_19332,N_18329);
xnor U20521 (N_20521,N_18167,N_18799);
and U20522 (N_20522,N_19655,N_18519);
nor U20523 (N_20523,N_19298,N_19540);
or U20524 (N_20524,N_19935,N_19272);
or U20525 (N_20525,N_18592,N_18187);
nand U20526 (N_20526,N_18068,N_19674);
nand U20527 (N_20527,N_18014,N_18094);
and U20528 (N_20528,N_18211,N_18702);
or U20529 (N_20529,N_18937,N_19234);
nand U20530 (N_20530,N_19662,N_19644);
xor U20531 (N_20531,N_18275,N_18059);
xor U20532 (N_20532,N_19327,N_19443);
nor U20533 (N_20533,N_19271,N_18853);
and U20534 (N_20534,N_18237,N_18279);
and U20535 (N_20535,N_19902,N_19937);
nand U20536 (N_20536,N_19127,N_19746);
nor U20537 (N_20537,N_19113,N_18792);
xor U20538 (N_20538,N_18228,N_18150);
and U20539 (N_20539,N_18206,N_19021);
nand U20540 (N_20540,N_19918,N_18951);
xor U20541 (N_20541,N_19744,N_19341);
xor U20542 (N_20542,N_18933,N_19908);
and U20543 (N_20543,N_19954,N_18189);
xor U20544 (N_20544,N_19105,N_18108);
nor U20545 (N_20545,N_18123,N_19513);
or U20546 (N_20546,N_19709,N_18175);
xnor U20547 (N_20547,N_18731,N_18847);
nand U20548 (N_20548,N_19382,N_18604);
xnor U20549 (N_20549,N_18306,N_19492);
xor U20550 (N_20550,N_18935,N_19618);
or U20551 (N_20551,N_19570,N_18541);
and U20552 (N_20552,N_19613,N_18235);
and U20553 (N_20553,N_19656,N_18551);
xor U20554 (N_20554,N_18287,N_19839);
and U20555 (N_20555,N_18924,N_19827);
and U20556 (N_20556,N_18617,N_19096);
or U20557 (N_20557,N_18565,N_18093);
nand U20558 (N_20558,N_19444,N_19912);
and U20559 (N_20559,N_18333,N_19704);
and U20560 (N_20560,N_19940,N_18527);
nand U20561 (N_20561,N_18432,N_19245);
nand U20562 (N_20562,N_18165,N_18291);
xor U20563 (N_20563,N_19819,N_18097);
xor U20564 (N_20564,N_19068,N_18988);
or U20565 (N_20565,N_18457,N_18864);
nand U20566 (N_20566,N_18966,N_18590);
nor U20567 (N_20567,N_19075,N_19756);
nand U20568 (N_20568,N_18160,N_18901);
nand U20569 (N_20569,N_18796,N_18121);
and U20570 (N_20570,N_19875,N_18552);
or U20571 (N_20571,N_18680,N_19916);
and U20572 (N_20572,N_19745,N_19451);
or U20573 (N_20573,N_18508,N_18124);
nand U20574 (N_20574,N_19410,N_18465);
nand U20575 (N_20575,N_19123,N_19798);
xor U20576 (N_20576,N_19983,N_19576);
or U20577 (N_20577,N_18213,N_18267);
nand U20578 (N_20578,N_18771,N_19976);
xor U20579 (N_20579,N_19297,N_19429);
or U20580 (N_20580,N_18374,N_19608);
xor U20581 (N_20581,N_19951,N_18596);
nand U20582 (N_20582,N_18496,N_18170);
nand U20583 (N_20583,N_18526,N_19381);
nand U20584 (N_20584,N_19577,N_18392);
xor U20585 (N_20585,N_19880,N_18399);
and U20586 (N_20586,N_19463,N_19428);
nand U20587 (N_20587,N_18789,N_19796);
nand U20588 (N_20588,N_18277,N_19889);
or U20589 (N_20589,N_18421,N_19692);
and U20590 (N_20590,N_19129,N_19848);
and U20591 (N_20591,N_18239,N_19251);
or U20592 (N_20592,N_18622,N_18606);
or U20593 (N_20593,N_19736,N_18513);
and U20594 (N_20594,N_18383,N_18260);
xor U20595 (N_20595,N_19027,N_19319);
nor U20596 (N_20596,N_18787,N_18658);
nand U20597 (N_20597,N_19458,N_18721);
xnor U20598 (N_20598,N_19958,N_18940);
xnor U20599 (N_20599,N_18203,N_18129);
nor U20600 (N_20600,N_19579,N_19734);
nand U20601 (N_20601,N_19138,N_18471);
nor U20602 (N_20602,N_19669,N_18411);
and U20603 (N_20603,N_19794,N_19557);
nand U20604 (N_20604,N_19402,N_18120);
and U20605 (N_20605,N_18882,N_18562);
xnor U20606 (N_20606,N_18699,N_19452);
or U20607 (N_20607,N_19727,N_19671);
xor U20608 (N_20608,N_18709,N_19216);
nor U20609 (N_20609,N_19079,N_18003);
nand U20610 (N_20610,N_19891,N_19841);
xnor U20611 (N_20611,N_19006,N_19190);
nand U20612 (N_20612,N_19166,N_19012);
nor U20613 (N_20613,N_18091,N_18487);
and U20614 (N_20614,N_19453,N_18673);
xnor U20615 (N_20615,N_19106,N_19666);
or U20616 (N_20616,N_19496,N_18443);
or U20617 (N_20617,N_18326,N_19649);
xnor U20618 (N_20618,N_19700,N_18949);
nor U20619 (N_20619,N_18712,N_19052);
and U20620 (N_20620,N_19659,N_19001);
xnor U20621 (N_20621,N_18481,N_18410);
nand U20622 (N_20622,N_19829,N_18396);
and U20623 (N_20623,N_19978,N_19498);
or U20624 (N_20624,N_18578,N_18936);
nor U20625 (N_20625,N_19260,N_19679);
or U20626 (N_20626,N_18661,N_19208);
nor U20627 (N_20627,N_19056,N_18838);
or U20628 (N_20628,N_19640,N_18013);
nand U20629 (N_20629,N_19401,N_18215);
nand U20630 (N_20630,N_18367,N_18430);
and U20631 (N_20631,N_18100,N_19317);
and U20632 (N_20632,N_18740,N_18594);
or U20633 (N_20633,N_19890,N_19294);
nor U20634 (N_20634,N_18479,N_19698);
and U20635 (N_20635,N_18101,N_19647);
nand U20636 (N_20636,N_18791,N_18690);
and U20637 (N_20637,N_19517,N_19037);
and U20638 (N_20638,N_18254,N_18589);
nor U20639 (N_20639,N_18265,N_18887);
and U20640 (N_20640,N_19676,N_19802);
nor U20641 (N_20641,N_18317,N_18879);
and U20642 (N_20642,N_18625,N_18691);
and U20643 (N_20643,N_19395,N_18482);
nor U20644 (N_20644,N_19605,N_19179);
and U20645 (N_20645,N_18010,N_19548);
nand U20646 (N_20646,N_18309,N_18507);
nand U20647 (N_20647,N_19256,N_19024);
and U20648 (N_20648,N_18149,N_18483);
and U20649 (N_20649,N_18646,N_18343);
nand U20650 (N_20650,N_19845,N_18802);
and U20651 (N_20651,N_18137,N_18968);
and U20652 (N_20652,N_18107,N_19323);
nand U20653 (N_20653,N_18103,N_18732);
xor U20654 (N_20654,N_18502,N_19071);
xnor U20655 (N_20655,N_18494,N_19070);
xnor U20656 (N_20656,N_19211,N_19485);
xor U20657 (N_20657,N_18764,N_18386);
nor U20658 (N_20658,N_19781,N_18591);
nand U20659 (N_20659,N_19711,N_19181);
or U20660 (N_20660,N_18992,N_18717);
nor U20661 (N_20661,N_18795,N_19900);
or U20662 (N_20662,N_19872,N_18453);
xor U20663 (N_20663,N_19715,N_19370);
nor U20664 (N_20664,N_19362,N_18974);
or U20665 (N_20665,N_18130,N_18779);
nand U20666 (N_20666,N_18282,N_18884);
nand U20667 (N_20667,N_19144,N_19749);
and U20668 (N_20668,N_19480,N_18414);
nand U20669 (N_20669,N_19299,N_18818);
xnor U20670 (N_20670,N_19406,N_19046);
or U20671 (N_20671,N_18114,N_19111);
xor U20672 (N_20672,N_18957,N_19214);
nand U20673 (N_20673,N_19014,N_18044);
nand U20674 (N_20674,N_18723,N_18086);
or U20675 (N_20675,N_19879,N_18023);
and U20676 (N_20676,N_19314,N_19831);
and U20677 (N_20677,N_19490,N_18446);
or U20678 (N_20678,N_19482,N_18083);
nor U20679 (N_20679,N_19550,N_19243);
xnor U20680 (N_20680,N_18047,N_19844);
xnor U20681 (N_20681,N_18049,N_18724);
or U20682 (N_20682,N_18140,N_18448);
nand U20683 (N_20683,N_18216,N_18704);
xnor U20684 (N_20684,N_19917,N_19814);
or U20685 (N_20685,N_18711,N_19642);
or U20686 (N_20686,N_18458,N_19167);
nor U20687 (N_20687,N_18863,N_19423);
and U20688 (N_20688,N_19472,N_18198);
nor U20689 (N_20689,N_19464,N_19602);
nand U20690 (N_20690,N_18980,N_18486);
and U20691 (N_20691,N_19077,N_19589);
nand U20692 (N_20692,N_19172,N_18316);
and U20693 (N_20693,N_19201,N_18172);
xnor U20694 (N_20694,N_19766,N_18875);
and U20695 (N_20695,N_19652,N_18132);
or U20696 (N_20696,N_19355,N_19039);
or U20697 (N_20697,N_19356,N_19774);
and U20698 (N_20698,N_19185,N_18393);
or U20699 (N_20699,N_18748,N_18659);
and U20700 (N_20700,N_18116,N_18181);
and U20701 (N_20701,N_19328,N_19554);
nand U20702 (N_20702,N_18031,N_19292);
nor U20703 (N_20703,N_19924,N_18580);
or U20704 (N_20704,N_19661,N_19007);
xor U20705 (N_20705,N_18574,N_19512);
and U20706 (N_20706,N_18208,N_19974);
nor U20707 (N_20707,N_18810,N_18256);
nor U20708 (N_20708,N_19544,N_19952);
xnor U20709 (N_20709,N_18926,N_18829);
xor U20710 (N_20710,N_18485,N_18813);
xnor U20711 (N_20711,N_18022,N_19120);
nor U20712 (N_20712,N_19927,N_19380);
or U20713 (N_20713,N_19224,N_19098);
nor U20714 (N_20714,N_18745,N_18205);
or U20715 (N_20715,N_19038,N_18307);
xor U20716 (N_20716,N_18159,N_19551);
nand U20717 (N_20717,N_19121,N_19687);
or U20718 (N_20718,N_18742,N_19018);
or U20719 (N_20719,N_19217,N_19808);
nor U20720 (N_20720,N_19147,N_18941);
and U20721 (N_20721,N_18152,N_18759);
or U20722 (N_20722,N_18783,N_19914);
or U20723 (N_20723,N_19963,N_18497);
xor U20724 (N_20724,N_18241,N_19375);
and U20725 (N_20725,N_18384,N_18401);
nand U20726 (N_20726,N_18284,N_19280);
or U20727 (N_20727,N_18846,N_18036);
nand U20728 (N_20728,N_19689,N_18142);
or U20729 (N_20729,N_18518,N_18782);
nand U20730 (N_20730,N_18310,N_18444);
or U20731 (N_20731,N_18823,N_18016);
nor U20732 (N_20732,N_19654,N_19556);
and U20733 (N_20733,N_19838,N_18515);
nor U20734 (N_20734,N_19536,N_18773);
nand U20735 (N_20735,N_19995,N_19945);
and U20736 (N_20736,N_19286,N_19365);
xor U20737 (N_20737,N_19588,N_18028);
and U20738 (N_20738,N_19281,N_18984);
nand U20739 (N_20739,N_19456,N_18655);
or U20740 (N_20740,N_19601,N_18973);
or U20741 (N_20741,N_18621,N_18372);
and U20742 (N_20742,N_19685,N_19369);
nor U20743 (N_20743,N_18351,N_19354);
or U20744 (N_20744,N_18178,N_19932);
nand U20745 (N_20745,N_18464,N_19543);
nor U20746 (N_20746,N_19739,N_19578);
nor U20747 (N_20747,N_18767,N_18322);
and U20748 (N_20748,N_19523,N_18366);
or U20749 (N_20749,N_18840,N_19567);
nor U20750 (N_20750,N_18741,N_19238);
or U20751 (N_20751,N_18469,N_19964);
nand U20752 (N_20752,N_19084,N_18131);
or U20753 (N_20753,N_18694,N_19218);
or U20754 (N_20754,N_19047,N_18710);
xor U20755 (N_20755,N_19582,N_18048);
xor U20756 (N_20756,N_18784,N_19233);
nor U20757 (N_20757,N_19388,N_19028);
or U20758 (N_20758,N_19117,N_19919);
or U20759 (N_20759,N_18546,N_18872);
nand U20760 (N_20760,N_18662,N_18171);
or U20761 (N_20761,N_19723,N_18057);
or U20762 (N_20762,N_19611,N_19493);
and U20763 (N_20763,N_18627,N_18751);
nor U20764 (N_20764,N_19680,N_18720);
nor U20765 (N_20765,N_18312,N_18605);
nand U20766 (N_20766,N_19837,N_19970);
nand U20767 (N_20767,N_19950,N_19510);
xor U20768 (N_20768,N_19302,N_18753);
xor U20769 (N_20769,N_19982,N_19705);
nand U20770 (N_20770,N_19742,N_19285);
and U20771 (N_20771,N_19645,N_19921);
nor U20772 (N_20772,N_18774,N_19594);
nand U20773 (N_20773,N_18387,N_19440);
nand U20774 (N_20774,N_18558,N_18379);
nand U20775 (N_20775,N_19101,N_18219);
nor U20776 (N_20776,N_19449,N_19939);
xor U20777 (N_20777,N_18041,N_18034);
nand U20778 (N_20778,N_19473,N_18024);
xnor U20779 (N_20779,N_18327,N_18581);
or U20780 (N_20780,N_18243,N_18332);
or U20781 (N_20781,N_19420,N_18412);
or U20782 (N_20782,N_18385,N_19758);
and U20783 (N_20783,N_19058,N_18299);
and U20784 (N_20784,N_18470,N_19633);
nand U20785 (N_20785,N_18406,N_19008);
nand U20786 (N_20786,N_19196,N_19519);
xor U20787 (N_20787,N_18896,N_18134);
nand U20788 (N_20788,N_18271,N_18033);
nand U20789 (N_20789,N_18425,N_19441);
xor U20790 (N_20790,N_18318,N_19082);
nor U20791 (N_20791,N_18447,N_19278);
or U20792 (N_20792,N_18999,N_18355);
nor U20793 (N_20793,N_19712,N_18579);
nor U20794 (N_20794,N_19786,N_18026);
nand U20795 (N_20795,N_19076,N_19977);
or U20796 (N_20796,N_19612,N_19800);
nor U20797 (N_20797,N_18827,N_18474);
or U20798 (N_20798,N_18157,N_19340);
and U20799 (N_20799,N_19158,N_18330);
nand U20800 (N_20800,N_19476,N_19104);
or U20801 (N_20801,N_19348,N_19338);
nor U20802 (N_20802,N_18626,N_18769);
nand U20803 (N_20803,N_19336,N_19267);
and U20804 (N_20804,N_19915,N_18255);
nand U20805 (N_20805,N_19481,N_19010);
and U20806 (N_20806,N_18637,N_18809);
nor U20807 (N_20807,N_19073,N_18682);
nor U20808 (N_20808,N_19944,N_19905);
nor U20809 (N_20809,N_19468,N_18503);
or U20810 (N_20810,N_18113,N_19708);
nor U20811 (N_20811,N_19508,N_19422);
xnor U20812 (N_20812,N_18357,N_18700);
nand U20813 (N_20813,N_19142,N_18880);
nor U20814 (N_20814,N_19145,N_19248);
or U20815 (N_20815,N_19042,N_19415);
nor U20816 (N_20816,N_18407,N_19762);
or U20817 (N_20817,N_18221,N_19542);
nand U20818 (N_20818,N_19220,N_19942);
xor U20819 (N_20819,N_19720,N_19495);
nand U20820 (N_20820,N_19187,N_18201);
or U20821 (N_20821,N_19202,N_18128);
nand U20822 (N_20822,N_19412,N_19719);
nand U20823 (N_20823,N_19511,N_18418);
and U20824 (N_20824,N_18249,N_18616);
xnor U20825 (N_20825,N_19139,N_18085);
or U20826 (N_20826,N_18427,N_19584);
xor U20827 (N_20827,N_18934,N_19696);
nand U20828 (N_20828,N_19486,N_19620);
and U20829 (N_20829,N_19973,N_18225);
nor U20830 (N_20830,N_19346,N_19979);
nand U20831 (N_20831,N_19585,N_19573);
nand U20832 (N_20832,N_18045,N_19291);
or U20833 (N_20833,N_19150,N_18075);
xor U20834 (N_20834,N_18985,N_19430);
and U20835 (N_20835,N_18843,N_19376);
and U20836 (N_20836,N_19274,N_19114);
and U20837 (N_20837,N_19433,N_18921);
nand U20838 (N_20838,N_18339,N_19450);
xnor U20839 (N_20839,N_19461,N_19026);
nand U20840 (N_20840,N_19013,N_18826);
or U20841 (N_20841,N_19784,N_18088);
nand U20842 (N_20842,N_18356,N_18964);
and U20843 (N_20843,N_18236,N_19732);
or U20844 (N_20844,N_19153,N_18173);
or U20845 (N_20845,N_19614,N_19522);
xnor U20846 (N_20846,N_19931,N_19960);
and U20847 (N_20847,N_18645,N_19128);
nor U20848 (N_20848,N_18716,N_19853);
and U20849 (N_20849,N_19045,N_18438);
xnor U20850 (N_20850,N_19629,N_19813);
nand U20851 (N_20851,N_18918,N_18588);
xnor U20852 (N_20852,N_18151,N_19032);
nor U20853 (N_20853,N_19180,N_19436);
and U20854 (N_20854,N_19499,N_18403);
nor U20855 (N_20855,N_18657,N_18193);
and U20856 (N_20856,N_19706,N_19821);
and U20857 (N_20857,N_18744,N_19025);
nor U20858 (N_20858,N_19209,N_19424);
or U20859 (N_20859,N_18676,N_18603);
and U20860 (N_20860,N_19497,N_19990);
nand U20861 (N_20861,N_18555,N_19830);
nand U20862 (N_20862,N_18834,N_18295);
or U20863 (N_20863,N_18359,N_18778);
nand U20864 (N_20864,N_18324,N_19125);
xor U20865 (N_20865,N_19200,N_19776);
and U20866 (N_20866,N_19112,N_18663);
and U20867 (N_20867,N_18328,N_18196);
nand U20868 (N_20868,N_19435,N_19868);
nor U20869 (N_20869,N_19862,N_19590);
nor U20870 (N_20870,N_19906,N_18529);
nor U20871 (N_20871,N_18874,N_19325);
xnor U20872 (N_20872,N_18897,N_19658);
xnor U20873 (N_20873,N_18501,N_18436);
nand U20874 (N_20874,N_18986,N_19475);
xor U20875 (N_20875,N_18270,N_19494);
nor U20876 (N_20876,N_18188,N_18856);
and U20877 (N_20877,N_19938,N_19398);
or U20878 (N_20878,N_19684,N_19988);
or U20879 (N_20879,N_19509,N_18460);
nor U20880 (N_20880,N_19537,N_19790);
or U20881 (N_20881,N_19538,N_18183);
xor U20882 (N_20882,N_18250,N_18733);
xor U20883 (N_20883,N_19198,N_19384);
or U20884 (N_20884,N_18292,N_18660);
and U20885 (N_20885,N_19303,N_18981);
xnor U20886 (N_20886,N_19833,N_18786);
and U20887 (N_20887,N_19764,N_18451);
nand U20888 (N_20888,N_18730,N_19947);
nand U20889 (N_20889,N_18423,N_18812);
nor U20890 (N_20890,N_19632,N_19396);
nor U20891 (N_20891,N_19624,N_19622);
or U20892 (N_20892,N_18850,N_18539);
or U20893 (N_20893,N_18671,N_19363);
nand U20894 (N_20894,N_19244,N_18692);
nand U20895 (N_20895,N_18349,N_19672);
nor U20896 (N_20896,N_19405,N_18242);
and U20897 (N_20897,N_18727,N_18046);
or U20898 (N_20898,N_18415,N_19427);
or U20899 (N_20899,N_19772,N_19331);
nand U20900 (N_20900,N_19627,N_18454);
nor U20901 (N_20901,N_18413,N_18672);
nand U20902 (N_20902,N_19541,N_18463);
or U20903 (N_20903,N_19206,N_19804);
nor U20904 (N_20904,N_18547,N_18099);
xnor U20905 (N_20905,N_18369,N_18693);
nand U20906 (N_20906,N_18304,N_18651);
xnor U20907 (N_20907,N_18825,N_19378);
nor U20908 (N_20908,N_19069,N_18002);
and U20909 (N_20909,N_18112,N_19969);
or U20910 (N_20910,N_18899,N_19253);
nand U20911 (N_20911,N_19741,N_19438);
nor U20912 (N_20912,N_19457,N_19791);
and U20913 (N_20913,N_19103,N_19599);
nand U20914 (N_20914,N_18923,N_18785);
or U20915 (N_20915,N_19311,N_19532);
and U20916 (N_20916,N_18056,N_18532);
nand U20917 (N_20917,N_18325,N_19865);
and U20918 (N_20918,N_18429,N_18668);
nor U20919 (N_20919,N_19133,N_18476);
or U20920 (N_20920,N_19115,N_19956);
xor U20921 (N_20921,N_19165,N_18535);
xor U20922 (N_20922,N_19717,N_19043);
nand U20923 (N_20923,N_19961,N_19525);
nor U20924 (N_20924,N_19020,N_18670);
and U20925 (N_20925,N_18758,N_19284);
or U20926 (N_20926,N_18248,N_18380);
and U20927 (N_20927,N_19306,N_19834);
nor U20928 (N_20928,N_19663,N_19783);
or U20929 (N_20929,N_19151,N_19825);
nor U20930 (N_20930,N_18920,N_18754);
xor U20931 (N_20931,N_18186,N_19835);
xnor U20932 (N_20932,N_19559,N_18258);
xor U20933 (N_20933,N_18191,N_19367);
xnor U20934 (N_20934,N_19930,N_19146);
nand U20935 (N_20935,N_18072,N_19044);
nor U20936 (N_20936,N_18969,N_18301);
nor U20937 (N_20937,N_19182,N_19571);
and U20938 (N_20938,N_19339,N_19566);
nand U20939 (N_20939,N_18293,N_18623);
nor U20940 (N_20940,N_19321,N_18192);
nand U20941 (N_20941,N_19628,N_18587);
and U20942 (N_20942,N_19320,N_18948);
xnor U20943 (N_20943,N_19194,N_18038);
and U20944 (N_20944,N_19801,N_19250);
nor U20945 (N_20945,N_18959,N_18768);
nor U20946 (N_20946,N_18550,N_18911);
nand U20947 (N_20947,N_18852,N_18006);
nor U20948 (N_20948,N_19846,N_18323);
or U20949 (N_20949,N_19426,N_18928);
nand U20950 (N_20950,N_19371,N_18197);
nand U20951 (N_20951,N_19345,N_19887);
and U20952 (N_20952,N_19343,N_18982);
and U20953 (N_20953,N_19353,N_19003);
xor U20954 (N_20954,N_18638,N_19413);
xor U20955 (N_20955,N_19847,N_19347);
and U20956 (N_20956,N_19088,N_19817);
and U20957 (N_20957,N_18223,N_18908);
xnor U20958 (N_20958,N_19000,N_18794);
or U20959 (N_20959,N_18439,N_19467);
nand U20960 (N_20960,N_18607,N_19269);
and U20961 (N_20961,N_19469,N_19483);
nor U20962 (N_20962,N_18798,N_18944);
and U20963 (N_20963,N_18305,N_18995);
nor U20964 (N_20964,N_18991,N_18841);
nand U20965 (N_20965,N_18859,N_19907);
nand U20966 (N_20966,N_19065,N_18967);
xnor U20967 (N_20967,N_19287,N_19855);
or U20968 (N_20968,N_18777,N_18521);
or U20969 (N_20969,N_18498,N_18450);
nand U20970 (N_20970,N_19809,N_18561);
or U20971 (N_20971,N_19531,N_19364);
xor U20972 (N_20972,N_19751,N_18919);
nand U20973 (N_20973,N_19229,N_18214);
and U20974 (N_20974,N_19061,N_19533);
nor U20975 (N_20975,N_18488,N_18353);
and U20976 (N_20976,N_19102,N_18064);
and U20977 (N_20977,N_18997,N_19262);
and U20978 (N_20978,N_18750,N_18569);
nor U20979 (N_20979,N_19683,N_19419);
or U20980 (N_20980,N_18417,N_18461);
and U20981 (N_20981,N_19725,N_18125);
xor U20982 (N_20982,N_18685,N_18428);
nor U20983 (N_20983,N_19265,N_18499);
xor U20984 (N_20984,N_19173,N_18628);
xnor U20985 (N_20985,N_19161,N_18477);
and U20986 (N_20986,N_18528,N_19418);
and U20987 (N_20987,N_19621,N_18738);
or U20988 (N_20988,N_18945,N_18531);
xnor U20989 (N_20989,N_18419,N_18218);
and U20990 (N_20990,N_18653,N_18212);
or U20991 (N_20991,N_19333,N_18177);
xor U20992 (N_20992,N_18473,N_18903);
xor U20993 (N_20993,N_18735,N_18734);
nor U20994 (N_20994,N_18746,N_19270);
or U20995 (N_20995,N_18025,N_19110);
or U20996 (N_20996,N_19897,N_19688);
nand U20997 (N_20997,N_18378,N_19002);
xnor U20998 (N_20998,N_19107,N_18475);
or U20999 (N_20999,N_18641,N_19851);
or U21000 (N_21000,N_19647,N_18891);
xnor U21001 (N_21001,N_19389,N_19876);
and U21002 (N_21002,N_18583,N_19422);
nand U21003 (N_21003,N_19380,N_18978);
nor U21004 (N_21004,N_18575,N_18559);
xnor U21005 (N_21005,N_19727,N_18179);
or U21006 (N_21006,N_19193,N_19375);
nand U21007 (N_21007,N_18445,N_18605);
nor U21008 (N_21008,N_18384,N_19688);
nand U21009 (N_21009,N_19036,N_18014);
nor U21010 (N_21010,N_18696,N_18723);
nand U21011 (N_21011,N_19351,N_18349);
nand U21012 (N_21012,N_19512,N_19822);
nor U21013 (N_21013,N_18455,N_19481);
and U21014 (N_21014,N_19998,N_19006);
xor U21015 (N_21015,N_18978,N_18476);
and U21016 (N_21016,N_18652,N_19329);
or U21017 (N_21017,N_19989,N_19690);
nor U21018 (N_21018,N_19264,N_19786);
nand U21019 (N_21019,N_18515,N_19772);
nor U21020 (N_21020,N_19172,N_19755);
and U21021 (N_21021,N_19078,N_18563);
nor U21022 (N_21022,N_19492,N_19789);
nor U21023 (N_21023,N_19171,N_18751);
and U21024 (N_21024,N_19099,N_19423);
xor U21025 (N_21025,N_19265,N_19453);
nor U21026 (N_21026,N_19721,N_18727);
or U21027 (N_21027,N_18295,N_18206);
nand U21028 (N_21028,N_18933,N_18309);
nand U21029 (N_21029,N_19065,N_18331);
nor U21030 (N_21030,N_18655,N_19806);
nor U21031 (N_21031,N_19465,N_18390);
nand U21032 (N_21032,N_19588,N_19790);
nand U21033 (N_21033,N_18250,N_19210);
and U21034 (N_21034,N_19108,N_18721);
nand U21035 (N_21035,N_18741,N_18562);
or U21036 (N_21036,N_18266,N_18229);
xnor U21037 (N_21037,N_18677,N_18579);
xnor U21038 (N_21038,N_18018,N_18508);
and U21039 (N_21039,N_19680,N_19519);
xor U21040 (N_21040,N_19728,N_18276);
or U21041 (N_21041,N_18492,N_18142);
and U21042 (N_21042,N_19779,N_18767);
nor U21043 (N_21043,N_18667,N_18394);
xor U21044 (N_21044,N_19096,N_19504);
xnor U21045 (N_21045,N_19993,N_19669);
or U21046 (N_21046,N_18494,N_19753);
or U21047 (N_21047,N_19046,N_19554);
and U21048 (N_21048,N_18132,N_19454);
and U21049 (N_21049,N_18276,N_19763);
nor U21050 (N_21050,N_18979,N_19727);
nor U21051 (N_21051,N_18028,N_19531);
or U21052 (N_21052,N_19188,N_18912);
xnor U21053 (N_21053,N_18256,N_19715);
xor U21054 (N_21054,N_18444,N_19386);
xor U21055 (N_21055,N_18898,N_18646);
and U21056 (N_21056,N_19484,N_19291);
nand U21057 (N_21057,N_18642,N_19408);
nor U21058 (N_21058,N_18873,N_19638);
and U21059 (N_21059,N_18653,N_19858);
or U21060 (N_21060,N_18434,N_18016);
nor U21061 (N_21061,N_19090,N_18058);
nor U21062 (N_21062,N_18686,N_18213);
or U21063 (N_21063,N_18355,N_18767);
nand U21064 (N_21064,N_18398,N_19875);
xnor U21065 (N_21065,N_18402,N_18836);
nand U21066 (N_21066,N_18402,N_18105);
nand U21067 (N_21067,N_18874,N_18899);
nand U21068 (N_21068,N_19158,N_18822);
or U21069 (N_21069,N_19691,N_19696);
xor U21070 (N_21070,N_19028,N_19095);
nor U21071 (N_21071,N_19833,N_19007);
nor U21072 (N_21072,N_18961,N_19021);
and U21073 (N_21073,N_19308,N_18733);
and U21074 (N_21074,N_18034,N_19896);
nand U21075 (N_21075,N_19536,N_18635);
nand U21076 (N_21076,N_19427,N_19711);
nor U21077 (N_21077,N_18341,N_19468);
nor U21078 (N_21078,N_18018,N_18084);
xnor U21079 (N_21079,N_19268,N_19579);
xnor U21080 (N_21080,N_18402,N_18227);
or U21081 (N_21081,N_18704,N_18472);
nor U21082 (N_21082,N_18759,N_19768);
xnor U21083 (N_21083,N_19096,N_18701);
nor U21084 (N_21084,N_18240,N_18297);
or U21085 (N_21085,N_18569,N_18735);
nor U21086 (N_21086,N_18423,N_19592);
or U21087 (N_21087,N_18184,N_18116);
nor U21088 (N_21088,N_19357,N_18139);
nand U21089 (N_21089,N_19234,N_19026);
nor U21090 (N_21090,N_18357,N_18289);
xor U21091 (N_21091,N_18158,N_19552);
nor U21092 (N_21092,N_18734,N_19743);
nor U21093 (N_21093,N_18392,N_18941);
nor U21094 (N_21094,N_18229,N_18660);
nor U21095 (N_21095,N_18643,N_18355);
nor U21096 (N_21096,N_18738,N_18117);
xnor U21097 (N_21097,N_18820,N_18386);
or U21098 (N_21098,N_18993,N_19579);
nand U21099 (N_21099,N_19400,N_18316);
nor U21100 (N_21100,N_18346,N_18866);
and U21101 (N_21101,N_18645,N_18036);
xnor U21102 (N_21102,N_19357,N_19246);
and U21103 (N_21103,N_18742,N_19614);
nor U21104 (N_21104,N_18136,N_18468);
or U21105 (N_21105,N_19385,N_18830);
xnor U21106 (N_21106,N_18462,N_18761);
nand U21107 (N_21107,N_18925,N_19158);
or U21108 (N_21108,N_19323,N_18756);
nand U21109 (N_21109,N_19417,N_19164);
xor U21110 (N_21110,N_19849,N_19351);
and U21111 (N_21111,N_18154,N_18218);
and U21112 (N_21112,N_18632,N_19334);
or U21113 (N_21113,N_18695,N_18708);
xnor U21114 (N_21114,N_19797,N_19191);
and U21115 (N_21115,N_18660,N_19821);
xnor U21116 (N_21116,N_19880,N_18427);
xor U21117 (N_21117,N_18754,N_18662);
and U21118 (N_21118,N_18862,N_19553);
nor U21119 (N_21119,N_18914,N_19021);
and U21120 (N_21120,N_19540,N_18896);
or U21121 (N_21121,N_19520,N_18770);
xnor U21122 (N_21122,N_18613,N_19224);
or U21123 (N_21123,N_19160,N_19398);
or U21124 (N_21124,N_18837,N_19204);
nor U21125 (N_21125,N_19186,N_18096);
nor U21126 (N_21126,N_19453,N_18543);
nand U21127 (N_21127,N_19570,N_19760);
nand U21128 (N_21128,N_18107,N_18110);
nor U21129 (N_21129,N_18150,N_19179);
nor U21130 (N_21130,N_19716,N_19085);
or U21131 (N_21131,N_19087,N_18996);
xnor U21132 (N_21132,N_19624,N_18463);
nor U21133 (N_21133,N_18442,N_18249);
xnor U21134 (N_21134,N_19130,N_19284);
nor U21135 (N_21135,N_19741,N_19787);
and U21136 (N_21136,N_19132,N_19531);
nand U21137 (N_21137,N_19787,N_18317);
nand U21138 (N_21138,N_19510,N_18089);
xnor U21139 (N_21139,N_19104,N_18524);
nand U21140 (N_21140,N_18050,N_18832);
nand U21141 (N_21141,N_19930,N_18450);
nand U21142 (N_21142,N_18352,N_19191);
xor U21143 (N_21143,N_18968,N_18268);
xnor U21144 (N_21144,N_19487,N_19493);
or U21145 (N_21145,N_19479,N_18514);
nand U21146 (N_21146,N_19760,N_19669);
xnor U21147 (N_21147,N_19383,N_18919);
or U21148 (N_21148,N_19904,N_19168);
xnor U21149 (N_21149,N_18916,N_18296);
xnor U21150 (N_21150,N_18424,N_18764);
xnor U21151 (N_21151,N_18055,N_18445);
xnor U21152 (N_21152,N_19358,N_19997);
nand U21153 (N_21153,N_18726,N_19421);
and U21154 (N_21154,N_19685,N_18997);
nand U21155 (N_21155,N_18276,N_18147);
nand U21156 (N_21156,N_18601,N_19697);
xor U21157 (N_21157,N_18475,N_18209);
and U21158 (N_21158,N_19750,N_18844);
xor U21159 (N_21159,N_19694,N_19113);
nor U21160 (N_21160,N_18858,N_18082);
xnor U21161 (N_21161,N_18573,N_18830);
nand U21162 (N_21162,N_19117,N_19292);
nor U21163 (N_21163,N_19521,N_19626);
xor U21164 (N_21164,N_19042,N_18630);
nor U21165 (N_21165,N_18373,N_18093);
nor U21166 (N_21166,N_19213,N_19234);
xnor U21167 (N_21167,N_18224,N_19000);
nor U21168 (N_21168,N_19754,N_19961);
nor U21169 (N_21169,N_19577,N_18012);
or U21170 (N_21170,N_18109,N_19878);
and U21171 (N_21171,N_18531,N_19643);
and U21172 (N_21172,N_19780,N_18842);
nand U21173 (N_21173,N_18615,N_18583);
or U21174 (N_21174,N_18703,N_19972);
xor U21175 (N_21175,N_18172,N_18153);
xnor U21176 (N_21176,N_19746,N_19985);
nor U21177 (N_21177,N_19378,N_18451);
nor U21178 (N_21178,N_18631,N_19464);
nor U21179 (N_21179,N_19810,N_18825);
nand U21180 (N_21180,N_19164,N_19551);
nor U21181 (N_21181,N_19919,N_19052);
nand U21182 (N_21182,N_18758,N_18566);
or U21183 (N_21183,N_19864,N_18395);
nand U21184 (N_21184,N_18520,N_18415);
or U21185 (N_21185,N_19303,N_18899);
nand U21186 (N_21186,N_19764,N_18773);
and U21187 (N_21187,N_18252,N_19884);
nor U21188 (N_21188,N_19557,N_18163);
nor U21189 (N_21189,N_18081,N_18430);
or U21190 (N_21190,N_18119,N_19906);
nand U21191 (N_21191,N_19528,N_19254);
or U21192 (N_21192,N_19988,N_19109);
and U21193 (N_21193,N_18201,N_18881);
xor U21194 (N_21194,N_19587,N_18313);
xnor U21195 (N_21195,N_19465,N_18428);
nand U21196 (N_21196,N_19302,N_19356);
nor U21197 (N_21197,N_18480,N_18365);
and U21198 (N_21198,N_19037,N_18959);
and U21199 (N_21199,N_19394,N_19483);
nor U21200 (N_21200,N_19649,N_19954);
nor U21201 (N_21201,N_18268,N_18896);
or U21202 (N_21202,N_18763,N_19512);
and U21203 (N_21203,N_19644,N_19162);
nor U21204 (N_21204,N_18951,N_18930);
and U21205 (N_21205,N_18248,N_19958);
nand U21206 (N_21206,N_18830,N_19941);
or U21207 (N_21207,N_19772,N_18443);
nor U21208 (N_21208,N_18069,N_19619);
nand U21209 (N_21209,N_19282,N_18905);
nand U21210 (N_21210,N_19337,N_19823);
nand U21211 (N_21211,N_19898,N_19320);
xor U21212 (N_21212,N_19924,N_19293);
nor U21213 (N_21213,N_19160,N_19161);
xor U21214 (N_21214,N_19230,N_19909);
xor U21215 (N_21215,N_18951,N_18708);
and U21216 (N_21216,N_18135,N_18491);
nor U21217 (N_21217,N_19455,N_18871);
or U21218 (N_21218,N_18349,N_18408);
and U21219 (N_21219,N_19091,N_18640);
or U21220 (N_21220,N_18719,N_18484);
nor U21221 (N_21221,N_19796,N_19937);
and U21222 (N_21222,N_18807,N_19635);
and U21223 (N_21223,N_18858,N_19909);
or U21224 (N_21224,N_18547,N_19235);
nor U21225 (N_21225,N_18010,N_19701);
and U21226 (N_21226,N_19828,N_19926);
nand U21227 (N_21227,N_18847,N_19559);
nor U21228 (N_21228,N_19348,N_19054);
nor U21229 (N_21229,N_19432,N_18375);
nand U21230 (N_21230,N_19353,N_18063);
and U21231 (N_21231,N_18205,N_18109);
and U21232 (N_21232,N_18496,N_19919);
xor U21233 (N_21233,N_19184,N_18567);
and U21234 (N_21234,N_19763,N_19469);
and U21235 (N_21235,N_18499,N_18707);
xor U21236 (N_21236,N_19522,N_18809);
and U21237 (N_21237,N_19244,N_18170);
and U21238 (N_21238,N_19368,N_19215);
and U21239 (N_21239,N_19200,N_18941);
xnor U21240 (N_21240,N_19839,N_19986);
or U21241 (N_21241,N_18272,N_18330);
xnor U21242 (N_21242,N_19655,N_19732);
xnor U21243 (N_21243,N_18646,N_19904);
xor U21244 (N_21244,N_19277,N_19325);
or U21245 (N_21245,N_19588,N_19999);
and U21246 (N_21246,N_19742,N_18730);
nor U21247 (N_21247,N_18358,N_19779);
xnor U21248 (N_21248,N_19577,N_19553);
xnor U21249 (N_21249,N_18539,N_19061);
nand U21250 (N_21250,N_18456,N_19890);
nand U21251 (N_21251,N_18794,N_18910);
nor U21252 (N_21252,N_18759,N_19022);
xor U21253 (N_21253,N_19232,N_19112);
or U21254 (N_21254,N_19592,N_18838);
and U21255 (N_21255,N_18513,N_19551);
nor U21256 (N_21256,N_18805,N_19827);
nor U21257 (N_21257,N_18027,N_19057);
xor U21258 (N_21258,N_19008,N_19866);
nand U21259 (N_21259,N_18089,N_19552);
nor U21260 (N_21260,N_19771,N_19032);
or U21261 (N_21261,N_19085,N_18123);
or U21262 (N_21262,N_18445,N_18371);
xor U21263 (N_21263,N_19762,N_18097);
or U21264 (N_21264,N_19978,N_18170);
nand U21265 (N_21265,N_18867,N_18354);
or U21266 (N_21266,N_18804,N_18891);
and U21267 (N_21267,N_19094,N_18522);
nor U21268 (N_21268,N_19070,N_19854);
or U21269 (N_21269,N_19328,N_19509);
xnor U21270 (N_21270,N_19395,N_19126);
nand U21271 (N_21271,N_18549,N_19090);
and U21272 (N_21272,N_19472,N_19888);
nand U21273 (N_21273,N_18934,N_19155);
nor U21274 (N_21274,N_18936,N_18510);
xnor U21275 (N_21275,N_19199,N_18106);
or U21276 (N_21276,N_19914,N_18801);
xnor U21277 (N_21277,N_18122,N_18003);
xnor U21278 (N_21278,N_18297,N_18076);
nand U21279 (N_21279,N_19434,N_19004);
or U21280 (N_21280,N_19444,N_19203);
xor U21281 (N_21281,N_18360,N_18435);
nand U21282 (N_21282,N_19560,N_19047);
or U21283 (N_21283,N_18368,N_18253);
xor U21284 (N_21284,N_19904,N_18662);
and U21285 (N_21285,N_19041,N_18215);
and U21286 (N_21286,N_19135,N_18460);
xor U21287 (N_21287,N_19978,N_18994);
or U21288 (N_21288,N_19858,N_18212);
nor U21289 (N_21289,N_18709,N_19721);
or U21290 (N_21290,N_18058,N_19720);
nor U21291 (N_21291,N_18511,N_18949);
nor U21292 (N_21292,N_18428,N_18690);
and U21293 (N_21293,N_18886,N_18081);
nand U21294 (N_21294,N_19338,N_18292);
nor U21295 (N_21295,N_19077,N_19869);
nor U21296 (N_21296,N_19976,N_18815);
nand U21297 (N_21297,N_19981,N_18513);
xnor U21298 (N_21298,N_18621,N_19972);
and U21299 (N_21299,N_19617,N_19253);
or U21300 (N_21300,N_19429,N_18206);
xnor U21301 (N_21301,N_19919,N_19256);
or U21302 (N_21302,N_19834,N_18254);
or U21303 (N_21303,N_19989,N_18398);
nand U21304 (N_21304,N_19399,N_19574);
and U21305 (N_21305,N_19864,N_19028);
and U21306 (N_21306,N_19814,N_18723);
xor U21307 (N_21307,N_18923,N_18050);
nor U21308 (N_21308,N_19894,N_19201);
nor U21309 (N_21309,N_18972,N_19552);
nor U21310 (N_21310,N_18604,N_19017);
and U21311 (N_21311,N_19999,N_18752);
nand U21312 (N_21312,N_19447,N_19199);
nor U21313 (N_21313,N_18959,N_19058);
xnor U21314 (N_21314,N_18749,N_19661);
xnor U21315 (N_21315,N_18533,N_19576);
or U21316 (N_21316,N_19905,N_19591);
or U21317 (N_21317,N_18296,N_19796);
nand U21318 (N_21318,N_18927,N_18369);
or U21319 (N_21319,N_18661,N_19232);
xor U21320 (N_21320,N_18646,N_19910);
or U21321 (N_21321,N_18482,N_19859);
xnor U21322 (N_21322,N_18973,N_18542);
and U21323 (N_21323,N_18773,N_19867);
nand U21324 (N_21324,N_18051,N_19331);
xnor U21325 (N_21325,N_19931,N_18973);
nor U21326 (N_21326,N_19503,N_18235);
xnor U21327 (N_21327,N_19745,N_19812);
and U21328 (N_21328,N_18417,N_19433);
xor U21329 (N_21329,N_18682,N_19299);
nor U21330 (N_21330,N_18407,N_19072);
and U21331 (N_21331,N_18400,N_18609);
nand U21332 (N_21332,N_19639,N_19816);
nor U21333 (N_21333,N_18933,N_18502);
and U21334 (N_21334,N_18218,N_19432);
or U21335 (N_21335,N_19858,N_18175);
xnor U21336 (N_21336,N_19749,N_19323);
or U21337 (N_21337,N_19050,N_19337);
nand U21338 (N_21338,N_18265,N_18704);
xor U21339 (N_21339,N_18208,N_19093);
or U21340 (N_21340,N_19632,N_18484);
and U21341 (N_21341,N_19324,N_18604);
xor U21342 (N_21342,N_19757,N_18072);
and U21343 (N_21343,N_19165,N_18257);
and U21344 (N_21344,N_19023,N_18124);
nor U21345 (N_21345,N_19907,N_18297);
xnor U21346 (N_21346,N_18032,N_19878);
nand U21347 (N_21347,N_18257,N_19185);
and U21348 (N_21348,N_18938,N_19416);
xor U21349 (N_21349,N_18816,N_18948);
xnor U21350 (N_21350,N_19128,N_19554);
nand U21351 (N_21351,N_19309,N_18433);
and U21352 (N_21352,N_19407,N_19232);
and U21353 (N_21353,N_19022,N_18360);
and U21354 (N_21354,N_18901,N_18187);
nand U21355 (N_21355,N_19258,N_18552);
nor U21356 (N_21356,N_19115,N_18467);
nor U21357 (N_21357,N_18979,N_19459);
nor U21358 (N_21358,N_19215,N_19540);
nand U21359 (N_21359,N_19172,N_18793);
or U21360 (N_21360,N_18176,N_18576);
xnor U21361 (N_21361,N_19448,N_19437);
and U21362 (N_21362,N_19116,N_18166);
or U21363 (N_21363,N_18099,N_18623);
nor U21364 (N_21364,N_19209,N_18290);
or U21365 (N_21365,N_18195,N_18678);
and U21366 (N_21366,N_19830,N_19998);
nor U21367 (N_21367,N_19393,N_19675);
or U21368 (N_21368,N_19936,N_18501);
xor U21369 (N_21369,N_18495,N_19359);
and U21370 (N_21370,N_18035,N_19960);
nor U21371 (N_21371,N_19913,N_18227);
nor U21372 (N_21372,N_18049,N_19887);
or U21373 (N_21373,N_19482,N_19537);
and U21374 (N_21374,N_18316,N_18383);
xnor U21375 (N_21375,N_19532,N_19126);
nor U21376 (N_21376,N_19911,N_18146);
and U21377 (N_21377,N_18649,N_18696);
nor U21378 (N_21378,N_19510,N_19875);
nor U21379 (N_21379,N_19598,N_18983);
nand U21380 (N_21380,N_18689,N_19988);
xor U21381 (N_21381,N_18356,N_18319);
or U21382 (N_21382,N_19826,N_19488);
nand U21383 (N_21383,N_18116,N_19051);
xnor U21384 (N_21384,N_19190,N_18676);
and U21385 (N_21385,N_18000,N_19225);
and U21386 (N_21386,N_18916,N_18906);
and U21387 (N_21387,N_18691,N_19172);
nand U21388 (N_21388,N_18018,N_18183);
xnor U21389 (N_21389,N_19378,N_19848);
or U21390 (N_21390,N_19989,N_19583);
and U21391 (N_21391,N_19510,N_18554);
nand U21392 (N_21392,N_19215,N_18688);
or U21393 (N_21393,N_19509,N_18074);
or U21394 (N_21394,N_18602,N_18310);
or U21395 (N_21395,N_19517,N_19817);
nor U21396 (N_21396,N_18094,N_19703);
xor U21397 (N_21397,N_18356,N_18148);
nor U21398 (N_21398,N_19006,N_18977);
and U21399 (N_21399,N_18563,N_18775);
nor U21400 (N_21400,N_18744,N_18725);
nand U21401 (N_21401,N_18310,N_18489);
xor U21402 (N_21402,N_18118,N_19003);
nand U21403 (N_21403,N_19733,N_18521);
nand U21404 (N_21404,N_18772,N_19502);
nor U21405 (N_21405,N_19248,N_19976);
or U21406 (N_21406,N_19743,N_18324);
nand U21407 (N_21407,N_18046,N_18424);
nor U21408 (N_21408,N_19535,N_18724);
nor U21409 (N_21409,N_18105,N_18891);
nor U21410 (N_21410,N_19050,N_19452);
nand U21411 (N_21411,N_19101,N_19512);
or U21412 (N_21412,N_18798,N_18503);
and U21413 (N_21413,N_19301,N_19489);
nand U21414 (N_21414,N_18829,N_19315);
nand U21415 (N_21415,N_19944,N_18154);
nor U21416 (N_21416,N_19256,N_19585);
nor U21417 (N_21417,N_19363,N_19259);
and U21418 (N_21418,N_18502,N_19997);
nand U21419 (N_21419,N_19279,N_19672);
and U21420 (N_21420,N_19603,N_19479);
nor U21421 (N_21421,N_19191,N_19063);
nand U21422 (N_21422,N_19415,N_19350);
nand U21423 (N_21423,N_19160,N_18543);
or U21424 (N_21424,N_19628,N_19122);
nor U21425 (N_21425,N_19313,N_19950);
nand U21426 (N_21426,N_19147,N_18507);
nand U21427 (N_21427,N_19937,N_19462);
nor U21428 (N_21428,N_19975,N_19737);
and U21429 (N_21429,N_18252,N_19541);
or U21430 (N_21430,N_18453,N_19278);
nor U21431 (N_21431,N_18143,N_18092);
nand U21432 (N_21432,N_19830,N_18545);
xnor U21433 (N_21433,N_18080,N_18899);
xor U21434 (N_21434,N_19241,N_19693);
or U21435 (N_21435,N_18085,N_19262);
xor U21436 (N_21436,N_18628,N_19671);
and U21437 (N_21437,N_18826,N_19295);
nor U21438 (N_21438,N_19611,N_18791);
xor U21439 (N_21439,N_18320,N_19266);
or U21440 (N_21440,N_18728,N_19473);
or U21441 (N_21441,N_19193,N_18265);
and U21442 (N_21442,N_18978,N_18531);
nand U21443 (N_21443,N_19652,N_19644);
xnor U21444 (N_21444,N_18378,N_18019);
nor U21445 (N_21445,N_18369,N_18051);
xor U21446 (N_21446,N_19305,N_19627);
or U21447 (N_21447,N_19809,N_18565);
nor U21448 (N_21448,N_18864,N_19958);
nor U21449 (N_21449,N_18942,N_18712);
and U21450 (N_21450,N_18002,N_18931);
nand U21451 (N_21451,N_18891,N_19326);
xor U21452 (N_21452,N_19365,N_19766);
nand U21453 (N_21453,N_19415,N_19978);
or U21454 (N_21454,N_19650,N_19998);
or U21455 (N_21455,N_19330,N_19524);
and U21456 (N_21456,N_18474,N_19426);
nand U21457 (N_21457,N_19885,N_19650);
and U21458 (N_21458,N_18836,N_18406);
or U21459 (N_21459,N_18618,N_19055);
xnor U21460 (N_21460,N_19039,N_18053);
xnor U21461 (N_21461,N_18706,N_18356);
xor U21462 (N_21462,N_18876,N_19590);
nor U21463 (N_21463,N_19574,N_19361);
nor U21464 (N_21464,N_19244,N_18976);
xor U21465 (N_21465,N_19089,N_19413);
nand U21466 (N_21466,N_19485,N_18699);
nand U21467 (N_21467,N_18440,N_19572);
xor U21468 (N_21468,N_18626,N_18823);
xnor U21469 (N_21469,N_18380,N_18063);
nand U21470 (N_21470,N_18988,N_18375);
nor U21471 (N_21471,N_19761,N_18543);
xnor U21472 (N_21472,N_18800,N_19706);
nor U21473 (N_21473,N_19135,N_18607);
xnor U21474 (N_21474,N_19056,N_19700);
nand U21475 (N_21475,N_19746,N_18221);
nor U21476 (N_21476,N_19082,N_19819);
nand U21477 (N_21477,N_19097,N_18230);
xor U21478 (N_21478,N_18288,N_19458);
xnor U21479 (N_21479,N_19988,N_19098);
nand U21480 (N_21480,N_18921,N_19101);
or U21481 (N_21481,N_19690,N_19655);
nand U21482 (N_21482,N_18653,N_18861);
nand U21483 (N_21483,N_18520,N_19978);
or U21484 (N_21484,N_18212,N_18889);
or U21485 (N_21485,N_19745,N_19287);
xnor U21486 (N_21486,N_19943,N_18072);
and U21487 (N_21487,N_18528,N_18165);
or U21488 (N_21488,N_19859,N_19078);
and U21489 (N_21489,N_18462,N_19040);
nand U21490 (N_21490,N_19465,N_19478);
xor U21491 (N_21491,N_18829,N_18392);
and U21492 (N_21492,N_18376,N_18430);
nor U21493 (N_21493,N_19876,N_19443);
nor U21494 (N_21494,N_18746,N_19599);
and U21495 (N_21495,N_18653,N_18223);
and U21496 (N_21496,N_19744,N_19689);
nor U21497 (N_21497,N_18677,N_18819);
xnor U21498 (N_21498,N_19313,N_19270);
and U21499 (N_21499,N_18031,N_18014);
and U21500 (N_21500,N_18555,N_19145);
nand U21501 (N_21501,N_19595,N_18800);
nor U21502 (N_21502,N_18374,N_19654);
nand U21503 (N_21503,N_18840,N_19733);
or U21504 (N_21504,N_19339,N_19749);
nor U21505 (N_21505,N_19047,N_19804);
and U21506 (N_21506,N_19974,N_19500);
and U21507 (N_21507,N_18647,N_18915);
nand U21508 (N_21508,N_19239,N_19214);
and U21509 (N_21509,N_18920,N_19856);
nor U21510 (N_21510,N_19079,N_19516);
and U21511 (N_21511,N_19795,N_18910);
nor U21512 (N_21512,N_18630,N_18843);
and U21513 (N_21513,N_19289,N_19446);
xor U21514 (N_21514,N_18208,N_19029);
xor U21515 (N_21515,N_18633,N_19561);
nand U21516 (N_21516,N_19730,N_19063);
and U21517 (N_21517,N_19632,N_19800);
or U21518 (N_21518,N_19221,N_18655);
or U21519 (N_21519,N_18366,N_18319);
and U21520 (N_21520,N_19693,N_19237);
and U21521 (N_21521,N_19320,N_18831);
or U21522 (N_21522,N_18404,N_19778);
xor U21523 (N_21523,N_18554,N_19626);
and U21524 (N_21524,N_18962,N_18861);
and U21525 (N_21525,N_18566,N_18325);
or U21526 (N_21526,N_19160,N_18244);
nor U21527 (N_21527,N_18042,N_18535);
xnor U21528 (N_21528,N_19102,N_18582);
or U21529 (N_21529,N_19911,N_19223);
nor U21530 (N_21530,N_19980,N_18639);
or U21531 (N_21531,N_19581,N_18047);
and U21532 (N_21532,N_18074,N_18331);
nand U21533 (N_21533,N_18139,N_19048);
nand U21534 (N_21534,N_18925,N_19744);
nor U21535 (N_21535,N_19909,N_18459);
xnor U21536 (N_21536,N_19986,N_18185);
or U21537 (N_21537,N_18663,N_19589);
nand U21538 (N_21538,N_19009,N_18601);
xnor U21539 (N_21539,N_18058,N_19178);
nor U21540 (N_21540,N_19368,N_18454);
and U21541 (N_21541,N_18034,N_18273);
or U21542 (N_21542,N_19202,N_19657);
nand U21543 (N_21543,N_19319,N_18270);
and U21544 (N_21544,N_18293,N_18382);
nor U21545 (N_21545,N_19039,N_19781);
nand U21546 (N_21546,N_18862,N_19614);
and U21547 (N_21547,N_18754,N_19836);
nand U21548 (N_21548,N_18849,N_18901);
and U21549 (N_21549,N_18374,N_18248);
xnor U21550 (N_21550,N_19156,N_18361);
or U21551 (N_21551,N_19959,N_19111);
nand U21552 (N_21552,N_18193,N_18189);
xnor U21553 (N_21553,N_19209,N_19062);
nor U21554 (N_21554,N_19846,N_19844);
or U21555 (N_21555,N_19293,N_19292);
xnor U21556 (N_21556,N_18055,N_19931);
nand U21557 (N_21557,N_18201,N_18363);
and U21558 (N_21558,N_18978,N_19891);
or U21559 (N_21559,N_18454,N_19244);
nor U21560 (N_21560,N_18208,N_19893);
nor U21561 (N_21561,N_19154,N_19708);
nand U21562 (N_21562,N_19179,N_19612);
and U21563 (N_21563,N_19840,N_19132);
xnor U21564 (N_21564,N_19239,N_19119);
nand U21565 (N_21565,N_19784,N_19286);
or U21566 (N_21566,N_18857,N_19785);
nor U21567 (N_21567,N_19979,N_18051);
xnor U21568 (N_21568,N_18544,N_18313);
and U21569 (N_21569,N_18278,N_19205);
and U21570 (N_21570,N_19339,N_19930);
or U21571 (N_21571,N_19050,N_19320);
and U21572 (N_21572,N_18239,N_19670);
and U21573 (N_21573,N_18620,N_19921);
or U21574 (N_21574,N_19452,N_19241);
xnor U21575 (N_21575,N_19233,N_18372);
nor U21576 (N_21576,N_19953,N_18544);
nor U21577 (N_21577,N_18162,N_19161);
nand U21578 (N_21578,N_19094,N_18449);
xor U21579 (N_21579,N_19997,N_18759);
and U21580 (N_21580,N_19216,N_19775);
nand U21581 (N_21581,N_19789,N_19156);
nor U21582 (N_21582,N_18450,N_19904);
or U21583 (N_21583,N_18268,N_19124);
nand U21584 (N_21584,N_18527,N_18882);
nand U21585 (N_21585,N_19515,N_18492);
nand U21586 (N_21586,N_18471,N_19081);
nor U21587 (N_21587,N_19640,N_19394);
xnor U21588 (N_21588,N_19587,N_19642);
or U21589 (N_21589,N_19853,N_18393);
and U21590 (N_21590,N_19546,N_18896);
and U21591 (N_21591,N_19444,N_19652);
nor U21592 (N_21592,N_18602,N_18573);
xor U21593 (N_21593,N_19362,N_19917);
and U21594 (N_21594,N_19028,N_19269);
nand U21595 (N_21595,N_18145,N_18033);
xnor U21596 (N_21596,N_18277,N_18188);
or U21597 (N_21597,N_19870,N_19721);
or U21598 (N_21598,N_19637,N_18883);
or U21599 (N_21599,N_18427,N_18164);
and U21600 (N_21600,N_18259,N_18040);
nand U21601 (N_21601,N_18353,N_18417);
nor U21602 (N_21602,N_18762,N_18454);
nor U21603 (N_21603,N_19788,N_18583);
or U21604 (N_21604,N_19536,N_18479);
nand U21605 (N_21605,N_18798,N_18258);
nand U21606 (N_21606,N_18426,N_18783);
or U21607 (N_21607,N_18779,N_19684);
nor U21608 (N_21608,N_19172,N_18714);
nor U21609 (N_21609,N_18469,N_18846);
nor U21610 (N_21610,N_18904,N_18883);
nand U21611 (N_21611,N_18426,N_18802);
xor U21612 (N_21612,N_19192,N_19834);
nor U21613 (N_21613,N_19641,N_18292);
and U21614 (N_21614,N_18606,N_19078);
and U21615 (N_21615,N_18231,N_18446);
or U21616 (N_21616,N_18657,N_18549);
xor U21617 (N_21617,N_19592,N_19191);
and U21618 (N_21618,N_18030,N_18777);
nor U21619 (N_21619,N_18705,N_18706);
and U21620 (N_21620,N_19369,N_19442);
nand U21621 (N_21621,N_19892,N_19949);
nor U21622 (N_21622,N_19347,N_18042);
xor U21623 (N_21623,N_19761,N_19082);
or U21624 (N_21624,N_19981,N_18822);
nand U21625 (N_21625,N_19589,N_19862);
nor U21626 (N_21626,N_19113,N_19700);
and U21627 (N_21627,N_19778,N_19332);
and U21628 (N_21628,N_19177,N_19175);
and U21629 (N_21629,N_19445,N_18379);
nor U21630 (N_21630,N_19829,N_19120);
nand U21631 (N_21631,N_19609,N_18651);
xnor U21632 (N_21632,N_18293,N_18826);
and U21633 (N_21633,N_18400,N_19678);
nand U21634 (N_21634,N_18163,N_19000);
nor U21635 (N_21635,N_19173,N_19419);
or U21636 (N_21636,N_18822,N_19500);
or U21637 (N_21637,N_19875,N_18021);
or U21638 (N_21638,N_19485,N_19000);
and U21639 (N_21639,N_18123,N_18549);
nor U21640 (N_21640,N_18458,N_19845);
nand U21641 (N_21641,N_19488,N_18238);
nor U21642 (N_21642,N_19444,N_18160);
nand U21643 (N_21643,N_19007,N_18065);
or U21644 (N_21644,N_18885,N_19139);
or U21645 (N_21645,N_18842,N_19395);
or U21646 (N_21646,N_19501,N_18623);
and U21647 (N_21647,N_19353,N_19818);
xor U21648 (N_21648,N_19968,N_19701);
xor U21649 (N_21649,N_18969,N_18048);
nor U21650 (N_21650,N_19939,N_19510);
or U21651 (N_21651,N_18858,N_19076);
xnor U21652 (N_21652,N_18260,N_18989);
nand U21653 (N_21653,N_19810,N_19419);
nor U21654 (N_21654,N_18379,N_18237);
nor U21655 (N_21655,N_18275,N_18889);
nor U21656 (N_21656,N_19353,N_19528);
or U21657 (N_21657,N_19987,N_19963);
xnor U21658 (N_21658,N_18503,N_18718);
xnor U21659 (N_21659,N_18647,N_19561);
and U21660 (N_21660,N_19975,N_19821);
or U21661 (N_21661,N_19895,N_19238);
and U21662 (N_21662,N_18828,N_19218);
xnor U21663 (N_21663,N_19006,N_19073);
or U21664 (N_21664,N_18595,N_18159);
or U21665 (N_21665,N_18011,N_18782);
xnor U21666 (N_21666,N_19339,N_18556);
and U21667 (N_21667,N_18206,N_18468);
xnor U21668 (N_21668,N_18231,N_19900);
and U21669 (N_21669,N_19583,N_19842);
nand U21670 (N_21670,N_18178,N_19987);
xor U21671 (N_21671,N_18786,N_18315);
xnor U21672 (N_21672,N_18531,N_19036);
or U21673 (N_21673,N_19890,N_19707);
and U21674 (N_21674,N_18449,N_19209);
or U21675 (N_21675,N_19229,N_19857);
xnor U21676 (N_21676,N_19114,N_18193);
or U21677 (N_21677,N_18083,N_19804);
xor U21678 (N_21678,N_19911,N_18819);
nor U21679 (N_21679,N_18260,N_19388);
or U21680 (N_21680,N_18248,N_18121);
nand U21681 (N_21681,N_19533,N_18974);
nand U21682 (N_21682,N_18122,N_19036);
xor U21683 (N_21683,N_18736,N_19594);
nor U21684 (N_21684,N_18284,N_18741);
xnor U21685 (N_21685,N_18155,N_19731);
and U21686 (N_21686,N_19516,N_18651);
nand U21687 (N_21687,N_18978,N_18685);
or U21688 (N_21688,N_19624,N_18065);
or U21689 (N_21689,N_18578,N_19037);
or U21690 (N_21690,N_19754,N_18643);
xor U21691 (N_21691,N_19505,N_18539);
and U21692 (N_21692,N_18375,N_18825);
xnor U21693 (N_21693,N_19813,N_19042);
xor U21694 (N_21694,N_18333,N_18837);
and U21695 (N_21695,N_18806,N_19590);
or U21696 (N_21696,N_18528,N_18828);
and U21697 (N_21697,N_19048,N_19079);
xor U21698 (N_21698,N_18101,N_19060);
nand U21699 (N_21699,N_19792,N_19297);
xor U21700 (N_21700,N_19367,N_18941);
xnor U21701 (N_21701,N_18537,N_19444);
or U21702 (N_21702,N_19765,N_19990);
xnor U21703 (N_21703,N_19572,N_18046);
nand U21704 (N_21704,N_19126,N_18417);
nand U21705 (N_21705,N_18369,N_18581);
xor U21706 (N_21706,N_19031,N_18652);
and U21707 (N_21707,N_18394,N_18856);
and U21708 (N_21708,N_19988,N_18925);
xor U21709 (N_21709,N_19789,N_19844);
or U21710 (N_21710,N_19537,N_19304);
and U21711 (N_21711,N_18409,N_19783);
nor U21712 (N_21712,N_19295,N_18706);
or U21713 (N_21713,N_18487,N_19947);
xor U21714 (N_21714,N_18153,N_18693);
or U21715 (N_21715,N_19142,N_19578);
and U21716 (N_21716,N_18006,N_19692);
or U21717 (N_21717,N_19186,N_19417);
nor U21718 (N_21718,N_19852,N_19990);
or U21719 (N_21719,N_19703,N_19621);
nand U21720 (N_21720,N_19281,N_18803);
nor U21721 (N_21721,N_18855,N_19980);
or U21722 (N_21722,N_18138,N_19856);
or U21723 (N_21723,N_19866,N_18134);
nand U21724 (N_21724,N_19767,N_18891);
and U21725 (N_21725,N_18511,N_19742);
or U21726 (N_21726,N_18879,N_18527);
nand U21727 (N_21727,N_18026,N_18898);
and U21728 (N_21728,N_18731,N_18098);
xnor U21729 (N_21729,N_19525,N_19600);
nor U21730 (N_21730,N_18298,N_19369);
and U21731 (N_21731,N_19784,N_18010);
xor U21732 (N_21732,N_19647,N_19775);
or U21733 (N_21733,N_18614,N_19498);
xor U21734 (N_21734,N_19070,N_18155);
or U21735 (N_21735,N_18542,N_18611);
nand U21736 (N_21736,N_19102,N_18251);
or U21737 (N_21737,N_18830,N_19104);
nor U21738 (N_21738,N_18545,N_19817);
nor U21739 (N_21739,N_19824,N_19048);
xnor U21740 (N_21740,N_18181,N_19909);
nor U21741 (N_21741,N_18223,N_19293);
xor U21742 (N_21742,N_19770,N_18153);
nor U21743 (N_21743,N_19223,N_19935);
nor U21744 (N_21744,N_18050,N_19995);
and U21745 (N_21745,N_19420,N_19378);
xnor U21746 (N_21746,N_19488,N_18112);
or U21747 (N_21747,N_19154,N_19307);
or U21748 (N_21748,N_18766,N_18343);
nor U21749 (N_21749,N_18241,N_18127);
xor U21750 (N_21750,N_19871,N_19044);
xor U21751 (N_21751,N_19689,N_18971);
xnor U21752 (N_21752,N_19349,N_18406);
nand U21753 (N_21753,N_18886,N_18101);
or U21754 (N_21754,N_19353,N_18122);
or U21755 (N_21755,N_19088,N_18834);
nor U21756 (N_21756,N_19043,N_18939);
nor U21757 (N_21757,N_19212,N_18490);
or U21758 (N_21758,N_19601,N_19188);
xnor U21759 (N_21759,N_19191,N_18410);
nor U21760 (N_21760,N_19865,N_18175);
xnor U21761 (N_21761,N_18880,N_19876);
nand U21762 (N_21762,N_19597,N_18709);
xor U21763 (N_21763,N_18742,N_19788);
nand U21764 (N_21764,N_18181,N_19105);
nand U21765 (N_21765,N_18992,N_19852);
nand U21766 (N_21766,N_19978,N_19164);
nand U21767 (N_21767,N_18498,N_18474);
nor U21768 (N_21768,N_19910,N_18503);
and U21769 (N_21769,N_19166,N_19146);
nor U21770 (N_21770,N_18227,N_18065);
and U21771 (N_21771,N_19220,N_18290);
nor U21772 (N_21772,N_19360,N_19973);
nor U21773 (N_21773,N_19730,N_19722);
nand U21774 (N_21774,N_19487,N_19447);
or U21775 (N_21775,N_19381,N_19090);
nand U21776 (N_21776,N_19547,N_18497);
xnor U21777 (N_21777,N_19178,N_18945);
xnor U21778 (N_21778,N_18783,N_18900);
xnor U21779 (N_21779,N_19654,N_18723);
nand U21780 (N_21780,N_18259,N_18064);
and U21781 (N_21781,N_18259,N_19806);
nand U21782 (N_21782,N_18700,N_19431);
nor U21783 (N_21783,N_18545,N_18334);
and U21784 (N_21784,N_19600,N_19902);
nor U21785 (N_21785,N_19666,N_19812);
and U21786 (N_21786,N_19605,N_18034);
nor U21787 (N_21787,N_19140,N_18182);
and U21788 (N_21788,N_18666,N_19667);
nand U21789 (N_21789,N_18566,N_18417);
xnor U21790 (N_21790,N_18076,N_18672);
or U21791 (N_21791,N_18630,N_19823);
nor U21792 (N_21792,N_19748,N_18654);
xor U21793 (N_21793,N_19837,N_18881);
nand U21794 (N_21794,N_18871,N_19051);
nand U21795 (N_21795,N_18244,N_18407);
nor U21796 (N_21796,N_18692,N_18451);
and U21797 (N_21797,N_19542,N_18605);
nor U21798 (N_21798,N_19945,N_19029);
nor U21799 (N_21799,N_18080,N_18030);
and U21800 (N_21800,N_19062,N_19613);
nor U21801 (N_21801,N_18944,N_18534);
and U21802 (N_21802,N_19039,N_19452);
nor U21803 (N_21803,N_19154,N_18008);
or U21804 (N_21804,N_19329,N_19916);
xnor U21805 (N_21805,N_19974,N_18088);
nand U21806 (N_21806,N_19969,N_18156);
xor U21807 (N_21807,N_19647,N_19985);
xnor U21808 (N_21808,N_19176,N_19610);
nor U21809 (N_21809,N_18789,N_19738);
xnor U21810 (N_21810,N_18850,N_18287);
and U21811 (N_21811,N_19610,N_18298);
and U21812 (N_21812,N_18582,N_18433);
or U21813 (N_21813,N_19246,N_19127);
xor U21814 (N_21814,N_18803,N_18576);
and U21815 (N_21815,N_19798,N_19809);
xnor U21816 (N_21816,N_18102,N_18275);
nand U21817 (N_21817,N_19141,N_18143);
nor U21818 (N_21818,N_18906,N_19327);
and U21819 (N_21819,N_19689,N_18613);
or U21820 (N_21820,N_19337,N_19689);
and U21821 (N_21821,N_19550,N_18292);
nor U21822 (N_21822,N_19707,N_18786);
nand U21823 (N_21823,N_18721,N_19238);
nor U21824 (N_21824,N_19862,N_19560);
and U21825 (N_21825,N_19310,N_18350);
xnor U21826 (N_21826,N_19593,N_19861);
and U21827 (N_21827,N_18226,N_18693);
and U21828 (N_21828,N_18189,N_19239);
nor U21829 (N_21829,N_19867,N_18814);
or U21830 (N_21830,N_18961,N_18722);
or U21831 (N_21831,N_19877,N_19664);
or U21832 (N_21832,N_19938,N_18679);
or U21833 (N_21833,N_18409,N_18538);
xor U21834 (N_21834,N_19041,N_18515);
xnor U21835 (N_21835,N_18160,N_18583);
and U21836 (N_21836,N_19033,N_18351);
nor U21837 (N_21837,N_18859,N_18144);
or U21838 (N_21838,N_19834,N_18603);
xor U21839 (N_21839,N_18644,N_18483);
nand U21840 (N_21840,N_19198,N_19566);
nand U21841 (N_21841,N_19025,N_18568);
nand U21842 (N_21842,N_19530,N_18663);
xor U21843 (N_21843,N_19490,N_19779);
nor U21844 (N_21844,N_18939,N_19173);
xnor U21845 (N_21845,N_19626,N_19007);
xnor U21846 (N_21846,N_18172,N_19628);
nand U21847 (N_21847,N_18018,N_19883);
xnor U21848 (N_21848,N_18114,N_18794);
and U21849 (N_21849,N_19212,N_19167);
and U21850 (N_21850,N_19272,N_19623);
or U21851 (N_21851,N_19075,N_18824);
nor U21852 (N_21852,N_19396,N_18284);
or U21853 (N_21853,N_18043,N_18667);
or U21854 (N_21854,N_18841,N_19992);
nor U21855 (N_21855,N_18885,N_18797);
and U21856 (N_21856,N_19737,N_18982);
or U21857 (N_21857,N_18910,N_19977);
or U21858 (N_21858,N_19800,N_18596);
nor U21859 (N_21859,N_18155,N_19323);
nand U21860 (N_21860,N_18642,N_19871);
or U21861 (N_21861,N_18649,N_18896);
nand U21862 (N_21862,N_19433,N_19773);
or U21863 (N_21863,N_18173,N_18654);
xnor U21864 (N_21864,N_18688,N_18539);
xor U21865 (N_21865,N_19725,N_19576);
nand U21866 (N_21866,N_18568,N_18230);
nand U21867 (N_21867,N_19437,N_18964);
xnor U21868 (N_21868,N_19142,N_18480);
nand U21869 (N_21869,N_19765,N_19903);
nor U21870 (N_21870,N_19093,N_18233);
or U21871 (N_21871,N_18868,N_19051);
nor U21872 (N_21872,N_18625,N_19448);
nor U21873 (N_21873,N_19061,N_18581);
or U21874 (N_21874,N_19307,N_19379);
xnor U21875 (N_21875,N_18681,N_18087);
nor U21876 (N_21876,N_18177,N_19842);
nor U21877 (N_21877,N_18150,N_18335);
or U21878 (N_21878,N_19540,N_19477);
or U21879 (N_21879,N_19777,N_19323);
or U21880 (N_21880,N_18040,N_18821);
or U21881 (N_21881,N_19626,N_18562);
xor U21882 (N_21882,N_19252,N_18842);
or U21883 (N_21883,N_18233,N_18965);
or U21884 (N_21884,N_19468,N_19636);
and U21885 (N_21885,N_18333,N_18593);
and U21886 (N_21886,N_19774,N_19592);
nand U21887 (N_21887,N_18830,N_18132);
nor U21888 (N_21888,N_18849,N_19325);
or U21889 (N_21889,N_18266,N_18275);
xnor U21890 (N_21890,N_18954,N_18242);
or U21891 (N_21891,N_19104,N_18456);
nor U21892 (N_21892,N_19470,N_19371);
xor U21893 (N_21893,N_19214,N_18252);
xnor U21894 (N_21894,N_18428,N_18619);
and U21895 (N_21895,N_19275,N_19244);
nand U21896 (N_21896,N_18120,N_19303);
or U21897 (N_21897,N_19022,N_19584);
and U21898 (N_21898,N_19002,N_18930);
or U21899 (N_21899,N_19059,N_18466);
xnor U21900 (N_21900,N_19789,N_18614);
and U21901 (N_21901,N_18780,N_19952);
xnor U21902 (N_21902,N_19954,N_19973);
nand U21903 (N_21903,N_18185,N_19493);
nor U21904 (N_21904,N_19442,N_19850);
nand U21905 (N_21905,N_19057,N_19261);
nand U21906 (N_21906,N_19383,N_19573);
or U21907 (N_21907,N_18982,N_18537);
nor U21908 (N_21908,N_19732,N_18363);
xor U21909 (N_21909,N_19874,N_18084);
xnor U21910 (N_21910,N_18982,N_18854);
nor U21911 (N_21911,N_19529,N_19916);
nor U21912 (N_21912,N_19066,N_19751);
xor U21913 (N_21913,N_19881,N_18535);
nand U21914 (N_21914,N_18395,N_19758);
and U21915 (N_21915,N_18374,N_19124);
xnor U21916 (N_21916,N_19242,N_19039);
nor U21917 (N_21917,N_18192,N_19465);
nor U21918 (N_21918,N_19709,N_18099);
xnor U21919 (N_21919,N_19588,N_19833);
or U21920 (N_21920,N_19670,N_19709);
or U21921 (N_21921,N_19089,N_18537);
xor U21922 (N_21922,N_18280,N_18582);
nor U21923 (N_21923,N_19981,N_18008);
and U21924 (N_21924,N_19512,N_19835);
nor U21925 (N_21925,N_18942,N_18953);
nor U21926 (N_21926,N_19953,N_19845);
or U21927 (N_21927,N_18186,N_18662);
nand U21928 (N_21928,N_18597,N_19296);
or U21929 (N_21929,N_19284,N_19465);
xor U21930 (N_21930,N_18029,N_19329);
or U21931 (N_21931,N_18261,N_18677);
xor U21932 (N_21932,N_18203,N_19479);
or U21933 (N_21933,N_18850,N_18833);
nand U21934 (N_21934,N_19543,N_19718);
or U21935 (N_21935,N_19791,N_18820);
and U21936 (N_21936,N_18459,N_19943);
and U21937 (N_21937,N_18720,N_18231);
nand U21938 (N_21938,N_19796,N_18206);
or U21939 (N_21939,N_19658,N_18500);
nand U21940 (N_21940,N_18046,N_19564);
and U21941 (N_21941,N_18095,N_19046);
xnor U21942 (N_21942,N_18678,N_18924);
nor U21943 (N_21943,N_19148,N_19035);
and U21944 (N_21944,N_19919,N_18057);
and U21945 (N_21945,N_18389,N_19831);
xnor U21946 (N_21946,N_19304,N_18756);
nand U21947 (N_21947,N_19625,N_18096);
and U21948 (N_21948,N_18364,N_18409);
or U21949 (N_21949,N_19817,N_18593);
nor U21950 (N_21950,N_18989,N_18377);
and U21951 (N_21951,N_19228,N_18005);
nor U21952 (N_21952,N_19193,N_19513);
and U21953 (N_21953,N_18232,N_19743);
nor U21954 (N_21954,N_18942,N_19644);
xor U21955 (N_21955,N_18670,N_19645);
and U21956 (N_21956,N_18852,N_18090);
nor U21957 (N_21957,N_18290,N_18825);
or U21958 (N_21958,N_18844,N_19031);
or U21959 (N_21959,N_18635,N_19772);
or U21960 (N_21960,N_18957,N_18636);
nand U21961 (N_21961,N_19227,N_18547);
and U21962 (N_21962,N_18002,N_19705);
or U21963 (N_21963,N_19769,N_18674);
nand U21964 (N_21964,N_18984,N_18502);
or U21965 (N_21965,N_19829,N_19780);
nand U21966 (N_21966,N_19722,N_18175);
nand U21967 (N_21967,N_19374,N_18991);
xnor U21968 (N_21968,N_18852,N_18626);
xnor U21969 (N_21969,N_18404,N_19736);
nor U21970 (N_21970,N_19053,N_18179);
and U21971 (N_21971,N_19337,N_18142);
nor U21972 (N_21972,N_19181,N_18127);
nand U21973 (N_21973,N_19475,N_18374);
xor U21974 (N_21974,N_19272,N_18160);
and U21975 (N_21975,N_19926,N_18925);
xor U21976 (N_21976,N_18280,N_18041);
and U21977 (N_21977,N_18409,N_18929);
xor U21978 (N_21978,N_18828,N_18837);
nand U21979 (N_21979,N_19728,N_19712);
nor U21980 (N_21980,N_19271,N_19156);
xnor U21981 (N_21981,N_19114,N_19316);
nand U21982 (N_21982,N_18517,N_19956);
nor U21983 (N_21983,N_19431,N_19328);
xor U21984 (N_21984,N_18093,N_19319);
or U21985 (N_21985,N_18029,N_18065);
nor U21986 (N_21986,N_18709,N_19868);
nor U21987 (N_21987,N_18283,N_18064);
and U21988 (N_21988,N_19148,N_19346);
nor U21989 (N_21989,N_18341,N_18736);
and U21990 (N_21990,N_19323,N_19238);
nand U21991 (N_21991,N_19199,N_19326);
and U21992 (N_21992,N_19275,N_19834);
xor U21993 (N_21993,N_19761,N_19635);
and U21994 (N_21994,N_19461,N_18943);
nand U21995 (N_21995,N_19636,N_19104);
and U21996 (N_21996,N_19440,N_19914);
or U21997 (N_21997,N_18623,N_19293);
xor U21998 (N_21998,N_18976,N_19759);
xnor U21999 (N_21999,N_19281,N_18751);
or U22000 (N_22000,N_20199,N_20428);
nand U22001 (N_22001,N_20554,N_21943);
xnor U22002 (N_22002,N_21307,N_21839);
nand U22003 (N_22003,N_20018,N_20780);
nor U22004 (N_22004,N_21893,N_21583);
nand U22005 (N_22005,N_21041,N_20241);
xor U22006 (N_22006,N_20253,N_21766);
nor U22007 (N_22007,N_20771,N_21762);
nand U22008 (N_22008,N_20161,N_21536);
nand U22009 (N_22009,N_21309,N_21894);
or U22010 (N_22010,N_20165,N_20297);
xnor U22011 (N_22011,N_21807,N_20633);
nor U22012 (N_22012,N_21021,N_21574);
or U22013 (N_22013,N_20107,N_20468);
nand U22014 (N_22014,N_21968,N_21280);
nand U22015 (N_22015,N_21055,N_20840);
or U22016 (N_22016,N_21863,N_21678);
nor U22017 (N_22017,N_21520,N_21936);
nor U22018 (N_22018,N_20869,N_21902);
nor U22019 (N_22019,N_21376,N_21578);
or U22020 (N_22020,N_20605,N_20630);
xor U22021 (N_22021,N_21587,N_20908);
or U22022 (N_22022,N_21764,N_21805);
nand U22023 (N_22023,N_21413,N_21684);
and U22024 (N_22024,N_20470,N_20155);
xnor U22025 (N_22025,N_20287,N_21328);
or U22026 (N_22026,N_21987,N_20369);
nor U22027 (N_22027,N_21469,N_20009);
and U22028 (N_22028,N_21551,N_21000);
nor U22029 (N_22029,N_21605,N_20601);
nand U22030 (N_22030,N_20613,N_20383);
and U22031 (N_22031,N_20117,N_20250);
nor U22032 (N_22032,N_20657,N_20964);
or U22033 (N_22033,N_21282,N_21478);
xor U22034 (N_22034,N_21316,N_20717);
or U22035 (N_22035,N_21142,N_20285);
nand U22036 (N_22036,N_20077,N_21734);
and U22037 (N_22037,N_20409,N_21366);
or U22038 (N_22038,N_20019,N_20041);
or U22039 (N_22039,N_21899,N_21339);
nand U22040 (N_22040,N_20776,N_20321);
nor U22041 (N_22041,N_21405,N_21354);
nand U22042 (N_22042,N_20288,N_20478);
xor U22043 (N_22043,N_20080,N_21873);
nor U22044 (N_22044,N_20184,N_20035);
or U22045 (N_22045,N_21849,N_20769);
or U22046 (N_22046,N_21862,N_20294);
nand U22047 (N_22047,N_20420,N_21927);
or U22048 (N_22048,N_21275,N_21278);
or U22049 (N_22049,N_21485,N_20812);
xor U22050 (N_22050,N_20538,N_20988);
or U22051 (N_22051,N_21080,N_21958);
and U22052 (N_22052,N_21804,N_20309);
xor U22053 (N_22053,N_20263,N_20786);
and U22054 (N_22054,N_20295,N_20759);
or U22055 (N_22055,N_21547,N_21130);
nand U22056 (N_22056,N_21812,N_21314);
xor U22057 (N_22057,N_20473,N_21815);
or U22058 (N_22058,N_20971,N_21263);
xor U22059 (N_22059,N_20389,N_21476);
and U22060 (N_22060,N_21452,N_21267);
nor U22061 (N_22061,N_20673,N_20900);
nand U22062 (N_22062,N_20083,N_21774);
and U22063 (N_22063,N_20331,N_21479);
and U22064 (N_22064,N_20247,N_20011);
or U22065 (N_22065,N_21090,N_21779);
nand U22066 (N_22066,N_21879,N_21922);
and U22067 (N_22067,N_21198,N_21036);
xor U22068 (N_22068,N_21778,N_21518);
or U22069 (N_22069,N_20274,N_20319);
and U22070 (N_22070,N_21072,N_21160);
or U22071 (N_22071,N_21477,N_20043);
nor U22072 (N_22072,N_20230,N_21591);
nor U22073 (N_22073,N_21269,N_20884);
nand U22074 (N_22074,N_21207,N_20562);
or U22075 (N_22075,N_21004,N_20976);
or U22076 (N_22076,N_20890,N_21357);
xnor U22077 (N_22077,N_21896,N_20355);
nor U22078 (N_22078,N_21486,N_20663);
nor U22079 (N_22079,N_21363,N_20111);
nand U22080 (N_22080,N_21049,N_20029);
or U22081 (N_22081,N_21881,N_21315);
xnor U22082 (N_22082,N_20645,N_21819);
nor U22083 (N_22083,N_20593,N_20940);
xor U22084 (N_22084,N_21277,N_21209);
and U22085 (N_22085,N_20387,N_21175);
or U22086 (N_22086,N_21064,N_21969);
xor U22087 (N_22087,N_21204,N_20201);
nor U22088 (N_22088,N_21631,N_21341);
or U22089 (N_22089,N_21996,N_21797);
or U22090 (N_22090,N_20815,N_20374);
xnor U22091 (N_22091,N_20008,N_21506);
nor U22092 (N_22092,N_20547,N_20179);
nand U22093 (N_22093,N_21830,N_20923);
nand U22094 (N_22094,N_21012,N_20053);
nand U22095 (N_22095,N_21388,N_20049);
xnor U22096 (N_22096,N_21622,N_20298);
or U22097 (N_22097,N_21870,N_20166);
nor U22098 (N_22098,N_21095,N_21763);
nor U22099 (N_22099,N_20436,N_21098);
nor U22100 (N_22100,N_21407,N_21818);
xnor U22101 (N_22101,N_20252,N_21116);
and U22102 (N_22102,N_21192,N_21777);
and U22103 (N_22103,N_20114,N_20454);
xor U22104 (N_22104,N_20664,N_20316);
or U22105 (N_22105,N_21153,N_21543);
and U22106 (N_22106,N_20157,N_20025);
nor U22107 (N_22107,N_21850,N_20723);
nor U22108 (N_22108,N_20343,N_20045);
xnor U22109 (N_22109,N_21361,N_21385);
xnor U22110 (N_22110,N_20079,N_20680);
nor U22111 (N_22111,N_21632,N_21032);
nor U22112 (N_22112,N_21473,N_21855);
and U22113 (N_22113,N_20956,N_21352);
or U22114 (N_22114,N_20609,N_21738);
nor U22115 (N_22115,N_21445,N_21458);
and U22116 (N_22116,N_20286,N_21402);
nor U22117 (N_22117,N_20983,N_20887);
nand U22118 (N_22118,N_21414,N_20540);
xnor U22119 (N_22119,N_21338,N_20856);
nor U22120 (N_22120,N_21063,N_20846);
nand U22121 (N_22121,N_20278,N_21441);
or U22122 (N_22122,N_21600,N_20792);
or U22123 (N_22123,N_21735,N_21795);
or U22124 (N_22124,N_21531,N_20365);
or U22125 (N_22125,N_20777,N_21725);
and U22126 (N_22126,N_20926,N_21723);
nand U22127 (N_22127,N_21444,N_21661);
nor U22128 (N_22128,N_20359,N_20406);
nor U22129 (N_22129,N_21107,N_20026);
nand U22130 (N_22130,N_20619,N_20655);
nor U22131 (N_22131,N_20262,N_20251);
nor U22132 (N_22132,N_21918,N_21742);
xnor U22133 (N_22133,N_21746,N_20283);
nor U22134 (N_22134,N_20575,N_20271);
and U22135 (N_22135,N_20174,N_21285);
xor U22136 (N_22136,N_20508,N_21966);
xnor U22137 (N_22137,N_21645,N_21718);
xnor U22138 (N_22138,N_21939,N_20266);
and U22139 (N_22139,N_20170,N_20830);
and U22140 (N_22140,N_20496,N_21369);
nand U22141 (N_22141,N_21471,N_21292);
xnor U22142 (N_22142,N_20967,N_20275);
nand U22143 (N_22143,N_21571,N_20751);
nor U22144 (N_22144,N_21279,N_21685);
nor U22145 (N_22145,N_20293,N_21644);
xor U22146 (N_22146,N_20537,N_21935);
and U22147 (N_22147,N_20465,N_20951);
nor U22148 (N_22148,N_21078,N_20906);
nor U22149 (N_22149,N_20950,N_21853);
and U22150 (N_22150,N_20914,N_21817);
and U22151 (N_22151,N_20353,N_21604);
and U22152 (N_22152,N_20513,N_20895);
nand U22153 (N_22153,N_20533,N_20329);
and U22154 (N_22154,N_20587,N_21878);
and U22155 (N_22155,N_21652,N_21650);
xnor U22156 (N_22156,N_21651,N_20373);
nor U22157 (N_22157,N_21491,N_21629);
nand U22158 (N_22158,N_20621,N_21861);
nand U22159 (N_22159,N_20440,N_20485);
or U22160 (N_22160,N_21877,N_20054);
or U22161 (N_22161,N_21362,N_20300);
xnor U22162 (N_22162,N_21851,N_20418);
nor U22163 (N_22163,N_21635,N_20238);
nor U22164 (N_22164,N_21865,N_20710);
xnor U22165 (N_22165,N_20958,N_21970);
or U22166 (N_22166,N_20231,N_21435);
and U22167 (N_22167,N_20809,N_20567);
nor U22168 (N_22168,N_20131,N_21433);
or U22169 (N_22169,N_20864,N_20385);
nand U22170 (N_22170,N_20367,N_21378);
and U22171 (N_22171,N_21769,N_21609);
xnor U22172 (N_22172,N_21731,N_20076);
nor U22173 (N_22173,N_21466,N_21711);
and U22174 (N_22174,N_20223,N_20731);
xnor U22175 (N_22175,N_20291,N_20909);
and U22176 (N_22176,N_20344,N_20039);
xnor U22177 (N_22177,N_20766,N_20475);
nor U22178 (N_22178,N_21581,N_20474);
or U22179 (N_22179,N_21132,N_20614);
xnor U22180 (N_22180,N_21229,N_20681);
xnor U22181 (N_22181,N_21082,N_20878);
nand U22182 (N_22182,N_21977,N_21391);
xnor U22183 (N_22183,N_20469,N_21736);
nor U22184 (N_22184,N_20948,N_21519);
nand U22185 (N_22185,N_20313,N_20433);
and U22186 (N_22186,N_21249,N_20563);
xor U22187 (N_22187,N_21416,N_20495);
xor U22188 (N_22188,N_21146,N_20590);
or U22189 (N_22189,N_21962,N_20596);
xor U22190 (N_22190,N_21166,N_20486);
or U22191 (N_22191,N_21748,N_20110);
nor U22192 (N_22192,N_21179,N_21035);
nor U22193 (N_22193,N_20396,N_20512);
nand U22194 (N_22194,N_21147,N_20328);
and U22195 (N_22195,N_21811,N_21342);
and U22196 (N_22196,N_20228,N_21755);
or U22197 (N_22197,N_21848,N_20397);
nor U22198 (N_22198,N_20637,N_21750);
nor U22199 (N_22199,N_21127,N_20943);
nor U22200 (N_22200,N_21905,N_21022);
or U22201 (N_22201,N_21462,N_21360);
nand U22202 (N_22202,N_20548,N_21323);
xor U22203 (N_22203,N_20591,N_21013);
xor U22204 (N_22204,N_21490,N_21601);
xor U22205 (N_22205,N_21525,N_21934);
nand U22206 (N_22206,N_21890,N_21505);
nor U22207 (N_22207,N_20569,N_20642);
nor U22208 (N_22208,N_20349,N_20330);
or U22209 (N_22209,N_20209,N_21657);
or U22210 (N_22210,N_20744,N_21251);
xnor U22211 (N_22211,N_21690,N_20518);
and U22212 (N_22212,N_20484,N_21659);
nor U22213 (N_22213,N_21771,N_20933);
xor U22214 (N_22214,N_21534,N_20280);
or U22215 (N_22215,N_20753,N_21548);
or U22216 (N_22216,N_20444,N_21387);
nor U22217 (N_22217,N_20629,N_21216);
and U22218 (N_22218,N_21410,N_21183);
or U22219 (N_22219,N_20075,N_20171);
and U22220 (N_22220,N_20212,N_21372);
xnor U22221 (N_22221,N_20868,N_21048);
nand U22222 (N_22222,N_21171,N_21232);
and U22223 (N_22223,N_20921,N_20739);
and U22224 (N_22224,N_20497,N_20380);
or U22225 (N_22225,N_20123,N_20765);
and U22226 (N_22226,N_20081,N_21170);
nand U22227 (N_22227,N_20880,N_20832);
and U22228 (N_22228,N_21060,N_21428);
xor U22229 (N_22229,N_21621,N_21973);
or U22230 (N_22230,N_20066,N_20381);
nor U22231 (N_22231,N_20222,N_21355);
and U22232 (N_22232,N_21038,N_20192);
nor U22233 (N_22233,N_20867,N_21240);
and U22234 (N_22234,N_21912,N_21886);
or U22235 (N_22235,N_21223,N_20233);
or U22236 (N_22236,N_20499,N_20694);
nor U22237 (N_22237,N_20748,N_20145);
or U22238 (N_22238,N_20997,N_20617);
and U22239 (N_22239,N_20762,N_21834);
xnor U22240 (N_22240,N_20189,N_20141);
xnor U22241 (N_22241,N_20795,N_21727);
xor U22242 (N_22242,N_20341,N_20531);
and U22243 (N_22243,N_21539,N_20656);
nor U22244 (N_22244,N_20112,N_20752);
nand U22245 (N_22245,N_21129,N_20873);
nor U22246 (N_22246,N_21510,N_20737);
nor U22247 (N_22247,N_21720,N_20437);
nand U22248 (N_22248,N_20952,N_21667);
nand U22249 (N_22249,N_20564,N_20793);
or U22250 (N_22250,N_21220,N_20552);
xnor U22251 (N_22251,N_20024,N_20897);
nand U22252 (N_22252,N_20398,N_21186);
xor U22253 (N_22253,N_21529,N_20292);
xor U22254 (N_22254,N_20536,N_21997);
or U22255 (N_22255,N_21188,N_21933);
or U22256 (N_22256,N_20524,N_20109);
nor U22257 (N_22257,N_20783,N_20987);
or U22258 (N_22258,N_20747,N_21713);
nand U22259 (N_22259,N_20185,N_20691);
nand U22260 (N_22260,N_21701,N_20682);
or U22261 (N_22261,N_21952,N_20425);
or U22262 (N_22262,N_21992,N_21665);
or U22263 (N_22263,N_20898,N_21683);
or U22264 (N_22264,N_20327,N_21381);
xnor U22265 (N_22265,N_20819,N_20289);
nor U22266 (N_22266,N_20730,N_21437);
nor U22267 (N_22267,N_21709,N_21616);
nor U22268 (N_22268,N_21852,N_20671);
nor U22269 (N_22269,N_21101,N_21754);
or U22270 (N_22270,N_21247,N_20727);
nor U22271 (N_22271,N_20116,N_20325);
and U22272 (N_22272,N_21396,N_20237);
xnor U22273 (N_22273,N_20050,N_21660);
nand U22274 (N_22274,N_20178,N_21532);
nor U22275 (N_22275,N_20726,N_21675);
xor U22276 (N_22276,N_20401,N_21365);
and U22277 (N_22277,N_21564,N_20410);
xnor U22278 (N_22278,N_20432,N_20103);
and U22279 (N_22279,N_21423,N_20172);
nand U22280 (N_22280,N_21859,N_21020);
or U22281 (N_22281,N_21030,N_21037);
nor U22282 (N_22282,N_21500,N_20362);
xnor U22283 (N_22283,N_20515,N_20057);
and U22284 (N_22284,N_20491,N_21453);
nand U22285 (N_22285,N_20942,N_21390);
xor U22286 (N_22286,N_20915,N_20729);
nand U22287 (N_22287,N_21882,N_21205);
and U22288 (N_22288,N_20087,N_21737);
or U22289 (N_22289,N_21891,N_20553);
or U22290 (N_22290,N_21799,N_21944);
nand U22291 (N_22291,N_20181,N_21122);
nand U22292 (N_22292,N_20799,N_21029);
nor U22293 (N_22293,N_21553,N_21150);
nand U22294 (N_22294,N_20265,N_20093);
xor U22295 (N_22295,N_20911,N_21955);
or U22296 (N_22296,N_20807,N_21245);
xor U22297 (N_22297,N_20870,N_21926);
xnor U22298 (N_22298,N_21302,N_21568);
or U22299 (N_22299,N_21813,N_21317);
nor U22300 (N_22300,N_21284,N_20743);
xor U22301 (N_22301,N_20528,N_20866);
or U22302 (N_22302,N_20980,N_21454);
and U22303 (N_22303,N_20217,N_21297);
nor U22304 (N_22304,N_21050,N_20048);
or U22305 (N_22305,N_20756,N_21034);
nor U22306 (N_22306,N_21347,N_21674);
nand U22307 (N_22307,N_20532,N_21480);
xnor U22308 (N_22308,N_21348,N_21888);
nor U22309 (N_22309,N_21124,N_21259);
nand U22310 (N_22310,N_21099,N_20232);
and U22311 (N_22311,N_21431,N_20599);
xor U22312 (N_22312,N_21349,N_21931);
xnor U22313 (N_22313,N_20290,N_20101);
nand U22314 (N_22314,N_20646,N_21869);
nor U22315 (N_22315,N_21904,N_20720);
xnor U22316 (N_22316,N_20416,N_21070);
nor U22317 (N_22317,N_20095,N_20476);
nand U22318 (N_22318,N_20074,N_20849);
xor U22319 (N_22319,N_21954,N_20333);
or U22320 (N_22320,N_20205,N_21011);
and U22321 (N_22321,N_20459,N_20768);
nand U22322 (N_22322,N_21028,N_21065);
or U22323 (N_22323,N_21679,N_20653);
nand U22324 (N_22324,N_21800,N_20733);
or U22325 (N_22325,N_21638,N_20628);
nand U22326 (N_22326,N_20749,N_20360);
nor U22327 (N_22327,N_20413,N_21461);
nand U22328 (N_22328,N_20424,N_21729);
or U22329 (N_22329,N_21273,N_21168);
xnor U22330 (N_22330,N_20998,N_21149);
or U22331 (N_22331,N_21427,N_21721);
nor U22332 (N_22332,N_20635,N_21619);
nor U22333 (N_22333,N_21177,N_21582);
or U22334 (N_22334,N_21906,N_21196);
and U22335 (N_22335,N_20198,N_20270);
nor U22336 (N_22336,N_20139,N_21375);
and U22337 (N_22337,N_20571,N_20072);
nor U22338 (N_22338,N_20696,N_20974);
nor U22339 (N_22339,N_21228,N_20623);
and U22340 (N_22340,N_21215,N_20535);
nor U22341 (N_22341,N_21219,N_20667);
nand U22342 (N_22342,N_20666,N_20032);
nand U22343 (N_22343,N_21088,N_20862);
nand U22344 (N_22344,N_20435,N_20326);
nand U22345 (N_22345,N_21182,N_21985);
xnor U22346 (N_22346,N_21403,N_20393);
nor U22347 (N_22347,N_20970,N_20917);
or U22348 (N_22348,N_21512,N_20620);
nand U22349 (N_22349,N_21102,N_21367);
xor U22350 (N_22350,N_21106,N_20368);
or U22351 (N_22351,N_20986,N_20005);
and U22352 (N_22352,N_21825,N_21380);
nand U22353 (N_22353,N_20565,N_20782);
or U22354 (N_22354,N_20930,N_21558);
xor U22355 (N_22355,N_21608,N_20888);
and U22356 (N_22356,N_20438,N_21501);
or U22357 (N_22357,N_21434,N_21187);
nor U22358 (N_22358,N_21504,N_20439);
nor U22359 (N_22359,N_21174,N_21698);
xnor U22360 (N_22360,N_20530,N_20242);
nor U22361 (N_22361,N_20460,N_21871);
nor U22362 (N_22362,N_21213,N_21509);
nor U22363 (N_22363,N_20858,N_21643);
nand U22364 (N_22364,N_21274,N_20255);
nand U22365 (N_22365,N_20597,N_20337);
or U22366 (N_22366,N_21076,N_21913);
and U22367 (N_22367,N_21611,N_20582);
xor U22368 (N_22368,N_20023,N_20276);
or U22369 (N_22369,N_21459,N_21717);
nand U22370 (N_22370,N_21960,N_20227);
or U22371 (N_22371,N_20218,N_20307);
or U22372 (N_22372,N_20527,N_21595);
xor U22373 (N_22373,N_21255,N_20644);
or U22374 (N_22374,N_20221,N_20665);
or U22375 (N_22375,N_21418,N_20254);
nor U22376 (N_22376,N_21991,N_21972);
nand U22377 (N_22377,N_20542,N_21982);
nand U22378 (N_22378,N_20322,N_21335);
nor U22379 (N_22379,N_20248,N_21658);
and U22380 (N_22380,N_20761,N_20312);
nand U22381 (N_22381,N_20455,N_20984);
nand U22382 (N_22382,N_21087,N_20264);
nor U22383 (N_22383,N_21753,N_20643);
nand U22384 (N_22384,N_20728,N_21897);
xor U22385 (N_22385,N_20384,N_21340);
nand U22386 (N_22386,N_20108,N_21345);
nor U22387 (N_22387,N_20850,N_20924);
nor U22388 (N_22388,N_21567,N_20994);
nand U22389 (N_22389,N_20467,N_21989);
and U22390 (N_22390,N_21114,N_21875);
and U22391 (N_22391,N_21468,N_20566);
and U22392 (N_22392,N_21549,N_21025);
xor U22393 (N_22393,N_20305,N_21686);
and U22394 (N_22394,N_20676,N_21704);
nor U22395 (N_22395,N_21814,N_21217);
xor U22396 (N_22396,N_20649,N_20995);
nand U22397 (N_22397,N_21647,N_21134);
or U22398 (N_22398,N_20708,N_20126);
nand U22399 (N_22399,N_20559,N_20966);
or U22400 (N_22400,N_21789,N_20183);
or U22401 (N_22401,N_21181,N_21353);
nor U22402 (N_22402,N_21597,N_21144);
or U22403 (N_22403,N_20245,N_20828);
xor U22404 (N_22404,N_21359,N_21593);
nand U22405 (N_22405,N_21190,N_20177);
xor U22406 (N_22406,N_20259,N_20732);
nor U22407 (N_22407,N_21233,N_21585);
nor U22408 (N_22408,N_20992,N_21295);
xor U22409 (N_22409,N_20938,N_21592);
nand U22410 (N_22410,N_21136,N_20854);
xnor U22411 (N_22411,N_21079,N_21253);
xnor U22412 (N_22412,N_21752,N_20618);
or U22413 (N_22413,N_21559,N_21820);
nor U22414 (N_22414,N_21829,N_20679);
xnor U22415 (N_22415,N_20860,N_20855);
nor U22416 (N_22416,N_21648,N_21422);
nor U22417 (N_22417,N_20981,N_20370);
nor U22418 (N_22418,N_21161,N_20338);
or U22419 (N_22419,N_20027,N_20471);
and U22420 (N_22420,N_20445,N_20507);
or U22421 (N_22421,N_20804,N_21759);
nor U22422 (N_22422,N_21606,N_20256);
and U22423 (N_22423,N_21563,N_20082);
nor U22424 (N_22424,N_20314,N_20394);
and U22425 (N_22425,N_20672,N_21266);
and U22426 (N_22426,N_21002,N_20447);
and U22427 (N_22427,N_20722,N_21425);
and U22428 (N_22428,N_21959,N_21451);
nand U22429 (N_22429,N_20260,N_20071);
or U22430 (N_22430,N_20876,N_20545);
nand U22431 (N_22431,N_21238,N_20088);
nand U22432 (N_22432,N_20417,N_21864);
xnor U22433 (N_22433,N_20704,N_20125);
nand U22434 (N_22434,N_21900,N_20169);
and U22435 (N_22435,N_21793,N_21537);
or U22436 (N_22436,N_21202,N_21162);
or U22437 (N_22437,N_20044,N_20006);
xnor U22438 (N_22438,N_21200,N_20544);
and U22439 (N_22439,N_21081,N_21054);
xnor U22440 (N_22440,N_21350,N_20905);
nor U22441 (N_22441,N_21515,N_21401);
nor U22442 (N_22442,N_20581,N_20686);
nand U22443 (N_22443,N_21042,N_21522);
nor U22444 (N_22444,N_21051,N_20640);
xor U22445 (N_22445,N_21838,N_20431);
and U22446 (N_22446,N_21892,N_21560);
nor U22447 (N_22447,N_20767,N_20706);
xor U22448 (N_22448,N_21967,N_20001);
xnor U22449 (N_22449,N_21916,N_20580);
or U22450 (N_22450,N_21151,N_21979);
nor U22451 (N_22451,N_20814,N_20197);
or U22452 (N_22452,N_20501,N_20607);
nor U22453 (N_22453,N_20346,N_21443);
nor U22454 (N_22454,N_20721,N_20584);
and U22455 (N_22455,N_21180,N_21271);
or U22456 (N_22456,N_20429,N_20962);
and U22457 (N_22457,N_21872,N_20464);
xnor U22458 (N_22458,N_20932,N_21184);
nor U22459 (N_22459,N_21715,N_20774);
or U22460 (N_22460,N_20918,N_20448);
nor U22461 (N_22461,N_21788,N_20687);
or U22462 (N_22462,N_20194,N_21995);
or U22463 (N_22463,N_20388,N_20272);
nand U22464 (N_22464,N_20558,N_20701);
xor U22465 (N_22465,N_21929,N_20579);
and U22466 (N_22466,N_20779,N_20574);
nor U22467 (N_22467,N_21724,N_21330);
or U22468 (N_22468,N_21374,N_21530);
nor U22469 (N_22469,N_21783,N_20120);
nor U22470 (N_22470,N_21222,N_20481);
nor U22471 (N_22471,N_20236,N_20848);
nand U22472 (N_22472,N_20022,N_21705);
nand U22473 (N_22473,N_21409,N_20415);
nand U22474 (N_22474,N_21336,N_20366);
nand U22475 (N_22475,N_20718,N_20763);
nand U22476 (N_22476,N_21324,N_20847);
or U22477 (N_22477,N_21696,N_20662);
nand U22478 (N_22478,N_20810,N_21033);
nor U22479 (N_22479,N_20106,N_20411);
or U22480 (N_22480,N_20820,N_20506);
nand U22481 (N_22481,N_21841,N_20159);
nand U22482 (N_22482,N_21760,N_21671);
xor U22483 (N_22483,N_21901,N_21516);
or U22484 (N_22484,N_21440,N_20592);
nor U22485 (N_22485,N_21682,N_21666);
xor U22486 (N_22486,N_20953,N_21923);
nor U22487 (N_22487,N_21688,N_21550);
nor U22488 (N_22488,N_20442,N_20955);
or U22489 (N_22489,N_20634,N_20806);
xor U22490 (N_22490,N_21482,N_21327);
nand U22491 (N_22491,N_20059,N_20094);
nor U22492 (N_22492,N_20422,N_20977);
nor U22493 (N_22493,N_21576,N_21538);
or U22494 (N_22494,N_20754,N_20047);
xnor U22495 (N_22495,N_20453,N_20816);
nand U22496 (N_22496,N_21903,N_20490);
xor U22497 (N_22497,N_21803,N_21128);
or U22498 (N_22498,N_21154,N_21670);
xor U22499 (N_22499,N_21007,N_20827);
xor U22500 (N_22500,N_21393,N_21046);
nor U22501 (N_22501,N_20606,N_20885);
nand U22502 (N_22502,N_21242,N_21806);
nor U22503 (N_22503,N_20736,N_21942);
xnor U22504 (N_22504,N_20239,N_21152);
and U22505 (N_22505,N_20570,N_21642);
xnor U22506 (N_22506,N_21356,N_20133);
and U22507 (N_22507,N_20735,N_20090);
or U22508 (N_22508,N_20208,N_20061);
or U22509 (N_22509,N_20719,N_21876);
nor U22510 (N_22510,N_20306,N_21001);
nand U22511 (N_22511,N_21399,N_20186);
and U22512 (N_22512,N_20235,N_21436);
nor U22513 (N_22513,N_21159,N_21843);
or U22514 (N_22514,N_20577,N_20449);
nand U22515 (N_22515,N_20427,N_20595);
or U22516 (N_22516,N_20556,N_21283);
or U22517 (N_22517,N_20037,N_20789);
nand U22518 (N_22518,N_20400,N_20978);
nor U22519 (N_22519,N_20119,N_21281);
nor U22520 (N_22520,N_20745,N_21062);
nand U22521 (N_22521,N_21999,N_21639);
and U22522 (N_22522,N_20352,N_21334);
xnor U22523 (N_22523,N_21824,N_21172);
or U22524 (N_22524,N_21481,N_20845);
nor U22525 (N_22525,N_20757,N_20969);
and U22526 (N_22526,N_20578,N_21782);
and U22527 (N_22527,N_20973,N_20990);
nand U22528 (N_22528,N_21212,N_21785);
or U22529 (N_22529,N_21694,N_21056);
nor U22530 (N_22530,N_21907,N_20523);
nor U22531 (N_22531,N_21237,N_21313);
nand U22532 (N_22532,N_20162,N_21276);
nand U22533 (N_22533,N_21662,N_20130);
or U22534 (N_22534,N_20461,N_21524);
nand U22535 (N_22535,N_21321,N_21026);
and U22536 (N_22536,N_20190,N_20703);
or U22537 (N_22537,N_21556,N_21236);
nor U22538 (N_22538,N_21579,N_20351);
and U22539 (N_22539,N_21917,N_20549);
nand U22540 (N_22540,N_20874,N_21421);
or U22541 (N_22541,N_20796,N_20902);
or U22542 (N_22542,N_20358,N_21010);
nor U22543 (N_22543,N_21291,N_20452);
nand U22544 (N_22544,N_20881,N_20138);
nor U22545 (N_22545,N_21669,N_21948);
xor U22546 (N_22546,N_21712,N_21191);
and U22547 (N_22547,N_20851,N_21681);
or U22548 (N_22548,N_21364,N_20308);
and U22549 (N_22549,N_21801,N_20573);
xnor U22550 (N_22550,N_20903,N_21018);
xor U22551 (N_22551,N_20839,N_21092);
nand U22552 (N_22552,N_20299,N_21496);
nand U22553 (N_22553,N_20963,N_21346);
nand U22554 (N_22554,N_21920,N_21111);
nand U22555 (N_22555,N_20891,N_21406);
or U22556 (N_22556,N_21758,N_20030);
xor U22557 (N_22557,N_21311,N_21075);
nor U22558 (N_22558,N_21265,N_21395);
xor U22559 (N_22559,N_21398,N_20750);
xnor U22560 (N_22560,N_20084,N_21924);
xnor U22561 (N_22561,N_21826,N_20229);
and U22562 (N_22562,N_20838,N_21975);
xnor U22563 (N_22563,N_21971,N_20372);
or U22564 (N_22564,N_20463,N_21017);
nor U22565 (N_22565,N_20833,N_21636);
xnor U22566 (N_22566,N_20781,N_20700);
nor U22567 (N_22567,N_20818,N_21668);
nand U22568 (N_22568,N_20939,N_20480);
xor U22569 (N_22569,N_21741,N_21497);
nor U22570 (N_22570,N_20945,N_21498);
and U22571 (N_22571,N_21695,N_20684);
and U22572 (N_22572,N_21911,N_21542);
or U22573 (N_22573,N_21728,N_21895);
nand U22574 (N_22574,N_20934,N_20068);
nand U22575 (N_22575,N_20405,N_21329);
xor U22576 (N_22576,N_21426,N_20975);
or U22577 (N_22577,N_20800,N_21513);
and U22578 (N_22578,N_20758,N_21415);
nor U22579 (N_22579,N_21540,N_20135);
xnor U22580 (N_22580,N_21842,N_20402);
nand U22581 (N_22581,N_21258,N_20598);
or U22582 (N_22582,N_20711,N_20498);
nand U22583 (N_22583,N_20028,N_20007);
or U22584 (N_22584,N_21858,N_20258);
nand U22585 (N_22585,N_20128,N_20692);
nand U22586 (N_22586,N_21331,N_20668);
and U22587 (N_22587,N_20697,N_21630);
or U22588 (N_22588,N_20509,N_20240);
nand U22589 (N_22589,N_21322,N_21653);
and U22590 (N_22590,N_21195,N_20521);
or U22591 (N_22591,N_21464,N_21446);
or U22592 (N_22592,N_21786,N_20853);
or U22593 (N_22593,N_20993,N_21333);
nor U22594 (N_22594,N_20382,N_20146);
nand U22595 (N_22595,N_21808,N_21301);
xor U22596 (N_22596,N_21185,N_21047);
xor U22597 (N_22597,N_20175,N_21163);
xor U22598 (N_22598,N_20551,N_20142);
xnor U22599 (N_22599,N_21620,N_20317);
and U22600 (N_22600,N_20137,N_21956);
nand U22601 (N_22601,N_20794,N_21118);
or U22602 (N_22602,N_20121,N_21103);
xnor U22603 (N_22603,N_20086,N_21577);
nor U22604 (N_22604,N_20296,N_21140);
xnor U22605 (N_22605,N_20514,N_20588);
xor U22606 (N_22606,N_20113,N_20775);
xnor U22607 (N_22607,N_21673,N_21928);
xor U22608 (N_22608,N_20919,N_20674);
or U22609 (N_22609,N_20482,N_20823);
xnor U22610 (N_22610,N_21304,N_20960);
or U22611 (N_22611,N_21472,N_20929);
nand U22612 (N_22612,N_20332,N_21066);
or U22613 (N_22613,N_21358,N_20699);
nor U22614 (N_22614,N_20654,N_21155);
nor U22615 (N_22615,N_21287,N_20705);
nand U22616 (N_22616,N_20941,N_21432);
nor U22617 (N_22617,N_20534,N_21133);
xor U22618 (N_22618,N_20709,N_21672);
nand U22619 (N_22619,N_21844,N_21332);
nor U22620 (N_22620,N_20724,N_21993);
nor U22621 (N_22621,N_20034,N_20857);
or U22622 (N_22622,N_20091,N_20979);
or U22623 (N_22623,N_21494,N_20064);
nand U22624 (N_22624,N_21566,N_21027);
or U22625 (N_22625,N_21747,N_20944);
nor U22626 (N_22626,N_21860,N_20503);
xor U22627 (N_22627,N_20784,N_21708);
and U22628 (N_22628,N_20631,N_20069);
nand U22629 (N_22629,N_20320,N_21751);
nand U22630 (N_22630,N_20583,N_20364);
xnor U22631 (N_22631,N_20844,N_21484);
xnor U22632 (N_22632,N_21833,N_20104);
xnor U22633 (N_22633,N_20213,N_21091);
and U22634 (N_22634,N_21914,N_21565);
xor U22635 (N_22635,N_21562,N_21572);
xnor U22636 (N_22636,N_20446,N_20014);
and U22637 (N_22637,N_20015,N_21950);
xor U22638 (N_22638,N_20092,N_21131);
nand U22639 (N_22639,N_20600,N_21389);
or U22640 (N_22640,N_21588,N_21294);
and U22641 (N_22641,N_20152,N_20685);
and U22642 (N_22642,N_20207,N_20156);
or U22643 (N_22643,N_21544,N_20912);
nor U22644 (N_22644,N_21009,N_21424);
and U22645 (N_22645,N_20922,N_20802);
and U22646 (N_22646,N_20811,N_20561);
xor U22647 (N_22647,N_21173,N_20318);
xor U22648 (N_22648,N_21663,N_20168);
xor U22649 (N_22649,N_20734,N_21039);
xor U22650 (N_22650,N_20746,N_20693);
nor U22651 (N_22651,N_21298,N_20651);
nor U22652 (N_22652,N_20920,N_20632);
xor U22653 (N_22653,N_21442,N_21823);
or U22654 (N_22654,N_21714,N_20067);
nand U22655 (N_22655,N_21257,N_21448);
xnor U22656 (N_22656,N_20279,N_21296);
nor U22657 (N_22657,N_21105,N_21379);
nor U22658 (N_22658,N_21626,N_20968);
xor U22659 (N_22659,N_21006,N_20102);
and U22660 (N_22660,N_21528,N_20714);
nor U22661 (N_22661,N_20825,N_21312);
and U22662 (N_22662,N_21641,N_21306);
xor U22663 (N_22663,N_21123,N_21523);
nor U22664 (N_22664,N_20257,N_21533);
xor U22665 (N_22665,N_21835,N_21419);
and U22666 (N_22666,N_20226,N_21787);
nand U22667 (N_22667,N_21980,N_21467);
and U22668 (N_22668,N_21083,N_20031);
xor U22669 (N_22669,N_20143,N_20829);
or U22670 (N_22670,N_21005,N_20462);
or U22671 (N_22671,N_21640,N_21945);
or U22672 (N_22672,N_20423,N_21053);
or U22673 (N_22673,N_20196,N_20954);
and U22674 (N_22674,N_20020,N_21261);
nor U22675 (N_22675,N_20822,N_20350);
and U22676 (N_22676,N_20716,N_20519);
and U22677 (N_22677,N_21487,N_20153);
nand U22678 (N_22678,N_20608,N_21988);
nand U22679 (N_22679,N_20284,N_20124);
nor U22680 (N_22680,N_20821,N_20817);
or U22681 (N_22681,N_21089,N_20773);
nand U22682 (N_22682,N_21854,N_20058);
xnor U22683 (N_22683,N_20893,N_21981);
xor U22684 (N_22684,N_21470,N_21974);
nor U22685 (N_22685,N_21596,N_20797);
nor U22686 (N_22686,N_20627,N_21503);
nand U22687 (N_22687,N_20335,N_21248);
nand U22688 (N_22688,N_21739,N_21885);
nand U22689 (N_22689,N_21097,N_21545);
or U22690 (N_22690,N_20798,N_20576);
and U22691 (N_22691,N_20033,N_21743);
or U22692 (N_22692,N_21874,N_21910);
and U22693 (N_22693,N_20493,N_21397);
or U22694 (N_22694,N_20339,N_20805);
xnor U22695 (N_22695,N_20688,N_21569);
nor U22696 (N_22696,N_20225,N_20489);
and U22697 (N_22697,N_20434,N_21137);
or U22698 (N_22698,N_20883,N_20010);
and U22699 (N_22699,N_20875,N_20354);
xor U22700 (N_22700,N_20202,N_20345);
nand U22701 (N_22701,N_21475,N_20038);
nand U22702 (N_22702,N_21288,N_20517);
or U22703 (N_22703,N_20154,N_21096);
nor U22704 (N_22704,N_21260,N_20062);
xnor U22705 (N_22705,N_21439,N_20639);
or U22706 (N_22706,N_21623,N_21460);
and U22707 (N_22707,N_21262,N_20557);
and U22708 (N_22708,N_21716,N_20210);
or U22709 (N_22709,N_20899,N_21610);
and U22710 (N_22710,N_20522,N_20012);
and U22711 (N_22711,N_21780,N_20220);
or U22712 (N_22712,N_21953,N_21932);
nand U22713 (N_22713,N_20214,N_21404);
nor U22714 (N_22714,N_20910,N_21493);
xor U22715 (N_22715,N_21624,N_21318);
or U22716 (N_22716,N_20712,N_21719);
nor U22717 (N_22717,N_20713,N_21802);
xnor U22718 (N_22718,N_20243,N_20787);
nand U22719 (N_22719,N_20658,N_20889);
nand U22720 (N_22720,N_21880,N_20457);
nor U22721 (N_22721,N_21889,N_21580);
nor U22722 (N_22722,N_21909,N_21589);
nand U22723 (N_22723,N_20347,N_20451);
xor U22724 (N_22724,N_20546,N_20760);
xor U22725 (N_22725,N_21791,N_20334);
xnor U22726 (N_22726,N_21816,N_21024);
xor U22727 (N_22727,N_21104,N_20375);
or U22728 (N_22728,N_20122,N_20982);
nor U22729 (N_22729,N_21126,N_21615);
nand U22730 (N_22730,N_20602,N_20511);
nand U22731 (N_22731,N_21377,N_21617);
nor U22732 (N_22732,N_21557,N_21700);
xnor U22733 (N_22733,N_21810,N_20879);
nand U22734 (N_22734,N_20831,N_20234);
or U22735 (N_22735,N_21319,N_21699);
xor U22736 (N_22736,N_20901,N_21867);
nor U22737 (N_22737,N_21634,N_21412);
nand U22738 (N_22738,N_21117,N_21649);
xor U22739 (N_22739,N_20755,N_21394);
and U22740 (N_22740,N_20834,N_21963);
nand U22741 (N_22741,N_20707,N_21687);
or U22742 (N_22742,N_21765,N_20195);
and U22743 (N_22743,N_20622,N_20675);
nor U22744 (N_22744,N_20648,N_20604);
or U22745 (N_22745,N_20363,N_21798);
and U22746 (N_22746,N_20134,N_20852);
nand U22747 (N_22747,N_20764,N_20650);
xor U22748 (N_22748,N_21003,N_21517);
xor U22749 (N_22749,N_20099,N_21637);
nor U22750 (N_22750,N_21457,N_21507);
and U22751 (N_22751,N_21086,N_21573);
or U22752 (N_22752,N_20589,N_20450);
xor U22753 (N_22753,N_21449,N_20097);
nor U22754 (N_22754,N_21264,N_21178);
or U22755 (N_22755,N_21241,N_20013);
or U22756 (N_22756,N_20129,N_21139);
and U22757 (N_22757,N_21112,N_20105);
or U22758 (N_22758,N_20040,N_20936);
and U22759 (N_22759,N_21949,N_21607);
nor U22760 (N_22760,N_21194,N_21234);
nor U22761 (N_22761,N_21703,N_21109);
nand U22762 (N_22762,N_20246,N_21463);
nand U22763 (N_22763,N_20526,N_20872);
and U22764 (N_22764,N_21535,N_20626);
and U22765 (N_22765,N_20340,N_20065);
nand U22766 (N_22766,N_20543,N_21511);
nand U22767 (N_22767,N_21773,N_21625);
or U22768 (N_22768,N_21286,N_20191);
xor U22769 (N_22769,N_20132,N_20443);
xnor U22770 (N_22770,N_20555,N_21120);
or U22771 (N_22771,N_21145,N_21857);
xnor U22772 (N_22772,N_21268,N_20395);
nand U22773 (N_22773,N_20624,N_20136);
nor U22774 (N_22774,N_21827,N_20430);
nor U22775 (N_22775,N_21386,N_21189);
nand U22776 (N_22776,N_21502,N_20310);
nand U22777 (N_22777,N_20055,N_20472);
or U22778 (N_22778,N_21937,N_21951);
nand U22779 (N_22779,N_20458,N_21148);
or U22780 (N_22780,N_20140,N_21045);
nor U22781 (N_22781,N_21836,N_21654);
nor U22782 (N_22782,N_20725,N_21337);
nand U22783 (N_22783,N_21868,N_20268);
and U22784 (N_22784,N_20859,N_20456);
and U22785 (N_22785,N_20483,N_20826);
nand U22786 (N_22786,N_20916,N_21068);
or U22787 (N_22787,N_21570,N_20078);
nor U22788 (N_22788,N_20813,N_20211);
and U22789 (N_22789,N_21594,N_21919);
xnor U22790 (N_22790,N_21211,N_20070);
or U22791 (N_22791,N_21084,N_20539);
nor U22792 (N_22792,N_20865,N_20660);
nor U22793 (N_22793,N_20991,N_21613);
or U22794 (N_22794,N_20999,N_21093);
or U22795 (N_22795,N_20738,N_21603);
nor U22796 (N_22796,N_20636,N_21508);
or U22797 (N_22797,N_21602,N_20386);
nor U22798 (N_22798,N_21990,N_21225);
or U22799 (N_22799,N_20996,N_21059);
nand U22800 (N_22800,N_21845,N_20541);
nor U22801 (N_22801,N_20638,N_20399);
and U22802 (N_22802,N_21115,N_20021);
nor U22803 (N_22803,N_20392,N_21244);
and U22804 (N_22804,N_20877,N_20269);
nor U22805 (N_22805,N_21256,N_21067);
xor U22806 (N_22806,N_21310,N_21726);
nand U22807 (N_22807,N_20407,N_20928);
nor U22808 (N_22808,N_21206,N_21697);
xnor U22809 (N_22809,N_20871,N_21438);
or U22810 (N_22810,N_21058,N_21392);
nand U22811 (N_22811,N_20488,N_21169);
nand U22812 (N_22812,N_21527,N_21744);
nand U22813 (N_22813,N_20158,N_20479);
and U22814 (N_22814,N_21775,N_20149);
and U22815 (N_22815,N_21351,N_21521);
and U22816 (N_22816,N_20167,N_21732);
and U22817 (N_22817,N_20935,N_20611);
nor U22818 (N_22818,N_20412,N_21552);
and U22819 (N_22819,N_21031,N_20127);
nand U22820 (N_22820,N_21898,N_21303);
or U22821 (N_22821,N_21371,N_21809);
nand U22822 (N_22822,N_20652,N_21599);
and U22823 (N_22823,N_21121,N_21840);
nand U22824 (N_22824,N_21794,N_21325);
and U22825 (N_22825,N_21796,N_20273);
and U22826 (N_22826,N_21300,N_21941);
or U22827 (N_22827,N_21450,N_21141);
xnor U22828 (N_22828,N_20390,N_20907);
nor U22829 (N_22829,N_21203,N_21408);
nor U22830 (N_22830,N_20200,N_21561);
and U22831 (N_22831,N_21976,N_21370);
xnor U22832 (N_22832,N_21947,N_21008);
or U22833 (N_22833,N_21846,N_21384);
nor U22834 (N_22834,N_20568,N_20529);
or U22835 (N_22835,N_21201,N_21946);
or U22836 (N_22836,N_21986,N_21614);
nand U22837 (N_22837,N_20788,N_20249);
nand U22838 (N_22838,N_20785,N_21138);
nand U22839 (N_22839,N_20182,N_21343);
or U22840 (N_22840,N_20615,N_20937);
and U22841 (N_22841,N_21023,N_20348);
or U22842 (N_22842,N_21250,N_20959);
or U22843 (N_22843,N_20147,N_20216);
and U22844 (N_22844,N_21167,N_20510);
nor U22845 (N_22845,N_21546,N_20100);
or U22846 (N_22846,N_21757,N_21702);
nor U22847 (N_22847,N_21043,N_20224);
or U22848 (N_22848,N_20824,N_21176);
nor U22849 (N_22849,N_21252,N_21135);
and U22850 (N_22850,N_20670,N_21113);
or U22851 (N_22851,N_20790,N_21157);
and U22852 (N_22852,N_21957,N_21383);
xnor U22853 (N_22853,N_20586,N_20487);
and U22854 (N_22854,N_20060,N_20403);
xor U22855 (N_22855,N_20379,N_20315);
and U22856 (N_22856,N_21689,N_21768);
xnor U22857 (N_22857,N_20215,N_20378);
xor U22858 (N_22858,N_20690,N_20803);
nand U22859 (N_22859,N_20377,N_21828);
xnor U22860 (N_22860,N_21243,N_20089);
xnor U22861 (N_22861,N_21015,N_20063);
nor U22862 (N_22862,N_21368,N_21586);
xnor U22863 (N_22863,N_20277,N_21733);
or U22864 (N_22864,N_21430,N_21730);
nor U22865 (N_22865,N_20324,N_21706);
nor U22866 (N_22866,N_21575,N_20560);
nor U22867 (N_22867,N_20808,N_21790);
nor U22868 (N_22868,N_20715,N_20204);
xnor U22869 (N_22869,N_20659,N_20801);
nor U22870 (N_22870,N_21921,N_20371);
or U22871 (N_22871,N_20421,N_20925);
nand U22872 (N_22872,N_20896,N_20516);
xor U22873 (N_22873,N_21908,N_20404);
or U22874 (N_22874,N_20500,N_21420);
xor U22875 (N_22875,N_21584,N_21984);
and U22876 (N_22876,N_20961,N_20206);
and U22877 (N_22877,N_21499,N_21837);
or U22878 (N_22878,N_21964,N_21119);
and U22879 (N_22879,N_20863,N_20882);
xor U22880 (N_22880,N_21680,N_21040);
and U22881 (N_22881,N_20203,N_21495);
xor U22882 (N_22882,N_21221,N_20244);
xnor U22883 (N_22883,N_20361,N_20414);
xor U22884 (N_22884,N_20585,N_20677);
nand U22885 (N_22885,N_21293,N_21961);
and U22886 (N_22886,N_20965,N_20336);
or U22887 (N_22887,N_20180,N_20342);
and U22888 (N_22888,N_21740,N_20000);
or U22889 (N_22889,N_21770,N_21930);
xnor U22890 (N_22890,N_20357,N_21231);
or U22891 (N_22891,N_21073,N_20669);
or U22892 (N_22892,N_20164,N_21998);
and U22893 (N_22893,N_20603,N_21710);
nand U22894 (N_22894,N_21158,N_20835);
xnor U22895 (N_22895,N_20904,N_21143);
or U22896 (N_22896,N_21745,N_21488);
or U22897 (N_22897,N_21514,N_20972);
nor U22898 (N_22898,N_21456,N_20572);
xnor U22899 (N_22899,N_21214,N_20525);
nor U22900 (N_22900,N_20894,N_21492);
or U22901 (N_22901,N_20520,N_21254);
nand U22902 (N_22902,N_21598,N_20742);
or U22903 (N_22903,N_21057,N_21052);
nor U22904 (N_22904,N_20946,N_21308);
nor U22905 (N_22905,N_20017,N_20770);
nor U22906 (N_22906,N_20193,N_20985);
nor U22907 (N_22907,N_21270,N_20115);
nand U22908 (N_22908,N_20927,N_21776);
xor U22909 (N_22909,N_21692,N_21227);
xor U22910 (N_22910,N_20098,N_20303);
nand U22911 (N_22911,N_21226,N_20281);
xnor U22912 (N_22912,N_21866,N_20150);
nand U22913 (N_22913,N_21772,N_20841);
xor U22914 (N_22914,N_21320,N_20085);
and U22915 (N_22915,N_20466,N_21085);
or U22916 (N_22916,N_21417,N_21382);
xnor U22917 (N_22917,N_21230,N_20504);
nor U22918 (N_22918,N_20282,N_21884);
nand U22919 (N_22919,N_20641,N_21627);
or U22920 (N_22920,N_20837,N_20426);
nor U22921 (N_22921,N_21994,N_21749);
and U22922 (N_22922,N_20836,N_20892);
or U22923 (N_22923,N_21100,N_21019);
nor U22924 (N_22924,N_20842,N_21541);
xor U22925 (N_22925,N_21664,N_20261);
nor U22926 (N_22926,N_21781,N_20772);
and U22927 (N_22927,N_21978,N_21210);
xnor U22928 (N_22928,N_20187,N_21305);
nand U22929 (N_22929,N_20610,N_20702);
xnor U22930 (N_22930,N_20408,N_20160);
nor U22931 (N_22931,N_21299,N_20051);
or U22932 (N_22932,N_21633,N_21110);
or U22933 (N_22933,N_20219,N_20016);
nor U22934 (N_22934,N_21676,N_20616);
xnor U22935 (N_22935,N_21061,N_20004);
xor U22936 (N_22936,N_21208,N_20913);
nor U22937 (N_22937,N_20144,N_20151);
nand U22938 (N_22938,N_20989,N_20304);
nor U22939 (N_22939,N_20625,N_20502);
nor U22940 (N_22940,N_21218,N_21767);
or U22941 (N_22941,N_20176,N_21272);
nand U22942 (N_22942,N_20689,N_21856);
nand U22943 (N_22943,N_20148,N_21646);
nand U22944 (N_22944,N_20492,N_21193);
and U22945 (N_22945,N_20056,N_21821);
or U22946 (N_22946,N_20042,N_20419);
nor U22947 (N_22947,N_21290,N_21074);
or U22948 (N_22948,N_21883,N_21199);
xor U22949 (N_22949,N_21618,N_20843);
or U22950 (N_22950,N_21822,N_21014);
xor U22951 (N_22951,N_21555,N_20647);
xnor U22952 (N_22952,N_21108,N_21691);
and U22953 (N_22953,N_20036,N_20594);
nand U22954 (N_22954,N_20957,N_21554);
and U22955 (N_22955,N_21965,N_20661);
nor U22956 (N_22956,N_21447,N_20741);
and U22957 (N_22957,N_20046,N_20698);
nor U22958 (N_22958,N_21831,N_21925);
or U22959 (N_22959,N_20173,N_21429);
nor U22960 (N_22960,N_21077,N_20441);
nand U22961 (N_22961,N_21655,N_21465);
nor U22962 (N_22962,N_20302,N_21224);
nor U22963 (N_22963,N_20163,N_21400);
nor U22964 (N_22964,N_20947,N_21239);
xnor U22965 (N_22965,N_21373,N_21344);
nand U22966 (N_22966,N_21761,N_20683);
xor U22967 (N_22967,N_21489,N_21612);
nor U22968 (N_22968,N_21235,N_21792);
nand U22969 (N_22969,N_20356,N_20886);
xnor U22970 (N_22970,N_21526,N_20003);
nand U22971 (N_22971,N_20861,N_20311);
and U22972 (N_22972,N_20096,N_21289);
nand U22973 (N_22973,N_21693,N_21069);
nand U22974 (N_22974,N_21474,N_21197);
xor U22975 (N_22975,N_21940,N_20494);
and U22976 (N_22976,N_21044,N_21628);
nor U22977 (N_22977,N_21071,N_20391);
or U22978 (N_22978,N_20695,N_21784);
nand U22979 (N_22979,N_21246,N_21165);
xor U22980 (N_22980,N_21847,N_20301);
and U22981 (N_22981,N_21722,N_20778);
or U22982 (N_22982,N_20949,N_21887);
nand U22983 (N_22983,N_20477,N_20740);
or U22984 (N_22984,N_21915,N_21707);
or U22985 (N_22985,N_21156,N_21677);
xor U22986 (N_22986,N_20118,N_21938);
and U22987 (N_22987,N_21326,N_20791);
or U22988 (N_22988,N_20052,N_20505);
xor U22989 (N_22989,N_21483,N_20323);
nand U22990 (N_22990,N_20931,N_20002);
and U22991 (N_22991,N_21411,N_21983);
and U22992 (N_22992,N_20188,N_21094);
xor U22993 (N_22993,N_20376,N_21590);
or U22994 (N_22994,N_21832,N_21164);
nand U22995 (N_22995,N_20267,N_20073);
xnor U22996 (N_22996,N_20550,N_21656);
nor U22997 (N_22997,N_21016,N_21125);
xnor U22998 (N_22998,N_21455,N_20612);
or U22999 (N_22999,N_20678,N_21756);
xnor U23000 (N_23000,N_21237,N_20339);
xor U23001 (N_23001,N_20446,N_20486);
and U23002 (N_23002,N_20350,N_20683);
and U23003 (N_23003,N_21474,N_20750);
and U23004 (N_23004,N_20218,N_21746);
or U23005 (N_23005,N_20535,N_20101);
xnor U23006 (N_23006,N_20414,N_21943);
and U23007 (N_23007,N_20097,N_20868);
or U23008 (N_23008,N_20626,N_21577);
or U23009 (N_23009,N_21979,N_20572);
xnor U23010 (N_23010,N_21780,N_21203);
nand U23011 (N_23011,N_20045,N_20125);
nor U23012 (N_23012,N_21076,N_20688);
or U23013 (N_23013,N_20511,N_20821);
or U23014 (N_23014,N_21910,N_21219);
or U23015 (N_23015,N_21813,N_20581);
and U23016 (N_23016,N_21088,N_20359);
nand U23017 (N_23017,N_21489,N_21773);
nand U23018 (N_23018,N_20840,N_21594);
or U23019 (N_23019,N_21349,N_21517);
xnor U23020 (N_23020,N_20639,N_20435);
nor U23021 (N_23021,N_20311,N_21130);
xnor U23022 (N_23022,N_20750,N_21359);
nand U23023 (N_23023,N_20975,N_20061);
and U23024 (N_23024,N_21948,N_20280);
nor U23025 (N_23025,N_21088,N_20004);
and U23026 (N_23026,N_21341,N_21946);
nor U23027 (N_23027,N_20501,N_20913);
and U23028 (N_23028,N_21493,N_21979);
xor U23029 (N_23029,N_21704,N_20621);
or U23030 (N_23030,N_21893,N_21890);
nor U23031 (N_23031,N_21278,N_20737);
or U23032 (N_23032,N_21637,N_21336);
nand U23033 (N_23033,N_20593,N_20146);
nand U23034 (N_23034,N_20672,N_20475);
nand U23035 (N_23035,N_21578,N_21956);
nor U23036 (N_23036,N_20901,N_21496);
nand U23037 (N_23037,N_21230,N_21959);
xor U23038 (N_23038,N_20393,N_21481);
xnor U23039 (N_23039,N_21396,N_21989);
and U23040 (N_23040,N_21920,N_21107);
xor U23041 (N_23041,N_21634,N_21227);
nand U23042 (N_23042,N_20364,N_20889);
nand U23043 (N_23043,N_21602,N_20713);
nor U23044 (N_23044,N_21054,N_21431);
nor U23045 (N_23045,N_21395,N_21061);
nand U23046 (N_23046,N_20995,N_21452);
or U23047 (N_23047,N_21372,N_20637);
nor U23048 (N_23048,N_20078,N_21251);
and U23049 (N_23049,N_21836,N_20710);
xor U23050 (N_23050,N_21464,N_21745);
nor U23051 (N_23051,N_20067,N_21244);
xnor U23052 (N_23052,N_21031,N_20176);
xnor U23053 (N_23053,N_20551,N_20725);
nand U23054 (N_23054,N_21879,N_21685);
or U23055 (N_23055,N_21840,N_20547);
and U23056 (N_23056,N_21392,N_21911);
nand U23057 (N_23057,N_21752,N_20074);
nand U23058 (N_23058,N_21910,N_21178);
xor U23059 (N_23059,N_21408,N_20643);
or U23060 (N_23060,N_20668,N_21965);
and U23061 (N_23061,N_20249,N_20299);
nor U23062 (N_23062,N_21596,N_20772);
nand U23063 (N_23063,N_21000,N_20520);
and U23064 (N_23064,N_20982,N_21214);
nor U23065 (N_23065,N_20773,N_20047);
nor U23066 (N_23066,N_20385,N_21377);
and U23067 (N_23067,N_21776,N_21482);
nand U23068 (N_23068,N_20373,N_20750);
nor U23069 (N_23069,N_21097,N_21481);
and U23070 (N_23070,N_21874,N_21246);
or U23071 (N_23071,N_21702,N_21484);
nand U23072 (N_23072,N_20765,N_20753);
nor U23073 (N_23073,N_21397,N_21523);
nor U23074 (N_23074,N_21983,N_20915);
xnor U23075 (N_23075,N_21336,N_20703);
nor U23076 (N_23076,N_20324,N_21033);
or U23077 (N_23077,N_20182,N_20483);
or U23078 (N_23078,N_21384,N_21281);
or U23079 (N_23079,N_20369,N_21478);
or U23080 (N_23080,N_20395,N_21743);
nand U23081 (N_23081,N_20294,N_21271);
xor U23082 (N_23082,N_21822,N_20049);
and U23083 (N_23083,N_21914,N_20419);
nor U23084 (N_23084,N_21099,N_21744);
or U23085 (N_23085,N_20119,N_20373);
nor U23086 (N_23086,N_20646,N_20135);
nand U23087 (N_23087,N_21698,N_21603);
xor U23088 (N_23088,N_21381,N_21905);
xnor U23089 (N_23089,N_20188,N_20135);
xnor U23090 (N_23090,N_21476,N_21043);
or U23091 (N_23091,N_21762,N_21766);
xor U23092 (N_23092,N_21015,N_20456);
nand U23093 (N_23093,N_20663,N_20617);
or U23094 (N_23094,N_20777,N_21841);
xor U23095 (N_23095,N_21424,N_20914);
and U23096 (N_23096,N_20891,N_21230);
and U23097 (N_23097,N_20328,N_20175);
or U23098 (N_23098,N_21178,N_21376);
or U23099 (N_23099,N_21808,N_21145);
and U23100 (N_23100,N_20377,N_21482);
nor U23101 (N_23101,N_21531,N_20989);
xnor U23102 (N_23102,N_21885,N_21208);
xnor U23103 (N_23103,N_21179,N_20474);
and U23104 (N_23104,N_21796,N_20598);
or U23105 (N_23105,N_21719,N_20253);
and U23106 (N_23106,N_21782,N_21338);
or U23107 (N_23107,N_21960,N_21566);
or U23108 (N_23108,N_20728,N_21127);
nor U23109 (N_23109,N_21388,N_21134);
and U23110 (N_23110,N_20550,N_20438);
nor U23111 (N_23111,N_20718,N_20775);
or U23112 (N_23112,N_20053,N_20037);
nor U23113 (N_23113,N_20042,N_20861);
nor U23114 (N_23114,N_21442,N_21936);
or U23115 (N_23115,N_21280,N_21164);
and U23116 (N_23116,N_21602,N_21334);
xnor U23117 (N_23117,N_21516,N_20415);
nand U23118 (N_23118,N_21346,N_21022);
xnor U23119 (N_23119,N_21656,N_20349);
nor U23120 (N_23120,N_20878,N_21089);
nor U23121 (N_23121,N_20888,N_21411);
nand U23122 (N_23122,N_21960,N_21287);
nor U23123 (N_23123,N_20901,N_21742);
xnor U23124 (N_23124,N_20323,N_21369);
xor U23125 (N_23125,N_21555,N_20247);
xor U23126 (N_23126,N_21993,N_20866);
xnor U23127 (N_23127,N_20804,N_20378);
or U23128 (N_23128,N_20594,N_21821);
nand U23129 (N_23129,N_21213,N_21715);
nand U23130 (N_23130,N_21704,N_21894);
and U23131 (N_23131,N_21951,N_20834);
and U23132 (N_23132,N_20010,N_21715);
xor U23133 (N_23133,N_21107,N_21401);
and U23134 (N_23134,N_20745,N_20954);
and U23135 (N_23135,N_21468,N_21068);
nand U23136 (N_23136,N_20616,N_21618);
and U23137 (N_23137,N_20454,N_20550);
nand U23138 (N_23138,N_20997,N_21852);
and U23139 (N_23139,N_20791,N_20189);
xor U23140 (N_23140,N_21880,N_21707);
and U23141 (N_23141,N_20189,N_20196);
or U23142 (N_23142,N_20519,N_21957);
nand U23143 (N_23143,N_20317,N_20682);
or U23144 (N_23144,N_20258,N_21792);
xnor U23145 (N_23145,N_21378,N_20983);
or U23146 (N_23146,N_20168,N_21362);
nor U23147 (N_23147,N_21452,N_20633);
and U23148 (N_23148,N_20380,N_20561);
nor U23149 (N_23149,N_20253,N_20519);
or U23150 (N_23150,N_20505,N_20194);
nor U23151 (N_23151,N_20887,N_21927);
nand U23152 (N_23152,N_20431,N_21002);
nor U23153 (N_23153,N_20412,N_20830);
or U23154 (N_23154,N_21699,N_21075);
xor U23155 (N_23155,N_21172,N_21155);
and U23156 (N_23156,N_21099,N_21434);
nand U23157 (N_23157,N_21011,N_21990);
xnor U23158 (N_23158,N_20377,N_20568);
or U23159 (N_23159,N_20321,N_21926);
nand U23160 (N_23160,N_20448,N_20369);
and U23161 (N_23161,N_20026,N_20964);
nor U23162 (N_23162,N_21861,N_20337);
and U23163 (N_23163,N_20336,N_20487);
or U23164 (N_23164,N_21024,N_21080);
or U23165 (N_23165,N_21071,N_21608);
and U23166 (N_23166,N_20301,N_21602);
and U23167 (N_23167,N_20263,N_20933);
nor U23168 (N_23168,N_21719,N_20007);
nor U23169 (N_23169,N_21500,N_20777);
xnor U23170 (N_23170,N_21684,N_20703);
xor U23171 (N_23171,N_21746,N_21445);
and U23172 (N_23172,N_21676,N_20229);
nor U23173 (N_23173,N_20994,N_21369);
and U23174 (N_23174,N_21499,N_20236);
and U23175 (N_23175,N_20744,N_20344);
or U23176 (N_23176,N_20624,N_21549);
xnor U23177 (N_23177,N_20744,N_21144);
or U23178 (N_23178,N_20059,N_21127);
nor U23179 (N_23179,N_21467,N_21762);
nand U23180 (N_23180,N_20135,N_20515);
nor U23181 (N_23181,N_20989,N_21571);
and U23182 (N_23182,N_20223,N_20065);
and U23183 (N_23183,N_21504,N_21757);
and U23184 (N_23184,N_20840,N_21216);
or U23185 (N_23185,N_21860,N_21256);
and U23186 (N_23186,N_20516,N_21924);
or U23187 (N_23187,N_21215,N_20413);
xor U23188 (N_23188,N_20919,N_20948);
and U23189 (N_23189,N_20232,N_20649);
or U23190 (N_23190,N_20004,N_21462);
nor U23191 (N_23191,N_21321,N_21806);
xnor U23192 (N_23192,N_20861,N_20870);
or U23193 (N_23193,N_20678,N_21414);
and U23194 (N_23194,N_21900,N_20758);
xnor U23195 (N_23195,N_20606,N_20303);
xnor U23196 (N_23196,N_21663,N_20843);
nand U23197 (N_23197,N_20246,N_20275);
nor U23198 (N_23198,N_21944,N_21263);
and U23199 (N_23199,N_21288,N_21624);
nor U23200 (N_23200,N_21929,N_21834);
nand U23201 (N_23201,N_20573,N_21529);
nor U23202 (N_23202,N_21217,N_20779);
nor U23203 (N_23203,N_21198,N_20234);
or U23204 (N_23204,N_20491,N_20402);
or U23205 (N_23205,N_21936,N_20927);
xor U23206 (N_23206,N_20195,N_21206);
nand U23207 (N_23207,N_21282,N_21714);
nor U23208 (N_23208,N_20817,N_21453);
or U23209 (N_23209,N_21229,N_20296);
nand U23210 (N_23210,N_21684,N_21557);
nor U23211 (N_23211,N_21137,N_20659);
and U23212 (N_23212,N_21150,N_21554);
nor U23213 (N_23213,N_21554,N_20147);
nor U23214 (N_23214,N_21270,N_21551);
xnor U23215 (N_23215,N_20162,N_21128);
or U23216 (N_23216,N_20963,N_20037);
nor U23217 (N_23217,N_21084,N_21562);
xor U23218 (N_23218,N_21401,N_21907);
or U23219 (N_23219,N_21369,N_20413);
or U23220 (N_23220,N_20816,N_20447);
nand U23221 (N_23221,N_20055,N_20751);
nor U23222 (N_23222,N_20419,N_20816);
xor U23223 (N_23223,N_21855,N_21123);
nand U23224 (N_23224,N_21517,N_20421);
or U23225 (N_23225,N_20736,N_21967);
nor U23226 (N_23226,N_21687,N_21042);
or U23227 (N_23227,N_21919,N_20976);
and U23228 (N_23228,N_21013,N_20927);
xor U23229 (N_23229,N_20244,N_21598);
xnor U23230 (N_23230,N_21959,N_21205);
or U23231 (N_23231,N_20153,N_21676);
xnor U23232 (N_23232,N_21452,N_20863);
or U23233 (N_23233,N_20479,N_21896);
and U23234 (N_23234,N_21081,N_20072);
or U23235 (N_23235,N_20998,N_20000);
nor U23236 (N_23236,N_21845,N_20307);
nand U23237 (N_23237,N_21786,N_20095);
and U23238 (N_23238,N_21080,N_20473);
and U23239 (N_23239,N_21831,N_21365);
or U23240 (N_23240,N_20025,N_20985);
xor U23241 (N_23241,N_20025,N_21972);
nand U23242 (N_23242,N_20293,N_21851);
or U23243 (N_23243,N_21679,N_20225);
and U23244 (N_23244,N_20260,N_21457);
or U23245 (N_23245,N_20404,N_21631);
and U23246 (N_23246,N_20830,N_20526);
or U23247 (N_23247,N_21090,N_20660);
xnor U23248 (N_23248,N_20721,N_20698);
nand U23249 (N_23249,N_20610,N_21875);
xnor U23250 (N_23250,N_20740,N_20523);
xor U23251 (N_23251,N_20355,N_21380);
xnor U23252 (N_23252,N_21169,N_21066);
nand U23253 (N_23253,N_20205,N_21305);
nand U23254 (N_23254,N_20860,N_20719);
xor U23255 (N_23255,N_20843,N_21431);
and U23256 (N_23256,N_20867,N_21494);
xor U23257 (N_23257,N_20556,N_20057);
or U23258 (N_23258,N_21432,N_21814);
nor U23259 (N_23259,N_20703,N_20759);
xor U23260 (N_23260,N_20738,N_20354);
nand U23261 (N_23261,N_21345,N_21532);
xnor U23262 (N_23262,N_20809,N_20883);
nand U23263 (N_23263,N_21407,N_21609);
xor U23264 (N_23264,N_21161,N_20353);
nor U23265 (N_23265,N_21839,N_20278);
nand U23266 (N_23266,N_21565,N_20278);
or U23267 (N_23267,N_20426,N_20716);
nor U23268 (N_23268,N_21649,N_21308);
nor U23269 (N_23269,N_20440,N_21445);
nand U23270 (N_23270,N_20949,N_20908);
nand U23271 (N_23271,N_21770,N_21445);
xor U23272 (N_23272,N_20432,N_21168);
nand U23273 (N_23273,N_20281,N_20445);
xor U23274 (N_23274,N_20813,N_21970);
and U23275 (N_23275,N_20133,N_20379);
and U23276 (N_23276,N_21121,N_20303);
or U23277 (N_23277,N_21778,N_21651);
nor U23278 (N_23278,N_21905,N_20277);
or U23279 (N_23279,N_20723,N_20544);
and U23280 (N_23280,N_20654,N_21388);
nand U23281 (N_23281,N_20566,N_21191);
and U23282 (N_23282,N_20975,N_20467);
xor U23283 (N_23283,N_20932,N_21335);
nor U23284 (N_23284,N_21630,N_20359);
nand U23285 (N_23285,N_21096,N_20242);
or U23286 (N_23286,N_20954,N_20848);
nand U23287 (N_23287,N_21693,N_20430);
xnor U23288 (N_23288,N_20405,N_20238);
nand U23289 (N_23289,N_20699,N_21237);
nor U23290 (N_23290,N_21735,N_20625);
xnor U23291 (N_23291,N_20800,N_21736);
and U23292 (N_23292,N_20466,N_20748);
nor U23293 (N_23293,N_20235,N_21798);
xnor U23294 (N_23294,N_20337,N_21181);
and U23295 (N_23295,N_21822,N_20419);
nor U23296 (N_23296,N_20506,N_21448);
nand U23297 (N_23297,N_21085,N_21645);
or U23298 (N_23298,N_21079,N_21035);
nand U23299 (N_23299,N_21765,N_20807);
xnor U23300 (N_23300,N_21771,N_20622);
and U23301 (N_23301,N_21997,N_21450);
or U23302 (N_23302,N_20337,N_21546);
xor U23303 (N_23303,N_21030,N_20769);
nor U23304 (N_23304,N_20819,N_21267);
nor U23305 (N_23305,N_21126,N_21762);
xnor U23306 (N_23306,N_21867,N_20774);
or U23307 (N_23307,N_21455,N_21809);
and U23308 (N_23308,N_20060,N_20710);
or U23309 (N_23309,N_21814,N_20464);
xnor U23310 (N_23310,N_21336,N_20551);
nor U23311 (N_23311,N_20119,N_20092);
xnor U23312 (N_23312,N_21417,N_21751);
nand U23313 (N_23313,N_20957,N_20266);
or U23314 (N_23314,N_21161,N_21691);
and U23315 (N_23315,N_21397,N_21187);
and U23316 (N_23316,N_21929,N_21931);
xnor U23317 (N_23317,N_20513,N_21544);
nor U23318 (N_23318,N_20509,N_20574);
or U23319 (N_23319,N_20040,N_20653);
xnor U23320 (N_23320,N_21846,N_21865);
nand U23321 (N_23321,N_21633,N_20665);
and U23322 (N_23322,N_21672,N_21428);
xor U23323 (N_23323,N_20443,N_20224);
nor U23324 (N_23324,N_20693,N_21274);
or U23325 (N_23325,N_20837,N_21722);
nand U23326 (N_23326,N_20554,N_21526);
and U23327 (N_23327,N_20792,N_21035);
nand U23328 (N_23328,N_21586,N_20757);
nor U23329 (N_23329,N_20284,N_20096);
and U23330 (N_23330,N_21859,N_20671);
or U23331 (N_23331,N_20174,N_21537);
nand U23332 (N_23332,N_21264,N_20904);
and U23333 (N_23333,N_20448,N_20175);
nand U23334 (N_23334,N_21689,N_21449);
nor U23335 (N_23335,N_21075,N_20858);
nand U23336 (N_23336,N_21715,N_21558);
nor U23337 (N_23337,N_21628,N_21548);
nand U23338 (N_23338,N_21619,N_21067);
and U23339 (N_23339,N_20069,N_21612);
or U23340 (N_23340,N_21050,N_21195);
or U23341 (N_23341,N_21890,N_20497);
and U23342 (N_23342,N_21222,N_20569);
nand U23343 (N_23343,N_21709,N_20809);
or U23344 (N_23344,N_21660,N_21612);
nor U23345 (N_23345,N_21839,N_20497);
xor U23346 (N_23346,N_21041,N_21568);
xor U23347 (N_23347,N_21984,N_21250);
nand U23348 (N_23348,N_21874,N_21575);
xnor U23349 (N_23349,N_21794,N_21436);
nand U23350 (N_23350,N_20549,N_21583);
xnor U23351 (N_23351,N_20242,N_21877);
and U23352 (N_23352,N_21774,N_20785);
xor U23353 (N_23353,N_20149,N_20771);
xnor U23354 (N_23354,N_21882,N_20343);
xnor U23355 (N_23355,N_20714,N_21456);
or U23356 (N_23356,N_21665,N_20692);
or U23357 (N_23357,N_21055,N_20985);
nor U23358 (N_23358,N_21924,N_20854);
xor U23359 (N_23359,N_20755,N_21130);
or U23360 (N_23360,N_20252,N_20249);
nor U23361 (N_23361,N_21560,N_20084);
and U23362 (N_23362,N_20719,N_20991);
nor U23363 (N_23363,N_21832,N_20527);
xnor U23364 (N_23364,N_20526,N_20704);
xor U23365 (N_23365,N_20197,N_21203);
nor U23366 (N_23366,N_21402,N_20265);
nand U23367 (N_23367,N_20459,N_21098);
nand U23368 (N_23368,N_21801,N_20561);
nand U23369 (N_23369,N_20833,N_20831);
xor U23370 (N_23370,N_20071,N_21830);
and U23371 (N_23371,N_21544,N_21968);
nor U23372 (N_23372,N_20067,N_21253);
nand U23373 (N_23373,N_21151,N_20066);
or U23374 (N_23374,N_21054,N_21231);
or U23375 (N_23375,N_21606,N_21191);
nand U23376 (N_23376,N_21164,N_21805);
nand U23377 (N_23377,N_20642,N_21064);
and U23378 (N_23378,N_21245,N_20120);
nand U23379 (N_23379,N_20019,N_21696);
or U23380 (N_23380,N_20223,N_20869);
nand U23381 (N_23381,N_21843,N_21965);
and U23382 (N_23382,N_21594,N_20339);
nor U23383 (N_23383,N_20805,N_20106);
nor U23384 (N_23384,N_20729,N_20609);
nor U23385 (N_23385,N_21663,N_20883);
and U23386 (N_23386,N_21268,N_20576);
or U23387 (N_23387,N_20440,N_20367);
nor U23388 (N_23388,N_21568,N_20876);
or U23389 (N_23389,N_21685,N_21781);
nor U23390 (N_23390,N_20742,N_20116);
and U23391 (N_23391,N_20763,N_21993);
and U23392 (N_23392,N_21831,N_21206);
nand U23393 (N_23393,N_21385,N_21289);
and U23394 (N_23394,N_21905,N_21975);
nand U23395 (N_23395,N_21508,N_21199);
xor U23396 (N_23396,N_21829,N_20899);
xor U23397 (N_23397,N_21387,N_20894);
nand U23398 (N_23398,N_21887,N_20230);
and U23399 (N_23399,N_21939,N_21352);
nor U23400 (N_23400,N_20613,N_21199);
nand U23401 (N_23401,N_20274,N_20937);
nand U23402 (N_23402,N_21688,N_21239);
xnor U23403 (N_23403,N_20630,N_21531);
nand U23404 (N_23404,N_21097,N_21134);
and U23405 (N_23405,N_20090,N_20672);
or U23406 (N_23406,N_20799,N_20667);
xor U23407 (N_23407,N_20418,N_21956);
and U23408 (N_23408,N_21608,N_20852);
nand U23409 (N_23409,N_21551,N_20292);
and U23410 (N_23410,N_20405,N_21832);
nand U23411 (N_23411,N_21650,N_20088);
and U23412 (N_23412,N_21698,N_21324);
nor U23413 (N_23413,N_21206,N_21153);
xnor U23414 (N_23414,N_20876,N_21337);
or U23415 (N_23415,N_20380,N_21173);
xnor U23416 (N_23416,N_21269,N_21942);
and U23417 (N_23417,N_21790,N_20359);
xor U23418 (N_23418,N_21842,N_20885);
nand U23419 (N_23419,N_21122,N_21278);
and U23420 (N_23420,N_21399,N_21262);
nand U23421 (N_23421,N_21417,N_21548);
nor U23422 (N_23422,N_21505,N_21488);
or U23423 (N_23423,N_21798,N_21285);
xor U23424 (N_23424,N_20800,N_21557);
nor U23425 (N_23425,N_20608,N_20011);
nand U23426 (N_23426,N_21552,N_20996);
nand U23427 (N_23427,N_21022,N_20775);
nand U23428 (N_23428,N_20791,N_21898);
or U23429 (N_23429,N_21096,N_21370);
and U23430 (N_23430,N_20368,N_20051);
nand U23431 (N_23431,N_21124,N_21756);
nand U23432 (N_23432,N_21653,N_21862);
and U23433 (N_23433,N_20931,N_21808);
or U23434 (N_23434,N_20848,N_21568);
and U23435 (N_23435,N_21463,N_21384);
or U23436 (N_23436,N_20008,N_21190);
and U23437 (N_23437,N_21659,N_21008);
nor U23438 (N_23438,N_21910,N_20777);
nor U23439 (N_23439,N_21123,N_20197);
and U23440 (N_23440,N_21567,N_20259);
xor U23441 (N_23441,N_21578,N_20043);
and U23442 (N_23442,N_20322,N_21792);
nor U23443 (N_23443,N_21943,N_20588);
nor U23444 (N_23444,N_20699,N_20920);
nor U23445 (N_23445,N_20428,N_21871);
xor U23446 (N_23446,N_21746,N_20244);
and U23447 (N_23447,N_21607,N_21095);
nand U23448 (N_23448,N_20278,N_20348);
nand U23449 (N_23449,N_21133,N_20064);
or U23450 (N_23450,N_21614,N_21050);
and U23451 (N_23451,N_21753,N_21550);
nand U23452 (N_23452,N_20360,N_20774);
nand U23453 (N_23453,N_21761,N_20754);
and U23454 (N_23454,N_21090,N_21859);
or U23455 (N_23455,N_20336,N_20061);
nor U23456 (N_23456,N_21904,N_20325);
nand U23457 (N_23457,N_21703,N_20309);
or U23458 (N_23458,N_21919,N_21552);
nand U23459 (N_23459,N_21403,N_20738);
xnor U23460 (N_23460,N_20449,N_21732);
and U23461 (N_23461,N_20108,N_20180);
nand U23462 (N_23462,N_21569,N_20736);
and U23463 (N_23463,N_20047,N_21717);
nand U23464 (N_23464,N_21089,N_21647);
nand U23465 (N_23465,N_20104,N_20501);
xor U23466 (N_23466,N_20609,N_21247);
nand U23467 (N_23467,N_20143,N_21198);
and U23468 (N_23468,N_21150,N_21692);
nor U23469 (N_23469,N_20198,N_21970);
and U23470 (N_23470,N_21046,N_21838);
nor U23471 (N_23471,N_20087,N_21181);
xor U23472 (N_23472,N_20477,N_20353);
xor U23473 (N_23473,N_20391,N_21896);
or U23474 (N_23474,N_20164,N_21555);
xnor U23475 (N_23475,N_20925,N_21147);
nor U23476 (N_23476,N_21954,N_21412);
nand U23477 (N_23477,N_20803,N_21572);
nor U23478 (N_23478,N_21508,N_21138);
nand U23479 (N_23479,N_21571,N_20386);
nor U23480 (N_23480,N_20104,N_20864);
and U23481 (N_23481,N_20756,N_21476);
xor U23482 (N_23482,N_20234,N_21902);
or U23483 (N_23483,N_20197,N_21441);
or U23484 (N_23484,N_20818,N_21043);
and U23485 (N_23485,N_20325,N_21718);
or U23486 (N_23486,N_20691,N_21494);
xnor U23487 (N_23487,N_20130,N_21825);
and U23488 (N_23488,N_21393,N_20243);
xor U23489 (N_23489,N_20430,N_20271);
xor U23490 (N_23490,N_20789,N_21705);
and U23491 (N_23491,N_20602,N_20397);
or U23492 (N_23492,N_20778,N_20196);
nor U23493 (N_23493,N_21272,N_21600);
xnor U23494 (N_23494,N_21778,N_20405);
xor U23495 (N_23495,N_21382,N_20785);
and U23496 (N_23496,N_20852,N_20232);
or U23497 (N_23497,N_20665,N_20974);
nor U23498 (N_23498,N_20115,N_20596);
and U23499 (N_23499,N_20155,N_20209);
nor U23500 (N_23500,N_21494,N_20671);
nor U23501 (N_23501,N_21487,N_21776);
nor U23502 (N_23502,N_21589,N_21557);
nand U23503 (N_23503,N_21369,N_20953);
xor U23504 (N_23504,N_21599,N_20790);
nand U23505 (N_23505,N_21221,N_20323);
and U23506 (N_23506,N_21422,N_21236);
or U23507 (N_23507,N_20888,N_21634);
nand U23508 (N_23508,N_21614,N_20747);
nor U23509 (N_23509,N_20802,N_20646);
nor U23510 (N_23510,N_20800,N_21974);
or U23511 (N_23511,N_21753,N_21790);
or U23512 (N_23512,N_21783,N_21636);
or U23513 (N_23513,N_20522,N_20084);
nor U23514 (N_23514,N_20004,N_21442);
nand U23515 (N_23515,N_20518,N_20465);
and U23516 (N_23516,N_20594,N_21329);
or U23517 (N_23517,N_20846,N_21665);
nor U23518 (N_23518,N_20447,N_21842);
and U23519 (N_23519,N_20655,N_20148);
nand U23520 (N_23520,N_20737,N_21160);
or U23521 (N_23521,N_20807,N_21335);
or U23522 (N_23522,N_21983,N_20849);
and U23523 (N_23523,N_21550,N_20122);
nor U23524 (N_23524,N_21591,N_20916);
and U23525 (N_23525,N_21875,N_20998);
or U23526 (N_23526,N_21983,N_20029);
nand U23527 (N_23527,N_21940,N_20096);
or U23528 (N_23528,N_20095,N_20377);
nand U23529 (N_23529,N_20699,N_20175);
and U23530 (N_23530,N_20175,N_20010);
and U23531 (N_23531,N_20468,N_21342);
or U23532 (N_23532,N_20151,N_20945);
or U23533 (N_23533,N_20535,N_21273);
or U23534 (N_23534,N_21063,N_20513);
nand U23535 (N_23535,N_20723,N_21891);
nand U23536 (N_23536,N_20038,N_20093);
nor U23537 (N_23537,N_21515,N_20662);
and U23538 (N_23538,N_20571,N_21061);
nor U23539 (N_23539,N_21351,N_21573);
or U23540 (N_23540,N_20301,N_21208);
xor U23541 (N_23541,N_20156,N_20801);
or U23542 (N_23542,N_20715,N_21006);
nor U23543 (N_23543,N_21429,N_20418);
and U23544 (N_23544,N_21314,N_20403);
nor U23545 (N_23545,N_20715,N_20401);
or U23546 (N_23546,N_20981,N_21525);
and U23547 (N_23547,N_21526,N_21918);
and U23548 (N_23548,N_20412,N_21566);
xnor U23549 (N_23549,N_21768,N_20683);
and U23550 (N_23550,N_20406,N_21470);
xor U23551 (N_23551,N_20565,N_20614);
or U23552 (N_23552,N_21942,N_21247);
xor U23553 (N_23553,N_20310,N_21808);
or U23554 (N_23554,N_20319,N_20226);
xnor U23555 (N_23555,N_21561,N_21471);
or U23556 (N_23556,N_20590,N_20736);
nand U23557 (N_23557,N_20279,N_20261);
and U23558 (N_23558,N_21699,N_21576);
xor U23559 (N_23559,N_20804,N_21926);
xor U23560 (N_23560,N_20130,N_20366);
and U23561 (N_23561,N_21152,N_21759);
xnor U23562 (N_23562,N_20818,N_21817);
xor U23563 (N_23563,N_21704,N_21473);
or U23564 (N_23564,N_21512,N_21158);
nor U23565 (N_23565,N_21550,N_21714);
xor U23566 (N_23566,N_20450,N_20824);
nor U23567 (N_23567,N_21501,N_21778);
nor U23568 (N_23568,N_21414,N_21888);
nor U23569 (N_23569,N_20108,N_20722);
xnor U23570 (N_23570,N_21863,N_20878);
nor U23571 (N_23571,N_21564,N_20165);
xor U23572 (N_23572,N_21494,N_21355);
and U23573 (N_23573,N_20673,N_20011);
nor U23574 (N_23574,N_21989,N_20312);
nand U23575 (N_23575,N_21677,N_21665);
nand U23576 (N_23576,N_21226,N_20903);
nor U23577 (N_23577,N_21330,N_21769);
nand U23578 (N_23578,N_20051,N_21791);
nand U23579 (N_23579,N_21929,N_21609);
nand U23580 (N_23580,N_20237,N_21742);
nand U23581 (N_23581,N_21530,N_21228);
or U23582 (N_23582,N_21863,N_21867);
nand U23583 (N_23583,N_21135,N_20219);
and U23584 (N_23584,N_20082,N_21321);
nand U23585 (N_23585,N_20841,N_20593);
and U23586 (N_23586,N_20917,N_21525);
and U23587 (N_23587,N_20525,N_21376);
xor U23588 (N_23588,N_21214,N_21795);
nor U23589 (N_23589,N_21291,N_20306);
xor U23590 (N_23590,N_21325,N_20772);
nand U23591 (N_23591,N_21227,N_21192);
xnor U23592 (N_23592,N_20767,N_21681);
xor U23593 (N_23593,N_20243,N_20632);
and U23594 (N_23594,N_20961,N_20157);
xor U23595 (N_23595,N_21656,N_21589);
xor U23596 (N_23596,N_21878,N_21203);
nor U23597 (N_23597,N_20630,N_20489);
or U23598 (N_23598,N_20710,N_21460);
xor U23599 (N_23599,N_21788,N_21662);
nand U23600 (N_23600,N_21285,N_21385);
xnor U23601 (N_23601,N_21939,N_20953);
nor U23602 (N_23602,N_21890,N_20272);
or U23603 (N_23603,N_21573,N_21164);
or U23604 (N_23604,N_21748,N_20330);
nor U23605 (N_23605,N_21450,N_20878);
nand U23606 (N_23606,N_20203,N_21652);
xor U23607 (N_23607,N_20029,N_21080);
or U23608 (N_23608,N_20883,N_21570);
xnor U23609 (N_23609,N_20574,N_21545);
or U23610 (N_23610,N_21936,N_21892);
and U23611 (N_23611,N_21830,N_21163);
and U23612 (N_23612,N_21644,N_20413);
nor U23613 (N_23613,N_20433,N_20575);
nand U23614 (N_23614,N_20045,N_21200);
nor U23615 (N_23615,N_21693,N_21808);
and U23616 (N_23616,N_20554,N_20567);
nor U23617 (N_23617,N_21055,N_21954);
nor U23618 (N_23618,N_20137,N_21067);
nand U23619 (N_23619,N_21756,N_20053);
xnor U23620 (N_23620,N_21348,N_20189);
nor U23621 (N_23621,N_21523,N_20366);
or U23622 (N_23622,N_21416,N_21649);
and U23623 (N_23623,N_21837,N_21030);
nand U23624 (N_23624,N_20139,N_21204);
nand U23625 (N_23625,N_20108,N_21630);
xor U23626 (N_23626,N_20778,N_20475);
nand U23627 (N_23627,N_20431,N_21452);
xor U23628 (N_23628,N_20496,N_20588);
or U23629 (N_23629,N_20591,N_20864);
or U23630 (N_23630,N_21891,N_20834);
nor U23631 (N_23631,N_20172,N_21394);
nand U23632 (N_23632,N_21750,N_21111);
or U23633 (N_23633,N_21780,N_20820);
and U23634 (N_23634,N_20588,N_20011);
xor U23635 (N_23635,N_20503,N_20323);
xor U23636 (N_23636,N_21344,N_20379);
or U23637 (N_23637,N_21128,N_21870);
nor U23638 (N_23638,N_21919,N_20405);
xor U23639 (N_23639,N_20853,N_20696);
and U23640 (N_23640,N_20657,N_21807);
or U23641 (N_23641,N_20108,N_20777);
xnor U23642 (N_23642,N_21240,N_20965);
xnor U23643 (N_23643,N_21499,N_21040);
and U23644 (N_23644,N_20669,N_21165);
xnor U23645 (N_23645,N_20399,N_21147);
xnor U23646 (N_23646,N_20587,N_21952);
and U23647 (N_23647,N_21517,N_21275);
nor U23648 (N_23648,N_21821,N_21278);
or U23649 (N_23649,N_20694,N_21824);
and U23650 (N_23650,N_20577,N_21143);
or U23651 (N_23651,N_20738,N_21656);
nor U23652 (N_23652,N_21214,N_20885);
nand U23653 (N_23653,N_20574,N_21369);
nand U23654 (N_23654,N_20448,N_21521);
and U23655 (N_23655,N_21923,N_20269);
nor U23656 (N_23656,N_21499,N_21244);
xnor U23657 (N_23657,N_21096,N_21611);
or U23658 (N_23658,N_21055,N_21181);
and U23659 (N_23659,N_20993,N_20557);
or U23660 (N_23660,N_21990,N_20600);
or U23661 (N_23661,N_20440,N_20396);
nand U23662 (N_23662,N_21513,N_21877);
nor U23663 (N_23663,N_20061,N_20111);
and U23664 (N_23664,N_21413,N_21005);
nor U23665 (N_23665,N_21776,N_20812);
or U23666 (N_23666,N_21515,N_20515);
or U23667 (N_23667,N_21254,N_21546);
xor U23668 (N_23668,N_21378,N_21411);
and U23669 (N_23669,N_20396,N_20106);
nor U23670 (N_23670,N_21458,N_20278);
or U23671 (N_23671,N_21608,N_21754);
xor U23672 (N_23672,N_20806,N_21316);
nand U23673 (N_23673,N_21522,N_20234);
and U23674 (N_23674,N_21008,N_21629);
nor U23675 (N_23675,N_21105,N_21111);
and U23676 (N_23676,N_21950,N_20103);
nand U23677 (N_23677,N_20328,N_21921);
nor U23678 (N_23678,N_21493,N_20731);
or U23679 (N_23679,N_20929,N_20809);
and U23680 (N_23680,N_21222,N_20301);
or U23681 (N_23681,N_21644,N_20817);
and U23682 (N_23682,N_20372,N_21285);
nor U23683 (N_23683,N_20187,N_20667);
and U23684 (N_23684,N_21605,N_21091);
xor U23685 (N_23685,N_21755,N_20202);
and U23686 (N_23686,N_21929,N_21829);
xnor U23687 (N_23687,N_20675,N_21699);
and U23688 (N_23688,N_21645,N_21204);
nor U23689 (N_23689,N_21069,N_20617);
and U23690 (N_23690,N_21305,N_20553);
xor U23691 (N_23691,N_20602,N_21127);
and U23692 (N_23692,N_21365,N_20033);
nand U23693 (N_23693,N_21656,N_21037);
nand U23694 (N_23694,N_21470,N_21796);
or U23695 (N_23695,N_20138,N_20363);
or U23696 (N_23696,N_21245,N_20982);
xor U23697 (N_23697,N_20731,N_21502);
xnor U23698 (N_23698,N_20823,N_21377);
xor U23699 (N_23699,N_21037,N_21520);
nand U23700 (N_23700,N_21243,N_20564);
xnor U23701 (N_23701,N_20729,N_21550);
or U23702 (N_23702,N_20773,N_20096);
xor U23703 (N_23703,N_21958,N_20991);
or U23704 (N_23704,N_21236,N_20276);
nand U23705 (N_23705,N_21551,N_21471);
nor U23706 (N_23706,N_20672,N_20072);
or U23707 (N_23707,N_21783,N_21859);
nor U23708 (N_23708,N_20525,N_21952);
or U23709 (N_23709,N_20432,N_21237);
nor U23710 (N_23710,N_21796,N_21711);
xnor U23711 (N_23711,N_21255,N_21048);
xor U23712 (N_23712,N_20334,N_21655);
nand U23713 (N_23713,N_21337,N_20028);
or U23714 (N_23714,N_20600,N_20662);
nand U23715 (N_23715,N_20012,N_21033);
xnor U23716 (N_23716,N_20834,N_21506);
nor U23717 (N_23717,N_20075,N_20616);
xor U23718 (N_23718,N_21463,N_21487);
nand U23719 (N_23719,N_20154,N_20275);
and U23720 (N_23720,N_20487,N_21779);
or U23721 (N_23721,N_21144,N_21548);
nand U23722 (N_23722,N_21144,N_20945);
nor U23723 (N_23723,N_20947,N_21523);
xor U23724 (N_23724,N_21911,N_20421);
nor U23725 (N_23725,N_20574,N_20576);
or U23726 (N_23726,N_20387,N_20224);
nor U23727 (N_23727,N_21849,N_20092);
nand U23728 (N_23728,N_21812,N_20834);
or U23729 (N_23729,N_21377,N_20464);
nor U23730 (N_23730,N_21885,N_21757);
nand U23731 (N_23731,N_21891,N_20238);
or U23732 (N_23732,N_20846,N_20724);
nor U23733 (N_23733,N_20155,N_20220);
nand U23734 (N_23734,N_21279,N_20936);
or U23735 (N_23735,N_21577,N_21052);
and U23736 (N_23736,N_21122,N_21901);
nor U23737 (N_23737,N_20571,N_21120);
nor U23738 (N_23738,N_21461,N_21746);
and U23739 (N_23739,N_21228,N_21639);
nand U23740 (N_23740,N_20947,N_20599);
nand U23741 (N_23741,N_20261,N_20636);
nor U23742 (N_23742,N_21000,N_20135);
and U23743 (N_23743,N_20195,N_21126);
and U23744 (N_23744,N_21417,N_21491);
or U23745 (N_23745,N_20328,N_21854);
nand U23746 (N_23746,N_20824,N_21490);
nand U23747 (N_23747,N_21094,N_20290);
or U23748 (N_23748,N_21348,N_21602);
or U23749 (N_23749,N_20976,N_21963);
or U23750 (N_23750,N_20849,N_21676);
and U23751 (N_23751,N_20271,N_20824);
nand U23752 (N_23752,N_21544,N_21019);
xor U23753 (N_23753,N_21285,N_20302);
nand U23754 (N_23754,N_20222,N_21101);
xnor U23755 (N_23755,N_20059,N_20738);
xnor U23756 (N_23756,N_21690,N_20693);
xnor U23757 (N_23757,N_20676,N_20086);
nor U23758 (N_23758,N_20082,N_20458);
nand U23759 (N_23759,N_20059,N_21750);
xnor U23760 (N_23760,N_21830,N_20025);
nor U23761 (N_23761,N_20712,N_21277);
xnor U23762 (N_23762,N_20944,N_21663);
and U23763 (N_23763,N_20126,N_21379);
xnor U23764 (N_23764,N_20701,N_20714);
xor U23765 (N_23765,N_21593,N_21836);
nand U23766 (N_23766,N_20285,N_20964);
xor U23767 (N_23767,N_21869,N_21380);
and U23768 (N_23768,N_21292,N_20294);
nand U23769 (N_23769,N_20566,N_20198);
nor U23770 (N_23770,N_21685,N_21065);
xor U23771 (N_23771,N_20634,N_20847);
and U23772 (N_23772,N_21651,N_21460);
or U23773 (N_23773,N_20266,N_20889);
xnor U23774 (N_23774,N_21173,N_20761);
and U23775 (N_23775,N_20296,N_20799);
and U23776 (N_23776,N_21947,N_20865);
and U23777 (N_23777,N_21000,N_21724);
and U23778 (N_23778,N_20480,N_21770);
or U23779 (N_23779,N_20314,N_21252);
nor U23780 (N_23780,N_21810,N_21806);
and U23781 (N_23781,N_20367,N_21482);
xnor U23782 (N_23782,N_20080,N_21865);
nor U23783 (N_23783,N_21376,N_20061);
nand U23784 (N_23784,N_21381,N_21174);
nand U23785 (N_23785,N_20695,N_20100);
nor U23786 (N_23786,N_20305,N_21413);
xnor U23787 (N_23787,N_21570,N_21017);
xnor U23788 (N_23788,N_20241,N_20617);
nand U23789 (N_23789,N_20439,N_20929);
xor U23790 (N_23790,N_21560,N_20927);
or U23791 (N_23791,N_21195,N_21915);
xor U23792 (N_23792,N_20951,N_21690);
xnor U23793 (N_23793,N_21350,N_21314);
nand U23794 (N_23794,N_21550,N_20865);
xor U23795 (N_23795,N_20362,N_21793);
nand U23796 (N_23796,N_20176,N_20795);
xnor U23797 (N_23797,N_21266,N_20401);
xnor U23798 (N_23798,N_21754,N_20365);
or U23799 (N_23799,N_20211,N_21651);
xor U23800 (N_23800,N_20691,N_20647);
nor U23801 (N_23801,N_20940,N_20506);
nand U23802 (N_23802,N_20182,N_21055);
or U23803 (N_23803,N_21263,N_21690);
nor U23804 (N_23804,N_20988,N_20980);
nand U23805 (N_23805,N_20047,N_20538);
xnor U23806 (N_23806,N_21738,N_21165);
xor U23807 (N_23807,N_21223,N_21686);
nor U23808 (N_23808,N_20975,N_21644);
nor U23809 (N_23809,N_20201,N_21432);
and U23810 (N_23810,N_21122,N_20067);
xor U23811 (N_23811,N_20989,N_21070);
and U23812 (N_23812,N_21787,N_21062);
and U23813 (N_23813,N_21247,N_20418);
or U23814 (N_23814,N_21284,N_21423);
and U23815 (N_23815,N_21419,N_21567);
or U23816 (N_23816,N_20326,N_20194);
xor U23817 (N_23817,N_21648,N_21763);
nor U23818 (N_23818,N_20333,N_21059);
xor U23819 (N_23819,N_20357,N_20942);
nor U23820 (N_23820,N_21757,N_21607);
xnor U23821 (N_23821,N_21342,N_21036);
and U23822 (N_23822,N_21803,N_21138);
xor U23823 (N_23823,N_20828,N_21170);
nand U23824 (N_23824,N_21407,N_21592);
and U23825 (N_23825,N_20782,N_21950);
or U23826 (N_23826,N_21821,N_21042);
and U23827 (N_23827,N_21645,N_20655);
xor U23828 (N_23828,N_20668,N_20155);
xor U23829 (N_23829,N_21397,N_20913);
nor U23830 (N_23830,N_20879,N_20361);
or U23831 (N_23831,N_20079,N_20015);
nor U23832 (N_23832,N_21264,N_21695);
nor U23833 (N_23833,N_21024,N_20058);
xor U23834 (N_23834,N_21352,N_21250);
nand U23835 (N_23835,N_21347,N_20499);
xnor U23836 (N_23836,N_21600,N_20512);
xor U23837 (N_23837,N_20659,N_21213);
nor U23838 (N_23838,N_20846,N_20977);
nand U23839 (N_23839,N_20261,N_20413);
and U23840 (N_23840,N_21348,N_20761);
or U23841 (N_23841,N_20118,N_21611);
nor U23842 (N_23842,N_21554,N_21673);
nor U23843 (N_23843,N_21097,N_20779);
nor U23844 (N_23844,N_20039,N_21259);
xor U23845 (N_23845,N_20384,N_20462);
or U23846 (N_23846,N_21102,N_20083);
and U23847 (N_23847,N_21527,N_20495);
or U23848 (N_23848,N_21975,N_20696);
or U23849 (N_23849,N_21407,N_21539);
nor U23850 (N_23850,N_20990,N_20701);
or U23851 (N_23851,N_20848,N_20019);
xnor U23852 (N_23852,N_21242,N_20914);
xnor U23853 (N_23853,N_21081,N_20762);
and U23854 (N_23854,N_20592,N_21581);
nand U23855 (N_23855,N_21624,N_20140);
xor U23856 (N_23856,N_21027,N_21492);
or U23857 (N_23857,N_20354,N_20852);
and U23858 (N_23858,N_20303,N_20286);
nand U23859 (N_23859,N_20371,N_20298);
nand U23860 (N_23860,N_20069,N_20346);
or U23861 (N_23861,N_21288,N_21762);
nand U23862 (N_23862,N_20177,N_20266);
nand U23863 (N_23863,N_20841,N_20993);
nand U23864 (N_23864,N_20982,N_21394);
nand U23865 (N_23865,N_20692,N_20099);
nor U23866 (N_23866,N_21948,N_21001);
or U23867 (N_23867,N_20252,N_20358);
and U23868 (N_23868,N_21207,N_21310);
and U23869 (N_23869,N_21538,N_21680);
xor U23870 (N_23870,N_20827,N_20622);
nor U23871 (N_23871,N_21641,N_20918);
or U23872 (N_23872,N_20276,N_20649);
nor U23873 (N_23873,N_20250,N_21310);
xor U23874 (N_23874,N_21223,N_21716);
nand U23875 (N_23875,N_20934,N_20026);
nor U23876 (N_23876,N_21175,N_21369);
nor U23877 (N_23877,N_20424,N_21278);
xnor U23878 (N_23878,N_21759,N_20379);
or U23879 (N_23879,N_20879,N_21123);
nor U23880 (N_23880,N_20766,N_20808);
or U23881 (N_23881,N_21802,N_20630);
nand U23882 (N_23882,N_20020,N_21906);
nand U23883 (N_23883,N_20217,N_20288);
nor U23884 (N_23884,N_20375,N_21023);
or U23885 (N_23885,N_21248,N_20846);
nand U23886 (N_23886,N_20326,N_21143);
and U23887 (N_23887,N_20646,N_20250);
nor U23888 (N_23888,N_20037,N_21191);
and U23889 (N_23889,N_21863,N_21662);
and U23890 (N_23890,N_21345,N_21303);
xnor U23891 (N_23891,N_20169,N_21105);
nor U23892 (N_23892,N_20206,N_20769);
xnor U23893 (N_23893,N_20553,N_20307);
xnor U23894 (N_23894,N_21647,N_21171);
and U23895 (N_23895,N_20326,N_20141);
nor U23896 (N_23896,N_21465,N_21601);
nand U23897 (N_23897,N_21002,N_20353);
xor U23898 (N_23898,N_21501,N_21369);
nand U23899 (N_23899,N_21781,N_20083);
nor U23900 (N_23900,N_20393,N_21823);
xor U23901 (N_23901,N_21905,N_21623);
xor U23902 (N_23902,N_20158,N_20598);
or U23903 (N_23903,N_20838,N_20723);
nor U23904 (N_23904,N_21787,N_20158);
xor U23905 (N_23905,N_20211,N_21367);
xor U23906 (N_23906,N_20899,N_21754);
nand U23907 (N_23907,N_21970,N_21784);
and U23908 (N_23908,N_20070,N_20124);
xor U23909 (N_23909,N_20085,N_21368);
nand U23910 (N_23910,N_20305,N_21308);
or U23911 (N_23911,N_20766,N_20825);
nand U23912 (N_23912,N_20681,N_21675);
nor U23913 (N_23913,N_20269,N_20326);
and U23914 (N_23914,N_20317,N_21851);
nor U23915 (N_23915,N_21913,N_20483);
and U23916 (N_23916,N_21990,N_20678);
or U23917 (N_23917,N_20953,N_20852);
xnor U23918 (N_23918,N_21695,N_20673);
xnor U23919 (N_23919,N_20528,N_21709);
xnor U23920 (N_23920,N_21189,N_20445);
xor U23921 (N_23921,N_20272,N_21469);
nor U23922 (N_23922,N_21955,N_21253);
and U23923 (N_23923,N_21189,N_20656);
nand U23924 (N_23924,N_21108,N_20582);
and U23925 (N_23925,N_21032,N_20572);
nor U23926 (N_23926,N_21252,N_21112);
nor U23927 (N_23927,N_20838,N_20560);
xnor U23928 (N_23928,N_21350,N_20939);
and U23929 (N_23929,N_21168,N_20606);
nand U23930 (N_23930,N_21270,N_20740);
xor U23931 (N_23931,N_21189,N_20123);
nor U23932 (N_23932,N_20180,N_20177);
xnor U23933 (N_23933,N_21116,N_21149);
xor U23934 (N_23934,N_20767,N_21162);
nor U23935 (N_23935,N_21417,N_20995);
nor U23936 (N_23936,N_21039,N_20888);
xnor U23937 (N_23937,N_21471,N_20313);
nor U23938 (N_23938,N_21663,N_21476);
or U23939 (N_23939,N_20527,N_20851);
xnor U23940 (N_23940,N_21793,N_20276);
xnor U23941 (N_23941,N_20057,N_20153);
nor U23942 (N_23942,N_20087,N_21784);
xnor U23943 (N_23943,N_20816,N_20294);
nor U23944 (N_23944,N_21811,N_21256);
and U23945 (N_23945,N_21161,N_21841);
nand U23946 (N_23946,N_21051,N_20139);
nand U23947 (N_23947,N_20653,N_20094);
nand U23948 (N_23948,N_21120,N_20520);
nand U23949 (N_23949,N_20937,N_21596);
nand U23950 (N_23950,N_21813,N_20181);
and U23951 (N_23951,N_21129,N_20601);
nand U23952 (N_23952,N_21891,N_21031);
or U23953 (N_23953,N_20631,N_21533);
or U23954 (N_23954,N_20273,N_20758);
nor U23955 (N_23955,N_21777,N_20424);
and U23956 (N_23956,N_21620,N_21137);
and U23957 (N_23957,N_21913,N_21711);
xnor U23958 (N_23958,N_21552,N_21180);
nand U23959 (N_23959,N_21698,N_21397);
nand U23960 (N_23960,N_20707,N_20570);
or U23961 (N_23961,N_20660,N_20185);
nor U23962 (N_23962,N_20045,N_21938);
xor U23963 (N_23963,N_21915,N_21037);
and U23964 (N_23964,N_20757,N_21749);
xnor U23965 (N_23965,N_20889,N_21414);
or U23966 (N_23966,N_20121,N_20443);
and U23967 (N_23967,N_20544,N_21147);
xor U23968 (N_23968,N_21016,N_20454);
and U23969 (N_23969,N_21723,N_21555);
xnor U23970 (N_23970,N_21797,N_21882);
xor U23971 (N_23971,N_20191,N_21892);
nor U23972 (N_23972,N_20596,N_21170);
and U23973 (N_23973,N_21002,N_20595);
xnor U23974 (N_23974,N_20777,N_21331);
or U23975 (N_23975,N_21300,N_21627);
and U23976 (N_23976,N_20440,N_20959);
or U23977 (N_23977,N_20488,N_21801);
or U23978 (N_23978,N_21798,N_21247);
xor U23979 (N_23979,N_21875,N_20928);
and U23980 (N_23980,N_20679,N_20298);
nor U23981 (N_23981,N_21574,N_20822);
nor U23982 (N_23982,N_21912,N_20746);
xnor U23983 (N_23983,N_20789,N_21065);
and U23984 (N_23984,N_20726,N_20931);
nor U23985 (N_23985,N_20788,N_20040);
nand U23986 (N_23986,N_20726,N_20267);
nand U23987 (N_23987,N_20460,N_20437);
nor U23988 (N_23988,N_21465,N_20837);
nand U23989 (N_23989,N_20484,N_20133);
and U23990 (N_23990,N_21300,N_21089);
or U23991 (N_23991,N_20008,N_21538);
xnor U23992 (N_23992,N_21685,N_20637);
and U23993 (N_23993,N_20395,N_20343);
xor U23994 (N_23994,N_21481,N_20225);
or U23995 (N_23995,N_20521,N_20948);
nor U23996 (N_23996,N_21004,N_20399);
nand U23997 (N_23997,N_21842,N_20442);
nand U23998 (N_23998,N_20723,N_20926);
xnor U23999 (N_23999,N_21230,N_20780);
or U24000 (N_24000,N_23234,N_23332);
nand U24001 (N_24001,N_23006,N_22735);
xor U24002 (N_24002,N_22853,N_23787);
or U24003 (N_24003,N_23430,N_22712);
and U24004 (N_24004,N_22102,N_22017);
xor U24005 (N_24005,N_22773,N_22750);
nor U24006 (N_24006,N_23194,N_23185);
or U24007 (N_24007,N_22622,N_23607);
nand U24008 (N_24008,N_22364,N_22611);
nand U24009 (N_24009,N_23986,N_23034);
xor U24010 (N_24010,N_23456,N_22020);
and U24011 (N_24011,N_23484,N_22846);
nor U24012 (N_24012,N_23261,N_23151);
xor U24013 (N_24013,N_22659,N_23934);
and U24014 (N_24014,N_23167,N_22461);
nand U24015 (N_24015,N_23641,N_23520);
xor U24016 (N_24016,N_23842,N_22627);
nor U24017 (N_24017,N_23319,N_23681);
nand U24018 (N_24018,N_22935,N_22673);
nor U24019 (N_24019,N_22909,N_22711);
or U24020 (N_24020,N_23438,N_22862);
xor U24021 (N_24021,N_23535,N_22011);
nand U24022 (N_24022,N_23246,N_22744);
or U24023 (N_24023,N_23798,N_23147);
nor U24024 (N_24024,N_22174,N_23389);
or U24025 (N_24025,N_23577,N_23997);
xor U24026 (N_24026,N_22021,N_22388);
nor U24027 (N_24027,N_23058,N_23476);
nand U24028 (N_24028,N_22427,N_22974);
and U24029 (N_24029,N_23932,N_22459);
nand U24030 (N_24030,N_23971,N_23875);
xnor U24031 (N_24031,N_23470,N_22262);
nand U24032 (N_24032,N_22182,N_23411);
or U24033 (N_24033,N_23899,N_22572);
and U24034 (N_24034,N_23214,N_23047);
or U24035 (N_24035,N_23462,N_23418);
nand U24036 (N_24036,N_22514,N_22534);
xnor U24037 (N_24037,N_23104,N_22844);
or U24038 (N_24038,N_22050,N_23489);
or U24039 (N_24039,N_23368,N_23890);
nand U24040 (N_24040,N_22809,N_23055);
or U24041 (N_24041,N_23662,N_22573);
nand U24042 (N_24042,N_23328,N_23514);
nand U24043 (N_24043,N_23386,N_22705);
xor U24044 (N_24044,N_23292,N_23019);
nor U24045 (N_24045,N_22400,N_23694);
and U24046 (N_24046,N_22192,N_23973);
nor U24047 (N_24047,N_23410,N_23102);
nor U24048 (N_24048,N_22793,N_23938);
xnor U24049 (N_24049,N_23682,N_23768);
xnor U24050 (N_24050,N_22679,N_23191);
xnor U24051 (N_24051,N_22361,N_23869);
and U24052 (N_24052,N_23242,N_22927);
xor U24053 (N_24053,N_22272,N_22522);
xor U24054 (N_24054,N_22430,N_22484);
or U24055 (N_24055,N_23892,N_23091);
or U24056 (N_24056,N_22617,N_23891);
nor U24057 (N_24057,N_23873,N_23747);
nor U24058 (N_24058,N_23830,N_22284);
or U24059 (N_24059,N_22785,N_23583);
nor U24060 (N_24060,N_23136,N_22390);
xor U24061 (N_24061,N_22051,N_23671);
or U24062 (N_24062,N_23209,N_23581);
or U24063 (N_24063,N_22910,N_23523);
or U24064 (N_24064,N_22741,N_23637);
nand U24065 (N_24065,N_23630,N_23981);
and U24066 (N_24066,N_23918,N_23316);
xnor U24067 (N_24067,N_22194,N_22520);
or U24068 (N_24068,N_22449,N_22307);
nor U24069 (N_24069,N_23353,N_23111);
and U24070 (N_24070,N_23059,N_22839);
nor U24071 (N_24071,N_22460,N_22168);
or U24072 (N_24072,N_22407,N_23341);
xor U24073 (N_24073,N_22571,N_22438);
or U24074 (N_24074,N_22782,N_22924);
nand U24075 (N_24075,N_23937,N_23850);
nand U24076 (N_24076,N_23582,N_22810);
xnor U24077 (N_24077,N_23571,N_23452);
nand U24078 (N_24078,N_22198,N_22893);
or U24079 (N_24079,N_22606,N_23122);
xnor U24080 (N_24080,N_23486,N_22420);
xnor U24081 (N_24081,N_22936,N_22513);
nor U24082 (N_24082,N_23553,N_22031);
and U24083 (N_24083,N_23958,N_22199);
and U24084 (N_24084,N_23082,N_22416);
nor U24085 (N_24085,N_22314,N_23874);
xnor U24086 (N_24086,N_22160,N_23084);
xor U24087 (N_24087,N_23815,N_22553);
and U24088 (N_24088,N_23701,N_23827);
or U24089 (N_24089,N_23161,N_22581);
or U24090 (N_24090,N_23363,N_23854);
and U24091 (N_24091,N_23615,N_22500);
nand U24092 (N_24092,N_22180,N_22405);
and U24093 (N_24093,N_22471,N_23680);
and U24094 (N_24094,N_23144,N_22638);
or U24095 (N_24095,N_22715,N_22653);
xnor U24096 (N_24096,N_23688,N_23362);
nand U24097 (N_24097,N_23197,N_23464);
or U24098 (N_24098,N_22319,N_23796);
nand U24099 (N_24099,N_23700,N_22803);
and U24100 (N_24100,N_23095,N_23016);
nor U24101 (N_24101,N_22290,N_22753);
and U24102 (N_24102,N_22315,N_23404);
nor U24103 (N_24103,N_22585,N_22246);
or U24104 (N_24104,N_22037,N_22652);
xnor U24105 (N_24105,N_23479,N_23644);
or U24106 (N_24106,N_23693,N_23859);
nand U24107 (N_24107,N_22225,N_23636);
nor U24108 (N_24108,N_23928,N_23769);
xnor U24109 (N_24109,N_23993,N_22523);
nand U24110 (N_24110,N_22219,N_22639);
or U24111 (N_24111,N_23924,N_23844);
nor U24112 (N_24112,N_22382,N_23865);
xor U24113 (N_24113,N_23647,N_23424);
xnor U24114 (N_24114,N_22857,N_23751);
nor U24115 (N_24115,N_22918,N_23218);
and U24116 (N_24116,N_23604,N_22850);
and U24117 (N_24117,N_23656,N_23601);
and U24118 (N_24118,N_23158,N_23534);
nor U24119 (N_24119,N_22740,N_23183);
nor U24120 (N_24120,N_23229,N_22669);
xnor U24121 (N_24121,N_22042,N_22961);
or U24122 (N_24122,N_23510,N_23879);
xor U24123 (N_24123,N_23379,N_23692);
nand U24124 (N_24124,N_23244,N_23902);
nor U24125 (N_24125,N_22426,N_22556);
nand U24126 (N_24126,N_23451,N_22871);
or U24127 (N_24127,N_22429,N_22739);
nand U24128 (N_24128,N_22047,N_23719);
nor U24129 (N_24129,N_23421,N_22879);
xor U24130 (N_24130,N_23922,N_22282);
xnor U24131 (N_24131,N_23549,N_22206);
or U24132 (N_24132,N_22408,N_22575);
nor U24133 (N_24133,N_22251,N_22165);
xnor U24134 (N_24134,N_22019,N_22335);
nor U24135 (N_24135,N_22997,N_22525);
or U24136 (N_24136,N_23409,N_23148);
and U24137 (N_24137,N_22445,N_22006);
xor U24138 (N_24138,N_22519,N_22104);
nor U24139 (N_24139,N_22079,N_22217);
or U24140 (N_24140,N_22466,N_23454);
nand U24141 (N_24141,N_22018,N_22759);
and U24142 (N_24142,N_23543,N_23750);
xor U24143 (N_24143,N_22529,N_23318);
and U24144 (N_24144,N_23267,N_23010);
or U24145 (N_24145,N_23202,N_22706);
or U24146 (N_24146,N_22350,N_22559);
nand U24147 (N_24147,N_23776,N_22898);
or U24148 (N_24148,N_22344,N_22130);
or U24149 (N_24149,N_23049,N_23393);
nand U24150 (N_24150,N_22355,N_23907);
xnor U24151 (N_24151,N_22213,N_22953);
nand U24152 (N_24152,N_22279,N_22097);
nand U24153 (N_24153,N_23299,N_23665);
and U24154 (N_24154,N_22332,N_23880);
and U24155 (N_24155,N_23491,N_23133);
and U24156 (N_24156,N_22324,N_23829);
or U24157 (N_24157,N_23172,N_22373);
or U24158 (N_24158,N_23337,N_23356);
nor U24159 (N_24159,N_23575,N_22316);
xnor U24160 (N_24160,N_22274,N_22641);
xor U24161 (N_24161,N_22504,N_22222);
or U24162 (N_24162,N_23434,N_22719);
and U24163 (N_24163,N_22788,N_22291);
xnor U24164 (N_24164,N_23324,N_22300);
xor U24165 (N_24165,N_22325,N_23858);
and U24166 (N_24166,N_22790,N_23274);
nor U24167 (N_24167,N_22542,N_22946);
and U24168 (N_24168,N_22583,N_23822);
and U24169 (N_24169,N_23303,N_22647);
nor U24170 (N_24170,N_22389,N_23635);
and U24171 (N_24171,N_23030,N_23640);
nand U24172 (N_24172,N_23139,N_23901);
nand U24173 (N_24173,N_23975,N_22465);
nand U24174 (N_24174,N_23287,N_22614);
nand U24175 (N_24175,N_23738,N_22494);
and U24176 (N_24176,N_23734,N_23812);
and U24177 (N_24177,N_22680,N_23990);
or U24178 (N_24178,N_22345,N_22477);
or U24179 (N_24179,N_22271,N_22989);
or U24180 (N_24180,N_22726,N_22045);
or U24181 (N_24181,N_23847,N_23391);
nand U24182 (N_24182,N_22040,N_22061);
xor U24183 (N_24183,N_23475,N_23849);
xnor U24184 (N_24184,N_23346,N_23243);
nor U24185 (N_24185,N_23173,N_22384);
xor U24186 (N_24186,N_23396,N_23749);
xor U24187 (N_24187,N_23895,N_22299);
nor U24188 (N_24188,N_22818,N_22721);
or U24189 (N_24189,N_23855,N_22895);
and U24190 (N_24190,N_23284,N_23995);
nand U24191 (N_24191,N_22036,N_23532);
or U24192 (N_24192,N_22624,N_23802);
and U24193 (N_24193,N_23281,N_22173);
nor U24194 (N_24194,N_23471,N_22922);
xnor U24195 (N_24195,N_23338,N_23011);
and U24196 (N_24196,N_22044,N_23283);
nand U24197 (N_24197,N_23558,N_22814);
nand U24198 (N_24198,N_23127,N_23293);
nor U24199 (N_24199,N_23227,N_22386);
nor U24200 (N_24200,N_22185,N_23645);
xor U24201 (N_24201,N_23951,N_22530);
nor U24202 (N_24202,N_22101,N_22088);
and U24203 (N_24203,N_23350,N_23729);
nor U24204 (N_24204,N_22055,N_23529);
nand U24205 (N_24205,N_23089,N_22428);
and U24206 (N_24206,N_22352,N_22550);
or U24207 (N_24207,N_23867,N_22904);
or U24208 (N_24208,N_23099,N_23355);
nand U24209 (N_24209,N_22693,N_22969);
or U24210 (N_24210,N_23717,N_22143);
and U24211 (N_24211,N_23461,N_23041);
xnor U24212 (N_24212,N_23807,N_23864);
nand U24213 (N_24213,N_23258,N_22781);
xor U24214 (N_24214,N_22096,N_23881);
and U24215 (N_24215,N_23005,N_23264);
and U24216 (N_24216,N_23509,N_22303);
and U24217 (N_24217,N_23126,N_22489);
or U24218 (N_24218,N_23224,N_22737);
nand U24219 (N_24219,N_22634,N_22787);
or U24220 (N_24220,N_23828,N_22837);
nor U24221 (N_24221,N_22586,N_22510);
nor U24222 (N_24222,N_22800,N_22865);
nor U24223 (N_24223,N_22066,N_22881);
xnor U24224 (N_24224,N_22674,N_22369);
or U24225 (N_24225,N_22457,N_23226);
or U24226 (N_24226,N_23129,N_22840);
or U24227 (N_24227,N_23265,N_23012);
or U24228 (N_24228,N_22661,N_23763);
nor U24229 (N_24229,N_22847,N_22435);
xor U24230 (N_24230,N_23256,N_23949);
or U24231 (N_24231,N_23070,N_23412);
and U24232 (N_24232,N_23652,N_23841);
xor U24233 (N_24233,N_23882,N_22568);
nand U24234 (N_24234,N_23695,N_22499);
xor U24235 (N_24235,N_22012,N_22650);
xor U24236 (N_24236,N_22610,N_23978);
and U24237 (N_24237,N_23706,N_22368);
or U24238 (N_24238,N_23629,N_23395);
nand U24239 (N_24239,N_22409,N_22188);
nand U24240 (N_24240,N_23320,N_22649);
xnor U24241 (N_24241,N_22376,N_23926);
and U24242 (N_24242,N_22630,N_22032);
or U24243 (N_24243,N_22343,N_22806);
or U24244 (N_24244,N_23323,N_23171);
xnor U24245 (N_24245,N_23247,N_22444);
and U24246 (N_24246,N_22270,N_23221);
and U24247 (N_24247,N_23440,N_23413);
nor U24248 (N_24248,N_23760,N_22779);
nor U24249 (N_24249,N_22545,N_22544);
or U24250 (N_24250,N_23966,N_22998);
and U24251 (N_24251,N_23754,N_23217);
and U24252 (N_24252,N_23810,N_22473);
and U24253 (N_24253,N_23764,N_22897);
and U24254 (N_24254,N_22498,N_22704);
nand U24255 (N_24255,N_22849,N_23568);
and U24256 (N_24256,N_22958,N_23616);
or U24257 (N_24257,N_22822,N_22038);
xor U24258 (N_24258,N_22629,N_22421);
or U24259 (N_24259,N_22132,N_23824);
nand U24260 (N_24260,N_22141,N_23081);
or U24261 (N_24261,N_22950,N_23033);
or U24262 (N_24262,N_23381,N_22472);
nor U24263 (N_24263,N_22099,N_22231);
nor U24264 (N_24264,N_23605,N_22215);
nor U24265 (N_24265,N_22298,N_23105);
nand U24266 (N_24266,N_23067,N_23117);
nand U24267 (N_24267,N_23388,N_23024);
xor U24268 (N_24268,N_23277,N_22713);
nand U24269 (N_24269,N_23118,N_23811);
and U24270 (N_24270,N_23758,N_22985);
and U24271 (N_24271,N_23083,N_23726);
xnor U24272 (N_24272,N_23985,N_22372);
nor U24273 (N_24273,N_23567,N_23519);
or U24274 (N_24274,N_22172,N_23051);
and U24275 (N_24275,N_23651,N_23482);
nor U24276 (N_24276,N_22524,N_23596);
and U24277 (N_24277,N_23294,N_22714);
nand U24278 (N_24278,N_22268,N_23757);
or U24279 (N_24279,N_22375,N_22452);
nor U24280 (N_24280,N_23715,N_23253);
and U24281 (N_24281,N_22242,N_23205);
xor U24282 (N_24282,N_22486,N_23301);
or U24283 (N_24283,N_23453,N_23296);
and U24284 (N_24284,N_22068,N_22570);
and U24285 (N_24285,N_23876,N_22505);
nor U24286 (N_24286,N_22532,N_22861);
and U24287 (N_24287,N_22701,N_23472);
xor U24288 (N_24288,N_22432,N_23074);
nand U24289 (N_24289,N_22593,N_22437);
nor U24290 (N_24290,N_22869,N_23298);
or U24291 (N_24291,N_22979,N_23943);
and U24292 (N_24292,N_23013,N_22128);
xnor U24293 (N_24293,N_23128,N_23150);
and U24294 (N_24294,N_23839,N_23383);
nand U24295 (N_24295,N_22076,N_23385);
nor U24296 (N_24296,N_22440,N_23496);
and U24297 (N_24297,N_23580,N_23257);
or U24298 (N_24298,N_22339,N_23003);
or U24299 (N_24299,N_23348,N_23886);
or U24300 (N_24300,N_22091,N_23029);
nor U24301 (N_24301,N_22451,N_22626);
nor U24302 (N_24302,N_23545,N_23213);
nand U24303 (N_24303,N_23357,N_23378);
nor U24304 (N_24304,N_22598,N_22124);
nor U24305 (N_24305,N_23911,N_22265);
xnor U24306 (N_24306,N_23427,N_23487);
and U24307 (N_24307,N_22763,N_23955);
xor U24308 (N_24308,N_23554,N_23326);
or U24309 (N_24309,N_22266,N_23976);
nand U24310 (N_24310,N_22882,N_23309);
nor U24311 (N_24311,N_23007,N_23727);
xnor U24312 (N_24312,N_22381,N_23774);
nand U24313 (N_24313,N_23746,N_23959);
xor U24314 (N_24314,N_23889,N_22395);
and U24315 (N_24315,N_22878,N_22289);
and U24316 (N_24316,N_22379,N_23790);
nand U24317 (N_24317,N_23617,N_23164);
xnor U24318 (N_24318,N_22948,N_22117);
or U24319 (N_24319,N_23050,N_23428);
nand U24320 (N_24320,N_23587,N_23480);
and U24321 (N_24321,N_22965,N_23062);
and U24322 (N_24322,N_23788,N_22476);
nor U24323 (N_24323,N_22819,N_22619);
nor U24324 (N_24324,N_22053,N_23908);
or U24325 (N_24325,N_23610,N_23942);
nor U24326 (N_24326,N_22092,N_23679);
nand U24327 (N_24327,N_23463,N_22880);
xnor U24328 (N_24328,N_22666,N_23220);
xnor U24329 (N_24329,N_22521,N_22905);
or U24330 (N_24330,N_22761,N_23149);
xor U24331 (N_24331,N_23836,N_22872);
and U24332 (N_24332,N_23336,N_22323);
and U24333 (N_24333,N_22596,N_22243);
or U24334 (N_24334,N_23238,N_22868);
xor U24335 (N_24335,N_23308,N_22731);
nand U24336 (N_24336,N_22007,N_22186);
nor U24337 (N_24337,N_22921,N_23579);
nor U24338 (N_24338,N_22866,N_22838);
nor U24339 (N_24339,N_22312,N_22588);
xnor U24340 (N_24340,N_22812,N_22118);
nor U24341 (N_24341,N_23056,N_23478);
xor U24342 (N_24342,N_23663,N_22930);
or U24343 (N_24343,N_22703,N_22054);
nor U24344 (N_24344,N_23916,N_22228);
nand U24345 (N_24345,N_23712,N_23702);
nand U24346 (N_24346,N_23075,N_23270);
or U24347 (N_24347,N_23069,N_22580);
nand U24348 (N_24348,N_23290,N_22260);
nor U24349 (N_24349,N_22720,N_23547);
or U24350 (N_24350,N_22082,N_23090);
or U24351 (N_24351,N_22587,N_23499);
nor U24352 (N_24352,N_23585,N_23408);
nor U24353 (N_24353,N_22968,N_22887);
xnor U24354 (N_24354,N_23952,N_22563);
or U24355 (N_24355,N_22676,N_22665);
nor U24356 (N_24356,N_23664,N_22135);
and U24357 (N_24357,N_22709,N_23762);
or U24358 (N_24358,N_22516,N_22483);
nand U24359 (N_24359,N_23944,N_23599);
and U24360 (N_24360,N_22972,N_23080);
nor U24361 (N_24361,N_23704,N_23015);
nor U24362 (N_24362,N_23957,N_22766);
and U24363 (N_24363,N_22977,N_23894);
and U24364 (N_24364,N_22727,N_22456);
nand U24365 (N_24365,N_23542,N_22827);
nand U24366 (N_24366,N_22526,N_23063);
nor U24367 (N_24367,N_22202,N_23494);
and U24368 (N_24368,N_23619,N_23513);
nor U24369 (N_24369,N_23207,N_23225);
and U24370 (N_24370,N_22468,N_23313);
nor U24371 (N_24371,N_22286,N_22728);
nor U24372 (N_24372,N_22631,N_23940);
nand U24373 (N_24373,N_23170,N_22710);
or U24374 (N_24374,N_22942,N_22043);
nor U24375 (N_24375,N_23590,N_23088);
xnor U24376 (N_24376,N_22919,N_22609);
nand U24377 (N_24377,N_23939,N_22116);
xnor U24378 (N_24378,N_22152,N_23736);
nor U24379 (N_24379,N_22334,N_23756);
or U24380 (N_24380,N_23797,N_23045);
nand U24381 (N_24381,N_23398,N_22537);
xor U24382 (N_24382,N_23493,N_23562);
nand U24383 (N_24383,N_22518,N_23273);
xnor U24384 (N_24384,N_23216,N_23160);
xnor U24385 (N_24385,N_22613,N_23689);
nand U24386 (N_24386,N_23569,N_23351);
or U24387 (N_24387,N_23646,N_22789);
xor U24388 (N_24388,N_22492,N_23743);
xnor U24389 (N_24389,N_23910,N_22797);
nand U24390 (N_24390,N_23250,N_23439);
nor U24391 (N_24391,N_23709,N_22167);
nor U24392 (N_24392,N_23373,N_22966);
or U24393 (N_24393,N_22595,N_23426);
xor U24394 (N_24394,N_22623,N_23655);
or U24395 (N_24395,N_22552,N_22001);
xnor U24396 (N_24396,N_22184,N_22149);
and U24397 (N_24397,N_23786,N_23638);
nor U24398 (N_24398,N_23598,N_22275);
xor U24399 (N_24399,N_22115,N_23626);
or U24400 (N_24400,N_23988,N_22798);
nor U24401 (N_24401,N_22221,N_22347);
xor U24402 (N_24402,N_22826,N_23322);
or U24403 (N_24403,N_22000,N_23823);
nor U24404 (N_24404,N_22467,N_22176);
nand U24405 (N_24405,N_23027,N_23512);
xnor U24406 (N_24406,N_23177,N_23608);
nor U24407 (N_24407,N_22327,N_22396);
or U24408 (N_24408,N_22398,N_23877);
nor U24409 (N_24409,N_23917,N_22259);
nand U24410 (N_24410,N_23135,N_23962);
and U24411 (N_24411,N_23086,N_23595);
nand U24412 (N_24412,N_23792,N_22008);
xnor U24413 (N_24413,N_23678,N_22073);
xor U24414 (N_24414,N_22236,N_23187);
nor U24415 (N_24415,N_22939,N_23584);
nor U24416 (N_24416,N_22917,N_23967);
nand U24417 (N_24417,N_23455,N_22069);
nor U24418 (N_24418,N_23371,N_23321);
nand U24419 (N_24419,N_23401,N_22424);
nand U24420 (N_24420,N_23036,N_23517);
xnor U24421 (N_24421,N_22297,N_23536);
or U24422 (N_24422,N_22658,N_23820);
xor U24423 (N_24423,N_22877,N_22178);
nand U24424 (N_24424,N_22696,N_22496);
or U24425 (N_24425,N_23208,N_22855);
nor U24426 (N_24426,N_22991,N_23132);
and U24427 (N_24427,N_23960,N_23929);
xor U24428 (N_24428,N_23870,N_23846);
xnor U24429 (N_24429,N_23745,N_22955);
nor U24430 (N_24430,N_23772,N_22825);
nand U24431 (N_24431,N_22589,N_23956);
nor U24432 (N_24432,N_23101,N_22913);
or U24433 (N_24433,N_22551,N_22663);
nand U24434 (N_24434,N_23146,N_22870);
and U24435 (N_24435,N_23537,N_22729);
or U24436 (N_24436,N_23528,N_22888);
nand U24437 (N_24437,N_23306,N_23643);
and U24438 (N_24438,N_22337,N_23449);
and U24439 (N_24439,N_23673,N_22628);
nand U24440 (N_24440,N_23269,N_23785);
nor U24441 (N_24441,N_23262,N_22511);
nand U24442 (N_24442,N_22828,N_22086);
or U24443 (N_24443,N_23705,N_23883);
or U24444 (N_24444,N_23525,N_22480);
nand U24445 (N_24445,N_22774,N_22675);
and U24446 (N_24446,N_23648,N_23904);
nand U24447 (N_24447,N_23707,N_23037);
nor U24448 (N_24448,N_23612,N_23420);
nand U24449 (N_24449,N_22603,N_22767);
xor U24450 (N_24450,N_22123,N_23884);
xor U24451 (N_24451,N_22817,N_23686);
nor U24452 (N_24452,N_22656,N_23233);
xor U24453 (N_24453,N_22931,N_22605);
and U24454 (N_24454,N_23983,N_23900);
or U24455 (N_24455,N_23950,N_23035);
and U24456 (N_24456,N_22683,N_22328);
xnor U24457 (N_24457,N_23838,N_22821);
or U24458 (N_24458,N_22144,N_22406);
nor U24459 (N_24459,N_23893,N_23502);
xor U24460 (N_24460,N_23609,N_23863);
nand U24461 (N_24461,N_22133,N_22891);
and U24462 (N_24462,N_22830,N_23941);
and U24463 (N_24463,N_22205,N_23994);
nand U24464 (N_24464,N_23739,N_22945);
and U24465 (N_24465,N_23564,N_23009);
xnor U24466 (N_24466,N_23022,N_22028);
xor U24467 (N_24467,N_23137,N_23659);
xor U24468 (N_24468,N_22775,N_23325);
or U24469 (N_24469,N_22240,N_23906);
nand U24470 (N_24470,N_23065,N_23675);
or U24471 (N_24471,N_23156,N_23302);
or U24472 (N_24472,N_22153,N_23186);
xor U24473 (N_24473,N_23223,N_22801);
nor U24474 (N_24474,N_23165,N_23175);
xor U24475 (N_24475,N_22899,N_22264);
or U24476 (N_24476,N_23661,N_23592);
xnor U24477 (N_24477,N_22064,N_23555);
nand U24478 (N_24478,N_23733,N_23563);
nand U24479 (N_24479,N_22170,N_22293);
or U24480 (N_24480,N_22121,N_23968);
and U24481 (N_24481,N_23488,N_22501);
or U24482 (N_24482,N_23422,N_22920);
or U24483 (N_24483,N_22311,N_22657);
nor U24484 (N_24484,N_23072,N_22851);
and U24485 (N_24485,N_23984,N_23115);
nor U24486 (N_24486,N_22377,N_22987);
xnor U24487 (N_24487,N_22755,N_23335);
or U24488 (N_24488,N_23108,N_23834);
xnor U24489 (N_24489,N_22313,N_23498);
xor U24490 (N_24490,N_23382,N_23199);
nand U24491 (N_24491,N_22214,N_23921);
nand U24492 (N_24492,N_22094,N_22248);
nand U24493 (N_24493,N_22621,N_22114);
or U24494 (N_24494,N_23766,N_22590);
xnor U24495 (N_24495,N_23189,N_23222);
xnor U24496 (N_24496,N_23597,N_23722);
or U24497 (N_24497,N_22479,N_22387);
and U24498 (N_24498,N_23506,N_23687);
nor U24499 (N_24499,N_23327,N_23711);
nand U24500 (N_24500,N_22738,N_22034);
nand U24501 (N_24501,N_23046,N_23896);
nand U24502 (N_24502,N_23288,N_22558);
nor U24503 (N_24503,N_22125,N_22495);
and U24504 (N_24504,N_23085,N_23219);
and U24505 (N_24505,N_23178,N_23145);
and U24506 (N_24506,N_23406,N_22363);
xnor U24507 (N_24507,N_23625,N_22276);
nand U24508 (N_24508,N_22383,N_22686);
and U24509 (N_24509,N_23992,N_23948);
or U24510 (N_24510,N_23359,N_23367);
or U24511 (N_24511,N_23215,N_22937);
and U24512 (N_24512,N_22633,N_22288);
nand U24513 (N_24513,N_22151,N_22155);
or U24514 (N_24514,N_22250,N_22554);
nor U24515 (N_24515,N_23031,N_22508);
or U24516 (N_24516,N_23969,N_22072);
nand U24517 (N_24517,N_22885,N_23914);
or U24518 (N_24518,N_22263,N_22642);
nor U24519 (N_24519,N_23370,N_23295);
and U24520 (N_24520,N_22422,N_22848);
nand U24521 (N_24521,N_22035,N_23813);
xnor U24522 (N_24522,N_23002,N_22805);
or U24523 (N_24523,N_22843,N_22067);
nor U24524 (N_24524,N_23755,N_23423);
nor U24525 (N_24525,N_23767,N_22964);
or U24526 (N_24526,N_23526,N_23166);
nor U24527 (N_24527,N_22089,N_23228);
nand U24528 (N_24528,N_22547,N_23252);
nor U24529 (N_24529,N_22829,N_22894);
and U24530 (N_24530,N_23354,N_22566);
or U24531 (N_24531,N_23140,N_22137);
or U24532 (N_24532,N_23843,N_22431);
nand U24533 (N_24533,N_22211,N_23996);
and U24534 (N_24534,N_22497,N_22212);
xor U24535 (N_24535,N_23885,N_23000);
xor U24536 (N_24536,N_22836,N_22158);
nand U24537 (N_24537,N_23759,N_23698);
or U24538 (N_24538,N_22697,N_23780);
nand U24539 (N_24539,N_22863,N_23920);
xnor U24540 (N_24540,N_23540,N_22503);
nand U24541 (N_24541,N_22309,N_22462);
or U24542 (N_24542,N_23100,N_22139);
nor U24543 (N_24543,N_22063,N_22730);
nand U24544 (N_24544,N_23946,N_22247);
nor U24545 (N_24545,N_22485,N_23039);
nor U24546 (N_24546,N_23544,N_22667);
and U24547 (N_24547,N_22120,N_22446);
or U24548 (N_24548,N_23485,N_22230);
xor U24549 (N_24549,N_22209,N_23181);
or U24550 (N_24550,N_22694,N_23465);
and U24551 (N_24551,N_22237,N_22684);
xnor U24552 (N_24552,N_23697,N_22986);
nor U24553 (N_24553,N_22954,N_23042);
nand U24554 (N_24554,N_22280,N_23497);
or U24555 (N_24555,N_23114,N_23445);
or U24556 (N_24556,N_23490,N_22983);
nor U24557 (N_24557,N_22370,N_22098);
xnor U24558 (N_24558,N_23188,N_22938);
nand U24559 (N_24559,N_23204,N_22039);
nor U24560 (N_24560,N_23347,N_23248);
nand U24561 (N_24561,N_22856,N_22835);
nor U24562 (N_24562,N_22695,N_22952);
and U24563 (N_24563,N_22304,N_22834);
and U24564 (N_24564,N_22253,N_23212);
and U24565 (N_24565,N_22346,N_22200);
xor U24566 (N_24566,N_23551,N_23866);
nor U24567 (N_24567,N_22340,N_22947);
or U24568 (N_24568,N_22052,N_23263);
nor U24569 (N_24569,N_23163,N_23550);
xnor U24570 (N_24570,N_22150,N_23268);
nor U24571 (N_24571,N_23400,N_22749);
and U24572 (N_24572,N_23315,N_23038);
nor U24573 (N_24573,N_23236,N_23116);
xnor U24574 (N_24574,N_22415,N_22533);
nor U24575 (N_24575,N_23286,N_23773);
nand U24576 (N_24576,N_22487,N_23182);
xor U24577 (N_24577,N_22366,N_22976);
xnor U24578 (N_24578,N_23106,N_22393);
or U24579 (N_24579,N_23380,N_23684);
nor U24580 (N_24580,N_23531,N_23254);
and U24581 (N_24581,N_22778,N_22794);
and U24582 (N_24582,N_22075,N_22682);
nor U24583 (N_24583,N_23913,N_22203);
nand U24584 (N_24584,N_22059,N_22320);
xor U24585 (N_24585,N_22769,N_23925);
or U24586 (N_24586,N_22463,N_22475);
or U24587 (N_24587,N_23691,N_23076);
nand U24588 (N_24588,N_23852,N_22724);
or U24589 (N_24589,N_22169,N_23657);
and U24590 (N_24590,N_22539,N_23699);
and U24591 (N_24591,N_23795,N_23176);
and U24592 (N_24592,N_22455,N_23991);
nand U24593 (N_24593,N_22470,N_22644);
xor U24594 (N_24594,N_22540,N_22002);
nor U24595 (N_24595,N_22757,N_22027);
nand U24596 (N_24596,N_23157,N_22391);
nand U24597 (N_24597,N_22717,N_22005);
nor U24598 (N_24598,N_23436,N_22014);
xor U24599 (N_24599,N_23043,N_22254);
and U24600 (N_24600,N_22159,N_23912);
nand U24601 (N_24601,N_22296,N_23203);
nand U24602 (N_24602,N_22338,N_23483);
nand U24603 (N_24603,N_23737,N_22241);
nor U24604 (N_24604,N_22980,N_22783);
and U24605 (N_24605,N_23862,N_23622);
or U24606 (N_24606,N_22784,N_22318);
or U24607 (N_24607,N_22103,N_23198);
or U24608 (N_24608,N_23402,N_23155);
or U24609 (N_24609,N_23061,N_22220);
and U24610 (N_24610,N_23632,N_23814);
xnor U24611 (N_24611,N_22057,N_22996);
xnor U24612 (N_24612,N_23387,N_22592);
nor U24613 (N_24613,N_23448,N_22978);
or U24614 (N_24614,N_22569,N_22085);
xnor U24615 (N_24615,N_22535,N_22698);
or U24616 (N_24616,N_22146,N_23159);
or U24617 (N_24617,N_22074,N_22808);
and U24618 (N_24618,N_23103,N_23153);
or U24619 (N_24619,N_22062,N_22515);
nor U24620 (N_24620,N_22777,N_22056);
and U24621 (N_24621,N_22916,N_22912);
nor U24622 (N_24622,N_22591,N_22423);
or U24623 (N_24623,N_23334,N_23271);
xnor U24624 (N_24624,N_22560,N_23057);
and U24625 (N_24625,N_22105,N_23077);
or U24626 (N_24626,N_22858,N_22394);
xor U24627 (N_24627,N_23565,N_23800);
nor U24628 (N_24628,N_22883,N_22671);
nand U24629 (N_24629,N_23546,N_23817);
or U24630 (N_24630,N_22295,N_23731);
xnor U24631 (N_24631,N_23724,N_23196);
nor U24632 (N_24632,N_22876,N_22411);
or U24633 (N_24633,N_22126,N_22078);
or U24634 (N_24634,N_23871,N_22030);
nand U24635 (N_24635,N_22517,N_23837);
nand U24636 (N_24636,N_22227,N_23779);
or U24637 (N_24637,N_23473,N_22681);
and U24638 (N_24638,N_23201,N_22163);
nor U24639 (N_24639,N_22745,N_22960);
and U24640 (N_24640,N_23477,N_22025);
or U24641 (N_24641,N_23376,N_22561);
and U24642 (N_24642,N_23539,N_23516);
or U24643 (N_24643,N_23138,N_23631);
nand U24644 (N_24644,N_23588,N_22110);
or U24645 (N_24645,N_23972,N_23765);
nand U24646 (N_24646,N_23113,N_23500);
nand U24647 (N_24647,N_22365,N_22065);
and U24648 (N_24648,N_22441,N_22349);
and U24649 (N_24649,N_23667,N_22329);
nor U24650 (N_24650,N_22138,N_23230);
nor U24651 (N_24651,N_23096,N_23753);
and U24652 (N_24652,N_22196,N_23560);
nor U24653 (N_24653,N_22443,N_23927);
and U24654 (N_24654,N_23312,N_22469);
or U24655 (N_24655,N_23653,N_22678);
or U24656 (N_24656,N_22833,N_22341);
xnor U24657 (N_24657,N_22235,N_22677);
and U24658 (N_24658,N_23481,N_22201);
and U24659 (N_24659,N_22725,N_22823);
and U24660 (N_24660,N_22336,N_23241);
or U24661 (N_24661,N_22354,N_23570);
nand U24662 (N_24662,N_23048,N_23405);
xnor U24663 (N_24663,N_22207,N_23831);
or U24664 (N_24664,N_23518,N_23818);
and U24665 (N_24665,N_23690,N_23669);
or U24666 (N_24666,N_22764,N_22397);
nor U24667 (N_24667,N_23979,N_23435);
nand U24668 (N_24668,N_22579,N_23331);
xnor U24669 (N_24669,N_22333,N_23441);
nor U24670 (N_24670,N_22439,N_22244);
nand U24671 (N_24671,N_22048,N_23340);
nor U24672 (N_24672,N_22832,N_22148);
xor U24673 (N_24673,N_22816,N_22004);
and U24674 (N_24674,N_22758,N_22908);
or U24675 (N_24675,N_22538,N_23639);
nor U24676 (N_24676,N_23300,N_22732);
or U24677 (N_24677,N_22903,N_23285);
nand U24678 (N_24678,N_22136,N_22807);
xnor U24679 (N_24679,N_22493,N_23375);
nand U24680 (N_24680,N_23566,N_22095);
nand U24681 (N_24681,N_23718,N_23963);
and U24682 (N_24682,N_22901,N_22702);
or U24683 (N_24683,N_22612,N_22013);
xor U24684 (N_24684,N_23696,N_22189);
and U24685 (N_24685,N_23190,N_23068);
xor U24686 (N_24686,N_22831,N_22578);
nor U24687 (N_24687,N_22070,N_22414);
nor U24688 (N_24688,N_22425,N_23443);
and U24689 (N_24689,N_22984,N_23469);
xor U24690 (N_24690,N_22860,N_23793);
xnor U24691 (N_24691,N_23064,N_22765);
nand U24692 (N_24692,N_23930,N_23620);
xor U24693 (N_24693,N_23603,N_23474);
nand U24694 (N_24694,N_23501,N_22302);
xor U24695 (N_24695,N_22142,N_23853);
xor U24696 (N_24696,N_22107,N_23314);
nand U24697 (N_24697,N_23018,N_22842);
nor U24698 (N_24698,N_22208,N_23778);
or U24699 (N_24699,N_22478,N_23710);
and U24700 (N_24700,N_22873,N_22360);
or U24701 (N_24701,N_22925,N_23977);
nand U24702 (N_24702,N_22768,N_23999);
nand U24703 (N_24703,N_23961,N_23771);
nor U24704 (N_24704,N_23032,N_23026);
or U24705 (N_24705,N_23447,N_22923);
xor U24706 (N_24706,N_22106,N_22273);
nor U24707 (N_24707,N_23344,N_23364);
nor U24708 (N_24708,N_23860,N_22562);
and U24709 (N_24709,N_22975,N_22464);
xnor U24710 (N_24710,N_23071,N_22670);
and U24711 (N_24711,N_23369,N_22957);
and U24712 (N_24712,N_22257,N_23414);
xnor U24713 (N_24713,N_23557,N_22353);
or U24714 (N_24714,N_22654,N_23982);
nand U24715 (N_24715,N_22245,N_23676);
or U24716 (N_24716,N_22016,N_23280);
nor U24717 (N_24717,N_23109,N_22867);
nor U24718 (N_24718,N_22081,N_23232);
or U24719 (N_24719,N_22864,N_22326);
nand U24720 (N_24720,N_23120,N_23131);
xor U24721 (N_24721,N_23192,N_22024);
nand U24722 (N_24722,N_23297,N_23174);
nand U24723 (N_24723,N_23134,N_22301);
xor U24724 (N_24724,N_22374,N_22308);
xor U24725 (N_24725,N_22454,N_23561);
or U24726 (N_24726,N_23527,N_22023);
and U24727 (N_24727,N_22292,N_23457);
xor U24728 (N_24728,N_23169,N_22140);
nor U24729 (N_24729,N_23432,N_22229);
nand U24730 (N_24730,N_22664,N_23425);
nor U24731 (N_24731,N_23372,N_23278);
nor U24732 (N_24732,N_23851,N_23442);
nor U24733 (N_24733,N_22963,N_23417);
and U24734 (N_24734,N_22699,N_22567);
xor U24735 (N_24735,N_23791,N_23602);
nor U24736 (N_24736,N_23279,N_23017);
and U24737 (N_24737,N_22358,N_22413);
or U24738 (N_24738,N_23361,N_23728);
and U24739 (N_24739,N_22640,N_22080);
or U24740 (N_24740,N_23317,N_23794);
or U24741 (N_24741,N_22646,N_22041);
and U24742 (N_24742,N_22772,N_22306);
nand U24743 (N_24743,N_23808,N_23624);
xnor U24744 (N_24744,N_23856,N_22928);
xnor U24745 (N_24745,N_22815,N_22362);
xor U24746 (N_24746,N_22607,N_23235);
or U24747 (N_24747,N_22100,N_23028);
nor U24748 (N_24748,N_23123,N_22058);
or U24749 (N_24749,N_23433,N_23458);
xnor U24750 (N_24750,N_23397,N_23008);
and U24751 (N_24751,N_22404,N_22604);
or U24752 (N_24752,N_23857,N_22410);
and U24753 (N_24753,N_22691,N_22278);
xor U24754 (N_24754,N_23923,N_22743);
and U24755 (N_24755,N_22700,N_22177);
nand U24756 (N_24756,N_22733,N_23628);
xnor U24757 (N_24757,N_23735,N_23600);
or U24758 (N_24758,N_23211,N_22204);
and U24759 (N_24759,N_22359,N_23720);
nand U24760 (N_24760,N_23130,N_22122);
and U24761 (N_24761,N_22643,N_22620);
and U24762 (N_24762,N_23541,N_23945);
nand U24763 (N_24763,N_22565,N_23044);
nand U24764 (N_24764,N_22956,N_22084);
or U24765 (N_24765,N_22734,N_23801);
nand U24766 (N_24766,N_23974,N_23674);
and U24767 (N_24767,N_23110,N_22776);
nor U24768 (N_24768,N_22884,N_22342);
xor U24769 (N_24769,N_23255,N_23366);
nand U24770 (N_24770,N_22399,N_22915);
or U24771 (N_24771,N_22283,N_22557);
nor U24772 (N_24772,N_22791,N_23495);
and U24773 (N_24773,N_23845,N_22754);
and U24774 (N_24774,N_22951,N_22597);
nor U24775 (N_24775,N_22608,N_23154);
or U24776 (N_24776,N_23730,N_23708);
nand U24777 (N_24777,N_22962,N_23761);
nor U24778 (N_24778,N_22549,N_23915);
nor U24779 (N_24779,N_23716,N_22179);
nand U24780 (N_24780,N_22156,N_22010);
nand U24781 (N_24781,N_23627,N_22294);
xor U24782 (N_24782,N_23060,N_23021);
nand U24783 (N_24783,N_22392,N_22305);
and U24784 (N_24784,N_23970,N_23001);
nand U24785 (N_24785,N_22418,N_23805);
xor U24786 (N_24786,N_23054,N_23713);
or U24787 (N_24787,N_22748,N_23832);
nand U24788 (N_24788,N_23505,N_22488);
or U24789 (N_24789,N_22886,N_22926);
nor U24790 (N_24790,N_23522,N_22796);
nor U24791 (N_24791,N_22746,N_23611);
nand U24792 (N_24792,N_23868,N_23349);
or U24793 (N_24793,N_23533,N_22351);
or U24794 (N_24794,N_23360,N_22959);
nand U24795 (N_24795,N_22491,N_23725);
xnor U24796 (N_24796,N_23594,N_23444);
xnor U24797 (N_24797,N_22685,N_23394);
nor U24798 (N_24798,N_22197,N_23887);
or U24799 (N_24799,N_23593,N_23685);
nand U24800 (N_24800,N_22442,N_22417);
xnor U24801 (N_24801,N_22281,N_22906);
and U24802 (N_24802,N_22820,N_22949);
nor U24803 (N_24803,N_22574,N_23840);
nand U24804 (N_24804,N_22481,N_23621);
xnor U24805 (N_24805,N_22434,N_22600);
or U24806 (N_24806,N_22929,N_23613);
xor U24807 (N_24807,N_23775,N_22655);
nand U24808 (N_24808,N_23239,N_23521);
nor U24809 (N_24809,N_22995,N_22403);
nand U24810 (N_24810,N_22269,N_22090);
and U24811 (N_24811,N_22722,N_22171);
xor U24812 (N_24812,N_22616,N_22166);
nand U24813 (N_24813,N_23732,N_22907);
or U24814 (N_24814,N_23092,N_23980);
xnor U24815 (N_24815,N_22648,N_23460);
or U24816 (N_24816,N_22747,N_22786);
nor U24817 (N_24817,N_23358,N_22736);
and U24818 (N_24818,N_23898,N_23826);
xor U24819 (N_24819,N_23272,N_22718);
and U24820 (N_24820,N_23740,N_22507);
xor U24821 (N_24821,N_22433,N_23141);
nor U24822 (N_24822,N_23618,N_22127);
and U24823 (N_24823,N_22999,N_23989);
nor U24824 (N_24824,N_22419,N_23650);
nand U24825 (N_24825,N_23249,N_22577);
nor U24826 (N_24826,N_22804,N_23282);
and U24827 (N_24827,N_22402,N_23342);
nand U24828 (N_24828,N_22584,N_22970);
or U24829 (N_24829,N_23508,N_22087);
or U24830 (N_24830,N_22022,N_23143);
or U24831 (N_24831,N_23429,N_22252);
and U24832 (N_24832,N_22071,N_23803);
and U24833 (N_24833,N_22119,N_23703);
xnor U24834 (N_24834,N_23804,N_22009);
nand U24835 (N_24835,N_22601,N_23572);
xnor U24836 (N_24836,N_23237,N_22811);
and U24837 (N_24837,N_23276,N_22474);
or U24838 (N_24838,N_23168,N_22482);
and U24839 (N_24839,N_23079,N_22967);
nand U24840 (N_24840,N_23589,N_23415);
xnor U24841 (N_24841,N_22147,N_23374);
nand U24842 (N_24842,N_22707,N_22458);
xnor U24843 (N_24843,N_23390,N_23781);
nand U24844 (N_24844,N_22933,N_23507);
and U24845 (N_24845,N_23200,N_23909);
nor U24846 (N_24846,N_22175,N_23446);
nor U24847 (N_24847,N_23744,N_22994);
or U24848 (N_24848,N_23552,N_23511);
and U24849 (N_24849,N_22111,N_23919);
nand U24850 (N_24850,N_23259,N_22564);
nand U24851 (N_24851,N_23107,N_23339);
or U24852 (N_24852,N_23658,N_23784);
nand U24853 (N_24853,N_22015,N_23574);
and U24854 (N_24854,N_22615,N_23591);
and U24855 (N_24855,N_22988,N_23677);
nand U24856 (N_24856,N_23097,N_23752);
or U24857 (N_24857,N_22049,N_23897);
nor U24858 (N_24858,N_22134,N_23586);
or U24859 (N_24859,N_23660,N_23121);
and U24860 (N_24860,N_23933,N_22723);
nor U24861 (N_24861,N_23683,N_23503);
nor U24862 (N_24862,N_22688,N_23634);
nand U24863 (N_24863,N_23275,N_23559);
and U24864 (N_24864,N_23672,N_22033);
or U24865 (N_24865,N_22841,N_22191);
nor U24866 (N_24866,N_22321,N_23467);
nor U24867 (N_24867,N_23935,N_23953);
xor U24868 (N_24868,N_22190,N_23210);
nor U24869 (N_24869,N_22509,N_23789);
nand U24870 (N_24870,N_23330,N_23782);
nand U24871 (N_24871,N_23094,N_23125);
nand U24872 (N_24872,N_22527,N_23649);
and U24873 (N_24873,N_23087,N_23392);
or U24874 (N_24874,N_22932,N_22093);
nand U24875 (N_24875,N_23642,N_22287);
xnor U24876 (N_24876,N_23142,N_23240);
and U24877 (N_24877,N_22310,N_23504);
nor U24878 (N_24878,N_23903,N_23614);
nand U24879 (N_24879,N_22060,N_23548);
nor U24880 (N_24880,N_22255,N_22129);
nand U24881 (N_24881,N_23020,N_23633);
and U24882 (N_24882,N_22356,N_23468);
and U24883 (N_24883,N_23437,N_22109);
xor U24884 (N_24884,N_22944,N_22914);
and U24885 (N_24885,N_22660,N_22162);
xor U24886 (N_24886,N_23180,N_22367);
and U24887 (N_24887,N_22651,N_22108);
nor U24888 (N_24888,N_23152,N_22943);
nand U24889 (N_24889,N_22512,N_23416);
xnor U24890 (N_24890,N_22385,N_22582);
nand U24891 (N_24891,N_22845,N_22599);
xor U24892 (N_24892,N_23816,N_23809);
nor U24893 (N_24893,N_22003,N_23947);
nand U24894 (N_24894,N_22795,N_22602);
nor U24895 (N_24895,N_23014,N_23833);
xnor U24896 (N_24896,N_22760,N_23419);
and U24897 (N_24897,N_22195,N_22183);
nand U24898 (N_24898,N_22672,N_23742);
nand U24899 (N_24899,N_22874,N_23112);
and U24900 (N_24900,N_22690,N_23714);
xor U24901 (N_24901,N_23799,N_23888);
or U24902 (N_24902,N_22026,N_22216);
xor U24903 (N_24903,N_22348,N_23777);
nand U24904 (N_24904,N_23343,N_22689);
xnor U24905 (N_24905,N_22543,N_23231);
nor U24906 (N_24906,N_23936,N_23819);
and U24907 (N_24907,N_22378,N_23260);
or U24908 (N_24908,N_22780,N_22157);
nand U24909 (N_24909,N_22852,N_22632);
and U24910 (N_24910,N_22625,N_22181);
nor U24911 (N_24911,N_22742,N_22618);
xor U24912 (N_24912,N_23399,N_23431);
xor U24913 (N_24913,N_23931,N_22824);
and U24914 (N_24914,N_23524,N_23723);
nor U24915 (N_24915,N_23783,N_23245);
nor U24916 (N_24916,N_23623,N_22322);
or U24917 (N_24917,N_23119,N_22239);
or U24918 (N_24918,N_22234,N_23098);
nand U24919 (N_24919,N_23954,N_23195);
xnor U24920 (N_24920,N_23450,N_22317);
nor U24921 (N_24921,N_22210,N_22161);
and U24922 (N_24922,N_22813,N_22802);
or U24923 (N_24923,N_22668,N_22502);
nand U24924 (N_24924,N_23606,N_22277);
xnor U24925 (N_24925,N_23998,N_23352);
nand U24926 (N_24926,N_22536,N_23459);
nand U24927 (N_24927,N_22635,N_23311);
or U24928 (N_24928,N_22261,N_22752);
nand U24929 (N_24929,N_22187,N_22771);
or U24930 (N_24930,N_23530,N_22528);
nor U24931 (N_24931,N_23573,N_22555);
or U24932 (N_24932,N_22875,N_22226);
nor U24933 (N_24933,N_23515,N_23179);
or U24934 (N_24934,N_22113,N_23251);
nand U24935 (N_24935,N_23466,N_23578);
nand U24936 (N_24936,N_22708,N_22692);
nor U24937 (N_24937,N_23666,N_22990);
nand U24938 (N_24938,N_23407,N_23305);
nor U24939 (N_24939,N_23835,N_22238);
and U24940 (N_24940,N_22973,N_22233);
xnor U24941 (N_24941,N_23333,N_23825);
or U24942 (N_24942,N_23025,N_22112);
and U24943 (N_24943,N_23654,N_22854);
nor U24944 (N_24944,N_23556,N_23073);
or U24945 (N_24945,N_22576,N_22371);
and U24946 (N_24946,N_22046,N_22662);
nor U24947 (N_24947,N_22131,N_22546);
xor U24948 (N_24948,N_22412,N_23023);
nand U24949 (N_24949,N_22249,N_22548);
or U24950 (N_24950,N_23365,N_22751);
and U24951 (N_24951,N_22792,N_23770);
xnor U24952 (N_24952,N_22232,N_22453);
or U24953 (N_24953,N_22762,N_22357);
nor U24954 (N_24954,N_23066,N_23403);
nand U24955 (N_24955,N_22218,N_23329);
nand U24956 (N_24956,N_23905,N_22256);
xor U24957 (N_24957,N_22594,N_22940);
nand U24958 (N_24958,N_22756,N_22330);
and U24959 (N_24959,N_23741,N_23964);
or U24960 (N_24960,N_22258,N_22436);
or U24961 (N_24961,N_22889,N_23861);
nor U24962 (N_24962,N_22224,N_23040);
or U24963 (N_24963,N_22145,N_22450);
xnor U24964 (N_24964,N_22911,N_23053);
xnor U24965 (N_24965,N_23052,N_22267);
nor U24966 (N_24966,N_22531,N_22637);
nor U24967 (N_24967,N_22993,N_23193);
xnor U24968 (N_24968,N_22892,N_22645);
nor U24969 (N_24969,N_23184,N_23291);
nor U24970 (N_24970,N_22506,N_22981);
and U24971 (N_24971,N_23377,N_22971);
xor U24972 (N_24972,N_22331,N_22285);
nor U24973 (N_24973,N_23576,N_22799);
or U24974 (N_24974,N_23965,N_22448);
or U24975 (N_24975,N_23304,N_23987);
nand U24976 (N_24976,N_22687,N_23872);
or U24977 (N_24977,N_23004,N_23721);
or U24978 (N_24978,N_22941,N_22902);
xor U24979 (N_24979,N_23162,N_23078);
xnor U24980 (N_24980,N_22934,N_22896);
or U24981 (N_24981,N_22770,N_23124);
or U24982 (N_24982,N_23821,N_23289);
nor U24983 (N_24983,N_22164,N_23310);
nand U24984 (N_24984,N_22716,N_22083);
and U24985 (N_24985,N_23266,N_23345);
or U24986 (N_24986,N_22636,N_23538);
nor U24987 (N_24987,N_23670,N_22490);
xnor U24988 (N_24988,N_22223,N_23307);
nor U24989 (N_24989,N_23206,N_23878);
or U24990 (N_24990,N_23848,N_22900);
and U24991 (N_24991,N_23806,N_23093);
nand U24992 (N_24992,N_22193,N_22890);
nand U24993 (N_24993,N_22982,N_22401);
and U24994 (N_24994,N_23748,N_22992);
and U24995 (N_24995,N_22077,N_23384);
or U24996 (N_24996,N_22859,N_22447);
nand U24997 (N_24997,N_23492,N_22154);
and U24998 (N_24998,N_23668,N_22541);
or U24999 (N_24999,N_22029,N_22380);
and U25000 (N_25000,N_23973,N_23175);
and U25001 (N_25001,N_22318,N_23431);
or U25002 (N_25002,N_23468,N_22403);
nor U25003 (N_25003,N_22903,N_23017);
or U25004 (N_25004,N_22213,N_22070);
nand U25005 (N_25005,N_23091,N_23920);
or U25006 (N_25006,N_23523,N_22944);
nor U25007 (N_25007,N_23601,N_22035);
nor U25008 (N_25008,N_23090,N_22115);
and U25009 (N_25009,N_22010,N_23641);
nor U25010 (N_25010,N_22112,N_23688);
xor U25011 (N_25011,N_22460,N_23416);
nor U25012 (N_25012,N_23586,N_23521);
xnor U25013 (N_25013,N_23867,N_23757);
nand U25014 (N_25014,N_22863,N_22400);
and U25015 (N_25015,N_23338,N_22404);
nand U25016 (N_25016,N_23478,N_22687);
nor U25017 (N_25017,N_23152,N_23017);
and U25018 (N_25018,N_23067,N_23004);
or U25019 (N_25019,N_23706,N_22273);
or U25020 (N_25020,N_23064,N_22003);
xor U25021 (N_25021,N_23218,N_22801);
nor U25022 (N_25022,N_23306,N_23516);
xor U25023 (N_25023,N_23806,N_23673);
and U25024 (N_25024,N_23991,N_22427);
nand U25025 (N_25025,N_23928,N_22443);
or U25026 (N_25026,N_22583,N_22600);
and U25027 (N_25027,N_22739,N_23115);
xor U25028 (N_25028,N_23199,N_23017);
nor U25029 (N_25029,N_23681,N_22974);
nor U25030 (N_25030,N_23423,N_22508);
or U25031 (N_25031,N_23163,N_22033);
and U25032 (N_25032,N_23743,N_22009);
nand U25033 (N_25033,N_22153,N_22446);
or U25034 (N_25034,N_23792,N_23839);
and U25035 (N_25035,N_23935,N_22163);
or U25036 (N_25036,N_23239,N_23006);
nor U25037 (N_25037,N_22507,N_22848);
nand U25038 (N_25038,N_23058,N_23779);
nor U25039 (N_25039,N_23936,N_22295);
or U25040 (N_25040,N_22518,N_23148);
and U25041 (N_25041,N_22810,N_23574);
nor U25042 (N_25042,N_23928,N_23454);
nand U25043 (N_25043,N_22390,N_22303);
xnor U25044 (N_25044,N_23957,N_22305);
nor U25045 (N_25045,N_22484,N_23721);
and U25046 (N_25046,N_23716,N_23885);
and U25047 (N_25047,N_22868,N_22908);
xor U25048 (N_25048,N_22542,N_23721);
nand U25049 (N_25049,N_23127,N_22912);
nor U25050 (N_25050,N_23260,N_22693);
xnor U25051 (N_25051,N_23965,N_22681);
xnor U25052 (N_25052,N_22820,N_23893);
nand U25053 (N_25053,N_23382,N_23619);
nor U25054 (N_25054,N_23024,N_23983);
nand U25055 (N_25055,N_22212,N_22653);
xnor U25056 (N_25056,N_23604,N_23736);
nor U25057 (N_25057,N_22687,N_22342);
and U25058 (N_25058,N_23480,N_22786);
nand U25059 (N_25059,N_23190,N_22560);
nand U25060 (N_25060,N_23750,N_23916);
nor U25061 (N_25061,N_22671,N_22869);
nand U25062 (N_25062,N_22183,N_23189);
xor U25063 (N_25063,N_22753,N_22835);
nor U25064 (N_25064,N_22005,N_22486);
xnor U25065 (N_25065,N_23261,N_23756);
xnor U25066 (N_25066,N_22805,N_22632);
nor U25067 (N_25067,N_22272,N_23476);
xor U25068 (N_25068,N_23264,N_22167);
or U25069 (N_25069,N_22677,N_22784);
or U25070 (N_25070,N_22433,N_23319);
nor U25071 (N_25071,N_23341,N_22346);
nand U25072 (N_25072,N_23852,N_23851);
nor U25073 (N_25073,N_23100,N_22282);
xor U25074 (N_25074,N_22936,N_22549);
nor U25075 (N_25075,N_23731,N_22169);
or U25076 (N_25076,N_23841,N_23810);
and U25077 (N_25077,N_23080,N_22251);
xnor U25078 (N_25078,N_22999,N_22362);
nor U25079 (N_25079,N_22060,N_22087);
or U25080 (N_25080,N_23379,N_22582);
and U25081 (N_25081,N_22708,N_22097);
and U25082 (N_25082,N_22162,N_22524);
xor U25083 (N_25083,N_23952,N_22965);
and U25084 (N_25084,N_22464,N_22788);
nor U25085 (N_25085,N_22259,N_22933);
nand U25086 (N_25086,N_23396,N_22109);
nor U25087 (N_25087,N_22819,N_22742);
and U25088 (N_25088,N_23652,N_22132);
nand U25089 (N_25089,N_23675,N_23070);
and U25090 (N_25090,N_22406,N_22348);
nor U25091 (N_25091,N_22346,N_23741);
and U25092 (N_25092,N_23903,N_22223);
xnor U25093 (N_25093,N_22464,N_23358);
and U25094 (N_25094,N_23351,N_23278);
nor U25095 (N_25095,N_22972,N_23227);
nand U25096 (N_25096,N_22170,N_23944);
nor U25097 (N_25097,N_23454,N_23505);
nand U25098 (N_25098,N_22984,N_22062);
nor U25099 (N_25099,N_23417,N_22765);
or U25100 (N_25100,N_22983,N_22318);
nand U25101 (N_25101,N_22897,N_22908);
xnor U25102 (N_25102,N_22864,N_22122);
nor U25103 (N_25103,N_23631,N_23135);
and U25104 (N_25104,N_22064,N_22273);
and U25105 (N_25105,N_23565,N_22422);
nor U25106 (N_25106,N_23678,N_23791);
xnor U25107 (N_25107,N_23449,N_22705);
nor U25108 (N_25108,N_22560,N_23142);
nand U25109 (N_25109,N_22298,N_23368);
xnor U25110 (N_25110,N_23165,N_22937);
nand U25111 (N_25111,N_23100,N_23182);
nor U25112 (N_25112,N_22910,N_23407);
xor U25113 (N_25113,N_23609,N_23909);
nor U25114 (N_25114,N_23596,N_23880);
xor U25115 (N_25115,N_22411,N_23625);
or U25116 (N_25116,N_22951,N_22817);
or U25117 (N_25117,N_23956,N_23547);
nor U25118 (N_25118,N_22594,N_22640);
or U25119 (N_25119,N_22780,N_22378);
and U25120 (N_25120,N_22926,N_22517);
nand U25121 (N_25121,N_22939,N_23284);
nand U25122 (N_25122,N_23128,N_22380);
or U25123 (N_25123,N_23539,N_22020);
and U25124 (N_25124,N_22868,N_23440);
and U25125 (N_25125,N_23458,N_23682);
xnor U25126 (N_25126,N_23055,N_23114);
nor U25127 (N_25127,N_23128,N_22367);
nor U25128 (N_25128,N_22559,N_23359);
nor U25129 (N_25129,N_23333,N_22267);
or U25130 (N_25130,N_22870,N_22227);
nor U25131 (N_25131,N_22436,N_23913);
nand U25132 (N_25132,N_22684,N_22130);
or U25133 (N_25133,N_22312,N_23139);
and U25134 (N_25134,N_22422,N_23471);
or U25135 (N_25135,N_23826,N_23563);
or U25136 (N_25136,N_22555,N_22839);
xnor U25137 (N_25137,N_22394,N_22036);
or U25138 (N_25138,N_23981,N_23680);
nor U25139 (N_25139,N_23962,N_22987);
xor U25140 (N_25140,N_22782,N_23369);
nor U25141 (N_25141,N_22965,N_23629);
and U25142 (N_25142,N_23798,N_23118);
xnor U25143 (N_25143,N_23153,N_22260);
or U25144 (N_25144,N_23139,N_22144);
nand U25145 (N_25145,N_22952,N_22663);
and U25146 (N_25146,N_23293,N_22287);
nand U25147 (N_25147,N_22554,N_22059);
xor U25148 (N_25148,N_23424,N_23955);
nor U25149 (N_25149,N_23888,N_23465);
nor U25150 (N_25150,N_23533,N_23975);
nor U25151 (N_25151,N_23122,N_22086);
and U25152 (N_25152,N_23571,N_23352);
nor U25153 (N_25153,N_23364,N_22574);
xnor U25154 (N_25154,N_23596,N_22820);
nor U25155 (N_25155,N_22556,N_22159);
xor U25156 (N_25156,N_23340,N_23489);
or U25157 (N_25157,N_23752,N_22097);
xnor U25158 (N_25158,N_22300,N_23570);
and U25159 (N_25159,N_23890,N_23986);
xnor U25160 (N_25160,N_23807,N_23292);
xor U25161 (N_25161,N_22187,N_22132);
nand U25162 (N_25162,N_22911,N_23382);
xnor U25163 (N_25163,N_22547,N_23501);
and U25164 (N_25164,N_22549,N_22252);
xnor U25165 (N_25165,N_23741,N_23427);
xor U25166 (N_25166,N_22144,N_22104);
and U25167 (N_25167,N_23378,N_22228);
nor U25168 (N_25168,N_22065,N_23884);
and U25169 (N_25169,N_23406,N_22288);
or U25170 (N_25170,N_22234,N_23992);
nor U25171 (N_25171,N_23823,N_22385);
and U25172 (N_25172,N_23381,N_23622);
and U25173 (N_25173,N_23572,N_22365);
and U25174 (N_25174,N_23778,N_23431);
and U25175 (N_25175,N_22411,N_22850);
and U25176 (N_25176,N_22925,N_23735);
nor U25177 (N_25177,N_23452,N_23855);
or U25178 (N_25178,N_23815,N_22670);
nand U25179 (N_25179,N_22668,N_23072);
xor U25180 (N_25180,N_23884,N_23419);
xnor U25181 (N_25181,N_22968,N_22446);
and U25182 (N_25182,N_22768,N_22740);
and U25183 (N_25183,N_23793,N_22240);
and U25184 (N_25184,N_23025,N_23609);
nand U25185 (N_25185,N_22996,N_22523);
nand U25186 (N_25186,N_23856,N_22502);
xor U25187 (N_25187,N_23585,N_23793);
nor U25188 (N_25188,N_23382,N_23047);
xor U25189 (N_25189,N_22581,N_22528);
nor U25190 (N_25190,N_22586,N_22561);
nand U25191 (N_25191,N_22066,N_22248);
nor U25192 (N_25192,N_23281,N_23479);
xor U25193 (N_25193,N_22645,N_22776);
nor U25194 (N_25194,N_23966,N_23372);
nand U25195 (N_25195,N_23568,N_22394);
or U25196 (N_25196,N_23635,N_23922);
xor U25197 (N_25197,N_22456,N_23910);
nor U25198 (N_25198,N_23936,N_23925);
nor U25199 (N_25199,N_23961,N_23989);
or U25200 (N_25200,N_23378,N_22976);
nand U25201 (N_25201,N_22557,N_22606);
or U25202 (N_25202,N_22244,N_22697);
or U25203 (N_25203,N_23764,N_22618);
nand U25204 (N_25204,N_22996,N_22738);
or U25205 (N_25205,N_23962,N_23144);
xor U25206 (N_25206,N_22070,N_23433);
xor U25207 (N_25207,N_23005,N_23298);
and U25208 (N_25208,N_22271,N_22992);
xor U25209 (N_25209,N_22709,N_22876);
and U25210 (N_25210,N_22146,N_23830);
xor U25211 (N_25211,N_22907,N_22497);
or U25212 (N_25212,N_23824,N_22740);
nor U25213 (N_25213,N_22774,N_23286);
and U25214 (N_25214,N_23981,N_23392);
nor U25215 (N_25215,N_22565,N_23833);
xor U25216 (N_25216,N_23892,N_22919);
xor U25217 (N_25217,N_23971,N_23945);
or U25218 (N_25218,N_22298,N_22769);
xnor U25219 (N_25219,N_22331,N_23686);
or U25220 (N_25220,N_23126,N_22436);
and U25221 (N_25221,N_23154,N_22843);
or U25222 (N_25222,N_23459,N_23340);
or U25223 (N_25223,N_22055,N_23103);
nand U25224 (N_25224,N_23493,N_23292);
or U25225 (N_25225,N_22500,N_23881);
and U25226 (N_25226,N_23163,N_22849);
nor U25227 (N_25227,N_22551,N_23020);
xor U25228 (N_25228,N_22885,N_22992);
nor U25229 (N_25229,N_23651,N_23734);
or U25230 (N_25230,N_23697,N_23017);
nor U25231 (N_25231,N_22098,N_23904);
nand U25232 (N_25232,N_22592,N_23764);
xor U25233 (N_25233,N_22734,N_22617);
or U25234 (N_25234,N_23961,N_23680);
and U25235 (N_25235,N_22734,N_22570);
xor U25236 (N_25236,N_23218,N_22485);
or U25237 (N_25237,N_23285,N_23742);
and U25238 (N_25238,N_23746,N_22520);
xor U25239 (N_25239,N_22554,N_23434);
and U25240 (N_25240,N_23240,N_23113);
or U25241 (N_25241,N_22295,N_23120);
or U25242 (N_25242,N_22517,N_23843);
or U25243 (N_25243,N_23985,N_22408);
nand U25244 (N_25244,N_22810,N_23320);
nor U25245 (N_25245,N_23748,N_22807);
and U25246 (N_25246,N_23429,N_23416);
xor U25247 (N_25247,N_22406,N_22557);
and U25248 (N_25248,N_22144,N_23434);
nand U25249 (N_25249,N_23001,N_22443);
and U25250 (N_25250,N_22646,N_22515);
nor U25251 (N_25251,N_22692,N_22775);
and U25252 (N_25252,N_23583,N_23461);
nor U25253 (N_25253,N_22084,N_23436);
and U25254 (N_25254,N_23612,N_23819);
nor U25255 (N_25255,N_22815,N_23147);
or U25256 (N_25256,N_22530,N_22984);
or U25257 (N_25257,N_22146,N_22728);
or U25258 (N_25258,N_23773,N_23768);
and U25259 (N_25259,N_22194,N_22737);
nor U25260 (N_25260,N_22666,N_22445);
or U25261 (N_25261,N_22451,N_22293);
nor U25262 (N_25262,N_22024,N_23391);
nor U25263 (N_25263,N_22818,N_23869);
xnor U25264 (N_25264,N_23408,N_23220);
and U25265 (N_25265,N_23689,N_23294);
and U25266 (N_25266,N_22453,N_22422);
nand U25267 (N_25267,N_23201,N_23949);
or U25268 (N_25268,N_22344,N_22170);
nand U25269 (N_25269,N_22303,N_23866);
or U25270 (N_25270,N_22800,N_23554);
nor U25271 (N_25271,N_23405,N_22280);
nand U25272 (N_25272,N_22797,N_22580);
or U25273 (N_25273,N_22700,N_23748);
xor U25274 (N_25274,N_23656,N_23723);
or U25275 (N_25275,N_23989,N_22122);
and U25276 (N_25276,N_23270,N_23205);
nand U25277 (N_25277,N_22225,N_23559);
and U25278 (N_25278,N_22001,N_22414);
nand U25279 (N_25279,N_22947,N_22633);
xor U25280 (N_25280,N_23516,N_22114);
xnor U25281 (N_25281,N_23598,N_22819);
and U25282 (N_25282,N_22272,N_22441);
nand U25283 (N_25283,N_23259,N_23084);
or U25284 (N_25284,N_23374,N_23054);
xnor U25285 (N_25285,N_22270,N_23735);
nand U25286 (N_25286,N_23277,N_23944);
xnor U25287 (N_25287,N_23405,N_23475);
or U25288 (N_25288,N_22779,N_23421);
nor U25289 (N_25289,N_23736,N_22715);
nand U25290 (N_25290,N_23151,N_22374);
and U25291 (N_25291,N_22067,N_22636);
and U25292 (N_25292,N_23844,N_23177);
or U25293 (N_25293,N_23644,N_23278);
nor U25294 (N_25294,N_22862,N_23792);
xnor U25295 (N_25295,N_22941,N_23464);
nor U25296 (N_25296,N_22267,N_22425);
or U25297 (N_25297,N_23943,N_23501);
nand U25298 (N_25298,N_23841,N_23586);
xnor U25299 (N_25299,N_22876,N_23641);
or U25300 (N_25300,N_23823,N_22846);
and U25301 (N_25301,N_23817,N_22418);
nand U25302 (N_25302,N_23892,N_22539);
and U25303 (N_25303,N_23784,N_23969);
nand U25304 (N_25304,N_22871,N_23023);
xor U25305 (N_25305,N_22161,N_22571);
nand U25306 (N_25306,N_23587,N_22695);
and U25307 (N_25307,N_22587,N_23899);
nor U25308 (N_25308,N_23807,N_22778);
or U25309 (N_25309,N_22380,N_23047);
nor U25310 (N_25310,N_23663,N_23496);
nor U25311 (N_25311,N_22213,N_23925);
or U25312 (N_25312,N_22479,N_23606);
or U25313 (N_25313,N_22649,N_23378);
xor U25314 (N_25314,N_23233,N_23870);
nor U25315 (N_25315,N_22550,N_23238);
nor U25316 (N_25316,N_23809,N_23570);
nand U25317 (N_25317,N_23912,N_22440);
nor U25318 (N_25318,N_23827,N_23942);
nor U25319 (N_25319,N_22825,N_23812);
nand U25320 (N_25320,N_23795,N_22335);
nand U25321 (N_25321,N_22638,N_22295);
and U25322 (N_25322,N_23114,N_22675);
or U25323 (N_25323,N_22852,N_22818);
or U25324 (N_25324,N_22121,N_22006);
or U25325 (N_25325,N_22820,N_23376);
xor U25326 (N_25326,N_22818,N_23062);
nand U25327 (N_25327,N_22238,N_22894);
xor U25328 (N_25328,N_22263,N_23031);
and U25329 (N_25329,N_22471,N_22450);
or U25330 (N_25330,N_23525,N_23170);
xor U25331 (N_25331,N_22396,N_23166);
and U25332 (N_25332,N_22851,N_23544);
xor U25333 (N_25333,N_23852,N_22553);
nand U25334 (N_25334,N_23062,N_23208);
nand U25335 (N_25335,N_22016,N_23616);
nand U25336 (N_25336,N_23290,N_22286);
and U25337 (N_25337,N_22352,N_23662);
nor U25338 (N_25338,N_22082,N_22217);
xor U25339 (N_25339,N_22562,N_22337);
nand U25340 (N_25340,N_22350,N_22376);
or U25341 (N_25341,N_22757,N_23964);
nor U25342 (N_25342,N_22623,N_22732);
nand U25343 (N_25343,N_22699,N_22439);
or U25344 (N_25344,N_23826,N_22955);
nand U25345 (N_25345,N_23771,N_23768);
or U25346 (N_25346,N_22342,N_23011);
or U25347 (N_25347,N_22887,N_22190);
nor U25348 (N_25348,N_23153,N_22590);
xnor U25349 (N_25349,N_23524,N_22168);
nand U25350 (N_25350,N_23847,N_23886);
nor U25351 (N_25351,N_23380,N_23782);
nand U25352 (N_25352,N_22259,N_23766);
and U25353 (N_25353,N_22492,N_23647);
and U25354 (N_25354,N_23002,N_23988);
and U25355 (N_25355,N_23995,N_22273);
xor U25356 (N_25356,N_22628,N_22541);
nor U25357 (N_25357,N_23297,N_22334);
nand U25358 (N_25358,N_22877,N_23240);
nand U25359 (N_25359,N_22358,N_23949);
xnor U25360 (N_25360,N_23078,N_22186);
xnor U25361 (N_25361,N_23859,N_23061);
nand U25362 (N_25362,N_22709,N_22300);
xor U25363 (N_25363,N_23806,N_23099);
xnor U25364 (N_25364,N_22266,N_23571);
or U25365 (N_25365,N_23101,N_23501);
nor U25366 (N_25366,N_23625,N_22793);
or U25367 (N_25367,N_23520,N_23673);
or U25368 (N_25368,N_22093,N_22069);
xnor U25369 (N_25369,N_23934,N_22510);
xnor U25370 (N_25370,N_23637,N_23838);
or U25371 (N_25371,N_23146,N_23235);
nor U25372 (N_25372,N_22408,N_22521);
nor U25373 (N_25373,N_23496,N_22739);
or U25374 (N_25374,N_23641,N_23045);
nand U25375 (N_25375,N_23922,N_23662);
or U25376 (N_25376,N_23913,N_23551);
or U25377 (N_25377,N_23139,N_23469);
or U25378 (N_25378,N_22557,N_23313);
nand U25379 (N_25379,N_22631,N_22231);
nand U25380 (N_25380,N_23248,N_22276);
nor U25381 (N_25381,N_23652,N_23332);
or U25382 (N_25382,N_23802,N_22401);
nand U25383 (N_25383,N_23106,N_23671);
and U25384 (N_25384,N_23973,N_23631);
nor U25385 (N_25385,N_23097,N_22784);
or U25386 (N_25386,N_23096,N_23552);
and U25387 (N_25387,N_23349,N_23564);
or U25388 (N_25388,N_22185,N_23568);
nor U25389 (N_25389,N_23466,N_22930);
nand U25390 (N_25390,N_22635,N_23779);
or U25391 (N_25391,N_22215,N_23744);
xor U25392 (N_25392,N_22985,N_22683);
and U25393 (N_25393,N_22408,N_23193);
nor U25394 (N_25394,N_23366,N_22541);
nand U25395 (N_25395,N_22324,N_23812);
and U25396 (N_25396,N_23902,N_22572);
nand U25397 (N_25397,N_22376,N_23656);
nand U25398 (N_25398,N_23346,N_22232);
xor U25399 (N_25399,N_22077,N_23947);
nand U25400 (N_25400,N_22830,N_23087);
or U25401 (N_25401,N_23176,N_22649);
nand U25402 (N_25402,N_22891,N_22292);
nor U25403 (N_25403,N_23090,N_22564);
or U25404 (N_25404,N_22804,N_22641);
nor U25405 (N_25405,N_23584,N_22122);
or U25406 (N_25406,N_23112,N_23398);
or U25407 (N_25407,N_23229,N_22009);
and U25408 (N_25408,N_22428,N_23205);
xor U25409 (N_25409,N_22945,N_23144);
and U25410 (N_25410,N_23115,N_23792);
nand U25411 (N_25411,N_22044,N_23890);
and U25412 (N_25412,N_22803,N_22620);
xor U25413 (N_25413,N_23142,N_23930);
xor U25414 (N_25414,N_22085,N_23760);
and U25415 (N_25415,N_23341,N_22121);
xnor U25416 (N_25416,N_23015,N_22713);
xor U25417 (N_25417,N_23925,N_22881);
or U25418 (N_25418,N_23502,N_23891);
and U25419 (N_25419,N_23940,N_23008);
or U25420 (N_25420,N_22575,N_22028);
nand U25421 (N_25421,N_23771,N_22682);
xor U25422 (N_25422,N_23592,N_22289);
and U25423 (N_25423,N_23024,N_23942);
and U25424 (N_25424,N_22490,N_23779);
nor U25425 (N_25425,N_22217,N_22035);
and U25426 (N_25426,N_23192,N_22041);
xnor U25427 (N_25427,N_22864,N_23320);
or U25428 (N_25428,N_23389,N_22139);
nor U25429 (N_25429,N_22036,N_23171);
nand U25430 (N_25430,N_22065,N_23807);
xor U25431 (N_25431,N_23735,N_22948);
or U25432 (N_25432,N_23059,N_23463);
or U25433 (N_25433,N_23964,N_23550);
nand U25434 (N_25434,N_22072,N_22231);
and U25435 (N_25435,N_22957,N_22920);
or U25436 (N_25436,N_22189,N_22525);
xor U25437 (N_25437,N_23155,N_23866);
nand U25438 (N_25438,N_23198,N_22291);
nor U25439 (N_25439,N_23375,N_23278);
nor U25440 (N_25440,N_23691,N_22249);
nor U25441 (N_25441,N_22280,N_22804);
xnor U25442 (N_25442,N_23916,N_22078);
nand U25443 (N_25443,N_22246,N_22089);
xor U25444 (N_25444,N_22882,N_23726);
nor U25445 (N_25445,N_23431,N_23438);
and U25446 (N_25446,N_23963,N_22007);
xnor U25447 (N_25447,N_23147,N_22116);
nand U25448 (N_25448,N_22507,N_22309);
nand U25449 (N_25449,N_23466,N_23760);
xor U25450 (N_25450,N_22417,N_23307);
and U25451 (N_25451,N_23693,N_22694);
or U25452 (N_25452,N_23454,N_22278);
nand U25453 (N_25453,N_23026,N_22822);
nand U25454 (N_25454,N_22054,N_23225);
and U25455 (N_25455,N_22860,N_23926);
xnor U25456 (N_25456,N_22154,N_22388);
or U25457 (N_25457,N_23806,N_22588);
nor U25458 (N_25458,N_22250,N_22174);
and U25459 (N_25459,N_22891,N_23736);
or U25460 (N_25460,N_23229,N_23455);
nand U25461 (N_25461,N_22598,N_22675);
xor U25462 (N_25462,N_22182,N_22916);
or U25463 (N_25463,N_23610,N_22370);
nand U25464 (N_25464,N_23348,N_23046);
xor U25465 (N_25465,N_23660,N_23589);
xor U25466 (N_25466,N_22882,N_22216);
or U25467 (N_25467,N_22288,N_22771);
nor U25468 (N_25468,N_23518,N_22087);
nand U25469 (N_25469,N_22570,N_22732);
nor U25470 (N_25470,N_23331,N_23682);
nor U25471 (N_25471,N_22283,N_23622);
and U25472 (N_25472,N_23961,N_23273);
or U25473 (N_25473,N_22737,N_22939);
nand U25474 (N_25474,N_23249,N_23814);
xor U25475 (N_25475,N_23146,N_22204);
and U25476 (N_25476,N_23583,N_23596);
or U25477 (N_25477,N_23725,N_22721);
nand U25478 (N_25478,N_22431,N_23176);
xor U25479 (N_25479,N_22552,N_23167);
nand U25480 (N_25480,N_23383,N_23748);
xor U25481 (N_25481,N_23048,N_22305);
nand U25482 (N_25482,N_23947,N_22046);
xnor U25483 (N_25483,N_23035,N_23946);
nor U25484 (N_25484,N_23880,N_22699);
xnor U25485 (N_25485,N_23828,N_23392);
xnor U25486 (N_25486,N_22632,N_22124);
nand U25487 (N_25487,N_23429,N_22089);
and U25488 (N_25488,N_22463,N_22552);
nand U25489 (N_25489,N_23263,N_22854);
xor U25490 (N_25490,N_23401,N_22429);
nand U25491 (N_25491,N_23131,N_23894);
nor U25492 (N_25492,N_22731,N_22684);
or U25493 (N_25493,N_22468,N_23504);
and U25494 (N_25494,N_23109,N_22080);
nand U25495 (N_25495,N_23133,N_23073);
or U25496 (N_25496,N_22247,N_23253);
or U25497 (N_25497,N_22516,N_23198);
or U25498 (N_25498,N_22110,N_22918);
nor U25499 (N_25499,N_23563,N_22798);
nor U25500 (N_25500,N_22362,N_22665);
nand U25501 (N_25501,N_23801,N_23806);
nand U25502 (N_25502,N_22269,N_23242);
xnor U25503 (N_25503,N_22301,N_23060);
or U25504 (N_25504,N_23770,N_23813);
or U25505 (N_25505,N_23264,N_23236);
and U25506 (N_25506,N_22641,N_22860);
and U25507 (N_25507,N_22896,N_22172);
or U25508 (N_25508,N_22755,N_23394);
xor U25509 (N_25509,N_22676,N_23303);
or U25510 (N_25510,N_22028,N_23489);
nor U25511 (N_25511,N_22812,N_22794);
nor U25512 (N_25512,N_22977,N_22117);
nand U25513 (N_25513,N_23352,N_22750);
xor U25514 (N_25514,N_23482,N_23253);
xnor U25515 (N_25515,N_22747,N_23654);
or U25516 (N_25516,N_23497,N_22919);
or U25517 (N_25517,N_22395,N_23112);
nor U25518 (N_25518,N_22871,N_23799);
nand U25519 (N_25519,N_22471,N_23032);
xnor U25520 (N_25520,N_22360,N_23901);
nor U25521 (N_25521,N_23069,N_23796);
and U25522 (N_25522,N_23978,N_22749);
xnor U25523 (N_25523,N_23445,N_22709);
nand U25524 (N_25524,N_22660,N_22044);
xnor U25525 (N_25525,N_23614,N_22972);
and U25526 (N_25526,N_23866,N_23264);
or U25527 (N_25527,N_23530,N_22908);
or U25528 (N_25528,N_23610,N_23785);
xnor U25529 (N_25529,N_23886,N_22360);
xor U25530 (N_25530,N_23499,N_22975);
xor U25531 (N_25531,N_23759,N_23417);
nand U25532 (N_25532,N_23833,N_22222);
nor U25533 (N_25533,N_23478,N_23667);
nand U25534 (N_25534,N_23788,N_22543);
or U25535 (N_25535,N_23475,N_22253);
or U25536 (N_25536,N_22129,N_23535);
nor U25537 (N_25537,N_23597,N_22873);
or U25538 (N_25538,N_23902,N_23176);
xor U25539 (N_25539,N_22895,N_23403);
or U25540 (N_25540,N_22720,N_22006);
or U25541 (N_25541,N_22485,N_23820);
xor U25542 (N_25542,N_22480,N_22580);
or U25543 (N_25543,N_22858,N_22156);
nor U25544 (N_25544,N_22662,N_22845);
or U25545 (N_25545,N_23659,N_23581);
nand U25546 (N_25546,N_23040,N_23219);
or U25547 (N_25547,N_23987,N_23233);
and U25548 (N_25548,N_22836,N_22635);
and U25549 (N_25549,N_23584,N_23237);
or U25550 (N_25550,N_23387,N_23526);
nand U25551 (N_25551,N_23347,N_23121);
or U25552 (N_25552,N_22692,N_23082);
and U25553 (N_25553,N_23213,N_23432);
xor U25554 (N_25554,N_22123,N_22920);
or U25555 (N_25555,N_22504,N_22578);
or U25556 (N_25556,N_22985,N_22025);
nand U25557 (N_25557,N_22485,N_23548);
or U25558 (N_25558,N_22708,N_23359);
nor U25559 (N_25559,N_22263,N_23395);
nor U25560 (N_25560,N_22969,N_22015);
xor U25561 (N_25561,N_23174,N_23035);
and U25562 (N_25562,N_22560,N_22572);
or U25563 (N_25563,N_22618,N_22527);
xor U25564 (N_25564,N_22534,N_23097);
xor U25565 (N_25565,N_23780,N_23268);
or U25566 (N_25566,N_23400,N_22327);
nor U25567 (N_25567,N_22254,N_23356);
xnor U25568 (N_25568,N_23904,N_23246);
nor U25569 (N_25569,N_22789,N_23119);
xor U25570 (N_25570,N_22975,N_23536);
xnor U25571 (N_25571,N_23074,N_22573);
nand U25572 (N_25572,N_22073,N_22368);
nor U25573 (N_25573,N_22156,N_22533);
and U25574 (N_25574,N_23652,N_22602);
and U25575 (N_25575,N_22156,N_23076);
nand U25576 (N_25576,N_23928,N_23031);
nor U25577 (N_25577,N_23236,N_23829);
nand U25578 (N_25578,N_23224,N_23317);
and U25579 (N_25579,N_23495,N_22850);
nor U25580 (N_25580,N_22631,N_23550);
xor U25581 (N_25581,N_22558,N_23393);
and U25582 (N_25582,N_22266,N_23143);
and U25583 (N_25583,N_22831,N_22658);
nor U25584 (N_25584,N_22160,N_23770);
nand U25585 (N_25585,N_23880,N_23316);
nand U25586 (N_25586,N_22080,N_23186);
xor U25587 (N_25587,N_23251,N_23426);
nor U25588 (N_25588,N_22974,N_23096);
nor U25589 (N_25589,N_22278,N_22636);
xnor U25590 (N_25590,N_23310,N_23855);
or U25591 (N_25591,N_22216,N_23475);
nor U25592 (N_25592,N_23923,N_23491);
and U25593 (N_25593,N_23648,N_22084);
nand U25594 (N_25594,N_23705,N_22699);
or U25595 (N_25595,N_22583,N_23194);
xnor U25596 (N_25596,N_22821,N_23571);
xnor U25597 (N_25597,N_23370,N_23257);
or U25598 (N_25598,N_23499,N_23221);
xor U25599 (N_25599,N_22248,N_23098);
xor U25600 (N_25600,N_22152,N_23017);
and U25601 (N_25601,N_22981,N_23500);
nor U25602 (N_25602,N_23416,N_23708);
and U25603 (N_25603,N_23544,N_23710);
nand U25604 (N_25604,N_23519,N_22355);
and U25605 (N_25605,N_23117,N_23848);
nand U25606 (N_25606,N_22849,N_23034);
or U25607 (N_25607,N_22482,N_23672);
nor U25608 (N_25608,N_22402,N_23032);
and U25609 (N_25609,N_23594,N_23235);
nand U25610 (N_25610,N_23376,N_22261);
nor U25611 (N_25611,N_23638,N_23169);
nand U25612 (N_25612,N_22543,N_22912);
nand U25613 (N_25613,N_22919,N_22694);
nor U25614 (N_25614,N_23479,N_22422);
and U25615 (N_25615,N_23092,N_22146);
xnor U25616 (N_25616,N_23759,N_22132);
xnor U25617 (N_25617,N_23070,N_22541);
and U25618 (N_25618,N_22270,N_22066);
nor U25619 (N_25619,N_23854,N_23131);
xnor U25620 (N_25620,N_23097,N_22008);
and U25621 (N_25621,N_22732,N_23788);
nand U25622 (N_25622,N_23123,N_22703);
and U25623 (N_25623,N_22157,N_23864);
or U25624 (N_25624,N_22763,N_22705);
nand U25625 (N_25625,N_23608,N_22760);
xor U25626 (N_25626,N_23262,N_23378);
nand U25627 (N_25627,N_23419,N_23885);
nor U25628 (N_25628,N_23494,N_23932);
nand U25629 (N_25629,N_23143,N_23668);
nand U25630 (N_25630,N_22536,N_23517);
nor U25631 (N_25631,N_22948,N_23146);
or U25632 (N_25632,N_22060,N_23578);
and U25633 (N_25633,N_23105,N_22430);
nand U25634 (N_25634,N_23998,N_22290);
xnor U25635 (N_25635,N_23833,N_23706);
xor U25636 (N_25636,N_22285,N_22569);
nor U25637 (N_25637,N_22729,N_22472);
and U25638 (N_25638,N_22395,N_22026);
nand U25639 (N_25639,N_23368,N_23367);
xnor U25640 (N_25640,N_23769,N_23891);
xnor U25641 (N_25641,N_22340,N_22707);
xnor U25642 (N_25642,N_23354,N_22450);
xor U25643 (N_25643,N_22506,N_23046);
and U25644 (N_25644,N_23312,N_22595);
and U25645 (N_25645,N_22620,N_23086);
nand U25646 (N_25646,N_23812,N_22368);
xor U25647 (N_25647,N_22906,N_23267);
nand U25648 (N_25648,N_23706,N_23101);
nor U25649 (N_25649,N_22609,N_23981);
nand U25650 (N_25650,N_22657,N_22992);
and U25651 (N_25651,N_23889,N_23469);
xor U25652 (N_25652,N_23660,N_23015);
and U25653 (N_25653,N_23479,N_22195);
and U25654 (N_25654,N_22315,N_23820);
or U25655 (N_25655,N_23824,N_23342);
nand U25656 (N_25656,N_22450,N_23025);
xnor U25657 (N_25657,N_22035,N_22776);
nand U25658 (N_25658,N_22802,N_23835);
or U25659 (N_25659,N_22503,N_23183);
nand U25660 (N_25660,N_22740,N_23177);
nor U25661 (N_25661,N_22435,N_23291);
xnor U25662 (N_25662,N_23338,N_22316);
and U25663 (N_25663,N_23743,N_23579);
nor U25664 (N_25664,N_23769,N_22199);
xnor U25665 (N_25665,N_23862,N_23394);
or U25666 (N_25666,N_22889,N_23949);
nand U25667 (N_25667,N_22889,N_23921);
xnor U25668 (N_25668,N_22280,N_22065);
xnor U25669 (N_25669,N_23360,N_23621);
nand U25670 (N_25670,N_23796,N_22762);
and U25671 (N_25671,N_22639,N_22041);
xnor U25672 (N_25672,N_23792,N_23990);
or U25673 (N_25673,N_23470,N_23237);
nand U25674 (N_25674,N_23366,N_22836);
and U25675 (N_25675,N_22447,N_22985);
nor U25676 (N_25676,N_23833,N_22770);
and U25677 (N_25677,N_22287,N_22455);
nor U25678 (N_25678,N_22887,N_23866);
nor U25679 (N_25679,N_22409,N_23665);
xor U25680 (N_25680,N_22800,N_23181);
xnor U25681 (N_25681,N_22758,N_23779);
or U25682 (N_25682,N_23456,N_23053);
nor U25683 (N_25683,N_22008,N_23968);
and U25684 (N_25684,N_23135,N_22171);
nor U25685 (N_25685,N_23730,N_23128);
or U25686 (N_25686,N_22325,N_23812);
xnor U25687 (N_25687,N_23562,N_22857);
or U25688 (N_25688,N_22844,N_23703);
nand U25689 (N_25689,N_23596,N_23059);
and U25690 (N_25690,N_23898,N_22069);
xor U25691 (N_25691,N_22056,N_22020);
xnor U25692 (N_25692,N_22189,N_22162);
xor U25693 (N_25693,N_22866,N_22698);
or U25694 (N_25694,N_22297,N_22959);
xor U25695 (N_25695,N_23564,N_22209);
and U25696 (N_25696,N_23679,N_22734);
or U25697 (N_25697,N_23686,N_23672);
nand U25698 (N_25698,N_22164,N_23420);
nor U25699 (N_25699,N_22071,N_22140);
and U25700 (N_25700,N_22528,N_22941);
nor U25701 (N_25701,N_22990,N_23862);
xnor U25702 (N_25702,N_23865,N_23434);
xnor U25703 (N_25703,N_22236,N_23619);
or U25704 (N_25704,N_22072,N_22089);
or U25705 (N_25705,N_22232,N_22144);
xor U25706 (N_25706,N_22083,N_23463);
nand U25707 (N_25707,N_23293,N_23491);
or U25708 (N_25708,N_23513,N_23246);
and U25709 (N_25709,N_22302,N_22459);
nand U25710 (N_25710,N_23818,N_23379);
or U25711 (N_25711,N_22985,N_22443);
xor U25712 (N_25712,N_22352,N_22127);
xnor U25713 (N_25713,N_23961,N_22389);
nand U25714 (N_25714,N_23549,N_23282);
and U25715 (N_25715,N_23337,N_23891);
nand U25716 (N_25716,N_23478,N_23265);
xnor U25717 (N_25717,N_22264,N_23642);
or U25718 (N_25718,N_22930,N_22363);
or U25719 (N_25719,N_23311,N_22956);
or U25720 (N_25720,N_22110,N_22806);
nand U25721 (N_25721,N_23582,N_22678);
nor U25722 (N_25722,N_22127,N_23865);
and U25723 (N_25723,N_23920,N_23414);
xnor U25724 (N_25724,N_23631,N_22911);
or U25725 (N_25725,N_22719,N_23906);
and U25726 (N_25726,N_22553,N_23136);
and U25727 (N_25727,N_23272,N_23128);
and U25728 (N_25728,N_22790,N_22116);
nand U25729 (N_25729,N_22918,N_23127);
or U25730 (N_25730,N_23083,N_23681);
and U25731 (N_25731,N_23897,N_23595);
or U25732 (N_25732,N_23440,N_23143);
xor U25733 (N_25733,N_22097,N_23497);
and U25734 (N_25734,N_23755,N_23280);
and U25735 (N_25735,N_23927,N_22028);
nor U25736 (N_25736,N_22305,N_22572);
or U25737 (N_25737,N_23825,N_23434);
nand U25738 (N_25738,N_22668,N_23363);
or U25739 (N_25739,N_23037,N_22269);
nor U25740 (N_25740,N_22469,N_22502);
and U25741 (N_25741,N_22583,N_23813);
and U25742 (N_25742,N_22094,N_23622);
and U25743 (N_25743,N_23820,N_22832);
or U25744 (N_25744,N_23002,N_22603);
nand U25745 (N_25745,N_22481,N_22727);
nor U25746 (N_25746,N_22752,N_22420);
nand U25747 (N_25747,N_22841,N_22029);
or U25748 (N_25748,N_22891,N_23657);
xnor U25749 (N_25749,N_23884,N_22762);
or U25750 (N_25750,N_23892,N_22223);
nor U25751 (N_25751,N_23783,N_23980);
xnor U25752 (N_25752,N_23875,N_22430);
or U25753 (N_25753,N_23630,N_22551);
or U25754 (N_25754,N_23333,N_22811);
nor U25755 (N_25755,N_22819,N_23133);
or U25756 (N_25756,N_22267,N_22259);
xor U25757 (N_25757,N_23698,N_23690);
nor U25758 (N_25758,N_23531,N_23400);
and U25759 (N_25759,N_22550,N_23355);
nand U25760 (N_25760,N_23895,N_22343);
and U25761 (N_25761,N_23144,N_22560);
xor U25762 (N_25762,N_23366,N_22368);
or U25763 (N_25763,N_23594,N_22815);
or U25764 (N_25764,N_23932,N_23165);
nor U25765 (N_25765,N_23615,N_22023);
nor U25766 (N_25766,N_23815,N_22401);
or U25767 (N_25767,N_22481,N_22596);
nor U25768 (N_25768,N_23778,N_22409);
nor U25769 (N_25769,N_23285,N_22902);
xor U25770 (N_25770,N_23915,N_22696);
and U25771 (N_25771,N_22080,N_23426);
xor U25772 (N_25772,N_23613,N_22108);
nand U25773 (N_25773,N_23495,N_22334);
xnor U25774 (N_25774,N_23026,N_22376);
or U25775 (N_25775,N_23973,N_22926);
nor U25776 (N_25776,N_23000,N_23347);
or U25777 (N_25777,N_23935,N_23518);
or U25778 (N_25778,N_22899,N_23433);
xnor U25779 (N_25779,N_23957,N_23663);
and U25780 (N_25780,N_23150,N_22340);
nor U25781 (N_25781,N_22557,N_23736);
and U25782 (N_25782,N_23049,N_23160);
nand U25783 (N_25783,N_22384,N_22481);
nand U25784 (N_25784,N_22484,N_23500);
xnor U25785 (N_25785,N_22428,N_23218);
or U25786 (N_25786,N_22705,N_23935);
and U25787 (N_25787,N_23798,N_22568);
nand U25788 (N_25788,N_22403,N_22910);
and U25789 (N_25789,N_23684,N_22318);
and U25790 (N_25790,N_23748,N_23257);
xnor U25791 (N_25791,N_22356,N_23036);
or U25792 (N_25792,N_22683,N_23134);
or U25793 (N_25793,N_23184,N_23507);
nand U25794 (N_25794,N_22222,N_22141);
and U25795 (N_25795,N_22831,N_22367);
and U25796 (N_25796,N_23963,N_23049);
nor U25797 (N_25797,N_23427,N_22325);
xnor U25798 (N_25798,N_22009,N_22915);
nand U25799 (N_25799,N_22815,N_22084);
and U25800 (N_25800,N_22874,N_23765);
nor U25801 (N_25801,N_22145,N_23108);
nor U25802 (N_25802,N_22948,N_22684);
xor U25803 (N_25803,N_23622,N_22772);
nand U25804 (N_25804,N_23966,N_22694);
nor U25805 (N_25805,N_23577,N_22094);
nand U25806 (N_25806,N_22765,N_23326);
xnor U25807 (N_25807,N_23297,N_23652);
or U25808 (N_25808,N_22367,N_22718);
nor U25809 (N_25809,N_22138,N_23596);
and U25810 (N_25810,N_23618,N_23394);
or U25811 (N_25811,N_23728,N_22892);
and U25812 (N_25812,N_22888,N_22825);
xnor U25813 (N_25813,N_23129,N_22138);
nand U25814 (N_25814,N_23309,N_22979);
nand U25815 (N_25815,N_22398,N_22737);
xor U25816 (N_25816,N_22993,N_23452);
nand U25817 (N_25817,N_23433,N_23240);
nor U25818 (N_25818,N_22805,N_22030);
and U25819 (N_25819,N_23059,N_22923);
or U25820 (N_25820,N_22524,N_23236);
and U25821 (N_25821,N_23902,N_23869);
nor U25822 (N_25822,N_22680,N_22708);
or U25823 (N_25823,N_22271,N_23716);
nand U25824 (N_25824,N_23963,N_22470);
nor U25825 (N_25825,N_23814,N_22682);
or U25826 (N_25826,N_23127,N_23454);
and U25827 (N_25827,N_23896,N_23145);
xnor U25828 (N_25828,N_22991,N_23546);
nand U25829 (N_25829,N_23243,N_23570);
xor U25830 (N_25830,N_22047,N_23468);
nor U25831 (N_25831,N_23923,N_22972);
nand U25832 (N_25832,N_22934,N_23339);
or U25833 (N_25833,N_22754,N_22362);
nor U25834 (N_25834,N_22741,N_23565);
and U25835 (N_25835,N_23697,N_23450);
nor U25836 (N_25836,N_22802,N_22669);
and U25837 (N_25837,N_22807,N_23074);
or U25838 (N_25838,N_22533,N_22027);
and U25839 (N_25839,N_23717,N_22191);
or U25840 (N_25840,N_23625,N_22382);
or U25841 (N_25841,N_23280,N_22657);
xnor U25842 (N_25842,N_23813,N_23187);
xor U25843 (N_25843,N_23937,N_23593);
nand U25844 (N_25844,N_23997,N_23003);
and U25845 (N_25845,N_23817,N_22488);
nand U25846 (N_25846,N_22978,N_22043);
nor U25847 (N_25847,N_23562,N_22225);
nand U25848 (N_25848,N_23294,N_22067);
or U25849 (N_25849,N_22436,N_22380);
nor U25850 (N_25850,N_23610,N_22666);
nand U25851 (N_25851,N_23592,N_22243);
or U25852 (N_25852,N_22986,N_23872);
nor U25853 (N_25853,N_23793,N_23487);
xor U25854 (N_25854,N_22700,N_23739);
or U25855 (N_25855,N_22257,N_22332);
and U25856 (N_25856,N_23003,N_23567);
nor U25857 (N_25857,N_23328,N_23682);
xor U25858 (N_25858,N_22401,N_23525);
nor U25859 (N_25859,N_23308,N_23462);
or U25860 (N_25860,N_23983,N_23906);
xnor U25861 (N_25861,N_22775,N_22456);
and U25862 (N_25862,N_23751,N_23115);
or U25863 (N_25863,N_23176,N_22933);
nor U25864 (N_25864,N_22555,N_23599);
nor U25865 (N_25865,N_23233,N_23139);
and U25866 (N_25866,N_23414,N_22674);
nand U25867 (N_25867,N_23749,N_22514);
nand U25868 (N_25868,N_22659,N_23201);
or U25869 (N_25869,N_22887,N_23927);
nand U25870 (N_25870,N_23315,N_22400);
and U25871 (N_25871,N_23402,N_23009);
nor U25872 (N_25872,N_22117,N_23997);
or U25873 (N_25873,N_23041,N_23825);
or U25874 (N_25874,N_22760,N_23306);
nand U25875 (N_25875,N_23750,N_22979);
or U25876 (N_25876,N_23861,N_22749);
nand U25877 (N_25877,N_22054,N_22155);
or U25878 (N_25878,N_23058,N_22423);
nor U25879 (N_25879,N_23880,N_22957);
xor U25880 (N_25880,N_22344,N_23456);
and U25881 (N_25881,N_22262,N_23473);
and U25882 (N_25882,N_23663,N_22807);
xnor U25883 (N_25883,N_22827,N_23363);
xor U25884 (N_25884,N_22489,N_23800);
and U25885 (N_25885,N_22232,N_22981);
and U25886 (N_25886,N_22639,N_22188);
nand U25887 (N_25887,N_23528,N_22857);
or U25888 (N_25888,N_22243,N_23421);
or U25889 (N_25889,N_22985,N_22604);
or U25890 (N_25890,N_23854,N_22495);
or U25891 (N_25891,N_23955,N_22063);
xnor U25892 (N_25892,N_23701,N_23380);
nand U25893 (N_25893,N_23939,N_23609);
or U25894 (N_25894,N_23618,N_23891);
nor U25895 (N_25895,N_23720,N_22172);
or U25896 (N_25896,N_23696,N_22623);
nor U25897 (N_25897,N_23188,N_23284);
nor U25898 (N_25898,N_23191,N_22272);
xor U25899 (N_25899,N_22806,N_23648);
or U25900 (N_25900,N_22903,N_22669);
and U25901 (N_25901,N_23262,N_23507);
and U25902 (N_25902,N_22272,N_23858);
xnor U25903 (N_25903,N_22984,N_22287);
nor U25904 (N_25904,N_22984,N_23965);
nor U25905 (N_25905,N_23381,N_22481);
or U25906 (N_25906,N_22856,N_23539);
nand U25907 (N_25907,N_22367,N_22792);
or U25908 (N_25908,N_22879,N_23062);
nor U25909 (N_25909,N_23612,N_23940);
or U25910 (N_25910,N_22968,N_23520);
or U25911 (N_25911,N_22068,N_22302);
xor U25912 (N_25912,N_22710,N_22332);
or U25913 (N_25913,N_22182,N_23834);
xnor U25914 (N_25914,N_23240,N_22931);
nand U25915 (N_25915,N_22447,N_23325);
nor U25916 (N_25916,N_22791,N_22605);
nand U25917 (N_25917,N_23531,N_23965);
or U25918 (N_25918,N_22381,N_23967);
nor U25919 (N_25919,N_22790,N_22154);
nor U25920 (N_25920,N_22595,N_23742);
nand U25921 (N_25921,N_22855,N_23032);
and U25922 (N_25922,N_23487,N_23998);
xor U25923 (N_25923,N_22966,N_23549);
nor U25924 (N_25924,N_22852,N_22685);
nand U25925 (N_25925,N_23770,N_23052);
xor U25926 (N_25926,N_23672,N_22541);
or U25927 (N_25927,N_22332,N_23904);
nor U25928 (N_25928,N_22534,N_22627);
and U25929 (N_25929,N_23466,N_22007);
or U25930 (N_25930,N_23435,N_22364);
nor U25931 (N_25931,N_22420,N_22747);
xor U25932 (N_25932,N_22339,N_23435);
or U25933 (N_25933,N_22340,N_23298);
nand U25934 (N_25934,N_23093,N_23976);
or U25935 (N_25935,N_23280,N_22385);
and U25936 (N_25936,N_23600,N_23239);
nand U25937 (N_25937,N_23011,N_23125);
or U25938 (N_25938,N_22840,N_22928);
nand U25939 (N_25939,N_23788,N_22947);
or U25940 (N_25940,N_23821,N_23056);
and U25941 (N_25941,N_23350,N_22521);
xnor U25942 (N_25942,N_23011,N_23911);
xor U25943 (N_25943,N_22656,N_23653);
xor U25944 (N_25944,N_22114,N_23606);
and U25945 (N_25945,N_23413,N_22699);
and U25946 (N_25946,N_23551,N_23601);
and U25947 (N_25947,N_23184,N_23966);
nor U25948 (N_25948,N_23373,N_22225);
xor U25949 (N_25949,N_23784,N_23266);
xor U25950 (N_25950,N_23984,N_22003);
nand U25951 (N_25951,N_23676,N_23258);
or U25952 (N_25952,N_22844,N_22951);
nand U25953 (N_25953,N_22938,N_23093);
nor U25954 (N_25954,N_23083,N_22248);
nor U25955 (N_25955,N_22070,N_22350);
xor U25956 (N_25956,N_22294,N_22288);
nand U25957 (N_25957,N_22795,N_22505);
xnor U25958 (N_25958,N_22474,N_23910);
nor U25959 (N_25959,N_23637,N_22315);
nand U25960 (N_25960,N_23969,N_23651);
nor U25961 (N_25961,N_23150,N_22072);
and U25962 (N_25962,N_23722,N_23602);
and U25963 (N_25963,N_22360,N_23616);
and U25964 (N_25964,N_22696,N_23441);
and U25965 (N_25965,N_23427,N_22388);
and U25966 (N_25966,N_23960,N_23582);
xor U25967 (N_25967,N_22898,N_23697);
nand U25968 (N_25968,N_22254,N_22955);
nand U25969 (N_25969,N_22790,N_22544);
nand U25970 (N_25970,N_22334,N_23731);
or U25971 (N_25971,N_23161,N_23282);
and U25972 (N_25972,N_22091,N_22007);
xor U25973 (N_25973,N_23980,N_22947);
nor U25974 (N_25974,N_23702,N_23323);
and U25975 (N_25975,N_22775,N_22123);
or U25976 (N_25976,N_22290,N_23557);
and U25977 (N_25977,N_23593,N_22510);
or U25978 (N_25978,N_22186,N_22224);
or U25979 (N_25979,N_22300,N_23246);
nand U25980 (N_25980,N_23342,N_23144);
nand U25981 (N_25981,N_23628,N_22199);
and U25982 (N_25982,N_23230,N_23194);
and U25983 (N_25983,N_23602,N_23221);
xnor U25984 (N_25984,N_23968,N_22956);
xnor U25985 (N_25985,N_22861,N_22511);
nand U25986 (N_25986,N_22259,N_22329);
nand U25987 (N_25987,N_22234,N_23412);
xor U25988 (N_25988,N_22622,N_23901);
or U25989 (N_25989,N_22001,N_23792);
and U25990 (N_25990,N_23262,N_23409);
nand U25991 (N_25991,N_23861,N_22691);
nand U25992 (N_25992,N_23592,N_23793);
nor U25993 (N_25993,N_22245,N_23308);
nor U25994 (N_25994,N_22331,N_22603);
or U25995 (N_25995,N_22152,N_22162);
nand U25996 (N_25996,N_22956,N_22215);
nand U25997 (N_25997,N_23014,N_22294);
or U25998 (N_25998,N_22983,N_22874);
nand U25999 (N_25999,N_22957,N_23460);
nand U26000 (N_26000,N_24401,N_25561);
nand U26001 (N_26001,N_24066,N_25374);
nand U26002 (N_26002,N_25282,N_24068);
xor U26003 (N_26003,N_24433,N_24287);
nor U26004 (N_26004,N_24713,N_25660);
nand U26005 (N_26005,N_25341,N_25782);
and U26006 (N_26006,N_25557,N_25210);
nand U26007 (N_26007,N_25335,N_25217);
nand U26008 (N_26008,N_25475,N_24708);
or U26009 (N_26009,N_24440,N_25906);
nand U26010 (N_26010,N_24795,N_24638);
nor U26011 (N_26011,N_24019,N_24434);
nand U26012 (N_26012,N_24823,N_25492);
nor U26013 (N_26013,N_25932,N_25257);
xor U26014 (N_26014,N_24047,N_25084);
and U26015 (N_26015,N_25170,N_24918);
nand U26016 (N_26016,N_25138,N_24611);
and U26017 (N_26017,N_25320,N_24787);
nand U26018 (N_26018,N_25748,N_24710);
and U26019 (N_26019,N_24303,N_24830);
nor U26020 (N_26020,N_25076,N_25490);
and U26021 (N_26021,N_25201,N_25423);
nor U26022 (N_26022,N_25162,N_24013);
and U26023 (N_26023,N_24547,N_24032);
xnor U26024 (N_26024,N_25908,N_25303);
or U26025 (N_26025,N_24635,N_24408);
and U26026 (N_26026,N_24188,N_25603);
xor U26027 (N_26027,N_25161,N_25781);
xor U26028 (N_26028,N_25096,N_25893);
nand U26029 (N_26029,N_24317,N_25025);
or U26030 (N_26030,N_25836,N_24285);
xnor U26031 (N_26031,N_24956,N_25516);
or U26032 (N_26032,N_24201,N_25078);
nand U26033 (N_26033,N_25410,N_24206);
and U26034 (N_26034,N_24102,N_25895);
nand U26035 (N_26035,N_24500,N_24124);
nor U26036 (N_26036,N_25165,N_24414);
nand U26037 (N_26037,N_24779,N_24809);
or U26038 (N_26038,N_25017,N_24577);
or U26039 (N_26039,N_25184,N_25474);
and U26040 (N_26040,N_25048,N_25702);
nand U26041 (N_26041,N_24734,N_24924);
or U26042 (N_26042,N_25209,N_25828);
nand U26043 (N_26043,N_25744,N_25769);
and U26044 (N_26044,N_25866,N_25284);
or U26045 (N_26045,N_24798,N_25566);
nor U26046 (N_26046,N_25415,N_25774);
and U26047 (N_26047,N_24714,N_25588);
or U26048 (N_26048,N_24136,N_24170);
nor U26049 (N_26049,N_24179,N_24235);
nand U26050 (N_26050,N_25226,N_25234);
xnor U26051 (N_26051,N_24112,N_24274);
or U26052 (N_26052,N_24101,N_25350);
nor U26053 (N_26053,N_25759,N_24103);
or U26054 (N_26054,N_24839,N_25259);
xor U26055 (N_26055,N_25397,N_24561);
nand U26056 (N_26056,N_25141,N_25526);
or U26057 (N_26057,N_25652,N_24400);
nand U26058 (N_26058,N_24145,N_24447);
nor U26059 (N_26059,N_24522,N_25331);
nor U26060 (N_26060,N_24624,N_25695);
nor U26061 (N_26061,N_25177,N_25658);
nand U26062 (N_26062,N_24749,N_24295);
or U26063 (N_26063,N_25730,N_25590);
xor U26064 (N_26064,N_24007,N_24546);
and U26065 (N_26065,N_25204,N_24904);
and U26066 (N_26066,N_24791,N_25124);
xor U26067 (N_26067,N_24644,N_24603);
nor U26068 (N_26068,N_25054,N_24261);
or U26069 (N_26069,N_25442,N_25145);
and U26070 (N_26070,N_24557,N_25596);
nor U26071 (N_26071,N_24754,N_24914);
xor U26072 (N_26072,N_24014,N_25384);
xor U26073 (N_26073,N_25619,N_25785);
nor U26074 (N_26074,N_25742,N_25462);
nand U26075 (N_26075,N_25496,N_24692);
and U26076 (N_26076,N_25876,N_25562);
xor U26077 (N_26077,N_25667,N_25768);
xor U26078 (N_26078,N_24467,N_25931);
or U26079 (N_26079,N_24580,N_24377);
nor U26080 (N_26080,N_24175,N_24027);
and U26081 (N_26081,N_24571,N_25352);
nand U26082 (N_26082,N_24521,N_25511);
or U26083 (N_26083,N_24227,N_24954);
nor U26084 (N_26084,N_25907,N_25718);
and U26085 (N_26085,N_24504,N_25479);
and U26086 (N_26086,N_24927,N_24606);
and U26087 (N_26087,N_24207,N_24177);
and U26088 (N_26088,N_25656,N_25349);
or U26089 (N_26089,N_24864,N_25669);
xor U26090 (N_26090,N_24879,N_24456);
and U26091 (N_26091,N_25224,N_24951);
and U26092 (N_26092,N_24543,N_24497);
nand U26093 (N_26093,N_24674,N_25687);
nor U26094 (N_26094,N_24816,N_24540);
xnor U26095 (N_26095,N_25589,N_24190);
nor U26096 (N_26096,N_25127,N_24132);
or U26097 (N_26097,N_25790,N_25533);
xnor U26098 (N_26098,N_25583,N_25011);
nor U26099 (N_26099,N_25073,N_25424);
xnor U26100 (N_26100,N_24121,N_24881);
or U26101 (N_26101,N_25091,N_24378);
xnor U26102 (N_26102,N_25498,N_25045);
xor U26103 (N_26103,N_24616,N_25435);
or U26104 (N_26104,N_25007,N_25304);
xnor U26105 (N_26105,N_25079,N_25875);
nor U26106 (N_26106,N_25524,N_24872);
and U26107 (N_26107,N_24618,N_24394);
nor U26108 (N_26108,N_25394,N_24720);
nor U26109 (N_26109,N_25501,N_25560);
and U26110 (N_26110,N_24001,N_25369);
xor U26111 (N_26111,N_25216,N_24490);
xor U26112 (N_26112,N_24367,N_24528);
and U26113 (N_26113,N_24129,N_25860);
nor U26114 (N_26114,N_25633,N_24473);
or U26115 (N_26115,N_25738,N_25543);
nor U26116 (N_26116,N_25044,N_25679);
nor U26117 (N_26117,N_25746,N_24096);
or U26118 (N_26118,N_25636,N_24948);
or U26119 (N_26119,N_25154,N_25684);
or U26120 (N_26120,N_24648,N_24189);
or U26121 (N_26121,N_25148,N_24759);
nor U26122 (N_26122,N_24925,N_25878);
nor U26123 (N_26123,N_25466,N_25572);
or U26124 (N_26124,N_25714,N_24488);
nor U26125 (N_26125,N_25586,N_25457);
and U26126 (N_26126,N_25649,N_24843);
xor U26127 (N_26127,N_25556,N_25723);
or U26128 (N_26128,N_24459,N_24994);
and U26129 (N_26129,N_25997,N_24991);
xor U26130 (N_26130,N_25346,N_24251);
xor U26131 (N_26131,N_25013,N_24181);
nand U26132 (N_26132,N_24614,N_25788);
nand U26133 (N_26133,N_24288,N_25842);
nor U26134 (N_26134,N_25082,N_24147);
and U26135 (N_26135,N_25637,N_24184);
or U26136 (N_26136,N_25061,N_24592);
or U26137 (N_26137,N_24671,N_24479);
or U26138 (N_26138,N_25092,N_24760);
nand U26139 (N_26139,N_25593,N_24219);
nand U26140 (N_26140,N_25326,N_24679);
xnor U26141 (N_26141,N_24584,N_25072);
nor U26142 (N_26142,N_24273,N_24984);
or U26143 (N_26143,N_25886,N_24628);
and U26144 (N_26144,N_25131,N_24142);
and U26145 (N_26145,N_24133,N_25814);
nand U26146 (N_26146,N_24666,N_24097);
nand U26147 (N_26147,N_24800,N_25775);
xor U26148 (N_26148,N_24595,N_24135);
and U26149 (N_26149,N_25916,N_24896);
and U26150 (N_26150,N_24043,N_24932);
xnor U26151 (N_26151,N_25239,N_25232);
or U26152 (N_26152,N_25806,N_25821);
nand U26153 (N_26153,N_25142,N_24079);
and U26154 (N_26154,N_25610,N_24726);
xnor U26155 (N_26155,N_25591,N_24141);
nor U26156 (N_26156,N_24339,N_24410);
and U26157 (N_26157,N_24641,N_25368);
and U26158 (N_26158,N_24765,N_25532);
or U26159 (N_26159,N_24822,N_25443);
nor U26160 (N_26160,N_25975,N_24238);
xnor U26161 (N_26161,N_24084,N_25164);
xnor U26162 (N_26162,N_25925,N_25202);
and U26163 (N_26163,N_25697,N_24536);
and U26164 (N_26164,N_25459,N_24398);
or U26165 (N_26165,N_24116,N_25758);
nand U26166 (N_26166,N_24368,N_24021);
and U26167 (N_26167,N_25578,N_25522);
and U26168 (N_26168,N_25707,N_24252);
or U26169 (N_26169,N_25481,N_25926);
or U26170 (N_26170,N_24267,N_25405);
nor U26171 (N_26171,N_24688,N_24418);
nor U26172 (N_26172,N_24890,N_25322);
xnor U26173 (N_26173,N_24423,N_24115);
xor U26174 (N_26174,N_25275,N_25733);
nor U26175 (N_26175,N_25467,N_24900);
nand U26176 (N_26176,N_25712,N_24723);
xor U26177 (N_26177,N_24045,N_24108);
nand U26178 (N_26178,N_25792,N_24137);
and U26179 (N_26179,N_24200,N_25432);
nand U26180 (N_26180,N_24750,N_25570);
nor U26181 (N_26181,N_25644,N_25632);
nor U26182 (N_26182,N_24392,N_24849);
and U26183 (N_26183,N_24877,N_24863);
and U26184 (N_26184,N_25230,N_25049);
and U26185 (N_26185,N_25100,N_24088);
xnor U26186 (N_26186,N_24581,N_24769);
nand U26187 (N_26187,N_24220,N_24861);
nor U26188 (N_26188,N_24685,N_25575);
nor U26189 (N_26189,N_25278,N_24080);
and U26190 (N_26190,N_25323,N_25949);
and U26191 (N_26191,N_25834,N_24582);
xnor U26192 (N_26192,N_24901,N_25212);
and U26193 (N_26193,N_24499,N_25118);
nor U26194 (N_26194,N_24348,N_24552);
or U26195 (N_26195,N_25678,N_25213);
xor U26196 (N_26196,N_25540,N_25653);
xnor U26197 (N_26197,N_24344,N_24366);
nand U26198 (N_26198,N_24551,N_24331);
nand U26199 (N_26199,N_24903,N_25175);
and U26200 (N_26200,N_24451,N_24967);
or U26201 (N_26201,N_25240,N_25430);
xnor U26202 (N_26202,N_24813,N_24269);
or U26203 (N_26203,N_24040,N_25081);
xor U26204 (N_26204,N_24248,N_24429);
or U26205 (N_26205,N_24144,N_24257);
nand U26206 (N_26206,N_25174,N_25298);
xor U26207 (N_26207,N_25190,N_25329);
xnor U26208 (N_26208,N_25178,N_24283);
or U26209 (N_26209,N_25456,N_25861);
nand U26210 (N_26210,N_25086,N_25675);
nor U26211 (N_26211,N_25668,N_24781);
or U26212 (N_26212,N_24656,N_25276);
or U26213 (N_26213,N_24544,N_24508);
xnor U26214 (N_26214,N_24690,N_25804);
and U26215 (N_26215,N_24887,N_24634);
and U26216 (N_26216,N_24977,N_24302);
and U26217 (N_26217,N_25225,N_25356);
or U26218 (N_26218,N_25183,N_24773);
xor U26219 (N_26219,N_24512,N_24352);
and U26220 (N_26220,N_24715,N_24069);
nor U26221 (N_26221,N_24597,N_25000);
nor U26222 (N_26222,N_24017,N_25534);
xnor U26223 (N_26223,N_24598,N_25710);
nand U26224 (N_26224,N_24381,N_24646);
xor U26225 (N_26225,N_25939,N_24286);
and U26226 (N_26226,N_24055,N_25465);
or U26227 (N_26227,N_24041,N_24844);
nor U26228 (N_26228,N_24262,N_24778);
nor U26229 (N_26229,N_24402,N_24695);
and U26230 (N_26230,N_25328,N_25783);
or U26231 (N_26231,N_25324,N_25905);
xnor U26232 (N_26232,N_24963,N_25681);
xor U26233 (N_26233,N_25943,N_24507);
nand U26234 (N_26234,N_25724,N_25327);
nor U26235 (N_26235,N_25961,N_24475);
and U26236 (N_26236,N_24593,N_25973);
nand U26237 (N_26237,N_25077,N_25252);
or U26238 (N_26238,N_24847,N_25268);
xnor U26239 (N_26239,N_24746,N_24961);
xor U26240 (N_26240,N_24403,N_25646);
or U26241 (N_26241,N_25223,N_25063);
xnor U26242 (N_26242,N_25885,N_24793);
nor U26243 (N_26243,N_25580,N_25109);
or U26244 (N_26244,N_24159,N_25321);
and U26245 (N_26245,N_25125,N_24139);
xor U26246 (N_26246,N_25046,N_25597);
and U26247 (N_26247,N_25699,N_24572);
nor U26248 (N_26248,N_24596,N_25186);
nand U26249 (N_26249,N_24659,N_24933);
or U26250 (N_26250,N_24675,N_24321);
xor U26251 (N_26251,N_25657,N_25477);
nand U26252 (N_26252,N_24217,N_25904);
xnor U26253 (N_26253,N_24386,N_25877);
xor U26254 (N_26254,N_24011,N_25140);
nand U26255 (N_26255,N_24929,N_24371);
nand U26256 (N_26256,N_24837,N_25717);
and U26257 (N_26257,N_24815,N_24763);
xnor U26258 (N_26258,N_24930,N_25791);
nand U26259 (N_26259,N_24199,N_24478);
xnor U26260 (N_26260,N_25446,N_24563);
and U26261 (N_26261,N_24875,N_25917);
xor U26262 (N_26262,N_24629,N_24247);
or U26263 (N_26263,N_24686,N_25808);
nand U26264 (N_26264,N_25110,N_24098);
xor U26265 (N_26265,N_25843,N_24335);
xor U26266 (N_26266,N_25277,N_24973);
xor U26267 (N_26267,N_24884,N_25848);
nor U26268 (N_26268,N_25311,N_24446);
nor U26269 (N_26269,N_24501,N_24486);
xor U26270 (N_26270,N_24256,N_24626);
and U26271 (N_26271,N_25691,N_24704);
xnor U26272 (N_26272,N_25281,N_24642);
xnor U26273 (N_26273,N_25012,N_24535);
nor U26274 (N_26274,N_24233,N_25255);
and U26275 (N_26275,N_24652,N_25030);
nand U26276 (N_26276,N_24856,N_24702);
xor U26277 (N_26277,N_24464,N_24030);
xnor U26278 (N_26278,N_24851,N_25295);
xor U26279 (N_26279,N_24766,N_24889);
xnor U26280 (N_26280,N_24026,N_25355);
xnor U26281 (N_26281,N_24637,N_25634);
and U26282 (N_26282,N_24384,N_25795);
or U26283 (N_26283,N_24353,N_24171);
and U26284 (N_26284,N_25599,N_25399);
nand U26285 (N_26285,N_24023,N_25999);
nand U26286 (N_26286,N_25813,N_25852);
xnor U26287 (N_26287,N_25302,N_24998);
nor U26288 (N_26288,N_24029,N_24073);
xnor U26289 (N_26289,N_25293,N_24910);
nor U26290 (N_26290,N_25801,N_25574);
nor U26291 (N_26291,N_24074,N_24018);
nor U26292 (N_26292,N_24050,N_24359);
xor U26293 (N_26293,N_25250,N_25229);
nor U26294 (N_26294,N_24509,N_24496);
nor U26295 (N_26295,N_24452,N_24495);
nor U26296 (N_26296,N_25071,N_24037);
or U26297 (N_26297,N_25732,N_24345);
nor U26298 (N_26298,N_25408,N_24525);
xnor U26299 (N_26299,N_24513,N_24134);
nor U26300 (N_26300,N_24942,N_24039);
and U26301 (N_26301,N_24873,N_25631);
or U26302 (N_26302,N_25470,N_24182);
and U26303 (N_26303,N_24485,N_24803);
or U26304 (N_26304,N_24911,N_25308);
and U26305 (N_26305,N_24539,N_25114);
xnor U26306 (N_26306,N_24064,N_25845);
nand U26307 (N_26307,N_25058,N_24833);
nor U26308 (N_26308,N_25090,N_25617);
or U26309 (N_26309,N_25854,N_24567);
or U26310 (N_26310,N_24310,N_25418);
nand U26311 (N_26311,N_25431,N_24448);
nand U26312 (N_26312,N_25559,N_25332);
nor U26313 (N_26313,N_25715,N_25409);
xor U26314 (N_26314,N_25864,N_24542);
nand U26315 (N_26315,N_25515,N_24154);
and U26316 (N_26316,N_25488,N_25246);
or U26317 (N_26317,N_24906,N_24117);
xor U26318 (N_26318,N_25620,N_25978);
nand U26319 (N_26319,N_25741,N_24640);
nor U26320 (N_26320,N_25129,N_25153);
nand U26321 (N_26321,N_24105,N_24304);
nor U26322 (N_26322,N_24458,N_24263);
and U26323 (N_26323,N_24387,N_24296);
and U26324 (N_26324,N_25334,N_25549);
and U26325 (N_26325,N_24426,N_25789);
or U26326 (N_26326,N_25510,N_25152);
nor U26327 (N_26327,N_24436,N_24774);
nand U26328 (N_26328,N_25215,N_24526);
and U26329 (N_26329,N_25936,N_24711);
or U26330 (N_26330,N_24314,N_25608);
and U26331 (N_26331,N_25087,N_25292);
nand U26332 (N_26332,N_24435,N_25553);
and U26333 (N_26333,N_25052,N_25353);
nand U26334 (N_26334,N_25976,N_25191);
nor U26335 (N_26335,N_24211,N_24768);
or U26336 (N_26336,N_24975,N_25780);
nor U26337 (N_26337,N_25060,N_24104);
xnor U26338 (N_26338,N_24559,N_25606);
xor U26339 (N_26339,N_24968,N_25338);
nand U26340 (N_26340,N_24550,N_24494);
xor U26341 (N_26341,N_24989,N_25538);
and U26342 (N_26342,N_25909,N_24369);
and U26343 (N_26343,N_24920,N_24338);
or U26344 (N_26344,N_25482,N_25527);
nor U26345 (N_26345,N_24143,N_24076);
nor U26346 (N_26346,N_25256,N_24917);
nor U26347 (N_26347,N_25506,N_25753);
nand U26348 (N_26348,N_25495,N_24246);
and U26349 (N_26349,N_24315,N_24748);
nor U26350 (N_26350,N_25417,N_25624);
nand U26351 (N_26351,N_25362,N_24309);
or U26352 (N_26352,N_24453,N_25371);
xnor U26353 (N_26353,N_25870,N_25600);
nand U26354 (N_26354,N_25584,N_25342);
nor U26355 (N_26355,N_24853,N_24300);
or U26356 (N_26356,N_25940,N_24301);
and U26357 (N_26357,N_24320,N_25771);
nand U26358 (N_26358,N_25440,N_24416);
or U26359 (N_26359,N_24916,N_25245);
or U26360 (N_26360,N_24430,N_24379);
and U26361 (N_26361,N_24958,N_25249);
nand U26362 (N_26362,N_25508,N_25144);
and U26363 (N_26363,N_24208,N_24940);
nand U26364 (N_26364,N_25247,N_24757);
nor U26365 (N_26365,N_24744,N_24293);
nor U26366 (N_26366,N_25763,N_25003);
nand U26367 (N_26367,N_25317,N_25413);
and U26368 (N_26368,N_25280,N_25289);
xor U26369 (N_26369,N_24683,N_24806);
or U26370 (N_26370,N_24196,N_24163);
and U26371 (N_26371,N_25163,N_25370);
nor U26372 (N_26372,N_25751,N_24937);
xnor U26373 (N_26373,N_24099,N_24297);
nor U26374 (N_26374,N_25396,N_25489);
or U26375 (N_26375,N_25571,N_24185);
xor U26376 (N_26376,N_25376,N_25523);
xnor U26377 (N_26377,N_25402,N_25502);
nand U26378 (N_26378,N_24305,N_24375);
nor U26379 (N_26379,N_24993,N_25244);
or U26380 (N_26380,N_25625,N_24623);
nand U26381 (N_26381,N_25964,N_25372);
nor U26382 (N_26382,N_25988,N_25703);
xnor U26383 (N_26383,N_25115,N_25406);
nor U26384 (N_26384,N_24341,N_24031);
and U26385 (N_26385,N_25261,N_24072);
nor U26386 (N_26386,N_25550,N_25798);
nor U26387 (N_26387,N_25812,N_25910);
nand U26388 (N_26388,N_25196,N_24980);
or U26389 (N_26389,N_25108,N_24239);
nand U26390 (N_26390,N_24653,N_25770);
nor U26391 (N_26391,N_25500,N_24838);
nor U26392 (N_26392,N_25472,N_25199);
or U26393 (N_26393,N_24004,N_24390);
nand U26394 (N_26394,N_24046,N_24056);
xnor U26395 (N_26395,N_24891,N_25220);
xor U26396 (N_26396,N_24531,N_25690);
nand U26397 (N_26397,N_25994,N_25043);
xnor U26398 (N_26398,N_24093,N_24484);
or U26399 (N_26399,N_24845,N_25139);
xnor U26400 (N_26400,N_25933,N_24931);
or U26401 (N_26401,N_25857,N_24785);
nor U26402 (N_26402,N_24034,N_24732);
xnor U26403 (N_26403,N_24575,N_24255);
nand U26404 (N_26404,N_25375,N_24568);
or U26405 (N_26405,N_24449,N_25883);
and U26406 (N_26406,N_24573,N_25521);
nor U26407 (N_26407,N_24681,N_24882);
or U26408 (N_26408,N_24608,N_24985);
or U26409 (N_26409,N_24747,N_24794);
and U26410 (N_26410,N_25080,N_25547);
or U26411 (N_26411,N_24583,N_25514);
nand U26412 (N_26412,N_25033,N_25944);
nand U26413 (N_26413,N_25412,N_25053);
or U26414 (N_26414,N_24682,N_24230);
nand U26415 (N_26415,N_25891,N_25429);
or U26416 (N_26416,N_25272,N_25680);
nand U26417 (N_26417,N_24601,N_25018);
nor U26418 (N_26418,N_25373,N_24558);
or U26419 (N_26419,N_24878,N_24389);
nand U26420 (N_26420,N_25552,N_25478);
xnor U26421 (N_26421,N_25065,N_25984);
or U26422 (N_26422,N_24498,N_24709);
nand U26423 (N_26423,N_25345,N_25366);
or U26424 (N_26424,N_24362,N_24393);
xnor U26425 (N_26425,N_25039,N_25378);
nor U26426 (N_26426,N_25157,N_24059);
and U26427 (N_26427,N_25051,N_24721);
nor U26428 (N_26428,N_25849,N_25387);
xor U26429 (N_26429,N_25688,N_24533);
nand U26430 (N_26430,N_25734,N_24992);
or U26431 (N_26431,N_25414,N_24388);
nand U26432 (N_26432,N_25601,N_24307);
and U26433 (N_26433,N_25727,N_25787);
xnor U26434 (N_26434,N_24204,N_24218);
or U26435 (N_26435,N_25149,N_24203);
and U26436 (N_26436,N_24454,N_24049);
nor U26437 (N_26437,N_25156,N_25582);
or U26438 (N_26438,N_24921,N_25517);
and U26439 (N_26439,N_25720,N_25513);
xnor U26440 (N_26440,N_24862,N_25403);
nand U26441 (N_26441,N_24926,N_25829);
and U26442 (N_26442,N_25546,N_25889);
or U26443 (N_26443,N_24158,N_25294);
or U26444 (N_26444,N_24999,N_25855);
or U26445 (N_26445,N_24894,N_24858);
xor U26446 (N_26446,N_24953,N_24176);
nor U26447 (N_26447,N_24249,N_25760);
xnor U26448 (N_26448,N_24413,N_24169);
or U26449 (N_26449,N_25833,N_25121);
xnor U26450 (N_26450,N_25683,N_25029);
and U26451 (N_26451,N_24758,N_24422);
and U26452 (N_26452,N_25006,N_24518);
or U26453 (N_26453,N_24783,N_24915);
xor U26454 (N_26454,N_24326,N_25535);
nand U26455 (N_26455,N_24519,N_24048);
xnor U26456 (N_26456,N_24660,N_24586);
nand U26457 (N_26457,N_25262,N_25626);
or U26458 (N_26458,N_24716,N_24537);
or U26459 (N_26459,N_25206,N_25594);
nand U26460 (N_26460,N_24865,N_24632);
and U26461 (N_26461,N_24399,N_24938);
or U26462 (N_26462,N_24155,N_25130);
and U26463 (N_26463,N_24358,N_24483);
nand U26464 (N_26464,N_24775,N_25444);
or U26465 (N_26465,N_24654,N_25010);
or U26466 (N_26466,N_25119,N_24852);
or U26467 (N_26467,N_25662,N_25200);
and U26468 (N_26468,N_24127,N_25872);
xnor U26469 (N_26469,N_25974,N_24052);
and U26470 (N_26470,N_24243,N_25612);
or U26471 (N_26471,N_24502,N_24780);
or U26472 (N_26472,N_25426,N_24782);
and U26473 (N_26473,N_25749,N_24346);
nor U26474 (N_26474,N_24223,N_24193);
xnor U26475 (N_26475,N_25111,N_24126);
nor U26476 (N_26476,N_25158,N_25197);
and U26477 (N_26477,N_25064,N_24123);
nor U26478 (N_26478,N_25981,N_24372);
nor U26479 (N_26479,N_25663,N_25260);
nor U26480 (N_26480,N_24612,N_25062);
nand U26481 (N_26481,N_25627,N_24324);
nand U26482 (N_26482,N_24665,N_24425);
nor U26483 (N_26483,N_24860,N_25831);
and U26484 (N_26484,N_25659,N_24161);
xor U26485 (N_26485,N_25301,N_24342);
nor U26486 (N_26486,N_24857,N_24538);
nor U26487 (N_26487,N_24187,N_24174);
nand U26488 (N_26488,N_24265,N_24357);
or U26489 (N_26489,N_25070,N_24028);
and U26490 (N_26490,N_25797,N_24736);
nand U26491 (N_26491,N_25309,N_25358);
or U26492 (N_26492,N_24836,N_24620);
xnor U26493 (N_26493,N_25023,N_24441);
nand U26494 (N_26494,N_24699,N_25469);
nand U26495 (N_26495,N_25454,N_24471);
or U26496 (N_26496,N_24354,N_25537);
and U26497 (N_26497,N_25095,N_25882);
nand U26498 (N_26498,N_25725,N_24489);
nand U26499 (N_26499,N_25728,N_25464);
or U26500 (N_26500,N_25764,N_25731);
or U26501 (N_26501,N_24730,N_24275);
xor U26502 (N_26502,N_25541,N_24202);
nand U26503 (N_26503,N_25271,N_24696);
xnor U26504 (N_26504,N_24808,N_25339);
nor U26505 (N_26505,N_24825,N_24867);
xor U26506 (N_26506,N_25015,N_25987);
and U26507 (N_26507,N_24470,N_25736);
or U26508 (N_26508,N_25841,N_24703);
and U26509 (N_26509,N_24812,N_25439);
nor U26510 (N_26510,N_24850,N_25238);
nor U26511 (N_26511,N_24491,N_24271);
nand U26512 (N_26512,N_24576,N_24974);
nor U26513 (N_26513,N_25844,N_24311);
nor U26514 (N_26514,N_24125,N_25173);
nor U26515 (N_26515,N_25923,N_24647);
nor U26516 (N_26516,N_24655,N_25057);
nand U26517 (N_26517,N_25390,N_25027);
nand U26518 (N_26518,N_24385,N_25313);
nor U26519 (N_26519,N_24070,N_24087);
nand U26520 (N_26520,N_25433,N_24109);
xor U26521 (N_26521,N_24336,N_25168);
nand U26522 (N_26522,N_24523,N_25512);
nor U26523 (N_26523,N_24415,N_25473);
nand U26524 (N_26524,N_24530,N_25607);
or U26525 (N_26525,N_24742,N_25069);
or U26526 (N_26526,N_25008,N_24090);
or U26527 (N_26527,N_25180,N_25705);
xnor U26528 (N_26528,N_24332,N_24667);
nor U26529 (N_26529,N_24365,N_25270);
xor U26530 (N_26530,N_25333,N_24691);
nand U26531 (N_26531,N_24636,N_24564);
xor U26532 (N_26532,N_25151,N_25265);
or U26533 (N_26533,N_24067,N_24591);
nand U26534 (N_26534,N_24111,N_24745);
xor U26535 (N_26535,N_24417,N_24361);
and U26536 (N_26536,N_25504,N_24284);
nor U26537 (N_26537,N_24673,N_25445);
and U26538 (N_26538,N_25604,N_25810);
nor U26539 (N_26539,N_25041,N_25776);
nor U26540 (N_26540,N_24549,N_24396);
nand U26541 (N_26541,N_24796,N_25026);
and U26542 (N_26542,N_25542,N_25894);
nand U26543 (N_26543,N_24329,N_25581);
nor U26544 (N_26544,N_24565,N_24630);
xnor U26545 (N_26545,N_25629,N_24038);
or U26546 (N_26546,N_25136,N_24898);
nor U26547 (N_26547,N_24566,N_24035);
or U26548 (N_26548,N_25316,N_24517);
and U26549 (N_26549,N_24290,N_24210);
xor U26550 (N_26550,N_25169,N_25851);
nand U26551 (N_26551,N_25134,N_24892);
and U26552 (N_26552,N_24015,N_24245);
nor U26553 (N_26553,N_24560,N_25743);
xnor U26554 (N_26554,N_24725,N_24002);
nand U26555 (N_26555,N_24083,N_25283);
nand U26556 (N_26556,N_25420,N_24016);
and U26557 (N_26557,N_24114,N_25921);
nand U26558 (N_26558,N_25530,N_25871);
nand U26559 (N_26559,N_24738,N_24053);
nor U26560 (N_26560,N_25159,N_25066);
xor U26561 (N_26561,N_24743,N_24131);
nor U26562 (N_26562,N_25651,N_24254);
nor U26563 (N_26563,N_24859,N_25471);
and U26564 (N_26564,N_24506,N_25098);
and U26565 (N_26565,N_25385,N_25336);
nor U26566 (N_26566,N_24854,N_24776);
or U26567 (N_26567,N_24717,N_25449);
xnor U26568 (N_26568,N_25647,N_24482);
nor U26569 (N_26569,N_25938,N_25116);
and U26570 (N_26570,N_25900,N_25747);
nor U26571 (N_26571,N_24602,N_25038);
nor U26572 (N_26572,N_25393,N_24649);
and U26573 (N_26573,N_24266,N_25105);
and U26574 (N_26574,N_24444,N_25056);
xor U26575 (N_26575,N_24874,N_24194);
or U26576 (N_26576,N_24827,N_24347);
nand U26577 (N_26577,N_24350,N_25991);
and U26578 (N_26578,N_24095,N_25945);
nand U26579 (N_26579,N_25615,N_25438);
nor U26580 (N_26580,N_25614,N_24986);
or U26581 (N_26581,N_24680,N_25266);
and U26582 (N_26582,N_24012,N_25243);
and U26583 (N_26583,N_24183,N_24777);
xnor U26584 (N_26584,N_24042,N_25097);
and U26585 (N_26585,N_25171,N_24191);
nand U26586 (N_26586,N_24545,N_24876);
nor U26587 (N_26587,N_24364,N_24427);
nand U26588 (N_26588,N_25416,N_25686);
and U26589 (N_26589,N_25761,N_24870);
nor U26590 (N_26590,N_24236,N_24804);
nand U26591 (N_26591,N_25953,N_25868);
nand U26592 (N_26592,N_25505,N_25595);
xor U26593 (N_26593,N_25959,N_25364);
xor U26594 (N_26594,N_25958,N_25419);
xor U26595 (N_26595,N_24645,N_24676);
nand U26596 (N_26596,N_25133,N_24455);
and U26597 (N_26597,N_25484,N_24472);
or U26598 (N_26598,N_24609,N_25859);
xor U26599 (N_26599,N_25509,N_25242);
nor U26600 (N_26600,N_24946,N_25989);
nor U26601 (N_26601,N_25640,N_25956);
nor U26602 (N_26602,N_25853,N_25696);
xnor U26603 (N_26603,N_25347,N_24173);
xnor U26604 (N_26604,N_24520,N_25458);
nor U26605 (N_26605,N_25865,N_25083);
or U26606 (N_26606,N_24790,N_25701);
xor U26607 (N_26607,N_25737,N_25367);
or U26608 (N_26608,N_24312,N_24751);
and U26609 (N_26609,N_24578,N_24619);
nor U26610 (N_26610,N_24316,N_25913);
nor U26611 (N_26611,N_24672,N_25726);
xnor U26612 (N_26612,N_24770,N_24888);
nor U26613 (N_26613,N_25862,N_24212);
and U26614 (N_26614,N_25912,N_25155);
and U26615 (N_26615,N_24149,N_25343);
or U26616 (N_26616,N_24832,N_24527);
nor U26617 (N_26617,N_24420,N_25740);
nor U26618 (N_26618,N_25765,N_24712);
xor U26619 (N_26619,N_25930,N_24835);
or U26620 (N_26620,N_25757,N_25185);
nand U26621 (N_26621,N_24281,N_25729);
or U26622 (N_26622,N_24051,N_24323);
xor U26623 (N_26623,N_24514,N_24363);
and U26624 (N_26624,N_25483,N_24268);
nand U26625 (N_26625,N_25363,N_25055);
or U26626 (N_26626,N_25040,N_25305);
xor U26627 (N_26627,N_25914,N_24009);
nor U26628 (N_26628,N_25207,N_25398);
nand U26629 (N_26629,N_25274,N_25545);
xor U26630 (N_26630,N_25085,N_24737);
xor U26631 (N_26631,N_24950,N_25968);
or U26632 (N_26632,N_24466,N_24981);
xor U26633 (N_26633,N_24270,N_25693);
xor U26634 (N_26634,N_25621,N_25670);
or U26635 (N_26635,N_24198,N_24298);
and U26636 (N_26636,N_25592,N_25383);
and U26637 (N_26637,N_24541,N_25227);
nand U26638 (N_26638,N_24282,N_25869);
nor U26639 (N_26639,N_24982,N_25901);
nand U26640 (N_26640,N_25195,N_24585);
xnor U26641 (N_26641,N_24741,N_24625);
and U26642 (N_26642,N_25643,N_25189);
xor U26643 (N_26643,N_24988,N_24569);
xnor U26644 (N_26644,N_24380,N_25379);
nor U26645 (N_26645,N_25979,N_24579);
nor U26646 (N_26646,N_25377,N_25248);
xor U26647 (N_26647,N_25618,N_24062);
or U26648 (N_26648,N_25579,N_24325);
xnor U26649 (N_26649,N_24658,N_25555);
and U26650 (N_26650,N_25692,N_24438);
xnor U26651 (N_26651,N_24272,N_25896);
or U26652 (N_26652,N_24771,N_25094);
or U26653 (N_26653,N_25969,N_25766);
xor U26654 (N_26654,N_24330,N_24792);
or U26655 (N_26655,N_25609,N_25059);
nor U26656 (N_26656,N_24292,N_24669);
nand U26657 (N_26657,N_25762,N_24221);
and U26658 (N_26658,N_25957,N_24532);
and U26659 (N_26659,N_24570,N_25287);
nand U26660 (N_26660,N_25031,N_25665);
or U26661 (N_26661,N_25650,N_24829);
nand U26662 (N_26662,N_25179,N_24590);
nor U26663 (N_26663,N_25359,N_24842);
nor U26664 (N_26664,N_25441,N_24562);
nand U26665 (N_26665,N_25539,N_24086);
or U26666 (N_26666,N_24356,N_25993);
xor U26667 (N_26667,N_25708,N_24106);
nand U26668 (N_26668,N_25682,N_25434);
xor U26669 (N_26669,N_25203,N_24197);
or U26670 (N_26670,N_24600,N_24727);
xor U26671 (N_26671,N_25779,N_24828);
nand U26672 (N_26672,N_25754,N_24664);
or U26673 (N_26673,N_25019,N_25273);
nand U26674 (N_26674,N_24821,N_25573);
nor U26675 (N_26675,N_25638,N_24006);
nor U26676 (N_26676,N_25948,N_24912);
nor U26677 (N_26677,N_25952,N_24319);
nand U26678 (N_26678,N_25767,N_24556);
nand U26679 (N_26679,N_24772,N_25167);
xnor U26680 (N_26680,N_25587,N_24972);
and U26681 (N_26681,N_24817,N_24529);
nand U26682 (N_26682,N_24633,N_25700);
xor U26683 (N_26683,N_25722,N_25671);
nor U26684 (N_26684,N_25137,N_24555);
xor U26685 (N_26685,N_24024,N_24995);
or U26686 (N_26686,N_25922,N_25721);
xor U26687 (N_26687,N_24701,N_24622);
and U26688 (N_26688,N_24391,N_25817);
nor U26689 (N_26689,N_24820,N_25068);
xor U26690 (N_26690,N_24008,N_25093);
or U26691 (N_26691,N_24697,N_24923);
xor U26692 (N_26692,N_24405,N_24264);
nand U26693 (N_26693,N_25300,N_25823);
and U26694 (N_26694,N_24662,N_24237);
or U26695 (N_26695,N_24395,N_25147);
xor U26696 (N_26696,N_24805,N_25123);
nor U26697 (N_26697,N_25194,N_25067);
or U26698 (N_26698,N_25918,N_24883);
nand U26699 (N_26699,N_25887,N_25146);
or U26700 (N_26700,N_24684,N_24719);
or U26701 (N_26701,N_24594,N_25622);
or U26702 (N_26702,N_24605,N_25296);
xor U26703 (N_26703,N_24242,N_25551);
xor U26704 (N_26704,N_25966,N_24503);
nand U26705 (N_26705,N_25800,N_25421);
xnor U26706 (N_26706,N_25847,N_24848);
and U26707 (N_26707,N_24060,N_24477);
or U26708 (N_26708,N_25404,N_24885);
or U26709 (N_26709,N_25306,N_25919);
nand U26710 (N_26710,N_25827,N_24661);
xor U26711 (N_26711,N_24318,N_24229);
or U26712 (N_26712,N_25354,N_24941);
nand U26713 (N_26713,N_25036,N_25635);
or U26714 (N_26714,N_24928,N_25529);
xnor U26715 (N_26715,N_24554,N_25839);
or U26716 (N_26716,N_24990,N_25407);
nand U26717 (N_26717,N_25351,N_25577);
nor U26718 (N_26718,N_24949,N_24959);
nor U26719 (N_26719,N_24278,N_25218);
xor U26720 (N_26720,N_25951,N_25856);
nor U26721 (N_26721,N_24919,N_24445);
nor U26722 (N_26722,N_24934,N_25480);
or U26723 (N_26723,N_25493,N_25735);
nand U26724 (N_26724,N_24152,N_24299);
xor U26725 (N_26725,N_24044,N_24607);
xnor U26726 (N_26726,N_24718,N_25929);
nand U26727 (N_26727,N_24764,N_25982);
nand U26728 (N_26728,N_24151,N_25568);
and U26729 (N_26729,N_25102,N_25824);
nand U26730 (N_26730,N_24058,N_24480);
and U26731 (N_26731,N_24908,N_24178);
or U26732 (N_26732,N_24668,N_25035);
or U26733 (N_26733,N_24966,N_25279);
nand U26734 (N_26734,N_25422,N_24786);
nor U26735 (N_26735,N_24244,N_24976);
nor U26736 (N_26736,N_24148,N_24869);
and U26737 (N_26737,N_24627,N_24957);
nor U26738 (N_26738,N_25400,N_25074);
xnor U26739 (N_26739,N_25507,N_24213);
xor U26740 (N_26740,N_24650,N_25803);
xnor U26741 (N_26741,N_24071,N_25009);
nor U26742 (N_26742,N_24003,N_25251);
or U26743 (N_26743,N_25585,N_25267);
or U26744 (N_26744,N_24831,N_24360);
and U26745 (N_26745,N_24437,N_25528);
xnor U26746 (N_26746,N_24788,N_24907);
nand U26747 (N_26747,N_25811,N_24524);
and U26748 (N_26748,N_24707,N_24553);
and U26749 (N_26749,N_24291,N_25641);
nor U26750 (N_26750,N_24728,N_24166);
nand U26751 (N_26751,N_25388,N_25330);
xor U26752 (N_26752,N_25694,N_25297);
xor U26753 (N_26753,N_24376,N_24327);
xnor U26754 (N_26754,N_24752,N_24228);
and U26755 (N_26755,N_24094,N_25554);
xor U26756 (N_26756,N_25996,N_24439);
xor U26757 (N_26757,N_24617,N_25548);
and U26758 (N_26758,N_24253,N_25395);
nand U26759 (N_26759,N_25709,N_25235);
nor U26760 (N_26760,N_25453,N_25772);
or U26761 (N_26761,N_24374,N_25846);
or U26762 (N_26762,N_24548,N_25193);
nand U26763 (N_26763,N_25777,N_25965);
nor U26764 (N_26764,N_24784,N_25676);
nor U26765 (N_26765,N_24308,N_25088);
nor U26766 (N_26766,N_24222,N_24706);
or U26767 (N_26767,N_25075,N_25182);
xnor U26768 (N_26768,N_24322,N_25386);
nand U26769 (N_26769,N_25898,N_24406);
xor U26770 (N_26770,N_24846,N_25630);
xor U26771 (N_26771,N_25450,N_25525);
and U26772 (N_26772,N_25835,N_25312);
and U26773 (N_26773,N_24947,N_25745);
and U26774 (N_26774,N_24826,N_25666);
nor U26775 (N_26775,N_24005,N_25315);
or U26776 (N_26776,N_25263,N_25253);
and U26777 (N_26777,N_25719,N_24476);
xor U26778 (N_26778,N_24899,N_25927);
or U26779 (N_26779,N_25962,N_24944);
or U26780 (N_26780,N_25357,N_24663);
nor U26781 (N_26781,N_25879,N_24866);
or U26782 (N_26782,N_24054,N_24419);
xor U26783 (N_26783,N_24373,N_24739);
xor U26784 (N_26784,N_25567,N_25863);
or U26785 (N_26785,N_24260,N_25897);
xor U26786 (N_26786,N_24687,N_25089);
nor U26787 (N_26787,N_24767,N_24935);
nor U26788 (N_26788,N_25487,N_25884);
xnor U26789 (N_26789,N_25995,N_24801);
or U26790 (N_26790,N_24960,N_24639);
nor U26791 (N_26791,N_24280,N_25269);
nand U26792 (N_26792,N_25628,N_25773);
or U26793 (N_26793,N_24334,N_24971);
xor U26794 (N_26794,N_24516,N_25106);
and U26795 (N_26795,N_25967,N_24240);
nand U26796 (N_26796,N_24411,N_25318);
nand U26797 (N_26797,N_24729,N_25739);
or U26798 (N_26798,N_25016,N_24962);
xor U26799 (N_26799,N_24755,N_24515);
nor U26800 (N_26800,N_24818,N_25576);
nor U26801 (N_26801,N_25494,N_25222);
nand U26802 (N_26802,N_24965,N_25361);
nand U26803 (N_26803,N_24057,N_24810);
nand U26804 (N_26804,N_25664,N_25971);
or U26805 (N_26805,N_25960,N_25452);
or U26806 (N_26806,N_25286,N_25947);
and U26807 (N_26807,N_25934,N_25192);
xor U26808 (N_26808,N_24061,N_25160);
or U26809 (N_26809,N_24355,N_25181);
xor U26810 (N_26810,N_24897,N_25219);
or U26811 (N_26811,N_25531,N_24807);
and U26812 (N_26812,N_25447,N_24020);
nand U26813 (N_26813,N_24631,N_24740);
or U26814 (N_26814,N_25211,N_24258);
nand U26815 (N_26815,N_25460,N_24172);
and U26816 (N_26816,N_25980,N_25463);
nand U26817 (N_26817,N_24893,N_25427);
xnor U26818 (N_26818,N_24983,N_24762);
nand U26819 (N_26819,N_25837,N_25569);
nor U26820 (N_26820,N_24969,N_25476);
nor U26821 (N_26821,N_25002,N_25005);
or U26822 (N_26822,N_25850,N_24340);
nor U26823 (N_26823,N_24621,N_25382);
nor U26824 (N_26824,N_25448,N_25858);
or U26825 (N_26825,N_25706,N_24442);
xnor U26826 (N_26826,N_25928,N_24978);
or U26827 (N_26827,N_24689,N_25838);
nor U26828 (N_26828,N_25381,N_25880);
and U26829 (N_26829,N_24036,N_24834);
nor U26830 (N_26830,N_25623,N_24075);
nand U26831 (N_26831,N_25655,N_25677);
and U26832 (N_26832,N_24000,N_24460);
and U26833 (N_26833,N_25314,N_25942);
nor U26834 (N_26834,N_24130,N_25558);
nand U26835 (N_26835,N_25613,N_25307);
and U26836 (N_26836,N_24333,N_25344);
xor U26837 (N_26837,N_25150,N_25611);
xor U26838 (N_26838,N_24164,N_25437);
or U26839 (N_26839,N_25802,N_25122);
nand U26840 (N_26840,N_24802,N_25365);
or U26841 (N_26841,N_25117,N_24604);
or U26842 (N_26842,N_25389,N_24880);
nor U26843 (N_26843,N_25107,N_25796);
nor U26844 (N_26844,N_25915,N_25654);
nor U26845 (N_26845,N_25673,N_24122);
nand U26846 (N_26846,N_24997,N_24670);
and U26847 (N_26847,N_25888,N_25135);
and U26848 (N_26848,N_24370,N_24250);
nand U26849 (N_26849,N_25786,N_25890);
nor U26850 (N_26850,N_24383,N_24231);
or U26851 (N_26851,N_24234,N_24481);
nand U26852 (N_26852,N_24214,N_25254);
nor U26853 (N_26853,N_25963,N_25380);
and U26854 (N_26854,N_24209,N_25941);
nor U26855 (N_26855,N_25867,N_25411);
nand U26856 (N_26856,N_25143,N_24469);
nor U26857 (N_26857,N_24615,N_25288);
or U26858 (N_26858,N_24081,N_24996);
nand U26859 (N_26859,N_25103,N_24328);
xor U26860 (N_26860,N_25101,N_25946);
nor U26861 (N_26861,N_25132,N_25519);
nor U26862 (N_26862,N_24922,N_25392);
or U26863 (N_26863,N_24468,N_25648);
and U26864 (N_26864,N_25176,N_24241);
and U26865 (N_26865,N_24110,N_25902);
xnor U26866 (N_26866,N_25935,N_24421);
and U26867 (N_26867,N_24033,N_24487);
and U26868 (N_26868,N_25674,N_25285);
nor U26869 (N_26869,N_24289,N_24107);
nor U26870 (N_26870,N_25598,N_24936);
nand U26871 (N_26871,N_24756,N_24085);
nor U26872 (N_26872,N_25903,N_25565);
xor U26873 (N_26873,N_25037,N_24895);
xnor U26874 (N_26874,N_24574,N_25325);
xnor U26875 (N_26875,N_25166,N_25820);
and U26876 (N_26876,N_24138,N_25698);
nand U26877 (N_26877,N_25099,N_24226);
xnor U26878 (N_26878,N_24128,N_24432);
xor U26879 (N_26879,N_25028,N_24078);
or U26880 (N_26880,N_24824,N_25290);
nor U26881 (N_26881,N_25711,N_25809);
nand U26882 (N_26882,N_25816,N_24160);
nand U26883 (N_26883,N_24216,N_24343);
or U26884 (N_26884,N_24259,N_24215);
or U26885 (N_26885,N_25172,N_25874);
nand U26886 (N_26886,N_24789,N_24677);
nor U26887 (N_26887,N_25661,N_24082);
or U26888 (N_26888,N_25187,N_24943);
nand U26889 (N_26889,N_25518,N_24162);
nand U26890 (N_26890,N_24457,N_24905);
or U26891 (N_26891,N_24511,N_25830);
nand U26892 (N_26892,N_24587,N_25899);
nand U26893 (N_26893,N_25992,N_25794);
or U26894 (N_26894,N_24294,N_25645);
nand U26895 (N_26895,N_25436,N_25825);
xnor U26896 (N_26896,N_25485,N_25616);
and U26897 (N_26897,N_25970,N_25236);
nor U26898 (N_26898,N_24276,N_25752);
or U26899 (N_26899,N_25793,N_24407);
nor U26900 (N_26900,N_25113,N_24939);
nand U26901 (N_26901,N_24902,N_24306);
nor U26902 (N_26902,N_25873,N_25881);
and U26903 (N_26903,N_25778,N_25998);
nor U26904 (N_26904,N_24431,N_25032);
xnor U26905 (N_26905,N_24022,N_25955);
nor U26906 (N_26906,N_25755,N_25807);
or U26907 (N_26907,N_24871,N_24814);
nand U26908 (N_26908,N_25704,N_25563);
or U26909 (N_26909,N_24091,N_24120);
nor U26910 (N_26910,N_25920,N_25985);
or U26911 (N_26911,N_24168,N_25024);
nand U26912 (N_26912,N_24694,N_24424);
nor U26913 (N_26913,N_24195,N_24678);
or U26914 (N_26914,N_24025,N_24913);
nand U26915 (N_26915,N_25499,N_24952);
and U26916 (N_26916,N_25716,N_25840);
or U26917 (N_26917,N_24693,N_24146);
or U26918 (N_26918,N_24722,N_25004);
and U26919 (N_26919,N_24092,N_25208);
or U26920 (N_26920,N_24979,N_24651);
nand U26921 (N_26921,N_24157,N_24461);
xnor U26922 (N_26922,N_25972,N_25241);
xnor U26923 (N_26923,N_25264,N_25340);
nor U26924 (N_26924,N_25205,N_25126);
nor U26925 (N_26925,N_25214,N_24599);
nand U26926 (N_26926,N_25104,N_24588);
xor U26927 (N_26927,N_24799,N_25689);
or U26928 (N_26928,N_24753,N_25310);
or U26929 (N_26929,N_24089,N_25503);
nor U26930 (N_26930,N_25892,N_25022);
nor U26931 (N_26931,N_24463,N_24412);
nand U26932 (N_26932,N_24855,N_25319);
and U26933 (N_26933,N_24409,N_25685);
nand U26934 (N_26934,N_25818,N_25819);
xnor U26935 (N_26935,N_25128,N_25428);
nor U26936 (N_26936,N_25120,N_25461);
or U26937 (N_26937,N_24698,N_25451);
nor U26938 (N_26938,N_25050,N_24113);
nor U26939 (N_26939,N_24987,N_24811);
xnor U26940 (N_26940,N_24192,N_24868);
nand U26941 (N_26941,N_24492,N_25990);
nor U26942 (N_26942,N_24205,N_24313);
xor U26943 (N_26943,N_24065,N_25954);
nand U26944 (N_26944,N_24140,N_25977);
nor U26945 (N_26945,N_25799,N_24909);
or U26946 (N_26946,N_25468,N_25784);
xnor U26947 (N_26947,N_25672,N_25805);
nor U26948 (N_26948,N_25642,N_24225);
or U26949 (N_26949,N_25455,N_24970);
nor U26950 (N_26950,N_24964,N_24119);
xnor U26951 (N_26951,N_25605,N_24643);
nor U26952 (N_26952,N_25983,N_25034);
nand U26953 (N_26953,N_25491,N_25602);
nor U26954 (N_26954,N_25348,N_24010);
nand U26955 (N_26955,N_25020,N_24819);
and U26956 (N_26956,N_25544,N_25047);
nor U26957 (N_26957,N_24841,N_24397);
nor U26958 (N_26958,N_25021,N_24510);
xor U26959 (N_26959,N_25425,N_25937);
nand U26960 (N_26960,N_25986,N_24450);
and U26961 (N_26961,N_25391,N_24610);
or U26962 (N_26962,N_25497,N_25291);
nand U26963 (N_26963,N_24153,N_24351);
nand U26964 (N_26964,N_24589,N_25042);
xnor U26965 (N_26965,N_24465,N_24063);
nor U26966 (N_26966,N_24657,N_25014);
nand U26967 (N_26967,N_25713,N_24700);
or U26968 (N_26968,N_25401,N_25112);
or U26969 (N_26969,N_25950,N_24705);
xnor U26970 (N_26970,N_25299,N_24761);
nand U26971 (N_26971,N_25564,N_25486);
and U26972 (N_26972,N_25822,N_25536);
and U26973 (N_26973,N_25198,N_24404);
or U26974 (N_26974,N_25337,N_25520);
nand U26975 (N_26975,N_24279,N_24731);
nor U26976 (N_26976,N_25231,N_24186);
nand U26977 (N_26977,N_24428,N_25188);
nor U26978 (N_26978,N_24232,N_24443);
and U26979 (N_26979,N_24613,N_24349);
or U26980 (N_26980,N_25360,N_24150);
xor U26981 (N_26981,N_25756,N_24382);
nor U26982 (N_26982,N_24474,N_25815);
or U26983 (N_26983,N_24735,N_25001);
or U26984 (N_26984,N_25924,N_24167);
or U26985 (N_26985,N_25228,N_25258);
nor U26986 (N_26986,N_25911,N_25832);
xnor U26987 (N_26987,N_24534,N_24165);
nand U26988 (N_26988,N_25221,N_24462);
and U26989 (N_26989,N_24955,N_24277);
nand U26990 (N_26990,N_24505,N_25750);
nor U26991 (N_26991,N_24724,N_24797);
xor U26992 (N_26992,N_25826,N_24493);
or U26993 (N_26993,N_24840,N_24100);
nand U26994 (N_26994,N_24945,N_25237);
xnor U26995 (N_26995,N_24118,N_24733);
xor U26996 (N_26996,N_24156,N_24886);
nor U26997 (N_26997,N_24180,N_25233);
nor U26998 (N_26998,N_24337,N_25639);
nor U26999 (N_26999,N_24224,N_24077);
or U27000 (N_27000,N_25075,N_24627);
xor U27001 (N_27001,N_25741,N_25453);
nor U27002 (N_27002,N_25959,N_25937);
xor U27003 (N_27003,N_24936,N_25881);
or U27004 (N_27004,N_25529,N_24884);
xnor U27005 (N_27005,N_24810,N_24911);
nor U27006 (N_27006,N_24892,N_24957);
nand U27007 (N_27007,N_25304,N_25104);
and U27008 (N_27008,N_24005,N_24214);
nand U27009 (N_27009,N_24549,N_25056);
and U27010 (N_27010,N_24859,N_24507);
or U27011 (N_27011,N_25892,N_24986);
or U27012 (N_27012,N_24637,N_24263);
nand U27013 (N_27013,N_24035,N_24334);
or U27014 (N_27014,N_25756,N_25659);
xnor U27015 (N_27015,N_25630,N_24745);
nor U27016 (N_27016,N_25284,N_25156);
nand U27017 (N_27017,N_24745,N_25019);
and U27018 (N_27018,N_25333,N_24695);
xnor U27019 (N_27019,N_24004,N_25800);
xor U27020 (N_27020,N_24617,N_25245);
and U27021 (N_27021,N_24227,N_24885);
nand U27022 (N_27022,N_25908,N_25619);
nand U27023 (N_27023,N_25661,N_25686);
and U27024 (N_27024,N_25316,N_25782);
xnor U27025 (N_27025,N_25349,N_25588);
nand U27026 (N_27026,N_25198,N_24552);
and U27027 (N_27027,N_24163,N_24153);
nand U27028 (N_27028,N_24689,N_24612);
and U27029 (N_27029,N_25425,N_24549);
or U27030 (N_27030,N_24829,N_25028);
nand U27031 (N_27031,N_25547,N_25684);
nand U27032 (N_27032,N_25163,N_24138);
or U27033 (N_27033,N_25729,N_25066);
nand U27034 (N_27034,N_24717,N_24123);
nand U27035 (N_27035,N_25489,N_24984);
xnor U27036 (N_27036,N_24831,N_25777);
or U27037 (N_27037,N_24657,N_24254);
xnor U27038 (N_27038,N_25720,N_24912);
nand U27039 (N_27039,N_25281,N_24151);
nand U27040 (N_27040,N_24994,N_25347);
xor U27041 (N_27041,N_25575,N_25278);
nor U27042 (N_27042,N_25120,N_25177);
or U27043 (N_27043,N_25053,N_25661);
or U27044 (N_27044,N_25178,N_24132);
nor U27045 (N_27045,N_25127,N_25032);
nor U27046 (N_27046,N_25718,N_25272);
nor U27047 (N_27047,N_25546,N_25352);
xor U27048 (N_27048,N_25143,N_25228);
nor U27049 (N_27049,N_24037,N_24909);
nand U27050 (N_27050,N_25382,N_25719);
xnor U27051 (N_27051,N_24103,N_24994);
or U27052 (N_27052,N_25097,N_24094);
or U27053 (N_27053,N_25727,N_25413);
and U27054 (N_27054,N_25625,N_25445);
xnor U27055 (N_27055,N_25845,N_24495);
or U27056 (N_27056,N_25128,N_24019);
xnor U27057 (N_27057,N_24343,N_25184);
xor U27058 (N_27058,N_24329,N_24667);
and U27059 (N_27059,N_24544,N_25069);
nor U27060 (N_27060,N_25238,N_24389);
nand U27061 (N_27061,N_25402,N_24036);
nand U27062 (N_27062,N_25587,N_24443);
and U27063 (N_27063,N_25884,N_25768);
xnor U27064 (N_27064,N_24877,N_24501);
nor U27065 (N_27065,N_25075,N_25426);
nand U27066 (N_27066,N_25085,N_24723);
nand U27067 (N_27067,N_24006,N_25733);
nor U27068 (N_27068,N_25104,N_24148);
xnor U27069 (N_27069,N_25929,N_24885);
nand U27070 (N_27070,N_24352,N_25099);
and U27071 (N_27071,N_24903,N_24310);
nor U27072 (N_27072,N_25317,N_25092);
and U27073 (N_27073,N_25270,N_24172);
and U27074 (N_27074,N_24074,N_25004);
and U27075 (N_27075,N_25843,N_24778);
and U27076 (N_27076,N_24257,N_24601);
or U27077 (N_27077,N_24032,N_24033);
and U27078 (N_27078,N_25843,N_25329);
or U27079 (N_27079,N_25014,N_25398);
nor U27080 (N_27080,N_25913,N_24136);
nor U27081 (N_27081,N_25240,N_24582);
xnor U27082 (N_27082,N_25317,N_24289);
xnor U27083 (N_27083,N_24159,N_25821);
nor U27084 (N_27084,N_24420,N_25972);
nor U27085 (N_27085,N_24693,N_25589);
or U27086 (N_27086,N_25067,N_25616);
or U27087 (N_27087,N_25102,N_25761);
nand U27088 (N_27088,N_24020,N_24693);
nor U27089 (N_27089,N_24244,N_24004);
nand U27090 (N_27090,N_25538,N_24142);
nor U27091 (N_27091,N_25080,N_25108);
nand U27092 (N_27092,N_25672,N_24909);
nand U27093 (N_27093,N_24331,N_25357);
nor U27094 (N_27094,N_25550,N_24535);
xnor U27095 (N_27095,N_25762,N_25742);
nand U27096 (N_27096,N_24550,N_25542);
xnor U27097 (N_27097,N_24991,N_25014);
xor U27098 (N_27098,N_24326,N_25473);
xor U27099 (N_27099,N_24636,N_24151);
xor U27100 (N_27100,N_25401,N_25535);
or U27101 (N_27101,N_25797,N_25984);
xor U27102 (N_27102,N_24268,N_24793);
xor U27103 (N_27103,N_24574,N_25942);
xnor U27104 (N_27104,N_24121,N_24834);
nand U27105 (N_27105,N_25991,N_24172);
or U27106 (N_27106,N_25299,N_25698);
nand U27107 (N_27107,N_25045,N_25951);
nand U27108 (N_27108,N_24801,N_24606);
xor U27109 (N_27109,N_25637,N_24371);
nor U27110 (N_27110,N_25958,N_25104);
nor U27111 (N_27111,N_24867,N_25404);
or U27112 (N_27112,N_25692,N_24960);
or U27113 (N_27113,N_25746,N_25502);
nand U27114 (N_27114,N_25672,N_25841);
nand U27115 (N_27115,N_24141,N_24800);
xor U27116 (N_27116,N_25715,N_25617);
or U27117 (N_27117,N_25146,N_25632);
and U27118 (N_27118,N_25820,N_24482);
and U27119 (N_27119,N_24363,N_25945);
nor U27120 (N_27120,N_25531,N_25292);
and U27121 (N_27121,N_24884,N_25126);
and U27122 (N_27122,N_24002,N_25093);
xor U27123 (N_27123,N_24287,N_24659);
nand U27124 (N_27124,N_24496,N_24559);
and U27125 (N_27125,N_24947,N_25731);
nor U27126 (N_27126,N_25151,N_24540);
or U27127 (N_27127,N_24179,N_25223);
nand U27128 (N_27128,N_25677,N_25235);
or U27129 (N_27129,N_24887,N_25432);
and U27130 (N_27130,N_24472,N_24424);
xnor U27131 (N_27131,N_25623,N_25545);
and U27132 (N_27132,N_25541,N_25374);
nor U27133 (N_27133,N_25188,N_25249);
nand U27134 (N_27134,N_24693,N_25822);
nor U27135 (N_27135,N_25163,N_25771);
nor U27136 (N_27136,N_25529,N_24458);
xor U27137 (N_27137,N_24851,N_25664);
xnor U27138 (N_27138,N_24064,N_24428);
or U27139 (N_27139,N_24062,N_24143);
nor U27140 (N_27140,N_24469,N_24725);
xor U27141 (N_27141,N_24580,N_25219);
and U27142 (N_27142,N_24591,N_24804);
nand U27143 (N_27143,N_24487,N_24999);
nor U27144 (N_27144,N_25726,N_25512);
nor U27145 (N_27145,N_25903,N_24833);
nor U27146 (N_27146,N_24992,N_24420);
xor U27147 (N_27147,N_24233,N_24845);
and U27148 (N_27148,N_24317,N_24206);
nor U27149 (N_27149,N_24002,N_24341);
and U27150 (N_27150,N_25374,N_25385);
and U27151 (N_27151,N_24702,N_24520);
nand U27152 (N_27152,N_25478,N_24540);
or U27153 (N_27153,N_24114,N_25152);
and U27154 (N_27154,N_24354,N_24668);
nor U27155 (N_27155,N_25060,N_25348);
nor U27156 (N_27156,N_25389,N_25882);
xor U27157 (N_27157,N_24581,N_25320);
or U27158 (N_27158,N_24337,N_24091);
nand U27159 (N_27159,N_24895,N_24201);
nand U27160 (N_27160,N_24921,N_25389);
or U27161 (N_27161,N_24112,N_25969);
nand U27162 (N_27162,N_25966,N_24044);
nor U27163 (N_27163,N_24200,N_24477);
nor U27164 (N_27164,N_25875,N_24864);
or U27165 (N_27165,N_24697,N_25353);
and U27166 (N_27166,N_24052,N_25837);
and U27167 (N_27167,N_25895,N_25777);
nor U27168 (N_27168,N_24341,N_25695);
xnor U27169 (N_27169,N_25468,N_24352);
nand U27170 (N_27170,N_25542,N_25087);
nor U27171 (N_27171,N_25101,N_24149);
nand U27172 (N_27172,N_25959,N_25631);
nor U27173 (N_27173,N_24180,N_25253);
nand U27174 (N_27174,N_25337,N_25007);
nor U27175 (N_27175,N_25915,N_25552);
nand U27176 (N_27176,N_25484,N_24375);
xnor U27177 (N_27177,N_24836,N_24977);
xnor U27178 (N_27178,N_25689,N_25507);
xor U27179 (N_27179,N_24661,N_25135);
and U27180 (N_27180,N_24565,N_25419);
and U27181 (N_27181,N_25115,N_25081);
and U27182 (N_27182,N_24999,N_24866);
xnor U27183 (N_27183,N_25752,N_25423);
nand U27184 (N_27184,N_24341,N_24961);
and U27185 (N_27185,N_25049,N_24607);
xnor U27186 (N_27186,N_25531,N_25666);
or U27187 (N_27187,N_25994,N_25606);
or U27188 (N_27188,N_24966,N_25248);
nand U27189 (N_27189,N_25382,N_24128);
nand U27190 (N_27190,N_24826,N_24733);
xor U27191 (N_27191,N_25469,N_24597);
and U27192 (N_27192,N_25221,N_24476);
and U27193 (N_27193,N_24488,N_24375);
nor U27194 (N_27194,N_25373,N_24978);
xor U27195 (N_27195,N_25413,N_25788);
nor U27196 (N_27196,N_24403,N_24237);
xnor U27197 (N_27197,N_25050,N_24865);
xor U27198 (N_27198,N_25386,N_25151);
xnor U27199 (N_27199,N_24631,N_24224);
nor U27200 (N_27200,N_25252,N_25719);
nor U27201 (N_27201,N_25191,N_24727);
nor U27202 (N_27202,N_24865,N_24611);
nor U27203 (N_27203,N_25702,N_24236);
nand U27204 (N_27204,N_24681,N_25380);
nor U27205 (N_27205,N_25830,N_25083);
nand U27206 (N_27206,N_24254,N_24763);
nand U27207 (N_27207,N_25799,N_24227);
or U27208 (N_27208,N_24308,N_25465);
nor U27209 (N_27209,N_24346,N_24653);
or U27210 (N_27210,N_25701,N_24495);
nor U27211 (N_27211,N_25715,N_24157);
nor U27212 (N_27212,N_24991,N_25371);
or U27213 (N_27213,N_24863,N_25197);
and U27214 (N_27214,N_24835,N_24799);
nor U27215 (N_27215,N_24389,N_24435);
or U27216 (N_27216,N_25290,N_24679);
nor U27217 (N_27217,N_25003,N_25327);
nor U27218 (N_27218,N_25402,N_25569);
nand U27219 (N_27219,N_24398,N_24268);
nor U27220 (N_27220,N_25159,N_24379);
nand U27221 (N_27221,N_24463,N_25269);
or U27222 (N_27222,N_25350,N_25632);
nor U27223 (N_27223,N_25046,N_24960);
xor U27224 (N_27224,N_25529,N_25664);
or U27225 (N_27225,N_25591,N_24291);
nand U27226 (N_27226,N_25689,N_24330);
xor U27227 (N_27227,N_25681,N_24391);
nor U27228 (N_27228,N_24683,N_24622);
nor U27229 (N_27229,N_25878,N_24224);
or U27230 (N_27230,N_25362,N_25313);
xor U27231 (N_27231,N_25411,N_25006);
xnor U27232 (N_27232,N_24247,N_24356);
nor U27233 (N_27233,N_24853,N_25860);
or U27234 (N_27234,N_24957,N_24308);
nand U27235 (N_27235,N_25619,N_24293);
nand U27236 (N_27236,N_24068,N_25706);
xnor U27237 (N_27237,N_24207,N_24025);
or U27238 (N_27238,N_24866,N_24822);
or U27239 (N_27239,N_25524,N_24719);
or U27240 (N_27240,N_25311,N_24901);
or U27241 (N_27241,N_24631,N_24859);
nor U27242 (N_27242,N_25148,N_25209);
or U27243 (N_27243,N_24722,N_24914);
nor U27244 (N_27244,N_24158,N_24698);
and U27245 (N_27245,N_25609,N_24449);
xor U27246 (N_27246,N_24570,N_25078);
xnor U27247 (N_27247,N_25829,N_24799);
or U27248 (N_27248,N_24607,N_25121);
and U27249 (N_27249,N_25048,N_25595);
nand U27250 (N_27250,N_24571,N_25973);
nor U27251 (N_27251,N_25732,N_25296);
xnor U27252 (N_27252,N_24680,N_25654);
or U27253 (N_27253,N_25622,N_24340);
nor U27254 (N_27254,N_25140,N_24081);
xnor U27255 (N_27255,N_25385,N_25167);
xnor U27256 (N_27256,N_25068,N_25606);
nand U27257 (N_27257,N_25655,N_24085);
and U27258 (N_27258,N_25510,N_25994);
xor U27259 (N_27259,N_24955,N_24507);
nor U27260 (N_27260,N_24820,N_25053);
xnor U27261 (N_27261,N_25726,N_24908);
xnor U27262 (N_27262,N_24406,N_24508);
or U27263 (N_27263,N_24176,N_24789);
and U27264 (N_27264,N_25004,N_25630);
nand U27265 (N_27265,N_25457,N_24358);
or U27266 (N_27266,N_25808,N_25469);
or U27267 (N_27267,N_24548,N_24150);
and U27268 (N_27268,N_24603,N_24859);
nand U27269 (N_27269,N_24860,N_25367);
and U27270 (N_27270,N_24287,N_25912);
nand U27271 (N_27271,N_25575,N_25693);
and U27272 (N_27272,N_24967,N_24692);
xor U27273 (N_27273,N_25737,N_25313);
xor U27274 (N_27274,N_25174,N_24851);
or U27275 (N_27275,N_24861,N_25934);
nor U27276 (N_27276,N_25077,N_24166);
nor U27277 (N_27277,N_24178,N_24405);
nand U27278 (N_27278,N_25223,N_24829);
and U27279 (N_27279,N_24303,N_24537);
or U27280 (N_27280,N_25449,N_25386);
nand U27281 (N_27281,N_25629,N_25758);
nor U27282 (N_27282,N_25488,N_24463);
and U27283 (N_27283,N_25314,N_25658);
and U27284 (N_27284,N_25213,N_24753);
or U27285 (N_27285,N_24923,N_24005);
nor U27286 (N_27286,N_25003,N_24321);
or U27287 (N_27287,N_24839,N_24219);
and U27288 (N_27288,N_25167,N_24764);
xor U27289 (N_27289,N_25981,N_25716);
or U27290 (N_27290,N_25140,N_25630);
xnor U27291 (N_27291,N_24925,N_25176);
or U27292 (N_27292,N_24830,N_25454);
nand U27293 (N_27293,N_24768,N_24820);
or U27294 (N_27294,N_24332,N_25980);
nand U27295 (N_27295,N_25464,N_25441);
or U27296 (N_27296,N_24203,N_24180);
nor U27297 (N_27297,N_24484,N_25763);
nor U27298 (N_27298,N_24466,N_24706);
nor U27299 (N_27299,N_24470,N_24159);
and U27300 (N_27300,N_25138,N_25171);
nand U27301 (N_27301,N_24754,N_25668);
xor U27302 (N_27302,N_25296,N_25214);
or U27303 (N_27303,N_24022,N_25581);
or U27304 (N_27304,N_24526,N_24393);
or U27305 (N_27305,N_25323,N_24688);
or U27306 (N_27306,N_25928,N_24931);
nor U27307 (N_27307,N_25792,N_25626);
nor U27308 (N_27308,N_24456,N_25088);
nand U27309 (N_27309,N_25235,N_25361);
or U27310 (N_27310,N_24143,N_25522);
and U27311 (N_27311,N_25691,N_25211);
xor U27312 (N_27312,N_24780,N_24175);
or U27313 (N_27313,N_24488,N_25680);
and U27314 (N_27314,N_24308,N_24692);
nand U27315 (N_27315,N_24314,N_24004);
or U27316 (N_27316,N_24192,N_24592);
or U27317 (N_27317,N_24833,N_25103);
and U27318 (N_27318,N_24229,N_24236);
and U27319 (N_27319,N_25900,N_25744);
and U27320 (N_27320,N_25155,N_24193);
nor U27321 (N_27321,N_25663,N_24825);
and U27322 (N_27322,N_24062,N_25056);
and U27323 (N_27323,N_24760,N_25326);
nor U27324 (N_27324,N_25024,N_24815);
nor U27325 (N_27325,N_25242,N_25861);
xnor U27326 (N_27326,N_25646,N_24589);
nand U27327 (N_27327,N_25499,N_24006);
or U27328 (N_27328,N_24129,N_25712);
and U27329 (N_27329,N_24089,N_25244);
and U27330 (N_27330,N_25402,N_25755);
nor U27331 (N_27331,N_24982,N_24340);
xnor U27332 (N_27332,N_24281,N_25052);
or U27333 (N_27333,N_25590,N_24323);
nand U27334 (N_27334,N_24810,N_25140);
nor U27335 (N_27335,N_25268,N_24614);
xnor U27336 (N_27336,N_24472,N_24540);
nand U27337 (N_27337,N_25317,N_25289);
and U27338 (N_27338,N_25111,N_24725);
xor U27339 (N_27339,N_25684,N_25437);
and U27340 (N_27340,N_24058,N_25833);
xnor U27341 (N_27341,N_24678,N_24942);
xor U27342 (N_27342,N_25885,N_25312);
xnor U27343 (N_27343,N_25255,N_24794);
or U27344 (N_27344,N_25158,N_25909);
nor U27345 (N_27345,N_24663,N_24441);
nand U27346 (N_27346,N_24825,N_25747);
xnor U27347 (N_27347,N_24646,N_25956);
nand U27348 (N_27348,N_24701,N_25330);
nor U27349 (N_27349,N_24637,N_25627);
nand U27350 (N_27350,N_24645,N_24815);
nor U27351 (N_27351,N_25912,N_24630);
and U27352 (N_27352,N_25287,N_24036);
nor U27353 (N_27353,N_24541,N_25531);
xor U27354 (N_27354,N_25198,N_25576);
nor U27355 (N_27355,N_24944,N_25845);
or U27356 (N_27356,N_24141,N_25407);
xnor U27357 (N_27357,N_24584,N_24261);
and U27358 (N_27358,N_24425,N_24875);
or U27359 (N_27359,N_24234,N_25716);
xnor U27360 (N_27360,N_24192,N_24328);
xnor U27361 (N_27361,N_24007,N_25884);
nor U27362 (N_27362,N_24374,N_24277);
nor U27363 (N_27363,N_24816,N_24211);
and U27364 (N_27364,N_24893,N_24629);
xnor U27365 (N_27365,N_24290,N_25042);
nor U27366 (N_27366,N_25694,N_24727);
or U27367 (N_27367,N_24538,N_24674);
and U27368 (N_27368,N_25307,N_25974);
or U27369 (N_27369,N_24033,N_25977);
and U27370 (N_27370,N_25881,N_24150);
and U27371 (N_27371,N_25962,N_25541);
nor U27372 (N_27372,N_24261,N_24273);
nor U27373 (N_27373,N_25530,N_24217);
or U27374 (N_27374,N_24575,N_25917);
or U27375 (N_27375,N_24699,N_24077);
xor U27376 (N_27376,N_25174,N_24291);
and U27377 (N_27377,N_24747,N_25388);
nor U27378 (N_27378,N_24806,N_25884);
nand U27379 (N_27379,N_25985,N_25984);
nor U27380 (N_27380,N_24952,N_24126);
and U27381 (N_27381,N_24809,N_24752);
nand U27382 (N_27382,N_24836,N_24027);
nor U27383 (N_27383,N_24860,N_25872);
xnor U27384 (N_27384,N_25543,N_25733);
or U27385 (N_27385,N_25323,N_25701);
and U27386 (N_27386,N_25810,N_24823);
nor U27387 (N_27387,N_25655,N_25350);
nor U27388 (N_27388,N_24131,N_24450);
and U27389 (N_27389,N_25195,N_25162);
xnor U27390 (N_27390,N_25032,N_25190);
and U27391 (N_27391,N_24316,N_25432);
nand U27392 (N_27392,N_24602,N_24270);
or U27393 (N_27393,N_24646,N_24133);
nand U27394 (N_27394,N_25536,N_25026);
nand U27395 (N_27395,N_25662,N_24746);
xor U27396 (N_27396,N_24747,N_25327);
and U27397 (N_27397,N_24366,N_24588);
and U27398 (N_27398,N_25612,N_25534);
and U27399 (N_27399,N_24698,N_24188);
or U27400 (N_27400,N_25488,N_24216);
and U27401 (N_27401,N_24770,N_25772);
nand U27402 (N_27402,N_25100,N_25706);
nor U27403 (N_27403,N_24304,N_25162);
xnor U27404 (N_27404,N_25006,N_25152);
xor U27405 (N_27405,N_25018,N_25435);
or U27406 (N_27406,N_24913,N_24483);
xor U27407 (N_27407,N_24088,N_24315);
or U27408 (N_27408,N_25356,N_24686);
xnor U27409 (N_27409,N_25482,N_24075);
nand U27410 (N_27410,N_24940,N_24623);
and U27411 (N_27411,N_24806,N_25525);
nand U27412 (N_27412,N_25592,N_24895);
or U27413 (N_27413,N_25621,N_24200);
nand U27414 (N_27414,N_25355,N_25642);
or U27415 (N_27415,N_25485,N_24717);
nor U27416 (N_27416,N_25165,N_25060);
nor U27417 (N_27417,N_24767,N_24222);
xor U27418 (N_27418,N_24915,N_25215);
nand U27419 (N_27419,N_24246,N_24615);
xor U27420 (N_27420,N_24124,N_24524);
nand U27421 (N_27421,N_24572,N_24374);
and U27422 (N_27422,N_25042,N_24128);
xnor U27423 (N_27423,N_25770,N_25010);
and U27424 (N_27424,N_24316,N_25525);
and U27425 (N_27425,N_24554,N_24482);
or U27426 (N_27426,N_25091,N_25200);
nor U27427 (N_27427,N_25291,N_25287);
xnor U27428 (N_27428,N_24988,N_25550);
and U27429 (N_27429,N_24619,N_24828);
and U27430 (N_27430,N_25314,N_25695);
nand U27431 (N_27431,N_25941,N_25448);
or U27432 (N_27432,N_24678,N_25304);
or U27433 (N_27433,N_24237,N_25272);
nor U27434 (N_27434,N_25719,N_24860);
nand U27435 (N_27435,N_24599,N_24486);
nand U27436 (N_27436,N_24861,N_25166);
or U27437 (N_27437,N_25914,N_25235);
and U27438 (N_27438,N_25131,N_25597);
or U27439 (N_27439,N_25956,N_25003);
and U27440 (N_27440,N_25258,N_24758);
nor U27441 (N_27441,N_24398,N_25205);
xnor U27442 (N_27442,N_24065,N_25044);
xor U27443 (N_27443,N_25702,N_25529);
nor U27444 (N_27444,N_25874,N_24285);
xor U27445 (N_27445,N_25321,N_25314);
or U27446 (N_27446,N_24012,N_24344);
nor U27447 (N_27447,N_24678,N_25780);
nor U27448 (N_27448,N_25059,N_24439);
xor U27449 (N_27449,N_25122,N_25537);
and U27450 (N_27450,N_24516,N_24434);
xnor U27451 (N_27451,N_25906,N_24753);
nor U27452 (N_27452,N_25478,N_24713);
and U27453 (N_27453,N_25607,N_25244);
nand U27454 (N_27454,N_24336,N_24524);
xnor U27455 (N_27455,N_25969,N_25085);
xnor U27456 (N_27456,N_25837,N_24563);
xnor U27457 (N_27457,N_25702,N_24483);
xor U27458 (N_27458,N_25442,N_24874);
nand U27459 (N_27459,N_24338,N_24082);
or U27460 (N_27460,N_25243,N_24736);
nor U27461 (N_27461,N_24799,N_24878);
nand U27462 (N_27462,N_24069,N_25386);
nor U27463 (N_27463,N_24690,N_25967);
xor U27464 (N_27464,N_25376,N_25398);
and U27465 (N_27465,N_24421,N_25477);
or U27466 (N_27466,N_24199,N_25122);
or U27467 (N_27467,N_25499,N_24436);
xnor U27468 (N_27468,N_24941,N_24623);
nand U27469 (N_27469,N_25186,N_24384);
nor U27470 (N_27470,N_25491,N_25562);
xnor U27471 (N_27471,N_25791,N_25442);
nor U27472 (N_27472,N_24579,N_24257);
nor U27473 (N_27473,N_25461,N_25479);
xor U27474 (N_27474,N_24066,N_24819);
nand U27475 (N_27475,N_24740,N_25642);
and U27476 (N_27476,N_25720,N_24854);
nand U27477 (N_27477,N_24865,N_25920);
xor U27478 (N_27478,N_24259,N_24522);
nor U27479 (N_27479,N_25536,N_25077);
nand U27480 (N_27480,N_24034,N_25677);
or U27481 (N_27481,N_24185,N_24518);
and U27482 (N_27482,N_25647,N_24728);
nor U27483 (N_27483,N_25660,N_25560);
nand U27484 (N_27484,N_25296,N_24884);
xnor U27485 (N_27485,N_25842,N_24174);
or U27486 (N_27486,N_24063,N_25477);
nor U27487 (N_27487,N_25952,N_25329);
xnor U27488 (N_27488,N_24972,N_25351);
and U27489 (N_27489,N_24392,N_25556);
nand U27490 (N_27490,N_25317,N_25462);
nand U27491 (N_27491,N_24990,N_24074);
and U27492 (N_27492,N_24464,N_24191);
nand U27493 (N_27493,N_24469,N_24348);
or U27494 (N_27494,N_24705,N_25444);
nand U27495 (N_27495,N_25435,N_24418);
or U27496 (N_27496,N_24092,N_25640);
and U27497 (N_27497,N_24363,N_25121);
xnor U27498 (N_27498,N_25699,N_24545);
nor U27499 (N_27499,N_24326,N_25915);
nand U27500 (N_27500,N_24498,N_24572);
and U27501 (N_27501,N_25706,N_24581);
xnor U27502 (N_27502,N_24173,N_24048);
xor U27503 (N_27503,N_25683,N_25855);
xnor U27504 (N_27504,N_24667,N_25266);
xnor U27505 (N_27505,N_24816,N_25841);
xnor U27506 (N_27506,N_25278,N_25064);
and U27507 (N_27507,N_25272,N_25003);
xor U27508 (N_27508,N_24397,N_25141);
nor U27509 (N_27509,N_24641,N_25018);
nand U27510 (N_27510,N_24955,N_25452);
nor U27511 (N_27511,N_24903,N_24375);
or U27512 (N_27512,N_25931,N_24364);
or U27513 (N_27513,N_24379,N_24001);
nand U27514 (N_27514,N_24214,N_25997);
xnor U27515 (N_27515,N_25216,N_24115);
and U27516 (N_27516,N_24342,N_25649);
and U27517 (N_27517,N_25545,N_25353);
and U27518 (N_27518,N_24704,N_24544);
xor U27519 (N_27519,N_25386,N_25408);
or U27520 (N_27520,N_25023,N_24381);
nand U27521 (N_27521,N_24729,N_24148);
or U27522 (N_27522,N_24425,N_24340);
nor U27523 (N_27523,N_24545,N_25379);
or U27524 (N_27524,N_25652,N_25817);
xnor U27525 (N_27525,N_25935,N_25748);
nand U27526 (N_27526,N_25895,N_25576);
nand U27527 (N_27527,N_25195,N_24953);
or U27528 (N_27528,N_24880,N_24968);
xor U27529 (N_27529,N_25696,N_24394);
or U27530 (N_27530,N_24575,N_25021);
or U27531 (N_27531,N_24913,N_24510);
and U27532 (N_27532,N_24977,N_24091);
nor U27533 (N_27533,N_24828,N_25492);
and U27534 (N_27534,N_25529,N_25022);
xnor U27535 (N_27535,N_25789,N_24602);
and U27536 (N_27536,N_24228,N_25643);
nor U27537 (N_27537,N_25501,N_25097);
xor U27538 (N_27538,N_24045,N_25766);
xnor U27539 (N_27539,N_24380,N_25342);
or U27540 (N_27540,N_25520,N_24731);
and U27541 (N_27541,N_24148,N_24684);
nor U27542 (N_27542,N_24152,N_24900);
or U27543 (N_27543,N_24945,N_25384);
nor U27544 (N_27544,N_25248,N_25831);
and U27545 (N_27545,N_24880,N_25035);
nand U27546 (N_27546,N_24137,N_24658);
or U27547 (N_27547,N_24028,N_25829);
and U27548 (N_27548,N_24226,N_25368);
nand U27549 (N_27549,N_24070,N_24297);
nor U27550 (N_27550,N_25602,N_25454);
and U27551 (N_27551,N_24716,N_25534);
xnor U27552 (N_27552,N_24664,N_24505);
nand U27553 (N_27553,N_25296,N_25543);
nor U27554 (N_27554,N_25653,N_25551);
and U27555 (N_27555,N_25714,N_25343);
nor U27556 (N_27556,N_25717,N_24841);
or U27557 (N_27557,N_24036,N_25128);
nor U27558 (N_27558,N_25061,N_25982);
nand U27559 (N_27559,N_24032,N_25819);
nand U27560 (N_27560,N_25418,N_25410);
xnor U27561 (N_27561,N_25283,N_25525);
and U27562 (N_27562,N_24528,N_24811);
nand U27563 (N_27563,N_25003,N_24675);
and U27564 (N_27564,N_25601,N_24272);
xnor U27565 (N_27565,N_25841,N_25479);
nor U27566 (N_27566,N_25098,N_25702);
nand U27567 (N_27567,N_25148,N_25247);
xnor U27568 (N_27568,N_25848,N_25629);
xor U27569 (N_27569,N_25791,N_25437);
and U27570 (N_27570,N_25335,N_24106);
nor U27571 (N_27571,N_24410,N_25341);
or U27572 (N_27572,N_25736,N_25274);
or U27573 (N_27573,N_25979,N_25028);
nor U27574 (N_27574,N_24229,N_25391);
nand U27575 (N_27575,N_24876,N_25442);
and U27576 (N_27576,N_25486,N_24108);
and U27577 (N_27577,N_25637,N_25725);
and U27578 (N_27578,N_25791,N_25208);
and U27579 (N_27579,N_25542,N_25533);
and U27580 (N_27580,N_25320,N_24289);
nor U27581 (N_27581,N_25829,N_25072);
xor U27582 (N_27582,N_25442,N_25516);
and U27583 (N_27583,N_24190,N_25659);
nand U27584 (N_27584,N_25986,N_24766);
and U27585 (N_27585,N_25647,N_24789);
and U27586 (N_27586,N_24923,N_25810);
xor U27587 (N_27587,N_25666,N_25003);
xnor U27588 (N_27588,N_24321,N_24712);
or U27589 (N_27589,N_25280,N_24351);
nor U27590 (N_27590,N_24712,N_24380);
nand U27591 (N_27591,N_24920,N_25629);
xor U27592 (N_27592,N_24649,N_25778);
or U27593 (N_27593,N_24329,N_24790);
and U27594 (N_27594,N_25227,N_24486);
xnor U27595 (N_27595,N_24040,N_24577);
nand U27596 (N_27596,N_24932,N_24490);
or U27597 (N_27597,N_25052,N_24487);
or U27598 (N_27598,N_25654,N_25220);
nor U27599 (N_27599,N_25326,N_25207);
or U27600 (N_27600,N_24241,N_24043);
nor U27601 (N_27601,N_25440,N_25026);
and U27602 (N_27602,N_24437,N_24692);
nor U27603 (N_27603,N_25966,N_25926);
or U27604 (N_27604,N_25612,N_25409);
nor U27605 (N_27605,N_25806,N_24758);
and U27606 (N_27606,N_24414,N_24920);
nand U27607 (N_27607,N_24655,N_24557);
nand U27608 (N_27608,N_24620,N_25306);
nor U27609 (N_27609,N_25195,N_25828);
xor U27610 (N_27610,N_25040,N_25274);
or U27611 (N_27611,N_25027,N_25400);
and U27612 (N_27612,N_25832,N_25295);
and U27613 (N_27613,N_25564,N_24041);
or U27614 (N_27614,N_25451,N_24494);
and U27615 (N_27615,N_24226,N_24925);
xnor U27616 (N_27616,N_25591,N_24848);
nand U27617 (N_27617,N_25246,N_24278);
or U27618 (N_27618,N_25556,N_25921);
or U27619 (N_27619,N_24306,N_24700);
and U27620 (N_27620,N_24147,N_24150);
xnor U27621 (N_27621,N_25700,N_25924);
xnor U27622 (N_27622,N_25553,N_24982);
xnor U27623 (N_27623,N_24493,N_25167);
nand U27624 (N_27624,N_24484,N_24510);
and U27625 (N_27625,N_24415,N_24760);
xor U27626 (N_27626,N_25865,N_24656);
xor U27627 (N_27627,N_25490,N_24500);
nand U27628 (N_27628,N_25881,N_25223);
and U27629 (N_27629,N_25862,N_25775);
and U27630 (N_27630,N_25151,N_24209);
and U27631 (N_27631,N_25019,N_24223);
nor U27632 (N_27632,N_24159,N_25610);
nor U27633 (N_27633,N_25529,N_24705);
nand U27634 (N_27634,N_24247,N_24351);
nand U27635 (N_27635,N_25135,N_24697);
or U27636 (N_27636,N_25963,N_25911);
xor U27637 (N_27637,N_24715,N_24926);
nand U27638 (N_27638,N_25903,N_24814);
nor U27639 (N_27639,N_24284,N_24472);
nor U27640 (N_27640,N_24165,N_25640);
or U27641 (N_27641,N_25228,N_24034);
nor U27642 (N_27642,N_25365,N_24545);
xnor U27643 (N_27643,N_25433,N_25681);
nand U27644 (N_27644,N_25271,N_25108);
or U27645 (N_27645,N_24747,N_25607);
nand U27646 (N_27646,N_24999,N_24543);
or U27647 (N_27647,N_24358,N_25607);
nor U27648 (N_27648,N_25302,N_24443);
nand U27649 (N_27649,N_24486,N_24602);
xnor U27650 (N_27650,N_24510,N_24631);
or U27651 (N_27651,N_25175,N_24549);
nor U27652 (N_27652,N_25702,N_24052);
nand U27653 (N_27653,N_24198,N_25106);
nor U27654 (N_27654,N_25189,N_24985);
xnor U27655 (N_27655,N_25151,N_25670);
xor U27656 (N_27656,N_25338,N_25223);
nand U27657 (N_27657,N_25280,N_24882);
nor U27658 (N_27658,N_25285,N_25819);
and U27659 (N_27659,N_25577,N_25658);
and U27660 (N_27660,N_25678,N_24341);
and U27661 (N_27661,N_25761,N_24978);
xor U27662 (N_27662,N_25648,N_25512);
and U27663 (N_27663,N_24740,N_24690);
or U27664 (N_27664,N_25253,N_24630);
nor U27665 (N_27665,N_24205,N_24145);
xnor U27666 (N_27666,N_25290,N_25497);
nor U27667 (N_27667,N_24596,N_24168);
nand U27668 (N_27668,N_25138,N_25651);
nand U27669 (N_27669,N_25126,N_24954);
or U27670 (N_27670,N_24091,N_24739);
nor U27671 (N_27671,N_24466,N_24010);
and U27672 (N_27672,N_24891,N_25102);
or U27673 (N_27673,N_25766,N_24037);
and U27674 (N_27674,N_24190,N_24382);
xor U27675 (N_27675,N_25296,N_24616);
or U27676 (N_27676,N_24139,N_25372);
and U27677 (N_27677,N_24018,N_24813);
or U27678 (N_27678,N_25117,N_24304);
or U27679 (N_27679,N_24736,N_25720);
or U27680 (N_27680,N_24751,N_25837);
or U27681 (N_27681,N_24456,N_24333);
and U27682 (N_27682,N_24976,N_24764);
xor U27683 (N_27683,N_25485,N_25910);
nand U27684 (N_27684,N_25167,N_24159);
nor U27685 (N_27685,N_24369,N_24487);
or U27686 (N_27686,N_25217,N_25865);
or U27687 (N_27687,N_25289,N_25738);
nand U27688 (N_27688,N_24959,N_25470);
xor U27689 (N_27689,N_24559,N_25490);
nor U27690 (N_27690,N_24446,N_25624);
nand U27691 (N_27691,N_24699,N_25378);
nor U27692 (N_27692,N_24544,N_25296);
or U27693 (N_27693,N_24927,N_24784);
nand U27694 (N_27694,N_25132,N_24294);
or U27695 (N_27695,N_25862,N_25912);
nor U27696 (N_27696,N_24644,N_24625);
or U27697 (N_27697,N_25072,N_24686);
nor U27698 (N_27698,N_25408,N_24361);
nand U27699 (N_27699,N_24881,N_25470);
nor U27700 (N_27700,N_25106,N_25620);
nand U27701 (N_27701,N_25880,N_25246);
and U27702 (N_27702,N_25021,N_24500);
xor U27703 (N_27703,N_24788,N_24139);
nand U27704 (N_27704,N_24857,N_24234);
xnor U27705 (N_27705,N_24046,N_25259);
or U27706 (N_27706,N_24853,N_25443);
xor U27707 (N_27707,N_24890,N_25299);
nand U27708 (N_27708,N_25990,N_24093);
or U27709 (N_27709,N_25415,N_24518);
or U27710 (N_27710,N_25837,N_25578);
nand U27711 (N_27711,N_25752,N_24015);
nand U27712 (N_27712,N_25941,N_24649);
and U27713 (N_27713,N_25544,N_24952);
xnor U27714 (N_27714,N_24663,N_24269);
or U27715 (N_27715,N_25687,N_24283);
or U27716 (N_27716,N_25220,N_24010);
xor U27717 (N_27717,N_24908,N_25612);
and U27718 (N_27718,N_25461,N_24510);
or U27719 (N_27719,N_25259,N_24058);
and U27720 (N_27720,N_25294,N_24212);
nor U27721 (N_27721,N_25858,N_25712);
or U27722 (N_27722,N_24066,N_25275);
and U27723 (N_27723,N_24229,N_25793);
nand U27724 (N_27724,N_24571,N_25951);
and U27725 (N_27725,N_24814,N_24506);
xnor U27726 (N_27726,N_24467,N_25752);
xnor U27727 (N_27727,N_24866,N_24962);
and U27728 (N_27728,N_24151,N_24015);
xor U27729 (N_27729,N_24851,N_24227);
nand U27730 (N_27730,N_24047,N_24599);
nor U27731 (N_27731,N_25388,N_24575);
or U27732 (N_27732,N_25283,N_24321);
nand U27733 (N_27733,N_25196,N_24379);
xor U27734 (N_27734,N_25637,N_24333);
and U27735 (N_27735,N_25057,N_24909);
and U27736 (N_27736,N_25068,N_25833);
and U27737 (N_27737,N_25231,N_24098);
nand U27738 (N_27738,N_25298,N_24158);
and U27739 (N_27739,N_24359,N_25753);
nor U27740 (N_27740,N_25822,N_24307);
nor U27741 (N_27741,N_24090,N_24634);
or U27742 (N_27742,N_24461,N_25611);
and U27743 (N_27743,N_24764,N_24587);
or U27744 (N_27744,N_25269,N_25686);
and U27745 (N_27745,N_24000,N_24950);
nand U27746 (N_27746,N_25757,N_24852);
or U27747 (N_27747,N_24826,N_25721);
and U27748 (N_27748,N_25828,N_24556);
or U27749 (N_27749,N_25862,N_25917);
xnor U27750 (N_27750,N_25439,N_24727);
xnor U27751 (N_27751,N_25817,N_24004);
or U27752 (N_27752,N_24314,N_25100);
and U27753 (N_27753,N_24322,N_25892);
and U27754 (N_27754,N_24358,N_25706);
or U27755 (N_27755,N_25116,N_25829);
and U27756 (N_27756,N_24673,N_25483);
and U27757 (N_27757,N_25633,N_24413);
nand U27758 (N_27758,N_24762,N_25376);
nor U27759 (N_27759,N_24443,N_25016);
nand U27760 (N_27760,N_24413,N_25132);
and U27761 (N_27761,N_25613,N_25341);
and U27762 (N_27762,N_25593,N_25945);
nor U27763 (N_27763,N_24231,N_25970);
xor U27764 (N_27764,N_25747,N_24699);
xnor U27765 (N_27765,N_24724,N_25953);
nor U27766 (N_27766,N_25237,N_25311);
and U27767 (N_27767,N_24289,N_25010);
or U27768 (N_27768,N_25725,N_24640);
nand U27769 (N_27769,N_24499,N_25110);
xnor U27770 (N_27770,N_24715,N_25438);
nand U27771 (N_27771,N_24372,N_24592);
nor U27772 (N_27772,N_24676,N_24219);
nand U27773 (N_27773,N_24315,N_24063);
nor U27774 (N_27774,N_25694,N_25076);
or U27775 (N_27775,N_25602,N_24841);
and U27776 (N_27776,N_25405,N_24329);
nand U27777 (N_27777,N_25239,N_24278);
nor U27778 (N_27778,N_24669,N_24126);
nor U27779 (N_27779,N_24789,N_25814);
nor U27780 (N_27780,N_25711,N_24871);
nand U27781 (N_27781,N_25327,N_25189);
and U27782 (N_27782,N_24148,N_25118);
and U27783 (N_27783,N_25093,N_25533);
nor U27784 (N_27784,N_25246,N_25951);
xnor U27785 (N_27785,N_24843,N_24394);
nor U27786 (N_27786,N_24232,N_25654);
and U27787 (N_27787,N_25369,N_25982);
and U27788 (N_27788,N_24442,N_24471);
xnor U27789 (N_27789,N_25048,N_25089);
nand U27790 (N_27790,N_24331,N_25317);
xor U27791 (N_27791,N_24956,N_24739);
nor U27792 (N_27792,N_24053,N_25105);
and U27793 (N_27793,N_25000,N_24087);
or U27794 (N_27794,N_24367,N_24904);
or U27795 (N_27795,N_24774,N_25686);
nand U27796 (N_27796,N_24909,N_25788);
or U27797 (N_27797,N_25081,N_24618);
or U27798 (N_27798,N_25217,N_24154);
and U27799 (N_27799,N_25671,N_25980);
nor U27800 (N_27800,N_25090,N_24545);
nand U27801 (N_27801,N_24696,N_25889);
xor U27802 (N_27802,N_25155,N_24213);
nor U27803 (N_27803,N_25355,N_25100);
xnor U27804 (N_27804,N_24710,N_24143);
and U27805 (N_27805,N_25817,N_25560);
and U27806 (N_27806,N_25702,N_25715);
xor U27807 (N_27807,N_25197,N_25254);
xnor U27808 (N_27808,N_25501,N_25200);
and U27809 (N_27809,N_24054,N_25438);
xnor U27810 (N_27810,N_25280,N_25291);
xor U27811 (N_27811,N_24319,N_24102);
and U27812 (N_27812,N_25134,N_24602);
and U27813 (N_27813,N_25000,N_24781);
and U27814 (N_27814,N_25992,N_25779);
nor U27815 (N_27815,N_25654,N_24356);
nor U27816 (N_27816,N_25700,N_24616);
or U27817 (N_27817,N_25435,N_25735);
nand U27818 (N_27818,N_25401,N_25193);
nand U27819 (N_27819,N_24215,N_24730);
and U27820 (N_27820,N_25793,N_25877);
nor U27821 (N_27821,N_25205,N_25867);
nand U27822 (N_27822,N_25905,N_25845);
or U27823 (N_27823,N_24862,N_25725);
nand U27824 (N_27824,N_24346,N_24983);
nor U27825 (N_27825,N_25763,N_25401);
or U27826 (N_27826,N_25444,N_25878);
nand U27827 (N_27827,N_24810,N_24538);
or U27828 (N_27828,N_25200,N_24855);
and U27829 (N_27829,N_25295,N_24687);
nand U27830 (N_27830,N_24231,N_25049);
nand U27831 (N_27831,N_24301,N_25124);
xnor U27832 (N_27832,N_24214,N_24606);
nor U27833 (N_27833,N_25847,N_24639);
and U27834 (N_27834,N_24713,N_24878);
nor U27835 (N_27835,N_24943,N_25585);
or U27836 (N_27836,N_25579,N_24651);
and U27837 (N_27837,N_25654,N_24801);
xor U27838 (N_27838,N_25598,N_25943);
or U27839 (N_27839,N_25068,N_24781);
nand U27840 (N_27840,N_25860,N_24203);
and U27841 (N_27841,N_24130,N_24919);
or U27842 (N_27842,N_25977,N_24275);
xnor U27843 (N_27843,N_25181,N_25561);
nand U27844 (N_27844,N_25941,N_25438);
and U27845 (N_27845,N_25291,N_25872);
nor U27846 (N_27846,N_24577,N_25126);
nor U27847 (N_27847,N_25850,N_24988);
nand U27848 (N_27848,N_24309,N_25531);
nor U27849 (N_27849,N_25962,N_25257);
or U27850 (N_27850,N_24230,N_24579);
and U27851 (N_27851,N_25056,N_24551);
nand U27852 (N_27852,N_24786,N_24937);
or U27853 (N_27853,N_24480,N_25358);
xnor U27854 (N_27854,N_24144,N_25387);
nand U27855 (N_27855,N_25995,N_25147);
nand U27856 (N_27856,N_24023,N_24329);
or U27857 (N_27857,N_25898,N_25177);
and U27858 (N_27858,N_24094,N_25276);
xnor U27859 (N_27859,N_25507,N_25348);
or U27860 (N_27860,N_24334,N_24194);
and U27861 (N_27861,N_25749,N_24434);
nand U27862 (N_27862,N_25135,N_25195);
nor U27863 (N_27863,N_24790,N_24361);
xor U27864 (N_27864,N_25767,N_25359);
or U27865 (N_27865,N_24488,N_24196);
and U27866 (N_27866,N_25798,N_24229);
and U27867 (N_27867,N_24893,N_24128);
nand U27868 (N_27868,N_24126,N_24815);
or U27869 (N_27869,N_24868,N_24864);
nor U27870 (N_27870,N_25837,N_24377);
xnor U27871 (N_27871,N_25904,N_24010);
and U27872 (N_27872,N_25339,N_24473);
xor U27873 (N_27873,N_25665,N_25750);
or U27874 (N_27874,N_24960,N_25108);
nand U27875 (N_27875,N_24866,N_25845);
nor U27876 (N_27876,N_24706,N_25236);
nor U27877 (N_27877,N_24770,N_24907);
nand U27878 (N_27878,N_24883,N_24516);
and U27879 (N_27879,N_25599,N_24245);
xor U27880 (N_27880,N_25947,N_24456);
and U27881 (N_27881,N_25545,N_24592);
and U27882 (N_27882,N_24888,N_24172);
xnor U27883 (N_27883,N_24553,N_25315);
nor U27884 (N_27884,N_24376,N_25914);
or U27885 (N_27885,N_24135,N_25012);
or U27886 (N_27886,N_25369,N_25303);
nand U27887 (N_27887,N_24494,N_24198);
and U27888 (N_27888,N_25512,N_25181);
and U27889 (N_27889,N_24032,N_24245);
xnor U27890 (N_27890,N_24202,N_25452);
and U27891 (N_27891,N_25600,N_24657);
nand U27892 (N_27892,N_25149,N_25971);
or U27893 (N_27893,N_25753,N_25442);
and U27894 (N_27894,N_25404,N_24026);
and U27895 (N_27895,N_24023,N_24879);
xor U27896 (N_27896,N_25858,N_24501);
or U27897 (N_27897,N_24454,N_24869);
or U27898 (N_27898,N_24903,N_24121);
nand U27899 (N_27899,N_24129,N_24594);
xor U27900 (N_27900,N_24136,N_24928);
nand U27901 (N_27901,N_25887,N_25414);
xnor U27902 (N_27902,N_25054,N_24804);
nand U27903 (N_27903,N_24262,N_25944);
or U27904 (N_27904,N_25466,N_24049);
nand U27905 (N_27905,N_24898,N_24700);
or U27906 (N_27906,N_25671,N_24878);
or U27907 (N_27907,N_25448,N_25007);
xor U27908 (N_27908,N_24675,N_24824);
nor U27909 (N_27909,N_25750,N_24653);
nand U27910 (N_27910,N_25501,N_25159);
nor U27911 (N_27911,N_25551,N_25073);
nor U27912 (N_27912,N_24373,N_25403);
nor U27913 (N_27913,N_24532,N_24690);
xnor U27914 (N_27914,N_24664,N_24300);
nand U27915 (N_27915,N_25219,N_25641);
and U27916 (N_27916,N_25818,N_25149);
and U27917 (N_27917,N_25639,N_24578);
or U27918 (N_27918,N_25564,N_25207);
or U27919 (N_27919,N_25030,N_24038);
and U27920 (N_27920,N_25062,N_24748);
or U27921 (N_27921,N_24235,N_24706);
nor U27922 (N_27922,N_25445,N_25299);
nor U27923 (N_27923,N_24429,N_25377);
nor U27924 (N_27924,N_24741,N_24339);
and U27925 (N_27925,N_25663,N_24385);
and U27926 (N_27926,N_25734,N_25506);
xor U27927 (N_27927,N_25277,N_25756);
xor U27928 (N_27928,N_24771,N_25554);
xor U27929 (N_27929,N_25406,N_24549);
nor U27930 (N_27930,N_25245,N_25427);
nand U27931 (N_27931,N_24024,N_24971);
and U27932 (N_27932,N_24598,N_25375);
nor U27933 (N_27933,N_24442,N_24394);
xnor U27934 (N_27934,N_25899,N_24041);
or U27935 (N_27935,N_25330,N_25489);
nor U27936 (N_27936,N_25401,N_24736);
xor U27937 (N_27937,N_24601,N_24229);
nand U27938 (N_27938,N_24602,N_25532);
nor U27939 (N_27939,N_24215,N_24345);
xor U27940 (N_27940,N_24777,N_25036);
nand U27941 (N_27941,N_25256,N_25444);
and U27942 (N_27942,N_24628,N_24641);
and U27943 (N_27943,N_24707,N_25715);
xor U27944 (N_27944,N_24605,N_25468);
nand U27945 (N_27945,N_25180,N_25710);
and U27946 (N_27946,N_25494,N_24078);
and U27947 (N_27947,N_24993,N_24033);
nor U27948 (N_27948,N_24849,N_25271);
and U27949 (N_27949,N_24970,N_25681);
nand U27950 (N_27950,N_25387,N_24966);
or U27951 (N_27951,N_25948,N_25537);
and U27952 (N_27952,N_25942,N_25813);
nand U27953 (N_27953,N_24593,N_24439);
xor U27954 (N_27954,N_24777,N_25913);
nor U27955 (N_27955,N_25570,N_24591);
and U27956 (N_27956,N_24637,N_25228);
and U27957 (N_27957,N_24090,N_24103);
xor U27958 (N_27958,N_24733,N_25003);
or U27959 (N_27959,N_24409,N_24976);
nor U27960 (N_27960,N_25630,N_24510);
xor U27961 (N_27961,N_24804,N_24225);
and U27962 (N_27962,N_24336,N_25704);
nand U27963 (N_27963,N_24972,N_24935);
or U27964 (N_27964,N_25955,N_24636);
nand U27965 (N_27965,N_24195,N_25136);
or U27966 (N_27966,N_24286,N_25861);
or U27967 (N_27967,N_25853,N_25935);
xnor U27968 (N_27968,N_25824,N_25084);
or U27969 (N_27969,N_24494,N_25627);
and U27970 (N_27970,N_25302,N_24732);
and U27971 (N_27971,N_25226,N_25957);
nand U27972 (N_27972,N_25001,N_24233);
or U27973 (N_27973,N_24459,N_25123);
nand U27974 (N_27974,N_24814,N_24619);
nor U27975 (N_27975,N_25231,N_24466);
or U27976 (N_27976,N_25075,N_25606);
or U27977 (N_27977,N_24305,N_25629);
xnor U27978 (N_27978,N_25086,N_25812);
nand U27979 (N_27979,N_24893,N_24087);
nor U27980 (N_27980,N_25973,N_24310);
or U27981 (N_27981,N_25501,N_25683);
xor U27982 (N_27982,N_24225,N_25270);
nor U27983 (N_27983,N_25913,N_24176);
and U27984 (N_27984,N_24346,N_25584);
xnor U27985 (N_27985,N_24881,N_24157);
or U27986 (N_27986,N_24692,N_24585);
xor U27987 (N_27987,N_24077,N_24902);
or U27988 (N_27988,N_25180,N_24426);
or U27989 (N_27989,N_24099,N_25420);
and U27990 (N_27990,N_24207,N_25082);
xnor U27991 (N_27991,N_24845,N_24666);
nand U27992 (N_27992,N_25192,N_25739);
and U27993 (N_27993,N_24913,N_25364);
xor U27994 (N_27994,N_24410,N_24676);
xnor U27995 (N_27995,N_25788,N_24619);
nor U27996 (N_27996,N_25180,N_25375);
xnor U27997 (N_27997,N_25747,N_24274);
xor U27998 (N_27998,N_24198,N_24908);
nand U27999 (N_27999,N_24040,N_24621);
or U28000 (N_28000,N_26678,N_26332);
nand U28001 (N_28001,N_27651,N_27600);
xor U28002 (N_28002,N_26037,N_26831);
xnor U28003 (N_28003,N_26185,N_27916);
nand U28004 (N_28004,N_27823,N_26344);
nor U28005 (N_28005,N_27720,N_26505);
and U28006 (N_28006,N_26713,N_26063);
xor U28007 (N_28007,N_26503,N_26543);
nor U28008 (N_28008,N_27398,N_26922);
nand U28009 (N_28009,N_26295,N_27509);
and U28010 (N_28010,N_26180,N_26387);
xor U28011 (N_28011,N_27147,N_26081);
nand U28012 (N_28012,N_26516,N_26253);
and U28013 (N_28013,N_26531,N_27322);
nand U28014 (N_28014,N_27145,N_27879);
nand U28015 (N_28015,N_26703,N_26080);
xnor U28016 (N_28016,N_26007,N_27781);
or U28017 (N_28017,N_27295,N_26345);
nand U28018 (N_28018,N_27779,N_27588);
or U28019 (N_28019,N_27456,N_26143);
xor U28020 (N_28020,N_26411,N_26167);
and U28021 (N_28021,N_27718,N_27457);
xnor U28022 (N_28022,N_26755,N_27925);
xnor U28023 (N_28023,N_27523,N_27783);
nor U28024 (N_28024,N_27043,N_26170);
nand U28025 (N_28025,N_26255,N_27655);
nor U28026 (N_28026,N_26719,N_26905);
xnor U28027 (N_28027,N_26529,N_26680);
or U28028 (N_28028,N_26055,N_27596);
and U28029 (N_28029,N_27510,N_27730);
or U28030 (N_28030,N_27172,N_27199);
or U28031 (N_28031,N_26202,N_26765);
or U28032 (N_28032,N_27135,N_27859);
nand U28033 (N_28033,N_26263,N_26864);
or U28034 (N_28034,N_26616,N_26168);
and U28035 (N_28035,N_27705,N_27118);
or U28036 (N_28036,N_26870,N_26547);
or U28037 (N_28037,N_26245,N_26177);
or U28038 (N_28038,N_26378,N_27763);
or U28039 (N_28039,N_27208,N_27958);
nand U28040 (N_28040,N_26735,N_27694);
nor U28041 (N_28041,N_27015,N_26053);
xor U28042 (N_28042,N_27978,N_27782);
xnor U28043 (N_28043,N_27418,N_26149);
xor U28044 (N_28044,N_26855,N_26268);
or U28045 (N_28045,N_27482,N_27557);
nor U28046 (N_28046,N_26985,N_26305);
nand U28047 (N_28047,N_26954,N_26209);
or U28048 (N_28048,N_27982,N_27613);
and U28049 (N_28049,N_26119,N_26714);
xnor U28050 (N_28050,N_27273,N_27011);
and U28051 (N_28051,N_27333,N_27049);
or U28052 (N_28052,N_26222,N_27461);
or U28053 (N_28053,N_27619,N_26301);
and U28054 (N_28054,N_27403,N_27451);
or U28055 (N_28055,N_26711,N_26339);
nor U28056 (N_28056,N_26402,N_27639);
or U28057 (N_28057,N_27381,N_27211);
xor U28058 (N_28058,N_26468,N_26465);
and U28059 (N_28059,N_26062,N_26051);
nand U28060 (N_28060,N_26901,N_26605);
and U28061 (N_28061,N_27165,N_27669);
and U28062 (N_28062,N_26558,N_26949);
xnor U28063 (N_28063,N_27238,N_26230);
nand U28064 (N_28064,N_26495,N_27814);
and U28065 (N_28065,N_26751,N_27968);
and U28066 (N_28066,N_27559,N_26834);
nor U28067 (N_28067,N_27259,N_27708);
and U28068 (N_28068,N_27649,N_26298);
or U28069 (N_28069,N_27047,N_26815);
nor U28070 (N_28070,N_27385,N_27817);
nor U28071 (N_28071,N_26647,N_26045);
or U28072 (N_28072,N_26115,N_27529);
and U28073 (N_28073,N_27120,N_27098);
xor U28074 (N_28074,N_26451,N_27949);
and U28075 (N_28075,N_27219,N_26218);
and U28076 (N_28076,N_26005,N_27653);
and U28077 (N_28077,N_27525,N_27101);
nand U28078 (N_28078,N_26234,N_27197);
nor U28079 (N_28079,N_26324,N_27928);
or U28080 (N_28080,N_27911,N_27836);
nor U28081 (N_28081,N_26319,N_27663);
nor U28082 (N_28082,N_27164,N_26692);
or U28083 (N_28083,N_26466,N_27533);
nor U28084 (N_28084,N_27325,N_26498);
and U28085 (N_28085,N_26667,N_27526);
and U28086 (N_28086,N_26764,N_27074);
or U28087 (N_28087,N_27413,N_27833);
nand U28088 (N_28088,N_27633,N_27511);
nor U28089 (N_28089,N_26530,N_27059);
nor U28090 (N_28090,N_27391,N_26244);
xor U28091 (N_28091,N_26092,N_26338);
and U28092 (N_28092,N_27767,N_27886);
and U28093 (N_28093,N_27582,N_26663);
nand U28094 (N_28094,N_27981,N_26658);
xnor U28095 (N_28095,N_26969,N_27269);
nand U28096 (N_28096,N_27213,N_27682);
nand U28097 (N_28097,N_27426,N_27931);
and U28098 (N_28098,N_26066,N_26389);
and U28099 (N_28099,N_27980,N_26563);
or U28100 (N_28100,N_27630,N_27173);
nand U28101 (N_28101,N_27412,N_27080);
or U28102 (N_28102,N_26984,N_26668);
nor U28103 (N_28103,N_27277,N_27698);
xor U28104 (N_28104,N_27122,N_26911);
nor U28105 (N_28105,N_27858,N_26512);
or U28106 (N_28106,N_26455,N_26621);
nand U28107 (N_28107,N_27434,N_26448);
nor U28108 (N_28108,N_26026,N_26721);
or U28109 (N_28109,N_27438,N_26067);
nor U28110 (N_28110,N_26031,N_27144);
nor U28111 (N_28111,N_27615,N_26043);
xor U28112 (N_28112,N_26163,N_27969);
xnor U28113 (N_28113,N_27713,N_26135);
nand U28114 (N_28114,N_27466,N_26296);
nor U28115 (N_28115,N_27866,N_26004);
xor U28116 (N_28116,N_26424,N_27857);
or U28117 (N_28117,N_26057,N_27553);
xor U28118 (N_28118,N_27745,N_27967);
or U28119 (N_28119,N_27977,N_27973);
nand U28120 (N_28120,N_27224,N_26259);
or U28121 (N_28121,N_26310,N_26110);
or U28122 (N_28122,N_26827,N_27787);
or U28123 (N_28123,N_26862,N_27174);
or U28124 (N_28124,N_27711,N_27107);
nor U28125 (N_28125,N_27493,N_26164);
and U28126 (N_28126,N_26173,N_27192);
xnor U28127 (N_28127,N_26609,N_26707);
nand U28128 (N_28128,N_27151,N_27139);
or U28129 (N_28129,N_27799,N_26361);
or U28130 (N_28130,N_27266,N_27260);
or U28131 (N_28131,N_26125,N_26229);
xor U28132 (N_28132,N_27640,N_27264);
or U28133 (N_28133,N_27784,N_27441);
nor U28134 (N_28134,N_26029,N_26236);
and U28135 (N_28135,N_27565,N_26737);
xnor U28136 (N_28136,N_27873,N_26859);
and U28137 (N_28137,N_27169,N_26644);
xor U28138 (N_28138,N_27484,N_26606);
and U28139 (N_28139,N_26603,N_26362);
and U28140 (N_28140,N_27296,N_27785);
nand U28141 (N_28141,N_26690,N_26824);
nand U28142 (N_28142,N_26286,N_26847);
nor U28143 (N_28143,N_27156,N_26307);
or U28144 (N_28144,N_27963,N_26910);
xor U28145 (N_28145,N_26844,N_27181);
nand U28146 (N_28146,N_27283,N_26629);
nand U28147 (N_28147,N_26419,N_26175);
and U28148 (N_28148,N_27016,N_27369);
xnor U28149 (N_28149,N_26688,N_26133);
xnor U28150 (N_28150,N_26270,N_26314);
nand U28151 (N_28151,N_26851,N_27222);
nand U28152 (N_28152,N_26211,N_26684);
and U28153 (N_28153,N_27922,N_26715);
xor U28154 (N_28154,N_26706,N_26857);
nand U28155 (N_28155,N_27951,N_27514);
or U28156 (N_28156,N_27474,N_27618);
xor U28157 (N_28157,N_26538,N_27472);
nor U28158 (N_28158,N_26878,N_27756);
nand U28159 (N_28159,N_26243,N_27513);
xor U28160 (N_28160,N_27584,N_26015);
nor U28161 (N_28161,N_26912,N_26687);
nor U28162 (N_28162,N_27303,N_27937);
nand U28163 (N_28163,N_27959,N_26034);
nor U28164 (N_28164,N_26930,N_27987);
xnor U28165 (N_28165,N_27485,N_26179);
nor U28166 (N_28166,N_26630,N_26665);
xnor U28167 (N_28167,N_26582,N_26552);
or U28168 (N_28168,N_26769,N_26872);
nor U28169 (N_28169,N_26291,N_26171);
or U28170 (N_28170,N_27180,N_27644);
nand U28171 (N_28171,N_27078,N_26743);
nand U28172 (N_28172,N_27998,N_27520);
and U28173 (N_28173,N_26739,N_26654);
xnor U28174 (N_28174,N_26427,N_27071);
nor U28175 (N_28175,N_26828,N_27979);
or U28176 (N_28176,N_27008,N_27309);
nand U28177 (N_28177,N_26377,N_27537);
xnor U28178 (N_28178,N_27750,N_27646);
or U28179 (N_28179,N_27668,N_27975);
xor U28180 (N_28180,N_27791,N_27091);
nor U28181 (N_28181,N_26748,N_27910);
or U28182 (N_28182,N_27923,N_26303);
xnor U28183 (N_28183,N_27251,N_26981);
nor U28184 (N_28184,N_26699,N_26601);
xnor U28185 (N_28185,N_26702,N_26823);
xor U28186 (N_28186,N_27683,N_26566);
or U28187 (N_28187,N_27638,N_27244);
or U28188 (N_28188,N_27163,N_26610);
and U28189 (N_28189,N_26726,N_26945);
or U28190 (N_28190,N_27865,N_26458);
xor U28191 (N_28191,N_27862,N_26783);
nand U28192 (N_28192,N_26897,N_26613);
and U28193 (N_28193,N_27941,N_26232);
nor U28194 (N_28194,N_26532,N_27747);
nor U28195 (N_28195,N_27373,N_26623);
nor U28196 (N_28196,N_26800,N_26681);
xor U28197 (N_28197,N_26830,N_27724);
or U28198 (N_28198,N_26423,N_26460);
nor U28199 (N_28199,N_27032,N_27505);
xor U28200 (N_28200,N_27943,N_27818);
nor U28201 (N_28201,N_27530,N_27377);
and U28202 (N_28202,N_27002,N_27214);
xnor U28203 (N_28203,N_27929,N_27367);
or U28204 (N_28204,N_27749,N_27035);
and U28205 (N_28205,N_26006,N_26808);
nor U28206 (N_28206,N_26876,N_26562);
or U28207 (N_28207,N_27193,N_26251);
xor U28208 (N_28208,N_26999,N_27366);
nand U28209 (N_28209,N_26317,N_26861);
xor U28210 (N_28210,N_26651,N_27989);
nand U28211 (N_28211,N_26725,N_26440);
nand U28212 (N_28212,N_27729,N_26369);
or U28213 (N_28213,N_27442,N_27661);
or U28214 (N_28214,N_26090,N_26968);
nand U28215 (N_28215,N_27888,N_27809);
or U28216 (N_28216,N_27946,N_27134);
and U28217 (N_28217,N_26289,N_26777);
xnor U28218 (N_28218,N_26429,N_27189);
xnor U28219 (N_28219,N_27587,N_26256);
nand U28220 (N_28220,N_27486,N_26447);
nor U28221 (N_28221,N_27837,N_27306);
nor U28222 (N_28222,N_27878,N_26269);
nor U28223 (N_28223,N_27938,N_26148);
and U28224 (N_28224,N_26089,N_26024);
or U28225 (N_28225,N_27345,N_26453);
nor U28226 (N_28226,N_27893,N_26152);
xnor U28227 (N_28227,N_26557,N_27632);
nor U28228 (N_28228,N_26759,N_27890);
or U28229 (N_28229,N_27437,N_27499);
nand U28230 (N_28230,N_27714,N_27570);
xnor U28231 (N_28231,N_27021,N_26600);
nand U28232 (N_28232,N_26250,N_26249);
xor U28233 (N_28233,N_26354,N_26444);
xor U28234 (N_28234,N_26524,N_26528);
and U28235 (N_28235,N_26576,N_26271);
nand U28236 (N_28236,N_27722,N_27246);
xor U28237 (N_28237,N_26627,N_27731);
nor U28238 (N_28238,N_27754,N_26716);
or U28239 (N_28239,N_26084,N_27849);
and U28240 (N_28240,N_27620,N_27334);
nor U28241 (N_28241,N_27871,N_26730);
nor U28242 (N_28242,N_26551,N_27906);
nand U28243 (N_28243,N_26363,N_26138);
or U28244 (N_28244,N_27512,N_27532);
xnor U28245 (N_28245,N_27734,N_27789);
xnor U28246 (N_28246,N_26340,N_26883);
and U28247 (N_28247,N_26020,N_26504);
or U28248 (N_28248,N_26477,N_27354);
or U28249 (N_28249,N_26103,N_26052);
and U28250 (N_28250,N_27292,N_26449);
nor U28251 (N_28251,N_27023,N_27517);
xnor U28252 (N_28252,N_27908,N_27067);
and U28253 (N_28253,N_26578,N_27397);
xor U28254 (N_28254,N_27489,N_26106);
xnor U28255 (N_28255,N_27880,N_26909);
xor U28256 (N_28256,N_26308,N_27490);
nor U28257 (N_28257,N_26728,N_27019);
or U28258 (N_28258,N_27313,N_26276);
nor U28259 (N_28259,N_27820,N_27498);
and U28260 (N_28260,N_27964,N_27786);
and U28261 (N_28261,N_27117,N_26881);
and U28262 (N_28262,N_27432,N_26100);
nor U28263 (N_28263,N_26000,N_26306);
nand U28264 (N_28264,N_27691,N_26195);
or U28265 (N_28265,N_27488,N_27300);
nor U28266 (N_28266,N_26920,N_27220);
nand U28267 (N_28267,N_27227,N_27875);
and U28268 (N_28268,N_26464,N_27966);
nor U28269 (N_28269,N_27436,N_27579);
nor U28270 (N_28270,N_27700,N_26235);
and U28271 (N_28271,N_26720,N_27390);
and U28272 (N_28272,N_26144,N_27518);
and U28273 (N_28273,N_26858,N_26973);
and U28274 (N_28274,N_26254,N_27723);
and U28275 (N_28275,N_26572,N_27703);
nor U28276 (N_28276,N_27806,N_26718);
nand U28277 (N_28277,N_27188,N_27918);
nor U28278 (N_28278,N_26522,N_27123);
xor U28279 (N_28279,N_26813,N_26372);
and U28280 (N_28280,N_26391,N_27136);
xnor U28281 (N_28281,N_27664,N_27113);
nand U28282 (N_28282,N_26581,N_27311);
nand U28283 (N_28283,N_26659,N_27468);
nand U28284 (N_28284,N_26047,N_26604);
or U28285 (N_28285,N_26262,N_27473);
or U28286 (N_28286,N_27109,N_27674);
and U28287 (N_28287,N_26187,N_26113);
xnor U28288 (N_28288,N_26096,N_27522);
or U28289 (N_28289,N_27801,N_26775);
or U28290 (N_28290,N_27932,N_27738);
xnor U28291 (N_28291,N_27770,N_27055);
nand U28292 (N_28292,N_27119,N_26788);
and U28293 (N_28293,N_27326,N_26575);
nand U28294 (N_28294,N_27344,N_26257);
xnor U28295 (N_28295,N_27240,N_26484);
or U28296 (N_28296,N_27036,N_26746);
and U28297 (N_28297,N_27231,N_26943);
nand U28298 (N_28298,N_27414,N_27765);
or U28299 (N_28299,N_27996,N_26799);
nor U28300 (N_28300,N_26889,N_27900);
xor U28301 (N_28301,N_26722,N_27678);
and U28302 (N_28302,N_26884,N_26474);
nor U28303 (N_28303,N_27527,N_27005);
xnor U28304 (N_28304,N_26842,N_27312);
xnor U28305 (N_28305,N_26513,N_26997);
nand U28306 (N_28306,N_26381,N_27131);
and U28307 (N_28307,N_26365,N_26592);
and U28308 (N_28308,N_26131,N_26717);
nor U28309 (N_28309,N_27406,N_26986);
xnor U28310 (N_28310,N_27508,N_26083);
and U28311 (N_28311,N_27874,N_27891);
xor U28312 (N_28312,N_26673,N_26213);
xor U28313 (N_28313,N_27764,N_27534);
nor U28314 (N_28314,N_27631,N_26614);
nand U28315 (N_28315,N_27606,N_26095);
nor U28316 (N_28316,N_27610,N_27170);
and U28317 (N_28317,N_27324,N_26591);
nand U28318 (N_28318,N_26698,N_27501);
nor U28319 (N_28319,N_26098,N_26560);
nor U28320 (N_28320,N_26502,N_26403);
and U28321 (N_28321,N_26742,N_27245);
and U28322 (N_28322,N_26450,N_26932);
nand U28323 (N_28323,N_26277,N_26261);
nor U28324 (N_28324,N_26147,N_26645);
or U28325 (N_28325,N_26960,N_26107);
and U28326 (N_28326,N_27168,N_27680);
xor U28327 (N_28327,N_27093,N_26380);
xor U28328 (N_28328,N_27645,N_27575);
nand U28329 (N_28329,N_27357,N_26805);
xor U28330 (N_28330,N_26485,N_26198);
nor U28331 (N_28331,N_27672,N_27449);
or U28332 (N_28332,N_27991,N_26472);
nor U28333 (N_28333,N_26669,N_27717);
xnor U28334 (N_28334,N_26955,N_26639);
nand U28335 (N_28335,N_26506,N_26046);
and U28336 (N_28336,N_27476,N_26763);
nand U28337 (N_28337,N_27177,N_26040);
nand U28338 (N_28338,N_26486,N_27298);
nor U28339 (N_28339,N_26567,N_26890);
nor U28340 (N_28340,N_27129,N_26297);
or U28341 (N_28341,N_27628,N_26944);
and U28342 (N_28342,N_27415,N_26694);
xor U28343 (N_28343,N_27375,N_26819);
or U28344 (N_28344,N_27018,N_26077);
nor U28345 (N_28345,N_27346,N_26546);
nand U28346 (N_28346,N_27627,N_27810);
and U28347 (N_28347,N_26772,N_26208);
and U28348 (N_28348,N_26685,N_27234);
or U28349 (N_28349,N_27323,N_27206);
nand U28350 (N_28350,N_26446,N_27743);
xnor U28351 (N_28351,N_27315,N_26555);
nand U28352 (N_28352,N_27241,N_26935);
xnor U28353 (N_28353,N_27110,N_26991);
xor U28354 (N_28354,N_27318,N_26456);
nor U28355 (N_28355,N_27429,N_27634);
xor U28356 (N_28356,N_27001,N_26686);
and U28357 (N_28357,N_26795,N_26892);
xnor U28358 (N_28358,N_26632,N_26416);
nand U28359 (N_28359,N_26846,N_26134);
and U28360 (N_28360,N_26525,N_27033);
nand U28361 (N_28361,N_27228,N_27250);
nor U28362 (N_28362,N_27453,N_26771);
xor U28363 (N_28363,N_27393,N_26165);
nand U28364 (N_28364,N_26508,N_26619);
xnor U28365 (N_28365,N_27540,N_27732);
and U28366 (N_28366,N_27190,N_27812);
nand U28367 (N_28367,N_27569,N_26696);
and U28368 (N_28368,N_26641,N_26540);
or U28369 (N_28369,N_27072,N_26397);
nor U28370 (N_28370,N_26215,N_27611);
and U28371 (N_28371,N_26197,N_26267);
and U28372 (N_28372,N_27469,N_26784);
nor U28373 (N_28373,N_27726,N_27636);
or U28374 (N_28374,N_26848,N_27503);
and U28375 (N_28375,N_26583,N_27902);
xnor U28376 (N_28376,N_27057,N_27758);
or U28377 (N_28377,N_27604,N_27341);
xor U28378 (N_28378,N_26754,N_26181);
or U28379 (N_28379,N_27811,N_27106);
and U28380 (N_28380,N_27045,N_27370);
nand U28381 (N_28381,N_26597,N_26059);
and U28382 (N_28382,N_27807,N_26833);
or U28383 (N_28383,N_27230,N_26050);
nand U28384 (N_28384,N_26526,N_27590);
nand U28385 (N_28385,N_27621,N_26829);
or U28386 (N_28386,N_26792,N_27007);
and U28387 (N_28387,N_26587,N_26602);
or U28388 (N_28388,N_27643,N_26894);
nand U28389 (N_28389,N_26396,N_26488);
or U28390 (N_28390,N_27719,N_26626);
nor U28391 (N_28391,N_27304,N_27601);
nand U28392 (N_28392,N_26490,N_26517);
nor U28393 (N_28393,N_27563,N_26060);
nand U28394 (N_28394,N_26018,N_26571);
and U28395 (N_28395,N_27372,N_27470);
nand U28396 (N_28396,N_27562,N_26278);
or U28397 (N_28397,N_26118,N_27755);
or U28398 (N_28398,N_27384,N_27710);
nand U28399 (N_28399,N_27157,N_26708);
nand U28400 (N_28400,N_26414,N_27020);
xor U28401 (N_28401,N_26153,N_27641);
and U28402 (N_28402,N_26430,N_26733);
and U28403 (N_28403,N_27475,N_26022);
nand U28404 (N_28404,N_26782,N_27210);
nand U28405 (N_28405,N_27970,N_27550);
xnor U28406 (N_28406,N_26674,N_26607);
nor U28407 (N_28407,N_27751,N_26412);
and U28408 (N_28408,N_26166,N_27592);
and U28409 (N_28409,N_27395,N_26789);
nand U28410 (N_28410,N_26642,N_27409);
nor U28411 (N_28411,N_27838,N_26976);
nor U28412 (N_28412,N_26328,N_26766);
xnor U28413 (N_28413,N_27077,N_27159);
nor U28414 (N_28414,N_26643,N_26589);
and U28415 (N_28415,N_26839,N_27102);
nor U28416 (N_28416,N_26407,N_26330);
xnor U28417 (N_28417,N_27348,N_27338);
xnor U28418 (N_28418,N_27774,N_27930);
nand U28419 (N_28419,N_26977,N_27660);
xnor U28420 (N_28420,N_27506,N_26902);
nand U28421 (N_28421,N_26679,N_27567);
nor U28422 (N_28422,N_27160,N_26071);
nor U28423 (N_28423,N_27362,N_27116);
xor U28424 (N_28424,N_27221,N_27564);
or U28425 (N_28425,N_26279,N_26938);
or U28426 (N_28426,N_27154,N_26671);
and U28427 (N_28427,N_26554,N_26142);
or U28428 (N_28428,N_26882,N_27337);
nand U28429 (N_28429,N_26288,N_27648);
xnor U28430 (N_28430,N_26041,N_27307);
nor U28431 (N_28431,N_26482,N_27748);
and U28432 (N_28432,N_26732,N_26770);
nor U28433 (N_28433,N_27196,N_27115);
or U28434 (N_28434,N_26539,N_26079);
nor U28435 (N_28435,N_27819,N_26467);
nor U28436 (N_28436,N_27647,N_27363);
nand U28437 (N_28437,N_27642,N_26193);
and U28438 (N_28438,N_27542,N_26996);
or U28439 (N_28439,N_27446,N_27531);
or U28440 (N_28440,N_27343,N_26404);
nand U28441 (N_28441,N_27138,N_26825);
or U28442 (N_28442,N_27090,N_26368);
nor U28443 (N_28443,N_27450,N_27876);
nand U28444 (N_28444,N_26917,N_27848);
nand U28445 (N_28445,N_27458,N_27697);
nor U28446 (N_28446,N_26201,N_27046);
xnor U28447 (N_28447,N_26023,N_26329);
and U28448 (N_28448,N_27671,N_26661);
nand U28449 (N_28449,N_27762,N_27447);
nor U28450 (N_28450,N_26373,N_27133);
and U28451 (N_28451,N_26660,N_26952);
xnor U28452 (N_28452,N_26014,N_26085);
and U28453 (N_28453,N_27773,N_26974);
nor U28454 (N_28454,N_26127,N_26240);
nand U28455 (N_28455,N_26394,N_26272);
and U28456 (N_28456,N_27608,N_26479);
and U28457 (N_28457,N_26433,N_26662);
nand U28458 (N_28458,N_26545,N_27798);
and U28459 (N_28459,N_26936,N_26599);
or U28460 (N_28460,N_26704,N_26896);
nor U28461 (N_28461,N_27321,N_27044);
or U28462 (N_28462,N_27287,N_26027);
xnor U28463 (N_28463,N_27268,N_26491);
or U28464 (N_28464,N_26379,N_26638);
and U28465 (N_28465,N_26341,N_26035);
nand U28466 (N_28466,N_27757,N_26835);
nor U28467 (N_28467,N_27431,N_27371);
and U28468 (N_28468,N_26961,N_27805);
nand U28469 (N_28469,N_27920,N_26388);
nand U28470 (N_28470,N_27616,N_27685);
xor U28471 (N_28471,N_27374,N_26248);
and U28472 (N_28472,N_27439,N_27712);
nand U28473 (N_28473,N_26044,N_26094);
nand U28474 (N_28474,N_26183,N_27659);
or U28475 (N_28475,N_26664,N_27428);
or U28476 (N_28476,N_27594,N_27576);
or U28477 (N_28477,N_27285,N_26360);
nand U28478 (N_28478,N_27884,N_27141);
and U28479 (N_28479,N_27423,N_27267);
or U28480 (N_28480,N_27793,N_27356);
nand U28481 (N_28481,N_26871,N_26785);
nor U28482 (N_28482,N_26773,N_27885);
and U28483 (N_28483,N_26536,N_27654);
nor U28484 (N_28484,N_27062,N_27185);
nand U28485 (N_28485,N_26797,N_26112);
or U28486 (N_28486,N_27280,N_27797);
or U28487 (N_28487,N_27637,N_27612);
and U28488 (N_28488,N_27706,N_26435);
or U28489 (N_28489,N_26778,N_26806);
or U28490 (N_28490,N_27972,N_27294);
and U28491 (N_28491,N_26192,N_27097);
or U28492 (N_28492,N_26975,N_26425);
xor U28493 (N_28493,N_27042,N_27974);
nand U28494 (N_28494,N_27236,N_26205);
nand U28495 (N_28495,N_27625,N_27463);
nor U28496 (N_28496,N_26573,N_27950);
and U28497 (N_28497,N_26224,N_26203);
and U28498 (N_28498,N_27105,N_26242);
or U28499 (N_28499,N_27607,N_27521);
or U28500 (N_28500,N_26724,N_26832);
nor U28501 (N_28501,N_27253,N_27417);
nor U28502 (N_28502,N_26321,N_27194);
nor U28503 (N_28503,N_27389,N_26499);
and U28504 (N_28504,N_27962,N_27912);
nor U28505 (N_28505,N_26786,N_26246);
and U28506 (N_28506,N_27889,N_27657);
xor U28507 (N_28507,N_27317,N_26155);
and U28508 (N_28508,N_26320,N_27670);
xnor U28509 (N_28509,N_26492,N_27877);
and U28510 (N_28510,N_26074,N_27556);
nor U28511 (N_28511,N_26212,N_26970);
xor U28512 (N_28512,N_26082,N_27815);
or U28513 (N_28513,N_26494,N_27985);
or U28514 (N_28514,N_27332,N_26712);
nand U28515 (N_28515,N_26877,N_26648);
or U28516 (N_28516,N_27954,N_26102);
and U28517 (N_28517,N_26518,N_26916);
nand U28518 (N_28518,N_27022,N_26011);
or U28519 (N_28519,N_26925,N_26519);
nand U28520 (N_28520,N_26221,N_26367);
or U28521 (N_28521,N_26334,N_27027);
or U28522 (N_28522,N_27919,N_26867);
or U28523 (N_28523,N_26570,N_27394);
nand U28524 (N_28524,N_27383,N_27212);
nand U28525 (N_28525,N_27014,N_26762);
xnor U28526 (N_28526,N_26845,N_27087);
nand U28527 (N_28527,N_26010,N_26946);
nor U28528 (N_28528,N_27103,N_26461);
or U28529 (N_28529,N_27955,N_27408);
and U28530 (N_28530,N_26086,N_27382);
nand U28531 (N_28531,N_27041,N_26070);
or U28532 (N_28532,N_27207,N_27746);
nand U28533 (N_28533,N_26906,N_26252);
and U28534 (N_28534,N_26207,N_27840);
nor U28535 (N_28535,N_27624,N_26853);
and U28536 (N_28536,N_26331,N_27992);
nor U28537 (N_28537,N_26875,N_27861);
and U28538 (N_28538,N_27166,N_27709);
nor U28539 (N_28539,N_27085,N_27860);
nor U28540 (N_28540,N_26352,N_26182);
nor U28541 (N_28541,N_26199,N_27626);
nor U28542 (N_28542,N_27715,N_27265);
xor U28543 (N_28543,N_27839,N_26942);
xor U28544 (N_28544,N_26312,N_27242);
xnor U28545 (N_28545,N_26415,N_26544);
nor U28546 (N_28546,N_27548,N_26967);
xor U28547 (N_28547,N_26200,N_26284);
nand U28548 (N_28548,N_27560,N_27328);
and U28549 (N_28549,N_27504,N_27095);
xnor U28550 (N_28550,N_27350,N_26959);
xnor U28551 (N_28551,N_26441,N_27320);
nor U28552 (N_28552,N_27351,N_26913);
xor U28553 (N_28553,N_27017,N_27617);
nand U28554 (N_28554,N_26965,N_26233);
nor U28555 (N_28555,N_26617,N_27687);
xnor U28556 (N_28556,N_27150,N_26439);
or U28557 (N_28557,N_26075,N_27702);
nand U28558 (N_28558,N_27716,N_27945);
nand U28559 (N_28559,N_26983,N_26395);
or U28560 (N_28560,N_26452,N_26431);
or U28561 (N_28561,N_27997,N_27552);
xor U28562 (N_28562,N_27030,N_26126);
or U28563 (N_28563,N_27605,N_27430);
nand U28564 (N_28564,N_26178,N_26744);
and U28565 (N_28565,N_26016,N_26756);
nor U28566 (N_28566,N_26781,N_26814);
xor U28567 (N_28567,N_26426,N_26141);
nand U28568 (N_28568,N_27898,N_27686);
xor U28569 (N_28569,N_27577,N_27176);
nor U28570 (N_28570,N_26693,N_26438);
nor U28571 (N_28571,N_27824,N_27183);
or U28572 (N_28572,N_26879,N_27155);
and U28573 (N_28573,N_27195,N_27462);
and U28574 (N_28574,N_27401,N_27247);
or U28575 (N_28575,N_27175,N_27761);
xor U28576 (N_28576,N_27235,N_26812);
nor U28577 (N_28577,N_27060,N_27330);
nand U28578 (N_28578,N_26520,N_27004);
xnor U28579 (N_28579,N_26817,N_26039);
nand U28580 (N_28580,N_26042,N_27727);
or U28581 (N_28581,N_26553,N_27068);
nor U28582 (N_28582,N_26370,N_26646);
nor U28583 (N_28583,N_27850,N_27127);
or U28584 (N_28584,N_27288,N_27179);
xor U28585 (N_28585,N_27209,N_27578);
nand U28586 (N_28586,N_27178,N_27379);
and U28587 (N_28587,N_27561,N_27843);
xnor U28588 (N_28588,N_26120,N_27065);
nor U28589 (N_28589,N_26934,N_26527);
and U28590 (N_28590,N_26316,N_26358);
nor U28591 (N_28591,N_27961,N_27031);
nand U28592 (N_28592,N_26802,N_26574);
and U28593 (N_28593,N_26768,N_27305);
xnor U28594 (N_28594,N_26962,N_27201);
and U28595 (N_28595,N_26371,N_26666);
or U28596 (N_28596,N_26150,N_27006);
xor U28597 (N_28597,N_27999,N_27662);
xor U28598 (N_28598,N_27844,N_26705);
or U28599 (N_28599,N_27842,N_27314);
nor U28600 (N_28600,N_27777,N_27568);
xnor U28601 (N_28601,N_26926,N_26710);
nand U28602 (N_28602,N_27854,N_27360);
and U28603 (N_28603,N_27289,N_26376);
nand U28604 (N_28604,N_27753,N_26869);
or U28605 (N_28605,N_27086,N_26542);
nand U28606 (N_28606,N_27826,N_27003);
or U28607 (N_28607,N_26758,N_26309);
nand U28608 (N_28608,N_26921,N_27400);
nor U28609 (N_28609,N_27566,N_26325);
or U28610 (N_28610,N_27465,N_26357);
or U28611 (N_28611,N_27831,N_26028);
nor U28612 (N_28612,N_27800,N_26470);
nor U28613 (N_28613,N_27009,N_27760);
or U28614 (N_28614,N_26670,N_27897);
nand U28615 (N_28615,N_27739,N_27342);
nor U28616 (N_28616,N_26631,N_26323);
or U28617 (N_28617,N_27913,N_27056);
nor U28618 (N_28618,N_26128,N_27775);
nand U28619 (N_28619,N_27507,N_26584);
or U28620 (N_28620,N_26480,N_27881);
xnor U28621 (N_28621,N_26580,N_26787);
xnor U28622 (N_28622,N_27496,N_26366);
xnor U28623 (N_28623,N_26108,N_27191);
nor U28624 (N_28624,N_27444,N_27420);
nor U28625 (N_28625,N_27203,N_26950);
nand U28626 (N_28626,N_26342,N_27917);
or U28627 (N_28627,N_27721,N_27993);
nor U28628 (N_28628,N_26675,N_27125);
nand U28629 (N_28629,N_27692,N_27158);
and U28630 (N_28630,N_26217,N_26683);
nand U28631 (N_28631,N_26393,N_27899);
and U28632 (N_28632,N_26349,N_26608);
nand U28633 (N_28633,N_26176,N_27574);
or U28634 (N_28634,N_27491,N_27232);
nand U28635 (N_28635,N_27539,N_26753);
or U28636 (N_28636,N_26327,N_27699);
nand U28637 (N_28637,N_27778,N_26117);
or U28638 (N_28638,N_27696,N_26682);
xnor U28639 (N_28639,N_27171,N_26548);
nor U28640 (N_28640,N_27558,N_27075);
xnor U28641 (N_28641,N_27088,N_27602);
xnor U28642 (N_28642,N_26247,N_27132);
and U28643 (N_28643,N_26826,N_27316);
nor U28644 (N_28644,N_27029,N_26953);
nor U28645 (N_28645,N_26190,N_27108);
nand U28646 (N_28646,N_26750,N_27467);
nand U28647 (N_28647,N_27053,N_26072);
nand U28648 (N_28648,N_27237,N_27376);
nor U28649 (N_28649,N_26514,N_27573);
nor U28650 (N_28650,N_27121,N_26907);
nand U28651 (N_28651,N_26337,N_27882);
nor U28652 (N_28652,N_27656,N_26137);
nor U28653 (N_28653,N_26392,N_27635);
xnor U28654 (N_28654,N_26091,N_26417);
xor U28655 (N_28655,N_27957,N_26274);
and U28656 (N_28656,N_26442,N_26030);
xnor U28657 (N_28657,N_26489,N_27847);
nand U28658 (N_28658,N_27863,N_26130);
nor U28659 (N_28659,N_26865,N_27276);
and U28660 (N_28660,N_26933,N_27544);
or U28661 (N_28661,N_27519,N_27435);
xor U28662 (N_28662,N_27089,N_26987);
nor U28663 (N_28663,N_27026,N_26174);
xor U28664 (N_28664,N_26677,N_27076);
nor U28665 (N_28665,N_26818,N_27248);
nor U28666 (N_28666,N_27492,N_27301);
nor U28667 (N_28667,N_26012,N_27652);
xnor U28668 (N_28668,N_26752,N_26887);
and U28669 (N_28669,N_26734,N_26428);
and U28670 (N_28670,N_27771,N_26569);
or U28671 (N_28671,N_27433,N_26634);
or U28672 (N_28672,N_27701,N_27976);
nand U28673 (N_28673,N_26918,N_27827);
nand U28674 (N_28674,N_27541,N_26798);
nor U28675 (N_28675,N_27153,N_26109);
nor U28676 (N_28676,N_27140,N_26238);
xnor U28677 (N_28677,N_27229,N_26124);
or U28678 (N_28678,N_27909,N_26219);
or U28679 (N_28679,N_27039,N_27665);
and U28680 (N_28680,N_26281,N_27443);
nor U28681 (N_28681,N_26672,N_27609);
or U28682 (N_28682,N_27984,N_26088);
nand U28683 (N_28683,N_26635,N_27856);
and U28684 (N_28684,N_26204,N_27361);
xor U28685 (N_28685,N_26947,N_27549);
xor U28686 (N_28686,N_27124,N_26564);
nor U28687 (N_28687,N_27104,N_27830);
xor U28688 (N_28688,N_27994,N_27892);
nand U28689 (N_28689,N_26836,N_27939);
xor U28690 (N_28690,N_27184,N_27995);
and U28691 (N_28691,N_26880,N_26535);
xor U28692 (N_28692,N_26405,N_26333);
or U28693 (N_28693,N_27258,N_26924);
nor U28694 (N_28694,N_27494,N_26409);
and U28695 (N_28695,N_27907,N_27853);
or U28696 (N_28696,N_26579,N_27536);
or U28697 (N_28697,N_26343,N_27790);
and U28698 (N_28698,N_26293,N_27516);
or U28699 (N_28699,N_27069,N_27404);
nor U28700 (N_28700,N_27364,N_26136);
and U28701 (N_28701,N_26701,N_26791);
nand U28702 (N_28702,N_26434,N_27742);
nor U28703 (N_28703,N_26061,N_27940);
nand U28704 (N_28704,N_27262,N_26069);
nand U28705 (N_28705,N_26145,N_27058);
or U28706 (N_28706,N_27825,N_26656);
or U28707 (N_28707,N_26355,N_26033);
and U28708 (N_28708,N_26577,N_27872);
and U28709 (N_28709,N_26228,N_27223);
xor U28710 (N_28710,N_27673,N_27788);
or U28711 (N_28711,N_26994,N_26140);
nor U28712 (N_28712,N_26723,N_27261);
nor U28713 (N_28713,N_26928,N_27971);
or U28714 (N_28714,N_27688,N_26898);
xnor U28715 (N_28715,N_26459,N_27274);
and U28716 (N_28716,N_27137,N_27319);
nand U28717 (N_28717,N_26893,N_26497);
or U28718 (N_28718,N_27835,N_27841);
or U28719 (N_28719,N_27883,N_26649);
nand U28720 (N_28720,N_27308,N_27419);
nor U28721 (N_28721,N_26958,N_27162);
or U28722 (N_28722,N_26172,N_27048);
nand U28723 (N_28723,N_26266,N_26473);
nand U28724 (N_28724,N_27769,N_26927);
or U28725 (N_28725,N_27452,N_27063);
nand U28726 (N_28726,N_26691,N_27421);
xor U28727 (N_28727,N_27339,N_27864);
or U28728 (N_28728,N_27792,N_26432);
or U28729 (N_28729,N_26809,N_27927);
nor U28730 (N_28730,N_27816,N_26873);
xnor U28731 (N_28731,N_27598,N_26534);
nand U28732 (N_28732,N_26908,N_26793);
or U28733 (N_28733,N_26191,N_26158);
xor U28734 (N_28734,N_27965,N_26837);
and U28735 (N_28735,N_27388,N_27064);
or U28736 (N_28736,N_27744,N_26038);
or U28737 (N_28737,N_27780,N_26273);
or U28738 (N_28738,N_26633,N_26929);
xnor U28739 (N_28739,N_27684,N_26874);
or U28740 (N_28740,N_27852,N_27832);
xor U28741 (N_28741,N_26840,N_27622);
nor U28742 (N_28742,N_27112,N_26820);
nand U28743 (N_28743,N_26227,N_26496);
and U28744 (N_28744,N_26017,N_27477);
nand U28745 (N_28745,N_27082,N_26931);
or U28746 (N_28746,N_26500,N_26287);
nor U28747 (N_28747,N_27281,N_26129);
nor U28748 (N_28748,N_26483,N_26625);
or U28749 (N_28749,N_27143,N_27290);
and U28750 (N_28750,N_27681,N_27733);
nor U28751 (N_28751,N_26383,N_26628);
and U28752 (N_28752,N_26462,N_26336);
nand U28753 (N_28753,N_27256,N_26585);
xor U28754 (N_28754,N_27040,N_26511);
or U28755 (N_28755,N_26533,N_27677);
xnor U28756 (N_28756,N_26283,N_27546);
xnor U28757 (N_28757,N_26774,N_27358);
nor U28758 (N_28758,N_26891,N_26541);
nand U28759 (N_28759,N_26993,N_26139);
xnor U28760 (N_28760,N_26008,N_26550);
nor U28761 (N_28761,N_26019,N_27768);
nand U28762 (N_28762,N_27182,N_27502);
xnor U28763 (N_28763,N_27051,N_27936);
and U28764 (N_28764,N_27218,N_27983);
or U28765 (N_28765,N_26549,N_27952);
and U28766 (N_28766,N_26990,N_26410);
nor U28767 (N_28767,N_27052,N_26225);
or U28768 (N_28768,N_27380,N_27901);
nand U28769 (N_28769,N_26655,N_26794);
or U28770 (N_28770,N_26804,N_26979);
or U28771 (N_28771,N_26471,N_27921);
or U28772 (N_28772,N_26637,N_27411);
nand U28773 (N_28773,N_26001,N_26111);
xnor U28774 (N_28774,N_27025,N_27948);
nor U28775 (N_28775,N_26940,N_27595);
xor U28776 (N_28776,N_26709,N_26400);
nor U28777 (N_28777,N_27695,N_27944);
and U28778 (N_28778,N_26700,N_26156);
nor U28779 (N_28779,N_26390,N_26241);
nor U28780 (N_28780,N_27740,N_27034);
or U28781 (N_28781,N_27092,N_26054);
or U28782 (N_28782,N_27986,N_26009);
nand U28783 (N_28783,N_27368,N_26013);
nand U28784 (N_28784,N_27378,N_27365);
xnor U28785 (N_28785,N_26184,N_27934);
xor U28786 (N_28786,N_27667,N_27215);
nand U28787 (N_28787,N_26956,N_27693);
or U28788 (N_28788,N_27591,N_27953);
nor U28789 (N_28789,N_27904,N_27083);
nand U28790 (N_28790,N_27243,N_27679);
xnor U28791 (N_28791,N_26104,N_26151);
and U28792 (N_28792,N_27355,N_26767);
nor U28793 (N_28793,N_27821,N_27073);
nand U28794 (N_28794,N_26903,N_27416);
nor U28795 (N_28795,N_27279,N_27352);
or U28796 (N_28796,N_26398,N_27855);
nor U28797 (N_28797,N_27422,N_26860);
nand U28798 (N_28798,N_27736,N_27867);
nor U28799 (N_28799,N_26885,N_27658);
nor U28800 (N_28800,N_26058,N_27725);
xnor U28801 (N_28801,N_26588,N_27942);
nor U28802 (N_28802,N_26807,N_26521);
nor U28803 (N_28803,N_26971,N_27445);
xnor U28804 (N_28804,N_26957,N_27571);
nand U28805 (N_28805,N_27500,N_27198);
xor U28806 (N_28806,N_26188,N_26078);
and U28807 (N_28807,N_26988,N_26622);
nand U28808 (N_28808,N_27407,N_27424);
nand U28809 (N_28809,N_27741,N_26816);
nand U28810 (N_28810,N_27000,N_27599);
xnor U28811 (N_28811,N_26729,N_26385);
or U28812 (N_28812,N_26123,N_26507);
nor U28813 (N_28813,N_27405,N_26036);
and U28814 (N_28814,N_27528,N_27666);
xnor U28815 (N_28815,N_26594,N_26736);
or U28816 (N_28816,N_26258,N_26568);
nand U28817 (N_28817,N_27111,N_27894);
or U28818 (N_28818,N_27096,N_26413);
xnor U28819 (N_28819,N_26821,N_27152);
or U28820 (N_28820,N_26326,N_27593);
xor U28821 (N_28821,N_26652,N_26657);
xnor U28822 (N_28822,N_26863,N_27795);
nand U28823 (N_28823,N_27167,N_27543);
and U28824 (N_28824,N_27161,N_27956);
nand U28825 (N_28825,N_26995,N_26226);
and U28826 (N_28826,N_27336,N_26206);
or U28827 (N_28827,N_27297,N_27263);
nor U28828 (N_28828,N_26856,N_26843);
nor U28829 (N_28829,N_27099,N_27728);
nand U28830 (N_28830,N_27028,N_26747);
xor U28831 (N_28831,N_27455,N_27829);
and U28832 (N_28832,N_26116,N_26294);
nor U28833 (N_28833,N_26868,N_27478);
or U28834 (N_28834,N_27597,N_26351);
or U28835 (N_28835,N_26593,N_26966);
or U28836 (N_28836,N_26941,N_26169);
nor U28837 (N_28837,N_27349,N_26216);
xor U28838 (N_28838,N_26194,N_26478);
nand U28839 (N_28839,N_27440,N_26849);
and U28840 (N_28840,N_27255,N_27257);
or U28841 (N_28841,N_27623,N_27310);
xnor U28842 (N_28842,N_27822,N_27583);
or U28843 (N_28843,N_26741,N_27226);
xnor U28844 (N_28844,N_27903,N_27960);
nor U28845 (N_28845,N_27538,N_27284);
xnor U28846 (N_28846,N_27216,N_26159);
nand U28847 (N_28847,N_27200,N_26220);
and U28848 (N_28848,N_26101,N_27870);
nand U28849 (N_28849,N_27481,N_26160);
nor U28850 (N_28850,N_27286,N_27128);
nor U28851 (N_28851,N_27586,N_27387);
nor U28852 (N_28852,N_26146,N_26523);
xnor U28853 (N_28853,N_27094,N_26676);
xor U28854 (N_28854,N_26304,N_26032);
nand U28855 (N_28855,N_26114,N_26299);
nand U28856 (N_28856,N_27487,N_26811);
xor U28857 (N_28857,N_26105,N_27803);
nand U28858 (N_28858,N_27233,N_27402);
and U28859 (N_28859,N_26065,N_27130);
nand U28860 (N_28860,N_26049,N_26923);
xor U28861 (N_28861,N_26021,N_26260);
nand U28862 (N_28862,N_26346,N_26420);
nand U28863 (N_28863,N_26122,N_26445);
and U28864 (N_28864,N_26375,N_26421);
or U28865 (N_28865,N_27515,N_26056);
or U28866 (N_28866,N_27580,N_27225);
and U28867 (N_28867,N_26239,N_26761);
nor U28868 (N_28868,N_26650,N_26841);
or U28869 (N_28869,N_27249,N_27545);
or U28870 (N_28870,N_26313,N_26437);
nand U28871 (N_28871,N_27834,N_27100);
and U28872 (N_28872,N_27079,N_27675);
nor U28873 (N_28873,N_26939,N_27802);
xor U28874 (N_28874,N_27359,N_27480);
or U28875 (N_28875,N_27868,N_26980);
xnor U28876 (N_28876,N_27146,N_26196);
xnor U28877 (N_28877,N_26886,N_26586);
nand U28878 (N_28878,N_26537,N_26854);
or U28879 (N_28879,N_27759,N_27081);
or U28880 (N_28880,N_26469,N_26282);
nor U28881 (N_28881,N_27869,N_26399);
and U28882 (N_28882,N_26322,N_27589);
and U28883 (N_28883,N_26275,N_27572);
nor U28884 (N_28884,N_27585,N_26210);
or U28885 (N_28885,N_26093,N_26481);
nand U28886 (N_28886,N_26302,N_26852);
nor U28887 (N_28887,N_26561,N_26989);
and U28888 (N_28888,N_26796,N_27013);
and U28889 (N_28889,N_26418,N_27766);
nor U28890 (N_28890,N_27126,N_26596);
and U28891 (N_28891,N_26915,N_26822);
and U28892 (N_28892,N_26475,N_27347);
and U28893 (N_28893,N_27614,N_27396);
and U28894 (N_28894,N_26476,N_27935);
nand U28895 (N_28895,N_27796,N_27933);
nand U28896 (N_28896,N_26695,N_27581);
and U28897 (N_28897,N_27340,N_26097);
or U28898 (N_28898,N_27271,N_26801);
nand U28899 (N_28899,N_27535,N_27554);
xnor U28900 (N_28900,N_26382,N_26214);
nor U28901 (N_28901,N_27037,N_26285);
nand U28902 (N_28902,N_27555,N_26760);
and U28903 (N_28903,N_26048,N_27142);
xnor U28904 (N_28904,N_26998,N_27813);
nand U28905 (N_28905,N_26335,N_26068);
or U28906 (N_28906,N_27186,N_26866);
xor U28907 (N_28907,N_26776,N_27293);
xnor U28908 (N_28908,N_27914,N_26265);
nand U28909 (N_28909,N_27254,N_26731);
or U28910 (N_28910,N_26838,N_27291);
or U28911 (N_28911,N_27704,N_27460);
xor U28912 (N_28912,N_26121,N_26501);
nand U28913 (N_28913,N_26757,N_26727);
xnor U28914 (N_28914,N_27329,N_26073);
and U28915 (N_28915,N_27114,N_27202);
nand U28916 (N_28916,N_26914,N_27464);
xor U28917 (N_28917,N_26132,N_27547);
and U28918 (N_28918,N_26359,N_26348);
nand U28919 (N_28919,N_26161,N_26002);
and U28920 (N_28920,N_27690,N_26895);
or U28921 (N_28921,N_26992,N_27425);
xor U28922 (N_28922,N_27828,N_27676);
nor U28923 (N_28923,N_27905,N_26436);
or U28924 (N_28924,N_26408,N_27915);
or U28925 (N_28925,N_27808,N_26850);
and U28926 (N_28926,N_27399,N_27689);
nor U28927 (N_28927,N_27988,N_27302);
nand U28928 (N_28928,N_26590,N_27148);
xor U28929 (N_28929,N_27335,N_27752);
nand U28930 (N_28930,N_26919,N_27272);
and U28931 (N_28931,N_26487,N_26595);
and U28932 (N_28932,N_26888,N_27524);
nand U28933 (N_28933,N_26689,N_26780);
nand U28934 (N_28934,N_27050,N_27024);
or U28935 (N_28935,N_26972,N_27275);
nor U28936 (N_28936,N_26099,N_26948);
xor U28937 (N_28937,N_26899,N_27495);
nor U28938 (N_28938,N_26900,N_26978);
nor U28939 (N_28939,N_27331,N_26937);
and U28940 (N_28940,N_27707,N_27204);
nor U28941 (N_28941,N_26612,N_27038);
nor U28942 (N_28942,N_27926,N_26463);
nand U28943 (N_28943,N_27895,N_26509);
nand U28944 (N_28944,N_27010,N_26223);
nor U28945 (N_28945,N_27427,N_26280);
nand U28946 (N_28946,N_26315,N_26640);
xor U28947 (N_28947,N_27737,N_26738);
nand U28948 (N_28948,N_26951,N_26749);
or U28949 (N_28949,N_26598,N_26064);
or U28950 (N_28950,N_27217,N_26624);
nor U28951 (N_28951,N_27804,N_27084);
or U28952 (N_28952,N_27845,N_27924);
nand U28953 (N_28953,N_27012,N_26350);
xor U28954 (N_28954,N_27794,N_26300);
xor U28955 (N_28955,N_27887,N_26803);
or U28956 (N_28956,N_26318,N_27282);
and U28957 (N_28957,N_27410,N_27629);
or U28958 (N_28958,N_26615,N_26515);
and U28959 (N_28959,N_26636,N_27386);
and U28960 (N_28960,N_27205,N_27776);
and U28961 (N_28961,N_26157,N_26565);
xnor U28962 (N_28962,N_26290,N_27851);
xor U28963 (N_28963,N_26154,N_27846);
nor U28964 (N_28964,N_26162,N_26003);
nand U28965 (N_28965,N_26264,N_27353);
or U28966 (N_28966,N_26443,N_27187);
nand U28967 (N_28967,N_27149,N_27947);
xor U28968 (N_28968,N_27066,N_26790);
xnor U28969 (N_28969,N_26779,N_26457);
or U28970 (N_28970,N_26364,N_27990);
xnor U28971 (N_28971,N_26454,N_27070);
nor U28972 (N_28972,N_26189,N_26556);
nor U28973 (N_28973,N_27327,N_26374);
nor U28974 (N_28974,N_26618,N_27896);
and U28975 (N_28975,N_27061,N_26697);
xnor U28976 (N_28976,N_26401,N_26087);
or U28977 (N_28977,N_26231,N_27650);
and U28978 (N_28978,N_26964,N_27054);
and U28979 (N_28979,N_27454,N_27551);
xor U28980 (N_28980,N_27239,N_26292);
and U28981 (N_28981,N_26510,N_27603);
and U28982 (N_28982,N_26237,N_27483);
or U28983 (N_28983,N_27270,N_26406);
nand U28984 (N_28984,N_26653,N_27252);
or U28985 (N_28985,N_26353,N_26810);
or U28986 (N_28986,N_26559,N_27479);
or U28987 (N_28987,N_26620,N_26186);
xor U28988 (N_28988,N_26386,N_27278);
nand U28989 (N_28989,N_26740,N_26422);
and U28990 (N_28990,N_26025,N_26982);
nor U28991 (N_28991,N_26347,N_27459);
or U28992 (N_28992,N_27772,N_26611);
or U28993 (N_28993,N_27735,N_26745);
xor U28994 (N_28994,N_26904,N_26384);
or U28995 (N_28995,N_26963,N_26356);
nor U28996 (N_28996,N_27448,N_27497);
and U28997 (N_28997,N_27299,N_27392);
nor U28998 (N_28998,N_26493,N_26076);
and U28999 (N_28999,N_26311,N_27471);
xnor U29000 (N_29000,N_26531,N_27812);
nand U29001 (N_29001,N_27148,N_27098);
xnor U29002 (N_29002,N_27668,N_27462);
and U29003 (N_29003,N_26160,N_27387);
and U29004 (N_29004,N_26164,N_27416);
or U29005 (N_29005,N_26153,N_27136);
or U29006 (N_29006,N_26493,N_27110);
nand U29007 (N_29007,N_27388,N_27408);
and U29008 (N_29008,N_27731,N_26552);
and U29009 (N_29009,N_27751,N_26427);
or U29010 (N_29010,N_27226,N_26954);
nor U29011 (N_29011,N_27104,N_26433);
nor U29012 (N_29012,N_26394,N_26161);
xnor U29013 (N_29013,N_27802,N_27983);
nor U29014 (N_29014,N_26973,N_27060);
nor U29015 (N_29015,N_27471,N_26383);
and U29016 (N_29016,N_27350,N_26472);
or U29017 (N_29017,N_26090,N_27324);
or U29018 (N_29018,N_27685,N_27484);
nor U29019 (N_29019,N_27631,N_26782);
xnor U29020 (N_29020,N_27219,N_27432);
nand U29021 (N_29021,N_27880,N_26441);
and U29022 (N_29022,N_27468,N_27799);
and U29023 (N_29023,N_26574,N_27562);
nor U29024 (N_29024,N_27330,N_27471);
nand U29025 (N_29025,N_27938,N_26337);
or U29026 (N_29026,N_26548,N_27776);
nand U29027 (N_29027,N_27914,N_26543);
and U29028 (N_29028,N_27611,N_27761);
nor U29029 (N_29029,N_26899,N_27501);
and U29030 (N_29030,N_26546,N_26397);
nand U29031 (N_29031,N_27172,N_26374);
and U29032 (N_29032,N_27971,N_26656);
xor U29033 (N_29033,N_26347,N_26285);
nor U29034 (N_29034,N_26747,N_26356);
nor U29035 (N_29035,N_27047,N_27650);
xor U29036 (N_29036,N_27604,N_26004);
nand U29037 (N_29037,N_26888,N_27636);
or U29038 (N_29038,N_26457,N_26721);
and U29039 (N_29039,N_26852,N_27524);
and U29040 (N_29040,N_26361,N_27503);
or U29041 (N_29041,N_27049,N_27504);
and U29042 (N_29042,N_26490,N_26200);
xnor U29043 (N_29043,N_27963,N_27074);
xnor U29044 (N_29044,N_27534,N_27931);
nand U29045 (N_29045,N_27360,N_26927);
xnor U29046 (N_29046,N_26761,N_26656);
or U29047 (N_29047,N_26519,N_26255);
or U29048 (N_29048,N_27059,N_26464);
nand U29049 (N_29049,N_27424,N_27509);
nor U29050 (N_29050,N_27576,N_27143);
nand U29051 (N_29051,N_27415,N_27586);
nor U29052 (N_29052,N_27855,N_27194);
or U29053 (N_29053,N_26000,N_26107);
nand U29054 (N_29054,N_26171,N_27703);
nor U29055 (N_29055,N_26458,N_26567);
and U29056 (N_29056,N_26622,N_27219);
nand U29057 (N_29057,N_26132,N_27522);
and U29058 (N_29058,N_26613,N_27409);
and U29059 (N_29059,N_26048,N_27167);
nand U29060 (N_29060,N_26894,N_27245);
or U29061 (N_29061,N_27432,N_26048);
nand U29062 (N_29062,N_27160,N_27297);
or U29063 (N_29063,N_26595,N_27315);
or U29064 (N_29064,N_27757,N_27972);
and U29065 (N_29065,N_26995,N_27888);
nand U29066 (N_29066,N_26747,N_26101);
nor U29067 (N_29067,N_26368,N_27834);
or U29068 (N_29068,N_27135,N_26753);
nand U29069 (N_29069,N_27518,N_26564);
nor U29070 (N_29070,N_27661,N_27963);
nand U29071 (N_29071,N_26797,N_27728);
or U29072 (N_29072,N_27787,N_27089);
xor U29073 (N_29073,N_26899,N_26549);
nand U29074 (N_29074,N_27343,N_26914);
nor U29075 (N_29075,N_26739,N_26908);
nor U29076 (N_29076,N_27545,N_26700);
or U29077 (N_29077,N_27529,N_26586);
or U29078 (N_29078,N_26147,N_26685);
nor U29079 (N_29079,N_26379,N_27514);
nor U29080 (N_29080,N_27288,N_27377);
and U29081 (N_29081,N_27345,N_27280);
nand U29082 (N_29082,N_26083,N_26524);
nor U29083 (N_29083,N_27519,N_27612);
nand U29084 (N_29084,N_27043,N_26977);
nor U29085 (N_29085,N_26968,N_27756);
xnor U29086 (N_29086,N_27977,N_27416);
nand U29087 (N_29087,N_26238,N_26893);
nand U29088 (N_29088,N_26849,N_27698);
and U29089 (N_29089,N_27848,N_26706);
nand U29090 (N_29090,N_26285,N_26716);
nor U29091 (N_29091,N_26552,N_27366);
nor U29092 (N_29092,N_26151,N_26608);
nor U29093 (N_29093,N_27717,N_27293);
nand U29094 (N_29094,N_27034,N_27607);
xnor U29095 (N_29095,N_27457,N_26086);
and U29096 (N_29096,N_27944,N_27826);
or U29097 (N_29097,N_26178,N_27480);
nand U29098 (N_29098,N_26961,N_26997);
xnor U29099 (N_29099,N_26392,N_26182);
or U29100 (N_29100,N_27121,N_26575);
nor U29101 (N_29101,N_26112,N_26628);
and U29102 (N_29102,N_27449,N_27660);
nand U29103 (N_29103,N_27975,N_27662);
nor U29104 (N_29104,N_27219,N_26337);
nand U29105 (N_29105,N_27061,N_26247);
or U29106 (N_29106,N_27085,N_26863);
nand U29107 (N_29107,N_27444,N_27308);
xor U29108 (N_29108,N_26255,N_27508);
xnor U29109 (N_29109,N_27997,N_27653);
xor U29110 (N_29110,N_27069,N_27241);
and U29111 (N_29111,N_26034,N_26221);
or U29112 (N_29112,N_27599,N_27636);
nand U29113 (N_29113,N_27319,N_27375);
xor U29114 (N_29114,N_27386,N_27887);
nand U29115 (N_29115,N_27164,N_27957);
xnor U29116 (N_29116,N_27709,N_27041);
or U29117 (N_29117,N_26524,N_26298);
nand U29118 (N_29118,N_26276,N_27037);
nor U29119 (N_29119,N_27708,N_26827);
and U29120 (N_29120,N_26120,N_26165);
nor U29121 (N_29121,N_26075,N_27486);
nor U29122 (N_29122,N_26856,N_26446);
nand U29123 (N_29123,N_27920,N_26604);
or U29124 (N_29124,N_27466,N_26510);
or U29125 (N_29125,N_26976,N_26326);
xnor U29126 (N_29126,N_26787,N_26264);
nor U29127 (N_29127,N_27564,N_27825);
nand U29128 (N_29128,N_26023,N_27255);
or U29129 (N_29129,N_26616,N_27744);
nor U29130 (N_29130,N_27989,N_26244);
xnor U29131 (N_29131,N_26133,N_26852);
nor U29132 (N_29132,N_26129,N_27765);
and U29133 (N_29133,N_26956,N_26167);
or U29134 (N_29134,N_27096,N_27288);
and U29135 (N_29135,N_27822,N_27923);
and U29136 (N_29136,N_27622,N_26941);
nor U29137 (N_29137,N_27125,N_26383);
and U29138 (N_29138,N_27868,N_26668);
or U29139 (N_29139,N_27206,N_26613);
xor U29140 (N_29140,N_26839,N_27756);
nor U29141 (N_29141,N_26090,N_27048);
nor U29142 (N_29142,N_27557,N_26118);
or U29143 (N_29143,N_27853,N_26914);
nand U29144 (N_29144,N_26871,N_26217);
and U29145 (N_29145,N_27481,N_26512);
nor U29146 (N_29146,N_27771,N_27048);
xor U29147 (N_29147,N_27476,N_26522);
xor U29148 (N_29148,N_27070,N_26188);
nand U29149 (N_29149,N_26861,N_27317);
nor U29150 (N_29150,N_27656,N_26745);
nand U29151 (N_29151,N_27306,N_27712);
and U29152 (N_29152,N_27369,N_26097);
xnor U29153 (N_29153,N_26653,N_26190);
or U29154 (N_29154,N_26005,N_27562);
nand U29155 (N_29155,N_27626,N_27152);
xnor U29156 (N_29156,N_27525,N_27365);
nand U29157 (N_29157,N_26617,N_27531);
nor U29158 (N_29158,N_27023,N_26906);
or U29159 (N_29159,N_27888,N_27760);
xnor U29160 (N_29160,N_26472,N_26161);
or U29161 (N_29161,N_26896,N_26181);
nor U29162 (N_29162,N_26343,N_26470);
or U29163 (N_29163,N_27206,N_27525);
and U29164 (N_29164,N_27232,N_26031);
and U29165 (N_29165,N_26506,N_27264);
nand U29166 (N_29166,N_26451,N_26802);
and U29167 (N_29167,N_26136,N_26993);
xnor U29168 (N_29168,N_26317,N_26656);
or U29169 (N_29169,N_27063,N_26479);
and U29170 (N_29170,N_26536,N_26726);
xor U29171 (N_29171,N_26388,N_26506);
nand U29172 (N_29172,N_27873,N_27056);
nand U29173 (N_29173,N_27970,N_26180);
nand U29174 (N_29174,N_27285,N_26820);
or U29175 (N_29175,N_26707,N_27333);
or U29176 (N_29176,N_26103,N_27300);
and U29177 (N_29177,N_26068,N_27446);
nor U29178 (N_29178,N_26955,N_26329);
or U29179 (N_29179,N_26274,N_26898);
or U29180 (N_29180,N_26984,N_27917);
or U29181 (N_29181,N_26002,N_26054);
and U29182 (N_29182,N_26819,N_27071);
xor U29183 (N_29183,N_27283,N_27688);
or U29184 (N_29184,N_27806,N_26684);
and U29185 (N_29185,N_26440,N_26711);
xor U29186 (N_29186,N_26878,N_27293);
and U29187 (N_29187,N_27044,N_26441);
nand U29188 (N_29188,N_26807,N_26829);
nor U29189 (N_29189,N_26127,N_26308);
nor U29190 (N_29190,N_26402,N_26880);
nor U29191 (N_29191,N_26550,N_27278);
nor U29192 (N_29192,N_27297,N_26815);
or U29193 (N_29193,N_27406,N_27682);
nor U29194 (N_29194,N_26980,N_26240);
xor U29195 (N_29195,N_26233,N_27426);
xnor U29196 (N_29196,N_27684,N_26590);
and U29197 (N_29197,N_26403,N_27474);
xnor U29198 (N_29198,N_27770,N_27687);
xor U29199 (N_29199,N_26161,N_27852);
and U29200 (N_29200,N_27145,N_26147);
and U29201 (N_29201,N_27838,N_27379);
and U29202 (N_29202,N_26775,N_26672);
nand U29203 (N_29203,N_27813,N_26947);
and U29204 (N_29204,N_27258,N_27034);
or U29205 (N_29205,N_27401,N_26034);
nor U29206 (N_29206,N_26222,N_27418);
and U29207 (N_29207,N_27536,N_27742);
or U29208 (N_29208,N_26153,N_26844);
xnor U29209 (N_29209,N_27386,N_27216);
nand U29210 (N_29210,N_26334,N_26758);
nand U29211 (N_29211,N_27050,N_26765);
xor U29212 (N_29212,N_27760,N_26046);
xor U29213 (N_29213,N_26598,N_26437);
and U29214 (N_29214,N_27819,N_26539);
or U29215 (N_29215,N_27883,N_27799);
xor U29216 (N_29216,N_26472,N_27741);
or U29217 (N_29217,N_27347,N_27435);
xor U29218 (N_29218,N_27178,N_27906);
or U29219 (N_29219,N_27783,N_27124);
or U29220 (N_29220,N_27455,N_27581);
nor U29221 (N_29221,N_26207,N_27291);
and U29222 (N_29222,N_27258,N_27399);
xor U29223 (N_29223,N_26818,N_27097);
or U29224 (N_29224,N_26447,N_27396);
nor U29225 (N_29225,N_27380,N_27374);
xnor U29226 (N_29226,N_27817,N_26659);
xor U29227 (N_29227,N_26335,N_26336);
or U29228 (N_29228,N_26571,N_27939);
nor U29229 (N_29229,N_27400,N_26003);
or U29230 (N_29230,N_26850,N_27813);
xor U29231 (N_29231,N_27516,N_26468);
xor U29232 (N_29232,N_26013,N_27871);
or U29233 (N_29233,N_26595,N_26818);
nor U29234 (N_29234,N_26427,N_27380);
and U29235 (N_29235,N_27963,N_26053);
or U29236 (N_29236,N_26073,N_26479);
nand U29237 (N_29237,N_27810,N_26222);
and U29238 (N_29238,N_27082,N_27803);
nor U29239 (N_29239,N_26675,N_26509);
or U29240 (N_29240,N_26791,N_27569);
and U29241 (N_29241,N_27468,N_27280);
and U29242 (N_29242,N_26791,N_27594);
or U29243 (N_29243,N_27718,N_26389);
or U29244 (N_29244,N_27085,N_27190);
and U29245 (N_29245,N_26526,N_26344);
nand U29246 (N_29246,N_27224,N_26396);
and U29247 (N_29247,N_26308,N_26674);
nand U29248 (N_29248,N_27732,N_27185);
nor U29249 (N_29249,N_27457,N_27331);
nand U29250 (N_29250,N_26216,N_27776);
and U29251 (N_29251,N_27387,N_26838);
nand U29252 (N_29252,N_26058,N_27311);
and U29253 (N_29253,N_27879,N_26601);
and U29254 (N_29254,N_27136,N_27250);
or U29255 (N_29255,N_27031,N_26496);
xor U29256 (N_29256,N_27797,N_26514);
nand U29257 (N_29257,N_27638,N_26722);
and U29258 (N_29258,N_27413,N_26225);
nor U29259 (N_29259,N_26898,N_27037);
xnor U29260 (N_29260,N_27660,N_26801);
and U29261 (N_29261,N_26647,N_27357);
or U29262 (N_29262,N_27039,N_26737);
or U29263 (N_29263,N_27994,N_26298);
xnor U29264 (N_29264,N_27022,N_26270);
nand U29265 (N_29265,N_26135,N_26607);
xnor U29266 (N_29266,N_26150,N_27236);
xnor U29267 (N_29267,N_26429,N_26397);
nand U29268 (N_29268,N_27614,N_26290);
and U29269 (N_29269,N_27392,N_26451);
nor U29270 (N_29270,N_27276,N_26281);
and U29271 (N_29271,N_26831,N_27202);
and U29272 (N_29272,N_27232,N_27794);
xnor U29273 (N_29273,N_27690,N_27421);
nor U29274 (N_29274,N_26413,N_27815);
nand U29275 (N_29275,N_27437,N_27298);
nor U29276 (N_29276,N_26641,N_27695);
or U29277 (N_29277,N_27830,N_26864);
nor U29278 (N_29278,N_27507,N_26019);
xnor U29279 (N_29279,N_26572,N_27714);
xnor U29280 (N_29280,N_27040,N_26935);
nand U29281 (N_29281,N_27592,N_27893);
nor U29282 (N_29282,N_27855,N_27050);
xor U29283 (N_29283,N_26108,N_26980);
nand U29284 (N_29284,N_26489,N_27262);
and U29285 (N_29285,N_27340,N_27842);
and U29286 (N_29286,N_27236,N_27887);
and U29287 (N_29287,N_26700,N_26382);
or U29288 (N_29288,N_27887,N_26469);
and U29289 (N_29289,N_26760,N_26813);
nand U29290 (N_29290,N_27678,N_26125);
nand U29291 (N_29291,N_27703,N_27974);
and U29292 (N_29292,N_26796,N_26221);
and U29293 (N_29293,N_27220,N_26017);
or U29294 (N_29294,N_27105,N_26561);
nand U29295 (N_29295,N_27146,N_27567);
or U29296 (N_29296,N_26026,N_27150);
or U29297 (N_29297,N_26255,N_26463);
nor U29298 (N_29298,N_26012,N_27163);
nor U29299 (N_29299,N_26322,N_27685);
nor U29300 (N_29300,N_27749,N_27513);
or U29301 (N_29301,N_27176,N_26880);
nand U29302 (N_29302,N_26748,N_26813);
xnor U29303 (N_29303,N_26255,N_27605);
nand U29304 (N_29304,N_26967,N_26868);
or U29305 (N_29305,N_26271,N_26315);
nand U29306 (N_29306,N_27974,N_27060);
nand U29307 (N_29307,N_27601,N_26852);
xor U29308 (N_29308,N_27913,N_27373);
or U29309 (N_29309,N_26603,N_26899);
or U29310 (N_29310,N_26173,N_26360);
or U29311 (N_29311,N_27063,N_27793);
nor U29312 (N_29312,N_26498,N_26080);
or U29313 (N_29313,N_26207,N_27242);
nand U29314 (N_29314,N_26044,N_26518);
or U29315 (N_29315,N_27524,N_26197);
nor U29316 (N_29316,N_27790,N_27985);
or U29317 (N_29317,N_27587,N_26375);
xnor U29318 (N_29318,N_27914,N_27980);
xor U29319 (N_29319,N_26486,N_27341);
xor U29320 (N_29320,N_26213,N_26846);
xnor U29321 (N_29321,N_26491,N_27888);
and U29322 (N_29322,N_27881,N_27795);
nor U29323 (N_29323,N_27472,N_26169);
or U29324 (N_29324,N_26317,N_27511);
or U29325 (N_29325,N_26809,N_26581);
xnor U29326 (N_29326,N_27792,N_26492);
and U29327 (N_29327,N_26625,N_27461);
and U29328 (N_29328,N_27965,N_27426);
nor U29329 (N_29329,N_27731,N_26621);
and U29330 (N_29330,N_26364,N_26225);
nand U29331 (N_29331,N_26579,N_27679);
and U29332 (N_29332,N_27480,N_26899);
or U29333 (N_29333,N_27937,N_26598);
or U29334 (N_29334,N_26882,N_27650);
nand U29335 (N_29335,N_26496,N_27257);
nor U29336 (N_29336,N_26832,N_26069);
or U29337 (N_29337,N_26173,N_27397);
nor U29338 (N_29338,N_26611,N_27338);
or U29339 (N_29339,N_27089,N_27800);
nor U29340 (N_29340,N_26903,N_27105);
nand U29341 (N_29341,N_26240,N_27100);
xnor U29342 (N_29342,N_26991,N_26450);
or U29343 (N_29343,N_26329,N_27688);
or U29344 (N_29344,N_27725,N_27638);
nand U29345 (N_29345,N_26955,N_27981);
nor U29346 (N_29346,N_26691,N_27949);
or U29347 (N_29347,N_27357,N_26579);
nor U29348 (N_29348,N_27124,N_26245);
and U29349 (N_29349,N_27268,N_27570);
or U29350 (N_29350,N_26353,N_27495);
nor U29351 (N_29351,N_27739,N_27359);
nor U29352 (N_29352,N_26576,N_27037);
xnor U29353 (N_29353,N_27313,N_26285);
nor U29354 (N_29354,N_26991,N_27664);
and U29355 (N_29355,N_27368,N_27347);
xor U29356 (N_29356,N_27274,N_27245);
nor U29357 (N_29357,N_27537,N_27250);
nor U29358 (N_29358,N_27991,N_26969);
and U29359 (N_29359,N_27928,N_26594);
xor U29360 (N_29360,N_26341,N_26966);
or U29361 (N_29361,N_26169,N_26142);
nand U29362 (N_29362,N_26301,N_27576);
nor U29363 (N_29363,N_26071,N_26099);
nor U29364 (N_29364,N_26149,N_26620);
nand U29365 (N_29365,N_27237,N_27141);
nand U29366 (N_29366,N_26376,N_26875);
xnor U29367 (N_29367,N_26971,N_26664);
xnor U29368 (N_29368,N_26660,N_27180);
and U29369 (N_29369,N_26717,N_27555);
nand U29370 (N_29370,N_27947,N_26015);
nand U29371 (N_29371,N_26137,N_26175);
or U29372 (N_29372,N_27187,N_26576);
xnor U29373 (N_29373,N_26707,N_27078);
xnor U29374 (N_29374,N_27900,N_27038);
nand U29375 (N_29375,N_26886,N_26003);
and U29376 (N_29376,N_27133,N_26600);
nor U29377 (N_29377,N_27063,N_26993);
and U29378 (N_29378,N_26023,N_26362);
nand U29379 (N_29379,N_27251,N_27417);
xnor U29380 (N_29380,N_26291,N_26562);
nand U29381 (N_29381,N_26591,N_27303);
nand U29382 (N_29382,N_27457,N_27669);
or U29383 (N_29383,N_26639,N_26656);
nand U29384 (N_29384,N_27980,N_27739);
xnor U29385 (N_29385,N_27453,N_27192);
xor U29386 (N_29386,N_26701,N_27762);
nand U29387 (N_29387,N_26571,N_27119);
and U29388 (N_29388,N_27008,N_26780);
nor U29389 (N_29389,N_27795,N_26331);
and U29390 (N_29390,N_26395,N_26132);
nor U29391 (N_29391,N_26276,N_27463);
nor U29392 (N_29392,N_27743,N_26069);
and U29393 (N_29393,N_27730,N_27974);
and U29394 (N_29394,N_27604,N_27448);
nand U29395 (N_29395,N_26374,N_26524);
xnor U29396 (N_29396,N_26464,N_27689);
nand U29397 (N_29397,N_26145,N_26811);
nor U29398 (N_29398,N_26761,N_27244);
xnor U29399 (N_29399,N_27716,N_27503);
nand U29400 (N_29400,N_26990,N_27188);
xor U29401 (N_29401,N_26692,N_26227);
nand U29402 (N_29402,N_27017,N_27442);
nor U29403 (N_29403,N_26894,N_26602);
and U29404 (N_29404,N_27778,N_26983);
nor U29405 (N_29405,N_26112,N_27681);
nor U29406 (N_29406,N_26553,N_27592);
or U29407 (N_29407,N_27899,N_27870);
and U29408 (N_29408,N_27939,N_26277);
and U29409 (N_29409,N_26603,N_27755);
and U29410 (N_29410,N_26904,N_26419);
nor U29411 (N_29411,N_26131,N_27020);
nor U29412 (N_29412,N_26160,N_26344);
or U29413 (N_29413,N_26423,N_27849);
nor U29414 (N_29414,N_26091,N_26403);
nand U29415 (N_29415,N_27406,N_26926);
and U29416 (N_29416,N_26164,N_27186);
nand U29417 (N_29417,N_26385,N_26101);
or U29418 (N_29418,N_26426,N_26758);
or U29419 (N_29419,N_26926,N_26618);
nand U29420 (N_29420,N_26698,N_27016);
and U29421 (N_29421,N_26648,N_26687);
nand U29422 (N_29422,N_27544,N_27558);
nand U29423 (N_29423,N_27790,N_27984);
or U29424 (N_29424,N_26120,N_27045);
or U29425 (N_29425,N_26489,N_26797);
nor U29426 (N_29426,N_27056,N_26126);
nor U29427 (N_29427,N_26587,N_26579);
nor U29428 (N_29428,N_26216,N_26499);
or U29429 (N_29429,N_26936,N_26844);
nand U29430 (N_29430,N_26738,N_27119);
or U29431 (N_29431,N_27502,N_26331);
or U29432 (N_29432,N_26681,N_27059);
xnor U29433 (N_29433,N_27066,N_27367);
nor U29434 (N_29434,N_26316,N_27654);
xnor U29435 (N_29435,N_27620,N_27850);
xor U29436 (N_29436,N_27908,N_27964);
xnor U29437 (N_29437,N_26782,N_26081);
xnor U29438 (N_29438,N_26009,N_26702);
xnor U29439 (N_29439,N_26759,N_26469);
or U29440 (N_29440,N_26313,N_26574);
and U29441 (N_29441,N_27413,N_27263);
nor U29442 (N_29442,N_27291,N_27337);
or U29443 (N_29443,N_27277,N_26347);
nor U29444 (N_29444,N_26062,N_26444);
or U29445 (N_29445,N_26075,N_27343);
or U29446 (N_29446,N_26169,N_26693);
or U29447 (N_29447,N_26967,N_26490);
or U29448 (N_29448,N_27433,N_26826);
nor U29449 (N_29449,N_26102,N_26741);
nand U29450 (N_29450,N_26052,N_26469);
nand U29451 (N_29451,N_27559,N_26639);
or U29452 (N_29452,N_27637,N_27226);
xor U29453 (N_29453,N_26260,N_26745);
nor U29454 (N_29454,N_27988,N_27881);
and U29455 (N_29455,N_27690,N_26745);
xor U29456 (N_29456,N_27724,N_27815);
xnor U29457 (N_29457,N_26690,N_27240);
nor U29458 (N_29458,N_26548,N_27325);
nand U29459 (N_29459,N_27229,N_27038);
xor U29460 (N_29460,N_27311,N_27368);
nor U29461 (N_29461,N_27930,N_27308);
nand U29462 (N_29462,N_27768,N_27887);
xnor U29463 (N_29463,N_27886,N_26363);
xor U29464 (N_29464,N_26382,N_26776);
xor U29465 (N_29465,N_26539,N_27078);
and U29466 (N_29466,N_27926,N_27531);
nor U29467 (N_29467,N_26893,N_26470);
nand U29468 (N_29468,N_27718,N_26693);
and U29469 (N_29469,N_26258,N_26301);
xnor U29470 (N_29470,N_27135,N_26373);
nand U29471 (N_29471,N_27466,N_26821);
or U29472 (N_29472,N_27426,N_26775);
and U29473 (N_29473,N_27261,N_27782);
xor U29474 (N_29474,N_27709,N_26650);
and U29475 (N_29475,N_26347,N_27169);
nor U29476 (N_29476,N_27900,N_26127);
and U29477 (N_29477,N_26782,N_26051);
and U29478 (N_29478,N_26202,N_26607);
or U29479 (N_29479,N_27855,N_27043);
nor U29480 (N_29480,N_26155,N_27593);
nor U29481 (N_29481,N_26942,N_27902);
xor U29482 (N_29482,N_27509,N_26840);
and U29483 (N_29483,N_27257,N_26901);
nand U29484 (N_29484,N_26057,N_26989);
and U29485 (N_29485,N_26971,N_26231);
nor U29486 (N_29486,N_26799,N_27168);
and U29487 (N_29487,N_27136,N_27805);
nand U29488 (N_29488,N_27096,N_27701);
xor U29489 (N_29489,N_26177,N_27937);
or U29490 (N_29490,N_26579,N_26262);
and U29491 (N_29491,N_26671,N_26236);
or U29492 (N_29492,N_27381,N_26681);
or U29493 (N_29493,N_27038,N_26915);
xnor U29494 (N_29494,N_27770,N_27709);
nor U29495 (N_29495,N_26437,N_26601);
and U29496 (N_29496,N_26357,N_27833);
nor U29497 (N_29497,N_27264,N_26084);
nor U29498 (N_29498,N_27666,N_26460);
nor U29499 (N_29499,N_26501,N_27057);
or U29500 (N_29500,N_26925,N_27364);
or U29501 (N_29501,N_27693,N_27354);
and U29502 (N_29502,N_27750,N_26679);
nor U29503 (N_29503,N_26130,N_26604);
or U29504 (N_29504,N_27283,N_27034);
nor U29505 (N_29505,N_26589,N_27127);
nand U29506 (N_29506,N_26406,N_27961);
and U29507 (N_29507,N_27444,N_26083);
xor U29508 (N_29508,N_26341,N_27561);
xor U29509 (N_29509,N_27586,N_26962);
xor U29510 (N_29510,N_27978,N_26430);
and U29511 (N_29511,N_27813,N_27316);
or U29512 (N_29512,N_26676,N_26768);
xnor U29513 (N_29513,N_27748,N_26546);
xnor U29514 (N_29514,N_27648,N_26938);
or U29515 (N_29515,N_26376,N_27465);
xnor U29516 (N_29516,N_27290,N_27042);
nor U29517 (N_29517,N_27695,N_26231);
and U29518 (N_29518,N_26812,N_27915);
nor U29519 (N_29519,N_27804,N_26834);
nand U29520 (N_29520,N_27779,N_26454);
xnor U29521 (N_29521,N_26465,N_27468);
nor U29522 (N_29522,N_26767,N_27095);
or U29523 (N_29523,N_27347,N_26866);
xor U29524 (N_29524,N_26230,N_26471);
xnor U29525 (N_29525,N_26153,N_26087);
xor U29526 (N_29526,N_26426,N_26599);
and U29527 (N_29527,N_26206,N_27449);
and U29528 (N_29528,N_26214,N_26888);
nand U29529 (N_29529,N_27915,N_27613);
nor U29530 (N_29530,N_26853,N_26665);
nor U29531 (N_29531,N_27197,N_27991);
nor U29532 (N_29532,N_27937,N_27967);
or U29533 (N_29533,N_26220,N_27748);
and U29534 (N_29534,N_26338,N_26622);
or U29535 (N_29535,N_26206,N_26919);
nand U29536 (N_29536,N_27698,N_26851);
nand U29537 (N_29537,N_27570,N_26323);
nand U29538 (N_29538,N_27575,N_27924);
xor U29539 (N_29539,N_26880,N_27498);
nand U29540 (N_29540,N_26172,N_26814);
nor U29541 (N_29541,N_26471,N_26033);
and U29542 (N_29542,N_27868,N_27148);
or U29543 (N_29543,N_26347,N_27738);
xnor U29544 (N_29544,N_27413,N_26154);
nor U29545 (N_29545,N_26665,N_27283);
nor U29546 (N_29546,N_27951,N_27039);
xor U29547 (N_29547,N_27460,N_26487);
nand U29548 (N_29548,N_26046,N_26701);
and U29549 (N_29549,N_26931,N_26653);
nand U29550 (N_29550,N_26078,N_26833);
or U29551 (N_29551,N_27274,N_26874);
nand U29552 (N_29552,N_27138,N_26611);
and U29553 (N_29553,N_27936,N_27909);
or U29554 (N_29554,N_26510,N_27822);
nand U29555 (N_29555,N_27879,N_26714);
nand U29556 (N_29556,N_27481,N_26866);
and U29557 (N_29557,N_27190,N_27377);
and U29558 (N_29558,N_26696,N_26968);
nor U29559 (N_29559,N_26552,N_27184);
and U29560 (N_29560,N_26385,N_27004);
nand U29561 (N_29561,N_27668,N_26441);
nand U29562 (N_29562,N_27351,N_26867);
and U29563 (N_29563,N_27963,N_27150);
xor U29564 (N_29564,N_27702,N_27235);
or U29565 (N_29565,N_27980,N_27959);
nand U29566 (N_29566,N_26352,N_27192);
nor U29567 (N_29567,N_26607,N_27533);
nand U29568 (N_29568,N_27890,N_27539);
and U29569 (N_29569,N_26851,N_26996);
xor U29570 (N_29570,N_26551,N_27581);
or U29571 (N_29571,N_26220,N_27614);
or U29572 (N_29572,N_26492,N_26830);
xor U29573 (N_29573,N_27236,N_26383);
nand U29574 (N_29574,N_26994,N_26879);
and U29575 (N_29575,N_27280,N_26345);
and U29576 (N_29576,N_27701,N_27897);
and U29577 (N_29577,N_27005,N_27610);
or U29578 (N_29578,N_26352,N_26779);
nor U29579 (N_29579,N_26355,N_26653);
nand U29580 (N_29580,N_26185,N_26552);
or U29581 (N_29581,N_27212,N_26772);
and U29582 (N_29582,N_26364,N_27008);
nand U29583 (N_29583,N_26361,N_27024);
nor U29584 (N_29584,N_27085,N_26657);
and U29585 (N_29585,N_27766,N_27199);
or U29586 (N_29586,N_27397,N_27078);
nor U29587 (N_29587,N_26374,N_26239);
and U29588 (N_29588,N_27133,N_26410);
xnor U29589 (N_29589,N_26217,N_26776);
or U29590 (N_29590,N_26779,N_27134);
and U29591 (N_29591,N_26004,N_26665);
nand U29592 (N_29592,N_26585,N_26467);
xnor U29593 (N_29593,N_26490,N_26764);
and U29594 (N_29594,N_27639,N_26783);
nor U29595 (N_29595,N_27674,N_26076);
nand U29596 (N_29596,N_27905,N_26050);
or U29597 (N_29597,N_26980,N_26086);
xnor U29598 (N_29598,N_26093,N_27406);
and U29599 (N_29599,N_26376,N_26430);
and U29600 (N_29600,N_27109,N_26948);
nor U29601 (N_29601,N_27216,N_26011);
and U29602 (N_29602,N_26333,N_26952);
and U29603 (N_29603,N_26068,N_26881);
and U29604 (N_29604,N_26873,N_26461);
xor U29605 (N_29605,N_26432,N_27196);
nor U29606 (N_29606,N_27034,N_27212);
and U29607 (N_29607,N_27490,N_27045);
nor U29608 (N_29608,N_26602,N_26330);
nand U29609 (N_29609,N_27696,N_27809);
xnor U29610 (N_29610,N_27174,N_26058);
xnor U29611 (N_29611,N_27162,N_27470);
nand U29612 (N_29612,N_27318,N_26196);
or U29613 (N_29613,N_26486,N_27056);
and U29614 (N_29614,N_26909,N_27839);
xor U29615 (N_29615,N_26839,N_27030);
nand U29616 (N_29616,N_27605,N_26737);
and U29617 (N_29617,N_26837,N_27850);
and U29618 (N_29618,N_27790,N_27889);
or U29619 (N_29619,N_27527,N_26745);
nand U29620 (N_29620,N_26598,N_26621);
nor U29621 (N_29621,N_27127,N_26823);
nor U29622 (N_29622,N_27579,N_26084);
nor U29623 (N_29623,N_26002,N_27046);
xnor U29624 (N_29624,N_27636,N_26445);
and U29625 (N_29625,N_27190,N_26412);
and U29626 (N_29626,N_26477,N_26396);
nand U29627 (N_29627,N_26928,N_26343);
xnor U29628 (N_29628,N_26903,N_27682);
and U29629 (N_29629,N_27057,N_26418);
xnor U29630 (N_29630,N_26459,N_26639);
or U29631 (N_29631,N_26891,N_26429);
or U29632 (N_29632,N_26091,N_27076);
xnor U29633 (N_29633,N_27342,N_26376);
or U29634 (N_29634,N_26607,N_26923);
and U29635 (N_29635,N_27717,N_27359);
nor U29636 (N_29636,N_27667,N_26120);
xnor U29637 (N_29637,N_26895,N_26863);
and U29638 (N_29638,N_27639,N_26658);
and U29639 (N_29639,N_27903,N_27831);
and U29640 (N_29640,N_26789,N_26401);
nor U29641 (N_29641,N_26723,N_26855);
nand U29642 (N_29642,N_26556,N_27217);
nand U29643 (N_29643,N_27128,N_27614);
or U29644 (N_29644,N_26820,N_27927);
and U29645 (N_29645,N_26549,N_26608);
xor U29646 (N_29646,N_26779,N_27369);
and U29647 (N_29647,N_27840,N_26985);
nor U29648 (N_29648,N_26507,N_26101);
xor U29649 (N_29649,N_26188,N_27789);
nand U29650 (N_29650,N_27428,N_26148);
and U29651 (N_29651,N_27040,N_27088);
nand U29652 (N_29652,N_26750,N_26518);
and U29653 (N_29653,N_27444,N_27732);
nor U29654 (N_29654,N_27854,N_27448);
or U29655 (N_29655,N_26807,N_26482);
nor U29656 (N_29656,N_26326,N_26610);
nor U29657 (N_29657,N_27092,N_26596);
xor U29658 (N_29658,N_26451,N_26352);
or U29659 (N_29659,N_27491,N_26066);
xor U29660 (N_29660,N_27456,N_26912);
nand U29661 (N_29661,N_26095,N_27836);
nor U29662 (N_29662,N_26662,N_27582);
and U29663 (N_29663,N_27720,N_26117);
and U29664 (N_29664,N_27555,N_27526);
or U29665 (N_29665,N_26412,N_26681);
nor U29666 (N_29666,N_27243,N_27447);
nand U29667 (N_29667,N_26242,N_26593);
or U29668 (N_29668,N_27964,N_26794);
nor U29669 (N_29669,N_26319,N_27571);
xnor U29670 (N_29670,N_26589,N_26818);
nor U29671 (N_29671,N_26455,N_26675);
and U29672 (N_29672,N_26457,N_26932);
xor U29673 (N_29673,N_27837,N_26068);
nor U29674 (N_29674,N_27695,N_27881);
nand U29675 (N_29675,N_27636,N_26900);
nor U29676 (N_29676,N_26260,N_26238);
nand U29677 (N_29677,N_26621,N_27772);
xor U29678 (N_29678,N_26797,N_26875);
or U29679 (N_29679,N_26209,N_27143);
or U29680 (N_29680,N_27670,N_26879);
nand U29681 (N_29681,N_27347,N_27579);
nand U29682 (N_29682,N_26680,N_27673);
and U29683 (N_29683,N_27431,N_26752);
nand U29684 (N_29684,N_26078,N_26741);
nand U29685 (N_29685,N_27495,N_26616);
or U29686 (N_29686,N_26864,N_26257);
xor U29687 (N_29687,N_27396,N_26537);
nand U29688 (N_29688,N_27513,N_26673);
xor U29689 (N_29689,N_27897,N_27542);
nand U29690 (N_29690,N_26064,N_27645);
nand U29691 (N_29691,N_27049,N_27260);
or U29692 (N_29692,N_27600,N_27991);
or U29693 (N_29693,N_27287,N_27365);
nand U29694 (N_29694,N_26429,N_26046);
and U29695 (N_29695,N_27283,N_27288);
or U29696 (N_29696,N_26211,N_27945);
or U29697 (N_29697,N_26786,N_26629);
or U29698 (N_29698,N_26146,N_27587);
and U29699 (N_29699,N_26919,N_27187);
xor U29700 (N_29700,N_26275,N_26929);
or U29701 (N_29701,N_26579,N_27398);
nand U29702 (N_29702,N_27469,N_26687);
or U29703 (N_29703,N_26332,N_27357);
and U29704 (N_29704,N_27259,N_27831);
and U29705 (N_29705,N_26391,N_26426);
or U29706 (N_29706,N_27988,N_26440);
nor U29707 (N_29707,N_27372,N_27225);
nand U29708 (N_29708,N_26384,N_26267);
nand U29709 (N_29709,N_26244,N_27439);
or U29710 (N_29710,N_26822,N_26386);
xnor U29711 (N_29711,N_26325,N_27991);
nor U29712 (N_29712,N_27591,N_26848);
nor U29713 (N_29713,N_27007,N_26476);
nor U29714 (N_29714,N_27067,N_26877);
nand U29715 (N_29715,N_27286,N_26218);
xor U29716 (N_29716,N_27477,N_27447);
nor U29717 (N_29717,N_26611,N_27916);
xor U29718 (N_29718,N_27760,N_26208);
nor U29719 (N_29719,N_27530,N_26531);
or U29720 (N_29720,N_27126,N_26893);
xnor U29721 (N_29721,N_27342,N_27306);
nand U29722 (N_29722,N_26653,N_27535);
nand U29723 (N_29723,N_27771,N_27464);
xor U29724 (N_29724,N_26760,N_27039);
and U29725 (N_29725,N_26773,N_27280);
or U29726 (N_29726,N_26581,N_26756);
nand U29727 (N_29727,N_26054,N_26434);
and U29728 (N_29728,N_26434,N_27740);
and U29729 (N_29729,N_26813,N_27519);
and U29730 (N_29730,N_26891,N_27843);
xnor U29731 (N_29731,N_26435,N_26107);
and U29732 (N_29732,N_27635,N_26239);
nor U29733 (N_29733,N_26212,N_26631);
nand U29734 (N_29734,N_26047,N_26861);
and U29735 (N_29735,N_27104,N_26249);
nand U29736 (N_29736,N_27220,N_27609);
and U29737 (N_29737,N_27088,N_26078);
nor U29738 (N_29738,N_27355,N_26237);
nor U29739 (N_29739,N_26272,N_26516);
or U29740 (N_29740,N_26607,N_26243);
xnor U29741 (N_29741,N_26436,N_27097);
or U29742 (N_29742,N_27254,N_26294);
xor U29743 (N_29743,N_27596,N_26380);
nand U29744 (N_29744,N_26363,N_26619);
or U29745 (N_29745,N_27359,N_27538);
xor U29746 (N_29746,N_26385,N_27305);
xnor U29747 (N_29747,N_27929,N_26871);
nand U29748 (N_29748,N_27225,N_27613);
and U29749 (N_29749,N_27809,N_27430);
xor U29750 (N_29750,N_26801,N_27171);
nand U29751 (N_29751,N_27725,N_26208);
or U29752 (N_29752,N_26101,N_27521);
or U29753 (N_29753,N_26627,N_26460);
and U29754 (N_29754,N_26443,N_27459);
and U29755 (N_29755,N_27034,N_26654);
or U29756 (N_29756,N_26499,N_27413);
and U29757 (N_29757,N_26489,N_26747);
and U29758 (N_29758,N_26411,N_26904);
nand U29759 (N_29759,N_26593,N_27444);
or U29760 (N_29760,N_26215,N_26418);
or U29761 (N_29761,N_27006,N_26181);
and U29762 (N_29762,N_26201,N_27394);
nor U29763 (N_29763,N_26375,N_27103);
xor U29764 (N_29764,N_26265,N_26540);
or U29765 (N_29765,N_26859,N_26205);
nor U29766 (N_29766,N_27194,N_27062);
or U29767 (N_29767,N_27486,N_26724);
xnor U29768 (N_29768,N_26133,N_26484);
nand U29769 (N_29769,N_27736,N_27630);
and U29770 (N_29770,N_27842,N_26886);
and U29771 (N_29771,N_26081,N_26660);
nor U29772 (N_29772,N_27925,N_26888);
or U29773 (N_29773,N_27432,N_26528);
nand U29774 (N_29774,N_27006,N_26515);
and U29775 (N_29775,N_27903,N_26376);
and U29776 (N_29776,N_27604,N_27478);
nand U29777 (N_29777,N_26568,N_27267);
xor U29778 (N_29778,N_27572,N_26587);
or U29779 (N_29779,N_27688,N_27033);
xor U29780 (N_29780,N_27070,N_27888);
and U29781 (N_29781,N_26813,N_26391);
nand U29782 (N_29782,N_26687,N_27287);
xnor U29783 (N_29783,N_26039,N_26272);
xor U29784 (N_29784,N_26189,N_26216);
or U29785 (N_29785,N_26179,N_26570);
nor U29786 (N_29786,N_26273,N_27945);
and U29787 (N_29787,N_27200,N_26692);
nor U29788 (N_29788,N_26321,N_27031);
xor U29789 (N_29789,N_26195,N_27712);
xnor U29790 (N_29790,N_26028,N_26822);
nor U29791 (N_29791,N_27205,N_27295);
nand U29792 (N_29792,N_27891,N_27574);
nand U29793 (N_29793,N_26800,N_27301);
nand U29794 (N_29794,N_26735,N_26829);
and U29795 (N_29795,N_26320,N_27917);
or U29796 (N_29796,N_26199,N_26819);
or U29797 (N_29797,N_27293,N_27876);
nand U29798 (N_29798,N_27156,N_27845);
nand U29799 (N_29799,N_27908,N_26751);
nor U29800 (N_29800,N_27936,N_26758);
nor U29801 (N_29801,N_26908,N_27958);
and U29802 (N_29802,N_27014,N_26064);
nand U29803 (N_29803,N_26048,N_27503);
nand U29804 (N_29804,N_27088,N_27106);
xnor U29805 (N_29805,N_27541,N_26659);
xnor U29806 (N_29806,N_26511,N_26071);
xor U29807 (N_29807,N_26673,N_26768);
and U29808 (N_29808,N_27109,N_26641);
xnor U29809 (N_29809,N_26407,N_26091);
and U29810 (N_29810,N_27210,N_27452);
or U29811 (N_29811,N_27916,N_27478);
nor U29812 (N_29812,N_26128,N_26624);
nand U29813 (N_29813,N_27538,N_27933);
nor U29814 (N_29814,N_27102,N_26928);
nand U29815 (N_29815,N_27987,N_26827);
or U29816 (N_29816,N_26122,N_26999);
and U29817 (N_29817,N_27734,N_26920);
and U29818 (N_29818,N_26014,N_27345);
nor U29819 (N_29819,N_26100,N_27458);
nand U29820 (N_29820,N_26138,N_26595);
or U29821 (N_29821,N_26613,N_27149);
nand U29822 (N_29822,N_26528,N_27109);
xor U29823 (N_29823,N_27749,N_26431);
xor U29824 (N_29824,N_26447,N_26703);
nor U29825 (N_29825,N_27051,N_26903);
nand U29826 (N_29826,N_27370,N_26798);
or U29827 (N_29827,N_27563,N_27919);
or U29828 (N_29828,N_26888,N_27442);
nand U29829 (N_29829,N_27147,N_26141);
and U29830 (N_29830,N_27580,N_27877);
xor U29831 (N_29831,N_26512,N_26138);
xnor U29832 (N_29832,N_26886,N_27004);
nand U29833 (N_29833,N_26928,N_27426);
nand U29834 (N_29834,N_27750,N_27592);
xnor U29835 (N_29835,N_27812,N_27187);
and U29836 (N_29836,N_26812,N_27939);
or U29837 (N_29837,N_26341,N_27818);
nand U29838 (N_29838,N_26641,N_26873);
xnor U29839 (N_29839,N_26878,N_27057);
nand U29840 (N_29840,N_26812,N_26378);
nor U29841 (N_29841,N_27590,N_27678);
nor U29842 (N_29842,N_26985,N_27469);
or U29843 (N_29843,N_27597,N_26184);
or U29844 (N_29844,N_26809,N_27233);
xor U29845 (N_29845,N_27219,N_27220);
nand U29846 (N_29846,N_27933,N_27945);
xnor U29847 (N_29847,N_26042,N_26416);
nand U29848 (N_29848,N_26690,N_27964);
xor U29849 (N_29849,N_27924,N_26400);
xor U29850 (N_29850,N_27623,N_27092);
xnor U29851 (N_29851,N_26749,N_26952);
nand U29852 (N_29852,N_27522,N_26419);
nor U29853 (N_29853,N_26082,N_26868);
nor U29854 (N_29854,N_26487,N_26116);
nand U29855 (N_29855,N_26383,N_27912);
nand U29856 (N_29856,N_27647,N_27588);
or U29857 (N_29857,N_27341,N_27702);
and U29858 (N_29858,N_27982,N_26679);
or U29859 (N_29859,N_27033,N_26895);
or U29860 (N_29860,N_26644,N_26122);
xnor U29861 (N_29861,N_26977,N_27169);
xnor U29862 (N_29862,N_27826,N_27383);
nand U29863 (N_29863,N_26644,N_26407);
or U29864 (N_29864,N_26580,N_26933);
xnor U29865 (N_29865,N_26258,N_27004);
and U29866 (N_29866,N_26884,N_26023);
nand U29867 (N_29867,N_27075,N_27363);
xnor U29868 (N_29868,N_27927,N_26621);
xnor U29869 (N_29869,N_27571,N_27904);
nor U29870 (N_29870,N_26893,N_27749);
nand U29871 (N_29871,N_27924,N_27142);
or U29872 (N_29872,N_26509,N_27776);
and U29873 (N_29873,N_27584,N_26918);
or U29874 (N_29874,N_27214,N_26649);
xnor U29875 (N_29875,N_27233,N_26866);
and U29876 (N_29876,N_27636,N_27680);
nor U29877 (N_29877,N_27935,N_27195);
and U29878 (N_29878,N_27981,N_27846);
and U29879 (N_29879,N_26801,N_27099);
nor U29880 (N_29880,N_26285,N_27055);
nand U29881 (N_29881,N_26563,N_27991);
nor U29882 (N_29882,N_27032,N_27755);
nand U29883 (N_29883,N_27401,N_26748);
or U29884 (N_29884,N_26389,N_27946);
xnor U29885 (N_29885,N_26480,N_26446);
xor U29886 (N_29886,N_27848,N_27899);
xor U29887 (N_29887,N_26883,N_26512);
or U29888 (N_29888,N_27319,N_26693);
or U29889 (N_29889,N_26038,N_27264);
and U29890 (N_29890,N_27560,N_26322);
nand U29891 (N_29891,N_27330,N_26914);
nor U29892 (N_29892,N_26276,N_27882);
xor U29893 (N_29893,N_26669,N_26433);
and U29894 (N_29894,N_26224,N_27388);
nor U29895 (N_29895,N_27072,N_27917);
xnor U29896 (N_29896,N_27345,N_26665);
or U29897 (N_29897,N_27775,N_27394);
or U29898 (N_29898,N_26433,N_26371);
nor U29899 (N_29899,N_27931,N_26474);
and U29900 (N_29900,N_27505,N_27670);
nor U29901 (N_29901,N_27637,N_26644);
or U29902 (N_29902,N_27192,N_26509);
nor U29903 (N_29903,N_27708,N_27512);
and U29904 (N_29904,N_26023,N_26999);
xor U29905 (N_29905,N_27136,N_26797);
and U29906 (N_29906,N_26856,N_26455);
nand U29907 (N_29907,N_26057,N_26757);
or U29908 (N_29908,N_27857,N_26825);
nand U29909 (N_29909,N_26936,N_26944);
xor U29910 (N_29910,N_26930,N_27445);
nand U29911 (N_29911,N_27734,N_26748);
nand U29912 (N_29912,N_26006,N_27497);
and U29913 (N_29913,N_26493,N_26742);
or U29914 (N_29914,N_27290,N_26619);
nand U29915 (N_29915,N_27698,N_27330);
xnor U29916 (N_29916,N_27259,N_26253);
nand U29917 (N_29917,N_26566,N_27966);
nor U29918 (N_29918,N_27702,N_27923);
or U29919 (N_29919,N_27514,N_26320);
and U29920 (N_29920,N_26862,N_26872);
nand U29921 (N_29921,N_27160,N_26803);
nor U29922 (N_29922,N_26045,N_26073);
or U29923 (N_29923,N_27861,N_27300);
and U29924 (N_29924,N_27322,N_26429);
xnor U29925 (N_29925,N_27610,N_26757);
nand U29926 (N_29926,N_26267,N_26792);
nor U29927 (N_29927,N_27957,N_27372);
nor U29928 (N_29928,N_26435,N_27462);
xor U29929 (N_29929,N_27574,N_26428);
and U29930 (N_29930,N_26740,N_26969);
or U29931 (N_29931,N_26231,N_27130);
nor U29932 (N_29932,N_27144,N_26798);
xor U29933 (N_29933,N_26736,N_26744);
nand U29934 (N_29934,N_27435,N_27623);
nor U29935 (N_29935,N_27644,N_27189);
and U29936 (N_29936,N_26745,N_27341);
and U29937 (N_29937,N_26587,N_26019);
xnor U29938 (N_29938,N_26062,N_27988);
or U29939 (N_29939,N_26507,N_27647);
nor U29940 (N_29940,N_27676,N_27053);
nand U29941 (N_29941,N_27030,N_26591);
nor U29942 (N_29942,N_26076,N_26088);
xnor U29943 (N_29943,N_27492,N_27053);
nor U29944 (N_29944,N_27173,N_27665);
xnor U29945 (N_29945,N_27514,N_27311);
nand U29946 (N_29946,N_26501,N_27061);
nand U29947 (N_29947,N_27861,N_26127);
xor U29948 (N_29948,N_26870,N_27952);
and U29949 (N_29949,N_27965,N_27597);
nand U29950 (N_29950,N_27904,N_26373);
or U29951 (N_29951,N_27202,N_26019);
nor U29952 (N_29952,N_27925,N_26411);
nor U29953 (N_29953,N_27807,N_26286);
xnor U29954 (N_29954,N_27004,N_27265);
xor U29955 (N_29955,N_26178,N_27877);
or U29956 (N_29956,N_27242,N_27480);
nor U29957 (N_29957,N_26871,N_27567);
xnor U29958 (N_29958,N_26033,N_27953);
nor U29959 (N_29959,N_26497,N_26042);
nand U29960 (N_29960,N_27261,N_26769);
xnor U29961 (N_29961,N_26367,N_27162);
xor U29962 (N_29962,N_27808,N_26480);
nand U29963 (N_29963,N_27875,N_26220);
xnor U29964 (N_29964,N_26302,N_26439);
nor U29965 (N_29965,N_27682,N_26017);
and U29966 (N_29966,N_27218,N_26897);
nor U29967 (N_29967,N_27982,N_26021);
nand U29968 (N_29968,N_27687,N_27936);
nand U29969 (N_29969,N_26991,N_27344);
xor U29970 (N_29970,N_27604,N_26743);
xor U29971 (N_29971,N_26209,N_27722);
or U29972 (N_29972,N_27683,N_27476);
xnor U29973 (N_29973,N_27151,N_26974);
nor U29974 (N_29974,N_26079,N_27122);
or U29975 (N_29975,N_27240,N_27446);
and U29976 (N_29976,N_26434,N_27289);
xnor U29977 (N_29977,N_27129,N_27888);
and U29978 (N_29978,N_27350,N_27418);
nand U29979 (N_29979,N_26662,N_27886);
xnor U29980 (N_29980,N_26344,N_27000);
nand U29981 (N_29981,N_26801,N_27823);
or U29982 (N_29982,N_27339,N_26422);
or U29983 (N_29983,N_26074,N_26041);
and U29984 (N_29984,N_27824,N_26126);
or U29985 (N_29985,N_26576,N_27203);
or U29986 (N_29986,N_27549,N_27569);
and U29987 (N_29987,N_26590,N_27130);
nor U29988 (N_29988,N_26036,N_27480);
and U29989 (N_29989,N_26954,N_27118);
nor U29990 (N_29990,N_26317,N_26947);
and U29991 (N_29991,N_26845,N_27581);
nor U29992 (N_29992,N_26790,N_27412);
nor U29993 (N_29993,N_26195,N_26227);
nor U29994 (N_29994,N_26599,N_27807);
and U29995 (N_29995,N_27364,N_27886);
and U29996 (N_29996,N_27485,N_26587);
or U29997 (N_29997,N_27792,N_27780);
nor U29998 (N_29998,N_26248,N_26986);
nor U29999 (N_29999,N_26258,N_26344);
nand UO_0 (O_0,N_29167,N_28728);
and UO_1 (O_1,N_29753,N_29342);
or UO_2 (O_2,N_29749,N_29098);
nor UO_3 (O_3,N_28659,N_29690);
xor UO_4 (O_4,N_28428,N_29919);
xnor UO_5 (O_5,N_29268,N_29818);
nand UO_6 (O_6,N_28518,N_29468);
or UO_7 (O_7,N_29909,N_28073);
or UO_8 (O_8,N_28657,N_28268);
or UO_9 (O_9,N_28893,N_28612);
nor UO_10 (O_10,N_28590,N_29899);
nor UO_11 (O_11,N_28743,N_29443);
nand UO_12 (O_12,N_28497,N_29787);
and UO_13 (O_13,N_29625,N_29374);
and UO_14 (O_14,N_28969,N_28228);
and UO_15 (O_15,N_29738,N_28062);
or UO_16 (O_16,N_28017,N_28187);
or UO_17 (O_17,N_29300,N_29571);
or UO_18 (O_18,N_28575,N_28248);
and UO_19 (O_19,N_28867,N_28795);
or UO_20 (O_20,N_29890,N_29339);
nand UO_21 (O_21,N_28512,N_28735);
xor UO_22 (O_22,N_29769,N_29981);
nor UO_23 (O_23,N_29553,N_28463);
nand UO_24 (O_24,N_28613,N_28899);
and UO_25 (O_25,N_29608,N_29499);
nor UO_26 (O_26,N_28255,N_28979);
and UO_27 (O_27,N_29770,N_29520);
nand UO_28 (O_28,N_28666,N_28888);
or UO_29 (O_29,N_28894,N_28176);
and UO_30 (O_30,N_28038,N_29146);
nor UO_31 (O_31,N_29014,N_29454);
nand UO_32 (O_32,N_28812,N_29871);
nand UO_33 (O_33,N_28045,N_29889);
and UO_34 (O_34,N_29228,N_28383);
xnor UO_35 (O_35,N_28593,N_28323);
or UO_36 (O_36,N_29123,N_29996);
nand UO_37 (O_37,N_29995,N_29324);
and UO_38 (O_38,N_29430,N_29376);
xnor UO_39 (O_39,N_28199,N_29309);
nand UO_40 (O_40,N_28909,N_28193);
nand UO_41 (O_41,N_29657,N_29286);
nand UO_42 (O_42,N_28422,N_28364);
nor UO_43 (O_43,N_29351,N_28142);
xnor UO_44 (O_44,N_28445,N_29932);
nor UO_45 (O_45,N_28389,N_28907);
or UO_46 (O_46,N_29370,N_28646);
nand UO_47 (O_47,N_28699,N_28799);
and UO_48 (O_48,N_29176,N_28037);
and UO_49 (O_49,N_29629,N_29857);
and UO_50 (O_50,N_29858,N_29706);
and UO_51 (O_51,N_29179,N_28970);
and UO_52 (O_52,N_29435,N_28656);
nor UO_53 (O_53,N_29739,N_28696);
and UO_54 (O_54,N_29208,N_29360);
nor UO_55 (O_55,N_29204,N_28610);
or UO_56 (O_56,N_29106,N_28502);
nand UO_57 (O_57,N_29137,N_29537);
nor UO_58 (O_58,N_29728,N_29810);
nand UO_59 (O_59,N_29955,N_28031);
and UO_60 (O_60,N_29595,N_29085);
or UO_61 (O_61,N_29646,N_28474);
or UO_62 (O_62,N_29425,N_28480);
nand UO_63 (O_63,N_28857,N_28379);
or UO_64 (O_64,N_28252,N_29698);
xor UO_65 (O_65,N_29424,N_28608);
nor UO_66 (O_66,N_28658,N_29659);
xor UO_67 (O_67,N_29515,N_29539);
or UO_68 (O_68,N_28604,N_28543);
nor UO_69 (O_69,N_29860,N_28594);
nand UO_70 (O_70,N_28546,N_28592);
or UO_71 (O_71,N_28082,N_28053);
or UO_72 (O_72,N_28623,N_28274);
xnor UO_73 (O_73,N_29131,N_28832);
and UO_74 (O_74,N_29357,N_29151);
and UO_75 (O_75,N_28689,N_28309);
nor UO_76 (O_76,N_29641,N_29777);
xor UO_77 (O_77,N_28436,N_29058);
or UO_78 (O_78,N_29241,N_28808);
or UO_79 (O_79,N_29980,N_29001);
or UO_80 (O_80,N_29295,N_29631);
and UO_81 (O_81,N_28457,N_28377);
nand UO_82 (O_82,N_29596,N_29516);
nor UO_83 (O_83,N_28516,N_29600);
and UO_84 (O_84,N_29437,N_28357);
or UO_85 (O_85,N_29110,N_28793);
and UO_86 (O_86,N_28317,N_29707);
xnor UO_87 (O_87,N_28103,N_29475);
and UO_88 (O_88,N_29648,N_29220);
nand UO_89 (O_89,N_28640,N_29051);
and UO_90 (O_90,N_29299,N_28151);
nand UO_91 (O_91,N_28353,N_28624);
or UO_92 (O_92,N_29733,N_28257);
xnor UO_93 (O_93,N_28496,N_28814);
nor UO_94 (O_94,N_29122,N_29675);
xor UO_95 (O_95,N_28711,N_29288);
and UO_96 (O_96,N_29103,N_28064);
xnor UO_97 (O_97,N_28634,N_28256);
nand UO_98 (O_98,N_29916,N_28720);
nor UO_99 (O_99,N_28788,N_29084);
and UO_100 (O_100,N_28966,N_28362);
nand UO_101 (O_101,N_29418,N_28755);
nand UO_102 (O_102,N_29081,N_29121);
xor UO_103 (O_103,N_29813,N_29958);
and UO_104 (O_104,N_29802,N_28527);
and UO_105 (O_105,N_29774,N_28181);
xnor UO_106 (O_106,N_28940,N_28475);
nor UO_107 (O_107,N_28765,N_29400);
xor UO_108 (O_108,N_28084,N_29908);
xor UO_109 (O_109,N_29509,N_28363);
nand UO_110 (O_110,N_29593,N_29464);
nand UO_111 (O_111,N_28169,N_29135);
nor UO_112 (O_112,N_28571,N_28669);
and UO_113 (O_113,N_28300,N_28579);
xnor UO_114 (O_114,N_28349,N_29136);
or UO_115 (O_115,N_29294,N_29594);
nand UO_116 (O_116,N_28304,N_28886);
nand UO_117 (O_117,N_29399,N_29394);
and UO_118 (O_118,N_28729,N_28553);
or UO_119 (O_119,N_29637,N_28416);
nand UO_120 (O_120,N_28750,N_28742);
or UO_121 (O_121,N_28314,N_29301);
xnor UO_122 (O_122,N_29969,N_28558);
xnor UO_123 (O_123,N_28227,N_29444);
nand UO_124 (O_124,N_29613,N_28850);
nand UO_125 (O_125,N_28266,N_28050);
or UO_126 (O_126,N_28506,N_29233);
nor UO_127 (O_127,N_28757,N_29460);
nand UO_128 (O_128,N_29002,N_28514);
or UO_129 (O_129,N_28954,N_29705);
and UO_130 (O_130,N_29822,N_28091);
nand UO_131 (O_131,N_28213,N_28431);
and UO_132 (O_132,N_28839,N_29589);
xor UO_133 (O_133,N_29512,N_28826);
and UO_134 (O_134,N_29927,N_28642);
xor UO_135 (O_135,N_29171,N_28901);
and UO_136 (O_136,N_29290,N_28712);
nor UO_137 (O_137,N_29582,N_29105);
nor UO_138 (O_138,N_29789,N_28411);
xor UO_139 (O_139,N_28110,N_28835);
or UO_140 (O_140,N_28589,N_29297);
or UO_141 (O_141,N_29853,N_28980);
nand UO_142 (O_142,N_28405,N_29148);
and UO_143 (O_143,N_28427,N_29074);
and UO_144 (O_144,N_29132,N_28987);
and UO_145 (O_145,N_29320,N_28773);
or UO_146 (O_146,N_29993,N_29611);
xnor UO_147 (O_147,N_29476,N_29481);
nor UO_148 (O_148,N_29238,N_28885);
nor UO_149 (O_149,N_28264,N_29182);
or UO_150 (O_150,N_28495,N_28399);
or UO_151 (O_151,N_29569,N_29108);
xor UO_152 (O_152,N_29771,N_28749);
and UO_153 (O_153,N_28925,N_29163);
nand UO_154 (O_154,N_28762,N_28845);
or UO_155 (O_155,N_28034,N_29727);
xnor UO_156 (O_156,N_29130,N_28004);
nand UO_157 (O_157,N_29213,N_28419);
nand UO_158 (O_158,N_28803,N_29172);
nor UO_159 (O_159,N_28680,N_28087);
nand UO_160 (O_160,N_29905,N_29579);
nor UO_161 (O_161,N_29005,N_29231);
nand UO_162 (O_162,N_29102,N_29494);
nand UO_163 (O_163,N_28129,N_28166);
xor UO_164 (O_164,N_29164,N_29111);
nor UO_165 (O_165,N_29284,N_29104);
nor UO_166 (O_166,N_29188,N_29057);
or UO_167 (O_167,N_28878,N_29990);
nor UO_168 (O_168,N_29925,N_28414);
or UO_169 (O_169,N_28770,N_28124);
or UO_170 (O_170,N_28697,N_29038);
nor UO_171 (O_171,N_28410,N_29948);
and UO_172 (O_172,N_28498,N_29071);
and UO_173 (O_173,N_29258,N_28439);
and UO_174 (O_174,N_29793,N_28133);
or UO_175 (O_175,N_28488,N_28171);
and UO_176 (O_176,N_28718,N_29183);
nand UO_177 (O_177,N_28535,N_29712);
xnor UO_178 (O_178,N_29851,N_29989);
nand UO_179 (O_179,N_29518,N_28811);
and UO_180 (O_180,N_29432,N_28225);
xnor UO_181 (O_181,N_28201,N_29830);
nor UO_182 (O_182,N_29279,N_29410);
nor UO_183 (O_183,N_28469,N_29350);
and UO_184 (O_184,N_29070,N_29879);
or UO_185 (O_185,N_29506,N_28334);
xnor UO_186 (O_186,N_29703,N_28797);
xor UO_187 (O_187,N_28898,N_28818);
nand UO_188 (O_188,N_28348,N_28632);
nand UO_189 (O_189,N_29129,N_28967);
xor UO_190 (O_190,N_28200,N_28306);
xnor UO_191 (O_191,N_28097,N_28597);
and UO_192 (O_192,N_29364,N_29797);
or UO_193 (O_193,N_28552,N_29940);
and UO_194 (O_194,N_29356,N_28965);
nor UO_195 (O_195,N_28173,N_29689);
or UO_196 (O_196,N_29904,N_29881);
or UO_197 (O_197,N_29758,N_29367);
and UO_198 (O_198,N_28574,N_28816);
or UO_199 (O_199,N_29722,N_28989);
or UO_200 (O_200,N_29549,N_29599);
xnor UO_201 (O_201,N_29216,N_29209);
nand UO_202 (O_202,N_29999,N_28260);
xor UO_203 (O_203,N_29974,N_29782);
or UO_204 (O_204,N_28329,N_29575);
nor UO_205 (O_205,N_28703,N_29406);
xnor UO_206 (O_206,N_28378,N_29732);
nor UO_207 (O_207,N_29679,N_29378);
or UO_208 (O_208,N_29704,N_28450);
and UO_209 (O_209,N_29710,N_28123);
nand UO_210 (O_210,N_29152,N_29282);
xnor UO_211 (O_211,N_29823,N_29740);
nand UO_212 (O_212,N_29363,N_29429);
nor UO_213 (O_213,N_28067,N_28607);
xor UO_214 (O_214,N_28690,N_28351);
or UO_215 (O_215,N_28057,N_28154);
and UO_216 (O_216,N_29413,N_29361);
nand UO_217 (O_217,N_28098,N_28043);
xor UO_218 (O_218,N_28111,N_28860);
nor UO_219 (O_219,N_28635,N_28510);
xor UO_220 (O_220,N_28000,N_28541);
nor UO_221 (O_221,N_29168,N_28483);
and UO_222 (O_222,N_29101,N_28930);
or UO_223 (O_223,N_28270,N_29820);
nor UO_224 (O_224,N_29161,N_28961);
nand UO_225 (O_225,N_29345,N_28112);
and UO_226 (O_226,N_29828,N_28320);
and UO_227 (O_227,N_28408,N_28752);
or UO_228 (O_228,N_29626,N_29480);
xnor UO_229 (O_229,N_28606,N_28233);
and UO_230 (O_230,N_28873,N_29191);
and UO_231 (O_231,N_29700,N_28239);
and UO_232 (O_232,N_28332,N_28008);
nand UO_233 (O_233,N_29692,N_28245);
xnor UO_234 (O_234,N_28948,N_29773);
nor UO_235 (O_235,N_28175,N_28707);
nand UO_236 (O_236,N_29040,N_28354);
nor UO_237 (O_237,N_29497,N_28605);
nor UO_238 (O_238,N_28356,N_28958);
or UO_239 (O_239,N_28501,N_28026);
xnor UO_240 (O_240,N_28714,N_28588);
nand UO_241 (O_241,N_29023,N_28372);
and UO_242 (O_242,N_28023,N_28149);
and UO_243 (O_243,N_29651,N_29620);
and UO_244 (O_244,N_28027,N_29786);
nand UO_245 (O_245,N_28157,N_28307);
nand UO_246 (O_246,N_28039,N_29165);
xor UO_247 (O_247,N_29293,N_29352);
nor UO_248 (O_248,N_29459,N_29697);
xor UO_249 (O_249,N_29859,N_28188);
or UO_250 (O_250,N_29368,N_29959);
nand UO_251 (O_251,N_28631,N_28207);
or UO_252 (O_252,N_29489,N_28459);
or UO_253 (O_253,N_28924,N_29092);
nand UO_254 (O_254,N_28681,N_28194);
xor UO_255 (O_255,N_29610,N_29551);
or UO_256 (O_256,N_28125,N_29100);
nor UO_257 (O_257,N_28993,N_29982);
nor UO_258 (O_258,N_28204,N_29125);
nand UO_259 (O_259,N_28550,N_28611);
nand UO_260 (O_260,N_28494,N_29457);
and UO_261 (O_261,N_29186,N_28345);
nand UO_262 (O_262,N_28517,N_29096);
nor UO_263 (O_263,N_29086,N_28929);
nor UO_264 (O_264,N_29484,N_28100);
and UO_265 (O_265,N_28366,N_29012);
nand UO_266 (O_266,N_29353,N_28020);
nor UO_267 (O_267,N_28025,N_29478);
or UO_268 (O_268,N_29112,N_29854);
nand UO_269 (O_269,N_28990,N_28708);
and UO_270 (O_270,N_29466,N_29650);
or UO_271 (O_271,N_29701,N_28880);
and UO_272 (O_272,N_28108,N_28802);
xnor UO_273 (O_273,N_28296,N_29546);
or UO_274 (O_274,N_28344,N_29614);
xor UO_275 (O_275,N_28400,N_29319);
or UO_276 (O_276,N_28406,N_28069);
nand UO_277 (O_277,N_29560,N_29415);
nand UO_278 (O_278,N_29045,N_29778);
nand UO_279 (O_279,N_28817,N_28163);
nand UO_280 (O_280,N_28944,N_29630);
nor UO_281 (O_281,N_28805,N_29225);
or UO_282 (O_282,N_29721,N_29482);
nor UO_283 (O_283,N_28784,N_28555);
xor UO_284 (O_284,N_29744,N_28991);
nand UO_285 (O_285,N_28210,N_29652);
xor UO_286 (O_286,N_29156,N_29331);
nor UO_287 (O_287,N_28614,N_29672);
nand UO_288 (O_288,N_29844,N_28758);
nor UO_289 (O_289,N_28951,N_28879);
nand UO_290 (O_290,N_28782,N_28912);
nor UO_291 (O_291,N_29662,N_29903);
nor UO_292 (O_292,N_28325,N_29195);
nor UO_293 (O_293,N_28197,N_29197);
or UO_294 (O_294,N_29775,N_28582);
nand UO_295 (O_295,N_28537,N_28783);
nand UO_296 (O_296,N_29387,N_29139);
or UO_297 (O_297,N_29262,N_28934);
nor UO_298 (O_298,N_28916,N_29267);
nand UO_299 (O_299,N_29439,N_28897);
xnor UO_300 (O_300,N_29465,N_28144);
and UO_301 (O_301,N_28823,N_28807);
nor UO_302 (O_302,N_29042,N_29063);
xor UO_303 (O_303,N_28074,N_28371);
nand UO_304 (O_304,N_29442,N_29649);
or UO_305 (O_305,N_29962,N_28745);
and UO_306 (O_306,N_29261,N_29952);
or UO_307 (O_307,N_28596,N_29335);
nor UO_308 (O_308,N_29619,N_29486);
nand UO_309 (O_309,N_28305,N_29886);
nor UO_310 (O_310,N_29597,N_29696);
and UO_311 (O_311,N_29142,N_28085);
nand UO_312 (O_312,N_29633,N_28763);
xor UO_313 (O_313,N_28336,N_28913);
nor UO_314 (O_314,N_28779,N_28206);
xnor UO_315 (O_315,N_28024,N_28337);
nand UO_316 (O_316,N_29311,N_28156);
nand UO_317 (O_317,N_29834,N_29150);
xor UO_318 (O_318,N_29380,N_29157);
or UO_319 (O_319,N_29665,N_28568);
xor UO_320 (O_320,N_28941,N_29615);
and UO_321 (O_321,N_28215,N_28504);
or UO_322 (O_322,N_28367,N_28395);
and UO_323 (O_323,N_28016,N_29862);
nor UO_324 (O_324,N_29408,N_28955);
xnor UO_325 (O_325,N_28704,N_29416);
or UO_326 (O_326,N_28397,N_29627);
and UO_327 (O_327,N_29166,N_29391);
nand UO_328 (O_328,N_28922,N_28633);
nor UO_329 (O_329,N_29711,N_29934);
nor UO_330 (O_330,N_28122,N_29799);
or UO_331 (O_331,N_28778,N_28937);
nand UO_332 (O_332,N_29354,N_29988);
and UO_333 (O_333,N_28781,N_29530);
nand UO_334 (O_334,N_29906,N_28855);
xor UO_335 (O_335,N_29073,N_29323);
and UO_336 (O_336,N_28468,N_29094);
nor UO_337 (O_337,N_29436,N_29382);
or UO_338 (O_338,N_29998,N_28645);
and UO_339 (O_339,N_29082,N_28914);
or UO_340 (O_340,N_29003,N_29894);
and UO_341 (O_341,N_28919,N_29237);
xnor UO_342 (O_342,N_29053,N_28287);
nor UO_343 (O_343,N_28977,N_29029);
and UO_344 (O_344,N_28787,N_28198);
nand UO_345 (O_345,N_28202,N_29762);
xnor UO_346 (O_346,N_28080,N_29419);
and UO_347 (O_347,N_29236,N_28903);
nor UO_348 (O_348,N_29963,N_28283);
nor UO_349 (O_349,N_28895,N_28375);
nor UO_350 (O_350,N_28716,N_28569);
xor UO_351 (O_351,N_28281,N_28828);
nand UO_352 (O_352,N_29017,N_29240);
xnor UO_353 (O_353,N_29785,N_28286);
or UO_354 (O_354,N_29020,N_28813);
or UO_355 (O_355,N_29984,N_29377);
nor UO_356 (O_356,N_28237,N_29717);
nand UO_357 (O_357,N_29992,N_29768);
xor UO_358 (O_358,N_29059,N_29117);
or UO_359 (O_359,N_29107,N_28259);
and UO_360 (O_360,N_29751,N_28838);
nor UO_361 (O_361,N_29557,N_28789);
nand UO_362 (O_362,N_29227,N_28627);
nand UO_363 (O_363,N_29067,N_28715);
nor UO_364 (O_364,N_29603,N_29937);
and UO_365 (O_365,N_28946,N_28126);
nor UO_366 (O_366,N_28524,N_29756);
nor UO_367 (O_367,N_28942,N_28923);
nand UO_368 (O_368,N_28282,N_29861);
nand UO_369 (O_369,N_28051,N_28682);
and UO_370 (O_370,N_28819,N_29542);
xnor UO_371 (O_371,N_28479,N_29495);
nand UO_372 (O_372,N_29477,N_29809);
nand UO_373 (O_373,N_28068,N_29907);
and UO_374 (O_374,N_28713,N_28675);
xor UO_375 (O_375,N_29901,N_29490);
and UO_376 (O_376,N_28908,N_29215);
or UO_377 (O_377,N_29099,N_29930);
or UO_378 (O_378,N_28920,N_29332);
xnor UO_379 (O_379,N_29694,N_29337);
nor UO_380 (O_380,N_29283,N_28858);
and UO_381 (O_381,N_28491,N_29461);
xor UO_382 (O_382,N_28285,N_28263);
xnor UO_383 (O_383,N_28983,N_29147);
or UO_384 (O_384,N_28476,N_29517);
xor UO_385 (O_385,N_28321,N_28036);
xnor UO_386 (O_386,N_29863,N_29018);
nor UO_387 (O_387,N_28721,N_29445);
nand UO_388 (O_388,N_29741,N_29845);
nand UO_389 (O_389,N_29050,N_28905);
nand UO_390 (O_390,N_29093,N_28441);
nand UO_391 (O_391,N_29688,N_28090);
and UO_392 (O_392,N_28709,N_29056);
xor UO_393 (O_393,N_29212,N_29522);
or UO_394 (O_394,N_28086,N_28978);
xnor UO_395 (O_395,N_28449,N_29421);
nor UO_396 (O_396,N_28297,N_28896);
xor UO_397 (O_397,N_28007,N_28220);
nand UO_398 (O_398,N_29158,N_29748);
nor UO_399 (O_399,N_28560,N_29805);
and UO_400 (O_400,N_28798,N_28780);
nor UO_401 (O_401,N_29848,N_29313);
xor UO_402 (O_402,N_28679,N_29961);
xor UO_403 (O_403,N_29849,N_29726);
xor UO_404 (O_404,N_29069,N_29316);
nor UO_405 (O_405,N_29398,N_29395);
xor UO_406 (O_406,N_29967,N_28028);
nand UO_407 (O_407,N_29973,N_29434);
nor UO_408 (O_408,N_29529,N_28078);
nor UO_409 (O_409,N_29054,N_28767);
nor UO_410 (O_410,N_28424,N_28710);
nor UO_411 (O_411,N_29022,N_28443);
or UO_412 (O_412,N_29184,N_28121);
nand UO_413 (O_413,N_29779,N_28644);
nand UO_414 (O_414,N_28677,N_29624);
xor UO_415 (O_415,N_29939,N_29878);
or UO_416 (O_416,N_29884,N_28727);
and UO_417 (O_417,N_28350,N_28327);
nor UO_418 (O_418,N_29587,N_28792);
nand UO_419 (O_419,N_28861,N_28927);
nor UO_420 (O_420,N_28018,N_28310);
and UO_421 (O_421,N_28576,N_28275);
nand UO_422 (O_422,N_28772,N_29177);
or UO_423 (O_423,N_29255,N_28380);
nor UO_424 (O_424,N_28869,N_29761);
and UO_425 (O_425,N_28161,N_29663);
nor UO_426 (O_426,N_29016,N_28686);
nand UO_427 (O_427,N_29329,N_29383);
xor UO_428 (O_428,N_28700,N_28047);
and UO_429 (O_429,N_29470,N_28153);
or UO_430 (O_430,N_28330,N_28326);
or UO_431 (O_431,N_28771,N_29302);
nand UO_432 (O_432,N_29997,N_29162);
or UO_433 (O_433,N_28670,N_28526);
or UO_434 (O_434,N_28949,N_29508);
nand UO_435 (O_435,N_29242,N_29766);
nand UO_436 (O_436,N_29680,N_28190);
nand UO_437 (O_437,N_29836,N_28209);
xor UO_438 (O_438,N_28600,N_29533);
or UO_439 (O_439,N_28598,N_29338);
or UO_440 (O_440,N_28661,N_28099);
xnor UO_441 (O_441,N_29348,N_29764);
nor UO_442 (O_442,N_29257,N_29221);
nand UO_443 (O_443,N_29790,N_28584);
xnor UO_444 (O_444,N_28691,N_29032);
or UO_445 (O_445,N_28877,N_29260);
xor UO_446 (O_446,N_29562,N_29666);
xnor UO_447 (O_447,N_29654,N_28820);
xnor UO_448 (O_448,N_29140,N_28196);
or UO_449 (O_449,N_28186,N_29089);
nand UO_450 (O_450,N_29501,N_28048);
xor UO_451 (O_451,N_28971,N_28261);
and UO_452 (O_452,N_28401,N_29676);
xor UO_453 (O_453,N_29826,N_28756);
nand UO_454 (O_454,N_28041,N_28972);
and UO_455 (O_455,N_28417,N_28254);
xor UO_456 (O_456,N_28938,N_29760);
nand UO_457 (O_457,N_29855,N_29691);
and UO_458 (O_458,N_28172,N_29133);
xor UO_459 (O_459,N_29341,N_29816);
nor UO_460 (O_460,N_29420,N_29923);
or UO_461 (O_461,N_29505,N_29735);
nand UO_462 (O_462,N_28164,N_28688);
or UO_463 (O_463,N_29892,N_28208);
or UO_464 (O_464,N_29276,N_29604);
or UO_465 (O_465,N_28231,N_29607);
xnor UO_466 (O_466,N_29540,N_29736);
nand UO_467 (O_467,N_29322,N_29548);
and UO_468 (O_468,N_28650,N_29713);
and UO_469 (O_469,N_28654,N_29746);
nand UO_470 (O_470,N_29660,N_28564);
xnor UO_471 (O_471,N_29314,N_28499);
xnor UO_472 (O_472,N_28794,N_28420);
nor UO_473 (O_473,N_29492,N_28015);
nand UO_474 (O_474,N_28141,N_28433);
xnor UO_475 (O_475,N_29547,N_29964);
or UO_476 (O_476,N_28625,N_29469);
and UO_477 (O_477,N_28250,N_29623);
nand UO_478 (O_478,N_28360,N_28071);
xnor UO_479 (O_479,N_28130,N_28019);
or UO_480 (O_480,N_29235,N_29971);
or UO_481 (O_481,N_29566,N_28238);
or UO_482 (O_482,N_29145,N_28148);
nand UO_483 (O_483,N_29839,N_29315);
and UO_484 (O_484,N_28002,N_29291);
nand UO_485 (O_485,N_28890,N_28759);
and UO_486 (O_486,N_28996,N_28132);
nand UO_487 (O_487,N_29372,N_29681);
nand UO_488 (O_488,N_29960,N_28089);
and UO_489 (O_489,N_28643,N_29882);
nor UO_490 (O_490,N_28822,N_28900);
xor UO_491 (O_491,N_28736,N_29577);
nor UO_492 (O_492,N_28009,N_28029);
nor UO_493 (O_493,N_28739,N_28548);
nand UO_494 (O_494,N_28521,N_28962);
nand UO_495 (O_495,N_28407,N_29815);
nor UO_496 (O_496,N_28482,N_28203);
nor UO_497 (O_497,N_29409,N_29333);
nor UO_498 (O_498,N_29921,N_28906);
or UO_499 (O_499,N_29896,N_29668);
nor UO_500 (O_500,N_29280,N_29827);
nand UO_501 (O_501,N_28726,N_29393);
or UO_502 (O_502,N_28603,N_28904);
xnor UO_503 (O_503,N_28288,N_28649);
or UO_504 (O_504,N_29814,N_28724);
xnor UO_505 (O_505,N_29504,N_28421);
nor UO_506 (O_506,N_29060,N_29556);
and UO_507 (O_507,N_29328,N_28134);
nor UO_508 (O_508,N_29519,N_29792);
or UO_509 (O_509,N_29891,N_29384);
and UO_510 (O_510,N_28453,N_29966);
and UO_511 (O_511,N_29065,N_28973);
or UO_512 (O_512,N_29895,N_28740);
nand UO_513 (O_513,N_29978,N_29682);
nand UO_514 (O_514,N_29527,N_28120);
xor UO_515 (O_515,N_28520,N_28313);
and UO_516 (O_516,N_29647,N_29015);
nor UO_517 (O_517,N_29965,N_28964);
xnor UO_518 (O_518,N_29423,N_29044);
xnor UO_519 (O_519,N_28581,N_28761);
nand UO_520 (O_520,N_28889,N_29745);
and UO_521 (O_521,N_29304,N_29450);
and UO_522 (O_522,N_28205,N_28106);
and UO_523 (O_523,N_28236,N_28396);
or UO_524 (O_524,N_29039,N_28101);
and UO_525 (O_525,N_28747,N_28044);
and UO_526 (O_526,N_28315,N_29385);
nor UO_527 (O_527,N_28840,N_28147);
nor UO_528 (O_528,N_29173,N_29244);
and UO_529 (O_529,N_28609,N_29277);
or UO_530 (O_530,N_29207,N_28533);
nor UO_531 (O_531,N_28540,N_29931);
and UO_532 (O_532,N_28005,N_29578);
or UO_533 (O_533,N_29496,N_28528);
and UO_534 (O_534,N_28931,N_29911);
nand UO_535 (O_535,N_28992,N_29000);
nand UO_536 (O_536,N_29609,N_29011);
xnor UO_537 (O_537,N_28769,N_28229);
and UO_538 (O_538,N_29234,N_28926);
xor UO_539 (O_539,N_29835,N_29239);
or UO_540 (O_540,N_29426,N_29194);
and UO_541 (O_541,N_29811,N_28694);
xnor UO_542 (O_542,N_29386,N_29946);
and UO_543 (O_543,N_28768,N_28947);
or UO_544 (O_544,N_28295,N_28525);
or UO_545 (O_545,N_29935,N_28279);
or UO_546 (O_546,N_28824,N_29521);
or UO_547 (O_547,N_29334,N_29767);
xor UO_548 (O_548,N_29252,N_28318);
or UO_549 (O_549,N_29189,N_29564);
xor UO_550 (O_550,N_28685,N_29287);
xor UO_551 (O_551,N_28470,N_29975);
xnor UO_552 (O_552,N_28425,N_28751);
nand UO_553 (O_553,N_29754,N_28791);
nor UO_554 (O_554,N_28549,N_29037);
xnor UO_555 (O_555,N_28131,N_28293);
or UO_556 (O_556,N_28738,N_28012);
and UO_557 (O_557,N_28626,N_29273);
xor UO_558 (O_558,N_28055,N_28114);
and UO_559 (O_559,N_29524,N_28663);
nor UO_560 (O_560,N_29513,N_29783);
and UO_561 (O_561,N_28539,N_28096);
nand UO_562 (O_562,N_28705,N_29957);
nor UO_563 (O_563,N_29699,N_29737);
xnor UO_564 (O_564,N_28722,N_28874);
nor UO_565 (O_565,N_28536,N_28311);
or UO_566 (O_566,N_29757,N_28587);
nor UO_567 (O_567,N_28562,N_29729);
or UO_568 (O_568,N_29601,N_29412);
nand UO_569 (O_569,N_28374,N_28219);
nand UO_570 (O_570,N_28719,N_29298);
nor UO_571 (O_571,N_29821,N_28815);
or UO_572 (O_572,N_28801,N_29715);
xor UO_573 (O_573,N_29265,N_28467);
xor UO_574 (O_574,N_28865,N_29035);
nor UO_575 (O_575,N_28246,N_28580);
or UO_576 (O_576,N_28692,N_28945);
xor UO_577 (O_577,N_28471,N_29526);
nor UO_578 (O_578,N_29584,N_28347);
nand UO_579 (O_579,N_28554,N_28853);
nand UO_580 (O_580,N_29214,N_28863);
or UO_581 (O_581,N_28534,N_28403);
or UO_582 (O_582,N_29365,N_29780);
nor UO_583 (O_583,N_29180,N_29772);
or UO_584 (O_584,N_29838,N_28243);
and UO_585 (O_585,N_28278,N_28075);
or UO_586 (O_586,N_28639,N_29635);
xnor UO_587 (O_587,N_29831,N_29318);
xnor UO_588 (O_588,N_28460,N_29369);
or UO_589 (O_589,N_28731,N_28628);
nand UO_590 (O_590,N_29644,N_29027);
nand UO_591 (O_591,N_29543,N_29642);
and UO_592 (O_592,N_29985,N_29272);
xnor UO_593 (O_593,N_28262,N_28185);
nor UO_594 (O_594,N_29281,N_29621);
xor UO_595 (O_595,N_28651,N_29266);
nor UO_596 (O_596,N_29076,N_28218);
nor UO_597 (O_597,N_28076,N_28490);
and UO_598 (O_598,N_29397,N_28871);
and UO_599 (O_599,N_28174,N_28328);
or UO_600 (O_600,N_28346,N_28150);
xnor UO_601 (O_601,N_29083,N_28072);
nand UO_602 (O_602,N_29472,N_29720);
or UO_603 (O_603,N_29572,N_29534);
xor UO_604 (O_604,N_28102,N_29062);
and UO_605 (O_605,N_28432,N_29563);
xor UO_606 (O_606,N_29095,N_29602);
xor UO_607 (O_607,N_29734,N_28104);
and UO_608 (O_608,N_28244,N_28415);
or UO_609 (O_609,N_28409,N_29674);
and UO_610 (O_610,N_29807,N_28162);
nor UO_611 (O_611,N_28585,N_28701);
xnor UO_612 (O_612,N_29928,N_29249);
and UO_613 (O_613,N_28253,N_29833);
and UO_614 (O_614,N_29024,N_29559);
and UO_615 (O_615,N_28145,N_28883);
xor UO_616 (O_616,N_28466,N_28387);
nand UO_617 (O_617,N_28559,N_28361);
nand UO_618 (O_618,N_28830,N_28676);
or UO_619 (O_619,N_28766,N_28061);
nor UO_620 (O_620,N_29887,N_28465);
xor UO_621 (O_621,N_28222,N_28331);
and UO_622 (O_622,N_28376,N_28247);
and UO_623 (O_623,N_28565,N_28664);
and UO_624 (O_624,N_28189,N_28402);
or UO_625 (O_625,N_28732,N_28277);
and UO_626 (O_626,N_29153,N_29924);
and UO_627 (O_627,N_28706,N_29573);
and UO_628 (O_628,N_28294,N_29586);
xnor UO_629 (O_629,N_29910,N_29075);
nor UO_630 (O_630,N_28667,N_28529);
and UO_631 (O_631,N_29446,N_29558);
or UO_632 (O_632,N_29580,N_28981);
xor UO_633 (O_633,N_29956,N_28423);
or UO_634 (O_634,N_29804,N_28982);
nand UO_635 (O_635,N_29243,N_29441);
or UO_636 (O_636,N_29224,N_29598);
xor UO_637 (O_637,N_29922,N_29327);
and UO_638 (O_638,N_29606,N_28505);
nor UO_639 (O_639,N_29683,N_28723);
nand UO_640 (O_640,N_29730,N_28806);
nand UO_641 (O_641,N_29321,N_29405);
and UO_642 (O_642,N_28006,N_28523);
nor UO_643 (O_643,N_29048,N_28968);
xnor UO_644 (O_644,N_29567,N_29856);
nand UO_645 (O_645,N_28183,N_28192);
xnor UO_646 (O_646,N_28875,N_29832);
nor UO_647 (O_647,N_29417,N_29968);
xor UO_648 (O_648,N_29041,N_29210);
or UO_649 (O_649,N_28754,N_29452);
or UO_650 (O_650,N_29574,N_28507);
or UO_651 (O_651,N_29841,N_29392);
nand UO_652 (O_652,N_28511,N_29077);
nand UO_653 (O_653,N_28458,N_28563);
and UO_654 (O_654,N_29535,N_29458);
or UO_655 (O_655,N_29864,N_29763);
nand UO_656 (O_656,N_29639,N_29817);
nor UO_657 (O_657,N_29976,N_28872);
nand UO_658 (O_658,N_29379,N_29256);
and UO_659 (O_659,N_28487,N_29920);
and UO_660 (O_660,N_29401,N_29192);
nand UO_661 (O_661,N_28093,N_29259);
nor UO_662 (O_662,N_29561,N_29428);
xor UO_663 (O_663,N_28660,N_29877);
xor UO_664 (O_664,N_28567,N_29091);
or UO_665 (O_665,N_28140,N_29875);
nor UO_666 (O_666,N_29565,N_28217);
and UO_667 (O_667,N_28083,N_28390);
xor UO_668 (O_668,N_28273,N_29819);
nor UO_669 (O_669,N_29525,N_28586);
xnor UO_670 (O_670,N_29453,N_29634);
and UO_671 (O_671,N_29203,N_29502);
or UO_672 (O_672,N_29473,N_28573);
nand UO_673 (O_673,N_29953,N_28868);
nor UO_674 (O_674,N_28342,N_29719);
or UO_675 (O_675,N_28003,N_29097);
or UO_676 (O_676,N_28876,N_28542);
nand UO_677 (O_677,N_28777,N_29585);
nor UO_678 (O_678,N_28760,N_28013);
and UO_679 (O_679,N_29159,N_28809);
or UO_680 (O_680,N_29883,N_28943);
nor UO_681 (O_681,N_29072,N_28095);
xor UO_682 (O_682,N_28046,N_29708);
nand UO_683 (O_683,N_29031,N_28352);
xor UO_684 (O_684,N_29791,N_29285);
and UO_685 (O_685,N_28444,N_29687);
or UO_686 (O_686,N_29340,N_29278);
nor UO_687 (O_687,N_29036,N_29190);
or UO_688 (O_688,N_28785,N_29116);
xor UO_689 (O_689,N_29004,N_28999);
xor UO_690 (O_690,N_28833,N_29034);
xor UO_691 (O_691,N_29033,N_29307);
and UO_692 (O_692,N_29196,N_28836);
and UO_693 (O_693,N_29912,N_29755);
nor UO_694 (O_694,N_28370,N_29433);
xor UO_695 (O_695,N_28851,N_28301);
and UO_696 (O_696,N_28456,N_28384);
nand UO_697 (O_697,N_28617,N_28412);
nand UO_698 (O_698,N_28339,N_29274);
and UO_699 (O_699,N_28052,N_28746);
xor UO_700 (O_700,N_29493,N_29205);
xnor UO_701 (O_701,N_28139,N_28340);
nor UO_702 (O_702,N_29143,N_29079);
xnor UO_703 (O_703,N_28155,N_28994);
and UO_704 (O_704,N_29296,N_29670);
nand UO_705 (O_705,N_28115,N_29784);
xor UO_706 (O_706,N_29009,N_29622);
or UO_707 (O_707,N_29500,N_28852);
and UO_708 (O_708,N_28088,N_28615);
or UO_709 (O_709,N_29926,N_29343);
nand UO_710 (O_710,N_29685,N_28796);
nor UO_711 (O_711,N_29202,N_29181);
nor UO_712 (O_712,N_28143,N_28519);
xnor UO_713 (O_713,N_28429,N_29375);
nor UO_714 (O_714,N_29149,N_28988);
or UO_715 (O_715,N_29972,N_28065);
nand UO_716 (O_716,N_28481,N_29068);
or UO_717 (O_717,N_29389,N_29918);
nor UO_718 (O_718,N_28269,N_29979);
and UO_719 (O_719,N_28864,N_28040);
nand UO_720 (O_720,N_29950,N_28077);
and UO_721 (O_721,N_28547,N_29568);
or UO_722 (O_722,N_28911,N_28641);
xnor UO_723 (O_723,N_29264,N_29824);
xor UO_724 (O_724,N_29223,N_28398);
or UO_725 (O_725,N_29951,N_28960);
nor UO_726 (O_726,N_29947,N_29531);
and UO_727 (O_727,N_29414,N_29226);
xnor UO_728 (O_728,N_28448,N_28234);
nand UO_729 (O_729,N_28776,N_28825);
or UO_730 (O_730,N_29632,N_29064);
or UO_731 (O_731,N_28011,N_29846);
and UO_732 (O_732,N_28935,N_29941);
and UO_733 (O_733,N_28442,N_28385);
and UO_734 (O_734,N_28462,N_29411);
and UO_735 (O_735,N_28870,N_28671);
nand UO_736 (O_736,N_28636,N_28184);
nor UO_737 (O_737,N_29115,N_28892);
xor UO_738 (O_738,N_29403,N_29684);
nor UO_739 (O_739,N_28251,N_29942);
xnor UO_740 (O_740,N_29938,N_29617);
and UO_741 (O_741,N_29806,N_28637);
nor UO_742 (O_742,N_28513,N_29678);
and UO_743 (O_743,N_29893,N_28241);
nand UO_744 (O_744,N_28753,N_28674);
xnor UO_745 (O_745,N_28918,N_28058);
and UO_746 (O_746,N_28319,N_28741);
nand UO_747 (O_747,N_29407,N_29590);
or UO_748 (O_748,N_28842,N_29640);
or UO_749 (O_749,N_29867,N_28455);
xnor UO_750 (O_750,N_28128,N_29127);
or UO_751 (O_751,N_29366,N_29987);
and UO_752 (O_752,N_29636,N_29025);
xor UO_753 (O_753,N_28928,N_28136);
and UO_754 (O_754,N_29876,N_29359);
nand UO_755 (O_755,N_28532,N_28744);
nand UO_756 (O_756,N_28515,N_29200);
or UO_757 (O_757,N_29667,N_29373);
and UO_758 (O_758,N_29438,N_28997);
or UO_759 (O_759,N_28995,N_29752);
or UO_760 (O_760,N_28341,N_28066);
nand UO_761 (O_761,N_28394,N_28804);
and UO_762 (O_762,N_29247,N_29552);
and UO_763 (O_763,N_28956,N_29028);
xor UO_764 (O_764,N_28733,N_29330);
and UO_765 (O_765,N_29868,N_28572);
xnor UO_766 (O_766,N_28212,N_28070);
nand UO_767 (O_767,N_29066,N_29462);
or UO_768 (O_768,N_28687,N_29795);
nor UO_769 (O_769,N_28556,N_29467);
nand UO_770 (O_770,N_29211,N_28655);
and UO_771 (O_771,N_29747,N_28373);
nand UO_772 (O_772,N_29030,N_29479);
nor UO_773 (O_773,N_29902,N_28662);
and UO_774 (O_774,N_29355,N_28289);
and UO_775 (O_775,N_28881,N_29528);
or UO_776 (O_776,N_29404,N_28223);
nand UO_777 (O_777,N_28561,N_28001);
xnor UO_778 (O_778,N_29592,N_28485);
xor UO_779 (O_779,N_29263,N_28665);
or UO_780 (O_780,N_28800,N_29605);
xnor UO_781 (O_781,N_28503,N_29723);
and UO_782 (O_782,N_28725,N_29628);
nor UO_783 (O_783,N_29275,N_28566);
nor UO_784 (O_784,N_28933,N_28265);
xor UO_785 (O_785,N_29914,N_28284);
or UO_786 (O_786,N_28333,N_29187);
or UO_787 (O_787,N_29174,N_28165);
and UO_788 (O_788,N_29402,N_28426);
and UO_789 (O_789,N_28437,N_29185);
or UO_790 (O_790,N_29750,N_28272);
and UO_791 (O_791,N_28774,N_29655);
nor UO_792 (O_792,N_29798,N_28698);
nor UO_793 (O_793,N_29347,N_29977);
xnor UO_794 (O_794,N_28079,N_29885);
and UO_795 (O_795,N_28619,N_29936);
nand UO_796 (O_796,N_29544,N_28290);
xor UO_797 (O_797,N_29325,N_29943);
and UO_798 (O_798,N_28359,N_28847);
and UO_799 (O_799,N_28060,N_29743);
nor UO_800 (O_800,N_29616,N_28369);
nor UO_801 (O_801,N_29289,N_28059);
nand UO_802 (O_802,N_28827,N_28683);
or UO_803 (O_803,N_28303,N_29796);
and UO_804 (O_804,N_29837,N_28530);
and UO_805 (O_805,N_29847,N_29230);
or UO_806 (O_806,N_28452,N_28884);
nor UO_807 (O_807,N_29759,N_29555);
nor UO_808 (O_808,N_28672,N_28538);
xor UO_809 (O_809,N_29046,N_29308);
xor UO_810 (O_810,N_28338,N_29488);
nor UO_811 (O_811,N_29217,N_29825);
nand UO_812 (O_812,N_29714,N_28551);
nand UO_813 (O_813,N_28014,N_29900);
nor UO_814 (O_814,N_28856,N_29349);
xnor UO_815 (O_815,N_29178,N_28473);
and UO_816 (O_816,N_28602,N_28936);
nand UO_817 (O_817,N_28601,N_29788);
nor UO_818 (O_818,N_29671,N_29114);
or UO_819 (O_819,N_28638,N_29326);
or UO_820 (O_820,N_28522,N_28921);
xor UO_821 (O_821,N_28392,N_29078);
nor UO_822 (O_822,N_29986,N_29010);
or UO_823 (O_823,N_28049,N_28324);
or UO_824 (O_824,N_28647,N_29532);
or UO_825 (O_825,N_28216,N_29794);
xnor UO_826 (O_826,N_29310,N_28478);
nand UO_827 (O_827,N_28298,N_28910);
xnor UO_828 (O_828,N_29451,N_28280);
nor UO_829 (O_829,N_28258,N_29491);
nand UO_830 (O_830,N_28695,N_28730);
nand UO_831 (O_831,N_28391,N_29253);
and UO_832 (O_832,N_28195,N_28435);
xor UO_833 (O_833,N_28146,N_29144);
nor UO_834 (O_834,N_29970,N_29155);
or UO_835 (O_835,N_28846,N_28180);
xor UO_836 (O_836,N_29483,N_29427);
or UO_837 (O_837,N_29169,N_29043);
nor UO_838 (O_838,N_29396,N_28135);
or UO_839 (O_839,N_29008,N_29866);
and UO_840 (O_840,N_28786,N_29913);
and UO_841 (O_841,N_28629,N_28578);
nand UO_842 (O_842,N_29583,N_28854);
nor UO_843 (O_843,N_29306,N_29199);
and UO_844 (O_844,N_29541,N_28388);
nand UO_845 (O_845,N_29006,N_29702);
or UO_846 (O_846,N_29312,N_29618);
nand UO_847 (O_847,N_28081,N_29206);
nor UO_848 (O_848,N_29872,N_28242);
xnor UO_849 (O_849,N_29431,N_29686);
nand UO_850 (O_850,N_29232,N_28975);
or UO_851 (O_851,N_28358,N_29695);
and UO_852 (O_852,N_29229,N_28063);
nand UO_853 (O_853,N_28382,N_28355);
nor UO_854 (O_854,N_29742,N_28447);
xor UO_855 (O_855,N_28214,N_29487);
xor UO_856 (O_856,N_29455,N_29852);
nand UO_857 (O_857,N_29254,N_28622);
or UO_858 (O_858,N_29270,N_29013);
and UO_859 (O_859,N_29422,N_29812);
xor UO_860 (O_860,N_28734,N_29915);
xnor UO_861 (O_861,N_29305,N_29944);
and UO_862 (O_862,N_28717,N_29052);
and UO_863 (O_863,N_28138,N_29160);
or UO_864 (O_864,N_29344,N_28430);
xnor UO_865 (O_865,N_29865,N_28545);
xor UO_866 (O_866,N_28952,N_28652);
and UO_867 (O_867,N_29303,N_29945);
nor UO_868 (O_868,N_29134,N_28693);
nor UO_869 (O_869,N_28464,N_28950);
nand UO_870 (O_870,N_28984,N_28167);
nand UO_871 (O_871,N_28493,N_28616);
nand UO_872 (O_872,N_28365,N_28117);
and UO_873 (O_873,N_29175,N_29120);
xnor UO_874 (O_874,N_29880,N_29661);
nand UO_875 (O_875,N_28790,N_29390);
nor UO_876 (O_876,N_29245,N_28957);
nand UO_877 (O_877,N_29047,N_28915);
xnor UO_878 (O_878,N_28291,N_28998);
nand UO_879 (O_879,N_29638,N_29829);
nand UO_880 (O_880,N_28843,N_29510);
and UO_881 (O_881,N_28413,N_28152);
and UO_882 (O_882,N_28492,N_28393);
or UO_883 (O_883,N_29917,N_28477);
nand UO_884 (O_884,N_29388,N_29949);
nor UO_885 (O_885,N_28160,N_28959);
or UO_886 (O_886,N_28748,N_28829);
xnor UO_887 (O_887,N_28544,N_28335);
nand UO_888 (O_888,N_28837,N_28191);
xor UO_889 (O_889,N_28461,N_28107);
or UO_890 (O_890,N_28056,N_28599);
or UO_891 (O_891,N_28308,N_28848);
and UO_892 (O_892,N_29049,N_29503);
and UO_893 (O_893,N_28022,N_28030);
xnor UO_894 (O_894,N_28118,N_28673);
nor UO_895 (O_895,N_28113,N_29193);
nand UO_896 (O_896,N_28322,N_29138);
nor UO_897 (O_897,N_28472,N_28010);
nor UO_898 (O_898,N_29507,N_29581);
or UO_899 (O_899,N_29119,N_29776);
or UO_900 (O_900,N_29447,N_29591);
and UO_901 (O_901,N_29485,N_29456);
and UO_902 (O_902,N_29576,N_29087);
and UO_903 (O_903,N_29498,N_29724);
nor UO_904 (O_904,N_28235,N_28974);
and UO_905 (O_905,N_28418,N_28882);
and UO_906 (O_906,N_29218,N_29693);
and UO_907 (O_907,N_29061,N_28033);
and UO_908 (O_908,N_29007,N_28831);
xnor UO_909 (O_909,N_29781,N_28891);
and UO_910 (O_910,N_28116,N_28866);
xnor UO_911 (O_911,N_28168,N_28887);
and UO_912 (O_912,N_28127,N_28451);
xor UO_913 (O_913,N_29718,N_29656);
nand UO_914 (O_914,N_28035,N_29870);
nor UO_915 (O_915,N_29840,N_28484);
or UO_916 (O_916,N_28531,N_29588);
and UO_917 (O_917,N_29716,N_29198);
or UO_918 (O_918,N_29709,N_28953);
nand UO_919 (O_919,N_29808,N_29292);
nor UO_920 (O_920,N_28404,N_28684);
and UO_921 (O_921,N_29219,N_29801);
and UO_922 (O_922,N_28343,N_28230);
nor UO_923 (O_923,N_28821,N_28119);
nor UO_924 (O_924,N_28440,N_29271);
or UO_925 (O_925,N_28591,N_29725);
and UO_926 (O_926,N_29570,N_28849);
and UO_927 (O_927,N_28032,N_29843);
nand UO_928 (O_928,N_28810,N_28042);
xor UO_929 (O_929,N_28249,N_28292);
xnor UO_930 (O_930,N_29021,N_29898);
nand UO_931 (O_931,N_28177,N_29933);
and UO_932 (O_932,N_28182,N_29463);
or UO_933 (O_933,N_28312,N_28844);
nand UO_934 (O_934,N_29850,N_29346);
xor UO_935 (O_935,N_28381,N_29731);
nor UO_936 (O_936,N_28583,N_28862);
and UO_937 (O_937,N_29449,N_28446);
nor UO_938 (O_938,N_29336,N_28917);
nand UO_939 (O_939,N_28092,N_28963);
xor UO_940 (O_940,N_28486,N_28211);
or UO_941 (O_941,N_29113,N_29118);
nor UO_942 (O_942,N_28630,N_29248);
nor UO_943 (O_943,N_29448,N_28299);
xor UO_944 (O_944,N_28170,N_28221);
nand UO_945 (O_945,N_28557,N_29929);
nor UO_946 (O_946,N_29269,N_29222);
nand UO_947 (O_947,N_29612,N_28158);
nor UO_948 (O_948,N_28094,N_29991);
nor UO_949 (O_949,N_28454,N_29545);
nor UO_950 (O_950,N_29842,N_28021);
nor UO_951 (O_951,N_28737,N_29765);
or UO_952 (O_952,N_29141,N_29983);
and UO_953 (O_953,N_29317,N_29090);
and UO_954 (O_954,N_29019,N_28178);
nand UO_955 (O_955,N_29124,N_29536);
nand UO_956 (O_956,N_28702,N_29514);
or UO_957 (O_957,N_28386,N_28137);
nand UO_958 (O_958,N_29440,N_29869);
nand UO_959 (O_959,N_29381,N_28775);
xnor UO_960 (O_960,N_29088,N_29251);
xnor UO_961 (O_961,N_28434,N_29677);
or UO_962 (O_962,N_28508,N_29154);
nor UO_963 (O_963,N_29653,N_28302);
and UO_964 (O_964,N_29954,N_29803);
and UO_965 (O_965,N_29523,N_29897);
or UO_966 (O_966,N_29673,N_29055);
xor UO_967 (O_967,N_28653,N_28232);
nor UO_968 (O_968,N_28764,N_29994);
xor UO_969 (O_969,N_28841,N_29080);
nor UO_970 (O_970,N_29873,N_29643);
xor UO_971 (O_971,N_28595,N_28489);
or UO_972 (O_972,N_28620,N_29550);
nor UO_973 (O_973,N_29128,N_29874);
or UO_974 (O_974,N_29658,N_29358);
and UO_975 (O_975,N_29201,N_29800);
nand UO_976 (O_976,N_28618,N_28986);
and UO_977 (O_977,N_28678,N_28932);
nor UO_978 (O_978,N_28570,N_29371);
and UO_979 (O_979,N_29170,N_29474);
nor UO_980 (O_980,N_28240,N_28500);
nand UO_981 (O_981,N_28179,N_28109);
and UO_982 (O_982,N_29362,N_28577);
and UO_983 (O_983,N_28985,N_29026);
and UO_984 (O_984,N_29126,N_28939);
nand UO_985 (O_985,N_29664,N_28224);
nor UO_986 (O_986,N_28276,N_29246);
and UO_987 (O_987,N_28859,N_29554);
and UO_988 (O_988,N_28271,N_28976);
or UO_989 (O_989,N_28621,N_28226);
and UO_990 (O_990,N_28438,N_29109);
nand UO_991 (O_991,N_29250,N_29511);
or UO_992 (O_992,N_28668,N_28902);
nand UO_993 (O_993,N_29471,N_28316);
nand UO_994 (O_994,N_29888,N_28159);
xor UO_995 (O_995,N_28368,N_29538);
or UO_996 (O_996,N_28509,N_29669);
or UO_997 (O_997,N_28834,N_28054);
or UO_998 (O_998,N_28267,N_28648);
or UO_999 (O_999,N_28105,N_29645);
or UO_1000 (O_1000,N_29626,N_28559);
xnor UO_1001 (O_1001,N_29317,N_28823);
xor UO_1002 (O_1002,N_28474,N_29452);
nor UO_1003 (O_1003,N_28991,N_28634);
and UO_1004 (O_1004,N_28085,N_29987);
and UO_1005 (O_1005,N_29879,N_28460);
xnor UO_1006 (O_1006,N_28470,N_28825);
nand UO_1007 (O_1007,N_28786,N_29455);
and UO_1008 (O_1008,N_29775,N_29334);
and UO_1009 (O_1009,N_28415,N_28180);
or UO_1010 (O_1010,N_29066,N_28094);
or UO_1011 (O_1011,N_28274,N_29836);
and UO_1012 (O_1012,N_29510,N_28285);
xnor UO_1013 (O_1013,N_29064,N_28671);
nand UO_1014 (O_1014,N_28787,N_28333);
xor UO_1015 (O_1015,N_28345,N_28772);
xor UO_1016 (O_1016,N_28570,N_28555);
nand UO_1017 (O_1017,N_28982,N_28049);
nand UO_1018 (O_1018,N_28213,N_29361);
and UO_1019 (O_1019,N_29449,N_28378);
or UO_1020 (O_1020,N_29766,N_29678);
or UO_1021 (O_1021,N_29576,N_28417);
or UO_1022 (O_1022,N_29882,N_29104);
xnor UO_1023 (O_1023,N_28348,N_29587);
nand UO_1024 (O_1024,N_28642,N_29296);
nand UO_1025 (O_1025,N_29916,N_28354);
nor UO_1026 (O_1026,N_29509,N_29540);
nand UO_1027 (O_1027,N_28515,N_29528);
or UO_1028 (O_1028,N_29949,N_28412);
and UO_1029 (O_1029,N_29632,N_29584);
xor UO_1030 (O_1030,N_29932,N_29751);
and UO_1031 (O_1031,N_29002,N_28298);
or UO_1032 (O_1032,N_28495,N_29155);
nor UO_1033 (O_1033,N_28968,N_29098);
and UO_1034 (O_1034,N_29701,N_29944);
nand UO_1035 (O_1035,N_28978,N_28056);
and UO_1036 (O_1036,N_29170,N_29793);
nand UO_1037 (O_1037,N_28592,N_28630);
xnor UO_1038 (O_1038,N_29903,N_29241);
and UO_1039 (O_1039,N_28631,N_29886);
or UO_1040 (O_1040,N_28944,N_28022);
nor UO_1041 (O_1041,N_29431,N_28902);
nor UO_1042 (O_1042,N_28354,N_28352);
nand UO_1043 (O_1043,N_29623,N_28070);
nor UO_1044 (O_1044,N_28876,N_29401);
and UO_1045 (O_1045,N_29925,N_29897);
xor UO_1046 (O_1046,N_29730,N_29640);
nand UO_1047 (O_1047,N_28898,N_29486);
and UO_1048 (O_1048,N_29962,N_29586);
nor UO_1049 (O_1049,N_28413,N_28700);
nand UO_1050 (O_1050,N_28042,N_28722);
and UO_1051 (O_1051,N_29187,N_28460);
xnor UO_1052 (O_1052,N_28976,N_29234);
nand UO_1053 (O_1053,N_28102,N_28517);
and UO_1054 (O_1054,N_29144,N_29641);
and UO_1055 (O_1055,N_28646,N_28959);
nand UO_1056 (O_1056,N_29712,N_28351);
xor UO_1057 (O_1057,N_29198,N_29896);
or UO_1058 (O_1058,N_28786,N_29814);
nand UO_1059 (O_1059,N_29206,N_28428);
and UO_1060 (O_1060,N_28042,N_29532);
or UO_1061 (O_1061,N_29354,N_29004);
xor UO_1062 (O_1062,N_28609,N_28051);
nand UO_1063 (O_1063,N_29701,N_28555);
or UO_1064 (O_1064,N_28127,N_28737);
nor UO_1065 (O_1065,N_28793,N_29574);
nor UO_1066 (O_1066,N_28852,N_28017);
nand UO_1067 (O_1067,N_28652,N_29658);
and UO_1068 (O_1068,N_28744,N_29960);
nor UO_1069 (O_1069,N_29303,N_29848);
and UO_1070 (O_1070,N_29503,N_29495);
xnor UO_1071 (O_1071,N_28174,N_28682);
nand UO_1072 (O_1072,N_28601,N_29820);
or UO_1073 (O_1073,N_28864,N_28645);
or UO_1074 (O_1074,N_28320,N_28371);
xor UO_1075 (O_1075,N_28402,N_28279);
nor UO_1076 (O_1076,N_29587,N_29724);
nor UO_1077 (O_1077,N_28937,N_29986);
nand UO_1078 (O_1078,N_28187,N_28023);
or UO_1079 (O_1079,N_29599,N_28150);
nor UO_1080 (O_1080,N_29726,N_29829);
xnor UO_1081 (O_1081,N_29322,N_29835);
and UO_1082 (O_1082,N_29332,N_28446);
and UO_1083 (O_1083,N_29937,N_28386);
and UO_1084 (O_1084,N_28092,N_28334);
and UO_1085 (O_1085,N_28867,N_28044);
nor UO_1086 (O_1086,N_29241,N_29822);
and UO_1087 (O_1087,N_28015,N_29250);
nor UO_1088 (O_1088,N_29116,N_29038);
nor UO_1089 (O_1089,N_29167,N_28229);
nand UO_1090 (O_1090,N_29363,N_29208);
or UO_1091 (O_1091,N_29153,N_29885);
or UO_1092 (O_1092,N_28393,N_29751);
xor UO_1093 (O_1093,N_29098,N_29742);
and UO_1094 (O_1094,N_28152,N_28731);
and UO_1095 (O_1095,N_29816,N_29269);
and UO_1096 (O_1096,N_28793,N_29982);
and UO_1097 (O_1097,N_29352,N_28950);
nand UO_1098 (O_1098,N_28221,N_28871);
nand UO_1099 (O_1099,N_28654,N_28385);
and UO_1100 (O_1100,N_29336,N_28299);
nand UO_1101 (O_1101,N_29170,N_28363);
or UO_1102 (O_1102,N_28606,N_28361);
nor UO_1103 (O_1103,N_28793,N_29493);
nor UO_1104 (O_1104,N_29929,N_28359);
xor UO_1105 (O_1105,N_29722,N_28927);
nor UO_1106 (O_1106,N_29111,N_29554);
and UO_1107 (O_1107,N_29529,N_28402);
or UO_1108 (O_1108,N_28304,N_29389);
or UO_1109 (O_1109,N_28584,N_29554);
or UO_1110 (O_1110,N_29189,N_28755);
xnor UO_1111 (O_1111,N_28142,N_28517);
xnor UO_1112 (O_1112,N_29896,N_28281);
and UO_1113 (O_1113,N_29988,N_29833);
or UO_1114 (O_1114,N_28859,N_29984);
or UO_1115 (O_1115,N_28142,N_29183);
nor UO_1116 (O_1116,N_28391,N_28982);
nor UO_1117 (O_1117,N_28534,N_29390);
or UO_1118 (O_1118,N_29628,N_28855);
xor UO_1119 (O_1119,N_29923,N_28892);
or UO_1120 (O_1120,N_28978,N_29821);
and UO_1121 (O_1121,N_28389,N_29345);
or UO_1122 (O_1122,N_28162,N_29137);
and UO_1123 (O_1123,N_29894,N_28484);
xnor UO_1124 (O_1124,N_28324,N_28740);
nor UO_1125 (O_1125,N_28505,N_29731);
and UO_1126 (O_1126,N_28055,N_28724);
nor UO_1127 (O_1127,N_29406,N_28673);
xor UO_1128 (O_1128,N_28364,N_29036);
nand UO_1129 (O_1129,N_28556,N_29753);
xor UO_1130 (O_1130,N_28422,N_28655);
xnor UO_1131 (O_1131,N_28879,N_28298);
nand UO_1132 (O_1132,N_29406,N_28082);
nand UO_1133 (O_1133,N_29205,N_29281);
and UO_1134 (O_1134,N_29296,N_29065);
or UO_1135 (O_1135,N_29288,N_29043);
xor UO_1136 (O_1136,N_28927,N_28081);
or UO_1137 (O_1137,N_29044,N_28723);
nor UO_1138 (O_1138,N_28179,N_29088);
nand UO_1139 (O_1139,N_29171,N_28293);
xnor UO_1140 (O_1140,N_28141,N_29653);
nor UO_1141 (O_1141,N_29312,N_28612);
nand UO_1142 (O_1142,N_29639,N_28958);
and UO_1143 (O_1143,N_28157,N_28055);
and UO_1144 (O_1144,N_28588,N_28010);
or UO_1145 (O_1145,N_28986,N_28728);
nor UO_1146 (O_1146,N_28942,N_28391);
nand UO_1147 (O_1147,N_28445,N_29754);
xor UO_1148 (O_1148,N_29520,N_29270);
nor UO_1149 (O_1149,N_28027,N_28044);
nand UO_1150 (O_1150,N_29610,N_28848);
or UO_1151 (O_1151,N_29580,N_29113);
and UO_1152 (O_1152,N_28657,N_29009);
xor UO_1153 (O_1153,N_29209,N_29637);
and UO_1154 (O_1154,N_28023,N_29722);
or UO_1155 (O_1155,N_28462,N_29573);
and UO_1156 (O_1156,N_29365,N_28895);
nand UO_1157 (O_1157,N_28591,N_29289);
xor UO_1158 (O_1158,N_29893,N_29304);
or UO_1159 (O_1159,N_28240,N_28771);
nor UO_1160 (O_1160,N_28696,N_28217);
and UO_1161 (O_1161,N_29900,N_29016);
nor UO_1162 (O_1162,N_29388,N_28870);
nor UO_1163 (O_1163,N_28312,N_29756);
and UO_1164 (O_1164,N_28844,N_28592);
and UO_1165 (O_1165,N_29040,N_28620);
xnor UO_1166 (O_1166,N_29762,N_29555);
xnor UO_1167 (O_1167,N_29713,N_29980);
nor UO_1168 (O_1168,N_29935,N_28652);
nor UO_1169 (O_1169,N_28316,N_29742);
nand UO_1170 (O_1170,N_28614,N_29011);
nor UO_1171 (O_1171,N_29293,N_28672);
nand UO_1172 (O_1172,N_29241,N_29239);
or UO_1173 (O_1173,N_28365,N_28579);
nand UO_1174 (O_1174,N_28465,N_28162);
xnor UO_1175 (O_1175,N_28589,N_29798);
nor UO_1176 (O_1176,N_28959,N_29997);
and UO_1177 (O_1177,N_28152,N_29711);
xor UO_1178 (O_1178,N_29648,N_29268);
and UO_1179 (O_1179,N_28786,N_28114);
nor UO_1180 (O_1180,N_28568,N_29940);
and UO_1181 (O_1181,N_28353,N_29442);
or UO_1182 (O_1182,N_29957,N_28306);
and UO_1183 (O_1183,N_28885,N_28970);
nand UO_1184 (O_1184,N_28561,N_29068);
nor UO_1185 (O_1185,N_28157,N_29550);
or UO_1186 (O_1186,N_29267,N_29839);
and UO_1187 (O_1187,N_28622,N_29887);
or UO_1188 (O_1188,N_29767,N_29323);
nor UO_1189 (O_1189,N_28868,N_28470);
nand UO_1190 (O_1190,N_28740,N_29622);
or UO_1191 (O_1191,N_28777,N_28017);
or UO_1192 (O_1192,N_28013,N_28852);
nor UO_1193 (O_1193,N_29890,N_29119);
nor UO_1194 (O_1194,N_29036,N_29354);
nand UO_1195 (O_1195,N_29419,N_28313);
and UO_1196 (O_1196,N_28053,N_28765);
nand UO_1197 (O_1197,N_29555,N_28979);
nand UO_1198 (O_1198,N_28612,N_28042);
nand UO_1199 (O_1199,N_29905,N_29655);
and UO_1200 (O_1200,N_28803,N_29276);
xor UO_1201 (O_1201,N_28517,N_29120);
or UO_1202 (O_1202,N_28053,N_28151);
or UO_1203 (O_1203,N_29948,N_28808);
nand UO_1204 (O_1204,N_28657,N_28586);
nand UO_1205 (O_1205,N_29441,N_29440);
nand UO_1206 (O_1206,N_29920,N_29769);
nor UO_1207 (O_1207,N_29302,N_29106);
and UO_1208 (O_1208,N_28468,N_29974);
and UO_1209 (O_1209,N_29511,N_28063);
nand UO_1210 (O_1210,N_29971,N_29794);
nand UO_1211 (O_1211,N_28018,N_29894);
nor UO_1212 (O_1212,N_28381,N_28862);
or UO_1213 (O_1213,N_29905,N_29638);
xor UO_1214 (O_1214,N_29826,N_28030);
nand UO_1215 (O_1215,N_28810,N_28837);
xnor UO_1216 (O_1216,N_29282,N_29408);
xnor UO_1217 (O_1217,N_29126,N_28413);
nor UO_1218 (O_1218,N_29968,N_28998);
xnor UO_1219 (O_1219,N_28487,N_29196);
and UO_1220 (O_1220,N_29215,N_29589);
nand UO_1221 (O_1221,N_28862,N_28289);
nand UO_1222 (O_1222,N_29106,N_29088);
nor UO_1223 (O_1223,N_28915,N_28036);
and UO_1224 (O_1224,N_28312,N_28879);
xor UO_1225 (O_1225,N_29882,N_29238);
or UO_1226 (O_1226,N_28673,N_29088);
nand UO_1227 (O_1227,N_28655,N_28411);
xor UO_1228 (O_1228,N_28693,N_28259);
or UO_1229 (O_1229,N_29081,N_28912);
xnor UO_1230 (O_1230,N_28371,N_28446);
or UO_1231 (O_1231,N_29632,N_28034);
and UO_1232 (O_1232,N_29815,N_29782);
or UO_1233 (O_1233,N_29495,N_28861);
nand UO_1234 (O_1234,N_28119,N_29860);
nand UO_1235 (O_1235,N_29629,N_28311);
and UO_1236 (O_1236,N_29162,N_29742);
or UO_1237 (O_1237,N_28116,N_28165);
and UO_1238 (O_1238,N_28824,N_28818);
nand UO_1239 (O_1239,N_29065,N_29192);
nor UO_1240 (O_1240,N_28600,N_28857);
nor UO_1241 (O_1241,N_29597,N_28354);
xor UO_1242 (O_1242,N_29272,N_29691);
and UO_1243 (O_1243,N_29631,N_28611);
or UO_1244 (O_1244,N_29670,N_28532);
nor UO_1245 (O_1245,N_28232,N_28743);
nand UO_1246 (O_1246,N_28523,N_28530);
nor UO_1247 (O_1247,N_28556,N_29628);
xnor UO_1248 (O_1248,N_28483,N_28288);
nand UO_1249 (O_1249,N_28491,N_29411);
and UO_1250 (O_1250,N_29536,N_28592);
nand UO_1251 (O_1251,N_28221,N_28386);
or UO_1252 (O_1252,N_28737,N_28425);
or UO_1253 (O_1253,N_28665,N_28011);
xnor UO_1254 (O_1254,N_29120,N_28872);
nand UO_1255 (O_1255,N_28852,N_28079);
or UO_1256 (O_1256,N_28085,N_29768);
or UO_1257 (O_1257,N_28122,N_28954);
nor UO_1258 (O_1258,N_28806,N_29761);
or UO_1259 (O_1259,N_29272,N_28398);
nor UO_1260 (O_1260,N_29697,N_29734);
nand UO_1261 (O_1261,N_29672,N_28552);
nor UO_1262 (O_1262,N_28939,N_28113);
nand UO_1263 (O_1263,N_29028,N_28906);
nand UO_1264 (O_1264,N_29185,N_29452);
or UO_1265 (O_1265,N_29194,N_29864);
xor UO_1266 (O_1266,N_28542,N_28196);
nand UO_1267 (O_1267,N_28183,N_29753);
xnor UO_1268 (O_1268,N_28843,N_29154);
nand UO_1269 (O_1269,N_28347,N_28741);
xnor UO_1270 (O_1270,N_29238,N_28199);
nand UO_1271 (O_1271,N_28865,N_28223);
xor UO_1272 (O_1272,N_28004,N_28579);
xnor UO_1273 (O_1273,N_28746,N_28230);
or UO_1274 (O_1274,N_29178,N_28020);
or UO_1275 (O_1275,N_29856,N_28471);
or UO_1276 (O_1276,N_28323,N_29805);
nand UO_1277 (O_1277,N_28683,N_29342);
or UO_1278 (O_1278,N_28966,N_29016);
and UO_1279 (O_1279,N_28830,N_28841);
xor UO_1280 (O_1280,N_29484,N_29937);
or UO_1281 (O_1281,N_29692,N_28826);
nor UO_1282 (O_1282,N_28488,N_28497);
or UO_1283 (O_1283,N_28669,N_29606);
nand UO_1284 (O_1284,N_29291,N_29284);
xor UO_1285 (O_1285,N_29383,N_28980);
and UO_1286 (O_1286,N_28518,N_28126);
nand UO_1287 (O_1287,N_29089,N_28350);
xor UO_1288 (O_1288,N_28673,N_28841);
and UO_1289 (O_1289,N_29209,N_28419);
or UO_1290 (O_1290,N_29210,N_29207);
xor UO_1291 (O_1291,N_28733,N_29605);
nand UO_1292 (O_1292,N_28666,N_29542);
nor UO_1293 (O_1293,N_28365,N_28544);
nand UO_1294 (O_1294,N_28622,N_29329);
or UO_1295 (O_1295,N_29954,N_29840);
xor UO_1296 (O_1296,N_28373,N_28463);
nand UO_1297 (O_1297,N_28079,N_28577);
nand UO_1298 (O_1298,N_28737,N_29863);
and UO_1299 (O_1299,N_28106,N_29909);
nand UO_1300 (O_1300,N_28154,N_29134);
nor UO_1301 (O_1301,N_28820,N_28561);
or UO_1302 (O_1302,N_29813,N_29152);
nand UO_1303 (O_1303,N_29390,N_28256);
xor UO_1304 (O_1304,N_29321,N_29437);
and UO_1305 (O_1305,N_29703,N_29145);
nor UO_1306 (O_1306,N_29843,N_28763);
and UO_1307 (O_1307,N_29669,N_28522);
nor UO_1308 (O_1308,N_28552,N_28954);
nor UO_1309 (O_1309,N_29576,N_28156);
nand UO_1310 (O_1310,N_29680,N_29195);
nand UO_1311 (O_1311,N_28857,N_28565);
xnor UO_1312 (O_1312,N_28636,N_28347);
xnor UO_1313 (O_1313,N_29348,N_29627);
and UO_1314 (O_1314,N_29648,N_28191);
or UO_1315 (O_1315,N_28838,N_28441);
or UO_1316 (O_1316,N_28184,N_28112);
nor UO_1317 (O_1317,N_28134,N_29849);
xor UO_1318 (O_1318,N_28145,N_28911);
nor UO_1319 (O_1319,N_29314,N_29749);
or UO_1320 (O_1320,N_29087,N_28209);
and UO_1321 (O_1321,N_29470,N_28659);
nand UO_1322 (O_1322,N_28563,N_29494);
nor UO_1323 (O_1323,N_29910,N_29169);
xnor UO_1324 (O_1324,N_29426,N_29106);
nand UO_1325 (O_1325,N_28187,N_29942);
and UO_1326 (O_1326,N_28049,N_28370);
nor UO_1327 (O_1327,N_29072,N_29137);
nor UO_1328 (O_1328,N_29989,N_28660);
or UO_1329 (O_1329,N_28254,N_29080);
nand UO_1330 (O_1330,N_29792,N_28810);
nor UO_1331 (O_1331,N_29974,N_28380);
xor UO_1332 (O_1332,N_29689,N_28138);
nand UO_1333 (O_1333,N_28466,N_28135);
nand UO_1334 (O_1334,N_29020,N_29972);
nand UO_1335 (O_1335,N_28237,N_29759);
or UO_1336 (O_1336,N_28063,N_28310);
or UO_1337 (O_1337,N_28474,N_28313);
or UO_1338 (O_1338,N_28583,N_29257);
nor UO_1339 (O_1339,N_28848,N_28614);
nor UO_1340 (O_1340,N_29560,N_28259);
xnor UO_1341 (O_1341,N_29355,N_28559);
xor UO_1342 (O_1342,N_29296,N_28831);
xor UO_1343 (O_1343,N_29332,N_28116);
nor UO_1344 (O_1344,N_29015,N_28898);
and UO_1345 (O_1345,N_29366,N_29676);
xnor UO_1346 (O_1346,N_28872,N_28796);
nor UO_1347 (O_1347,N_29004,N_29323);
or UO_1348 (O_1348,N_28404,N_29998);
xnor UO_1349 (O_1349,N_28547,N_29510);
nand UO_1350 (O_1350,N_29185,N_28038);
nand UO_1351 (O_1351,N_29680,N_28076);
or UO_1352 (O_1352,N_29959,N_29913);
or UO_1353 (O_1353,N_28137,N_29366);
nor UO_1354 (O_1354,N_29696,N_29999);
or UO_1355 (O_1355,N_29092,N_29349);
nor UO_1356 (O_1356,N_29054,N_28514);
and UO_1357 (O_1357,N_29816,N_28314);
nor UO_1358 (O_1358,N_28318,N_28081);
and UO_1359 (O_1359,N_28376,N_29656);
nor UO_1360 (O_1360,N_28760,N_28949);
and UO_1361 (O_1361,N_29738,N_29114);
or UO_1362 (O_1362,N_28873,N_29261);
or UO_1363 (O_1363,N_29110,N_29480);
and UO_1364 (O_1364,N_28957,N_29139);
and UO_1365 (O_1365,N_29696,N_29140);
nor UO_1366 (O_1366,N_28848,N_29318);
nand UO_1367 (O_1367,N_29066,N_29303);
xor UO_1368 (O_1368,N_29387,N_28715);
or UO_1369 (O_1369,N_29024,N_28010);
or UO_1370 (O_1370,N_28351,N_28618);
xor UO_1371 (O_1371,N_28708,N_28590);
and UO_1372 (O_1372,N_29462,N_29829);
xor UO_1373 (O_1373,N_28765,N_28177);
or UO_1374 (O_1374,N_28590,N_29859);
nand UO_1375 (O_1375,N_28689,N_29679);
or UO_1376 (O_1376,N_29120,N_29389);
and UO_1377 (O_1377,N_28323,N_29997);
or UO_1378 (O_1378,N_29348,N_28076);
xnor UO_1379 (O_1379,N_29019,N_29323);
or UO_1380 (O_1380,N_28905,N_29491);
nand UO_1381 (O_1381,N_28031,N_28464);
and UO_1382 (O_1382,N_28482,N_29191);
and UO_1383 (O_1383,N_29566,N_28472);
xnor UO_1384 (O_1384,N_28997,N_28470);
xnor UO_1385 (O_1385,N_28202,N_28413);
xor UO_1386 (O_1386,N_28970,N_29245);
nor UO_1387 (O_1387,N_28904,N_29207);
or UO_1388 (O_1388,N_28779,N_28190);
and UO_1389 (O_1389,N_29576,N_29045);
or UO_1390 (O_1390,N_28957,N_29203);
nand UO_1391 (O_1391,N_29255,N_29563);
nor UO_1392 (O_1392,N_29614,N_29519);
nand UO_1393 (O_1393,N_28390,N_29321);
nand UO_1394 (O_1394,N_29626,N_29594);
xor UO_1395 (O_1395,N_29461,N_29606);
or UO_1396 (O_1396,N_28986,N_28650);
or UO_1397 (O_1397,N_29195,N_28882);
nor UO_1398 (O_1398,N_29432,N_29259);
nand UO_1399 (O_1399,N_28985,N_29965);
and UO_1400 (O_1400,N_28559,N_28762);
nand UO_1401 (O_1401,N_28312,N_28478);
or UO_1402 (O_1402,N_28334,N_29820);
xor UO_1403 (O_1403,N_29651,N_28911);
nor UO_1404 (O_1404,N_28887,N_28248);
xor UO_1405 (O_1405,N_29005,N_29500);
xnor UO_1406 (O_1406,N_29809,N_28384);
and UO_1407 (O_1407,N_28281,N_29566);
nor UO_1408 (O_1408,N_28140,N_29672);
nor UO_1409 (O_1409,N_28083,N_28474);
nand UO_1410 (O_1410,N_29737,N_28309);
nand UO_1411 (O_1411,N_28112,N_28487);
and UO_1412 (O_1412,N_28644,N_29045);
xnor UO_1413 (O_1413,N_28070,N_28181);
and UO_1414 (O_1414,N_29084,N_29398);
and UO_1415 (O_1415,N_29690,N_28023);
and UO_1416 (O_1416,N_28343,N_28384);
or UO_1417 (O_1417,N_29709,N_29907);
xnor UO_1418 (O_1418,N_29830,N_29105);
or UO_1419 (O_1419,N_29377,N_29848);
nor UO_1420 (O_1420,N_28411,N_28745);
nand UO_1421 (O_1421,N_29451,N_29650);
nor UO_1422 (O_1422,N_29913,N_29575);
nand UO_1423 (O_1423,N_28917,N_29824);
xor UO_1424 (O_1424,N_29225,N_29084);
or UO_1425 (O_1425,N_29262,N_28110);
xor UO_1426 (O_1426,N_28012,N_28963);
nand UO_1427 (O_1427,N_28137,N_28110);
and UO_1428 (O_1428,N_29194,N_29766);
and UO_1429 (O_1429,N_28039,N_28742);
and UO_1430 (O_1430,N_28689,N_28680);
nand UO_1431 (O_1431,N_28430,N_29038);
or UO_1432 (O_1432,N_29381,N_29837);
xnor UO_1433 (O_1433,N_28060,N_28553);
nor UO_1434 (O_1434,N_29292,N_29642);
nor UO_1435 (O_1435,N_29247,N_28750);
and UO_1436 (O_1436,N_29177,N_28686);
nand UO_1437 (O_1437,N_29742,N_29040);
nor UO_1438 (O_1438,N_28362,N_28221);
xor UO_1439 (O_1439,N_28251,N_29795);
and UO_1440 (O_1440,N_28194,N_28365);
and UO_1441 (O_1441,N_29518,N_29660);
xnor UO_1442 (O_1442,N_29693,N_28140);
or UO_1443 (O_1443,N_28824,N_29538);
nor UO_1444 (O_1444,N_29119,N_28062);
and UO_1445 (O_1445,N_29593,N_29610);
nor UO_1446 (O_1446,N_29317,N_28256);
xnor UO_1447 (O_1447,N_29727,N_28108);
xnor UO_1448 (O_1448,N_28390,N_28884);
nor UO_1449 (O_1449,N_28863,N_28835);
nand UO_1450 (O_1450,N_28979,N_28869);
and UO_1451 (O_1451,N_28113,N_28604);
xnor UO_1452 (O_1452,N_29059,N_28203);
and UO_1453 (O_1453,N_28136,N_28756);
xnor UO_1454 (O_1454,N_29887,N_29428);
and UO_1455 (O_1455,N_29940,N_29124);
xnor UO_1456 (O_1456,N_29170,N_29554);
nand UO_1457 (O_1457,N_28216,N_28825);
or UO_1458 (O_1458,N_28804,N_29345);
nor UO_1459 (O_1459,N_29012,N_29797);
or UO_1460 (O_1460,N_29612,N_29108);
or UO_1461 (O_1461,N_28206,N_28272);
nor UO_1462 (O_1462,N_29179,N_28120);
or UO_1463 (O_1463,N_29867,N_28348);
and UO_1464 (O_1464,N_28382,N_28256);
and UO_1465 (O_1465,N_28156,N_29175);
nor UO_1466 (O_1466,N_28215,N_28248);
or UO_1467 (O_1467,N_29914,N_29892);
nor UO_1468 (O_1468,N_28945,N_28376);
and UO_1469 (O_1469,N_28135,N_28372);
and UO_1470 (O_1470,N_29584,N_28865);
nor UO_1471 (O_1471,N_28183,N_29313);
nand UO_1472 (O_1472,N_29939,N_29223);
nor UO_1473 (O_1473,N_29269,N_29500);
xnor UO_1474 (O_1474,N_28033,N_28189);
or UO_1475 (O_1475,N_29208,N_29736);
nand UO_1476 (O_1476,N_28917,N_28598);
nor UO_1477 (O_1477,N_29831,N_28809);
nor UO_1478 (O_1478,N_29249,N_28811);
and UO_1479 (O_1479,N_28763,N_29649);
and UO_1480 (O_1480,N_29791,N_29799);
nor UO_1481 (O_1481,N_28768,N_29266);
or UO_1482 (O_1482,N_28055,N_28674);
or UO_1483 (O_1483,N_28808,N_29343);
nand UO_1484 (O_1484,N_29444,N_29071);
and UO_1485 (O_1485,N_29483,N_29841);
xnor UO_1486 (O_1486,N_28840,N_28622);
or UO_1487 (O_1487,N_28952,N_28316);
nor UO_1488 (O_1488,N_28420,N_29569);
or UO_1489 (O_1489,N_28324,N_28092);
nor UO_1490 (O_1490,N_29986,N_28319);
nor UO_1491 (O_1491,N_29296,N_28351);
and UO_1492 (O_1492,N_29828,N_28819);
xor UO_1493 (O_1493,N_29720,N_29788);
xnor UO_1494 (O_1494,N_28877,N_28004);
or UO_1495 (O_1495,N_29284,N_28009);
nor UO_1496 (O_1496,N_28726,N_28099);
xor UO_1497 (O_1497,N_29916,N_29104);
or UO_1498 (O_1498,N_28129,N_29471);
nand UO_1499 (O_1499,N_29424,N_29351);
nand UO_1500 (O_1500,N_29531,N_28592);
nand UO_1501 (O_1501,N_28800,N_29582);
or UO_1502 (O_1502,N_29011,N_28831);
nand UO_1503 (O_1503,N_28367,N_29758);
or UO_1504 (O_1504,N_29262,N_28614);
and UO_1505 (O_1505,N_28392,N_29978);
and UO_1506 (O_1506,N_29958,N_29518);
nand UO_1507 (O_1507,N_29050,N_28311);
xnor UO_1508 (O_1508,N_29857,N_28029);
nand UO_1509 (O_1509,N_29170,N_28900);
nand UO_1510 (O_1510,N_29018,N_29437);
nand UO_1511 (O_1511,N_28470,N_29617);
nor UO_1512 (O_1512,N_29059,N_28972);
xor UO_1513 (O_1513,N_28063,N_29922);
nor UO_1514 (O_1514,N_28163,N_29189);
and UO_1515 (O_1515,N_28229,N_28510);
nor UO_1516 (O_1516,N_29959,N_28057);
and UO_1517 (O_1517,N_29674,N_28093);
and UO_1518 (O_1518,N_29226,N_28762);
nor UO_1519 (O_1519,N_28730,N_29582);
and UO_1520 (O_1520,N_28658,N_29940);
and UO_1521 (O_1521,N_29362,N_28879);
and UO_1522 (O_1522,N_29118,N_28680);
xnor UO_1523 (O_1523,N_28614,N_28202);
and UO_1524 (O_1524,N_29487,N_29461);
and UO_1525 (O_1525,N_29764,N_28013);
nor UO_1526 (O_1526,N_29617,N_29778);
nor UO_1527 (O_1527,N_29321,N_29443);
xor UO_1528 (O_1528,N_28661,N_28629);
xnor UO_1529 (O_1529,N_28396,N_29859);
nand UO_1530 (O_1530,N_29335,N_29629);
nand UO_1531 (O_1531,N_28359,N_28137);
or UO_1532 (O_1532,N_28940,N_28722);
nand UO_1533 (O_1533,N_29603,N_29300);
nor UO_1534 (O_1534,N_28099,N_28970);
nand UO_1535 (O_1535,N_29229,N_28008);
or UO_1536 (O_1536,N_28494,N_28344);
nor UO_1537 (O_1537,N_28221,N_28638);
xnor UO_1538 (O_1538,N_29492,N_29940);
nor UO_1539 (O_1539,N_29864,N_28786);
nor UO_1540 (O_1540,N_28001,N_28070);
nor UO_1541 (O_1541,N_28653,N_29765);
and UO_1542 (O_1542,N_29956,N_29812);
or UO_1543 (O_1543,N_29437,N_28508);
nor UO_1544 (O_1544,N_28273,N_28572);
xnor UO_1545 (O_1545,N_29529,N_29037);
nor UO_1546 (O_1546,N_29649,N_29580);
nor UO_1547 (O_1547,N_28520,N_29423);
and UO_1548 (O_1548,N_29468,N_29315);
nor UO_1549 (O_1549,N_29204,N_29155);
or UO_1550 (O_1550,N_29756,N_28767);
nor UO_1551 (O_1551,N_28504,N_28809);
and UO_1552 (O_1552,N_29682,N_28043);
nor UO_1553 (O_1553,N_29480,N_29500);
nand UO_1554 (O_1554,N_28407,N_28207);
nand UO_1555 (O_1555,N_28681,N_29840);
xnor UO_1556 (O_1556,N_29053,N_28691);
xnor UO_1557 (O_1557,N_29643,N_28749);
and UO_1558 (O_1558,N_29007,N_29403);
nand UO_1559 (O_1559,N_29059,N_29865);
xnor UO_1560 (O_1560,N_28413,N_29555);
and UO_1561 (O_1561,N_29270,N_29887);
or UO_1562 (O_1562,N_28165,N_29094);
nor UO_1563 (O_1563,N_28582,N_28725);
and UO_1564 (O_1564,N_29328,N_28825);
and UO_1565 (O_1565,N_29276,N_28437);
or UO_1566 (O_1566,N_28868,N_28226);
nor UO_1567 (O_1567,N_28184,N_29298);
or UO_1568 (O_1568,N_29892,N_28395);
xnor UO_1569 (O_1569,N_28435,N_28128);
or UO_1570 (O_1570,N_28368,N_28293);
nand UO_1571 (O_1571,N_28363,N_28817);
xor UO_1572 (O_1572,N_28839,N_28840);
or UO_1573 (O_1573,N_29476,N_28326);
or UO_1574 (O_1574,N_29735,N_29016);
or UO_1575 (O_1575,N_28785,N_28002);
xnor UO_1576 (O_1576,N_28231,N_29524);
nand UO_1577 (O_1577,N_29118,N_28472);
and UO_1578 (O_1578,N_29218,N_28175);
xor UO_1579 (O_1579,N_29492,N_29545);
or UO_1580 (O_1580,N_28761,N_29025);
and UO_1581 (O_1581,N_28402,N_29472);
nor UO_1582 (O_1582,N_29657,N_28783);
or UO_1583 (O_1583,N_28390,N_28127);
and UO_1584 (O_1584,N_29935,N_28319);
nor UO_1585 (O_1585,N_28561,N_28925);
nand UO_1586 (O_1586,N_29725,N_28611);
and UO_1587 (O_1587,N_29461,N_28246);
xor UO_1588 (O_1588,N_28759,N_29698);
or UO_1589 (O_1589,N_28825,N_28460);
nor UO_1590 (O_1590,N_29326,N_29887);
or UO_1591 (O_1591,N_28206,N_29014);
nor UO_1592 (O_1592,N_29024,N_28293);
and UO_1593 (O_1593,N_28519,N_29716);
nand UO_1594 (O_1594,N_28648,N_29591);
xnor UO_1595 (O_1595,N_28380,N_29530);
nand UO_1596 (O_1596,N_28541,N_28108);
nor UO_1597 (O_1597,N_29379,N_29904);
xnor UO_1598 (O_1598,N_29835,N_29069);
xnor UO_1599 (O_1599,N_29928,N_29741);
xor UO_1600 (O_1600,N_28699,N_28922);
or UO_1601 (O_1601,N_28525,N_28066);
or UO_1602 (O_1602,N_28614,N_28997);
and UO_1603 (O_1603,N_28326,N_28133);
nor UO_1604 (O_1604,N_29373,N_29690);
nand UO_1605 (O_1605,N_28761,N_29798);
or UO_1606 (O_1606,N_29643,N_29903);
nand UO_1607 (O_1607,N_29057,N_29196);
nor UO_1608 (O_1608,N_29584,N_28205);
or UO_1609 (O_1609,N_28074,N_28187);
nand UO_1610 (O_1610,N_28132,N_29673);
nand UO_1611 (O_1611,N_28901,N_28395);
or UO_1612 (O_1612,N_28741,N_29011);
nor UO_1613 (O_1613,N_29598,N_28397);
nor UO_1614 (O_1614,N_29529,N_28022);
nand UO_1615 (O_1615,N_29038,N_28768);
nand UO_1616 (O_1616,N_29623,N_29679);
and UO_1617 (O_1617,N_29987,N_29161);
nor UO_1618 (O_1618,N_29443,N_28990);
and UO_1619 (O_1619,N_28454,N_29760);
and UO_1620 (O_1620,N_29888,N_28219);
xnor UO_1621 (O_1621,N_29483,N_29869);
and UO_1622 (O_1622,N_28920,N_29025);
nor UO_1623 (O_1623,N_29586,N_28760);
nand UO_1624 (O_1624,N_28919,N_29928);
or UO_1625 (O_1625,N_28778,N_28358);
nor UO_1626 (O_1626,N_29687,N_28818);
xnor UO_1627 (O_1627,N_29847,N_29896);
nand UO_1628 (O_1628,N_29479,N_28916);
or UO_1629 (O_1629,N_29489,N_28396);
xnor UO_1630 (O_1630,N_28190,N_29497);
nor UO_1631 (O_1631,N_29586,N_28954);
and UO_1632 (O_1632,N_28183,N_28067);
nor UO_1633 (O_1633,N_29322,N_29264);
xnor UO_1634 (O_1634,N_28288,N_29313);
xor UO_1635 (O_1635,N_29485,N_28669);
and UO_1636 (O_1636,N_29336,N_29616);
nand UO_1637 (O_1637,N_28657,N_29564);
and UO_1638 (O_1638,N_29303,N_28180);
nand UO_1639 (O_1639,N_28591,N_29495);
nand UO_1640 (O_1640,N_28807,N_29442);
or UO_1641 (O_1641,N_29002,N_29947);
and UO_1642 (O_1642,N_28831,N_28648);
xnor UO_1643 (O_1643,N_29057,N_28750);
nand UO_1644 (O_1644,N_29998,N_29326);
xor UO_1645 (O_1645,N_29832,N_29332);
and UO_1646 (O_1646,N_28781,N_29753);
nand UO_1647 (O_1647,N_29782,N_28323);
nor UO_1648 (O_1648,N_28782,N_29385);
and UO_1649 (O_1649,N_29254,N_28136);
nor UO_1650 (O_1650,N_29246,N_29773);
nand UO_1651 (O_1651,N_28195,N_29934);
and UO_1652 (O_1652,N_28490,N_29892);
and UO_1653 (O_1653,N_29880,N_28388);
and UO_1654 (O_1654,N_29537,N_28781);
nand UO_1655 (O_1655,N_29119,N_29399);
and UO_1656 (O_1656,N_28054,N_29868);
or UO_1657 (O_1657,N_28889,N_29408);
or UO_1658 (O_1658,N_29627,N_28307);
or UO_1659 (O_1659,N_28614,N_29889);
nor UO_1660 (O_1660,N_28970,N_28890);
xor UO_1661 (O_1661,N_28505,N_29371);
xor UO_1662 (O_1662,N_28605,N_28613);
nand UO_1663 (O_1663,N_28232,N_29769);
or UO_1664 (O_1664,N_29387,N_29981);
xor UO_1665 (O_1665,N_29059,N_29890);
nand UO_1666 (O_1666,N_29711,N_28804);
and UO_1667 (O_1667,N_29304,N_28603);
nor UO_1668 (O_1668,N_28444,N_28074);
and UO_1669 (O_1669,N_28283,N_29789);
nand UO_1670 (O_1670,N_29814,N_28884);
or UO_1671 (O_1671,N_29775,N_29227);
nand UO_1672 (O_1672,N_28164,N_29186);
xor UO_1673 (O_1673,N_28044,N_28905);
and UO_1674 (O_1674,N_29365,N_29137);
xnor UO_1675 (O_1675,N_29106,N_29527);
nor UO_1676 (O_1676,N_28393,N_28833);
nor UO_1677 (O_1677,N_29345,N_28504);
nand UO_1678 (O_1678,N_28794,N_29715);
nand UO_1679 (O_1679,N_29891,N_29452);
xor UO_1680 (O_1680,N_29388,N_28488);
nor UO_1681 (O_1681,N_28210,N_29481);
xor UO_1682 (O_1682,N_28411,N_29784);
xor UO_1683 (O_1683,N_29974,N_29204);
nor UO_1684 (O_1684,N_29221,N_29773);
and UO_1685 (O_1685,N_29866,N_29777);
nor UO_1686 (O_1686,N_29231,N_29766);
or UO_1687 (O_1687,N_28848,N_28200);
nand UO_1688 (O_1688,N_29052,N_29431);
or UO_1689 (O_1689,N_29415,N_28579);
nand UO_1690 (O_1690,N_28808,N_29595);
or UO_1691 (O_1691,N_29474,N_29263);
nor UO_1692 (O_1692,N_28182,N_29002);
or UO_1693 (O_1693,N_28431,N_28474);
nand UO_1694 (O_1694,N_29706,N_28214);
or UO_1695 (O_1695,N_29985,N_28756);
nand UO_1696 (O_1696,N_29375,N_28998);
or UO_1697 (O_1697,N_28772,N_29216);
xnor UO_1698 (O_1698,N_28881,N_29002);
and UO_1699 (O_1699,N_29717,N_29275);
or UO_1700 (O_1700,N_29018,N_28244);
nand UO_1701 (O_1701,N_28248,N_28551);
nand UO_1702 (O_1702,N_28642,N_29541);
or UO_1703 (O_1703,N_28326,N_28342);
and UO_1704 (O_1704,N_28097,N_28114);
xor UO_1705 (O_1705,N_29019,N_29732);
and UO_1706 (O_1706,N_29218,N_28703);
or UO_1707 (O_1707,N_29279,N_29553);
and UO_1708 (O_1708,N_29375,N_28663);
xor UO_1709 (O_1709,N_29053,N_29444);
nand UO_1710 (O_1710,N_28393,N_29931);
xnor UO_1711 (O_1711,N_28436,N_29767);
and UO_1712 (O_1712,N_28032,N_29457);
nor UO_1713 (O_1713,N_29714,N_29300);
or UO_1714 (O_1714,N_28730,N_28645);
nor UO_1715 (O_1715,N_28911,N_29044);
and UO_1716 (O_1716,N_29548,N_28787);
and UO_1717 (O_1717,N_29390,N_28718);
nand UO_1718 (O_1718,N_28702,N_28407);
or UO_1719 (O_1719,N_29654,N_29163);
or UO_1720 (O_1720,N_28338,N_29554);
nor UO_1721 (O_1721,N_29249,N_29646);
xnor UO_1722 (O_1722,N_28030,N_29634);
nand UO_1723 (O_1723,N_29692,N_28122);
or UO_1724 (O_1724,N_29319,N_28328);
xnor UO_1725 (O_1725,N_29890,N_29674);
nor UO_1726 (O_1726,N_29332,N_28175);
nand UO_1727 (O_1727,N_29514,N_29267);
nand UO_1728 (O_1728,N_28778,N_28000);
nand UO_1729 (O_1729,N_28085,N_28489);
xor UO_1730 (O_1730,N_29956,N_29552);
nor UO_1731 (O_1731,N_28022,N_29838);
xor UO_1732 (O_1732,N_28446,N_28983);
and UO_1733 (O_1733,N_28172,N_29758);
nand UO_1734 (O_1734,N_29600,N_29006);
xor UO_1735 (O_1735,N_28099,N_28194);
nor UO_1736 (O_1736,N_29284,N_28076);
xnor UO_1737 (O_1737,N_28172,N_28673);
nor UO_1738 (O_1738,N_28963,N_29678);
nand UO_1739 (O_1739,N_29912,N_29818);
or UO_1740 (O_1740,N_29116,N_29588);
nand UO_1741 (O_1741,N_28006,N_29344);
xnor UO_1742 (O_1742,N_28488,N_29792);
and UO_1743 (O_1743,N_29064,N_29198);
nand UO_1744 (O_1744,N_28800,N_29544);
xor UO_1745 (O_1745,N_29419,N_29561);
nor UO_1746 (O_1746,N_29264,N_29654);
nand UO_1747 (O_1747,N_29432,N_28946);
nand UO_1748 (O_1748,N_28059,N_29788);
nor UO_1749 (O_1749,N_28268,N_28822);
nor UO_1750 (O_1750,N_29831,N_28475);
or UO_1751 (O_1751,N_28471,N_29050);
nand UO_1752 (O_1752,N_28590,N_29250);
nor UO_1753 (O_1753,N_28199,N_28630);
and UO_1754 (O_1754,N_29496,N_28166);
xor UO_1755 (O_1755,N_28959,N_28421);
nand UO_1756 (O_1756,N_28588,N_29890);
xnor UO_1757 (O_1757,N_28515,N_29071);
or UO_1758 (O_1758,N_28938,N_28104);
and UO_1759 (O_1759,N_28975,N_28324);
xnor UO_1760 (O_1760,N_28824,N_29773);
and UO_1761 (O_1761,N_28056,N_29269);
nand UO_1762 (O_1762,N_29145,N_29012);
or UO_1763 (O_1763,N_29863,N_28446);
nor UO_1764 (O_1764,N_29640,N_28111);
and UO_1765 (O_1765,N_29379,N_28822);
xnor UO_1766 (O_1766,N_29261,N_29282);
xor UO_1767 (O_1767,N_28126,N_29420);
xor UO_1768 (O_1768,N_28007,N_28974);
or UO_1769 (O_1769,N_29399,N_29510);
nand UO_1770 (O_1770,N_28048,N_29419);
nand UO_1771 (O_1771,N_29997,N_28239);
or UO_1772 (O_1772,N_28913,N_28166);
nor UO_1773 (O_1773,N_29395,N_28633);
xnor UO_1774 (O_1774,N_28637,N_29223);
xor UO_1775 (O_1775,N_28934,N_29998);
nor UO_1776 (O_1776,N_29087,N_29200);
nand UO_1777 (O_1777,N_29830,N_29349);
and UO_1778 (O_1778,N_29590,N_29720);
or UO_1779 (O_1779,N_29844,N_28673);
and UO_1780 (O_1780,N_29003,N_29270);
nor UO_1781 (O_1781,N_29965,N_28286);
nor UO_1782 (O_1782,N_29026,N_28045);
nor UO_1783 (O_1783,N_28142,N_29804);
nor UO_1784 (O_1784,N_29246,N_28073);
nand UO_1785 (O_1785,N_29548,N_28056);
nand UO_1786 (O_1786,N_29539,N_29758);
xnor UO_1787 (O_1787,N_28286,N_28644);
nand UO_1788 (O_1788,N_29997,N_29431);
nor UO_1789 (O_1789,N_28573,N_29049);
or UO_1790 (O_1790,N_29720,N_28550);
xor UO_1791 (O_1791,N_28628,N_28715);
or UO_1792 (O_1792,N_28666,N_28041);
or UO_1793 (O_1793,N_29213,N_28330);
xor UO_1794 (O_1794,N_28993,N_28614);
and UO_1795 (O_1795,N_28045,N_29377);
or UO_1796 (O_1796,N_28703,N_29725);
nand UO_1797 (O_1797,N_28582,N_29592);
or UO_1798 (O_1798,N_29254,N_28323);
or UO_1799 (O_1799,N_29735,N_29444);
nand UO_1800 (O_1800,N_29635,N_28367);
nand UO_1801 (O_1801,N_29069,N_29059);
xor UO_1802 (O_1802,N_28405,N_28332);
nor UO_1803 (O_1803,N_29195,N_28903);
or UO_1804 (O_1804,N_29392,N_28852);
nand UO_1805 (O_1805,N_28651,N_28269);
xor UO_1806 (O_1806,N_28360,N_29498);
nor UO_1807 (O_1807,N_29632,N_28947);
and UO_1808 (O_1808,N_28607,N_28097);
nand UO_1809 (O_1809,N_29979,N_29308);
nor UO_1810 (O_1810,N_29136,N_28340);
nor UO_1811 (O_1811,N_28888,N_28931);
nand UO_1812 (O_1812,N_28551,N_29978);
xnor UO_1813 (O_1813,N_28708,N_28368);
nand UO_1814 (O_1814,N_28509,N_29079);
and UO_1815 (O_1815,N_28451,N_28721);
and UO_1816 (O_1816,N_28134,N_29281);
and UO_1817 (O_1817,N_28885,N_29274);
xor UO_1818 (O_1818,N_29577,N_28581);
or UO_1819 (O_1819,N_29081,N_28790);
nor UO_1820 (O_1820,N_29534,N_29225);
nor UO_1821 (O_1821,N_29264,N_29700);
nor UO_1822 (O_1822,N_28124,N_29320);
nand UO_1823 (O_1823,N_28388,N_28262);
or UO_1824 (O_1824,N_28344,N_28789);
nand UO_1825 (O_1825,N_28922,N_28917);
or UO_1826 (O_1826,N_29368,N_28125);
or UO_1827 (O_1827,N_29654,N_28687);
nor UO_1828 (O_1828,N_29456,N_28990);
nor UO_1829 (O_1829,N_29335,N_28517);
nand UO_1830 (O_1830,N_28922,N_29065);
or UO_1831 (O_1831,N_28277,N_29523);
xor UO_1832 (O_1832,N_28372,N_29847);
or UO_1833 (O_1833,N_29987,N_29095);
xnor UO_1834 (O_1834,N_28712,N_29134);
xnor UO_1835 (O_1835,N_29113,N_28288);
nor UO_1836 (O_1836,N_29169,N_28853);
nand UO_1837 (O_1837,N_28518,N_28336);
nor UO_1838 (O_1838,N_29762,N_29870);
nor UO_1839 (O_1839,N_29742,N_28891);
or UO_1840 (O_1840,N_29817,N_28874);
or UO_1841 (O_1841,N_29015,N_28079);
nand UO_1842 (O_1842,N_28997,N_28521);
or UO_1843 (O_1843,N_29145,N_28985);
or UO_1844 (O_1844,N_29103,N_29640);
xor UO_1845 (O_1845,N_28934,N_28697);
or UO_1846 (O_1846,N_28404,N_28282);
nand UO_1847 (O_1847,N_29042,N_28632);
xnor UO_1848 (O_1848,N_28811,N_28948);
or UO_1849 (O_1849,N_29961,N_29348);
or UO_1850 (O_1850,N_29536,N_28442);
and UO_1851 (O_1851,N_28856,N_29764);
nor UO_1852 (O_1852,N_28799,N_29047);
xnor UO_1853 (O_1853,N_28412,N_28596);
and UO_1854 (O_1854,N_28235,N_29603);
nor UO_1855 (O_1855,N_28302,N_28819);
and UO_1856 (O_1856,N_28924,N_28459);
nand UO_1857 (O_1857,N_28523,N_29184);
nand UO_1858 (O_1858,N_28514,N_28122);
xor UO_1859 (O_1859,N_29331,N_28464);
xor UO_1860 (O_1860,N_28949,N_28094);
and UO_1861 (O_1861,N_29460,N_29358);
xor UO_1862 (O_1862,N_29832,N_28587);
nor UO_1863 (O_1863,N_29880,N_29328);
nor UO_1864 (O_1864,N_28391,N_28374);
and UO_1865 (O_1865,N_28770,N_29708);
xnor UO_1866 (O_1866,N_28695,N_28338);
and UO_1867 (O_1867,N_29548,N_29605);
and UO_1868 (O_1868,N_29949,N_29307);
nor UO_1869 (O_1869,N_28995,N_28356);
nor UO_1870 (O_1870,N_29286,N_29742);
nor UO_1871 (O_1871,N_29181,N_29919);
or UO_1872 (O_1872,N_29092,N_29627);
or UO_1873 (O_1873,N_29181,N_28508);
or UO_1874 (O_1874,N_29655,N_29472);
nor UO_1875 (O_1875,N_29130,N_29224);
or UO_1876 (O_1876,N_28962,N_28916);
or UO_1877 (O_1877,N_28200,N_28024);
or UO_1878 (O_1878,N_28680,N_28036);
nor UO_1879 (O_1879,N_29953,N_29363);
or UO_1880 (O_1880,N_28849,N_28396);
and UO_1881 (O_1881,N_29295,N_28343);
and UO_1882 (O_1882,N_29012,N_28316);
and UO_1883 (O_1883,N_29557,N_28447);
or UO_1884 (O_1884,N_29973,N_28011);
nor UO_1885 (O_1885,N_29675,N_29757);
nor UO_1886 (O_1886,N_28527,N_28947);
and UO_1887 (O_1887,N_29190,N_28251);
nor UO_1888 (O_1888,N_28207,N_29753);
and UO_1889 (O_1889,N_28699,N_29578);
nand UO_1890 (O_1890,N_28687,N_28904);
and UO_1891 (O_1891,N_29799,N_29852);
nand UO_1892 (O_1892,N_29508,N_29687);
nor UO_1893 (O_1893,N_29154,N_28333);
xor UO_1894 (O_1894,N_29089,N_28222);
or UO_1895 (O_1895,N_28379,N_29805);
or UO_1896 (O_1896,N_28294,N_29569);
xnor UO_1897 (O_1897,N_28100,N_29783);
nor UO_1898 (O_1898,N_29151,N_28305);
and UO_1899 (O_1899,N_29090,N_29220);
nand UO_1900 (O_1900,N_28298,N_29908);
xor UO_1901 (O_1901,N_29048,N_29840);
nand UO_1902 (O_1902,N_28765,N_28261);
nor UO_1903 (O_1903,N_28975,N_29158);
nand UO_1904 (O_1904,N_28983,N_28508);
nor UO_1905 (O_1905,N_28667,N_29513);
nand UO_1906 (O_1906,N_28695,N_29755);
xor UO_1907 (O_1907,N_28828,N_28174);
and UO_1908 (O_1908,N_29096,N_29725);
xor UO_1909 (O_1909,N_28294,N_29737);
nor UO_1910 (O_1910,N_29227,N_29557);
nand UO_1911 (O_1911,N_28425,N_28650);
xor UO_1912 (O_1912,N_28624,N_29655);
nor UO_1913 (O_1913,N_28628,N_29323);
and UO_1914 (O_1914,N_28556,N_28620);
nor UO_1915 (O_1915,N_29255,N_29579);
nor UO_1916 (O_1916,N_29004,N_28786);
nand UO_1917 (O_1917,N_28036,N_28136);
and UO_1918 (O_1918,N_29425,N_29618);
nand UO_1919 (O_1919,N_29365,N_29155);
xnor UO_1920 (O_1920,N_28716,N_28723);
and UO_1921 (O_1921,N_28322,N_28935);
xnor UO_1922 (O_1922,N_29262,N_29212);
or UO_1923 (O_1923,N_29702,N_28211);
nor UO_1924 (O_1924,N_28651,N_29370);
nor UO_1925 (O_1925,N_28125,N_28663);
xnor UO_1926 (O_1926,N_29395,N_29834);
xor UO_1927 (O_1927,N_28360,N_29659);
xnor UO_1928 (O_1928,N_28790,N_29610);
xor UO_1929 (O_1929,N_28201,N_29587);
nor UO_1930 (O_1930,N_29352,N_28423);
or UO_1931 (O_1931,N_29352,N_29801);
nand UO_1932 (O_1932,N_28689,N_29747);
and UO_1933 (O_1933,N_28633,N_29375);
nand UO_1934 (O_1934,N_28296,N_29191);
xnor UO_1935 (O_1935,N_28507,N_28893);
or UO_1936 (O_1936,N_28615,N_29366);
nor UO_1937 (O_1937,N_29564,N_29260);
and UO_1938 (O_1938,N_29884,N_29340);
nor UO_1939 (O_1939,N_29351,N_28732);
and UO_1940 (O_1940,N_29675,N_28000);
nand UO_1941 (O_1941,N_29807,N_28571);
or UO_1942 (O_1942,N_28338,N_28226);
xnor UO_1943 (O_1943,N_28179,N_29423);
and UO_1944 (O_1944,N_29528,N_29775);
or UO_1945 (O_1945,N_29445,N_29564);
nand UO_1946 (O_1946,N_28778,N_28810);
xnor UO_1947 (O_1947,N_29173,N_28438);
nand UO_1948 (O_1948,N_28780,N_28302);
and UO_1949 (O_1949,N_28760,N_28810);
or UO_1950 (O_1950,N_28932,N_28994);
xnor UO_1951 (O_1951,N_29162,N_29308);
nor UO_1952 (O_1952,N_28146,N_28467);
xor UO_1953 (O_1953,N_28512,N_28610);
nand UO_1954 (O_1954,N_29500,N_29572);
and UO_1955 (O_1955,N_28853,N_28867);
xor UO_1956 (O_1956,N_28966,N_29838);
and UO_1957 (O_1957,N_29742,N_29696);
and UO_1958 (O_1958,N_28477,N_29725);
nand UO_1959 (O_1959,N_28155,N_29534);
xor UO_1960 (O_1960,N_29367,N_29018);
and UO_1961 (O_1961,N_29520,N_28530);
nand UO_1962 (O_1962,N_28182,N_28569);
and UO_1963 (O_1963,N_29779,N_29754);
and UO_1964 (O_1964,N_29604,N_28490);
or UO_1965 (O_1965,N_29401,N_28632);
xor UO_1966 (O_1966,N_29656,N_29081);
xor UO_1967 (O_1967,N_28483,N_28480);
xnor UO_1968 (O_1968,N_29553,N_28428);
xor UO_1969 (O_1969,N_29202,N_28479);
nand UO_1970 (O_1970,N_28936,N_29992);
nor UO_1971 (O_1971,N_28258,N_29088);
and UO_1972 (O_1972,N_28577,N_28882);
nand UO_1973 (O_1973,N_28789,N_29945);
or UO_1974 (O_1974,N_28538,N_28078);
xor UO_1975 (O_1975,N_28901,N_28917);
xor UO_1976 (O_1976,N_29956,N_28571);
xor UO_1977 (O_1977,N_28917,N_28100);
xor UO_1978 (O_1978,N_28349,N_28752);
or UO_1979 (O_1979,N_29103,N_28352);
or UO_1980 (O_1980,N_28822,N_28469);
nor UO_1981 (O_1981,N_29969,N_28193);
nand UO_1982 (O_1982,N_29240,N_28982);
nor UO_1983 (O_1983,N_29006,N_29671);
xor UO_1984 (O_1984,N_29055,N_29733);
and UO_1985 (O_1985,N_29678,N_28211);
xor UO_1986 (O_1986,N_28677,N_29333);
xor UO_1987 (O_1987,N_29603,N_28996);
nand UO_1988 (O_1988,N_28963,N_28851);
nand UO_1989 (O_1989,N_28788,N_29896);
nor UO_1990 (O_1990,N_28279,N_29028);
and UO_1991 (O_1991,N_28515,N_28781);
and UO_1992 (O_1992,N_28332,N_28763);
nor UO_1993 (O_1993,N_28737,N_29170);
nor UO_1994 (O_1994,N_29965,N_29376);
and UO_1995 (O_1995,N_28933,N_28663);
and UO_1996 (O_1996,N_28289,N_29604);
nand UO_1997 (O_1997,N_29662,N_29484);
nor UO_1998 (O_1998,N_28446,N_29964);
nor UO_1999 (O_1999,N_28328,N_28796);
and UO_2000 (O_2000,N_28372,N_28621);
nor UO_2001 (O_2001,N_28609,N_28141);
and UO_2002 (O_2002,N_29631,N_29769);
or UO_2003 (O_2003,N_28875,N_28097);
or UO_2004 (O_2004,N_29065,N_28371);
and UO_2005 (O_2005,N_29935,N_28257);
and UO_2006 (O_2006,N_29425,N_29080);
xnor UO_2007 (O_2007,N_28310,N_29652);
and UO_2008 (O_2008,N_29725,N_28219);
and UO_2009 (O_2009,N_28287,N_29161);
nor UO_2010 (O_2010,N_28999,N_28822);
or UO_2011 (O_2011,N_29406,N_28554);
nor UO_2012 (O_2012,N_29805,N_28953);
and UO_2013 (O_2013,N_28721,N_28354);
xnor UO_2014 (O_2014,N_28506,N_29515);
and UO_2015 (O_2015,N_29870,N_29673);
nand UO_2016 (O_2016,N_28557,N_29359);
and UO_2017 (O_2017,N_29688,N_29965);
nor UO_2018 (O_2018,N_28836,N_29777);
or UO_2019 (O_2019,N_29960,N_28746);
xnor UO_2020 (O_2020,N_29464,N_28818);
and UO_2021 (O_2021,N_28077,N_28939);
nor UO_2022 (O_2022,N_29359,N_29521);
nor UO_2023 (O_2023,N_28454,N_28273);
and UO_2024 (O_2024,N_28049,N_28586);
or UO_2025 (O_2025,N_29237,N_28760);
nor UO_2026 (O_2026,N_28296,N_28947);
and UO_2027 (O_2027,N_28273,N_29829);
nor UO_2028 (O_2028,N_29206,N_28361);
nor UO_2029 (O_2029,N_28790,N_28342);
nand UO_2030 (O_2030,N_29071,N_29109);
or UO_2031 (O_2031,N_28136,N_29120);
and UO_2032 (O_2032,N_28230,N_28506);
nand UO_2033 (O_2033,N_28096,N_29860);
nor UO_2034 (O_2034,N_28946,N_28491);
and UO_2035 (O_2035,N_29075,N_29220);
nor UO_2036 (O_2036,N_28699,N_29992);
nor UO_2037 (O_2037,N_28829,N_28097);
nor UO_2038 (O_2038,N_29012,N_29633);
or UO_2039 (O_2039,N_28188,N_28182);
xnor UO_2040 (O_2040,N_29738,N_29577);
xor UO_2041 (O_2041,N_28422,N_28090);
nor UO_2042 (O_2042,N_28092,N_28672);
and UO_2043 (O_2043,N_29147,N_28339);
nand UO_2044 (O_2044,N_28446,N_28460);
xnor UO_2045 (O_2045,N_29449,N_28043);
xor UO_2046 (O_2046,N_29809,N_29643);
nand UO_2047 (O_2047,N_29122,N_28101);
and UO_2048 (O_2048,N_28970,N_29788);
nand UO_2049 (O_2049,N_29890,N_29173);
nand UO_2050 (O_2050,N_29391,N_29812);
nor UO_2051 (O_2051,N_29731,N_28233);
nand UO_2052 (O_2052,N_29590,N_29908);
or UO_2053 (O_2053,N_29929,N_28501);
nor UO_2054 (O_2054,N_28496,N_28925);
nand UO_2055 (O_2055,N_28223,N_28227);
and UO_2056 (O_2056,N_28065,N_29375);
and UO_2057 (O_2057,N_28044,N_28541);
nor UO_2058 (O_2058,N_29790,N_29850);
nand UO_2059 (O_2059,N_28623,N_28179);
xor UO_2060 (O_2060,N_29261,N_28259);
nand UO_2061 (O_2061,N_28347,N_29297);
or UO_2062 (O_2062,N_28613,N_28522);
and UO_2063 (O_2063,N_29061,N_29075);
xnor UO_2064 (O_2064,N_28610,N_28880);
nor UO_2065 (O_2065,N_29873,N_28890);
xor UO_2066 (O_2066,N_29214,N_28735);
or UO_2067 (O_2067,N_29760,N_28917);
or UO_2068 (O_2068,N_28204,N_28021);
and UO_2069 (O_2069,N_29984,N_28970);
nor UO_2070 (O_2070,N_29505,N_29554);
nand UO_2071 (O_2071,N_28143,N_29072);
nand UO_2072 (O_2072,N_29679,N_28329);
xnor UO_2073 (O_2073,N_29985,N_29804);
and UO_2074 (O_2074,N_28034,N_29750);
xor UO_2075 (O_2075,N_29183,N_29350);
nor UO_2076 (O_2076,N_29167,N_28703);
or UO_2077 (O_2077,N_29208,N_28835);
nand UO_2078 (O_2078,N_29275,N_28273);
nand UO_2079 (O_2079,N_29722,N_29084);
nand UO_2080 (O_2080,N_28810,N_29831);
nor UO_2081 (O_2081,N_28913,N_29889);
nand UO_2082 (O_2082,N_28530,N_29845);
and UO_2083 (O_2083,N_29208,N_29963);
nand UO_2084 (O_2084,N_29090,N_28875);
nand UO_2085 (O_2085,N_29133,N_28187);
or UO_2086 (O_2086,N_28235,N_28333);
nor UO_2087 (O_2087,N_29213,N_28807);
xnor UO_2088 (O_2088,N_28756,N_28687);
xnor UO_2089 (O_2089,N_28306,N_29255);
nor UO_2090 (O_2090,N_29784,N_29041);
nor UO_2091 (O_2091,N_28882,N_29772);
and UO_2092 (O_2092,N_29900,N_29518);
nand UO_2093 (O_2093,N_29704,N_28353);
or UO_2094 (O_2094,N_28732,N_28229);
or UO_2095 (O_2095,N_29808,N_28398);
xnor UO_2096 (O_2096,N_28800,N_28376);
xnor UO_2097 (O_2097,N_28471,N_28932);
or UO_2098 (O_2098,N_28491,N_29750);
nor UO_2099 (O_2099,N_28855,N_29796);
and UO_2100 (O_2100,N_28179,N_28723);
nand UO_2101 (O_2101,N_29869,N_29173);
nand UO_2102 (O_2102,N_28967,N_29696);
xor UO_2103 (O_2103,N_29666,N_29781);
nand UO_2104 (O_2104,N_28270,N_29982);
or UO_2105 (O_2105,N_28611,N_29258);
or UO_2106 (O_2106,N_29553,N_28155);
xor UO_2107 (O_2107,N_29719,N_29813);
nor UO_2108 (O_2108,N_29679,N_29546);
and UO_2109 (O_2109,N_28336,N_28400);
nor UO_2110 (O_2110,N_29259,N_28952);
nand UO_2111 (O_2111,N_28202,N_29541);
nand UO_2112 (O_2112,N_28334,N_29572);
nand UO_2113 (O_2113,N_29949,N_28844);
xnor UO_2114 (O_2114,N_28499,N_28884);
xnor UO_2115 (O_2115,N_28781,N_28145);
nor UO_2116 (O_2116,N_28802,N_28933);
or UO_2117 (O_2117,N_28527,N_28789);
nand UO_2118 (O_2118,N_28035,N_29466);
and UO_2119 (O_2119,N_28918,N_29114);
nand UO_2120 (O_2120,N_29289,N_28759);
or UO_2121 (O_2121,N_29906,N_29933);
or UO_2122 (O_2122,N_29440,N_29406);
xnor UO_2123 (O_2123,N_28281,N_28904);
nor UO_2124 (O_2124,N_29910,N_28629);
and UO_2125 (O_2125,N_29488,N_29005);
or UO_2126 (O_2126,N_29230,N_28543);
and UO_2127 (O_2127,N_29825,N_29198);
nand UO_2128 (O_2128,N_29400,N_29675);
nand UO_2129 (O_2129,N_28849,N_28002);
and UO_2130 (O_2130,N_28643,N_28586);
or UO_2131 (O_2131,N_29927,N_29497);
nand UO_2132 (O_2132,N_29114,N_29485);
xor UO_2133 (O_2133,N_29496,N_28361);
or UO_2134 (O_2134,N_28384,N_28903);
and UO_2135 (O_2135,N_29048,N_29620);
or UO_2136 (O_2136,N_29449,N_29367);
and UO_2137 (O_2137,N_29227,N_28463);
nor UO_2138 (O_2138,N_28449,N_29888);
and UO_2139 (O_2139,N_29246,N_29306);
nor UO_2140 (O_2140,N_29707,N_29647);
xnor UO_2141 (O_2141,N_28485,N_29664);
or UO_2142 (O_2142,N_28028,N_28651);
nor UO_2143 (O_2143,N_28249,N_28610);
and UO_2144 (O_2144,N_28175,N_29800);
or UO_2145 (O_2145,N_29183,N_29444);
and UO_2146 (O_2146,N_29802,N_28485);
nand UO_2147 (O_2147,N_29853,N_28473);
and UO_2148 (O_2148,N_29143,N_29126);
or UO_2149 (O_2149,N_28987,N_29129);
nor UO_2150 (O_2150,N_28183,N_28584);
xnor UO_2151 (O_2151,N_29206,N_29681);
xnor UO_2152 (O_2152,N_29285,N_29276);
or UO_2153 (O_2153,N_28015,N_29124);
and UO_2154 (O_2154,N_28677,N_28839);
or UO_2155 (O_2155,N_28540,N_29543);
xor UO_2156 (O_2156,N_29680,N_28483);
xnor UO_2157 (O_2157,N_29056,N_29797);
xnor UO_2158 (O_2158,N_28234,N_28471);
xor UO_2159 (O_2159,N_28758,N_28095);
or UO_2160 (O_2160,N_28402,N_29332);
and UO_2161 (O_2161,N_28759,N_28850);
nand UO_2162 (O_2162,N_28807,N_28735);
and UO_2163 (O_2163,N_28296,N_29155);
nand UO_2164 (O_2164,N_29820,N_29493);
and UO_2165 (O_2165,N_29989,N_28057);
xnor UO_2166 (O_2166,N_28808,N_29624);
nand UO_2167 (O_2167,N_28117,N_28153);
or UO_2168 (O_2168,N_29587,N_29306);
xnor UO_2169 (O_2169,N_29204,N_28243);
and UO_2170 (O_2170,N_29384,N_29533);
and UO_2171 (O_2171,N_29977,N_28008);
xor UO_2172 (O_2172,N_28077,N_29526);
and UO_2173 (O_2173,N_28697,N_28155);
or UO_2174 (O_2174,N_29532,N_29195);
xor UO_2175 (O_2175,N_28462,N_29847);
or UO_2176 (O_2176,N_28478,N_28330);
and UO_2177 (O_2177,N_29547,N_29853);
nor UO_2178 (O_2178,N_28217,N_28177);
nand UO_2179 (O_2179,N_29676,N_29661);
nand UO_2180 (O_2180,N_28893,N_28051);
or UO_2181 (O_2181,N_29555,N_29398);
nand UO_2182 (O_2182,N_28381,N_29009);
xnor UO_2183 (O_2183,N_28229,N_28086);
nor UO_2184 (O_2184,N_29370,N_28763);
xnor UO_2185 (O_2185,N_29337,N_29558);
xor UO_2186 (O_2186,N_29415,N_28156);
nor UO_2187 (O_2187,N_28729,N_29724);
and UO_2188 (O_2188,N_28389,N_29439);
or UO_2189 (O_2189,N_28323,N_28374);
xor UO_2190 (O_2190,N_29300,N_28338);
and UO_2191 (O_2191,N_29158,N_28980);
and UO_2192 (O_2192,N_28351,N_28986);
xnor UO_2193 (O_2193,N_28520,N_28556);
nor UO_2194 (O_2194,N_29239,N_28130);
nor UO_2195 (O_2195,N_29046,N_28394);
or UO_2196 (O_2196,N_28094,N_29400);
nor UO_2197 (O_2197,N_29620,N_29380);
and UO_2198 (O_2198,N_29041,N_28936);
nand UO_2199 (O_2199,N_28585,N_28515);
nand UO_2200 (O_2200,N_28466,N_29680);
nor UO_2201 (O_2201,N_29176,N_29174);
or UO_2202 (O_2202,N_29148,N_28125);
nor UO_2203 (O_2203,N_28980,N_28060);
or UO_2204 (O_2204,N_29382,N_28586);
nand UO_2205 (O_2205,N_29421,N_29750);
or UO_2206 (O_2206,N_28042,N_29757);
or UO_2207 (O_2207,N_29000,N_28837);
or UO_2208 (O_2208,N_29892,N_28244);
and UO_2209 (O_2209,N_28268,N_28371);
xnor UO_2210 (O_2210,N_29319,N_29044);
and UO_2211 (O_2211,N_29362,N_28233);
nand UO_2212 (O_2212,N_28606,N_28352);
xor UO_2213 (O_2213,N_28181,N_29353);
and UO_2214 (O_2214,N_28380,N_28477);
or UO_2215 (O_2215,N_29766,N_28776);
or UO_2216 (O_2216,N_28182,N_29025);
or UO_2217 (O_2217,N_29703,N_28416);
and UO_2218 (O_2218,N_29931,N_28131);
nand UO_2219 (O_2219,N_28533,N_29714);
nor UO_2220 (O_2220,N_29158,N_28312);
nand UO_2221 (O_2221,N_28638,N_28630);
and UO_2222 (O_2222,N_28407,N_28518);
xor UO_2223 (O_2223,N_28391,N_28488);
xor UO_2224 (O_2224,N_29997,N_29411);
or UO_2225 (O_2225,N_29892,N_28392);
xor UO_2226 (O_2226,N_28828,N_29581);
or UO_2227 (O_2227,N_28868,N_28102);
nand UO_2228 (O_2228,N_28015,N_28234);
nand UO_2229 (O_2229,N_28353,N_29341);
or UO_2230 (O_2230,N_29198,N_28549);
nand UO_2231 (O_2231,N_29873,N_28539);
and UO_2232 (O_2232,N_29903,N_28780);
and UO_2233 (O_2233,N_28833,N_29688);
xor UO_2234 (O_2234,N_28849,N_28214);
nand UO_2235 (O_2235,N_29436,N_28750);
nand UO_2236 (O_2236,N_28818,N_28287);
nor UO_2237 (O_2237,N_28294,N_29164);
and UO_2238 (O_2238,N_28174,N_29561);
xnor UO_2239 (O_2239,N_29825,N_29157);
or UO_2240 (O_2240,N_28294,N_29832);
nor UO_2241 (O_2241,N_29632,N_28008);
and UO_2242 (O_2242,N_29597,N_29298);
or UO_2243 (O_2243,N_28265,N_29173);
and UO_2244 (O_2244,N_29326,N_28432);
or UO_2245 (O_2245,N_28636,N_29320);
nand UO_2246 (O_2246,N_29092,N_28355);
and UO_2247 (O_2247,N_28202,N_29432);
and UO_2248 (O_2248,N_28918,N_29357);
and UO_2249 (O_2249,N_28863,N_28544);
nor UO_2250 (O_2250,N_28595,N_29740);
xor UO_2251 (O_2251,N_29050,N_28281);
and UO_2252 (O_2252,N_28149,N_28550);
or UO_2253 (O_2253,N_29724,N_29074);
xor UO_2254 (O_2254,N_28234,N_28018);
or UO_2255 (O_2255,N_28288,N_28327);
nand UO_2256 (O_2256,N_28300,N_29237);
nor UO_2257 (O_2257,N_28025,N_29458);
nor UO_2258 (O_2258,N_28558,N_28117);
or UO_2259 (O_2259,N_28362,N_28733);
nor UO_2260 (O_2260,N_29471,N_28372);
nand UO_2261 (O_2261,N_29568,N_28391);
nor UO_2262 (O_2262,N_29715,N_28367);
and UO_2263 (O_2263,N_29980,N_29021);
nand UO_2264 (O_2264,N_28463,N_29424);
or UO_2265 (O_2265,N_29190,N_28339);
nand UO_2266 (O_2266,N_28853,N_28907);
xor UO_2267 (O_2267,N_29754,N_28657);
or UO_2268 (O_2268,N_29520,N_28248);
nand UO_2269 (O_2269,N_29998,N_28497);
nor UO_2270 (O_2270,N_29173,N_28859);
nor UO_2271 (O_2271,N_28743,N_29971);
nor UO_2272 (O_2272,N_28064,N_28377);
or UO_2273 (O_2273,N_29064,N_29454);
or UO_2274 (O_2274,N_28244,N_29857);
xor UO_2275 (O_2275,N_29836,N_28710);
xnor UO_2276 (O_2276,N_29274,N_29701);
nor UO_2277 (O_2277,N_29212,N_28682);
and UO_2278 (O_2278,N_28489,N_28488);
or UO_2279 (O_2279,N_29099,N_29093);
xnor UO_2280 (O_2280,N_29770,N_29005);
xor UO_2281 (O_2281,N_29667,N_28737);
xnor UO_2282 (O_2282,N_28091,N_28487);
nand UO_2283 (O_2283,N_28021,N_28920);
or UO_2284 (O_2284,N_29339,N_28692);
xor UO_2285 (O_2285,N_28995,N_29785);
xnor UO_2286 (O_2286,N_28969,N_28541);
nand UO_2287 (O_2287,N_28106,N_28402);
and UO_2288 (O_2288,N_29714,N_29193);
or UO_2289 (O_2289,N_28991,N_28369);
nor UO_2290 (O_2290,N_28283,N_29952);
xor UO_2291 (O_2291,N_29862,N_29038);
nor UO_2292 (O_2292,N_28593,N_28103);
nor UO_2293 (O_2293,N_29258,N_29016);
nand UO_2294 (O_2294,N_28950,N_29520);
nand UO_2295 (O_2295,N_28475,N_28417);
or UO_2296 (O_2296,N_29676,N_29001);
nor UO_2297 (O_2297,N_29911,N_29329);
nor UO_2298 (O_2298,N_29866,N_28642);
xor UO_2299 (O_2299,N_28760,N_29252);
and UO_2300 (O_2300,N_28156,N_29918);
nand UO_2301 (O_2301,N_28999,N_28659);
or UO_2302 (O_2302,N_29751,N_28524);
xor UO_2303 (O_2303,N_29075,N_29299);
nor UO_2304 (O_2304,N_28069,N_29255);
nand UO_2305 (O_2305,N_29416,N_28459);
nor UO_2306 (O_2306,N_29341,N_28618);
xor UO_2307 (O_2307,N_28993,N_29735);
nor UO_2308 (O_2308,N_29637,N_28781);
nor UO_2309 (O_2309,N_28428,N_28764);
xor UO_2310 (O_2310,N_28704,N_29807);
and UO_2311 (O_2311,N_29204,N_29471);
and UO_2312 (O_2312,N_28940,N_29455);
and UO_2313 (O_2313,N_29038,N_29839);
nand UO_2314 (O_2314,N_28537,N_29737);
and UO_2315 (O_2315,N_29781,N_28329);
nor UO_2316 (O_2316,N_29088,N_28562);
nor UO_2317 (O_2317,N_28134,N_29226);
nand UO_2318 (O_2318,N_29374,N_29341);
or UO_2319 (O_2319,N_28892,N_29737);
nand UO_2320 (O_2320,N_29475,N_28418);
or UO_2321 (O_2321,N_28534,N_28957);
xnor UO_2322 (O_2322,N_28446,N_28105);
or UO_2323 (O_2323,N_29755,N_28582);
nand UO_2324 (O_2324,N_28118,N_28174);
nor UO_2325 (O_2325,N_29424,N_29010);
nand UO_2326 (O_2326,N_29862,N_29302);
nand UO_2327 (O_2327,N_28044,N_28006);
and UO_2328 (O_2328,N_29537,N_28148);
nor UO_2329 (O_2329,N_28038,N_28947);
and UO_2330 (O_2330,N_28351,N_28734);
or UO_2331 (O_2331,N_29602,N_29224);
nor UO_2332 (O_2332,N_29772,N_28393);
and UO_2333 (O_2333,N_28427,N_28166);
xor UO_2334 (O_2334,N_29788,N_28113);
xnor UO_2335 (O_2335,N_28504,N_29797);
xor UO_2336 (O_2336,N_29779,N_28696);
or UO_2337 (O_2337,N_28006,N_28031);
nand UO_2338 (O_2338,N_28093,N_28374);
and UO_2339 (O_2339,N_29539,N_28188);
xnor UO_2340 (O_2340,N_28336,N_29090);
nand UO_2341 (O_2341,N_29756,N_28340);
and UO_2342 (O_2342,N_29112,N_28066);
nand UO_2343 (O_2343,N_28834,N_29816);
and UO_2344 (O_2344,N_28958,N_29737);
or UO_2345 (O_2345,N_28070,N_28003);
and UO_2346 (O_2346,N_29997,N_29165);
and UO_2347 (O_2347,N_28815,N_28717);
xor UO_2348 (O_2348,N_29874,N_28054);
xor UO_2349 (O_2349,N_28888,N_28007);
and UO_2350 (O_2350,N_29495,N_28139);
nor UO_2351 (O_2351,N_29219,N_28841);
or UO_2352 (O_2352,N_28696,N_29287);
xnor UO_2353 (O_2353,N_29946,N_28332);
and UO_2354 (O_2354,N_29796,N_29067);
nor UO_2355 (O_2355,N_28834,N_29938);
nor UO_2356 (O_2356,N_28282,N_28598);
nor UO_2357 (O_2357,N_29887,N_29939);
nand UO_2358 (O_2358,N_28760,N_28539);
or UO_2359 (O_2359,N_29376,N_28451);
nand UO_2360 (O_2360,N_28321,N_29893);
and UO_2361 (O_2361,N_28406,N_29898);
or UO_2362 (O_2362,N_29526,N_28081);
nor UO_2363 (O_2363,N_29596,N_29165);
or UO_2364 (O_2364,N_28486,N_29734);
or UO_2365 (O_2365,N_28608,N_28824);
and UO_2366 (O_2366,N_29229,N_28454);
nor UO_2367 (O_2367,N_28606,N_28282);
nand UO_2368 (O_2368,N_28641,N_28208);
xor UO_2369 (O_2369,N_29730,N_28894);
xor UO_2370 (O_2370,N_29979,N_28945);
nor UO_2371 (O_2371,N_29614,N_29962);
or UO_2372 (O_2372,N_29483,N_29492);
xnor UO_2373 (O_2373,N_28780,N_29079);
xnor UO_2374 (O_2374,N_29788,N_29763);
nand UO_2375 (O_2375,N_28677,N_28631);
xnor UO_2376 (O_2376,N_29382,N_29055);
nand UO_2377 (O_2377,N_29021,N_29472);
xor UO_2378 (O_2378,N_28119,N_28340);
and UO_2379 (O_2379,N_28347,N_28572);
and UO_2380 (O_2380,N_28454,N_28117);
or UO_2381 (O_2381,N_28227,N_29072);
nor UO_2382 (O_2382,N_29402,N_28111);
or UO_2383 (O_2383,N_29658,N_28622);
or UO_2384 (O_2384,N_28325,N_28130);
xor UO_2385 (O_2385,N_28384,N_29742);
nand UO_2386 (O_2386,N_28097,N_28749);
or UO_2387 (O_2387,N_29783,N_29984);
nand UO_2388 (O_2388,N_29764,N_28455);
xnor UO_2389 (O_2389,N_28388,N_29342);
or UO_2390 (O_2390,N_29228,N_29995);
xor UO_2391 (O_2391,N_29339,N_28337);
nor UO_2392 (O_2392,N_29264,N_29534);
xor UO_2393 (O_2393,N_28866,N_29457);
nand UO_2394 (O_2394,N_28709,N_29756);
and UO_2395 (O_2395,N_28235,N_28684);
and UO_2396 (O_2396,N_28672,N_28185);
and UO_2397 (O_2397,N_29329,N_29166);
xnor UO_2398 (O_2398,N_29441,N_29795);
nand UO_2399 (O_2399,N_28317,N_29088);
nor UO_2400 (O_2400,N_28691,N_28192);
nor UO_2401 (O_2401,N_29040,N_28891);
or UO_2402 (O_2402,N_28347,N_28302);
and UO_2403 (O_2403,N_28789,N_28369);
nand UO_2404 (O_2404,N_29755,N_29671);
xnor UO_2405 (O_2405,N_28827,N_29138);
nand UO_2406 (O_2406,N_28928,N_29819);
nor UO_2407 (O_2407,N_29370,N_29058);
nand UO_2408 (O_2408,N_29814,N_28465);
nor UO_2409 (O_2409,N_29128,N_29189);
nor UO_2410 (O_2410,N_29901,N_28091);
nor UO_2411 (O_2411,N_28962,N_29848);
or UO_2412 (O_2412,N_28205,N_29793);
xor UO_2413 (O_2413,N_29797,N_29124);
and UO_2414 (O_2414,N_29407,N_29372);
and UO_2415 (O_2415,N_28990,N_28885);
and UO_2416 (O_2416,N_29928,N_29932);
and UO_2417 (O_2417,N_28957,N_29577);
nand UO_2418 (O_2418,N_28432,N_29232);
and UO_2419 (O_2419,N_28525,N_29952);
nor UO_2420 (O_2420,N_28997,N_29545);
and UO_2421 (O_2421,N_28548,N_28095);
nand UO_2422 (O_2422,N_29000,N_28706);
nor UO_2423 (O_2423,N_28048,N_29622);
or UO_2424 (O_2424,N_29042,N_29552);
nor UO_2425 (O_2425,N_28840,N_28040);
nor UO_2426 (O_2426,N_29306,N_28422);
nand UO_2427 (O_2427,N_29022,N_29297);
and UO_2428 (O_2428,N_29147,N_29424);
or UO_2429 (O_2429,N_29014,N_28420);
or UO_2430 (O_2430,N_28775,N_28598);
or UO_2431 (O_2431,N_29223,N_29091);
xor UO_2432 (O_2432,N_29366,N_28702);
and UO_2433 (O_2433,N_29561,N_28693);
nor UO_2434 (O_2434,N_28368,N_28609);
nand UO_2435 (O_2435,N_28074,N_28659);
or UO_2436 (O_2436,N_29000,N_29964);
xor UO_2437 (O_2437,N_29242,N_29748);
nor UO_2438 (O_2438,N_28775,N_28213);
or UO_2439 (O_2439,N_29750,N_29188);
nor UO_2440 (O_2440,N_29825,N_28449);
xnor UO_2441 (O_2441,N_28412,N_29617);
and UO_2442 (O_2442,N_29672,N_29547);
xor UO_2443 (O_2443,N_28156,N_28699);
and UO_2444 (O_2444,N_29778,N_29562);
xnor UO_2445 (O_2445,N_28399,N_28652);
or UO_2446 (O_2446,N_29141,N_28467);
or UO_2447 (O_2447,N_29542,N_28089);
nand UO_2448 (O_2448,N_29850,N_28745);
nand UO_2449 (O_2449,N_29547,N_28479);
xor UO_2450 (O_2450,N_29860,N_28793);
and UO_2451 (O_2451,N_28525,N_29470);
nand UO_2452 (O_2452,N_29980,N_28348);
nor UO_2453 (O_2453,N_29275,N_29033);
and UO_2454 (O_2454,N_28527,N_28872);
or UO_2455 (O_2455,N_28018,N_29629);
xor UO_2456 (O_2456,N_29797,N_28677);
xor UO_2457 (O_2457,N_29798,N_29176);
or UO_2458 (O_2458,N_28659,N_29614);
and UO_2459 (O_2459,N_28410,N_29560);
or UO_2460 (O_2460,N_29981,N_29468);
xor UO_2461 (O_2461,N_29150,N_29654);
nor UO_2462 (O_2462,N_28025,N_29411);
nand UO_2463 (O_2463,N_28828,N_28116);
and UO_2464 (O_2464,N_29494,N_29821);
and UO_2465 (O_2465,N_29486,N_28729);
nor UO_2466 (O_2466,N_29272,N_28132);
nor UO_2467 (O_2467,N_28651,N_28835);
nor UO_2468 (O_2468,N_28367,N_29443);
or UO_2469 (O_2469,N_29315,N_29812);
nand UO_2470 (O_2470,N_29336,N_29730);
nand UO_2471 (O_2471,N_29560,N_29612);
nand UO_2472 (O_2472,N_29329,N_29695);
xor UO_2473 (O_2473,N_28031,N_29369);
nor UO_2474 (O_2474,N_28930,N_28739);
and UO_2475 (O_2475,N_29738,N_29318);
and UO_2476 (O_2476,N_29880,N_29223);
and UO_2477 (O_2477,N_29759,N_29732);
nand UO_2478 (O_2478,N_29322,N_28676);
nand UO_2479 (O_2479,N_29108,N_29434);
and UO_2480 (O_2480,N_29652,N_28369);
or UO_2481 (O_2481,N_29129,N_29486);
nand UO_2482 (O_2482,N_29921,N_29200);
and UO_2483 (O_2483,N_28339,N_28438);
and UO_2484 (O_2484,N_28644,N_28076);
or UO_2485 (O_2485,N_29551,N_28237);
xnor UO_2486 (O_2486,N_29460,N_28404);
nand UO_2487 (O_2487,N_28822,N_28722);
or UO_2488 (O_2488,N_28175,N_29685);
xnor UO_2489 (O_2489,N_28414,N_28356);
nand UO_2490 (O_2490,N_28211,N_29661);
nand UO_2491 (O_2491,N_28487,N_29568);
or UO_2492 (O_2492,N_28473,N_28106);
or UO_2493 (O_2493,N_29286,N_28008);
xor UO_2494 (O_2494,N_28505,N_29298);
or UO_2495 (O_2495,N_29851,N_29190);
nor UO_2496 (O_2496,N_28678,N_28371);
nand UO_2497 (O_2497,N_28075,N_29678);
nor UO_2498 (O_2498,N_28566,N_28048);
nor UO_2499 (O_2499,N_29103,N_28676);
xnor UO_2500 (O_2500,N_28790,N_28963);
nand UO_2501 (O_2501,N_29218,N_29304);
and UO_2502 (O_2502,N_29118,N_29484);
or UO_2503 (O_2503,N_29979,N_29611);
or UO_2504 (O_2504,N_28708,N_28415);
nand UO_2505 (O_2505,N_28902,N_29888);
xnor UO_2506 (O_2506,N_28826,N_29476);
or UO_2507 (O_2507,N_29414,N_29960);
nor UO_2508 (O_2508,N_28698,N_28121);
and UO_2509 (O_2509,N_29139,N_29839);
or UO_2510 (O_2510,N_29794,N_28948);
or UO_2511 (O_2511,N_29244,N_28571);
nor UO_2512 (O_2512,N_29718,N_28027);
xor UO_2513 (O_2513,N_28129,N_29048);
or UO_2514 (O_2514,N_29888,N_28769);
nand UO_2515 (O_2515,N_29856,N_28989);
xor UO_2516 (O_2516,N_28512,N_28552);
nand UO_2517 (O_2517,N_28642,N_29992);
and UO_2518 (O_2518,N_28834,N_29849);
or UO_2519 (O_2519,N_29341,N_28741);
nand UO_2520 (O_2520,N_28953,N_29596);
nand UO_2521 (O_2521,N_29425,N_28387);
nor UO_2522 (O_2522,N_28846,N_29435);
nor UO_2523 (O_2523,N_28798,N_29704);
or UO_2524 (O_2524,N_29605,N_28030);
xor UO_2525 (O_2525,N_28563,N_28693);
nand UO_2526 (O_2526,N_29462,N_29987);
or UO_2527 (O_2527,N_28824,N_28196);
or UO_2528 (O_2528,N_29772,N_29916);
or UO_2529 (O_2529,N_28649,N_28847);
xor UO_2530 (O_2530,N_28757,N_28302);
nand UO_2531 (O_2531,N_28945,N_28853);
and UO_2532 (O_2532,N_29937,N_28620);
nor UO_2533 (O_2533,N_29902,N_29327);
xnor UO_2534 (O_2534,N_29567,N_28004);
xor UO_2535 (O_2535,N_28130,N_29659);
or UO_2536 (O_2536,N_28940,N_29582);
or UO_2537 (O_2537,N_28301,N_29621);
or UO_2538 (O_2538,N_29127,N_28106);
nand UO_2539 (O_2539,N_29095,N_28961);
nor UO_2540 (O_2540,N_29494,N_29128);
xor UO_2541 (O_2541,N_28345,N_29219);
nand UO_2542 (O_2542,N_28278,N_28917);
xnor UO_2543 (O_2543,N_29780,N_28447);
nor UO_2544 (O_2544,N_28146,N_28488);
xor UO_2545 (O_2545,N_29048,N_29600);
nor UO_2546 (O_2546,N_28892,N_29405);
or UO_2547 (O_2547,N_29412,N_29162);
nor UO_2548 (O_2548,N_29826,N_28076);
nor UO_2549 (O_2549,N_29805,N_29048);
xor UO_2550 (O_2550,N_28003,N_28941);
nor UO_2551 (O_2551,N_29229,N_29897);
xor UO_2552 (O_2552,N_28144,N_29112);
xor UO_2553 (O_2553,N_29824,N_28748);
xor UO_2554 (O_2554,N_28482,N_29831);
nor UO_2555 (O_2555,N_29823,N_29736);
nor UO_2556 (O_2556,N_29939,N_29482);
nor UO_2557 (O_2557,N_29209,N_28000);
and UO_2558 (O_2558,N_28537,N_28078);
xor UO_2559 (O_2559,N_28706,N_28320);
and UO_2560 (O_2560,N_28721,N_29079);
nor UO_2561 (O_2561,N_29243,N_29435);
and UO_2562 (O_2562,N_28794,N_28526);
or UO_2563 (O_2563,N_28015,N_28237);
and UO_2564 (O_2564,N_28751,N_29492);
xor UO_2565 (O_2565,N_28291,N_29737);
xor UO_2566 (O_2566,N_28247,N_29636);
nor UO_2567 (O_2567,N_28106,N_28450);
nand UO_2568 (O_2568,N_28193,N_29373);
and UO_2569 (O_2569,N_29820,N_28860);
xor UO_2570 (O_2570,N_28839,N_28503);
or UO_2571 (O_2571,N_28231,N_28409);
xnor UO_2572 (O_2572,N_28200,N_29591);
nand UO_2573 (O_2573,N_29313,N_28529);
nand UO_2574 (O_2574,N_28912,N_28183);
and UO_2575 (O_2575,N_28163,N_28132);
and UO_2576 (O_2576,N_29013,N_28162);
or UO_2577 (O_2577,N_29710,N_28165);
nor UO_2578 (O_2578,N_29897,N_28227);
nor UO_2579 (O_2579,N_29265,N_28663);
and UO_2580 (O_2580,N_29231,N_28642);
nor UO_2581 (O_2581,N_28998,N_29259);
and UO_2582 (O_2582,N_28217,N_29106);
xor UO_2583 (O_2583,N_28195,N_28728);
and UO_2584 (O_2584,N_28551,N_28077);
xnor UO_2585 (O_2585,N_28382,N_28425);
nand UO_2586 (O_2586,N_29591,N_29705);
and UO_2587 (O_2587,N_28753,N_28389);
nor UO_2588 (O_2588,N_28158,N_28052);
and UO_2589 (O_2589,N_28909,N_29321);
nor UO_2590 (O_2590,N_28258,N_29243);
and UO_2591 (O_2591,N_28509,N_29524);
or UO_2592 (O_2592,N_29186,N_28830);
or UO_2593 (O_2593,N_29827,N_29007);
nor UO_2594 (O_2594,N_29800,N_28241);
nor UO_2595 (O_2595,N_29509,N_29914);
or UO_2596 (O_2596,N_28886,N_29971);
and UO_2597 (O_2597,N_29345,N_29717);
and UO_2598 (O_2598,N_29265,N_28068);
or UO_2599 (O_2599,N_28608,N_28378);
xor UO_2600 (O_2600,N_29890,N_29088);
nand UO_2601 (O_2601,N_28273,N_28617);
and UO_2602 (O_2602,N_29383,N_28638);
nor UO_2603 (O_2603,N_28662,N_29926);
and UO_2604 (O_2604,N_28803,N_28844);
nor UO_2605 (O_2605,N_29835,N_28416);
nand UO_2606 (O_2606,N_28161,N_28033);
xor UO_2607 (O_2607,N_28526,N_28826);
nor UO_2608 (O_2608,N_28843,N_28172);
nor UO_2609 (O_2609,N_28021,N_28383);
or UO_2610 (O_2610,N_29895,N_28167);
nand UO_2611 (O_2611,N_29540,N_29174);
nor UO_2612 (O_2612,N_29708,N_29496);
nand UO_2613 (O_2613,N_28512,N_29779);
and UO_2614 (O_2614,N_29458,N_28682);
nor UO_2615 (O_2615,N_29641,N_28118);
or UO_2616 (O_2616,N_29185,N_28308);
nand UO_2617 (O_2617,N_29114,N_29790);
nand UO_2618 (O_2618,N_28265,N_28433);
xnor UO_2619 (O_2619,N_28057,N_29251);
nor UO_2620 (O_2620,N_29699,N_28360);
xor UO_2621 (O_2621,N_29469,N_28997);
nor UO_2622 (O_2622,N_28830,N_29550);
nor UO_2623 (O_2623,N_29494,N_28042);
nor UO_2624 (O_2624,N_29061,N_29621);
or UO_2625 (O_2625,N_29846,N_29513);
and UO_2626 (O_2626,N_29507,N_28229);
nor UO_2627 (O_2627,N_29368,N_28073);
xnor UO_2628 (O_2628,N_29344,N_28520);
nand UO_2629 (O_2629,N_29431,N_28666);
and UO_2630 (O_2630,N_29878,N_29955);
xor UO_2631 (O_2631,N_28049,N_29482);
nor UO_2632 (O_2632,N_28799,N_28387);
nand UO_2633 (O_2633,N_29305,N_29280);
and UO_2634 (O_2634,N_28504,N_29681);
nand UO_2635 (O_2635,N_28548,N_28501);
and UO_2636 (O_2636,N_28940,N_29522);
or UO_2637 (O_2637,N_29652,N_28796);
nand UO_2638 (O_2638,N_28159,N_28098);
xor UO_2639 (O_2639,N_29478,N_29711);
nor UO_2640 (O_2640,N_28698,N_28330);
nand UO_2641 (O_2641,N_28852,N_29092);
and UO_2642 (O_2642,N_29254,N_28124);
and UO_2643 (O_2643,N_28555,N_28316);
nand UO_2644 (O_2644,N_28867,N_28673);
nor UO_2645 (O_2645,N_29767,N_29302);
xnor UO_2646 (O_2646,N_29589,N_28147);
nor UO_2647 (O_2647,N_28562,N_28216);
xnor UO_2648 (O_2648,N_29826,N_28157);
nor UO_2649 (O_2649,N_28482,N_28846);
and UO_2650 (O_2650,N_29699,N_29026);
xnor UO_2651 (O_2651,N_29177,N_29987);
nor UO_2652 (O_2652,N_28461,N_29436);
xor UO_2653 (O_2653,N_29299,N_28279);
xor UO_2654 (O_2654,N_29566,N_28484);
and UO_2655 (O_2655,N_28254,N_29298);
xnor UO_2656 (O_2656,N_28832,N_29506);
nor UO_2657 (O_2657,N_29539,N_28216);
xnor UO_2658 (O_2658,N_28831,N_28631);
nand UO_2659 (O_2659,N_28564,N_28929);
or UO_2660 (O_2660,N_28377,N_29967);
xnor UO_2661 (O_2661,N_28906,N_28358);
nand UO_2662 (O_2662,N_28824,N_29332);
nor UO_2663 (O_2663,N_28177,N_29565);
nand UO_2664 (O_2664,N_29042,N_28410);
or UO_2665 (O_2665,N_28626,N_28133);
and UO_2666 (O_2666,N_28511,N_28069);
and UO_2667 (O_2667,N_28986,N_28256);
or UO_2668 (O_2668,N_29023,N_28395);
nor UO_2669 (O_2669,N_28048,N_28086);
or UO_2670 (O_2670,N_28600,N_29978);
nor UO_2671 (O_2671,N_28368,N_29340);
nor UO_2672 (O_2672,N_29740,N_29593);
nand UO_2673 (O_2673,N_29917,N_29878);
xnor UO_2674 (O_2674,N_29684,N_28337);
or UO_2675 (O_2675,N_29742,N_28345);
nand UO_2676 (O_2676,N_28875,N_28695);
xnor UO_2677 (O_2677,N_28040,N_29268);
xnor UO_2678 (O_2678,N_29990,N_29073);
nand UO_2679 (O_2679,N_29107,N_29562);
nand UO_2680 (O_2680,N_29318,N_29743);
xor UO_2681 (O_2681,N_28187,N_28103);
and UO_2682 (O_2682,N_29911,N_28866);
or UO_2683 (O_2683,N_28579,N_28883);
and UO_2684 (O_2684,N_28935,N_29809);
nand UO_2685 (O_2685,N_29870,N_29908);
xnor UO_2686 (O_2686,N_28980,N_29673);
xnor UO_2687 (O_2687,N_28898,N_28785);
or UO_2688 (O_2688,N_28834,N_29662);
or UO_2689 (O_2689,N_28528,N_28441);
or UO_2690 (O_2690,N_29081,N_29813);
nand UO_2691 (O_2691,N_28721,N_29551);
and UO_2692 (O_2692,N_29507,N_28964);
xnor UO_2693 (O_2693,N_28525,N_28044);
or UO_2694 (O_2694,N_29042,N_29721);
and UO_2695 (O_2695,N_29974,N_29017);
xor UO_2696 (O_2696,N_28676,N_29548);
xnor UO_2697 (O_2697,N_28977,N_28613);
or UO_2698 (O_2698,N_29078,N_29952);
and UO_2699 (O_2699,N_29879,N_28203);
and UO_2700 (O_2700,N_28399,N_28890);
nor UO_2701 (O_2701,N_29296,N_28749);
nor UO_2702 (O_2702,N_29075,N_28314);
nand UO_2703 (O_2703,N_28211,N_28081);
and UO_2704 (O_2704,N_28776,N_28270);
nand UO_2705 (O_2705,N_28205,N_28153);
nor UO_2706 (O_2706,N_29348,N_28318);
or UO_2707 (O_2707,N_28803,N_28408);
and UO_2708 (O_2708,N_28617,N_29403);
xor UO_2709 (O_2709,N_28169,N_28916);
nand UO_2710 (O_2710,N_29942,N_29201);
or UO_2711 (O_2711,N_29745,N_29839);
or UO_2712 (O_2712,N_28159,N_28923);
nor UO_2713 (O_2713,N_29581,N_28159);
nor UO_2714 (O_2714,N_29349,N_28550);
or UO_2715 (O_2715,N_29984,N_29497);
xor UO_2716 (O_2716,N_28324,N_29853);
xor UO_2717 (O_2717,N_28262,N_29490);
or UO_2718 (O_2718,N_29645,N_29998);
nand UO_2719 (O_2719,N_29396,N_28247);
xnor UO_2720 (O_2720,N_29635,N_28214);
or UO_2721 (O_2721,N_29423,N_29991);
nand UO_2722 (O_2722,N_28226,N_28211);
and UO_2723 (O_2723,N_29344,N_29617);
nand UO_2724 (O_2724,N_28160,N_29344);
nor UO_2725 (O_2725,N_28392,N_28069);
or UO_2726 (O_2726,N_28897,N_29576);
and UO_2727 (O_2727,N_29930,N_28662);
xnor UO_2728 (O_2728,N_29956,N_29629);
or UO_2729 (O_2729,N_28806,N_28313);
nand UO_2730 (O_2730,N_29905,N_29598);
or UO_2731 (O_2731,N_29022,N_29287);
xnor UO_2732 (O_2732,N_29440,N_29150);
xor UO_2733 (O_2733,N_28490,N_29874);
xnor UO_2734 (O_2734,N_29412,N_29586);
and UO_2735 (O_2735,N_28940,N_29344);
xnor UO_2736 (O_2736,N_28608,N_29263);
nor UO_2737 (O_2737,N_28366,N_28403);
and UO_2738 (O_2738,N_29455,N_28189);
nor UO_2739 (O_2739,N_29485,N_29660);
nor UO_2740 (O_2740,N_29218,N_28741);
nand UO_2741 (O_2741,N_29175,N_28902);
or UO_2742 (O_2742,N_28256,N_28060);
nand UO_2743 (O_2743,N_29907,N_28253);
or UO_2744 (O_2744,N_29451,N_28672);
or UO_2745 (O_2745,N_29569,N_28150);
and UO_2746 (O_2746,N_28724,N_29563);
and UO_2747 (O_2747,N_28907,N_29976);
or UO_2748 (O_2748,N_28946,N_28746);
or UO_2749 (O_2749,N_29886,N_29814);
xnor UO_2750 (O_2750,N_29349,N_28582);
nand UO_2751 (O_2751,N_29987,N_28318);
xnor UO_2752 (O_2752,N_29670,N_29564);
or UO_2753 (O_2753,N_29659,N_28776);
and UO_2754 (O_2754,N_29360,N_29308);
nand UO_2755 (O_2755,N_28145,N_28240);
or UO_2756 (O_2756,N_29016,N_29633);
or UO_2757 (O_2757,N_28777,N_28876);
or UO_2758 (O_2758,N_28568,N_28302);
nor UO_2759 (O_2759,N_29332,N_29998);
and UO_2760 (O_2760,N_28109,N_28989);
nor UO_2761 (O_2761,N_29132,N_29465);
nor UO_2762 (O_2762,N_28118,N_28264);
nand UO_2763 (O_2763,N_29663,N_28674);
nand UO_2764 (O_2764,N_29024,N_29174);
and UO_2765 (O_2765,N_29863,N_29190);
and UO_2766 (O_2766,N_28364,N_28174);
or UO_2767 (O_2767,N_28482,N_28997);
xnor UO_2768 (O_2768,N_28089,N_29902);
nand UO_2769 (O_2769,N_28930,N_28887);
and UO_2770 (O_2770,N_29595,N_28738);
nand UO_2771 (O_2771,N_28829,N_28211);
or UO_2772 (O_2772,N_29597,N_29875);
and UO_2773 (O_2773,N_28461,N_29154);
nand UO_2774 (O_2774,N_28292,N_29476);
and UO_2775 (O_2775,N_28850,N_29139);
and UO_2776 (O_2776,N_28140,N_28571);
nor UO_2777 (O_2777,N_28684,N_28424);
nor UO_2778 (O_2778,N_28374,N_28655);
nand UO_2779 (O_2779,N_28855,N_28182);
xor UO_2780 (O_2780,N_29771,N_28673);
or UO_2781 (O_2781,N_29487,N_29381);
nor UO_2782 (O_2782,N_29440,N_28534);
nor UO_2783 (O_2783,N_29588,N_29460);
nand UO_2784 (O_2784,N_29988,N_29363);
and UO_2785 (O_2785,N_29125,N_28986);
nor UO_2786 (O_2786,N_28749,N_28608);
nor UO_2787 (O_2787,N_28419,N_29253);
nor UO_2788 (O_2788,N_29637,N_28684);
nor UO_2789 (O_2789,N_29894,N_28396);
or UO_2790 (O_2790,N_28771,N_28945);
xor UO_2791 (O_2791,N_29157,N_28339);
xor UO_2792 (O_2792,N_28137,N_29059);
nand UO_2793 (O_2793,N_29822,N_29467);
or UO_2794 (O_2794,N_28907,N_28080);
and UO_2795 (O_2795,N_29158,N_29856);
xnor UO_2796 (O_2796,N_28075,N_29832);
or UO_2797 (O_2797,N_29328,N_28737);
nor UO_2798 (O_2798,N_28952,N_28513);
nand UO_2799 (O_2799,N_29507,N_29696);
or UO_2800 (O_2800,N_28590,N_28552);
nor UO_2801 (O_2801,N_29743,N_28204);
and UO_2802 (O_2802,N_28996,N_29647);
xor UO_2803 (O_2803,N_28006,N_29784);
nor UO_2804 (O_2804,N_29778,N_29800);
xor UO_2805 (O_2805,N_29848,N_29843);
nand UO_2806 (O_2806,N_28926,N_28561);
nor UO_2807 (O_2807,N_29842,N_28125);
nor UO_2808 (O_2808,N_28236,N_29202);
nand UO_2809 (O_2809,N_29049,N_29400);
nand UO_2810 (O_2810,N_29530,N_28298);
and UO_2811 (O_2811,N_28954,N_29005);
nor UO_2812 (O_2812,N_29711,N_29004);
or UO_2813 (O_2813,N_29310,N_28138);
and UO_2814 (O_2814,N_29703,N_28866);
nor UO_2815 (O_2815,N_28707,N_29432);
xor UO_2816 (O_2816,N_29694,N_28935);
nor UO_2817 (O_2817,N_29807,N_29135);
or UO_2818 (O_2818,N_28831,N_28694);
nor UO_2819 (O_2819,N_29175,N_29229);
or UO_2820 (O_2820,N_28758,N_28315);
xor UO_2821 (O_2821,N_29072,N_29601);
or UO_2822 (O_2822,N_29931,N_28093);
xor UO_2823 (O_2823,N_29627,N_29199);
xnor UO_2824 (O_2824,N_29477,N_28332);
and UO_2825 (O_2825,N_29867,N_28713);
or UO_2826 (O_2826,N_28673,N_28450);
nand UO_2827 (O_2827,N_29753,N_29709);
xnor UO_2828 (O_2828,N_29073,N_29763);
and UO_2829 (O_2829,N_29399,N_28769);
or UO_2830 (O_2830,N_29697,N_29631);
and UO_2831 (O_2831,N_29724,N_28821);
nor UO_2832 (O_2832,N_28972,N_28172);
nor UO_2833 (O_2833,N_28157,N_28053);
or UO_2834 (O_2834,N_29853,N_29030);
or UO_2835 (O_2835,N_28524,N_28825);
xor UO_2836 (O_2836,N_29249,N_29731);
or UO_2837 (O_2837,N_28930,N_28869);
xor UO_2838 (O_2838,N_28511,N_29968);
nor UO_2839 (O_2839,N_28593,N_29078);
nor UO_2840 (O_2840,N_29396,N_28782);
xor UO_2841 (O_2841,N_29638,N_28487);
or UO_2842 (O_2842,N_29414,N_28156);
nand UO_2843 (O_2843,N_29725,N_28667);
xnor UO_2844 (O_2844,N_28973,N_29889);
xnor UO_2845 (O_2845,N_29941,N_29850);
or UO_2846 (O_2846,N_28029,N_29331);
and UO_2847 (O_2847,N_29775,N_29367);
nor UO_2848 (O_2848,N_29537,N_29666);
nand UO_2849 (O_2849,N_28087,N_28063);
or UO_2850 (O_2850,N_28140,N_28417);
nor UO_2851 (O_2851,N_29595,N_29288);
xor UO_2852 (O_2852,N_29180,N_28309);
and UO_2853 (O_2853,N_28575,N_29495);
nand UO_2854 (O_2854,N_28627,N_29296);
nor UO_2855 (O_2855,N_28032,N_28206);
or UO_2856 (O_2856,N_29465,N_28388);
nor UO_2857 (O_2857,N_28095,N_29125);
nor UO_2858 (O_2858,N_28044,N_28492);
and UO_2859 (O_2859,N_29136,N_29267);
nand UO_2860 (O_2860,N_28836,N_29154);
or UO_2861 (O_2861,N_29383,N_28808);
nand UO_2862 (O_2862,N_28107,N_29294);
or UO_2863 (O_2863,N_28290,N_29758);
and UO_2864 (O_2864,N_28978,N_28291);
or UO_2865 (O_2865,N_28542,N_28374);
nand UO_2866 (O_2866,N_28010,N_29224);
nor UO_2867 (O_2867,N_28840,N_28000);
nor UO_2868 (O_2868,N_28808,N_29586);
nor UO_2869 (O_2869,N_29873,N_28001);
nor UO_2870 (O_2870,N_28223,N_29935);
or UO_2871 (O_2871,N_29409,N_29326);
xnor UO_2872 (O_2872,N_28283,N_28544);
xnor UO_2873 (O_2873,N_29443,N_29439);
xnor UO_2874 (O_2874,N_28991,N_28303);
nor UO_2875 (O_2875,N_29299,N_29246);
nand UO_2876 (O_2876,N_29266,N_28793);
xor UO_2877 (O_2877,N_28732,N_28745);
and UO_2878 (O_2878,N_29309,N_29156);
nor UO_2879 (O_2879,N_28124,N_28337);
and UO_2880 (O_2880,N_28903,N_28048);
xor UO_2881 (O_2881,N_29124,N_29905);
and UO_2882 (O_2882,N_28850,N_28389);
and UO_2883 (O_2883,N_29517,N_29430);
xnor UO_2884 (O_2884,N_28956,N_28410);
nor UO_2885 (O_2885,N_29712,N_28770);
nor UO_2886 (O_2886,N_28363,N_28490);
nand UO_2887 (O_2887,N_29380,N_28988);
nand UO_2888 (O_2888,N_29070,N_28816);
nand UO_2889 (O_2889,N_28046,N_28574);
xnor UO_2890 (O_2890,N_29538,N_29641);
or UO_2891 (O_2891,N_28114,N_28681);
nor UO_2892 (O_2892,N_29597,N_29012);
nand UO_2893 (O_2893,N_29259,N_28094);
or UO_2894 (O_2894,N_28904,N_29849);
xor UO_2895 (O_2895,N_29267,N_29657);
and UO_2896 (O_2896,N_29386,N_28809);
or UO_2897 (O_2897,N_28801,N_29456);
or UO_2898 (O_2898,N_29451,N_28334);
or UO_2899 (O_2899,N_28904,N_28040);
nand UO_2900 (O_2900,N_28420,N_28655);
xor UO_2901 (O_2901,N_29432,N_28410);
xnor UO_2902 (O_2902,N_29467,N_28872);
or UO_2903 (O_2903,N_28382,N_29736);
and UO_2904 (O_2904,N_28255,N_29681);
xnor UO_2905 (O_2905,N_29683,N_28639);
or UO_2906 (O_2906,N_29272,N_28939);
nor UO_2907 (O_2907,N_28963,N_29189);
and UO_2908 (O_2908,N_29869,N_29122);
and UO_2909 (O_2909,N_28705,N_29576);
and UO_2910 (O_2910,N_28693,N_29121);
and UO_2911 (O_2911,N_28276,N_29496);
xnor UO_2912 (O_2912,N_29984,N_29453);
xnor UO_2913 (O_2913,N_28689,N_28901);
nor UO_2914 (O_2914,N_28936,N_29547);
or UO_2915 (O_2915,N_28684,N_28890);
nor UO_2916 (O_2916,N_28933,N_29511);
nor UO_2917 (O_2917,N_28875,N_28854);
nand UO_2918 (O_2918,N_28136,N_28415);
nor UO_2919 (O_2919,N_28954,N_29474);
or UO_2920 (O_2920,N_29233,N_29323);
nor UO_2921 (O_2921,N_29237,N_28531);
xor UO_2922 (O_2922,N_29060,N_28309);
nand UO_2923 (O_2923,N_29934,N_28188);
nand UO_2924 (O_2924,N_29876,N_28208);
nand UO_2925 (O_2925,N_29407,N_29442);
or UO_2926 (O_2926,N_28967,N_28428);
or UO_2927 (O_2927,N_29480,N_29693);
xor UO_2928 (O_2928,N_29186,N_29436);
and UO_2929 (O_2929,N_29676,N_28481);
and UO_2930 (O_2930,N_29000,N_28717);
nor UO_2931 (O_2931,N_28820,N_28791);
xor UO_2932 (O_2932,N_29726,N_28859);
and UO_2933 (O_2933,N_29438,N_29688);
or UO_2934 (O_2934,N_28039,N_28567);
xor UO_2935 (O_2935,N_29577,N_28433);
nor UO_2936 (O_2936,N_29848,N_29763);
nor UO_2937 (O_2937,N_28173,N_29661);
and UO_2938 (O_2938,N_29753,N_29722);
nand UO_2939 (O_2939,N_29459,N_29669);
xnor UO_2940 (O_2940,N_28588,N_28596);
nand UO_2941 (O_2941,N_29586,N_29829);
xnor UO_2942 (O_2942,N_28743,N_28559);
xor UO_2943 (O_2943,N_29106,N_29678);
and UO_2944 (O_2944,N_28051,N_29091);
nor UO_2945 (O_2945,N_28389,N_29722);
nand UO_2946 (O_2946,N_28382,N_29543);
and UO_2947 (O_2947,N_28560,N_29305);
nor UO_2948 (O_2948,N_29809,N_28852);
and UO_2949 (O_2949,N_29174,N_29679);
xnor UO_2950 (O_2950,N_28956,N_29693);
nor UO_2951 (O_2951,N_29283,N_29858);
or UO_2952 (O_2952,N_28200,N_29061);
or UO_2953 (O_2953,N_29197,N_28535);
and UO_2954 (O_2954,N_28250,N_29129);
xnor UO_2955 (O_2955,N_29140,N_28047);
and UO_2956 (O_2956,N_29866,N_29892);
nor UO_2957 (O_2957,N_28859,N_28108);
nand UO_2958 (O_2958,N_29389,N_28999);
or UO_2959 (O_2959,N_29407,N_28291);
and UO_2960 (O_2960,N_28679,N_28248);
nand UO_2961 (O_2961,N_28403,N_28581);
nand UO_2962 (O_2962,N_28433,N_29190);
nand UO_2963 (O_2963,N_29351,N_28902);
nor UO_2964 (O_2964,N_28530,N_28506);
or UO_2965 (O_2965,N_28265,N_29087);
or UO_2966 (O_2966,N_28279,N_29605);
xnor UO_2967 (O_2967,N_29807,N_29824);
nor UO_2968 (O_2968,N_28419,N_29286);
and UO_2969 (O_2969,N_29616,N_28911);
nor UO_2970 (O_2970,N_29175,N_29419);
nand UO_2971 (O_2971,N_29489,N_29696);
nand UO_2972 (O_2972,N_28906,N_29381);
and UO_2973 (O_2973,N_29017,N_28004);
or UO_2974 (O_2974,N_28126,N_28880);
nand UO_2975 (O_2975,N_29322,N_29928);
and UO_2976 (O_2976,N_29425,N_29934);
nand UO_2977 (O_2977,N_28232,N_28688);
or UO_2978 (O_2978,N_28233,N_29291);
and UO_2979 (O_2979,N_28346,N_28817);
nand UO_2980 (O_2980,N_29970,N_29574);
nand UO_2981 (O_2981,N_29955,N_28236);
nor UO_2982 (O_2982,N_28511,N_29198);
nand UO_2983 (O_2983,N_28135,N_29659);
and UO_2984 (O_2984,N_29459,N_28251);
and UO_2985 (O_2985,N_28016,N_28737);
xor UO_2986 (O_2986,N_28213,N_28516);
or UO_2987 (O_2987,N_28850,N_29662);
or UO_2988 (O_2988,N_28548,N_29376);
nand UO_2989 (O_2989,N_29954,N_29978);
nor UO_2990 (O_2990,N_29203,N_28531);
or UO_2991 (O_2991,N_28197,N_29641);
and UO_2992 (O_2992,N_28575,N_29899);
xnor UO_2993 (O_2993,N_28536,N_28133);
nand UO_2994 (O_2994,N_28263,N_29106);
xnor UO_2995 (O_2995,N_28365,N_29678);
xor UO_2996 (O_2996,N_28422,N_29556);
nor UO_2997 (O_2997,N_29555,N_28192);
xor UO_2998 (O_2998,N_28893,N_28491);
nand UO_2999 (O_2999,N_29181,N_28762);
and UO_3000 (O_3000,N_29766,N_28476);
and UO_3001 (O_3001,N_29571,N_29931);
and UO_3002 (O_3002,N_28192,N_29872);
xnor UO_3003 (O_3003,N_29905,N_29373);
or UO_3004 (O_3004,N_29146,N_29173);
nand UO_3005 (O_3005,N_29578,N_29020);
or UO_3006 (O_3006,N_29990,N_28951);
or UO_3007 (O_3007,N_29401,N_29701);
xnor UO_3008 (O_3008,N_28692,N_29393);
nand UO_3009 (O_3009,N_28950,N_29472);
nor UO_3010 (O_3010,N_28142,N_29980);
or UO_3011 (O_3011,N_28914,N_29052);
xor UO_3012 (O_3012,N_29546,N_28529);
or UO_3013 (O_3013,N_29033,N_29151);
xor UO_3014 (O_3014,N_29371,N_29990);
or UO_3015 (O_3015,N_29633,N_28691);
nand UO_3016 (O_3016,N_29260,N_28470);
nand UO_3017 (O_3017,N_29105,N_28510);
and UO_3018 (O_3018,N_28263,N_29666);
nor UO_3019 (O_3019,N_28938,N_29602);
nor UO_3020 (O_3020,N_28240,N_28251);
or UO_3021 (O_3021,N_29528,N_29012);
xnor UO_3022 (O_3022,N_29753,N_28018);
nor UO_3023 (O_3023,N_28916,N_29275);
and UO_3024 (O_3024,N_28971,N_28302);
or UO_3025 (O_3025,N_29829,N_28566);
or UO_3026 (O_3026,N_28273,N_28980);
nand UO_3027 (O_3027,N_28144,N_28140);
nand UO_3028 (O_3028,N_28632,N_28258);
nor UO_3029 (O_3029,N_28699,N_28672);
and UO_3030 (O_3030,N_29601,N_28568);
or UO_3031 (O_3031,N_29764,N_28464);
nor UO_3032 (O_3032,N_28706,N_29621);
or UO_3033 (O_3033,N_28297,N_28864);
or UO_3034 (O_3034,N_28035,N_29387);
nand UO_3035 (O_3035,N_29505,N_28913);
or UO_3036 (O_3036,N_29903,N_28785);
xor UO_3037 (O_3037,N_28672,N_28214);
or UO_3038 (O_3038,N_29536,N_28461);
xor UO_3039 (O_3039,N_28500,N_28115);
nor UO_3040 (O_3040,N_29705,N_29881);
xnor UO_3041 (O_3041,N_29693,N_28041);
nor UO_3042 (O_3042,N_28301,N_28350);
nor UO_3043 (O_3043,N_29246,N_29284);
or UO_3044 (O_3044,N_28043,N_29750);
nand UO_3045 (O_3045,N_29599,N_28223);
nor UO_3046 (O_3046,N_29535,N_29891);
or UO_3047 (O_3047,N_29217,N_28816);
nor UO_3048 (O_3048,N_28398,N_29713);
xor UO_3049 (O_3049,N_29347,N_28474);
and UO_3050 (O_3050,N_29436,N_29371);
and UO_3051 (O_3051,N_28116,N_28973);
and UO_3052 (O_3052,N_28255,N_28113);
nor UO_3053 (O_3053,N_29226,N_28774);
nor UO_3054 (O_3054,N_29667,N_29302);
xor UO_3055 (O_3055,N_28017,N_29942);
nor UO_3056 (O_3056,N_29356,N_29367);
xnor UO_3057 (O_3057,N_28397,N_29710);
xnor UO_3058 (O_3058,N_29089,N_29472);
nand UO_3059 (O_3059,N_28498,N_29422);
or UO_3060 (O_3060,N_28680,N_28433);
nor UO_3061 (O_3061,N_29204,N_28679);
xor UO_3062 (O_3062,N_29133,N_28790);
and UO_3063 (O_3063,N_29080,N_28456);
and UO_3064 (O_3064,N_28970,N_29860);
and UO_3065 (O_3065,N_28815,N_28496);
xor UO_3066 (O_3066,N_28996,N_28493);
nor UO_3067 (O_3067,N_29482,N_29135);
nand UO_3068 (O_3068,N_28433,N_29923);
and UO_3069 (O_3069,N_28629,N_29931);
xor UO_3070 (O_3070,N_28444,N_29190);
nor UO_3071 (O_3071,N_28593,N_28128);
nor UO_3072 (O_3072,N_29105,N_28160);
and UO_3073 (O_3073,N_28858,N_29768);
and UO_3074 (O_3074,N_29421,N_28931);
and UO_3075 (O_3075,N_29340,N_29071);
nor UO_3076 (O_3076,N_28517,N_28664);
xor UO_3077 (O_3077,N_28352,N_28015);
xnor UO_3078 (O_3078,N_28949,N_29730);
or UO_3079 (O_3079,N_28455,N_29325);
nor UO_3080 (O_3080,N_28512,N_29563);
nand UO_3081 (O_3081,N_28696,N_29910);
xor UO_3082 (O_3082,N_29264,N_29514);
nand UO_3083 (O_3083,N_28929,N_28305);
and UO_3084 (O_3084,N_29776,N_29976);
or UO_3085 (O_3085,N_29100,N_28726);
or UO_3086 (O_3086,N_28675,N_28050);
nor UO_3087 (O_3087,N_29255,N_28048);
or UO_3088 (O_3088,N_29990,N_28083);
nand UO_3089 (O_3089,N_29622,N_29907);
or UO_3090 (O_3090,N_28984,N_29707);
or UO_3091 (O_3091,N_29039,N_28759);
xor UO_3092 (O_3092,N_29980,N_28673);
xnor UO_3093 (O_3093,N_29766,N_28494);
nor UO_3094 (O_3094,N_28862,N_29106);
nand UO_3095 (O_3095,N_29168,N_29482);
and UO_3096 (O_3096,N_28964,N_28717);
nand UO_3097 (O_3097,N_28886,N_28048);
and UO_3098 (O_3098,N_29862,N_28546);
nand UO_3099 (O_3099,N_28635,N_28028);
nor UO_3100 (O_3100,N_28202,N_29611);
nand UO_3101 (O_3101,N_29430,N_28378);
and UO_3102 (O_3102,N_29204,N_29641);
nand UO_3103 (O_3103,N_29030,N_28891);
nand UO_3104 (O_3104,N_28288,N_28325);
nor UO_3105 (O_3105,N_28818,N_29371);
and UO_3106 (O_3106,N_28334,N_29287);
nor UO_3107 (O_3107,N_29062,N_28274);
xnor UO_3108 (O_3108,N_28218,N_29822);
xnor UO_3109 (O_3109,N_29677,N_28156);
or UO_3110 (O_3110,N_28523,N_29269);
xnor UO_3111 (O_3111,N_29664,N_29112);
and UO_3112 (O_3112,N_29135,N_28993);
nor UO_3113 (O_3113,N_28901,N_29044);
xor UO_3114 (O_3114,N_28296,N_29209);
nand UO_3115 (O_3115,N_29554,N_28988);
nand UO_3116 (O_3116,N_29105,N_28679);
and UO_3117 (O_3117,N_28128,N_29585);
and UO_3118 (O_3118,N_29079,N_29210);
and UO_3119 (O_3119,N_28565,N_28039);
nand UO_3120 (O_3120,N_29527,N_29729);
xnor UO_3121 (O_3121,N_29334,N_28373);
and UO_3122 (O_3122,N_28361,N_29929);
and UO_3123 (O_3123,N_28920,N_28147);
nor UO_3124 (O_3124,N_29618,N_29541);
or UO_3125 (O_3125,N_29009,N_28733);
xnor UO_3126 (O_3126,N_29249,N_28554);
xor UO_3127 (O_3127,N_29539,N_28116);
xor UO_3128 (O_3128,N_29270,N_29665);
nor UO_3129 (O_3129,N_28194,N_28978);
nor UO_3130 (O_3130,N_29454,N_28972);
and UO_3131 (O_3131,N_28065,N_28720);
xnor UO_3132 (O_3132,N_28110,N_28349);
and UO_3133 (O_3133,N_29522,N_28946);
and UO_3134 (O_3134,N_28436,N_29465);
xor UO_3135 (O_3135,N_28659,N_28104);
or UO_3136 (O_3136,N_28095,N_29611);
nand UO_3137 (O_3137,N_29358,N_28453);
or UO_3138 (O_3138,N_29861,N_29904);
xnor UO_3139 (O_3139,N_29778,N_29431);
or UO_3140 (O_3140,N_28243,N_28778);
xnor UO_3141 (O_3141,N_28303,N_29139);
nor UO_3142 (O_3142,N_29758,N_29937);
xnor UO_3143 (O_3143,N_29429,N_29349);
xnor UO_3144 (O_3144,N_29337,N_28353);
nand UO_3145 (O_3145,N_28345,N_28951);
nand UO_3146 (O_3146,N_28772,N_28534);
nor UO_3147 (O_3147,N_29658,N_29051);
nand UO_3148 (O_3148,N_28796,N_28203);
nor UO_3149 (O_3149,N_29444,N_28995);
or UO_3150 (O_3150,N_28473,N_28400);
and UO_3151 (O_3151,N_29445,N_29441);
and UO_3152 (O_3152,N_29517,N_29747);
xnor UO_3153 (O_3153,N_29295,N_28946);
xor UO_3154 (O_3154,N_28411,N_28012);
xor UO_3155 (O_3155,N_28194,N_29587);
nand UO_3156 (O_3156,N_28603,N_29245);
nand UO_3157 (O_3157,N_29310,N_28366);
xor UO_3158 (O_3158,N_28317,N_28895);
xnor UO_3159 (O_3159,N_28284,N_29747);
or UO_3160 (O_3160,N_29480,N_28123);
xor UO_3161 (O_3161,N_28532,N_29183);
xnor UO_3162 (O_3162,N_28354,N_29356);
nand UO_3163 (O_3163,N_28686,N_29919);
nor UO_3164 (O_3164,N_29885,N_28423);
nand UO_3165 (O_3165,N_28379,N_28798);
nor UO_3166 (O_3166,N_29675,N_28006);
nand UO_3167 (O_3167,N_28413,N_29226);
nand UO_3168 (O_3168,N_29550,N_29903);
or UO_3169 (O_3169,N_29334,N_29802);
and UO_3170 (O_3170,N_28614,N_29104);
xnor UO_3171 (O_3171,N_29934,N_28725);
nor UO_3172 (O_3172,N_29420,N_29721);
or UO_3173 (O_3173,N_28220,N_28964);
xnor UO_3174 (O_3174,N_28454,N_29397);
nor UO_3175 (O_3175,N_28896,N_28113);
nor UO_3176 (O_3176,N_28780,N_29928);
or UO_3177 (O_3177,N_28300,N_29401);
nor UO_3178 (O_3178,N_29591,N_29344);
nand UO_3179 (O_3179,N_28985,N_29704);
and UO_3180 (O_3180,N_28250,N_29905);
nor UO_3181 (O_3181,N_28698,N_28300);
nor UO_3182 (O_3182,N_29363,N_29856);
nor UO_3183 (O_3183,N_28325,N_29692);
and UO_3184 (O_3184,N_28812,N_29667);
and UO_3185 (O_3185,N_29117,N_28581);
nor UO_3186 (O_3186,N_28866,N_28403);
nand UO_3187 (O_3187,N_28716,N_29074);
xor UO_3188 (O_3188,N_29329,N_28875);
nand UO_3189 (O_3189,N_29873,N_28775);
xnor UO_3190 (O_3190,N_29681,N_29904);
nor UO_3191 (O_3191,N_29918,N_29262);
xnor UO_3192 (O_3192,N_28295,N_28956);
nand UO_3193 (O_3193,N_29297,N_28692);
or UO_3194 (O_3194,N_29624,N_29034);
nor UO_3195 (O_3195,N_28851,N_28211);
or UO_3196 (O_3196,N_28255,N_29496);
xor UO_3197 (O_3197,N_29420,N_28795);
xnor UO_3198 (O_3198,N_28128,N_28795);
xor UO_3199 (O_3199,N_29119,N_28578);
nand UO_3200 (O_3200,N_29347,N_29134);
nand UO_3201 (O_3201,N_29293,N_28573);
nand UO_3202 (O_3202,N_28669,N_28033);
xor UO_3203 (O_3203,N_29798,N_29300);
xnor UO_3204 (O_3204,N_29569,N_28803);
or UO_3205 (O_3205,N_29236,N_28825);
and UO_3206 (O_3206,N_28004,N_29615);
or UO_3207 (O_3207,N_28105,N_29016);
nand UO_3208 (O_3208,N_28239,N_29209);
nand UO_3209 (O_3209,N_29579,N_28698);
or UO_3210 (O_3210,N_28043,N_29627);
or UO_3211 (O_3211,N_28657,N_29714);
xnor UO_3212 (O_3212,N_28888,N_29409);
and UO_3213 (O_3213,N_28856,N_29916);
and UO_3214 (O_3214,N_29605,N_29118);
nand UO_3215 (O_3215,N_29886,N_28140);
and UO_3216 (O_3216,N_28895,N_29930);
or UO_3217 (O_3217,N_29158,N_28918);
nor UO_3218 (O_3218,N_28614,N_28917);
xnor UO_3219 (O_3219,N_29962,N_28936);
nor UO_3220 (O_3220,N_28722,N_28088);
xor UO_3221 (O_3221,N_28495,N_29110);
nor UO_3222 (O_3222,N_28255,N_28863);
nor UO_3223 (O_3223,N_29692,N_29191);
or UO_3224 (O_3224,N_29705,N_29076);
xor UO_3225 (O_3225,N_28643,N_29514);
xor UO_3226 (O_3226,N_29161,N_28432);
nor UO_3227 (O_3227,N_29963,N_28738);
nor UO_3228 (O_3228,N_28300,N_29172);
xor UO_3229 (O_3229,N_29833,N_29650);
nor UO_3230 (O_3230,N_29731,N_29388);
xor UO_3231 (O_3231,N_29275,N_29372);
nor UO_3232 (O_3232,N_29761,N_29000);
xnor UO_3233 (O_3233,N_29647,N_29039);
or UO_3234 (O_3234,N_29627,N_29172);
or UO_3235 (O_3235,N_29746,N_28220);
nor UO_3236 (O_3236,N_29663,N_28657);
and UO_3237 (O_3237,N_28304,N_29281);
nor UO_3238 (O_3238,N_29735,N_29548);
xnor UO_3239 (O_3239,N_29087,N_28924);
and UO_3240 (O_3240,N_28501,N_29663);
nand UO_3241 (O_3241,N_29423,N_28805);
xor UO_3242 (O_3242,N_29147,N_29031);
and UO_3243 (O_3243,N_28413,N_29106);
nand UO_3244 (O_3244,N_28379,N_28446);
nand UO_3245 (O_3245,N_29573,N_28888);
nor UO_3246 (O_3246,N_28606,N_28873);
and UO_3247 (O_3247,N_28669,N_29747);
and UO_3248 (O_3248,N_28667,N_29006);
nand UO_3249 (O_3249,N_28611,N_29334);
or UO_3250 (O_3250,N_28515,N_28596);
and UO_3251 (O_3251,N_28669,N_29120);
and UO_3252 (O_3252,N_29204,N_28097);
xor UO_3253 (O_3253,N_29849,N_29444);
or UO_3254 (O_3254,N_28019,N_29322);
nor UO_3255 (O_3255,N_28549,N_28650);
xor UO_3256 (O_3256,N_29274,N_28734);
xnor UO_3257 (O_3257,N_29283,N_29415);
xor UO_3258 (O_3258,N_28124,N_28366);
nor UO_3259 (O_3259,N_29459,N_29340);
nor UO_3260 (O_3260,N_29400,N_28328);
nor UO_3261 (O_3261,N_29012,N_29498);
nand UO_3262 (O_3262,N_28856,N_29312);
nand UO_3263 (O_3263,N_29960,N_29881);
nand UO_3264 (O_3264,N_28771,N_28795);
nand UO_3265 (O_3265,N_28905,N_28736);
or UO_3266 (O_3266,N_28522,N_29327);
nor UO_3267 (O_3267,N_29677,N_28195);
nand UO_3268 (O_3268,N_29892,N_29533);
nand UO_3269 (O_3269,N_28878,N_29053);
and UO_3270 (O_3270,N_28585,N_28487);
and UO_3271 (O_3271,N_28131,N_28842);
nor UO_3272 (O_3272,N_28455,N_28669);
nand UO_3273 (O_3273,N_29757,N_29044);
nand UO_3274 (O_3274,N_28356,N_29656);
xnor UO_3275 (O_3275,N_28415,N_29850);
nor UO_3276 (O_3276,N_29415,N_28171);
or UO_3277 (O_3277,N_29361,N_28701);
or UO_3278 (O_3278,N_29435,N_29429);
and UO_3279 (O_3279,N_28235,N_29658);
nand UO_3280 (O_3280,N_29126,N_29431);
nand UO_3281 (O_3281,N_28390,N_29762);
nor UO_3282 (O_3282,N_28812,N_28065);
and UO_3283 (O_3283,N_29202,N_29854);
nand UO_3284 (O_3284,N_29982,N_29020);
and UO_3285 (O_3285,N_29235,N_28885);
xor UO_3286 (O_3286,N_28143,N_29452);
xnor UO_3287 (O_3287,N_28605,N_28797);
xnor UO_3288 (O_3288,N_28495,N_28308);
xnor UO_3289 (O_3289,N_28330,N_29005);
and UO_3290 (O_3290,N_28359,N_28373);
nand UO_3291 (O_3291,N_29195,N_29664);
xnor UO_3292 (O_3292,N_28494,N_29844);
xnor UO_3293 (O_3293,N_29510,N_28971);
and UO_3294 (O_3294,N_28682,N_29143);
xor UO_3295 (O_3295,N_29772,N_29374);
nand UO_3296 (O_3296,N_28075,N_29674);
nor UO_3297 (O_3297,N_28623,N_28208);
or UO_3298 (O_3298,N_28026,N_28601);
or UO_3299 (O_3299,N_28199,N_29103);
nor UO_3300 (O_3300,N_29758,N_29400);
nor UO_3301 (O_3301,N_29769,N_29540);
or UO_3302 (O_3302,N_28228,N_29827);
nor UO_3303 (O_3303,N_29883,N_29082);
or UO_3304 (O_3304,N_29443,N_28494);
nand UO_3305 (O_3305,N_29428,N_29191);
nor UO_3306 (O_3306,N_28944,N_28125);
or UO_3307 (O_3307,N_28711,N_28996);
nor UO_3308 (O_3308,N_29060,N_28841);
nand UO_3309 (O_3309,N_28479,N_28133);
nand UO_3310 (O_3310,N_28498,N_29490);
or UO_3311 (O_3311,N_28251,N_28910);
and UO_3312 (O_3312,N_28134,N_28309);
or UO_3313 (O_3313,N_28113,N_28832);
nor UO_3314 (O_3314,N_29873,N_29864);
nor UO_3315 (O_3315,N_29767,N_28437);
and UO_3316 (O_3316,N_28493,N_28959);
xnor UO_3317 (O_3317,N_29475,N_29451);
nand UO_3318 (O_3318,N_28949,N_28808);
or UO_3319 (O_3319,N_28900,N_29727);
and UO_3320 (O_3320,N_29498,N_29185);
nand UO_3321 (O_3321,N_28941,N_29471);
nand UO_3322 (O_3322,N_28553,N_29369);
xnor UO_3323 (O_3323,N_28109,N_28350);
or UO_3324 (O_3324,N_28318,N_29418);
nor UO_3325 (O_3325,N_29357,N_29406);
and UO_3326 (O_3326,N_29641,N_28785);
nand UO_3327 (O_3327,N_29924,N_29285);
xor UO_3328 (O_3328,N_28265,N_28046);
or UO_3329 (O_3329,N_28496,N_29469);
and UO_3330 (O_3330,N_29731,N_28448);
nand UO_3331 (O_3331,N_28168,N_29510);
and UO_3332 (O_3332,N_28364,N_29703);
nor UO_3333 (O_3333,N_29995,N_29893);
nand UO_3334 (O_3334,N_28281,N_29683);
nand UO_3335 (O_3335,N_28691,N_29938);
and UO_3336 (O_3336,N_29340,N_28474);
xnor UO_3337 (O_3337,N_29508,N_28678);
or UO_3338 (O_3338,N_28183,N_28429);
xnor UO_3339 (O_3339,N_29982,N_28588);
xor UO_3340 (O_3340,N_29687,N_28436);
or UO_3341 (O_3341,N_29326,N_28063);
nand UO_3342 (O_3342,N_28539,N_28724);
or UO_3343 (O_3343,N_28877,N_29041);
or UO_3344 (O_3344,N_29471,N_28310);
and UO_3345 (O_3345,N_29064,N_29808);
xor UO_3346 (O_3346,N_28127,N_29343);
nand UO_3347 (O_3347,N_29898,N_29034);
nand UO_3348 (O_3348,N_28292,N_28047);
nand UO_3349 (O_3349,N_29857,N_29766);
nor UO_3350 (O_3350,N_28343,N_29335);
or UO_3351 (O_3351,N_29480,N_28945);
or UO_3352 (O_3352,N_28287,N_29657);
xnor UO_3353 (O_3353,N_29649,N_28748);
xnor UO_3354 (O_3354,N_28664,N_29462);
or UO_3355 (O_3355,N_29921,N_29690);
or UO_3356 (O_3356,N_29636,N_28861);
or UO_3357 (O_3357,N_29891,N_28073);
nor UO_3358 (O_3358,N_28713,N_29125);
or UO_3359 (O_3359,N_29144,N_28704);
and UO_3360 (O_3360,N_28213,N_28308);
xor UO_3361 (O_3361,N_28875,N_29548);
and UO_3362 (O_3362,N_28852,N_29766);
xor UO_3363 (O_3363,N_29654,N_29247);
nor UO_3364 (O_3364,N_28541,N_29906);
nand UO_3365 (O_3365,N_28854,N_28411);
nand UO_3366 (O_3366,N_29788,N_29584);
nor UO_3367 (O_3367,N_29714,N_28444);
and UO_3368 (O_3368,N_28045,N_28508);
and UO_3369 (O_3369,N_28674,N_29481);
and UO_3370 (O_3370,N_29550,N_28324);
xor UO_3371 (O_3371,N_28283,N_28401);
nand UO_3372 (O_3372,N_29837,N_28336);
nor UO_3373 (O_3373,N_28157,N_29355);
or UO_3374 (O_3374,N_28276,N_28449);
xnor UO_3375 (O_3375,N_28883,N_29434);
nor UO_3376 (O_3376,N_28398,N_28739);
and UO_3377 (O_3377,N_29465,N_28010);
nand UO_3378 (O_3378,N_29609,N_29278);
nand UO_3379 (O_3379,N_29277,N_29088);
xnor UO_3380 (O_3380,N_29923,N_28916);
nor UO_3381 (O_3381,N_28978,N_28272);
nor UO_3382 (O_3382,N_29076,N_28232);
nor UO_3383 (O_3383,N_29862,N_28749);
nor UO_3384 (O_3384,N_29435,N_29549);
nor UO_3385 (O_3385,N_28105,N_28040);
or UO_3386 (O_3386,N_29528,N_29683);
and UO_3387 (O_3387,N_28817,N_28237);
nand UO_3388 (O_3388,N_29382,N_29366);
xnor UO_3389 (O_3389,N_29652,N_29189);
and UO_3390 (O_3390,N_28764,N_28048);
nand UO_3391 (O_3391,N_28406,N_28563);
xnor UO_3392 (O_3392,N_28774,N_28656);
nor UO_3393 (O_3393,N_28735,N_29881);
and UO_3394 (O_3394,N_28412,N_29131);
xnor UO_3395 (O_3395,N_29515,N_28688);
xnor UO_3396 (O_3396,N_28904,N_28802);
or UO_3397 (O_3397,N_29264,N_28791);
and UO_3398 (O_3398,N_29733,N_29467);
xnor UO_3399 (O_3399,N_29119,N_29690);
or UO_3400 (O_3400,N_28005,N_29744);
nand UO_3401 (O_3401,N_28597,N_28418);
or UO_3402 (O_3402,N_28906,N_28849);
nand UO_3403 (O_3403,N_28724,N_28649);
nor UO_3404 (O_3404,N_28173,N_28472);
nor UO_3405 (O_3405,N_29685,N_29994);
and UO_3406 (O_3406,N_29120,N_28392);
xnor UO_3407 (O_3407,N_28904,N_28868);
and UO_3408 (O_3408,N_28696,N_29376);
and UO_3409 (O_3409,N_29957,N_29011);
and UO_3410 (O_3410,N_28183,N_28023);
nor UO_3411 (O_3411,N_28426,N_29621);
xor UO_3412 (O_3412,N_28646,N_29483);
xor UO_3413 (O_3413,N_28335,N_29148);
or UO_3414 (O_3414,N_28028,N_29862);
nand UO_3415 (O_3415,N_28976,N_29912);
and UO_3416 (O_3416,N_28158,N_29532);
xnor UO_3417 (O_3417,N_28477,N_29393);
or UO_3418 (O_3418,N_28633,N_28530);
or UO_3419 (O_3419,N_28646,N_29589);
xnor UO_3420 (O_3420,N_29121,N_28698);
and UO_3421 (O_3421,N_29477,N_28426);
xor UO_3422 (O_3422,N_28957,N_28073);
and UO_3423 (O_3423,N_29692,N_29871);
nand UO_3424 (O_3424,N_28168,N_28497);
nor UO_3425 (O_3425,N_28175,N_29276);
xnor UO_3426 (O_3426,N_29819,N_28514);
nor UO_3427 (O_3427,N_28583,N_29749);
nor UO_3428 (O_3428,N_29339,N_29057);
or UO_3429 (O_3429,N_29108,N_29007);
nand UO_3430 (O_3430,N_29799,N_29798);
or UO_3431 (O_3431,N_29989,N_28963);
or UO_3432 (O_3432,N_28464,N_28886);
xor UO_3433 (O_3433,N_29203,N_28575);
nor UO_3434 (O_3434,N_28345,N_28185);
nor UO_3435 (O_3435,N_29599,N_28608);
nor UO_3436 (O_3436,N_29588,N_28748);
xnor UO_3437 (O_3437,N_28410,N_29887);
or UO_3438 (O_3438,N_29411,N_29648);
nand UO_3439 (O_3439,N_29860,N_28424);
or UO_3440 (O_3440,N_29915,N_29347);
xor UO_3441 (O_3441,N_29173,N_28957);
nor UO_3442 (O_3442,N_29989,N_28770);
or UO_3443 (O_3443,N_29216,N_29148);
and UO_3444 (O_3444,N_28411,N_28585);
nand UO_3445 (O_3445,N_29359,N_28036);
and UO_3446 (O_3446,N_29302,N_29532);
and UO_3447 (O_3447,N_29741,N_29983);
xnor UO_3448 (O_3448,N_29772,N_29339);
xor UO_3449 (O_3449,N_28125,N_28683);
nor UO_3450 (O_3450,N_28818,N_28553);
nand UO_3451 (O_3451,N_28859,N_28492);
nand UO_3452 (O_3452,N_28638,N_28871);
nor UO_3453 (O_3453,N_29425,N_29161);
xnor UO_3454 (O_3454,N_28537,N_28811);
xnor UO_3455 (O_3455,N_28329,N_28290);
or UO_3456 (O_3456,N_28793,N_29163);
and UO_3457 (O_3457,N_29546,N_29688);
or UO_3458 (O_3458,N_29613,N_29506);
xnor UO_3459 (O_3459,N_28407,N_29607);
nand UO_3460 (O_3460,N_29389,N_29640);
and UO_3461 (O_3461,N_29336,N_29032);
nor UO_3462 (O_3462,N_29369,N_28779);
nor UO_3463 (O_3463,N_28542,N_28167);
or UO_3464 (O_3464,N_29417,N_29450);
or UO_3465 (O_3465,N_28601,N_28396);
xnor UO_3466 (O_3466,N_28931,N_28207);
or UO_3467 (O_3467,N_28960,N_28231);
nor UO_3468 (O_3468,N_28595,N_29833);
or UO_3469 (O_3469,N_29504,N_28511);
nor UO_3470 (O_3470,N_29387,N_29893);
xnor UO_3471 (O_3471,N_28829,N_28907);
and UO_3472 (O_3472,N_29569,N_28611);
nand UO_3473 (O_3473,N_29627,N_29703);
or UO_3474 (O_3474,N_28219,N_28965);
xnor UO_3475 (O_3475,N_28235,N_29338);
and UO_3476 (O_3476,N_28421,N_28559);
xor UO_3477 (O_3477,N_29919,N_28617);
xnor UO_3478 (O_3478,N_29609,N_29180);
xor UO_3479 (O_3479,N_28439,N_28574);
nor UO_3480 (O_3480,N_29217,N_29884);
or UO_3481 (O_3481,N_29312,N_29789);
and UO_3482 (O_3482,N_29377,N_29803);
xor UO_3483 (O_3483,N_29779,N_28326);
and UO_3484 (O_3484,N_29776,N_28386);
and UO_3485 (O_3485,N_28462,N_29287);
nor UO_3486 (O_3486,N_28383,N_29702);
nor UO_3487 (O_3487,N_29792,N_29248);
xnor UO_3488 (O_3488,N_29813,N_28028);
or UO_3489 (O_3489,N_29604,N_29196);
or UO_3490 (O_3490,N_28619,N_29236);
nand UO_3491 (O_3491,N_29209,N_28713);
nor UO_3492 (O_3492,N_29956,N_28778);
nand UO_3493 (O_3493,N_28182,N_29940);
xnor UO_3494 (O_3494,N_29554,N_28896);
and UO_3495 (O_3495,N_28527,N_28584);
or UO_3496 (O_3496,N_28729,N_28444);
or UO_3497 (O_3497,N_29026,N_29939);
nor UO_3498 (O_3498,N_29409,N_29163);
and UO_3499 (O_3499,N_29846,N_28153);
endmodule