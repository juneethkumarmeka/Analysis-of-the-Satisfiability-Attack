module basic_500_3000_500_15_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_200,In_418);
and U1 (N_1,In_179,In_100);
or U2 (N_2,In_135,In_91);
nand U3 (N_3,In_244,In_103);
nand U4 (N_4,In_34,In_389);
nor U5 (N_5,In_214,In_366);
nand U6 (N_6,In_133,In_449);
and U7 (N_7,In_263,In_27);
and U8 (N_8,In_309,In_480);
nor U9 (N_9,In_481,In_232);
and U10 (N_10,In_382,In_443);
or U11 (N_11,In_196,In_437);
nand U12 (N_12,In_291,In_140);
nand U13 (N_13,In_413,In_126);
nor U14 (N_14,In_411,In_493);
and U15 (N_15,In_280,In_296);
nor U16 (N_16,In_203,In_262);
and U17 (N_17,In_99,In_221);
xnor U18 (N_18,In_304,In_465);
nor U19 (N_19,In_85,In_236);
and U20 (N_20,In_453,In_329);
and U21 (N_21,In_233,In_294);
nor U22 (N_22,In_249,In_386);
or U23 (N_23,In_312,In_79);
and U24 (N_24,In_234,In_80);
and U25 (N_25,In_384,In_485);
nor U26 (N_26,In_141,In_388);
and U27 (N_27,In_160,In_152);
and U28 (N_28,In_459,In_416);
or U29 (N_29,In_57,In_143);
nand U30 (N_30,In_295,In_467);
nand U31 (N_31,In_204,In_302);
and U32 (N_32,In_156,In_151);
or U33 (N_33,In_377,In_54);
and U34 (N_34,In_260,In_48);
or U35 (N_35,In_408,In_168);
or U36 (N_36,In_169,In_243);
or U37 (N_37,In_345,In_300);
nand U38 (N_38,In_115,In_446);
nor U39 (N_39,In_158,In_440);
or U40 (N_40,In_123,In_139);
and U41 (N_41,In_414,In_347);
and U42 (N_42,In_166,In_7);
nand U43 (N_43,In_252,In_49);
or U44 (N_44,In_201,In_466);
and U45 (N_45,In_474,In_219);
or U46 (N_46,In_438,In_44);
or U47 (N_47,In_404,In_182);
or U48 (N_48,In_318,In_239);
and U49 (N_49,In_375,In_476);
nor U50 (N_50,In_195,In_12);
nand U51 (N_51,In_484,In_487);
nor U52 (N_52,In_253,In_495);
or U53 (N_53,In_194,In_56);
nor U54 (N_54,In_87,In_489);
nor U55 (N_55,In_350,In_137);
or U56 (N_56,In_275,In_258);
nor U57 (N_57,In_469,In_316);
or U58 (N_58,In_314,In_351);
xnor U59 (N_59,In_305,In_211);
and U60 (N_60,In_72,In_266);
nand U61 (N_61,In_371,In_340);
and U62 (N_62,In_497,In_199);
nor U63 (N_63,In_146,In_272);
and U64 (N_64,In_400,In_172);
or U65 (N_65,In_349,In_149);
or U66 (N_66,In_407,In_59);
or U67 (N_67,In_421,In_401);
nand U68 (N_68,In_83,In_429);
nor U69 (N_69,In_30,In_215);
and U70 (N_70,In_282,In_251);
or U71 (N_71,In_320,In_176);
nand U72 (N_72,In_101,In_125);
xnor U73 (N_73,In_15,In_71);
nand U74 (N_74,In_220,In_207);
and U75 (N_75,In_119,In_448);
or U76 (N_76,In_35,In_120);
nand U77 (N_77,In_276,In_422);
or U78 (N_78,In_324,In_74);
nor U79 (N_79,In_230,In_257);
or U80 (N_80,In_227,In_55);
and U81 (N_81,In_150,In_372);
xnor U82 (N_82,In_97,In_228);
or U83 (N_83,In_278,In_391);
nor U84 (N_84,In_337,In_193);
nor U85 (N_85,In_14,In_483);
nor U86 (N_86,In_33,In_490);
nand U87 (N_87,In_188,In_104);
nor U88 (N_88,In_299,In_202);
or U89 (N_89,In_164,In_341);
nor U90 (N_90,In_23,In_353);
nand U91 (N_91,In_468,In_310);
nand U92 (N_92,In_147,In_477);
nand U93 (N_93,In_167,In_6);
and U94 (N_94,In_430,In_267);
and U95 (N_95,In_105,In_82);
nor U96 (N_96,In_297,In_491);
nand U97 (N_97,In_197,In_464);
and U98 (N_98,In_110,In_406);
nor U99 (N_99,In_362,In_245);
or U100 (N_100,In_261,In_129);
xor U101 (N_101,In_315,In_292);
or U102 (N_102,In_248,In_18);
nor U103 (N_103,In_289,In_1);
nor U104 (N_104,In_136,In_361);
or U105 (N_105,In_383,In_369);
nand U106 (N_106,In_427,In_183);
nor U107 (N_107,In_321,In_445);
and U108 (N_108,In_360,In_235);
and U109 (N_109,In_488,In_281);
or U110 (N_110,In_387,In_352);
nand U111 (N_111,In_417,In_118);
or U112 (N_112,In_162,In_475);
nand U113 (N_113,In_165,In_394);
nand U114 (N_114,In_271,In_333);
and U115 (N_115,In_43,In_94);
and U116 (N_116,In_61,In_58);
nor U117 (N_117,In_303,In_277);
or U118 (N_118,In_51,In_113);
nor U119 (N_119,In_462,In_247);
nor U120 (N_120,In_279,In_45);
nand U121 (N_121,In_157,In_460);
nand U122 (N_122,In_81,In_67);
and U123 (N_123,In_225,In_38);
or U124 (N_124,In_98,In_50);
nor U125 (N_125,In_210,In_308);
nor U126 (N_126,In_36,In_37);
and U127 (N_127,In_171,In_128);
and U128 (N_128,In_175,In_287);
nor U129 (N_129,In_288,In_216);
nand U130 (N_130,In_224,In_301);
or U131 (N_131,In_395,In_191);
nor U132 (N_132,In_451,In_26);
or U133 (N_133,In_356,In_174);
and U134 (N_134,In_223,In_492);
nor U135 (N_135,In_264,In_397);
or U136 (N_136,In_189,In_250);
and U137 (N_137,In_2,In_322);
and U138 (N_138,In_454,In_330);
xor U139 (N_139,In_425,In_90);
nor U140 (N_140,In_131,In_381);
or U141 (N_141,In_355,In_270);
or U142 (N_142,In_335,In_66);
nor U143 (N_143,In_117,In_238);
nor U144 (N_144,In_364,In_10);
or U145 (N_145,In_86,In_457);
or U146 (N_146,In_205,In_432);
nor U147 (N_147,In_265,In_499);
nand U148 (N_148,In_285,In_92);
nand U149 (N_149,In_69,In_343);
and U150 (N_150,In_76,In_284);
nor U151 (N_151,In_28,In_331);
or U152 (N_152,In_319,In_415);
and U153 (N_153,In_231,In_374);
nand U154 (N_154,In_431,In_269);
nor U155 (N_155,In_112,In_392);
nor U156 (N_156,In_471,In_463);
and U157 (N_157,In_478,In_144);
nor U158 (N_158,In_461,In_63);
or U159 (N_159,In_19,In_134);
nand U160 (N_160,In_246,In_9);
nor U161 (N_161,In_93,In_5);
nor U162 (N_162,In_102,In_426);
or U163 (N_163,In_357,In_84);
and U164 (N_164,In_428,In_111);
nor U165 (N_165,In_209,In_452);
and U166 (N_166,In_89,In_254);
nor U167 (N_167,In_178,In_218);
and U168 (N_168,In_52,In_479);
and U169 (N_169,In_379,In_154);
nand U170 (N_170,In_0,In_336);
nor U171 (N_171,In_42,In_420);
nand U172 (N_172,In_198,In_456);
nand U173 (N_173,In_273,In_241);
and U174 (N_174,In_313,In_450);
or U175 (N_175,In_46,In_433);
nand U176 (N_176,In_393,In_402);
or U177 (N_177,In_325,In_328);
nand U178 (N_178,In_334,In_368);
and U179 (N_179,In_3,In_217);
nand U180 (N_180,In_494,In_41);
or U181 (N_181,In_403,In_16);
nor U182 (N_182,In_96,In_208);
nand U183 (N_183,In_121,In_177);
and U184 (N_184,In_436,In_181);
or U185 (N_185,In_185,In_434);
nor U186 (N_186,In_163,In_354);
nor U187 (N_187,In_65,In_290);
nand U188 (N_188,In_222,In_73);
nor U189 (N_189,In_106,In_109);
nor U190 (N_190,In_286,In_373);
nand U191 (N_191,In_8,In_323);
or U192 (N_192,In_419,In_255);
or U193 (N_193,In_4,In_206);
nand U194 (N_194,In_13,In_127);
and U195 (N_195,In_95,In_486);
nor U196 (N_196,In_25,In_229);
nand U197 (N_197,In_439,In_317);
nor U198 (N_198,In_47,In_180);
xor U199 (N_199,In_107,In_70);
or U200 (N_200,In_20,N_84);
or U201 (N_201,N_148,N_101);
and U202 (N_202,In_145,N_20);
nand U203 (N_203,N_146,N_87);
and U204 (N_204,In_142,N_49);
nand U205 (N_205,In_424,In_412);
or U206 (N_206,In_256,In_344);
nand U207 (N_207,N_182,N_193);
and U208 (N_208,N_11,N_110);
or U209 (N_209,In_380,N_39);
nand U210 (N_210,N_57,N_3);
or U211 (N_211,N_134,In_396);
nand U212 (N_212,N_192,In_75);
nand U213 (N_213,N_109,In_132);
nand U214 (N_214,N_119,In_17);
nor U215 (N_215,N_53,N_33);
nor U216 (N_216,N_77,N_198);
and U217 (N_217,N_56,N_25);
nand U218 (N_218,N_183,N_23);
nor U219 (N_219,N_105,In_153);
nor U220 (N_220,In_268,N_165);
xor U221 (N_221,In_21,N_122);
or U222 (N_222,N_79,In_148);
or U223 (N_223,In_186,N_75);
or U224 (N_224,N_12,In_306);
nand U225 (N_225,N_114,N_47);
nand U226 (N_226,N_136,N_97);
xnor U227 (N_227,In_358,N_6);
or U228 (N_228,In_458,N_14);
and U229 (N_229,N_70,In_410);
and U230 (N_230,N_85,In_442);
nand U231 (N_231,N_178,N_13);
or U232 (N_232,In_365,In_242);
or U233 (N_233,N_113,N_120);
nor U234 (N_234,N_132,In_240);
or U235 (N_235,N_52,N_65);
and U236 (N_236,N_155,N_115);
nor U237 (N_237,N_4,In_399);
and U238 (N_238,N_126,N_187);
or U239 (N_239,N_8,N_141);
nor U240 (N_240,In_327,N_22);
or U241 (N_241,N_83,N_43);
and U242 (N_242,N_30,N_177);
nor U243 (N_243,N_194,N_55);
nand U244 (N_244,N_94,N_157);
nand U245 (N_245,N_104,N_166);
nor U246 (N_246,N_171,N_59);
nor U247 (N_247,N_44,In_68);
or U248 (N_248,N_27,In_390);
nor U249 (N_249,N_176,N_17);
or U250 (N_250,N_159,N_153);
nand U251 (N_251,N_93,N_123);
xor U252 (N_252,N_156,In_114);
or U253 (N_253,In_482,N_31);
nand U254 (N_254,N_127,N_48);
and U255 (N_255,N_175,N_139);
and U256 (N_256,In_116,In_11);
nand U257 (N_257,N_71,In_122);
nor U258 (N_258,N_181,N_89);
or U259 (N_259,N_32,In_363);
nand U260 (N_260,N_9,N_143);
and U261 (N_261,In_138,N_131);
or U262 (N_262,In_338,N_106);
nor U263 (N_263,N_138,N_66);
nor U264 (N_264,In_259,In_124);
nor U265 (N_265,N_18,N_158);
nand U266 (N_266,N_111,N_0);
nand U267 (N_267,In_64,N_160);
xnor U268 (N_268,In_24,N_149);
or U269 (N_269,N_98,N_170);
nor U270 (N_270,N_99,In_346);
nand U271 (N_271,N_189,N_86);
nand U272 (N_272,In_40,In_32);
and U273 (N_273,N_144,N_169);
and U274 (N_274,In_184,In_237);
nor U275 (N_275,In_370,N_10);
xor U276 (N_276,N_26,N_15);
or U277 (N_277,N_135,In_409);
or U278 (N_278,N_161,N_38);
or U279 (N_279,In_274,N_37);
xor U280 (N_280,N_167,N_80);
or U281 (N_281,N_191,In_78);
and U282 (N_282,N_34,In_441);
nor U283 (N_283,N_96,In_326);
nand U284 (N_284,In_339,N_41);
and U285 (N_285,In_378,N_54);
or U286 (N_286,In_192,In_444);
or U287 (N_287,N_62,N_7);
and U288 (N_288,N_173,N_174);
or U289 (N_289,N_117,In_173);
nor U290 (N_290,N_164,N_142);
nor U291 (N_291,In_342,N_112);
or U292 (N_292,N_19,In_447);
nor U293 (N_293,N_64,N_67);
nor U294 (N_294,N_128,N_107);
nor U295 (N_295,In_39,N_147);
or U296 (N_296,N_151,N_133);
or U297 (N_297,In_159,N_68);
nand U298 (N_298,In_332,In_348);
nand U299 (N_299,N_190,N_199);
and U300 (N_300,N_129,In_293);
or U301 (N_301,N_90,In_472);
or U302 (N_302,N_150,N_35);
nor U303 (N_303,N_145,N_121);
and U304 (N_304,In_283,N_50);
and U305 (N_305,N_184,N_2);
and U306 (N_306,In_496,N_172);
nor U307 (N_307,N_103,N_180);
nor U308 (N_308,N_73,N_168);
and U309 (N_309,N_95,In_423);
nand U310 (N_310,N_81,N_188);
nand U311 (N_311,N_116,N_179);
and U312 (N_312,N_100,N_5);
nand U313 (N_313,N_195,In_405);
or U314 (N_314,In_359,In_470);
and U315 (N_315,In_435,N_40);
or U316 (N_316,N_61,In_473);
nor U317 (N_317,In_62,In_77);
or U318 (N_318,N_46,In_455);
nand U319 (N_319,In_376,N_163);
and U320 (N_320,N_196,In_53);
xor U321 (N_321,In_187,N_36);
or U322 (N_322,N_74,In_498);
or U323 (N_323,N_137,N_45);
and U324 (N_324,N_92,N_21);
or U325 (N_325,N_186,In_213);
nor U326 (N_326,In_31,In_88);
nand U327 (N_327,N_82,In_29);
nand U328 (N_328,N_124,In_130);
nor U329 (N_329,In_22,N_108);
nand U330 (N_330,N_140,N_29);
or U331 (N_331,N_1,In_161);
nand U332 (N_332,N_51,N_162);
nand U333 (N_333,N_91,In_155);
and U334 (N_334,In_311,N_154);
nand U335 (N_335,N_185,In_170);
xor U336 (N_336,In_385,N_42);
nand U337 (N_337,In_60,N_102);
nor U338 (N_338,In_398,In_108);
and U339 (N_339,In_298,N_88);
nor U340 (N_340,N_60,N_63);
or U341 (N_341,N_118,In_307);
or U342 (N_342,N_28,In_367);
nand U343 (N_343,N_76,N_16);
nor U344 (N_344,N_78,N_69);
or U345 (N_345,In_190,In_212);
or U346 (N_346,N_24,N_152);
or U347 (N_347,N_72,N_58);
nand U348 (N_348,N_197,N_125);
and U349 (N_349,N_130,In_226);
and U350 (N_350,N_153,N_113);
nand U351 (N_351,N_111,In_399);
or U352 (N_352,In_259,N_117);
or U353 (N_353,In_256,N_136);
or U354 (N_354,N_36,In_367);
or U355 (N_355,In_226,N_71);
or U356 (N_356,N_123,N_59);
nor U357 (N_357,In_259,N_81);
nor U358 (N_358,In_410,In_116);
xor U359 (N_359,N_155,In_64);
nand U360 (N_360,In_190,N_195);
nor U361 (N_361,In_441,N_158);
nand U362 (N_362,N_82,In_237);
or U363 (N_363,In_259,N_136);
nor U364 (N_364,In_458,N_119);
and U365 (N_365,N_190,N_113);
nand U366 (N_366,In_108,In_447);
and U367 (N_367,N_69,In_31);
nand U368 (N_368,In_240,In_385);
and U369 (N_369,N_59,In_363);
and U370 (N_370,In_472,In_242);
nand U371 (N_371,N_100,N_143);
xnor U372 (N_372,In_306,N_52);
or U373 (N_373,N_106,N_133);
nor U374 (N_374,N_56,In_78);
nor U375 (N_375,In_326,N_143);
nand U376 (N_376,N_2,N_21);
and U377 (N_377,N_176,N_196);
nor U378 (N_378,N_65,In_268);
or U379 (N_379,N_5,In_142);
and U380 (N_380,N_16,N_142);
nor U381 (N_381,N_128,In_326);
or U382 (N_382,In_75,In_122);
or U383 (N_383,In_124,In_298);
nor U384 (N_384,N_154,N_100);
or U385 (N_385,N_24,In_307);
nand U386 (N_386,In_130,N_186);
nor U387 (N_387,In_370,N_158);
nor U388 (N_388,N_157,N_23);
or U389 (N_389,N_95,N_89);
or U390 (N_390,N_49,In_358);
or U391 (N_391,In_423,N_169);
nor U392 (N_392,N_164,N_160);
nand U393 (N_393,N_194,N_80);
nor U394 (N_394,N_108,N_73);
nand U395 (N_395,N_66,N_94);
or U396 (N_396,N_56,N_63);
or U397 (N_397,N_13,In_412);
nor U398 (N_398,N_19,N_174);
nand U399 (N_399,N_102,N_31);
or U400 (N_400,N_296,N_305);
or U401 (N_401,N_205,N_304);
nor U402 (N_402,N_203,N_387);
nor U403 (N_403,N_307,N_301);
or U404 (N_404,N_397,N_264);
nand U405 (N_405,N_204,N_249);
and U406 (N_406,N_314,N_270);
nand U407 (N_407,N_297,N_321);
and U408 (N_408,N_347,N_200);
and U409 (N_409,N_219,N_253);
or U410 (N_410,N_309,N_280);
nor U411 (N_411,N_241,N_386);
nand U412 (N_412,N_247,N_229);
nor U413 (N_413,N_266,N_260);
and U414 (N_414,N_306,N_292);
and U415 (N_415,N_256,N_371);
nor U416 (N_416,N_238,N_283);
nand U417 (N_417,N_245,N_394);
or U418 (N_418,N_393,N_272);
and U419 (N_419,N_202,N_355);
and U420 (N_420,N_322,N_334);
nor U421 (N_421,N_366,N_230);
nor U422 (N_422,N_330,N_285);
nor U423 (N_423,N_207,N_348);
nor U424 (N_424,N_251,N_328);
or U425 (N_425,N_233,N_237);
and U426 (N_426,N_317,N_399);
and U427 (N_427,N_224,N_212);
and U428 (N_428,N_290,N_255);
and U429 (N_429,N_345,N_268);
or U430 (N_430,N_375,N_263);
nor U431 (N_431,N_385,N_356);
and U432 (N_432,N_335,N_396);
and U433 (N_433,N_358,N_392);
and U434 (N_434,N_242,N_332);
nand U435 (N_435,N_395,N_300);
or U436 (N_436,N_370,N_228);
and U437 (N_437,N_338,N_291);
or U438 (N_438,N_352,N_248);
and U439 (N_439,N_362,N_384);
nand U440 (N_440,N_258,N_302);
xnor U441 (N_441,N_380,N_210);
or U442 (N_442,N_331,N_326);
and U443 (N_443,N_226,N_252);
nor U444 (N_444,N_214,N_350);
nor U445 (N_445,N_367,N_372);
xnor U446 (N_446,N_340,N_343);
and U447 (N_447,N_286,N_262);
nor U448 (N_448,N_299,N_231);
xnor U449 (N_449,N_303,N_379);
and U450 (N_450,N_254,N_389);
or U451 (N_451,N_383,N_312);
nand U452 (N_452,N_323,N_341);
and U453 (N_453,N_276,N_381);
and U454 (N_454,N_261,N_209);
or U455 (N_455,N_277,N_320);
and U456 (N_456,N_329,N_391);
and U457 (N_457,N_227,N_208);
nor U458 (N_458,N_271,N_222);
nand U459 (N_459,N_333,N_374);
and U460 (N_460,N_315,N_287);
nand U461 (N_461,N_310,N_278);
and U462 (N_462,N_308,N_239);
and U463 (N_463,N_357,N_243);
or U464 (N_464,N_295,N_319);
nor U465 (N_465,N_279,N_311);
and U466 (N_466,N_388,N_217);
nand U467 (N_467,N_339,N_235);
or U468 (N_468,N_225,N_349);
and U469 (N_469,N_382,N_346);
and U470 (N_470,N_359,N_267);
or U471 (N_471,N_365,N_259);
nand U472 (N_472,N_234,N_223);
nor U473 (N_473,N_363,N_216);
xor U474 (N_474,N_289,N_316);
or U475 (N_475,N_294,N_327);
nor U476 (N_476,N_274,N_273);
nand U477 (N_477,N_213,N_232);
nand U478 (N_478,N_344,N_220);
and U479 (N_479,N_282,N_373);
and U480 (N_480,N_257,N_390);
and U481 (N_481,N_281,N_361);
or U482 (N_482,N_201,N_215);
nand U483 (N_483,N_398,N_211);
or U484 (N_484,N_325,N_250);
nor U485 (N_485,N_376,N_369);
or U486 (N_486,N_377,N_313);
nor U487 (N_487,N_351,N_269);
or U488 (N_488,N_246,N_360);
and U489 (N_489,N_364,N_337);
xnor U490 (N_490,N_378,N_293);
and U491 (N_491,N_265,N_288);
nand U492 (N_492,N_221,N_342);
xnor U493 (N_493,N_318,N_284);
nand U494 (N_494,N_236,N_298);
nor U495 (N_495,N_324,N_275);
and U496 (N_496,N_353,N_206);
and U497 (N_497,N_244,N_240);
nor U498 (N_498,N_336,N_354);
nand U499 (N_499,N_218,N_368);
or U500 (N_500,N_221,N_371);
nor U501 (N_501,N_298,N_303);
and U502 (N_502,N_227,N_329);
nor U503 (N_503,N_285,N_205);
or U504 (N_504,N_307,N_232);
or U505 (N_505,N_251,N_211);
nor U506 (N_506,N_342,N_329);
nand U507 (N_507,N_362,N_255);
and U508 (N_508,N_377,N_200);
and U509 (N_509,N_234,N_348);
nand U510 (N_510,N_314,N_292);
or U511 (N_511,N_329,N_350);
nand U512 (N_512,N_326,N_274);
and U513 (N_513,N_346,N_213);
and U514 (N_514,N_205,N_392);
and U515 (N_515,N_277,N_250);
and U516 (N_516,N_351,N_297);
and U517 (N_517,N_387,N_242);
and U518 (N_518,N_387,N_265);
or U519 (N_519,N_286,N_205);
nand U520 (N_520,N_321,N_324);
nor U521 (N_521,N_320,N_200);
or U522 (N_522,N_315,N_265);
and U523 (N_523,N_235,N_223);
or U524 (N_524,N_367,N_351);
or U525 (N_525,N_391,N_292);
nand U526 (N_526,N_277,N_358);
or U527 (N_527,N_353,N_393);
and U528 (N_528,N_217,N_350);
or U529 (N_529,N_230,N_308);
nor U530 (N_530,N_268,N_239);
xnor U531 (N_531,N_247,N_281);
nor U532 (N_532,N_256,N_213);
and U533 (N_533,N_268,N_204);
and U534 (N_534,N_309,N_207);
or U535 (N_535,N_293,N_258);
nand U536 (N_536,N_335,N_270);
or U537 (N_537,N_235,N_270);
nor U538 (N_538,N_309,N_314);
nand U539 (N_539,N_345,N_395);
or U540 (N_540,N_340,N_381);
nor U541 (N_541,N_377,N_309);
nand U542 (N_542,N_246,N_253);
nand U543 (N_543,N_334,N_237);
nor U544 (N_544,N_207,N_303);
nand U545 (N_545,N_370,N_259);
and U546 (N_546,N_332,N_200);
or U547 (N_547,N_330,N_311);
and U548 (N_548,N_237,N_234);
nor U549 (N_549,N_285,N_243);
nand U550 (N_550,N_379,N_287);
nand U551 (N_551,N_327,N_356);
nor U552 (N_552,N_399,N_308);
nor U553 (N_553,N_331,N_267);
nor U554 (N_554,N_348,N_375);
and U555 (N_555,N_264,N_298);
and U556 (N_556,N_318,N_313);
and U557 (N_557,N_228,N_344);
nand U558 (N_558,N_240,N_209);
and U559 (N_559,N_304,N_342);
and U560 (N_560,N_376,N_323);
and U561 (N_561,N_310,N_288);
nand U562 (N_562,N_225,N_286);
nor U563 (N_563,N_216,N_383);
nor U564 (N_564,N_373,N_302);
or U565 (N_565,N_318,N_293);
nand U566 (N_566,N_203,N_327);
nand U567 (N_567,N_340,N_385);
and U568 (N_568,N_360,N_359);
or U569 (N_569,N_357,N_387);
or U570 (N_570,N_378,N_299);
and U571 (N_571,N_363,N_267);
nand U572 (N_572,N_322,N_288);
and U573 (N_573,N_371,N_203);
nand U574 (N_574,N_386,N_276);
or U575 (N_575,N_301,N_296);
and U576 (N_576,N_279,N_211);
and U577 (N_577,N_313,N_254);
nor U578 (N_578,N_286,N_245);
or U579 (N_579,N_380,N_204);
nor U580 (N_580,N_323,N_207);
nand U581 (N_581,N_272,N_274);
nand U582 (N_582,N_306,N_323);
and U583 (N_583,N_212,N_369);
and U584 (N_584,N_247,N_236);
nor U585 (N_585,N_220,N_380);
nor U586 (N_586,N_203,N_284);
and U587 (N_587,N_279,N_381);
and U588 (N_588,N_207,N_374);
nand U589 (N_589,N_313,N_300);
or U590 (N_590,N_240,N_273);
and U591 (N_591,N_258,N_237);
nor U592 (N_592,N_325,N_311);
nand U593 (N_593,N_388,N_301);
or U594 (N_594,N_346,N_324);
nor U595 (N_595,N_316,N_339);
nor U596 (N_596,N_330,N_277);
or U597 (N_597,N_337,N_392);
nand U598 (N_598,N_263,N_304);
nand U599 (N_599,N_335,N_274);
or U600 (N_600,N_446,N_401);
nor U601 (N_601,N_519,N_518);
nor U602 (N_602,N_570,N_591);
nand U603 (N_603,N_583,N_474);
nand U604 (N_604,N_454,N_440);
nor U605 (N_605,N_433,N_434);
or U606 (N_606,N_540,N_409);
and U607 (N_607,N_595,N_414);
nor U608 (N_608,N_533,N_564);
nor U609 (N_609,N_491,N_547);
and U610 (N_610,N_527,N_508);
nor U611 (N_611,N_456,N_435);
nor U612 (N_612,N_539,N_457);
or U613 (N_613,N_438,N_576);
nand U614 (N_614,N_526,N_536);
and U615 (N_615,N_571,N_530);
or U616 (N_616,N_534,N_580);
and U617 (N_617,N_575,N_509);
or U618 (N_618,N_554,N_562);
or U619 (N_619,N_579,N_480);
or U620 (N_620,N_450,N_555);
and U621 (N_621,N_402,N_451);
nand U622 (N_622,N_411,N_468);
and U623 (N_623,N_592,N_478);
nor U624 (N_624,N_462,N_475);
and U625 (N_625,N_502,N_432);
nor U626 (N_626,N_546,N_460);
or U627 (N_627,N_593,N_514);
nor U628 (N_628,N_485,N_493);
nor U629 (N_629,N_560,N_503);
nand U630 (N_630,N_543,N_447);
nand U631 (N_631,N_467,N_538);
nand U632 (N_632,N_558,N_515);
or U633 (N_633,N_477,N_511);
or U634 (N_634,N_582,N_531);
and U635 (N_635,N_469,N_429);
nand U636 (N_636,N_501,N_537);
and U637 (N_637,N_415,N_466);
nand U638 (N_638,N_542,N_507);
and U639 (N_639,N_492,N_461);
and U640 (N_640,N_463,N_528);
nand U641 (N_641,N_529,N_541);
or U642 (N_642,N_489,N_589);
or U643 (N_643,N_594,N_445);
nor U644 (N_644,N_545,N_471);
nor U645 (N_645,N_506,N_407);
and U646 (N_646,N_520,N_586);
nand U647 (N_647,N_522,N_439);
or U648 (N_648,N_549,N_500);
and U649 (N_649,N_421,N_452);
nor U650 (N_650,N_426,N_431);
or U651 (N_651,N_557,N_585);
and U652 (N_652,N_524,N_479);
nand U653 (N_653,N_568,N_486);
nand U654 (N_654,N_550,N_484);
and U655 (N_655,N_494,N_517);
or U656 (N_656,N_416,N_443);
nand U657 (N_657,N_470,N_553);
nor U658 (N_658,N_504,N_598);
nand U659 (N_659,N_510,N_563);
nand U660 (N_660,N_472,N_430);
and U661 (N_661,N_497,N_490);
and U662 (N_662,N_496,N_476);
and U663 (N_663,N_464,N_544);
and U664 (N_664,N_404,N_488);
and U665 (N_665,N_577,N_423);
and U666 (N_666,N_495,N_551);
nand U667 (N_667,N_444,N_573);
xnor U668 (N_668,N_513,N_561);
and U669 (N_669,N_574,N_588);
nand U670 (N_670,N_556,N_448);
nand U671 (N_671,N_532,N_425);
nor U672 (N_672,N_482,N_597);
nand U673 (N_673,N_596,N_420);
nor U674 (N_674,N_442,N_428);
nand U675 (N_675,N_459,N_400);
or U676 (N_676,N_405,N_566);
nor U677 (N_677,N_406,N_412);
or U678 (N_678,N_584,N_599);
and U679 (N_679,N_552,N_413);
nand U680 (N_680,N_572,N_523);
nor U681 (N_681,N_473,N_465);
nand U682 (N_682,N_516,N_505);
nand U683 (N_683,N_449,N_424);
or U684 (N_684,N_487,N_483);
or U685 (N_685,N_569,N_565);
and U686 (N_686,N_419,N_436);
and U687 (N_687,N_567,N_418);
and U688 (N_688,N_548,N_403);
xnor U689 (N_689,N_455,N_408);
nor U690 (N_690,N_559,N_427);
nor U691 (N_691,N_521,N_437);
nor U692 (N_692,N_512,N_587);
and U693 (N_693,N_422,N_535);
nor U694 (N_694,N_410,N_578);
xnor U695 (N_695,N_417,N_458);
or U696 (N_696,N_481,N_581);
and U697 (N_697,N_498,N_453);
or U698 (N_698,N_525,N_499);
nand U699 (N_699,N_441,N_590);
nand U700 (N_700,N_418,N_513);
or U701 (N_701,N_492,N_459);
and U702 (N_702,N_402,N_415);
and U703 (N_703,N_457,N_456);
xor U704 (N_704,N_484,N_555);
and U705 (N_705,N_482,N_537);
or U706 (N_706,N_535,N_568);
nand U707 (N_707,N_552,N_495);
nand U708 (N_708,N_475,N_469);
or U709 (N_709,N_453,N_443);
and U710 (N_710,N_499,N_510);
or U711 (N_711,N_554,N_592);
and U712 (N_712,N_550,N_405);
xnor U713 (N_713,N_454,N_449);
xor U714 (N_714,N_413,N_468);
nor U715 (N_715,N_454,N_529);
or U716 (N_716,N_542,N_501);
or U717 (N_717,N_582,N_522);
or U718 (N_718,N_514,N_595);
nand U719 (N_719,N_413,N_509);
and U720 (N_720,N_455,N_562);
nand U721 (N_721,N_572,N_479);
nor U722 (N_722,N_440,N_530);
nor U723 (N_723,N_583,N_418);
and U724 (N_724,N_468,N_446);
or U725 (N_725,N_496,N_515);
nor U726 (N_726,N_427,N_537);
or U727 (N_727,N_563,N_553);
nor U728 (N_728,N_585,N_437);
or U729 (N_729,N_446,N_510);
nor U730 (N_730,N_567,N_545);
nand U731 (N_731,N_473,N_464);
nand U732 (N_732,N_549,N_410);
and U733 (N_733,N_585,N_486);
nor U734 (N_734,N_472,N_553);
or U735 (N_735,N_439,N_469);
nor U736 (N_736,N_532,N_595);
nor U737 (N_737,N_455,N_501);
or U738 (N_738,N_468,N_428);
nand U739 (N_739,N_520,N_446);
nor U740 (N_740,N_437,N_431);
nor U741 (N_741,N_502,N_538);
nor U742 (N_742,N_546,N_406);
nor U743 (N_743,N_478,N_483);
nand U744 (N_744,N_587,N_416);
or U745 (N_745,N_483,N_579);
or U746 (N_746,N_589,N_454);
or U747 (N_747,N_442,N_571);
or U748 (N_748,N_450,N_504);
nand U749 (N_749,N_449,N_537);
nor U750 (N_750,N_510,N_541);
xor U751 (N_751,N_519,N_572);
or U752 (N_752,N_483,N_501);
nor U753 (N_753,N_549,N_595);
xor U754 (N_754,N_599,N_466);
and U755 (N_755,N_510,N_487);
nand U756 (N_756,N_487,N_545);
nor U757 (N_757,N_559,N_551);
xor U758 (N_758,N_486,N_407);
or U759 (N_759,N_475,N_451);
nor U760 (N_760,N_401,N_513);
nand U761 (N_761,N_549,N_559);
nand U762 (N_762,N_537,N_452);
and U763 (N_763,N_494,N_552);
or U764 (N_764,N_571,N_523);
nor U765 (N_765,N_400,N_552);
or U766 (N_766,N_444,N_586);
or U767 (N_767,N_566,N_515);
nor U768 (N_768,N_594,N_498);
nand U769 (N_769,N_415,N_509);
nand U770 (N_770,N_414,N_515);
or U771 (N_771,N_595,N_513);
and U772 (N_772,N_419,N_402);
and U773 (N_773,N_592,N_528);
and U774 (N_774,N_444,N_539);
nor U775 (N_775,N_428,N_476);
or U776 (N_776,N_587,N_441);
nand U777 (N_777,N_430,N_578);
nand U778 (N_778,N_587,N_499);
and U779 (N_779,N_519,N_466);
nor U780 (N_780,N_568,N_589);
nand U781 (N_781,N_446,N_478);
nand U782 (N_782,N_527,N_432);
nor U783 (N_783,N_502,N_436);
or U784 (N_784,N_582,N_447);
nand U785 (N_785,N_526,N_559);
or U786 (N_786,N_455,N_561);
and U787 (N_787,N_401,N_487);
or U788 (N_788,N_589,N_595);
nor U789 (N_789,N_565,N_464);
xor U790 (N_790,N_567,N_477);
nor U791 (N_791,N_481,N_443);
and U792 (N_792,N_537,N_504);
or U793 (N_793,N_534,N_469);
nand U794 (N_794,N_547,N_503);
nor U795 (N_795,N_572,N_401);
and U796 (N_796,N_584,N_535);
nand U797 (N_797,N_435,N_497);
or U798 (N_798,N_481,N_473);
nand U799 (N_799,N_442,N_492);
and U800 (N_800,N_631,N_658);
or U801 (N_801,N_627,N_669);
nor U802 (N_802,N_655,N_661);
and U803 (N_803,N_788,N_608);
and U804 (N_804,N_626,N_730);
or U805 (N_805,N_664,N_654);
nand U806 (N_806,N_764,N_671);
or U807 (N_807,N_681,N_614);
nand U808 (N_808,N_683,N_732);
xor U809 (N_809,N_686,N_757);
xor U810 (N_810,N_635,N_715);
and U811 (N_811,N_691,N_756);
nor U812 (N_812,N_697,N_785);
or U813 (N_813,N_659,N_620);
and U814 (N_814,N_721,N_679);
xor U815 (N_815,N_607,N_726);
xor U816 (N_816,N_769,N_710);
nor U817 (N_817,N_616,N_653);
or U818 (N_818,N_703,N_676);
nor U819 (N_819,N_656,N_753);
nor U820 (N_820,N_749,N_624);
and U821 (N_821,N_644,N_690);
or U822 (N_822,N_763,N_602);
and U823 (N_823,N_734,N_634);
nand U824 (N_824,N_613,N_706);
nor U825 (N_825,N_696,N_748);
nor U826 (N_826,N_792,N_758);
nand U827 (N_827,N_695,N_615);
or U828 (N_828,N_707,N_724);
and U829 (N_829,N_688,N_633);
xor U830 (N_830,N_733,N_740);
xnor U831 (N_831,N_651,N_713);
nand U832 (N_832,N_791,N_719);
nand U833 (N_833,N_781,N_742);
or U834 (N_834,N_760,N_660);
nor U835 (N_835,N_657,N_702);
nor U836 (N_836,N_622,N_650);
nand U837 (N_837,N_762,N_798);
and U838 (N_838,N_725,N_637);
and U839 (N_839,N_708,N_663);
and U840 (N_840,N_797,N_623);
and U841 (N_841,N_646,N_766);
or U842 (N_842,N_630,N_772);
nand U843 (N_843,N_744,N_793);
or U844 (N_844,N_723,N_776);
nand U845 (N_845,N_773,N_771);
and U846 (N_846,N_639,N_751);
nor U847 (N_847,N_611,N_605);
and U848 (N_848,N_752,N_712);
nand U849 (N_849,N_689,N_648);
nor U850 (N_850,N_778,N_665);
nor U851 (N_851,N_684,N_794);
nor U852 (N_852,N_728,N_694);
nor U853 (N_853,N_700,N_632);
nand U854 (N_854,N_601,N_609);
or U855 (N_855,N_625,N_698);
and U856 (N_856,N_612,N_674);
or U857 (N_857,N_722,N_747);
or U858 (N_858,N_704,N_600);
or U859 (N_859,N_685,N_768);
and U860 (N_860,N_693,N_666);
nand U861 (N_861,N_714,N_606);
or U862 (N_862,N_770,N_617);
nand U863 (N_863,N_692,N_652);
or U864 (N_864,N_699,N_731);
nor U865 (N_865,N_672,N_750);
nor U866 (N_866,N_717,N_636);
nor U867 (N_867,N_799,N_619);
or U868 (N_868,N_711,N_640);
and U869 (N_869,N_739,N_643);
nand U870 (N_870,N_662,N_735);
nor U871 (N_871,N_610,N_796);
nor U872 (N_872,N_754,N_774);
or U873 (N_873,N_787,N_784);
nand U874 (N_874,N_677,N_705);
and U875 (N_875,N_737,N_729);
and U876 (N_876,N_628,N_777);
nand U877 (N_877,N_645,N_775);
nand U878 (N_878,N_789,N_783);
nor U879 (N_879,N_746,N_668);
and U880 (N_880,N_604,N_701);
nor U881 (N_881,N_673,N_649);
or U882 (N_882,N_720,N_761);
nor U883 (N_883,N_641,N_642);
nor U884 (N_884,N_718,N_782);
nor U885 (N_885,N_743,N_727);
nor U886 (N_886,N_786,N_741);
nand U887 (N_887,N_618,N_795);
or U888 (N_888,N_755,N_647);
and U889 (N_889,N_621,N_736);
nor U890 (N_890,N_678,N_687);
or U891 (N_891,N_716,N_790);
nor U892 (N_892,N_682,N_603);
nand U893 (N_893,N_675,N_765);
or U894 (N_894,N_759,N_638);
nor U895 (N_895,N_670,N_629);
and U896 (N_896,N_738,N_745);
and U897 (N_897,N_680,N_709);
or U898 (N_898,N_667,N_779);
or U899 (N_899,N_767,N_780);
or U900 (N_900,N_689,N_711);
or U901 (N_901,N_646,N_758);
and U902 (N_902,N_618,N_652);
and U903 (N_903,N_643,N_651);
or U904 (N_904,N_794,N_647);
nand U905 (N_905,N_653,N_697);
or U906 (N_906,N_710,N_714);
and U907 (N_907,N_668,N_642);
and U908 (N_908,N_666,N_742);
or U909 (N_909,N_657,N_611);
and U910 (N_910,N_766,N_645);
nand U911 (N_911,N_623,N_609);
nand U912 (N_912,N_618,N_783);
or U913 (N_913,N_624,N_797);
and U914 (N_914,N_664,N_695);
and U915 (N_915,N_745,N_754);
and U916 (N_916,N_769,N_653);
nand U917 (N_917,N_764,N_684);
nand U918 (N_918,N_688,N_634);
nand U919 (N_919,N_616,N_657);
or U920 (N_920,N_603,N_639);
and U921 (N_921,N_635,N_704);
or U922 (N_922,N_751,N_706);
nand U923 (N_923,N_697,N_726);
and U924 (N_924,N_676,N_614);
and U925 (N_925,N_648,N_772);
and U926 (N_926,N_783,N_745);
nand U927 (N_927,N_749,N_787);
and U928 (N_928,N_716,N_784);
or U929 (N_929,N_631,N_647);
or U930 (N_930,N_621,N_645);
or U931 (N_931,N_708,N_627);
and U932 (N_932,N_670,N_749);
nor U933 (N_933,N_649,N_792);
and U934 (N_934,N_674,N_767);
and U935 (N_935,N_718,N_739);
and U936 (N_936,N_726,N_759);
and U937 (N_937,N_696,N_722);
nand U938 (N_938,N_751,N_752);
nor U939 (N_939,N_652,N_679);
nor U940 (N_940,N_760,N_718);
and U941 (N_941,N_617,N_789);
nand U942 (N_942,N_770,N_781);
nor U943 (N_943,N_616,N_794);
nor U944 (N_944,N_724,N_746);
xor U945 (N_945,N_609,N_743);
nand U946 (N_946,N_762,N_780);
nand U947 (N_947,N_612,N_676);
or U948 (N_948,N_731,N_663);
nor U949 (N_949,N_783,N_717);
nand U950 (N_950,N_663,N_676);
and U951 (N_951,N_790,N_673);
or U952 (N_952,N_717,N_702);
and U953 (N_953,N_758,N_716);
nor U954 (N_954,N_799,N_638);
nor U955 (N_955,N_706,N_655);
nand U956 (N_956,N_661,N_679);
or U957 (N_957,N_765,N_603);
and U958 (N_958,N_754,N_798);
and U959 (N_959,N_768,N_789);
xnor U960 (N_960,N_608,N_609);
or U961 (N_961,N_739,N_723);
nor U962 (N_962,N_764,N_733);
and U963 (N_963,N_732,N_607);
nor U964 (N_964,N_736,N_784);
nor U965 (N_965,N_738,N_788);
nand U966 (N_966,N_710,N_677);
or U967 (N_967,N_672,N_719);
nand U968 (N_968,N_718,N_626);
or U969 (N_969,N_607,N_637);
and U970 (N_970,N_775,N_774);
and U971 (N_971,N_741,N_637);
nor U972 (N_972,N_754,N_739);
or U973 (N_973,N_657,N_665);
and U974 (N_974,N_628,N_744);
nor U975 (N_975,N_667,N_605);
nand U976 (N_976,N_699,N_797);
and U977 (N_977,N_781,N_707);
nor U978 (N_978,N_701,N_794);
and U979 (N_979,N_779,N_625);
and U980 (N_980,N_620,N_686);
nor U981 (N_981,N_628,N_787);
nor U982 (N_982,N_751,N_691);
and U983 (N_983,N_617,N_677);
and U984 (N_984,N_769,N_788);
or U985 (N_985,N_769,N_778);
nand U986 (N_986,N_779,N_739);
or U987 (N_987,N_775,N_614);
nand U988 (N_988,N_721,N_613);
nor U989 (N_989,N_755,N_655);
nand U990 (N_990,N_725,N_671);
nand U991 (N_991,N_629,N_794);
and U992 (N_992,N_646,N_745);
or U993 (N_993,N_611,N_640);
nor U994 (N_994,N_685,N_757);
and U995 (N_995,N_661,N_672);
or U996 (N_996,N_748,N_666);
and U997 (N_997,N_726,N_762);
nand U998 (N_998,N_706,N_626);
nand U999 (N_999,N_689,N_640);
and U1000 (N_1000,N_855,N_945);
nand U1001 (N_1001,N_981,N_983);
nand U1002 (N_1002,N_825,N_996);
nand U1003 (N_1003,N_958,N_940);
nand U1004 (N_1004,N_821,N_876);
nor U1005 (N_1005,N_897,N_913);
and U1006 (N_1006,N_954,N_872);
or U1007 (N_1007,N_870,N_874);
and U1008 (N_1008,N_888,N_801);
or U1009 (N_1009,N_829,N_950);
nand U1010 (N_1010,N_863,N_849);
and U1011 (N_1011,N_815,N_808);
nor U1012 (N_1012,N_916,N_973);
or U1013 (N_1013,N_967,N_809);
or U1014 (N_1014,N_988,N_959);
nand U1015 (N_1015,N_850,N_978);
or U1016 (N_1016,N_957,N_938);
or U1017 (N_1017,N_997,N_928);
or U1018 (N_1018,N_917,N_846);
xnor U1019 (N_1019,N_856,N_949);
nor U1020 (N_1020,N_841,N_814);
or U1021 (N_1021,N_898,N_867);
or U1022 (N_1022,N_971,N_823);
nor U1023 (N_1023,N_925,N_882);
or U1024 (N_1024,N_820,N_879);
nor U1025 (N_1025,N_826,N_941);
or U1026 (N_1026,N_896,N_862);
or U1027 (N_1027,N_933,N_901);
or U1028 (N_1028,N_805,N_861);
or U1029 (N_1029,N_935,N_868);
nand U1030 (N_1030,N_934,N_974);
xor U1031 (N_1031,N_847,N_830);
and U1032 (N_1032,N_889,N_946);
nand U1033 (N_1033,N_903,N_900);
or U1034 (N_1034,N_836,N_985);
and U1035 (N_1035,N_979,N_892);
nand U1036 (N_1036,N_811,N_812);
nand U1037 (N_1037,N_911,N_895);
or U1038 (N_1038,N_852,N_869);
nor U1039 (N_1039,N_839,N_998);
or U1040 (N_1040,N_926,N_924);
nor U1041 (N_1041,N_822,N_920);
nand U1042 (N_1042,N_956,N_833);
or U1043 (N_1043,N_854,N_838);
nor U1044 (N_1044,N_929,N_878);
nand U1045 (N_1045,N_851,N_877);
nor U1046 (N_1046,N_976,N_918);
and U1047 (N_1047,N_904,N_943);
nand U1048 (N_1048,N_845,N_964);
and U1049 (N_1049,N_902,N_816);
and U1050 (N_1050,N_914,N_884);
nand U1051 (N_1051,N_939,N_802);
nor U1052 (N_1052,N_969,N_894);
nor U1053 (N_1053,N_936,N_932);
and U1054 (N_1054,N_963,N_899);
nand U1055 (N_1055,N_887,N_990);
nand U1056 (N_1056,N_953,N_960);
and U1057 (N_1057,N_944,N_858);
or U1058 (N_1058,N_986,N_875);
nand U1059 (N_1059,N_927,N_968);
nor U1060 (N_1060,N_912,N_893);
nor U1061 (N_1061,N_961,N_952);
nor U1062 (N_1062,N_885,N_837);
or U1063 (N_1063,N_871,N_819);
xor U1064 (N_1064,N_804,N_915);
or U1065 (N_1065,N_857,N_947);
nor U1066 (N_1066,N_866,N_970);
nand U1067 (N_1067,N_864,N_860);
or U1068 (N_1068,N_853,N_818);
nand U1069 (N_1069,N_827,N_831);
and U1070 (N_1070,N_890,N_992);
nand U1071 (N_1071,N_919,N_994);
and U1072 (N_1072,N_859,N_806);
and U1073 (N_1073,N_828,N_930);
and U1074 (N_1074,N_993,N_977);
or U1075 (N_1075,N_907,N_922);
nand U1076 (N_1076,N_965,N_848);
nor U1077 (N_1077,N_999,N_800);
and U1078 (N_1078,N_835,N_931);
xnor U1079 (N_1079,N_937,N_865);
xor U1080 (N_1080,N_921,N_982);
xnor U1081 (N_1081,N_807,N_813);
nand U1082 (N_1082,N_980,N_906);
or U1083 (N_1083,N_995,N_817);
nor U1084 (N_1084,N_975,N_908);
nand U1085 (N_1085,N_923,N_984);
nand U1086 (N_1086,N_803,N_972);
and U1087 (N_1087,N_948,N_810);
or U1088 (N_1088,N_873,N_962);
nor U1089 (N_1089,N_886,N_942);
nand U1090 (N_1090,N_840,N_834);
nand U1091 (N_1091,N_843,N_832);
and U1092 (N_1092,N_891,N_881);
or U1093 (N_1093,N_989,N_824);
nand U1094 (N_1094,N_987,N_951);
or U1095 (N_1095,N_883,N_844);
or U1096 (N_1096,N_905,N_880);
nor U1097 (N_1097,N_842,N_955);
nand U1098 (N_1098,N_910,N_909);
nor U1099 (N_1099,N_966,N_991);
and U1100 (N_1100,N_841,N_971);
nand U1101 (N_1101,N_880,N_813);
or U1102 (N_1102,N_957,N_992);
and U1103 (N_1103,N_954,N_992);
or U1104 (N_1104,N_886,N_828);
nand U1105 (N_1105,N_961,N_836);
or U1106 (N_1106,N_885,N_859);
or U1107 (N_1107,N_901,N_802);
and U1108 (N_1108,N_802,N_985);
or U1109 (N_1109,N_943,N_978);
nor U1110 (N_1110,N_839,N_853);
nor U1111 (N_1111,N_890,N_891);
nor U1112 (N_1112,N_922,N_959);
and U1113 (N_1113,N_905,N_803);
nand U1114 (N_1114,N_844,N_878);
or U1115 (N_1115,N_967,N_995);
nor U1116 (N_1116,N_889,N_837);
and U1117 (N_1117,N_866,N_902);
and U1118 (N_1118,N_937,N_809);
nor U1119 (N_1119,N_990,N_867);
and U1120 (N_1120,N_818,N_913);
or U1121 (N_1121,N_984,N_935);
or U1122 (N_1122,N_812,N_809);
nor U1123 (N_1123,N_819,N_844);
and U1124 (N_1124,N_915,N_983);
nand U1125 (N_1125,N_973,N_809);
nand U1126 (N_1126,N_981,N_807);
nand U1127 (N_1127,N_957,N_962);
nand U1128 (N_1128,N_858,N_852);
or U1129 (N_1129,N_834,N_915);
nand U1130 (N_1130,N_928,N_911);
and U1131 (N_1131,N_950,N_969);
or U1132 (N_1132,N_833,N_869);
and U1133 (N_1133,N_976,N_841);
and U1134 (N_1134,N_916,N_893);
or U1135 (N_1135,N_946,N_836);
or U1136 (N_1136,N_974,N_800);
and U1137 (N_1137,N_920,N_891);
and U1138 (N_1138,N_979,N_829);
or U1139 (N_1139,N_917,N_894);
and U1140 (N_1140,N_942,N_826);
and U1141 (N_1141,N_962,N_985);
or U1142 (N_1142,N_806,N_977);
or U1143 (N_1143,N_878,N_811);
nand U1144 (N_1144,N_974,N_984);
or U1145 (N_1145,N_963,N_812);
and U1146 (N_1146,N_858,N_969);
or U1147 (N_1147,N_858,N_836);
nand U1148 (N_1148,N_944,N_928);
nor U1149 (N_1149,N_940,N_819);
xnor U1150 (N_1150,N_821,N_819);
and U1151 (N_1151,N_829,N_910);
and U1152 (N_1152,N_983,N_841);
nand U1153 (N_1153,N_867,N_953);
or U1154 (N_1154,N_974,N_879);
or U1155 (N_1155,N_927,N_895);
and U1156 (N_1156,N_911,N_933);
or U1157 (N_1157,N_894,N_949);
nor U1158 (N_1158,N_838,N_967);
and U1159 (N_1159,N_899,N_983);
nor U1160 (N_1160,N_998,N_858);
and U1161 (N_1161,N_958,N_952);
or U1162 (N_1162,N_814,N_827);
nor U1163 (N_1163,N_954,N_922);
nand U1164 (N_1164,N_829,N_915);
or U1165 (N_1165,N_991,N_881);
nor U1166 (N_1166,N_921,N_875);
and U1167 (N_1167,N_822,N_881);
nor U1168 (N_1168,N_862,N_966);
and U1169 (N_1169,N_830,N_876);
nor U1170 (N_1170,N_896,N_837);
nor U1171 (N_1171,N_836,N_863);
or U1172 (N_1172,N_853,N_934);
nand U1173 (N_1173,N_931,N_864);
nor U1174 (N_1174,N_826,N_863);
nand U1175 (N_1175,N_959,N_984);
or U1176 (N_1176,N_872,N_814);
and U1177 (N_1177,N_862,N_804);
or U1178 (N_1178,N_966,N_893);
or U1179 (N_1179,N_871,N_836);
nor U1180 (N_1180,N_830,N_881);
nor U1181 (N_1181,N_976,N_962);
or U1182 (N_1182,N_914,N_957);
and U1183 (N_1183,N_885,N_831);
or U1184 (N_1184,N_935,N_954);
nor U1185 (N_1185,N_979,N_857);
or U1186 (N_1186,N_824,N_811);
and U1187 (N_1187,N_932,N_866);
or U1188 (N_1188,N_965,N_903);
or U1189 (N_1189,N_829,N_930);
nand U1190 (N_1190,N_805,N_851);
or U1191 (N_1191,N_811,N_865);
nor U1192 (N_1192,N_936,N_805);
and U1193 (N_1193,N_998,N_920);
or U1194 (N_1194,N_944,N_892);
nor U1195 (N_1195,N_952,N_862);
or U1196 (N_1196,N_954,N_911);
nor U1197 (N_1197,N_970,N_804);
and U1198 (N_1198,N_880,N_891);
and U1199 (N_1199,N_814,N_934);
or U1200 (N_1200,N_1099,N_1040);
or U1201 (N_1201,N_1146,N_1137);
and U1202 (N_1202,N_1078,N_1135);
nor U1203 (N_1203,N_1134,N_1126);
nand U1204 (N_1204,N_1162,N_1022);
and U1205 (N_1205,N_1064,N_1149);
nand U1206 (N_1206,N_1110,N_1142);
nand U1207 (N_1207,N_1106,N_1088);
nor U1208 (N_1208,N_1143,N_1176);
nor U1209 (N_1209,N_1029,N_1198);
nand U1210 (N_1210,N_1168,N_1023);
or U1211 (N_1211,N_1079,N_1053);
or U1212 (N_1212,N_1151,N_1034);
or U1213 (N_1213,N_1130,N_1039);
nor U1214 (N_1214,N_1189,N_1132);
nand U1215 (N_1215,N_1157,N_1036);
nor U1216 (N_1216,N_1046,N_1052);
nor U1217 (N_1217,N_1083,N_1159);
or U1218 (N_1218,N_1101,N_1073);
or U1219 (N_1219,N_1165,N_1153);
and U1220 (N_1220,N_1058,N_1115);
or U1221 (N_1221,N_1035,N_1103);
and U1222 (N_1222,N_1090,N_1139);
nor U1223 (N_1223,N_1048,N_1019);
and U1224 (N_1224,N_1155,N_1171);
or U1225 (N_1225,N_1102,N_1014);
or U1226 (N_1226,N_1147,N_1108);
nand U1227 (N_1227,N_1123,N_1156);
or U1228 (N_1228,N_1131,N_1133);
nand U1229 (N_1229,N_1150,N_1051);
or U1230 (N_1230,N_1028,N_1017);
nor U1231 (N_1231,N_1075,N_1077);
or U1232 (N_1232,N_1169,N_1182);
nor U1233 (N_1233,N_1027,N_1031);
nand U1234 (N_1234,N_1175,N_1122);
or U1235 (N_1235,N_1093,N_1127);
or U1236 (N_1236,N_1091,N_1063);
nor U1237 (N_1237,N_1117,N_1094);
and U1238 (N_1238,N_1125,N_1013);
nand U1239 (N_1239,N_1170,N_1164);
nor U1240 (N_1240,N_1066,N_1100);
and U1241 (N_1241,N_1119,N_1181);
or U1242 (N_1242,N_1057,N_1059);
or U1243 (N_1243,N_1166,N_1005);
and U1244 (N_1244,N_1192,N_1196);
or U1245 (N_1245,N_1054,N_1113);
or U1246 (N_1246,N_1007,N_1067);
nor U1247 (N_1247,N_1177,N_1163);
nand U1248 (N_1248,N_1193,N_1081);
nand U1249 (N_1249,N_1140,N_1138);
and U1250 (N_1250,N_1178,N_1076);
or U1251 (N_1251,N_1037,N_1174);
nand U1252 (N_1252,N_1030,N_1118);
xor U1253 (N_1253,N_1085,N_1105);
nand U1254 (N_1254,N_1097,N_1129);
or U1255 (N_1255,N_1050,N_1070);
and U1256 (N_1256,N_1011,N_1199);
and U1257 (N_1257,N_1111,N_1179);
or U1258 (N_1258,N_1009,N_1089);
nand U1259 (N_1259,N_1056,N_1041);
nor U1260 (N_1260,N_1161,N_1074);
nor U1261 (N_1261,N_1060,N_1069);
nor U1262 (N_1262,N_1012,N_1187);
and U1263 (N_1263,N_1032,N_1044);
nor U1264 (N_1264,N_1104,N_1158);
and U1265 (N_1265,N_1194,N_1062);
nand U1266 (N_1266,N_1114,N_1141);
nor U1267 (N_1267,N_1121,N_1095);
and U1268 (N_1268,N_1092,N_1107);
or U1269 (N_1269,N_1003,N_1082);
nor U1270 (N_1270,N_1144,N_1043);
or U1271 (N_1271,N_1098,N_1109);
nor U1272 (N_1272,N_1190,N_1049);
and U1273 (N_1273,N_1152,N_1055);
nor U1274 (N_1274,N_1038,N_1096);
nand U1275 (N_1275,N_1180,N_1148);
and U1276 (N_1276,N_1015,N_1124);
xnor U1277 (N_1277,N_1010,N_1002);
or U1278 (N_1278,N_1128,N_1160);
or U1279 (N_1279,N_1016,N_1086);
and U1280 (N_1280,N_1000,N_1065);
nand U1281 (N_1281,N_1008,N_1068);
or U1282 (N_1282,N_1195,N_1001);
and U1283 (N_1283,N_1145,N_1025);
nand U1284 (N_1284,N_1047,N_1197);
nor U1285 (N_1285,N_1184,N_1167);
nand U1286 (N_1286,N_1188,N_1042);
or U1287 (N_1287,N_1112,N_1072);
nand U1288 (N_1288,N_1173,N_1120);
nand U1289 (N_1289,N_1006,N_1191);
xor U1290 (N_1290,N_1026,N_1018);
nor U1291 (N_1291,N_1020,N_1080);
or U1292 (N_1292,N_1136,N_1045);
nor U1293 (N_1293,N_1084,N_1186);
nand U1294 (N_1294,N_1024,N_1087);
and U1295 (N_1295,N_1116,N_1071);
nand U1296 (N_1296,N_1033,N_1154);
or U1297 (N_1297,N_1185,N_1183);
and U1298 (N_1298,N_1172,N_1004);
and U1299 (N_1299,N_1021,N_1061);
and U1300 (N_1300,N_1050,N_1019);
and U1301 (N_1301,N_1149,N_1142);
nand U1302 (N_1302,N_1036,N_1196);
xor U1303 (N_1303,N_1015,N_1076);
or U1304 (N_1304,N_1156,N_1032);
nand U1305 (N_1305,N_1156,N_1096);
or U1306 (N_1306,N_1180,N_1119);
nor U1307 (N_1307,N_1190,N_1175);
nor U1308 (N_1308,N_1121,N_1192);
or U1309 (N_1309,N_1163,N_1140);
or U1310 (N_1310,N_1142,N_1141);
nand U1311 (N_1311,N_1079,N_1061);
xnor U1312 (N_1312,N_1193,N_1143);
or U1313 (N_1313,N_1094,N_1024);
or U1314 (N_1314,N_1164,N_1102);
or U1315 (N_1315,N_1069,N_1030);
nor U1316 (N_1316,N_1033,N_1172);
and U1317 (N_1317,N_1168,N_1107);
nor U1318 (N_1318,N_1117,N_1182);
and U1319 (N_1319,N_1144,N_1185);
nor U1320 (N_1320,N_1011,N_1157);
nand U1321 (N_1321,N_1001,N_1107);
nor U1322 (N_1322,N_1156,N_1113);
and U1323 (N_1323,N_1059,N_1120);
nand U1324 (N_1324,N_1078,N_1116);
nor U1325 (N_1325,N_1193,N_1053);
and U1326 (N_1326,N_1038,N_1050);
and U1327 (N_1327,N_1000,N_1091);
nand U1328 (N_1328,N_1198,N_1013);
nor U1329 (N_1329,N_1142,N_1036);
or U1330 (N_1330,N_1037,N_1118);
nor U1331 (N_1331,N_1144,N_1192);
and U1332 (N_1332,N_1180,N_1037);
and U1333 (N_1333,N_1180,N_1120);
nand U1334 (N_1334,N_1044,N_1163);
and U1335 (N_1335,N_1037,N_1108);
nor U1336 (N_1336,N_1157,N_1050);
or U1337 (N_1337,N_1035,N_1048);
or U1338 (N_1338,N_1069,N_1127);
and U1339 (N_1339,N_1084,N_1121);
and U1340 (N_1340,N_1088,N_1003);
nor U1341 (N_1341,N_1036,N_1171);
and U1342 (N_1342,N_1018,N_1029);
nand U1343 (N_1343,N_1023,N_1114);
nand U1344 (N_1344,N_1150,N_1037);
nand U1345 (N_1345,N_1100,N_1042);
or U1346 (N_1346,N_1197,N_1005);
and U1347 (N_1347,N_1004,N_1065);
or U1348 (N_1348,N_1055,N_1143);
or U1349 (N_1349,N_1113,N_1034);
or U1350 (N_1350,N_1167,N_1104);
or U1351 (N_1351,N_1054,N_1064);
xnor U1352 (N_1352,N_1054,N_1105);
or U1353 (N_1353,N_1015,N_1187);
xnor U1354 (N_1354,N_1035,N_1174);
or U1355 (N_1355,N_1182,N_1023);
and U1356 (N_1356,N_1098,N_1023);
and U1357 (N_1357,N_1067,N_1130);
and U1358 (N_1358,N_1110,N_1023);
and U1359 (N_1359,N_1064,N_1138);
nor U1360 (N_1360,N_1084,N_1172);
or U1361 (N_1361,N_1058,N_1126);
or U1362 (N_1362,N_1153,N_1189);
nor U1363 (N_1363,N_1029,N_1111);
nand U1364 (N_1364,N_1177,N_1113);
or U1365 (N_1365,N_1069,N_1174);
or U1366 (N_1366,N_1008,N_1054);
and U1367 (N_1367,N_1135,N_1015);
xnor U1368 (N_1368,N_1199,N_1114);
and U1369 (N_1369,N_1109,N_1087);
or U1370 (N_1370,N_1121,N_1103);
or U1371 (N_1371,N_1197,N_1038);
or U1372 (N_1372,N_1062,N_1179);
nand U1373 (N_1373,N_1081,N_1163);
or U1374 (N_1374,N_1179,N_1199);
nand U1375 (N_1375,N_1061,N_1163);
nand U1376 (N_1376,N_1085,N_1103);
nand U1377 (N_1377,N_1131,N_1011);
or U1378 (N_1378,N_1081,N_1022);
and U1379 (N_1379,N_1102,N_1179);
nand U1380 (N_1380,N_1086,N_1096);
nand U1381 (N_1381,N_1116,N_1127);
nor U1382 (N_1382,N_1163,N_1057);
xnor U1383 (N_1383,N_1153,N_1107);
nor U1384 (N_1384,N_1050,N_1009);
nand U1385 (N_1385,N_1105,N_1017);
and U1386 (N_1386,N_1148,N_1120);
nand U1387 (N_1387,N_1058,N_1196);
or U1388 (N_1388,N_1065,N_1003);
or U1389 (N_1389,N_1146,N_1174);
nor U1390 (N_1390,N_1088,N_1183);
and U1391 (N_1391,N_1194,N_1134);
nand U1392 (N_1392,N_1059,N_1101);
nand U1393 (N_1393,N_1172,N_1185);
and U1394 (N_1394,N_1131,N_1028);
xnor U1395 (N_1395,N_1155,N_1199);
nand U1396 (N_1396,N_1082,N_1173);
or U1397 (N_1397,N_1179,N_1121);
nand U1398 (N_1398,N_1065,N_1197);
nor U1399 (N_1399,N_1029,N_1017);
xnor U1400 (N_1400,N_1373,N_1359);
nor U1401 (N_1401,N_1376,N_1386);
nand U1402 (N_1402,N_1260,N_1274);
and U1403 (N_1403,N_1207,N_1202);
or U1404 (N_1404,N_1328,N_1203);
nand U1405 (N_1405,N_1278,N_1242);
or U1406 (N_1406,N_1313,N_1388);
and U1407 (N_1407,N_1234,N_1356);
nand U1408 (N_1408,N_1251,N_1349);
nand U1409 (N_1409,N_1364,N_1222);
nand U1410 (N_1410,N_1302,N_1389);
nand U1411 (N_1411,N_1390,N_1221);
and U1412 (N_1412,N_1214,N_1231);
nor U1413 (N_1413,N_1334,N_1295);
nand U1414 (N_1414,N_1200,N_1263);
or U1415 (N_1415,N_1246,N_1369);
nor U1416 (N_1416,N_1285,N_1336);
nor U1417 (N_1417,N_1235,N_1227);
or U1418 (N_1418,N_1385,N_1283);
nand U1419 (N_1419,N_1316,N_1252);
nor U1420 (N_1420,N_1280,N_1267);
nor U1421 (N_1421,N_1395,N_1332);
or U1422 (N_1422,N_1250,N_1318);
nor U1423 (N_1423,N_1317,N_1290);
and U1424 (N_1424,N_1394,N_1237);
nand U1425 (N_1425,N_1345,N_1309);
nand U1426 (N_1426,N_1387,N_1220);
and U1427 (N_1427,N_1211,N_1284);
nor U1428 (N_1428,N_1218,N_1230);
or U1429 (N_1429,N_1398,N_1350);
nand U1430 (N_1430,N_1253,N_1311);
or U1431 (N_1431,N_1338,N_1396);
nor U1432 (N_1432,N_1357,N_1206);
and U1433 (N_1433,N_1303,N_1301);
and U1434 (N_1434,N_1383,N_1341);
or U1435 (N_1435,N_1312,N_1233);
nor U1436 (N_1436,N_1346,N_1216);
nor U1437 (N_1437,N_1293,N_1205);
and U1438 (N_1438,N_1210,N_1380);
nand U1439 (N_1439,N_1339,N_1322);
and U1440 (N_1440,N_1340,N_1297);
nand U1441 (N_1441,N_1367,N_1370);
and U1442 (N_1442,N_1372,N_1358);
nand U1443 (N_1443,N_1254,N_1259);
xor U1444 (N_1444,N_1375,N_1308);
or U1445 (N_1445,N_1307,N_1265);
nand U1446 (N_1446,N_1391,N_1262);
nand U1447 (N_1447,N_1273,N_1219);
and U1448 (N_1448,N_1229,N_1298);
and U1449 (N_1449,N_1314,N_1279);
nand U1450 (N_1450,N_1392,N_1217);
and U1451 (N_1451,N_1296,N_1365);
nand U1452 (N_1452,N_1304,N_1384);
and U1453 (N_1453,N_1258,N_1324);
and U1454 (N_1454,N_1330,N_1323);
or U1455 (N_1455,N_1226,N_1368);
or U1456 (N_1456,N_1277,N_1294);
and U1457 (N_1457,N_1288,N_1257);
nor U1458 (N_1458,N_1393,N_1321);
nand U1459 (N_1459,N_1282,N_1249);
or U1460 (N_1460,N_1300,N_1382);
or U1461 (N_1461,N_1272,N_1377);
or U1462 (N_1462,N_1232,N_1271);
nand U1463 (N_1463,N_1256,N_1223);
or U1464 (N_1464,N_1244,N_1239);
and U1465 (N_1465,N_1363,N_1329);
nor U1466 (N_1466,N_1354,N_1289);
and U1467 (N_1467,N_1268,N_1224);
nand U1468 (N_1468,N_1204,N_1291);
nand U1469 (N_1469,N_1326,N_1360);
nor U1470 (N_1470,N_1299,N_1261);
and U1471 (N_1471,N_1243,N_1236);
and U1472 (N_1472,N_1361,N_1335);
and U1473 (N_1473,N_1347,N_1362);
nand U1474 (N_1474,N_1238,N_1270);
and U1475 (N_1475,N_1247,N_1348);
nor U1476 (N_1476,N_1325,N_1351);
nand U1477 (N_1477,N_1381,N_1213);
and U1478 (N_1478,N_1266,N_1344);
nand U1479 (N_1479,N_1276,N_1371);
or U1480 (N_1480,N_1355,N_1281);
nor U1481 (N_1481,N_1209,N_1212);
nor U1482 (N_1482,N_1315,N_1399);
nand U1483 (N_1483,N_1245,N_1269);
nand U1484 (N_1484,N_1333,N_1327);
nor U1485 (N_1485,N_1306,N_1374);
nor U1486 (N_1486,N_1319,N_1342);
and U1487 (N_1487,N_1264,N_1215);
nor U1488 (N_1488,N_1379,N_1397);
or U1489 (N_1489,N_1353,N_1310);
or U1490 (N_1490,N_1320,N_1331);
and U1491 (N_1491,N_1378,N_1366);
nor U1492 (N_1492,N_1352,N_1225);
or U1493 (N_1493,N_1337,N_1275);
and U1494 (N_1494,N_1343,N_1305);
and U1495 (N_1495,N_1292,N_1255);
or U1496 (N_1496,N_1241,N_1228);
and U1497 (N_1497,N_1208,N_1201);
nor U1498 (N_1498,N_1240,N_1286);
nand U1499 (N_1499,N_1248,N_1287);
and U1500 (N_1500,N_1310,N_1345);
or U1501 (N_1501,N_1237,N_1293);
or U1502 (N_1502,N_1290,N_1265);
nand U1503 (N_1503,N_1301,N_1227);
nand U1504 (N_1504,N_1372,N_1277);
and U1505 (N_1505,N_1317,N_1249);
and U1506 (N_1506,N_1239,N_1218);
or U1507 (N_1507,N_1318,N_1299);
or U1508 (N_1508,N_1396,N_1318);
nand U1509 (N_1509,N_1343,N_1321);
or U1510 (N_1510,N_1394,N_1331);
nand U1511 (N_1511,N_1230,N_1388);
nor U1512 (N_1512,N_1237,N_1225);
nand U1513 (N_1513,N_1376,N_1294);
nand U1514 (N_1514,N_1396,N_1229);
nor U1515 (N_1515,N_1313,N_1252);
nand U1516 (N_1516,N_1215,N_1270);
nand U1517 (N_1517,N_1342,N_1385);
nor U1518 (N_1518,N_1341,N_1331);
nor U1519 (N_1519,N_1364,N_1289);
and U1520 (N_1520,N_1304,N_1238);
nand U1521 (N_1521,N_1339,N_1385);
or U1522 (N_1522,N_1356,N_1278);
nor U1523 (N_1523,N_1230,N_1287);
xnor U1524 (N_1524,N_1251,N_1337);
or U1525 (N_1525,N_1318,N_1262);
nor U1526 (N_1526,N_1254,N_1264);
nand U1527 (N_1527,N_1334,N_1315);
and U1528 (N_1528,N_1314,N_1316);
xor U1529 (N_1529,N_1368,N_1328);
and U1530 (N_1530,N_1328,N_1319);
nor U1531 (N_1531,N_1302,N_1336);
nand U1532 (N_1532,N_1321,N_1269);
nand U1533 (N_1533,N_1351,N_1220);
nor U1534 (N_1534,N_1349,N_1317);
and U1535 (N_1535,N_1314,N_1237);
nor U1536 (N_1536,N_1320,N_1304);
nand U1537 (N_1537,N_1264,N_1312);
nor U1538 (N_1538,N_1297,N_1397);
nand U1539 (N_1539,N_1215,N_1250);
or U1540 (N_1540,N_1289,N_1285);
and U1541 (N_1541,N_1366,N_1344);
and U1542 (N_1542,N_1280,N_1273);
nor U1543 (N_1543,N_1305,N_1203);
nor U1544 (N_1544,N_1370,N_1289);
or U1545 (N_1545,N_1345,N_1370);
nand U1546 (N_1546,N_1358,N_1288);
and U1547 (N_1547,N_1367,N_1210);
nor U1548 (N_1548,N_1305,N_1239);
or U1549 (N_1549,N_1304,N_1211);
and U1550 (N_1550,N_1295,N_1218);
nor U1551 (N_1551,N_1383,N_1334);
nor U1552 (N_1552,N_1278,N_1340);
and U1553 (N_1553,N_1306,N_1202);
or U1554 (N_1554,N_1329,N_1341);
nor U1555 (N_1555,N_1256,N_1209);
nand U1556 (N_1556,N_1282,N_1311);
and U1557 (N_1557,N_1383,N_1387);
nand U1558 (N_1558,N_1323,N_1291);
and U1559 (N_1559,N_1249,N_1387);
and U1560 (N_1560,N_1291,N_1252);
nor U1561 (N_1561,N_1340,N_1389);
nor U1562 (N_1562,N_1355,N_1216);
xnor U1563 (N_1563,N_1357,N_1218);
nand U1564 (N_1564,N_1290,N_1232);
nor U1565 (N_1565,N_1373,N_1321);
or U1566 (N_1566,N_1365,N_1368);
and U1567 (N_1567,N_1227,N_1315);
xor U1568 (N_1568,N_1206,N_1399);
xnor U1569 (N_1569,N_1333,N_1297);
nand U1570 (N_1570,N_1285,N_1301);
or U1571 (N_1571,N_1249,N_1307);
and U1572 (N_1572,N_1269,N_1250);
nand U1573 (N_1573,N_1259,N_1358);
nor U1574 (N_1574,N_1290,N_1376);
nand U1575 (N_1575,N_1211,N_1255);
or U1576 (N_1576,N_1335,N_1294);
or U1577 (N_1577,N_1286,N_1386);
nor U1578 (N_1578,N_1307,N_1368);
nor U1579 (N_1579,N_1381,N_1374);
nand U1580 (N_1580,N_1381,N_1386);
nor U1581 (N_1581,N_1393,N_1283);
nor U1582 (N_1582,N_1329,N_1259);
xnor U1583 (N_1583,N_1292,N_1336);
and U1584 (N_1584,N_1216,N_1347);
nor U1585 (N_1585,N_1223,N_1341);
nor U1586 (N_1586,N_1388,N_1315);
nand U1587 (N_1587,N_1348,N_1347);
and U1588 (N_1588,N_1257,N_1208);
nand U1589 (N_1589,N_1256,N_1326);
nand U1590 (N_1590,N_1245,N_1293);
and U1591 (N_1591,N_1298,N_1293);
or U1592 (N_1592,N_1306,N_1365);
nand U1593 (N_1593,N_1379,N_1366);
nand U1594 (N_1594,N_1275,N_1298);
nor U1595 (N_1595,N_1238,N_1393);
and U1596 (N_1596,N_1300,N_1250);
xor U1597 (N_1597,N_1390,N_1392);
nand U1598 (N_1598,N_1236,N_1220);
or U1599 (N_1599,N_1399,N_1355);
xnor U1600 (N_1600,N_1467,N_1464);
or U1601 (N_1601,N_1454,N_1522);
and U1602 (N_1602,N_1421,N_1460);
nand U1603 (N_1603,N_1448,N_1491);
nor U1604 (N_1604,N_1543,N_1596);
xor U1605 (N_1605,N_1499,N_1412);
or U1606 (N_1606,N_1413,N_1564);
or U1607 (N_1607,N_1514,N_1580);
or U1608 (N_1608,N_1561,N_1417);
nor U1609 (N_1609,N_1461,N_1584);
nor U1610 (N_1610,N_1541,N_1453);
nand U1611 (N_1611,N_1443,N_1599);
nor U1612 (N_1612,N_1469,N_1503);
xnor U1613 (N_1613,N_1478,N_1505);
nor U1614 (N_1614,N_1536,N_1486);
and U1615 (N_1615,N_1513,N_1550);
or U1616 (N_1616,N_1459,N_1493);
and U1617 (N_1617,N_1515,N_1587);
nor U1618 (N_1618,N_1558,N_1476);
and U1619 (N_1619,N_1487,N_1583);
nand U1620 (N_1620,N_1456,N_1559);
nand U1621 (N_1621,N_1437,N_1405);
or U1622 (N_1622,N_1468,N_1555);
nor U1623 (N_1623,N_1579,N_1542);
and U1624 (N_1624,N_1425,N_1597);
nor U1625 (N_1625,N_1576,N_1511);
or U1626 (N_1626,N_1444,N_1409);
and U1627 (N_1627,N_1483,N_1552);
and U1628 (N_1628,N_1560,N_1427);
and U1629 (N_1629,N_1482,N_1481);
nor U1630 (N_1630,N_1535,N_1598);
and U1631 (N_1631,N_1532,N_1423);
nand U1632 (N_1632,N_1498,N_1573);
xor U1633 (N_1633,N_1537,N_1553);
xor U1634 (N_1634,N_1591,N_1508);
and U1635 (N_1635,N_1529,N_1449);
nand U1636 (N_1636,N_1512,N_1489);
nor U1637 (N_1637,N_1402,N_1502);
nor U1638 (N_1638,N_1458,N_1588);
and U1639 (N_1639,N_1432,N_1490);
xor U1640 (N_1640,N_1465,N_1420);
or U1641 (N_1641,N_1477,N_1582);
or U1642 (N_1642,N_1457,N_1414);
nor U1643 (N_1643,N_1434,N_1504);
nor U1644 (N_1644,N_1523,N_1403);
and U1645 (N_1645,N_1571,N_1439);
nand U1646 (N_1646,N_1452,N_1494);
nor U1647 (N_1647,N_1418,N_1521);
nor U1648 (N_1648,N_1581,N_1518);
xor U1649 (N_1649,N_1530,N_1475);
nor U1650 (N_1650,N_1426,N_1435);
and U1651 (N_1651,N_1431,N_1416);
or U1652 (N_1652,N_1455,N_1497);
and U1653 (N_1653,N_1479,N_1411);
nor U1654 (N_1654,N_1472,N_1544);
and U1655 (N_1655,N_1540,N_1506);
and U1656 (N_1656,N_1492,N_1520);
nand U1657 (N_1657,N_1546,N_1401);
nand U1658 (N_1658,N_1562,N_1575);
nor U1659 (N_1659,N_1501,N_1570);
and U1660 (N_1660,N_1462,N_1507);
or U1661 (N_1661,N_1488,N_1586);
and U1662 (N_1662,N_1408,N_1572);
nand U1663 (N_1663,N_1567,N_1473);
nor U1664 (N_1664,N_1406,N_1525);
and U1665 (N_1665,N_1419,N_1450);
nand U1666 (N_1666,N_1484,N_1415);
nand U1667 (N_1667,N_1436,N_1451);
nand U1668 (N_1668,N_1429,N_1474);
nor U1669 (N_1669,N_1595,N_1430);
nand U1670 (N_1670,N_1500,N_1404);
or U1671 (N_1671,N_1446,N_1480);
or U1672 (N_1672,N_1549,N_1539);
nand U1673 (N_1673,N_1438,N_1548);
and U1674 (N_1674,N_1566,N_1551);
nand U1675 (N_1675,N_1422,N_1594);
or U1676 (N_1676,N_1574,N_1533);
and U1677 (N_1677,N_1568,N_1545);
or U1678 (N_1678,N_1441,N_1485);
or U1679 (N_1679,N_1578,N_1440);
and U1680 (N_1680,N_1424,N_1516);
nand U1681 (N_1681,N_1534,N_1554);
xnor U1682 (N_1682,N_1442,N_1428);
xnor U1683 (N_1683,N_1557,N_1531);
and U1684 (N_1684,N_1556,N_1593);
and U1685 (N_1685,N_1517,N_1495);
nor U1686 (N_1686,N_1519,N_1527);
nor U1687 (N_1687,N_1592,N_1445);
or U1688 (N_1688,N_1410,N_1528);
and U1689 (N_1689,N_1590,N_1433);
and U1690 (N_1690,N_1538,N_1471);
or U1691 (N_1691,N_1470,N_1589);
and U1692 (N_1692,N_1463,N_1524);
nand U1693 (N_1693,N_1509,N_1569);
or U1694 (N_1694,N_1547,N_1407);
nor U1695 (N_1695,N_1510,N_1447);
and U1696 (N_1696,N_1585,N_1496);
and U1697 (N_1697,N_1563,N_1400);
and U1698 (N_1698,N_1577,N_1526);
or U1699 (N_1699,N_1565,N_1466);
and U1700 (N_1700,N_1485,N_1476);
nor U1701 (N_1701,N_1527,N_1475);
nand U1702 (N_1702,N_1422,N_1465);
nand U1703 (N_1703,N_1449,N_1455);
xnor U1704 (N_1704,N_1532,N_1442);
nand U1705 (N_1705,N_1579,N_1535);
and U1706 (N_1706,N_1422,N_1463);
nor U1707 (N_1707,N_1513,N_1449);
and U1708 (N_1708,N_1477,N_1560);
nand U1709 (N_1709,N_1503,N_1477);
nand U1710 (N_1710,N_1440,N_1453);
or U1711 (N_1711,N_1412,N_1526);
nor U1712 (N_1712,N_1452,N_1473);
and U1713 (N_1713,N_1448,N_1579);
nor U1714 (N_1714,N_1536,N_1471);
xor U1715 (N_1715,N_1590,N_1456);
or U1716 (N_1716,N_1460,N_1564);
or U1717 (N_1717,N_1470,N_1527);
nand U1718 (N_1718,N_1557,N_1516);
or U1719 (N_1719,N_1412,N_1548);
nand U1720 (N_1720,N_1450,N_1432);
nand U1721 (N_1721,N_1503,N_1493);
nand U1722 (N_1722,N_1529,N_1557);
nor U1723 (N_1723,N_1505,N_1587);
nand U1724 (N_1724,N_1585,N_1587);
nor U1725 (N_1725,N_1589,N_1525);
nor U1726 (N_1726,N_1421,N_1528);
or U1727 (N_1727,N_1517,N_1537);
nand U1728 (N_1728,N_1497,N_1525);
xnor U1729 (N_1729,N_1559,N_1547);
nor U1730 (N_1730,N_1424,N_1453);
xnor U1731 (N_1731,N_1476,N_1436);
nor U1732 (N_1732,N_1410,N_1554);
nand U1733 (N_1733,N_1544,N_1594);
nor U1734 (N_1734,N_1461,N_1407);
nand U1735 (N_1735,N_1434,N_1598);
nand U1736 (N_1736,N_1486,N_1573);
or U1737 (N_1737,N_1414,N_1446);
or U1738 (N_1738,N_1572,N_1465);
or U1739 (N_1739,N_1548,N_1531);
or U1740 (N_1740,N_1476,N_1517);
or U1741 (N_1741,N_1543,N_1582);
nor U1742 (N_1742,N_1540,N_1406);
and U1743 (N_1743,N_1437,N_1596);
nor U1744 (N_1744,N_1569,N_1431);
nand U1745 (N_1745,N_1401,N_1562);
nor U1746 (N_1746,N_1461,N_1495);
nand U1747 (N_1747,N_1465,N_1599);
and U1748 (N_1748,N_1480,N_1598);
or U1749 (N_1749,N_1423,N_1560);
or U1750 (N_1750,N_1589,N_1410);
and U1751 (N_1751,N_1455,N_1575);
xor U1752 (N_1752,N_1472,N_1416);
nand U1753 (N_1753,N_1504,N_1409);
or U1754 (N_1754,N_1417,N_1487);
and U1755 (N_1755,N_1499,N_1423);
and U1756 (N_1756,N_1578,N_1402);
nand U1757 (N_1757,N_1527,N_1431);
nor U1758 (N_1758,N_1460,N_1429);
xnor U1759 (N_1759,N_1431,N_1451);
and U1760 (N_1760,N_1548,N_1592);
nor U1761 (N_1761,N_1525,N_1483);
or U1762 (N_1762,N_1443,N_1531);
or U1763 (N_1763,N_1404,N_1522);
and U1764 (N_1764,N_1496,N_1409);
and U1765 (N_1765,N_1489,N_1485);
or U1766 (N_1766,N_1568,N_1417);
and U1767 (N_1767,N_1508,N_1460);
nand U1768 (N_1768,N_1535,N_1403);
nand U1769 (N_1769,N_1532,N_1485);
or U1770 (N_1770,N_1410,N_1467);
or U1771 (N_1771,N_1407,N_1433);
nand U1772 (N_1772,N_1464,N_1469);
nand U1773 (N_1773,N_1587,N_1565);
nor U1774 (N_1774,N_1454,N_1573);
or U1775 (N_1775,N_1513,N_1469);
nand U1776 (N_1776,N_1435,N_1552);
nand U1777 (N_1777,N_1469,N_1555);
and U1778 (N_1778,N_1494,N_1499);
or U1779 (N_1779,N_1402,N_1425);
nand U1780 (N_1780,N_1537,N_1454);
nand U1781 (N_1781,N_1559,N_1458);
nand U1782 (N_1782,N_1431,N_1504);
and U1783 (N_1783,N_1414,N_1507);
nor U1784 (N_1784,N_1404,N_1529);
and U1785 (N_1785,N_1535,N_1522);
and U1786 (N_1786,N_1575,N_1472);
or U1787 (N_1787,N_1585,N_1423);
and U1788 (N_1788,N_1451,N_1506);
nand U1789 (N_1789,N_1434,N_1454);
nor U1790 (N_1790,N_1592,N_1573);
or U1791 (N_1791,N_1547,N_1539);
and U1792 (N_1792,N_1446,N_1474);
nand U1793 (N_1793,N_1532,N_1502);
nand U1794 (N_1794,N_1591,N_1489);
nand U1795 (N_1795,N_1403,N_1470);
nand U1796 (N_1796,N_1573,N_1414);
nand U1797 (N_1797,N_1453,N_1400);
and U1798 (N_1798,N_1484,N_1416);
or U1799 (N_1799,N_1558,N_1553);
and U1800 (N_1800,N_1667,N_1710);
or U1801 (N_1801,N_1654,N_1784);
nand U1802 (N_1802,N_1697,N_1670);
and U1803 (N_1803,N_1721,N_1712);
and U1804 (N_1804,N_1612,N_1780);
nor U1805 (N_1805,N_1762,N_1658);
nor U1806 (N_1806,N_1602,N_1788);
nand U1807 (N_1807,N_1662,N_1791);
or U1808 (N_1808,N_1778,N_1707);
and U1809 (N_1809,N_1643,N_1649);
nand U1810 (N_1810,N_1717,N_1674);
and U1811 (N_1811,N_1629,N_1641);
and U1812 (N_1812,N_1793,N_1601);
or U1813 (N_1813,N_1769,N_1720);
or U1814 (N_1814,N_1698,N_1764);
or U1815 (N_1815,N_1648,N_1668);
and U1816 (N_1816,N_1747,N_1759);
or U1817 (N_1817,N_1690,N_1789);
nand U1818 (N_1818,N_1651,N_1770);
and U1819 (N_1819,N_1718,N_1619);
xor U1820 (N_1820,N_1645,N_1708);
and U1821 (N_1821,N_1683,N_1615);
or U1822 (N_1822,N_1603,N_1610);
nor U1823 (N_1823,N_1618,N_1725);
and U1824 (N_1824,N_1751,N_1736);
nor U1825 (N_1825,N_1699,N_1761);
nand U1826 (N_1826,N_1626,N_1653);
or U1827 (N_1827,N_1608,N_1728);
or U1828 (N_1828,N_1605,N_1739);
and U1829 (N_1829,N_1774,N_1607);
nand U1830 (N_1830,N_1790,N_1692);
nand U1831 (N_1831,N_1659,N_1614);
and U1832 (N_1832,N_1628,N_1672);
or U1833 (N_1833,N_1685,N_1777);
nand U1834 (N_1834,N_1729,N_1743);
nor U1835 (N_1835,N_1624,N_1765);
nor U1836 (N_1836,N_1679,N_1611);
or U1837 (N_1837,N_1663,N_1622);
or U1838 (N_1838,N_1640,N_1745);
or U1839 (N_1839,N_1660,N_1688);
nor U1840 (N_1840,N_1782,N_1700);
and U1841 (N_1841,N_1726,N_1750);
or U1842 (N_1842,N_1706,N_1763);
and U1843 (N_1843,N_1732,N_1642);
nor U1844 (N_1844,N_1766,N_1703);
or U1845 (N_1845,N_1773,N_1673);
nand U1846 (N_1846,N_1731,N_1755);
nor U1847 (N_1847,N_1664,N_1696);
or U1848 (N_1848,N_1600,N_1635);
or U1849 (N_1849,N_1606,N_1689);
nor U1850 (N_1850,N_1634,N_1768);
nor U1851 (N_1851,N_1631,N_1735);
nor U1852 (N_1852,N_1695,N_1677);
and U1853 (N_1853,N_1709,N_1678);
nand U1854 (N_1854,N_1734,N_1633);
and U1855 (N_1855,N_1644,N_1785);
and U1856 (N_1856,N_1727,N_1702);
and U1857 (N_1857,N_1752,N_1730);
nand U1858 (N_1858,N_1617,N_1616);
and U1859 (N_1859,N_1627,N_1711);
nand U1860 (N_1860,N_1680,N_1613);
nand U1861 (N_1861,N_1771,N_1630);
nor U1862 (N_1862,N_1681,N_1657);
nand U1863 (N_1863,N_1738,N_1676);
or U1864 (N_1864,N_1723,N_1772);
and U1865 (N_1865,N_1715,N_1691);
or U1866 (N_1866,N_1737,N_1748);
xor U1867 (N_1867,N_1671,N_1779);
and U1868 (N_1868,N_1713,N_1705);
nor U1869 (N_1869,N_1693,N_1655);
and U1870 (N_1870,N_1756,N_1656);
or U1871 (N_1871,N_1632,N_1798);
nand U1872 (N_1872,N_1647,N_1701);
or U1873 (N_1873,N_1636,N_1795);
and U1874 (N_1874,N_1650,N_1661);
or U1875 (N_1875,N_1687,N_1754);
nand U1876 (N_1876,N_1799,N_1669);
nand U1877 (N_1877,N_1719,N_1637);
nor U1878 (N_1878,N_1746,N_1665);
and U1879 (N_1879,N_1652,N_1675);
or U1880 (N_1880,N_1722,N_1792);
or U1881 (N_1881,N_1786,N_1794);
and U1882 (N_1882,N_1623,N_1744);
nor U1883 (N_1883,N_1716,N_1742);
nand U1884 (N_1884,N_1760,N_1775);
or U1885 (N_1885,N_1609,N_1682);
nand U1886 (N_1886,N_1757,N_1767);
nand U1887 (N_1887,N_1620,N_1781);
xor U1888 (N_1888,N_1740,N_1758);
or U1889 (N_1889,N_1638,N_1733);
nor U1890 (N_1890,N_1684,N_1796);
nand U1891 (N_1891,N_1686,N_1704);
and U1892 (N_1892,N_1753,N_1621);
and U1893 (N_1893,N_1714,N_1741);
nand U1894 (N_1894,N_1646,N_1639);
or U1895 (N_1895,N_1783,N_1694);
and U1896 (N_1896,N_1787,N_1749);
nor U1897 (N_1897,N_1724,N_1625);
nor U1898 (N_1898,N_1797,N_1604);
and U1899 (N_1899,N_1776,N_1666);
nand U1900 (N_1900,N_1675,N_1791);
and U1901 (N_1901,N_1765,N_1629);
nor U1902 (N_1902,N_1655,N_1640);
or U1903 (N_1903,N_1610,N_1762);
and U1904 (N_1904,N_1709,N_1775);
xor U1905 (N_1905,N_1737,N_1652);
and U1906 (N_1906,N_1654,N_1715);
nor U1907 (N_1907,N_1696,N_1734);
or U1908 (N_1908,N_1677,N_1682);
nand U1909 (N_1909,N_1689,N_1639);
xnor U1910 (N_1910,N_1610,N_1715);
nor U1911 (N_1911,N_1738,N_1761);
nand U1912 (N_1912,N_1707,N_1691);
or U1913 (N_1913,N_1752,N_1719);
nor U1914 (N_1914,N_1769,N_1749);
xor U1915 (N_1915,N_1696,N_1679);
nor U1916 (N_1916,N_1612,N_1671);
xnor U1917 (N_1917,N_1681,N_1610);
and U1918 (N_1918,N_1794,N_1651);
or U1919 (N_1919,N_1727,N_1729);
and U1920 (N_1920,N_1627,N_1742);
and U1921 (N_1921,N_1738,N_1693);
nand U1922 (N_1922,N_1625,N_1611);
or U1923 (N_1923,N_1609,N_1751);
and U1924 (N_1924,N_1645,N_1741);
nand U1925 (N_1925,N_1743,N_1715);
nor U1926 (N_1926,N_1651,N_1747);
nand U1927 (N_1927,N_1605,N_1619);
nor U1928 (N_1928,N_1650,N_1667);
and U1929 (N_1929,N_1789,N_1619);
nand U1930 (N_1930,N_1638,N_1750);
or U1931 (N_1931,N_1732,N_1758);
and U1932 (N_1932,N_1706,N_1657);
or U1933 (N_1933,N_1688,N_1609);
and U1934 (N_1934,N_1671,N_1638);
or U1935 (N_1935,N_1745,N_1635);
and U1936 (N_1936,N_1645,N_1632);
nor U1937 (N_1937,N_1669,N_1648);
nand U1938 (N_1938,N_1755,N_1671);
nor U1939 (N_1939,N_1666,N_1668);
xor U1940 (N_1940,N_1602,N_1620);
nor U1941 (N_1941,N_1625,N_1717);
nand U1942 (N_1942,N_1623,N_1755);
nand U1943 (N_1943,N_1650,N_1720);
nor U1944 (N_1944,N_1747,N_1790);
nor U1945 (N_1945,N_1765,N_1714);
nor U1946 (N_1946,N_1654,N_1783);
nand U1947 (N_1947,N_1625,N_1658);
nor U1948 (N_1948,N_1745,N_1732);
and U1949 (N_1949,N_1679,N_1782);
nand U1950 (N_1950,N_1769,N_1656);
or U1951 (N_1951,N_1756,N_1716);
nand U1952 (N_1952,N_1662,N_1671);
nand U1953 (N_1953,N_1686,N_1672);
and U1954 (N_1954,N_1661,N_1770);
or U1955 (N_1955,N_1772,N_1752);
and U1956 (N_1956,N_1798,N_1765);
nor U1957 (N_1957,N_1705,N_1768);
or U1958 (N_1958,N_1681,N_1671);
and U1959 (N_1959,N_1692,N_1792);
nor U1960 (N_1960,N_1657,N_1703);
nor U1961 (N_1961,N_1771,N_1681);
or U1962 (N_1962,N_1697,N_1620);
and U1963 (N_1963,N_1736,N_1606);
nand U1964 (N_1964,N_1786,N_1695);
nand U1965 (N_1965,N_1660,N_1609);
and U1966 (N_1966,N_1696,N_1627);
and U1967 (N_1967,N_1738,N_1627);
or U1968 (N_1968,N_1715,N_1612);
and U1969 (N_1969,N_1721,N_1781);
nand U1970 (N_1970,N_1601,N_1778);
nand U1971 (N_1971,N_1748,N_1617);
nor U1972 (N_1972,N_1793,N_1710);
nor U1973 (N_1973,N_1660,N_1639);
nor U1974 (N_1974,N_1788,N_1757);
or U1975 (N_1975,N_1756,N_1741);
nand U1976 (N_1976,N_1614,N_1745);
or U1977 (N_1977,N_1776,N_1726);
or U1978 (N_1978,N_1611,N_1727);
and U1979 (N_1979,N_1639,N_1713);
and U1980 (N_1980,N_1626,N_1793);
or U1981 (N_1981,N_1741,N_1787);
and U1982 (N_1982,N_1747,N_1734);
or U1983 (N_1983,N_1671,N_1655);
nor U1984 (N_1984,N_1775,N_1700);
nor U1985 (N_1985,N_1799,N_1756);
and U1986 (N_1986,N_1770,N_1712);
nor U1987 (N_1987,N_1615,N_1657);
xor U1988 (N_1988,N_1725,N_1600);
or U1989 (N_1989,N_1700,N_1776);
nor U1990 (N_1990,N_1654,N_1752);
and U1991 (N_1991,N_1666,N_1650);
nand U1992 (N_1992,N_1692,N_1748);
nor U1993 (N_1993,N_1739,N_1735);
or U1994 (N_1994,N_1606,N_1627);
nor U1995 (N_1995,N_1690,N_1791);
nor U1996 (N_1996,N_1679,N_1728);
nand U1997 (N_1997,N_1696,N_1689);
nand U1998 (N_1998,N_1620,N_1754);
and U1999 (N_1999,N_1751,N_1738);
nand U2000 (N_2000,N_1834,N_1811);
nand U2001 (N_2001,N_1994,N_1916);
and U2002 (N_2002,N_1991,N_1995);
nand U2003 (N_2003,N_1851,N_1883);
or U2004 (N_2004,N_1908,N_1902);
or U2005 (N_2005,N_1817,N_1868);
and U2006 (N_2006,N_1803,N_1903);
nor U2007 (N_2007,N_1836,N_1959);
or U2008 (N_2008,N_1873,N_1978);
or U2009 (N_2009,N_1806,N_1900);
and U2010 (N_2010,N_1905,N_1906);
xor U2011 (N_2011,N_1897,N_1996);
nor U2012 (N_2012,N_1824,N_1935);
and U2013 (N_2013,N_1950,N_1945);
and U2014 (N_2014,N_1878,N_1909);
nor U2015 (N_2015,N_1933,N_1997);
and U2016 (N_2016,N_1813,N_1939);
nand U2017 (N_2017,N_1907,N_1827);
and U2018 (N_2018,N_1964,N_1967);
nand U2019 (N_2019,N_1852,N_1960);
or U2020 (N_2020,N_1999,N_1802);
nand U2021 (N_2021,N_1826,N_1853);
and U2022 (N_2022,N_1890,N_1872);
or U2023 (N_2023,N_1987,N_1914);
and U2024 (N_2024,N_1957,N_1923);
nor U2025 (N_2025,N_1892,N_1835);
and U2026 (N_2026,N_1877,N_1989);
nor U2027 (N_2027,N_1814,N_1915);
nand U2028 (N_2028,N_1816,N_1972);
nand U2029 (N_2029,N_1937,N_1855);
or U2030 (N_2030,N_1910,N_1893);
and U2031 (N_2031,N_1986,N_1912);
or U2032 (N_2032,N_1979,N_1831);
nor U2033 (N_2033,N_1988,N_1849);
and U2034 (N_2034,N_1946,N_1885);
nor U2035 (N_2035,N_1875,N_1940);
and U2036 (N_2036,N_1918,N_1975);
and U2037 (N_2037,N_1830,N_1861);
or U2038 (N_2038,N_1854,N_1936);
nand U2039 (N_2039,N_1932,N_1841);
nor U2040 (N_2040,N_1938,N_1840);
and U2041 (N_2041,N_1808,N_1931);
nand U2042 (N_2042,N_1842,N_1815);
nor U2043 (N_2043,N_1825,N_1823);
nand U2044 (N_2044,N_1862,N_1800);
nor U2045 (N_2045,N_1822,N_1969);
and U2046 (N_2046,N_1970,N_1981);
nand U2047 (N_2047,N_1819,N_1904);
nor U2048 (N_2048,N_1886,N_1829);
or U2049 (N_2049,N_1930,N_1913);
or U2050 (N_2050,N_1866,N_1838);
nand U2051 (N_2051,N_1901,N_1867);
nor U2052 (N_2052,N_1884,N_1954);
nor U2053 (N_2053,N_1899,N_1948);
nor U2054 (N_2054,N_1856,N_1980);
xor U2055 (N_2055,N_1846,N_1833);
or U2056 (N_2056,N_1828,N_1805);
and U2057 (N_2057,N_1882,N_1898);
nand U2058 (N_2058,N_1949,N_1821);
nor U2059 (N_2059,N_1865,N_1993);
or U2060 (N_2060,N_1810,N_1863);
and U2061 (N_2061,N_1801,N_1911);
nor U2062 (N_2062,N_1844,N_1845);
and U2063 (N_2063,N_1998,N_1818);
and U2064 (N_2064,N_1807,N_1924);
nand U2065 (N_2065,N_1887,N_1976);
nand U2066 (N_2066,N_1990,N_1966);
and U2067 (N_2067,N_1858,N_1926);
and U2068 (N_2068,N_1889,N_1971);
or U2069 (N_2069,N_1895,N_1984);
nor U2070 (N_2070,N_1963,N_1860);
nand U2071 (N_2071,N_1874,N_1837);
or U2072 (N_2072,N_1942,N_1961);
or U2073 (N_2073,N_1974,N_1820);
nor U2074 (N_2074,N_1894,N_1944);
nor U2075 (N_2075,N_1843,N_1925);
nand U2076 (N_2076,N_1992,N_1982);
and U2077 (N_2077,N_1857,N_1919);
nor U2078 (N_2078,N_1956,N_1922);
nand U2079 (N_2079,N_1864,N_1934);
or U2080 (N_2080,N_1958,N_1896);
and U2081 (N_2081,N_1921,N_1876);
nand U2082 (N_2082,N_1983,N_1977);
or U2083 (N_2083,N_1869,N_1973);
or U2084 (N_2084,N_1952,N_1847);
nor U2085 (N_2085,N_1968,N_1985);
or U2086 (N_2086,N_1812,N_1870);
or U2087 (N_2087,N_1891,N_1871);
and U2088 (N_2088,N_1928,N_1809);
nor U2089 (N_2089,N_1832,N_1879);
or U2090 (N_2090,N_1917,N_1951);
nor U2091 (N_2091,N_1955,N_1839);
xnor U2092 (N_2092,N_1929,N_1943);
nand U2093 (N_2093,N_1947,N_1888);
nor U2094 (N_2094,N_1920,N_1965);
nand U2095 (N_2095,N_1848,N_1953);
and U2096 (N_2096,N_1927,N_1850);
or U2097 (N_2097,N_1962,N_1859);
and U2098 (N_2098,N_1804,N_1941);
or U2099 (N_2099,N_1880,N_1881);
and U2100 (N_2100,N_1880,N_1892);
nand U2101 (N_2101,N_1822,N_1925);
nand U2102 (N_2102,N_1856,N_1938);
and U2103 (N_2103,N_1855,N_1801);
and U2104 (N_2104,N_1893,N_1816);
and U2105 (N_2105,N_1971,N_1925);
nor U2106 (N_2106,N_1896,N_1964);
or U2107 (N_2107,N_1966,N_1921);
and U2108 (N_2108,N_1836,N_1832);
xnor U2109 (N_2109,N_1955,N_1987);
nand U2110 (N_2110,N_1934,N_1844);
nand U2111 (N_2111,N_1920,N_1940);
nor U2112 (N_2112,N_1997,N_1976);
nor U2113 (N_2113,N_1802,N_1918);
nor U2114 (N_2114,N_1884,N_1895);
and U2115 (N_2115,N_1967,N_1809);
nand U2116 (N_2116,N_1902,N_1897);
and U2117 (N_2117,N_1818,N_1978);
and U2118 (N_2118,N_1842,N_1831);
or U2119 (N_2119,N_1973,N_1925);
nand U2120 (N_2120,N_1880,N_1864);
nand U2121 (N_2121,N_1990,N_1832);
or U2122 (N_2122,N_1833,N_1903);
or U2123 (N_2123,N_1823,N_1919);
and U2124 (N_2124,N_1805,N_1873);
nor U2125 (N_2125,N_1899,N_1977);
nand U2126 (N_2126,N_1980,N_1832);
and U2127 (N_2127,N_1833,N_1969);
nor U2128 (N_2128,N_1920,N_1913);
nor U2129 (N_2129,N_1931,N_1978);
or U2130 (N_2130,N_1894,N_1873);
nand U2131 (N_2131,N_1806,N_1978);
nor U2132 (N_2132,N_1890,N_1969);
nand U2133 (N_2133,N_1855,N_1830);
or U2134 (N_2134,N_1855,N_1892);
nand U2135 (N_2135,N_1846,N_1839);
and U2136 (N_2136,N_1859,N_1806);
and U2137 (N_2137,N_1891,N_1937);
or U2138 (N_2138,N_1908,N_1812);
or U2139 (N_2139,N_1880,N_1915);
nand U2140 (N_2140,N_1951,N_1851);
nand U2141 (N_2141,N_1843,N_1836);
nand U2142 (N_2142,N_1818,N_1892);
or U2143 (N_2143,N_1989,N_1833);
nor U2144 (N_2144,N_1907,N_1920);
nor U2145 (N_2145,N_1936,N_1850);
nor U2146 (N_2146,N_1893,N_1885);
nor U2147 (N_2147,N_1973,N_1980);
nand U2148 (N_2148,N_1822,N_1873);
nor U2149 (N_2149,N_1813,N_1842);
nand U2150 (N_2150,N_1929,N_1863);
and U2151 (N_2151,N_1838,N_1834);
and U2152 (N_2152,N_1952,N_1831);
nor U2153 (N_2153,N_1992,N_1864);
or U2154 (N_2154,N_1932,N_1885);
or U2155 (N_2155,N_1831,N_1868);
nand U2156 (N_2156,N_1804,N_1958);
nand U2157 (N_2157,N_1993,N_1855);
and U2158 (N_2158,N_1968,N_1967);
nor U2159 (N_2159,N_1870,N_1810);
or U2160 (N_2160,N_1804,N_1864);
and U2161 (N_2161,N_1880,N_1971);
and U2162 (N_2162,N_1900,N_1926);
nand U2163 (N_2163,N_1965,N_1847);
nand U2164 (N_2164,N_1979,N_1845);
or U2165 (N_2165,N_1929,N_1978);
or U2166 (N_2166,N_1894,N_1869);
nand U2167 (N_2167,N_1807,N_1944);
nor U2168 (N_2168,N_1973,N_1883);
xor U2169 (N_2169,N_1993,N_1911);
and U2170 (N_2170,N_1862,N_1854);
nand U2171 (N_2171,N_1926,N_1945);
nor U2172 (N_2172,N_1844,N_1927);
or U2173 (N_2173,N_1925,N_1946);
nand U2174 (N_2174,N_1869,N_1949);
or U2175 (N_2175,N_1883,N_1979);
and U2176 (N_2176,N_1889,N_1873);
nand U2177 (N_2177,N_1931,N_1811);
nand U2178 (N_2178,N_1936,N_1947);
or U2179 (N_2179,N_1989,N_1856);
or U2180 (N_2180,N_1956,N_1930);
and U2181 (N_2181,N_1946,N_1911);
nor U2182 (N_2182,N_1884,N_1921);
nand U2183 (N_2183,N_1838,N_1844);
nor U2184 (N_2184,N_1949,N_1842);
or U2185 (N_2185,N_1951,N_1849);
or U2186 (N_2186,N_1904,N_1859);
and U2187 (N_2187,N_1856,N_1981);
or U2188 (N_2188,N_1867,N_1954);
nand U2189 (N_2189,N_1809,N_1851);
and U2190 (N_2190,N_1934,N_1909);
nand U2191 (N_2191,N_1957,N_1992);
or U2192 (N_2192,N_1959,N_1946);
nand U2193 (N_2193,N_1980,N_1981);
and U2194 (N_2194,N_1890,N_1964);
nand U2195 (N_2195,N_1810,N_1935);
and U2196 (N_2196,N_1958,N_1999);
nor U2197 (N_2197,N_1881,N_1889);
and U2198 (N_2198,N_1805,N_1880);
nor U2199 (N_2199,N_1881,N_1990);
nor U2200 (N_2200,N_2102,N_2142);
xor U2201 (N_2201,N_2103,N_2121);
and U2202 (N_2202,N_2174,N_2050);
or U2203 (N_2203,N_2030,N_2026);
nor U2204 (N_2204,N_2053,N_2078);
nor U2205 (N_2205,N_2006,N_2060);
and U2206 (N_2206,N_2119,N_2074);
and U2207 (N_2207,N_2129,N_2004);
or U2208 (N_2208,N_2034,N_2143);
or U2209 (N_2209,N_2140,N_2032);
nand U2210 (N_2210,N_2123,N_2017);
nor U2211 (N_2211,N_2197,N_2101);
nand U2212 (N_2212,N_2010,N_2173);
or U2213 (N_2213,N_2138,N_2095);
and U2214 (N_2214,N_2183,N_2021);
nor U2215 (N_2215,N_2008,N_2007);
nand U2216 (N_2216,N_2000,N_2109);
nor U2217 (N_2217,N_2136,N_2066);
and U2218 (N_2218,N_2011,N_2016);
and U2219 (N_2219,N_2199,N_2064);
nor U2220 (N_2220,N_2118,N_2194);
and U2221 (N_2221,N_2156,N_2077);
nand U2222 (N_2222,N_2153,N_2039);
and U2223 (N_2223,N_2012,N_2167);
nand U2224 (N_2224,N_2133,N_2029);
nand U2225 (N_2225,N_2106,N_2155);
nor U2226 (N_2226,N_2161,N_2009);
nor U2227 (N_2227,N_2058,N_2145);
and U2228 (N_2228,N_2131,N_2170);
nor U2229 (N_2229,N_2023,N_2180);
nand U2230 (N_2230,N_2185,N_2148);
or U2231 (N_2231,N_2091,N_2024);
nor U2232 (N_2232,N_2019,N_2038);
and U2233 (N_2233,N_2144,N_2195);
nor U2234 (N_2234,N_2176,N_2188);
or U2235 (N_2235,N_2114,N_2149);
nor U2236 (N_2236,N_2125,N_2020);
xnor U2237 (N_2237,N_2163,N_2001);
nand U2238 (N_2238,N_2189,N_2067);
and U2239 (N_2239,N_2152,N_2098);
or U2240 (N_2240,N_2087,N_2073);
nand U2241 (N_2241,N_2147,N_2100);
nor U2242 (N_2242,N_2093,N_2122);
and U2243 (N_2243,N_2169,N_2097);
nor U2244 (N_2244,N_2094,N_2028);
nor U2245 (N_2245,N_2191,N_2126);
nor U2246 (N_2246,N_2177,N_2134);
and U2247 (N_2247,N_2107,N_2061);
nor U2248 (N_2248,N_2088,N_2048);
nand U2249 (N_2249,N_2022,N_2049);
nand U2250 (N_2250,N_2083,N_2154);
and U2251 (N_2251,N_2042,N_2193);
or U2252 (N_2252,N_2003,N_2057);
nor U2253 (N_2253,N_2166,N_2070);
and U2254 (N_2254,N_2130,N_2165);
and U2255 (N_2255,N_2027,N_2045);
and U2256 (N_2256,N_2116,N_2041);
or U2257 (N_2257,N_2076,N_2099);
or U2258 (N_2258,N_2090,N_2184);
nor U2259 (N_2259,N_2059,N_2192);
and U2260 (N_2260,N_2096,N_2141);
and U2261 (N_2261,N_2002,N_2159);
nor U2262 (N_2262,N_2047,N_2105);
or U2263 (N_2263,N_2127,N_2187);
nor U2264 (N_2264,N_2110,N_2052);
nand U2265 (N_2265,N_2117,N_2068);
and U2266 (N_2266,N_2162,N_2113);
and U2267 (N_2267,N_2085,N_2115);
and U2268 (N_2268,N_2054,N_2135);
nand U2269 (N_2269,N_2111,N_2089);
nand U2270 (N_2270,N_2015,N_2037);
xor U2271 (N_2271,N_2072,N_2175);
or U2272 (N_2272,N_2104,N_2086);
and U2273 (N_2273,N_2080,N_2124);
nor U2274 (N_2274,N_2018,N_2084);
and U2275 (N_2275,N_2065,N_2160);
nor U2276 (N_2276,N_2182,N_2079);
nor U2277 (N_2277,N_2040,N_2137);
nor U2278 (N_2278,N_2196,N_2157);
nand U2279 (N_2279,N_2128,N_2146);
nor U2280 (N_2280,N_2112,N_2178);
nand U2281 (N_2281,N_2092,N_2013);
xor U2282 (N_2282,N_2139,N_2151);
or U2283 (N_2283,N_2190,N_2035);
nand U2284 (N_2284,N_2044,N_2164);
or U2285 (N_2285,N_2186,N_2063);
nand U2286 (N_2286,N_2056,N_2150);
or U2287 (N_2287,N_2031,N_2051);
nor U2288 (N_2288,N_2005,N_2082);
or U2289 (N_2289,N_2198,N_2171);
nand U2290 (N_2290,N_2055,N_2046);
nand U2291 (N_2291,N_2179,N_2071);
nor U2292 (N_2292,N_2033,N_2081);
nor U2293 (N_2293,N_2108,N_2025);
nand U2294 (N_2294,N_2075,N_2172);
or U2295 (N_2295,N_2181,N_2014);
nand U2296 (N_2296,N_2043,N_2036);
xnor U2297 (N_2297,N_2158,N_2132);
nor U2298 (N_2298,N_2062,N_2168);
or U2299 (N_2299,N_2069,N_2120);
or U2300 (N_2300,N_2166,N_2031);
and U2301 (N_2301,N_2157,N_2012);
and U2302 (N_2302,N_2171,N_2120);
and U2303 (N_2303,N_2016,N_2139);
nand U2304 (N_2304,N_2180,N_2108);
and U2305 (N_2305,N_2183,N_2128);
or U2306 (N_2306,N_2079,N_2086);
nand U2307 (N_2307,N_2162,N_2032);
or U2308 (N_2308,N_2133,N_2006);
and U2309 (N_2309,N_2024,N_2075);
nand U2310 (N_2310,N_2055,N_2095);
nor U2311 (N_2311,N_2062,N_2041);
and U2312 (N_2312,N_2097,N_2100);
nand U2313 (N_2313,N_2112,N_2030);
and U2314 (N_2314,N_2072,N_2199);
nor U2315 (N_2315,N_2084,N_2131);
nor U2316 (N_2316,N_2118,N_2052);
or U2317 (N_2317,N_2145,N_2057);
nand U2318 (N_2318,N_2157,N_2040);
nand U2319 (N_2319,N_2033,N_2049);
nand U2320 (N_2320,N_2048,N_2198);
and U2321 (N_2321,N_2065,N_2151);
nand U2322 (N_2322,N_2033,N_2158);
nor U2323 (N_2323,N_2172,N_2071);
xor U2324 (N_2324,N_2185,N_2056);
nor U2325 (N_2325,N_2121,N_2074);
and U2326 (N_2326,N_2173,N_2138);
xor U2327 (N_2327,N_2029,N_2069);
and U2328 (N_2328,N_2091,N_2084);
nand U2329 (N_2329,N_2128,N_2114);
nand U2330 (N_2330,N_2139,N_2193);
nor U2331 (N_2331,N_2123,N_2008);
nor U2332 (N_2332,N_2065,N_2087);
or U2333 (N_2333,N_2090,N_2061);
or U2334 (N_2334,N_2134,N_2046);
or U2335 (N_2335,N_2148,N_2143);
or U2336 (N_2336,N_2020,N_2071);
or U2337 (N_2337,N_2134,N_2097);
nor U2338 (N_2338,N_2154,N_2168);
xnor U2339 (N_2339,N_2183,N_2036);
nand U2340 (N_2340,N_2146,N_2096);
or U2341 (N_2341,N_2013,N_2054);
nor U2342 (N_2342,N_2100,N_2151);
nor U2343 (N_2343,N_2080,N_2101);
nand U2344 (N_2344,N_2100,N_2165);
nand U2345 (N_2345,N_2136,N_2040);
and U2346 (N_2346,N_2056,N_2126);
nand U2347 (N_2347,N_2192,N_2199);
and U2348 (N_2348,N_2005,N_2039);
nor U2349 (N_2349,N_2150,N_2098);
or U2350 (N_2350,N_2120,N_2002);
nor U2351 (N_2351,N_2141,N_2091);
or U2352 (N_2352,N_2174,N_2180);
nor U2353 (N_2353,N_2142,N_2010);
nand U2354 (N_2354,N_2098,N_2167);
and U2355 (N_2355,N_2151,N_2172);
nor U2356 (N_2356,N_2135,N_2074);
or U2357 (N_2357,N_2178,N_2135);
xor U2358 (N_2358,N_2046,N_2010);
and U2359 (N_2359,N_2047,N_2160);
or U2360 (N_2360,N_2105,N_2054);
and U2361 (N_2361,N_2050,N_2031);
and U2362 (N_2362,N_2002,N_2079);
nor U2363 (N_2363,N_2147,N_2099);
or U2364 (N_2364,N_2165,N_2117);
nor U2365 (N_2365,N_2161,N_2064);
or U2366 (N_2366,N_2168,N_2117);
nand U2367 (N_2367,N_2078,N_2103);
nor U2368 (N_2368,N_2106,N_2031);
and U2369 (N_2369,N_2104,N_2134);
nand U2370 (N_2370,N_2133,N_2110);
nor U2371 (N_2371,N_2027,N_2142);
and U2372 (N_2372,N_2114,N_2058);
and U2373 (N_2373,N_2065,N_2107);
nand U2374 (N_2374,N_2080,N_2045);
or U2375 (N_2375,N_2189,N_2018);
or U2376 (N_2376,N_2090,N_2079);
or U2377 (N_2377,N_2131,N_2028);
or U2378 (N_2378,N_2127,N_2045);
and U2379 (N_2379,N_2018,N_2179);
and U2380 (N_2380,N_2186,N_2065);
xor U2381 (N_2381,N_2057,N_2038);
and U2382 (N_2382,N_2177,N_2019);
nand U2383 (N_2383,N_2093,N_2074);
or U2384 (N_2384,N_2104,N_2179);
and U2385 (N_2385,N_2088,N_2117);
or U2386 (N_2386,N_2160,N_2033);
and U2387 (N_2387,N_2003,N_2190);
nand U2388 (N_2388,N_2131,N_2149);
and U2389 (N_2389,N_2125,N_2006);
nand U2390 (N_2390,N_2133,N_2094);
and U2391 (N_2391,N_2049,N_2199);
nand U2392 (N_2392,N_2117,N_2034);
nand U2393 (N_2393,N_2167,N_2064);
and U2394 (N_2394,N_2123,N_2146);
and U2395 (N_2395,N_2003,N_2068);
nor U2396 (N_2396,N_2009,N_2054);
nand U2397 (N_2397,N_2047,N_2024);
nand U2398 (N_2398,N_2190,N_2174);
nor U2399 (N_2399,N_2078,N_2130);
nand U2400 (N_2400,N_2313,N_2237);
and U2401 (N_2401,N_2362,N_2223);
or U2402 (N_2402,N_2325,N_2368);
or U2403 (N_2403,N_2384,N_2342);
and U2404 (N_2404,N_2281,N_2338);
and U2405 (N_2405,N_2245,N_2373);
and U2406 (N_2406,N_2304,N_2346);
nor U2407 (N_2407,N_2321,N_2328);
and U2408 (N_2408,N_2225,N_2207);
or U2409 (N_2409,N_2234,N_2331);
and U2410 (N_2410,N_2280,N_2246);
nand U2411 (N_2411,N_2303,N_2269);
xnor U2412 (N_2412,N_2290,N_2244);
nand U2413 (N_2413,N_2359,N_2263);
nor U2414 (N_2414,N_2205,N_2274);
and U2415 (N_2415,N_2228,N_2337);
xor U2416 (N_2416,N_2397,N_2387);
or U2417 (N_2417,N_2332,N_2267);
or U2418 (N_2418,N_2247,N_2270);
nand U2419 (N_2419,N_2309,N_2218);
nor U2420 (N_2420,N_2382,N_2227);
and U2421 (N_2421,N_2353,N_2305);
nor U2422 (N_2422,N_2302,N_2284);
nor U2423 (N_2423,N_2286,N_2312);
xnor U2424 (N_2424,N_2398,N_2258);
or U2425 (N_2425,N_2344,N_2236);
or U2426 (N_2426,N_2334,N_2272);
and U2427 (N_2427,N_2335,N_2255);
or U2428 (N_2428,N_2377,N_2220);
nor U2429 (N_2429,N_2354,N_2233);
and U2430 (N_2430,N_2385,N_2379);
or U2431 (N_2431,N_2327,N_2333);
nand U2432 (N_2432,N_2367,N_2355);
nor U2433 (N_2433,N_2288,N_2381);
and U2434 (N_2434,N_2378,N_2215);
or U2435 (N_2435,N_2252,N_2210);
and U2436 (N_2436,N_2349,N_2307);
or U2437 (N_2437,N_2243,N_2213);
nor U2438 (N_2438,N_2294,N_2260);
or U2439 (N_2439,N_2226,N_2316);
nor U2440 (N_2440,N_2285,N_2230);
and U2441 (N_2441,N_2395,N_2217);
and U2442 (N_2442,N_2300,N_2229);
nor U2443 (N_2443,N_2278,N_2311);
and U2444 (N_2444,N_2340,N_2358);
nor U2445 (N_2445,N_2256,N_2329);
or U2446 (N_2446,N_2265,N_2323);
and U2447 (N_2447,N_2277,N_2360);
nand U2448 (N_2448,N_2296,N_2389);
or U2449 (N_2449,N_2211,N_2356);
xor U2450 (N_2450,N_2299,N_2212);
nand U2451 (N_2451,N_2241,N_2364);
nor U2452 (N_2452,N_2259,N_2208);
or U2453 (N_2453,N_2239,N_2390);
nand U2454 (N_2454,N_2380,N_2314);
and U2455 (N_2455,N_2283,N_2348);
nor U2456 (N_2456,N_2320,N_2295);
and U2457 (N_2457,N_2238,N_2254);
nand U2458 (N_2458,N_2279,N_2357);
nor U2459 (N_2459,N_2392,N_2248);
or U2460 (N_2460,N_2350,N_2232);
and U2461 (N_2461,N_2365,N_2372);
and U2462 (N_2462,N_2324,N_2253);
and U2463 (N_2463,N_2315,N_2363);
or U2464 (N_2464,N_2366,N_2240);
and U2465 (N_2465,N_2231,N_2266);
nor U2466 (N_2466,N_2257,N_2250);
nand U2467 (N_2467,N_2287,N_2202);
nand U2468 (N_2468,N_2235,N_2216);
nor U2469 (N_2469,N_2370,N_2391);
nand U2470 (N_2470,N_2319,N_2273);
nor U2471 (N_2471,N_2339,N_2308);
nor U2472 (N_2472,N_2276,N_2271);
nor U2473 (N_2473,N_2376,N_2251);
or U2474 (N_2474,N_2383,N_2204);
or U2475 (N_2475,N_2343,N_2399);
nor U2476 (N_2476,N_2209,N_2396);
or U2477 (N_2477,N_2275,N_2297);
nor U2478 (N_2478,N_2282,N_2261);
nand U2479 (N_2479,N_2393,N_2200);
and U2480 (N_2480,N_2291,N_2219);
and U2481 (N_2481,N_2224,N_2317);
and U2482 (N_2482,N_2206,N_2352);
or U2483 (N_2483,N_2388,N_2386);
nand U2484 (N_2484,N_2345,N_2222);
or U2485 (N_2485,N_2264,N_2301);
and U2486 (N_2486,N_2203,N_2289);
nor U2487 (N_2487,N_2242,N_2371);
or U2488 (N_2488,N_2322,N_2351);
nand U2489 (N_2489,N_2292,N_2326);
and U2490 (N_2490,N_2394,N_2375);
and U2491 (N_2491,N_2262,N_2369);
and U2492 (N_2492,N_2214,N_2249);
nand U2493 (N_2493,N_2336,N_2361);
nand U2494 (N_2494,N_2347,N_2268);
or U2495 (N_2495,N_2318,N_2330);
nor U2496 (N_2496,N_2306,N_2293);
or U2497 (N_2497,N_2221,N_2201);
or U2498 (N_2498,N_2374,N_2298);
nand U2499 (N_2499,N_2341,N_2310);
nand U2500 (N_2500,N_2347,N_2393);
or U2501 (N_2501,N_2273,N_2364);
nor U2502 (N_2502,N_2292,N_2355);
nor U2503 (N_2503,N_2237,N_2294);
or U2504 (N_2504,N_2242,N_2298);
or U2505 (N_2505,N_2365,N_2333);
xor U2506 (N_2506,N_2305,N_2354);
nand U2507 (N_2507,N_2266,N_2372);
or U2508 (N_2508,N_2335,N_2229);
nor U2509 (N_2509,N_2339,N_2272);
nand U2510 (N_2510,N_2370,N_2289);
or U2511 (N_2511,N_2210,N_2325);
nand U2512 (N_2512,N_2228,N_2262);
nor U2513 (N_2513,N_2353,N_2226);
and U2514 (N_2514,N_2394,N_2281);
or U2515 (N_2515,N_2271,N_2208);
or U2516 (N_2516,N_2276,N_2316);
nor U2517 (N_2517,N_2310,N_2380);
nor U2518 (N_2518,N_2357,N_2216);
and U2519 (N_2519,N_2263,N_2229);
or U2520 (N_2520,N_2350,N_2229);
nand U2521 (N_2521,N_2367,N_2383);
nor U2522 (N_2522,N_2350,N_2360);
or U2523 (N_2523,N_2261,N_2218);
xnor U2524 (N_2524,N_2211,N_2299);
nand U2525 (N_2525,N_2207,N_2304);
nand U2526 (N_2526,N_2340,N_2357);
and U2527 (N_2527,N_2336,N_2250);
nand U2528 (N_2528,N_2391,N_2383);
and U2529 (N_2529,N_2239,N_2255);
or U2530 (N_2530,N_2313,N_2327);
or U2531 (N_2531,N_2391,N_2247);
and U2532 (N_2532,N_2368,N_2397);
and U2533 (N_2533,N_2351,N_2329);
xor U2534 (N_2534,N_2394,N_2222);
nand U2535 (N_2535,N_2241,N_2225);
and U2536 (N_2536,N_2242,N_2347);
nor U2537 (N_2537,N_2314,N_2213);
nor U2538 (N_2538,N_2351,N_2218);
and U2539 (N_2539,N_2294,N_2329);
nor U2540 (N_2540,N_2203,N_2260);
nor U2541 (N_2541,N_2309,N_2369);
or U2542 (N_2542,N_2368,N_2274);
and U2543 (N_2543,N_2229,N_2360);
nor U2544 (N_2544,N_2274,N_2237);
or U2545 (N_2545,N_2286,N_2308);
or U2546 (N_2546,N_2304,N_2282);
nor U2547 (N_2547,N_2293,N_2212);
nor U2548 (N_2548,N_2359,N_2365);
nand U2549 (N_2549,N_2380,N_2244);
nor U2550 (N_2550,N_2242,N_2372);
xor U2551 (N_2551,N_2274,N_2217);
xnor U2552 (N_2552,N_2236,N_2331);
or U2553 (N_2553,N_2320,N_2205);
nor U2554 (N_2554,N_2397,N_2365);
nand U2555 (N_2555,N_2298,N_2201);
or U2556 (N_2556,N_2337,N_2365);
nor U2557 (N_2557,N_2353,N_2271);
nor U2558 (N_2558,N_2377,N_2366);
or U2559 (N_2559,N_2328,N_2388);
nand U2560 (N_2560,N_2339,N_2226);
or U2561 (N_2561,N_2397,N_2275);
nor U2562 (N_2562,N_2330,N_2200);
nand U2563 (N_2563,N_2263,N_2236);
and U2564 (N_2564,N_2269,N_2233);
and U2565 (N_2565,N_2255,N_2269);
and U2566 (N_2566,N_2372,N_2302);
nand U2567 (N_2567,N_2265,N_2387);
xnor U2568 (N_2568,N_2284,N_2398);
or U2569 (N_2569,N_2354,N_2398);
nor U2570 (N_2570,N_2281,N_2237);
nand U2571 (N_2571,N_2344,N_2254);
nand U2572 (N_2572,N_2278,N_2370);
and U2573 (N_2573,N_2277,N_2315);
or U2574 (N_2574,N_2337,N_2307);
and U2575 (N_2575,N_2263,N_2285);
nor U2576 (N_2576,N_2348,N_2220);
and U2577 (N_2577,N_2331,N_2256);
nand U2578 (N_2578,N_2200,N_2270);
and U2579 (N_2579,N_2377,N_2373);
and U2580 (N_2580,N_2262,N_2263);
or U2581 (N_2581,N_2255,N_2248);
nand U2582 (N_2582,N_2356,N_2336);
or U2583 (N_2583,N_2365,N_2393);
nor U2584 (N_2584,N_2398,N_2346);
nor U2585 (N_2585,N_2341,N_2235);
or U2586 (N_2586,N_2251,N_2222);
and U2587 (N_2587,N_2341,N_2372);
nor U2588 (N_2588,N_2257,N_2211);
or U2589 (N_2589,N_2217,N_2253);
or U2590 (N_2590,N_2289,N_2233);
or U2591 (N_2591,N_2264,N_2206);
or U2592 (N_2592,N_2300,N_2382);
or U2593 (N_2593,N_2366,N_2394);
or U2594 (N_2594,N_2244,N_2353);
or U2595 (N_2595,N_2370,N_2384);
nor U2596 (N_2596,N_2346,N_2311);
nand U2597 (N_2597,N_2202,N_2251);
nand U2598 (N_2598,N_2247,N_2348);
nand U2599 (N_2599,N_2354,N_2364);
or U2600 (N_2600,N_2558,N_2497);
and U2601 (N_2601,N_2554,N_2427);
and U2602 (N_2602,N_2403,N_2498);
xor U2603 (N_2603,N_2541,N_2425);
or U2604 (N_2604,N_2408,N_2571);
or U2605 (N_2605,N_2527,N_2522);
and U2606 (N_2606,N_2583,N_2597);
and U2607 (N_2607,N_2595,N_2576);
or U2608 (N_2608,N_2422,N_2453);
and U2609 (N_2609,N_2437,N_2480);
or U2610 (N_2610,N_2441,N_2575);
and U2611 (N_2611,N_2410,N_2517);
nor U2612 (N_2612,N_2481,N_2566);
nand U2613 (N_2613,N_2516,N_2432);
or U2614 (N_2614,N_2569,N_2449);
nand U2615 (N_2615,N_2417,N_2539);
or U2616 (N_2616,N_2460,N_2452);
xnor U2617 (N_2617,N_2540,N_2526);
nand U2618 (N_2618,N_2489,N_2542);
nand U2619 (N_2619,N_2400,N_2486);
nor U2620 (N_2620,N_2545,N_2579);
and U2621 (N_2621,N_2471,N_2572);
nand U2622 (N_2622,N_2419,N_2520);
nor U2623 (N_2623,N_2538,N_2515);
nand U2624 (N_2624,N_2501,N_2530);
and U2625 (N_2625,N_2508,N_2531);
and U2626 (N_2626,N_2519,N_2567);
and U2627 (N_2627,N_2447,N_2411);
and U2628 (N_2628,N_2429,N_2555);
nand U2629 (N_2629,N_2568,N_2415);
and U2630 (N_2630,N_2465,N_2454);
nand U2631 (N_2631,N_2467,N_2534);
nand U2632 (N_2632,N_2469,N_2491);
nor U2633 (N_2633,N_2547,N_2433);
or U2634 (N_2634,N_2563,N_2536);
and U2635 (N_2635,N_2475,N_2533);
xor U2636 (N_2636,N_2412,N_2468);
or U2637 (N_2637,N_2406,N_2476);
nand U2638 (N_2638,N_2477,N_2496);
and U2639 (N_2639,N_2524,N_2559);
and U2640 (N_2640,N_2493,N_2591);
and U2641 (N_2641,N_2420,N_2435);
nor U2642 (N_2642,N_2470,N_2580);
or U2643 (N_2643,N_2443,N_2532);
nor U2644 (N_2644,N_2577,N_2506);
and U2645 (N_2645,N_2413,N_2528);
or U2646 (N_2646,N_2464,N_2593);
or U2647 (N_2647,N_2537,N_2431);
nor U2648 (N_2648,N_2535,N_2436);
nand U2649 (N_2649,N_2473,N_2502);
nand U2650 (N_2650,N_2484,N_2416);
and U2651 (N_2651,N_2434,N_2456);
nand U2652 (N_2652,N_2457,N_2500);
and U2653 (N_2653,N_2488,N_2439);
nand U2654 (N_2654,N_2483,N_2478);
and U2655 (N_2655,N_2551,N_2553);
or U2656 (N_2656,N_2585,N_2560);
xor U2657 (N_2657,N_2461,N_2564);
nand U2658 (N_2658,N_2414,N_2459);
and U2659 (N_2659,N_2523,N_2466);
or U2660 (N_2660,N_2582,N_2450);
and U2661 (N_2661,N_2548,N_2462);
and U2662 (N_2662,N_2598,N_2529);
or U2663 (N_2663,N_2556,N_2423);
nor U2664 (N_2664,N_2474,N_2552);
nand U2665 (N_2665,N_2581,N_2421);
nand U2666 (N_2666,N_2578,N_2505);
nor U2667 (N_2667,N_2512,N_2446);
nor U2668 (N_2668,N_2409,N_2587);
nand U2669 (N_2669,N_2599,N_2546);
nor U2670 (N_2670,N_2445,N_2424);
and U2671 (N_2671,N_2544,N_2574);
or U2672 (N_2672,N_2444,N_2549);
nand U2673 (N_2673,N_2402,N_2428);
nor U2674 (N_2674,N_2458,N_2588);
or U2675 (N_2675,N_2550,N_2573);
or U2676 (N_2676,N_2430,N_2504);
and U2677 (N_2677,N_2407,N_2592);
nand U2678 (N_2678,N_2570,N_2494);
nor U2679 (N_2679,N_2594,N_2525);
and U2680 (N_2680,N_2513,N_2586);
xor U2681 (N_2681,N_2485,N_2418);
and U2682 (N_2682,N_2404,N_2510);
and U2683 (N_2683,N_2514,N_2589);
and U2684 (N_2684,N_2590,N_2499);
or U2685 (N_2685,N_2451,N_2440);
or U2686 (N_2686,N_2490,N_2596);
nor U2687 (N_2687,N_2518,N_2448);
nand U2688 (N_2688,N_2584,N_2507);
nand U2689 (N_2689,N_2562,N_2487);
nor U2690 (N_2690,N_2561,N_2521);
nor U2691 (N_2691,N_2455,N_2472);
nand U2692 (N_2692,N_2482,N_2463);
and U2693 (N_2693,N_2543,N_2479);
and U2694 (N_2694,N_2503,N_2492);
or U2695 (N_2695,N_2442,N_2401);
nor U2696 (N_2696,N_2565,N_2438);
or U2697 (N_2697,N_2557,N_2405);
nand U2698 (N_2698,N_2495,N_2511);
and U2699 (N_2699,N_2509,N_2426);
nor U2700 (N_2700,N_2463,N_2529);
or U2701 (N_2701,N_2470,N_2506);
nand U2702 (N_2702,N_2497,N_2572);
nor U2703 (N_2703,N_2419,N_2561);
or U2704 (N_2704,N_2573,N_2479);
nand U2705 (N_2705,N_2567,N_2498);
nand U2706 (N_2706,N_2575,N_2520);
nand U2707 (N_2707,N_2499,N_2496);
nor U2708 (N_2708,N_2556,N_2572);
xor U2709 (N_2709,N_2546,N_2442);
nand U2710 (N_2710,N_2453,N_2405);
or U2711 (N_2711,N_2475,N_2556);
nand U2712 (N_2712,N_2482,N_2523);
or U2713 (N_2713,N_2539,N_2484);
nand U2714 (N_2714,N_2444,N_2594);
nor U2715 (N_2715,N_2564,N_2589);
or U2716 (N_2716,N_2526,N_2531);
and U2717 (N_2717,N_2514,N_2423);
and U2718 (N_2718,N_2587,N_2412);
and U2719 (N_2719,N_2532,N_2504);
and U2720 (N_2720,N_2521,N_2421);
and U2721 (N_2721,N_2480,N_2568);
and U2722 (N_2722,N_2421,N_2568);
or U2723 (N_2723,N_2569,N_2402);
and U2724 (N_2724,N_2484,N_2458);
xor U2725 (N_2725,N_2422,N_2562);
nand U2726 (N_2726,N_2518,N_2536);
and U2727 (N_2727,N_2544,N_2521);
or U2728 (N_2728,N_2431,N_2554);
or U2729 (N_2729,N_2425,N_2479);
nand U2730 (N_2730,N_2595,N_2539);
and U2731 (N_2731,N_2468,N_2493);
nand U2732 (N_2732,N_2486,N_2549);
nor U2733 (N_2733,N_2574,N_2514);
and U2734 (N_2734,N_2543,N_2489);
nor U2735 (N_2735,N_2506,N_2478);
and U2736 (N_2736,N_2591,N_2495);
and U2737 (N_2737,N_2546,N_2497);
or U2738 (N_2738,N_2535,N_2545);
nor U2739 (N_2739,N_2509,N_2467);
nand U2740 (N_2740,N_2493,N_2492);
or U2741 (N_2741,N_2458,N_2441);
or U2742 (N_2742,N_2547,N_2506);
and U2743 (N_2743,N_2514,N_2401);
or U2744 (N_2744,N_2449,N_2545);
nor U2745 (N_2745,N_2494,N_2476);
nor U2746 (N_2746,N_2535,N_2536);
and U2747 (N_2747,N_2434,N_2515);
nor U2748 (N_2748,N_2517,N_2533);
nand U2749 (N_2749,N_2553,N_2545);
nor U2750 (N_2750,N_2538,N_2457);
or U2751 (N_2751,N_2566,N_2543);
or U2752 (N_2752,N_2506,N_2462);
nor U2753 (N_2753,N_2462,N_2434);
and U2754 (N_2754,N_2575,N_2579);
nand U2755 (N_2755,N_2441,N_2545);
and U2756 (N_2756,N_2497,N_2439);
or U2757 (N_2757,N_2471,N_2561);
nor U2758 (N_2758,N_2504,N_2401);
nor U2759 (N_2759,N_2400,N_2431);
or U2760 (N_2760,N_2423,N_2467);
or U2761 (N_2761,N_2463,N_2471);
nand U2762 (N_2762,N_2583,N_2574);
and U2763 (N_2763,N_2480,N_2487);
nand U2764 (N_2764,N_2543,N_2410);
nand U2765 (N_2765,N_2537,N_2599);
and U2766 (N_2766,N_2503,N_2491);
nand U2767 (N_2767,N_2467,N_2571);
or U2768 (N_2768,N_2487,N_2553);
nand U2769 (N_2769,N_2564,N_2517);
or U2770 (N_2770,N_2513,N_2542);
nand U2771 (N_2771,N_2521,N_2502);
nand U2772 (N_2772,N_2447,N_2562);
nand U2773 (N_2773,N_2576,N_2498);
and U2774 (N_2774,N_2533,N_2555);
nand U2775 (N_2775,N_2525,N_2450);
nor U2776 (N_2776,N_2512,N_2519);
and U2777 (N_2777,N_2577,N_2442);
and U2778 (N_2778,N_2453,N_2528);
and U2779 (N_2779,N_2490,N_2595);
nand U2780 (N_2780,N_2524,N_2485);
nand U2781 (N_2781,N_2429,N_2595);
nand U2782 (N_2782,N_2450,N_2407);
or U2783 (N_2783,N_2501,N_2461);
nor U2784 (N_2784,N_2453,N_2455);
and U2785 (N_2785,N_2515,N_2457);
nand U2786 (N_2786,N_2442,N_2504);
nor U2787 (N_2787,N_2422,N_2568);
nor U2788 (N_2788,N_2516,N_2505);
nor U2789 (N_2789,N_2465,N_2592);
or U2790 (N_2790,N_2598,N_2411);
nor U2791 (N_2791,N_2500,N_2595);
and U2792 (N_2792,N_2569,N_2552);
nand U2793 (N_2793,N_2549,N_2563);
or U2794 (N_2794,N_2400,N_2501);
and U2795 (N_2795,N_2408,N_2509);
nand U2796 (N_2796,N_2509,N_2450);
nand U2797 (N_2797,N_2403,N_2411);
nor U2798 (N_2798,N_2499,N_2464);
nand U2799 (N_2799,N_2493,N_2437);
nand U2800 (N_2800,N_2706,N_2709);
and U2801 (N_2801,N_2679,N_2770);
nand U2802 (N_2802,N_2731,N_2760);
nand U2803 (N_2803,N_2718,N_2708);
xnor U2804 (N_2804,N_2705,N_2636);
or U2805 (N_2805,N_2632,N_2626);
nor U2806 (N_2806,N_2604,N_2689);
nor U2807 (N_2807,N_2752,N_2673);
nand U2808 (N_2808,N_2627,N_2733);
nand U2809 (N_2809,N_2790,N_2773);
nor U2810 (N_2810,N_2640,N_2743);
or U2811 (N_2811,N_2781,N_2786);
or U2812 (N_2812,N_2797,N_2623);
nand U2813 (N_2813,N_2625,N_2764);
or U2814 (N_2814,N_2602,N_2605);
or U2815 (N_2815,N_2700,N_2693);
nor U2816 (N_2816,N_2748,N_2724);
and U2817 (N_2817,N_2732,N_2739);
nand U2818 (N_2818,N_2682,N_2758);
nor U2819 (N_2819,N_2657,N_2792);
nand U2820 (N_2820,N_2698,N_2609);
nand U2821 (N_2821,N_2630,N_2727);
and U2822 (N_2822,N_2675,N_2753);
nor U2823 (N_2823,N_2777,N_2658);
and U2824 (N_2824,N_2791,N_2644);
or U2825 (N_2825,N_2769,N_2788);
nor U2826 (N_2826,N_2795,N_2738);
or U2827 (N_2827,N_2701,N_2650);
or U2828 (N_2828,N_2611,N_2717);
nor U2829 (N_2829,N_2639,N_2635);
nor U2830 (N_2830,N_2610,N_2685);
nand U2831 (N_2831,N_2697,N_2683);
and U2832 (N_2832,N_2735,N_2723);
nand U2833 (N_2833,N_2613,N_2745);
nor U2834 (N_2834,N_2695,N_2671);
and U2835 (N_2835,N_2710,N_2634);
and U2836 (N_2836,N_2798,N_2756);
and U2837 (N_2837,N_2734,N_2722);
nand U2838 (N_2838,N_2768,N_2621);
and U2839 (N_2839,N_2603,N_2742);
nor U2840 (N_2840,N_2656,N_2721);
nor U2841 (N_2841,N_2707,N_2755);
and U2842 (N_2842,N_2789,N_2651);
and U2843 (N_2843,N_2662,N_2641);
or U2844 (N_2844,N_2606,N_2772);
and U2845 (N_2845,N_2729,N_2703);
and U2846 (N_2846,N_2643,N_2600);
nand U2847 (N_2847,N_2746,N_2666);
xor U2848 (N_2848,N_2665,N_2784);
or U2849 (N_2849,N_2750,N_2648);
and U2850 (N_2850,N_2677,N_2642);
nor U2851 (N_2851,N_2796,N_2680);
or U2852 (N_2852,N_2749,N_2688);
nor U2853 (N_2853,N_2660,N_2687);
and U2854 (N_2854,N_2670,N_2765);
xnor U2855 (N_2855,N_2715,N_2653);
or U2856 (N_2856,N_2645,N_2669);
or U2857 (N_2857,N_2761,N_2637);
xnor U2858 (N_2858,N_2618,N_2607);
nand U2859 (N_2859,N_2751,N_2690);
nand U2860 (N_2860,N_2664,N_2667);
and U2861 (N_2861,N_2787,N_2766);
or U2862 (N_2862,N_2763,N_2785);
or U2863 (N_2863,N_2676,N_2713);
and U2864 (N_2864,N_2711,N_2681);
or U2865 (N_2865,N_2771,N_2759);
nor U2866 (N_2866,N_2646,N_2712);
nand U2867 (N_2867,N_2779,N_2612);
nor U2868 (N_2868,N_2730,N_2747);
or U2869 (N_2869,N_2654,N_2659);
or U2870 (N_2870,N_2633,N_2744);
and U2871 (N_2871,N_2601,N_2619);
or U2872 (N_2872,N_2622,N_2684);
or U2873 (N_2873,N_2793,N_2776);
or U2874 (N_2874,N_2617,N_2691);
nor U2875 (N_2875,N_2678,N_2741);
or U2876 (N_2876,N_2624,N_2620);
xor U2877 (N_2877,N_2736,N_2702);
nand U2878 (N_2878,N_2672,N_2615);
nand U2879 (N_2879,N_2794,N_2663);
nor U2880 (N_2880,N_2655,N_2647);
and U2881 (N_2881,N_2652,N_2696);
or U2882 (N_2882,N_2783,N_2686);
or U2883 (N_2883,N_2767,N_2614);
and U2884 (N_2884,N_2628,N_2699);
and U2885 (N_2885,N_2694,N_2714);
nor U2886 (N_2886,N_2780,N_2616);
xnor U2887 (N_2887,N_2754,N_2725);
nand U2888 (N_2888,N_2782,N_2774);
and U2889 (N_2889,N_2629,N_2638);
nor U2890 (N_2890,N_2726,N_2720);
and U2891 (N_2891,N_2757,N_2631);
or U2892 (N_2892,N_2674,N_2737);
nand U2893 (N_2893,N_2740,N_2799);
or U2894 (N_2894,N_2716,N_2704);
or U2895 (N_2895,N_2775,N_2661);
or U2896 (N_2896,N_2728,N_2692);
nand U2897 (N_2897,N_2719,N_2649);
and U2898 (N_2898,N_2762,N_2668);
or U2899 (N_2899,N_2608,N_2778);
nor U2900 (N_2900,N_2669,N_2615);
xor U2901 (N_2901,N_2705,N_2759);
nand U2902 (N_2902,N_2782,N_2716);
nand U2903 (N_2903,N_2773,N_2688);
or U2904 (N_2904,N_2691,N_2785);
and U2905 (N_2905,N_2774,N_2773);
or U2906 (N_2906,N_2669,N_2756);
nand U2907 (N_2907,N_2648,N_2700);
and U2908 (N_2908,N_2799,N_2658);
nand U2909 (N_2909,N_2720,N_2775);
or U2910 (N_2910,N_2683,N_2710);
or U2911 (N_2911,N_2639,N_2760);
and U2912 (N_2912,N_2624,N_2730);
nor U2913 (N_2913,N_2791,N_2655);
nor U2914 (N_2914,N_2620,N_2687);
nor U2915 (N_2915,N_2666,N_2681);
and U2916 (N_2916,N_2785,N_2740);
nand U2917 (N_2917,N_2762,N_2731);
and U2918 (N_2918,N_2735,N_2730);
and U2919 (N_2919,N_2704,N_2690);
nor U2920 (N_2920,N_2747,N_2718);
xor U2921 (N_2921,N_2664,N_2748);
nor U2922 (N_2922,N_2716,N_2744);
nand U2923 (N_2923,N_2796,N_2608);
and U2924 (N_2924,N_2732,N_2685);
or U2925 (N_2925,N_2707,N_2710);
or U2926 (N_2926,N_2670,N_2605);
nor U2927 (N_2927,N_2615,N_2732);
and U2928 (N_2928,N_2717,N_2640);
nand U2929 (N_2929,N_2712,N_2613);
nor U2930 (N_2930,N_2782,N_2749);
nand U2931 (N_2931,N_2625,N_2787);
nand U2932 (N_2932,N_2658,N_2601);
and U2933 (N_2933,N_2652,N_2663);
or U2934 (N_2934,N_2686,N_2735);
nand U2935 (N_2935,N_2617,N_2751);
or U2936 (N_2936,N_2718,N_2686);
and U2937 (N_2937,N_2750,N_2737);
nand U2938 (N_2938,N_2661,N_2793);
or U2939 (N_2939,N_2748,N_2707);
nand U2940 (N_2940,N_2662,N_2796);
and U2941 (N_2941,N_2661,N_2678);
nand U2942 (N_2942,N_2650,N_2622);
nor U2943 (N_2943,N_2721,N_2784);
and U2944 (N_2944,N_2715,N_2692);
nand U2945 (N_2945,N_2784,N_2782);
nand U2946 (N_2946,N_2625,N_2646);
nor U2947 (N_2947,N_2758,N_2716);
and U2948 (N_2948,N_2617,N_2736);
xnor U2949 (N_2949,N_2716,N_2614);
and U2950 (N_2950,N_2792,N_2661);
and U2951 (N_2951,N_2794,N_2712);
and U2952 (N_2952,N_2727,N_2670);
nand U2953 (N_2953,N_2606,N_2794);
and U2954 (N_2954,N_2678,N_2636);
nand U2955 (N_2955,N_2617,N_2694);
and U2956 (N_2956,N_2765,N_2690);
nor U2957 (N_2957,N_2751,N_2654);
nor U2958 (N_2958,N_2634,N_2786);
xor U2959 (N_2959,N_2642,N_2664);
and U2960 (N_2960,N_2656,N_2605);
and U2961 (N_2961,N_2750,N_2794);
nor U2962 (N_2962,N_2630,N_2667);
and U2963 (N_2963,N_2769,N_2629);
or U2964 (N_2964,N_2731,N_2655);
nor U2965 (N_2965,N_2611,N_2793);
and U2966 (N_2966,N_2783,N_2638);
or U2967 (N_2967,N_2768,N_2657);
or U2968 (N_2968,N_2632,N_2624);
and U2969 (N_2969,N_2610,N_2624);
or U2970 (N_2970,N_2695,N_2782);
nor U2971 (N_2971,N_2638,N_2630);
or U2972 (N_2972,N_2770,N_2775);
nand U2973 (N_2973,N_2790,N_2634);
and U2974 (N_2974,N_2771,N_2686);
nand U2975 (N_2975,N_2690,N_2650);
nand U2976 (N_2976,N_2655,N_2785);
nor U2977 (N_2977,N_2737,N_2693);
nor U2978 (N_2978,N_2689,N_2729);
or U2979 (N_2979,N_2611,N_2772);
nand U2980 (N_2980,N_2615,N_2734);
and U2981 (N_2981,N_2617,N_2659);
nor U2982 (N_2982,N_2718,N_2672);
and U2983 (N_2983,N_2794,N_2691);
nand U2984 (N_2984,N_2739,N_2617);
nand U2985 (N_2985,N_2662,N_2625);
and U2986 (N_2986,N_2703,N_2750);
or U2987 (N_2987,N_2719,N_2653);
nand U2988 (N_2988,N_2630,N_2734);
xnor U2989 (N_2989,N_2657,N_2756);
or U2990 (N_2990,N_2761,N_2729);
or U2991 (N_2991,N_2729,N_2606);
nand U2992 (N_2992,N_2705,N_2785);
nor U2993 (N_2993,N_2660,N_2678);
nand U2994 (N_2994,N_2792,N_2738);
nand U2995 (N_2995,N_2682,N_2710);
or U2996 (N_2996,N_2721,N_2799);
or U2997 (N_2997,N_2612,N_2742);
and U2998 (N_2998,N_2602,N_2655);
or U2999 (N_2999,N_2708,N_2799);
and UO_0 (O_0,N_2822,N_2839);
and UO_1 (O_1,N_2854,N_2857);
nor UO_2 (O_2,N_2877,N_2969);
nand UO_3 (O_3,N_2992,N_2812);
nor UO_4 (O_4,N_2830,N_2801);
nor UO_5 (O_5,N_2970,N_2913);
nand UO_6 (O_6,N_2880,N_2894);
and UO_7 (O_7,N_2864,N_2820);
nand UO_8 (O_8,N_2907,N_2829);
nand UO_9 (O_9,N_2999,N_2917);
nand UO_10 (O_10,N_2901,N_2995);
nor UO_11 (O_11,N_2998,N_2942);
nand UO_12 (O_12,N_2902,N_2978);
nand UO_13 (O_13,N_2938,N_2851);
or UO_14 (O_14,N_2911,N_2900);
nand UO_15 (O_15,N_2834,N_2989);
or UO_16 (O_16,N_2955,N_2856);
or UO_17 (O_17,N_2879,N_2804);
nor UO_18 (O_18,N_2840,N_2946);
nor UO_19 (O_19,N_2965,N_2975);
or UO_20 (O_20,N_2843,N_2990);
nand UO_21 (O_21,N_2903,N_2884);
and UO_22 (O_22,N_2943,N_2929);
nand UO_23 (O_23,N_2906,N_2927);
nor UO_24 (O_24,N_2944,N_2997);
nor UO_25 (O_25,N_2850,N_2899);
and UO_26 (O_26,N_2859,N_2832);
or UO_27 (O_27,N_2984,N_2972);
nor UO_28 (O_28,N_2996,N_2953);
nand UO_29 (O_29,N_2883,N_2865);
nand UO_30 (O_30,N_2905,N_2823);
nand UO_31 (O_31,N_2861,N_2808);
nor UO_32 (O_32,N_2814,N_2968);
and UO_33 (O_33,N_2920,N_2961);
nor UO_34 (O_34,N_2803,N_2979);
and UO_35 (O_35,N_2841,N_2921);
or UO_36 (O_36,N_2912,N_2811);
and UO_37 (O_37,N_2909,N_2915);
or UO_38 (O_38,N_2826,N_2891);
and UO_39 (O_39,N_2849,N_2806);
and UO_40 (O_40,N_2816,N_2982);
nand UO_41 (O_41,N_2827,N_2926);
or UO_42 (O_42,N_2828,N_2948);
nand UO_43 (O_43,N_2870,N_2817);
and UO_44 (O_44,N_2874,N_2838);
or UO_45 (O_45,N_2813,N_2872);
or UO_46 (O_46,N_2881,N_2833);
nand UO_47 (O_47,N_2868,N_2976);
or UO_48 (O_48,N_2888,N_2924);
nand UO_49 (O_49,N_2914,N_2886);
and UO_50 (O_50,N_2896,N_2980);
nor UO_51 (O_51,N_2985,N_2964);
and UO_52 (O_52,N_2956,N_2889);
or UO_53 (O_53,N_2876,N_2986);
or UO_54 (O_54,N_2957,N_2895);
and UO_55 (O_55,N_2893,N_2866);
nor UO_56 (O_56,N_2918,N_2802);
nor UO_57 (O_57,N_2950,N_2878);
nand UO_58 (O_58,N_2869,N_2935);
nor UO_59 (O_59,N_2885,N_2815);
or UO_60 (O_60,N_2852,N_2867);
xnor UO_61 (O_61,N_2819,N_2977);
or UO_62 (O_62,N_2846,N_2898);
xor UO_63 (O_63,N_2871,N_2892);
nand UO_64 (O_64,N_2988,N_2821);
and UO_65 (O_65,N_2937,N_2940);
or UO_66 (O_66,N_2862,N_2919);
nor UO_67 (O_67,N_2983,N_2951);
or UO_68 (O_68,N_2936,N_2994);
nand UO_69 (O_69,N_2845,N_2908);
and UO_70 (O_70,N_2863,N_2939);
xnor UO_71 (O_71,N_2991,N_2923);
nor UO_72 (O_72,N_2875,N_2810);
or UO_73 (O_73,N_2831,N_2932);
and UO_74 (O_74,N_2860,N_2855);
or UO_75 (O_75,N_2809,N_2945);
and UO_76 (O_76,N_2933,N_2910);
nand UO_77 (O_77,N_2847,N_2922);
xnor UO_78 (O_78,N_2800,N_2837);
and UO_79 (O_79,N_2818,N_2966);
or UO_80 (O_80,N_2887,N_2882);
nand UO_81 (O_81,N_2952,N_2897);
and UO_82 (O_82,N_2842,N_2904);
nor UO_83 (O_83,N_2930,N_2805);
nand UO_84 (O_84,N_2835,N_2825);
and UO_85 (O_85,N_2973,N_2853);
or UO_86 (O_86,N_2934,N_2971);
or UO_87 (O_87,N_2949,N_2958);
or UO_88 (O_88,N_2963,N_2993);
nand UO_89 (O_89,N_2916,N_2925);
nand UO_90 (O_90,N_2960,N_2974);
nand UO_91 (O_91,N_2890,N_2959);
and UO_92 (O_92,N_2844,N_2824);
nand UO_93 (O_93,N_2941,N_2848);
nand UO_94 (O_94,N_2807,N_2954);
nand UO_95 (O_95,N_2931,N_2928);
or UO_96 (O_96,N_2967,N_2873);
or UO_97 (O_97,N_2987,N_2962);
and UO_98 (O_98,N_2981,N_2858);
and UO_99 (O_99,N_2947,N_2836);
nand UO_100 (O_100,N_2901,N_2877);
nor UO_101 (O_101,N_2809,N_2868);
or UO_102 (O_102,N_2849,N_2857);
nor UO_103 (O_103,N_2966,N_2971);
and UO_104 (O_104,N_2828,N_2954);
nand UO_105 (O_105,N_2972,N_2858);
nand UO_106 (O_106,N_2831,N_2973);
nand UO_107 (O_107,N_2848,N_2806);
nor UO_108 (O_108,N_2842,N_2908);
nand UO_109 (O_109,N_2834,N_2952);
nand UO_110 (O_110,N_2821,N_2975);
or UO_111 (O_111,N_2824,N_2936);
and UO_112 (O_112,N_2843,N_2805);
nand UO_113 (O_113,N_2978,N_2944);
and UO_114 (O_114,N_2909,N_2822);
and UO_115 (O_115,N_2936,N_2972);
nor UO_116 (O_116,N_2864,N_2808);
or UO_117 (O_117,N_2932,N_2981);
and UO_118 (O_118,N_2947,N_2935);
nand UO_119 (O_119,N_2926,N_2896);
nor UO_120 (O_120,N_2831,N_2817);
nand UO_121 (O_121,N_2872,N_2969);
nand UO_122 (O_122,N_2856,N_2975);
and UO_123 (O_123,N_2820,N_2939);
nor UO_124 (O_124,N_2985,N_2954);
and UO_125 (O_125,N_2959,N_2818);
or UO_126 (O_126,N_2807,N_2937);
or UO_127 (O_127,N_2909,N_2853);
and UO_128 (O_128,N_2951,N_2961);
or UO_129 (O_129,N_2945,N_2860);
and UO_130 (O_130,N_2907,N_2863);
and UO_131 (O_131,N_2876,N_2886);
or UO_132 (O_132,N_2863,N_2876);
nor UO_133 (O_133,N_2947,N_2823);
xor UO_134 (O_134,N_2877,N_2832);
and UO_135 (O_135,N_2909,N_2992);
and UO_136 (O_136,N_2899,N_2901);
or UO_137 (O_137,N_2914,N_2852);
nor UO_138 (O_138,N_2927,N_2815);
nand UO_139 (O_139,N_2969,N_2997);
or UO_140 (O_140,N_2935,N_2916);
nor UO_141 (O_141,N_2912,N_2844);
or UO_142 (O_142,N_2830,N_2845);
and UO_143 (O_143,N_2986,N_2803);
nor UO_144 (O_144,N_2960,N_2910);
and UO_145 (O_145,N_2920,N_2877);
nand UO_146 (O_146,N_2812,N_2855);
nor UO_147 (O_147,N_2876,N_2930);
and UO_148 (O_148,N_2874,N_2944);
and UO_149 (O_149,N_2928,N_2884);
nand UO_150 (O_150,N_2892,N_2881);
xor UO_151 (O_151,N_2811,N_2935);
and UO_152 (O_152,N_2934,N_2858);
and UO_153 (O_153,N_2965,N_2883);
nor UO_154 (O_154,N_2878,N_2850);
nand UO_155 (O_155,N_2816,N_2824);
nor UO_156 (O_156,N_2999,N_2891);
nand UO_157 (O_157,N_2833,N_2911);
or UO_158 (O_158,N_2898,N_2981);
nor UO_159 (O_159,N_2855,N_2942);
and UO_160 (O_160,N_2843,N_2884);
nor UO_161 (O_161,N_2829,N_2999);
nand UO_162 (O_162,N_2860,N_2886);
or UO_163 (O_163,N_2809,N_2926);
nor UO_164 (O_164,N_2890,N_2923);
nand UO_165 (O_165,N_2946,N_2830);
nand UO_166 (O_166,N_2966,N_2936);
and UO_167 (O_167,N_2859,N_2978);
or UO_168 (O_168,N_2985,N_2848);
and UO_169 (O_169,N_2819,N_2836);
xor UO_170 (O_170,N_2845,N_2937);
nand UO_171 (O_171,N_2902,N_2810);
xnor UO_172 (O_172,N_2922,N_2807);
or UO_173 (O_173,N_2841,N_2883);
nand UO_174 (O_174,N_2800,N_2908);
nor UO_175 (O_175,N_2997,N_2833);
or UO_176 (O_176,N_2915,N_2946);
and UO_177 (O_177,N_2994,N_2911);
or UO_178 (O_178,N_2987,N_2931);
or UO_179 (O_179,N_2901,N_2956);
or UO_180 (O_180,N_2906,N_2978);
or UO_181 (O_181,N_2942,N_2835);
or UO_182 (O_182,N_2816,N_2954);
nor UO_183 (O_183,N_2969,N_2880);
or UO_184 (O_184,N_2818,N_2864);
nor UO_185 (O_185,N_2957,N_2910);
or UO_186 (O_186,N_2921,N_2830);
or UO_187 (O_187,N_2890,N_2810);
nand UO_188 (O_188,N_2919,N_2821);
nor UO_189 (O_189,N_2822,N_2875);
and UO_190 (O_190,N_2964,N_2882);
and UO_191 (O_191,N_2817,N_2892);
and UO_192 (O_192,N_2983,N_2889);
nand UO_193 (O_193,N_2859,N_2878);
nand UO_194 (O_194,N_2945,N_2851);
nor UO_195 (O_195,N_2831,N_2933);
nand UO_196 (O_196,N_2937,N_2907);
nand UO_197 (O_197,N_2956,N_2980);
and UO_198 (O_198,N_2853,N_2810);
nor UO_199 (O_199,N_2981,N_2859);
or UO_200 (O_200,N_2852,N_2918);
or UO_201 (O_201,N_2929,N_2967);
or UO_202 (O_202,N_2979,N_2916);
nand UO_203 (O_203,N_2884,N_2958);
and UO_204 (O_204,N_2977,N_2979);
nor UO_205 (O_205,N_2978,N_2937);
nand UO_206 (O_206,N_2970,N_2879);
nor UO_207 (O_207,N_2878,N_2893);
nor UO_208 (O_208,N_2981,N_2871);
or UO_209 (O_209,N_2969,N_2911);
nand UO_210 (O_210,N_2926,N_2807);
and UO_211 (O_211,N_2916,N_2893);
and UO_212 (O_212,N_2801,N_2874);
nand UO_213 (O_213,N_2968,N_2872);
or UO_214 (O_214,N_2915,N_2825);
nor UO_215 (O_215,N_2895,N_2894);
or UO_216 (O_216,N_2870,N_2916);
nand UO_217 (O_217,N_2867,N_2969);
or UO_218 (O_218,N_2960,N_2917);
nor UO_219 (O_219,N_2853,N_2917);
or UO_220 (O_220,N_2871,N_2979);
and UO_221 (O_221,N_2875,N_2974);
nor UO_222 (O_222,N_2965,N_2964);
and UO_223 (O_223,N_2948,N_2901);
or UO_224 (O_224,N_2841,N_2895);
and UO_225 (O_225,N_2945,N_2850);
or UO_226 (O_226,N_2811,N_2888);
xor UO_227 (O_227,N_2943,N_2874);
or UO_228 (O_228,N_2922,N_2937);
or UO_229 (O_229,N_2861,N_2909);
and UO_230 (O_230,N_2877,N_2925);
nor UO_231 (O_231,N_2981,N_2810);
nand UO_232 (O_232,N_2993,N_2930);
and UO_233 (O_233,N_2876,N_2852);
or UO_234 (O_234,N_2945,N_2827);
or UO_235 (O_235,N_2810,N_2865);
nor UO_236 (O_236,N_2879,N_2871);
nand UO_237 (O_237,N_2925,N_2853);
nor UO_238 (O_238,N_2986,N_2972);
nand UO_239 (O_239,N_2807,N_2987);
nand UO_240 (O_240,N_2898,N_2830);
nor UO_241 (O_241,N_2862,N_2831);
or UO_242 (O_242,N_2834,N_2908);
nor UO_243 (O_243,N_2957,N_2845);
nand UO_244 (O_244,N_2846,N_2892);
nor UO_245 (O_245,N_2865,N_2994);
xnor UO_246 (O_246,N_2853,N_2878);
and UO_247 (O_247,N_2939,N_2880);
and UO_248 (O_248,N_2856,N_2922);
nand UO_249 (O_249,N_2967,N_2972);
nand UO_250 (O_250,N_2909,N_2919);
or UO_251 (O_251,N_2945,N_2922);
nor UO_252 (O_252,N_2810,N_2868);
and UO_253 (O_253,N_2913,N_2881);
or UO_254 (O_254,N_2957,N_2815);
or UO_255 (O_255,N_2905,N_2883);
and UO_256 (O_256,N_2980,N_2897);
nand UO_257 (O_257,N_2972,N_2839);
and UO_258 (O_258,N_2853,N_2944);
and UO_259 (O_259,N_2826,N_2856);
and UO_260 (O_260,N_2876,N_2807);
nor UO_261 (O_261,N_2818,N_2918);
nand UO_262 (O_262,N_2882,N_2892);
and UO_263 (O_263,N_2884,N_2983);
or UO_264 (O_264,N_2972,N_2863);
nand UO_265 (O_265,N_2995,N_2829);
or UO_266 (O_266,N_2804,N_2980);
nor UO_267 (O_267,N_2979,N_2816);
nand UO_268 (O_268,N_2967,N_2966);
nor UO_269 (O_269,N_2836,N_2808);
nand UO_270 (O_270,N_2857,N_2926);
nand UO_271 (O_271,N_2869,N_2930);
nand UO_272 (O_272,N_2987,N_2826);
xnor UO_273 (O_273,N_2814,N_2994);
or UO_274 (O_274,N_2839,N_2948);
nor UO_275 (O_275,N_2876,N_2978);
nand UO_276 (O_276,N_2918,N_2854);
xor UO_277 (O_277,N_2934,N_2807);
and UO_278 (O_278,N_2891,N_2896);
or UO_279 (O_279,N_2896,N_2952);
nand UO_280 (O_280,N_2930,N_2954);
and UO_281 (O_281,N_2853,N_2970);
and UO_282 (O_282,N_2952,N_2820);
nand UO_283 (O_283,N_2814,N_2969);
or UO_284 (O_284,N_2868,N_2954);
and UO_285 (O_285,N_2905,N_2934);
nor UO_286 (O_286,N_2988,N_2893);
or UO_287 (O_287,N_2889,N_2920);
nor UO_288 (O_288,N_2986,N_2877);
or UO_289 (O_289,N_2915,N_2990);
nor UO_290 (O_290,N_2984,N_2929);
or UO_291 (O_291,N_2819,N_2867);
and UO_292 (O_292,N_2946,N_2895);
nand UO_293 (O_293,N_2911,N_2946);
xnor UO_294 (O_294,N_2801,N_2816);
nor UO_295 (O_295,N_2924,N_2951);
and UO_296 (O_296,N_2973,N_2870);
xor UO_297 (O_297,N_2983,N_2897);
and UO_298 (O_298,N_2851,N_2885);
or UO_299 (O_299,N_2957,N_2981);
nand UO_300 (O_300,N_2821,N_2851);
or UO_301 (O_301,N_2805,N_2902);
nor UO_302 (O_302,N_2915,N_2988);
and UO_303 (O_303,N_2954,N_2896);
or UO_304 (O_304,N_2972,N_2868);
or UO_305 (O_305,N_2879,N_2933);
and UO_306 (O_306,N_2824,N_2973);
and UO_307 (O_307,N_2803,N_2872);
and UO_308 (O_308,N_2838,N_2906);
nor UO_309 (O_309,N_2960,N_2916);
and UO_310 (O_310,N_2954,N_2999);
nand UO_311 (O_311,N_2839,N_2852);
nor UO_312 (O_312,N_2834,N_2896);
and UO_313 (O_313,N_2835,N_2875);
nand UO_314 (O_314,N_2985,N_2935);
nor UO_315 (O_315,N_2942,N_2808);
nor UO_316 (O_316,N_2804,N_2835);
nor UO_317 (O_317,N_2960,N_2928);
or UO_318 (O_318,N_2852,N_2830);
and UO_319 (O_319,N_2829,N_2819);
or UO_320 (O_320,N_2928,N_2839);
and UO_321 (O_321,N_2964,N_2811);
nand UO_322 (O_322,N_2860,N_2803);
nand UO_323 (O_323,N_2874,N_2806);
and UO_324 (O_324,N_2805,N_2994);
xor UO_325 (O_325,N_2875,N_2876);
nand UO_326 (O_326,N_2931,N_2968);
and UO_327 (O_327,N_2989,N_2855);
or UO_328 (O_328,N_2972,N_2949);
nand UO_329 (O_329,N_2977,N_2857);
and UO_330 (O_330,N_2985,N_2902);
nand UO_331 (O_331,N_2991,N_2999);
and UO_332 (O_332,N_2801,N_2825);
and UO_333 (O_333,N_2994,N_2879);
nor UO_334 (O_334,N_2861,N_2819);
nor UO_335 (O_335,N_2839,N_2926);
and UO_336 (O_336,N_2888,N_2973);
nor UO_337 (O_337,N_2958,N_2945);
nand UO_338 (O_338,N_2985,N_2934);
nor UO_339 (O_339,N_2875,N_2847);
and UO_340 (O_340,N_2849,N_2980);
or UO_341 (O_341,N_2904,N_2955);
and UO_342 (O_342,N_2881,N_2978);
or UO_343 (O_343,N_2854,N_2848);
nand UO_344 (O_344,N_2933,N_2874);
or UO_345 (O_345,N_2832,N_2861);
xnor UO_346 (O_346,N_2919,N_2949);
and UO_347 (O_347,N_2845,N_2898);
nand UO_348 (O_348,N_2936,N_2886);
nor UO_349 (O_349,N_2975,N_2876);
nand UO_350 (O_350,N_2994,N_2966);
and UO_351 (O_351,N_2876,N_2961);
and UO_352 (O_352,N_2835,N_2956);
and UO_353 (O_353,N_2808,N_2885);
or UO_354 (O_354,N_2924,N_2911);
and UO_355 (O_355,N_2974,N_2897);
nand UO_356 (O_356,N_2955,N_2868);
nand UO_357 (O_357,N_2847,N_2953);
and UO_358 (O_358,N_2848,N_2819);
nor UO_359 (O_359,N_2896,N_2829);
nor UO_360 (O_360,N_2878,N_2928);
nand UO_361 (O_361,N_2854,N_2871);
nor UO_362 (O_362,N_2938,N_2934);
nor UO_363 (O_363,N_2963,N_2857);
nor UO_364 (O_364,N_2843,N_2853);
or UO_365 (O_365,N_2997,N_2862);
and UO_366 (O_366,N_2896,N_2929);
nand UO_367 (O_367,N_2817,N_2871);
nor UO_368 (O_368,N_2972,N_2855);
nand UO_369 (O_369,N_2959,N_2989);
or UO_370 (O_370,N_2994,N_2836);
and UO_371 (O_371,N_2882,N_2942);
xnor UO_372 (O_372,N_2936,N_2984);
nor UO_373 (O_373,N_2867,N_2920);
nand UO_374 (O_374,N_2905,N_2973);
nor UO_375 (O_375,N_2820,N_2980);
nand UO_376 (O_376,N_2994,N_2940);
xor UO_377 (O_377,N_2899,N_2869);
or UO_378 (O_378,N_2974,N_2892);
and UO_379 (O_379,N_2811,N_2982);
and UO_380 (O_380,N_2940,N_2962);
and UO_381 (O_381,N_2903,N_2932);
nor UO_382 (O_382,N_2822,N_2952);
and UO_383 (O_383,N_2924,N_2821);
or UO_384 (O_384,N_2865,N_2982);
nand UO_385 (O_385,N_2884,N_2924);
nor UO_386 (O_386,N_2980,N_2869);
or UO_387 (O_387,N_2942,N_2925);
or UO_388 (O_388,N_2862,N_2918);
and UO_389 (O_389,N_2827,N_2844);
and UO_390 (O_390,N_2954,N_2967);
and UO_391 (O_391,N_2862,N_2815);
nand UO_392 (O_392,N_2959,N_2847);
or UO_393 (O_393,N_2959,N_2849);
or UO_394 (O_394,N_2971,N_2865);
or UO_395 (O_395,N_2809,N_2874);
xor UO_396 (O_396,N_2916,N_2816);
and UO_397 (O_397,N_2828,N_2842);
nor UO_398 (O_398,N_2926,N_2989);
nand UO_399 (O_399,N_2804,N_2999);
and UO_400 (O_400,N_2895,N_2808);
and UO_401 (O_401,N_2863,N_2995);
and UO_402 (O_402,N_2915,N_2994);
nor UO_403 (O_403,N_2896,N_2934);
and UO_404 (O_404,N_2862,N_2935);
nor UO_405 (O_405,N_2816,N_2874);
nor UO_406 (O_406,N_2913,N_2961);
and UO_407 (O_407,N_2921,N_2811);
nor UO_408 (O_408,N_2945,N_2848);
and UO_409 (O_409,N_2920,N_2885);
or UO_410 (O_410,N_2827,N_2931);
and UO_411 (O_411,N_2972,N_2964);
nor UO_412 (O_412,N_2994,N_2970);
nor UO_413 (O_413,N_2890,N_2896);
or UO_414 (O_414,N_2859,N_2940);
or UO_415 (O_415,N_2915,N_2984);
nor UO_416 (O_416,N_2812,N_2933);
and UO_417 (O_417,N_2871,N_2988);
and UO_418 (O_418,N_2809,N_2899);
and UO_419 (O_419,N_2981,N_2921);
or UO_420 (O_420,N_2954,N_2806);
nand UO_421 (O_421,N_2887,N_2961);
nor UO_422 (O_422,N_2922,N_2862);
nand UO_423 (O_423,N_2922,N_2999);
or UO_424 (O_424,N_2849,N_2845);
nor UO_425 (O_425,N_2801,N_2903);
and UO_426 (O_426,N_2821,N_2866);
and UO_427 (O_427,N_2874,N_2889);
and UO_428 (O_428,N_2864,N_2981);
and UO_429 (O_429,N_2992,N_2919);
and UO_430 (O_430,N_2952,N_2922);
nand UO_431 (O_431,N_2950,N_2920);
or UO_432 (O_432,N_2881,N_2920);
and UO_433 (O_433,N_2973,N_2812);
and UO_434 (O_434,N_2896,N_2849);
or UO_435 (O_435,N_2994,N_2989);
nor UO_436 (O_436,N_2862,N_2965);
or UO_437 (O_437,N_2921,N_2951);
nor UO_438 (O_438,N_2837,N_2918);
nor UO_439 (O_439,N_2905,N_2972);
and UO_440 (O_440,N_2878,N_2819);
and UO_441 (O_441,N_2951,N_2845);
or UO_442 (O_442,N_2954,N_2865);
nor UO_443 (O_443,N_2818,N_2962);
nor UO_444 (O_444,N_2802,N_2958);
or UO_445 (O_445,N_2919,N_2976);
nand UO_446 (O_446,N_2953,N_2969);
xor UO_447 (O_447,N_2871,N_2902);
nor UO_448 (O_448,N_2803,N_2822);
nor UO_449 (O_449,N_2877,N_2823);
nand UO_450 (O_450,N_2909,N_2989);
nor UO_451 (O_451,N_2804,N_2891);
or UO_452 (O_452,N_2800,N_2954);
nand UO_453 (O_453,N_2847,N_2885);
nor UO_454 (O_454,N_2900,N_2863);
and UO_455 (O_455,N_2951,N_2972);
nand UO_456 (O_456,N_2808,N_2876);
nand UO_457 (O_457,N_2957,N_2908);
nor UO_458 (O_458,N_2844,N_2959);
and UO_459 (O_459,N_2933,N_2946);
nand UO_460 (O_460,N_2920,N_2842);
xor UO_461 (O_461,N_2977,N_2823);
xnor UO_462 (O_462,N_2996,N_2943);
nand UO_463 (O_463,N_2830,N_2893);
and UO_464 (O_464,N_2897,N_2966);
nor UO_465 (O_465,N_2951,N_2906);
nand UO_466 (O_466,N_2827,N_2996);
nor UO_467 (O_467,N_2982,N_2831);
and UO_468 (O_468,N_2933,N_2972);
nor UO_469 (O_469,N_2899,N_2946);
nor UO_470 (O_470,N_2892,N_2920);
nand UO_471 (O_471,N_2879,N_2861);
nand UO_472 (O_472,N_2864,N_2933);
and UO_473 (O_473,N_2854,N_2990);
nor UO_474 (O_474,N_2885,N_2902);
or UO_475 (O_475,N_2812,N_2962);
and UO_476 (O_476,N_2881,N_2976);
and UO_477 (O_477,N_2902,N_2941);
or UO_478 (O_478,N_2846,N_2875);
nor UO_479 (O_479,N_2914,N_2854);
and UO_480 (O_480,N_2980,N_2821);
and UO_481 (O_481,N_2822,N_2979);
nor UO_482 (O_482,N_2933,N_2987);
nor UO_483 (O_483,N_2840,N_2823);
nand UO_484 (O_484,N_2931,N_2808);
or UO_485 (O_485,N_2893,N_2873);
nor UO_486 (O_486,N_2976,N_2885);
and UO_487 (O_487,N_2924,N_2936);
xor UO_488 (O_488,N_2857,N_2833);
or UO_489 (O_489,N_2875,N_2993);
nor UO_490 (O_490,N_2892,N_2995);
or UO_491 (O_491,N_2958,N_2891);
nor UO_492 (O_492,N_2992,N_2999);
and UO_493 (O_493,N_2960,N_2955);
xor UO_494 (O_494,N_2984,N_2974);
xor UO_495 (O_495,N_2953,N_2862);
or UO_496 (O_496,N_2968,N_2967);
nor UO_497 (O_497,N_2855,N_2996);
nor UO_498 (O_498,N_2948,N_2832);
and UO_499 (O_499,N_2959,N_2889);
endmodule