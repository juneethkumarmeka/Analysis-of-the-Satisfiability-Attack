module basic_1500_15000_2000_5_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_268,In_1156);
and U1 (N_1,In_1086,In_71);
nand U2 (N_2,In_783,In_1246);
nand U3 (N_3,In_453,In_951);
xnor U4 (N_4,In_290,In_1336);
nand U5 (N_5,In_807,In_657);
or U6 (N_6,In_53,In_140);
nand U7 (N_7,In_407,In_690);
nand U8 (N_8,In_991,In_653);
nand U9 (N_9,In_232,In_808);
or U10 (N_10,In_1461,In_1280);
or U11 (N_11,In_100,In_239);
and U12 (N_12,In_874,In_1266);
nand U13 (N_13,In_1173,In_1359);
and U14 (N_14,In_174,In_405);
nand U15 (N_15,In_1157,In_1161);
nand U16 (N_16,In_236,In_1357);
nor U17 (N_17,In_257,In_1333);
nor U18 (N_18,In_686,In_785);
and U19 (N_19,In_856,In_1282);
nor U20 (N_20,In_162,In_312);
or U21 (N_21,In_203,In_86);
or U22 (N_22,In_637,In_17);
nor U23 (N_23,In_635,In_885);
or U24 (N_24,In_883,In_612);
nor U25 (N_25,In_1315,In_1164);
nor U26 (N_26,In_1253,In_1181);
nand U27 (N_27,In_1002,In_1220);
nand U28 (N_28,In_551,In_25);
or U29 (N_29,In_795,In_869);
and U30 (N_30,In_24,In_650);
or U31 (N_31,In_1343,In_1327);
nand U32 (N_32,In_459,In_786);
nand U33 (N_33,In_226,In_1152);
or U34 (N_34,In_1414,In_1473);
nor U35 (N_35,In_995,In_1175);
or U36 (N_36,In_1272,In_1234);
and U37 (N_37,In_1393,In_332);
and U38 (N_38,In_594,In_397);
nand U39 (N_39,In_97,In_1205);
nand U40 (N_40,In_1021,In_321);
or U41 (N_41,In_1119,In_942);
and U42 (N_42,In_306,In_730);
nor U43 (N_43,In_633,In_1305);
or U44 (N_44,In_1385,In_171);
nand U45 (N_45,In_1478,In_393);
nand U46 (N_46,In_648,In_725);
and U47 (N_47,In_1448,In_1381);
nand U48 (N_48,In_1443,In_875);
nor U49 (N_49,In_994,In_779);
and U50 (N_50,In_978,In_1212);
or U51 (N_51,In_1050,In_514);
and U52 (N_52,In_178,In_1129);
nand U53 (N_53,In_406,In_1241);
nand U54 (N_54,In_982,In_917);
or U55 (N_55,In_112,In_679);
and U56 (N_56,In_32,In_992);
nor U57 (N_57,In_173,In_894);
nand U58 (N_58,In_1043,In_699);
or U59 (N_59,In_1260,In_1293);
and U60 (N_60,In_930,In_614);
xor U61 (N_61,In_673,In_664);
and U62 (N_62,In_1047,In_1436);
nand U63 (N_63,In_1072,In_844);
nor U64 (N_64,In_77,In_237);
nand U65 (N_65,In_150,In_1070);
nand U66 (N_66,In_52,In_202);
or U67 (N_67,In_1178,In_1243);
nand U68 (N_68,In_1471,In_928);
or U69 (N_69,In_1362,In_1488);
nor U70 (N_70,In_1341,In_1142);
nand U71 (N_71,In_955,In_1318);
nor U72 (N_72,In_1494,In_608);
and U73 (N_73,In_265,In_766);
nor U74 (N_74,In_889,In_80);
nor U75 (N_75,In_880,In_146);
or U76 (N_76,In_1447,In_910);
nand U77 (N_77,In_584,In_768);
and U78 (N_78,In_1289,In_1466);
nand U79 (N_79,In_967,In_461);
nor U80 (N_80,In_1171,In_909);
nand U81 (N_81,In_1369,In_139);
and U82 (N_82,In_1268,In_697);
nor U83 (N_83,In_313,In_1223);
or U84 (N_84,In_383,In_1027);
or U85 (N_85,In_297,In_552);
or U86 (N_86,In_570,In_247);
xnor U87 (N_87,In_1373,In_1022);
and U88 (N_88,In_610,In_661);
nor U89 (N_89,In_677,In_634);
or U90 (N_90,In_1041,In_182);
and U91 (N_91,In_1138,In_255);
or U92 (N_92,In_548,In_742);
nor U93 (N_93,In_1109,In_51);
or U94 (N_94,In_1489,In_451);
and U95 (N_95,In_1299,In_1163);
or U96 (N_96,In_1019,In_330);
and U97 (N_97,In_1190,In_912);
or U98 (N_98,In_1232,In_1079);
nor U99 (N_99,In_342,In_349);
xor U100 (N_100,In_1356,In_390);
nand U101 (N_101,In_719,In_274);
nor U102 (N_102,In_138,In_621);
nand U103 (N_103,In_573,In_1186);
nor U104 (N_104,In_263,In_241);
and U105 (N_105,In_127,In_827);
or U106 (N_106,In_746,In_1035);
nor U107 (N_107,In_1355,In_1487);
nand U108 (N_108,In_901,In_936);
or U109 (N_109,In_974,In_423);
or U110 (N_110,In_137,In_1049);
or U111 (N_111,In_749,In_1255);
nand U112 (N_112,In_945,In_997);
nor U113 (N_113,In_5,In_606);
nor U114 (N_114,In_771,In_1291);
and U115 (N_115,In_483,In_74);
nand U116 (N_116,In_281,In_1402);
and U117 (N_117,In_553,In_660);
nor U118 (N_118,In_222,In_817);
and U119 (N_119,In_683,In_476);
and U120 (N_120,In_12,In_152);
and U121 (N_121,In_1475,In_916);
and U122 (N_122,In_1,In_1092);
nor U123 (N_123,In_1094,In_975);
nor U124 (N_124,In_198,In_4);
nor U125 (N_125,In_1238,In_1184);
nand U126 (N_126,In_854,In_859);
nor U127 (N_127,In_1498,In_791);
and U128 (N_128,In_161,In_591);
or U129 (N_129,In_401,In_1206);
nand U130 (N_130,In_744,In_356);
and U131 (N_131,In_1392,In_1115);
nor U132 (N_132,In_72,In_82);
and U133 (N_133,In_214,In_1245);
nor U134 (N_134,In_1329,In_495);
and U135 (N_135,In_234,In_1091);
nor U136 (N_136,In_1066,In_258);
or U137 (N_137,In_961,In_688);
or U138 (N_138,In_1382,In_1139);
nor U139 (N_139,In_491,In_141);
nand U140 (N_140,In_564,In_309);
nor U141 (N_141,In_111,In_799);
nor U142 (N_142,In_1000,In_177);
nand U143 (N_143,In_831,In_1100);
nand U144 (N_144,In_520,In_478);
nand U145 (N_145,In_529,In_430);
or U146 (N_146,In_388,In_615);
nand U147 (N_147,In_1445,In_156);
xnor U148 (N_148,In_1203,In_632);
or U149 (N_149,In_1344,In_337);
nand U150 (N_150,In_877,In_1411);
nor U151 (N_151,In_1044,In_607);
nand U152 (N_152,In_1389,In_1211);
and U153 (N_153,In_801,In_1217);
nand U154 (N_154,In_48,In_30);
nor U155 (N_155,In_809,In_1406);
nand U156 (N_156,In_474,In_1176);
and U157 (N_157,In_240,In_1192);
or U158 (N_158,In_344,In_1400);
and U159 (N_159,In_946,In_754);
or U160 (N_160,In_1365,In_1360);
nand U161 (N_161,In_829,In_745);
nand U162 (N_162,In_1010,In_578);
nand U163 (N_163,In_521,In_914);
nor U164 (N_164,In_1292,In_1391);
or U165 (N_165,In_1383,In_184);
and U166 (N_166,In_1170,In_1463);
nor U167 (N_167,In_557,In_467);
and U168 (N_168,In_42,In_1014);
and U169 (N_169,In_618,In_409);
nor U170 (N_170,In_1148,In_1482);
nand U171 (N_171,In_921,In_675);
and U172 (N_172,In_443,In_480);
nand U173 (N_173,In_286,In_549);
nand U174 (N_174,In_1024,In_130);
or U175 (N_175,In_1427,In_1226);
nor U176 (N_176,In_1177,In_19);
nor U177 (N_177,In_1194,In_66);
nor U178 (N_178,In_373,In_119);
and U179 (N_179,In_229,In_698);
or U180 (N_180,In_887,In_282);
nor U181 (N_181,In_1229,In_1334);
nor U182 (N_182,In_643,In_92);
nand U183 (N_183,In_1440,In_1368);
or U184 (N_184,In_1009,In_1419);
and U185 (N_185,In_1252,In_194);
nand U186 (N_186,In_362,In_800);
and U187 (N_187,In_1030,In_825);
nor U188 (N_188,In_903,In_1317);
and U189 (N_189,In_1496,In_711);
and U190 (N_190,In_398,In_1444);
and U191 (N_191,In_68,In_195);
nor U192 (N_192,In_276,In_568);
nor U193 (N_193,In_539,In_843);
or U194 (N_194,In_213,In_419);
nand U195 (N_195,In_506,In_485);
nor U196 (N_196,In_235,In_33);
nor U197 (N_197,In_1042,In_693);
and U198 (N_198,In_810,In_837);
nand U199 (N_199,In_728,In_335);
nand U200 (N_200,In_1080,In_970);
nor U201 (N_201,In_798,In_849);
xor U202 (N_202,In_986,In_598);
nor U203 (N_203,In_492,In_1429);
or U204 (N_204,In_538,In_31);
nor U205 (N_205,In_600,In_1283);
nor U206 (N_206,In_76,In_987);
or U207 (N_207,In_1430,In_1218);
nand U208 (N_208,In_781,In_210);
or U209 (N_209,In_283,In_326);
or U210 (N_210,In_189,In_753);
or U211 (N_211,In_1040,In_700);
nor U212 (N_212,In_583,In_1201);
or U213 (N_213,In_750,In_45);
and U214 (N_214,In_852,In_338);
nor U215 (N_215,In_1418,In_1497);
nor U216 (N_216,In_314,In_590);
or U217 (N_217,In_888,In_731);
nor U218 (N_218,In_627,In_1055);
nor U219 (N_219,In_1099,In_120);
nand U220 (N_220,In_709,In_864);
and U221 (N_221,In_823,In_463);
nor U222 (N_222,In_1376,In_935);
or U223 (N_223,In_28,In_1209);
nor U224 (N_224,In_319,In_145);
or U225 (N_225,In_10,In_1451);
or U226 (N_226,In_1169,In_687);
and U227 (N_227,In_300,In_1380);
and U228 (N_228,In_1254,In_1480);
nor U229 (N_229,In_715,In_1345);
nand U230 (N_230,In_116,In_915);
and U231 (N_231,In_1278,In_70);
nor U232 (N_232,In_895,In_1256);
nand U233 (N_233,In_1339,In_842);
or U234 (N_234,In_1367,In_372);
and U235 (N_235,In_508,In_109);
nor U236 (N_236,In_206,In_269);
or U237 (N_237,In_878,In_611);
or U238 (N_238,In_18,In_1250);
nor U239 (N_239,In_998,In_11);
and U240 (N_240,In_681,In_976);
or U241 (N_241,In_380,In_248);
nor U242 (N_242,In_117,In_62);
or U243 (N_243,In_432,In_1191);
nand U244 (N_244,In_190,In_710);
or U245 (N_245,In_481,In_1207);
or U246 (N_246,In_47,In_528);
nor U247 (N_247,In_543,In_1200);
or U248 (N_248,In_1063,In_91);
nor U249 (N_249,In_850,In_365);
or U250 (N_250,In_378,In_299);
nor U251 (N_251,In_487,In_431);
nand U252 (N_252,In_1455,In_617);
nand U253 (N_253,In_587,In_426);
and U254 (N_254,In_550,In_706);
xnor U255 (N_255,In_75,In_579);
and U256 (N_256,In_567,In_1265);
nor U257 (N_257,In_447,In_1294);
nor U258 (N_258,In_848,In_158);
nand U259 (N_259,In_1490,In_597);
nand U260 (N_260,In_905,In_651);
and U261 (N_261,In_1015,In_1076);
and U262 (N_262,In_756,In_84);
nand U263 (N_263,In_641,In_1111);
and U264 (N_264,In_165,In_381);
or U265 (N_265,In_1090,In_948);
nand U266 (N_266,In_176,In_1249);
and U267 (N_267,In_1240,In_1467);
or U268 (N_268,In_1350,In_736);
and U269 (N_269,In_1059,In_435);
and U270 (N_270,In_294,In_1384);
and U271 (N_271,In_737,In_656);
and U272 (N_272,In_892,In_1133);
and U273 (N_273,In_369,In_384);
nor U274 (N_274,In_302,In_609);
or U275 (N_275,In_1394,In_622);
or U276 (N_276,In_104,In_1395);
nor U277 (N_277,In_839,In_628);
nor U278 (N_278,In_180,In_454);
or U279 (N_279,In_544,In_1031);
or U280 (N_280,In_93,In_322);
and U281 (N_281,In_586,In_505);
nand U282 (N_282,In_713,In_834);
and U283 (N_283,In_954,In_1352);
nand U284 (N_284,In_493,In_14);
nor U285 (N_285,In_392,In_26);
nand U286 (N_286,In_703,In_1012);
xnor U287 (N_287,In_947,In_863);
and U288 (N_288,In_1311,In_164);
nand U289 (N_289,In_264,In_1037);
nand U290 (N_290,In_36,In_1065);
or U291 (N_291,In_973,In_762);
nor U292 (N_292,In_1262,In_1363);
and U293 (N_293,In_1263,In_207);
nor U294 (N_294,In_375,In_882);
nand U295 (N_295,In_347,In_1499);
xnor U296 (N_296,In_167,In_1314);
nor U297 (N_297,In_437,In_537);
and U298 (N_298,In_1147,In_64);
nor U299 (N_299,In_1008,In_1005);
nand U300 (N_300,In_1013,In_811);
and U301 (N_301,In_655,In_1468);
nand U302 (N_302,In_1259,In_865);
or U303 (N_303,In_1308,In_941);
and U304 (N_304,In_971,In_488);
or U305 (N_305,In_106,In_1273);
nand U306 (N_306,In_1144,In_1174);
xnor U307 (N_307,In_1306,In_284);
and U308 (N_308,In_751,In_1085);
nor U309 (N_309,In_833,In_1088);
nor U310 (N_310,In_761,In_99);
and U311 (N_311,In_556,In_475);
nand U312 (N_312,In_1056,In_354);
xnor U313 (N_313,In_630,In_1183);
and U314 (N_314,In_867,In_603);
nor U315 (N_315,In_272,In_1302);
nor U316 (N_316,In_266,In_359);
or U317 (N_317,In_1348,In_417);
and U318 (N_318,In_562,In_379);
or U319 (N_319,In_331,In_580);
nand U320 (N_320,In_1208,In_102);
nand U321 (N_321,In_434,In_386);
nor U322 (N_322,In_1004,In_1123);
nor U323 (N_323,In_355,In_1185);
nand U324 (N_324,In_1449,In_471);
nand U325 (N_325,In_1247,In_1319);
nor U326 (N_326,In_462,In_1151);
or U327 (N_327,In_812,In_403);
or U328 (N_328,In_1387,In_1146);
nand U329 (N_329,In_950,In_1310);
or U330 (N_330,In_866,In_918);
nor U331 (N_331,In_394,In_1285);
nand U332 (N_332,In_58,In_374);
nand U333 (N_333,In_636,In_1264);
nor U334 (N_334,In_1267,In_1269);
and U335 (N_335,In_1470,In_1286);
xor U336 (N_336,In_327,In_1347);
nor U337 (N_337,In_1081,In_740);
and U338 (N_338,In_211,In_328);
or U339 (N_339,In_270,In_1126);
nand U340 (N_340,In_1162,In_581);
nor U341 (N_341,In_1221,In_1195);
nand U342 (N_342,In_712,In_530);
or U343 (N_343,In_696,In_1160);
nor U344 (N_344,In_1016,In_873);
nor U345 (N_345,In_911,In_3);
and U346 (N_346,In_90,In_490);
and U347 (N_347,In_503,In_1069);
and U348 (N_348,In_765,In_814);
nand U349 (N_349,In_1154,In_1346);
nand U350 (N_350,In_962,In_399);
and U351 (N_351,In_1073,In_1068);
and U352 (N_352,In_6,In_1023);
nand U353 (N_353,In_774,In_535);
nand U354 (N_354,In_575,In_340);
and U355 (N_355,In_204,In_1075);
or U356 (N_356,In_1197,In_1460);
or U357 (N_357,In_254,In_589);
or U358 (N_358,In_1295,In_1454);
nand U359 (N_359,In_620,In_1242);
nand U360 (N_360,In_671,In_1231);
nand U361 (N_361,In_436,In_943);
or U362 (N_362,In_420,In_183);
nand U363 (N_363,In_22,In_7);
or U364 (N_364,In_1053,In_563);
and U365 (N_365,In_46,In_747);
nor U366 (N_366,In_225,In_1420);
nor U367 (N_367,In_1301,In_1052);
and U368 (N_368,In_1116,In_1407);
or U369 (N_369,In_1127,In_716);
nor U370 (N_370,In_1431,In_40);
nand U371 (N_371,In_536,In_107);
or U372 (N_372,In_124,In_1364);
or U373 (N_373,In_507,In_1219);
or U374 (N_374,In_1222,In_69);
or U375 (N_375,In_217,In_1017);
or U376 (N_376,In_416,In_1189);
nor U377 (N_377,In_411,In_191);
nor U378 (N_378,In_1408,In_574);
or U379 (N_379,In_1335,In_244);
or U380 (N_380,In_1300,In_775);
nor U381 (N_381,In_625,In_305);
and U382 (N_382,In_125,In_701);
and U383 (N_383,In_502,In_350);
and U384 (N_384,In_1456,In_855);
and U385 (N_385,In_275,In_168);
or U386 (N_386,In_1216,In_246);
and U387 (N_387,In_816,In_65);
and U388 (N_388,In_1464,In_857);
and U389 (N_389,In_477,In_870);
nor U390 (N_390,In_512,In_1337);
and U391 (N_391,In_924,In_38);
nand U392 (N_392,In_1312,In_1424);
nand U393 (N_393,In_619,In_793);
nand U394 (N_394,In_50,In_694);
or U395 (N_395,In_1297,In_1484);
nor U396 (N_396,In_148,In_1492);
nor U397 (N_397,In_320,In_1150);
and U398 (N_398,In_197,In_638);
nor U399 (N_399,In_440,In_972);
or U400 (N_400,In_218,In_446);
nand U401 (N_401,In_85,In_554);
nor U402 (N_402,In_692,In_1491);
and U403 (N_403,In_1134,In_259);
or U404 (N_404,In_1304,In_593);
nor U405 (N_405,In_1415,In_67);
xor U406 (N_406,In_832,In_1349);
or U407 (N_407,In_588,In_789);
or U408 (N_408,In_517,In_389);
or U409 (N_409,In_219,In_223);
and U410 (N_410,In_851,In_469);
nor U411 (N_411,In_1034,In_377);
nand U412 (N_412,In_602,In_893);
nor U413 (N_413,In_441,In_876);
xor U414 (N_414,In_187,In_558);
or U415 (N_415,In_402,In_134);
or U416 (N_416,In_1159,In_640);
nor U417 (N_417,In_1379,In_346);
nor U418 (N_418,In_101,In_722);
and U419 (N_419,In_665,In_1257);
or U420 (N_420,In_123,In_316);
nand U421 (N_421,In_813,In_1244);
nand U422 (N_422,In_1130,In_1450);
or U423 (N_423,In_199,In_623);
or U424 (N_424,In_601,In_726);
nor U425 (N_425,In_1153,In_1353);
and U426 (N_426,In_404,In_639);
or U427 (N_427,In_1323,In_797);
or U428 (N_428,In_464,In_245);
and U429 (N_429,In_105,In_37);
or U430 (N_430,In_663,In_324);
nand U431 (N_431,In_999,In_1168);
nor U432 (N_432,In_279,In_958);
nor U433 (N_433,In_662,In_498);
and U434 (N_434,In_996,In_794);
and U435 (N_435,In_691,In_121);
and U436 (N_436,In_395,In_391);
or U437 (N_437,In_1199,In_776);
and U438 (N_438,In_427,In_522);
nand U439 (N_439,In_702,In_513);
nor U440 (N_440,In_678,In_1340);
and U441 (N_441,In_757,In_43);
nand U442 (N_442,In_1105,In_186);
xnor U443 (N_443,In_1366,In_1481);
nor U444 (N_444,In_718,In_136);
nand U445 (N_445,In_790,In_460);
nand U446 (N_446,In_1103,In_767);
and U447 (N_447,In_1439,In_504);
or U448 (N_448,In_175,In_547);
nor U449 (N_449,In_1288,In_624);
and U450 (N_450,In_1377,In_592);
and U451 (N_451,In_34,In_647);
nor U452 (N_452,In_868,In_16);
nor U453 (N_453,In_1422,In_1128);
and U454 (N_454,In_1277,In_1321);
nand U455 (N_455,In_1413,In_1077);
and U456 (N_456,In_271,In_1082);
nand U457 (N_457,In_1108,In_79);
nor U458 (N_458,In_201,In_29);
or U459 (N_459,In_285,In_497);
and U460 (N_460,In_500,In_805);
and U461 (N_461,In_287,In_1230);
nor U462 (N_462,In_489,In_1370);
or U463 (N_463,In_576,In_748);
or U464 (N_464,In_585,In_366);
nor U465 (N_465,In_527,In_523);
nand U466 (N_466,In_1320,In_993);
or U467 (N_467,In_988,In_329);
nor U468 (N_468,In_23,In_689);
nor U469 (N_469,In_674,In_645);
and U470 (N_470,In_308,In_913);
nor U471 (N_471,In_1074,In_1452);
and U472 (N_472,In_343,In_114);
or U473 (N_473,In_953,In_129);
nor U474 (N_474,In_1224,In_1372);
and U475 (N_475,In_1071,In_8);
and U476 (N_476,In_778,In_519);
or U477 (N_477,In_1064,In_468);
nand U478 (N_478,In_904,In_1417);
xor U479 (N_479,In_1110,In_115);
nand U480 (N_480,In_561,In_452);
and U481 (N_481,In_1061,In_1172);
nand U482 (N_482,In_1358,In_1296);
nor U483 (N_483,In_1479,In_752);
nand U484 (N_484,In_1274,In_231);
and U485 (N_485,In_243,In_667);
nor U486 (N_486,In_929,In_387);
nand U487 (N_487,In_172,In_473);
and U488 (N_488,In_458,In_1087);
and U489 (N_489,In_1095,In_723);
or U490 (N_490,In_193,In_605);
or U491 (N_491,In_1107,In_658);
and U492 (N_492,In_1290,In_1437);
nor U493 (N_493,In_1316,In_542);
nand U494 (N_494,In_1214,In_1330);
nand U495 (N_495,In_295,In_919);
nor U496 (N_496,In_414,In_524);
or U497 (N_497,In_815,In_896);
nor U498 (N_498,In_1029,In_261);
or U499 (N_499,In_1118,In_442);
and U500 (N_500,In_734,In_169);
nor U501 (N_501,In_965,In_940);
and U502 (N_502,In_1281,In_931);
xnor U503 (N_503,In_1298,In_298);
or U504 (N_504,In_163,In_858);
and U505 (N_505,In_1438,In_1442);
and U506 (N_506,In_154,In_293);
and U507 (N_507,In_456,In_780);
nand U508 (N_508,In_15,In_1018);
and U509 (N_509,In_759,In_1182);
nor U510 (N_510,In_385,In_773);
or U511 (N_511,In_1276,In_415);
nor U512 (N_512,In_361,In_1404);
or U513 (N_513,In_249,In_631);
nor U514 (N_514,In_932,In_1403);
and U515 (N_515,In_131,In_421);
or U516 (N_516,In_371,In_1058);
or U517 (N_517,In_804,In_981);
or U518 (N_518,In_902,In_835);
or U519 (N_519,In_1046,In_13);
or U520 (N_520,In_1453,In_135);
nor U521 (N_521,In_358,In_1233);
or U522 (N_522,In_1441,In_224);
nand U523 (N_523,In_59,In_920);
and U524 (N_524,In_339,In_672);
nand U525 (N_525,In_820,In_484);
nor U526 (N_526,In_989,In_352);
and U527 (N_527,In_729,In_55);
nor U528 (N_528,In_56,In_63);
and U529 (N_529,In_1477,In_57);
and U530 (N_530,In_1006,In_705);
xnor U531 (N_531,In_310,In_979);
or U532 (N_532,In_153,In_466);
nand U533 (N_533,In_1067,In_360);
or U534 (N_534,In_185,In_457);
nand U535 (N_535,In_763,In_1434);
nand U536 (N_536,In_1104,In_196);
nor U537 (N_537,In_1033,In_534);
nor U538 (N_538,In_291,In_438);
nand U539 (N_539,In_311,In_367);
nand U540 (N_540,In_1140,In_1235);
nand U541 (N_541,In_907,In_410);
and U542 (N_542,In_532,In_846);
or U543 (N_543,In_555,In_1432);
and U544 (N_544,In_1007,In_1045);
and U545 (N_545,In_215,In_652);
nand U546 (N_546,In_984,In_1057);
and U547 (N_547,In_155,In_1378);
and U548 (N_548,In_629,In_482);
and U549 (N_549,In_668,In_826);
nor U550 (N_550,In_307,In_1210);
nor U551 (N_551,In_1398,In_792);
or U552 (N_552,In_301,In_1275);
nor U553 (N_553,In_368,In_144);
xnor U554 (N_554,In_853,In_828);
and U555 (N_555,In_1493,In_1457);
or U556 (N_556,In_960,In_418);
xor U557 (N_557,In_1399,In_1435);
nand U558 (N_558,In_260,In_83);
nor U559 (N_559,In_784,In_228);
and U560 (N_560,In_739,In_424);
nor U561 (N_561,In_891,In_566);
nor U562 (N_562,In_44,In_108);
and U563 (N_563,In_871,In_1428);
and U564 (N_564,In_1465,In_450);
nor U565 (N_565,In_1462,In_304);
nor U566 (N_566,In_35,In_518);
and U567 (N_567,In_1131,In_1322);
and U568 (N_568,In_1188,In_782);
or U569 (N_569,In_830,In_596);
nor U570 (N_570,In_1228,In_925);
nand U571 (N_571,In_160,In_755);
nand U572 (N_572,In_879,In_1412);
or U573 (N_573,In_267,In_433);
nor U574 (N_574,In_428,In_1351);
and U575 (N_575,In_1374,In_1409);
xor U576 (N_576,In_444,In_714);
and U577 (N_577,In_1405,In_990);
or U578 (N_578,In_934,In_670);
nor U579 (N_579,In_1287,In_351);
or U580 (N_580,In_1303,In_230);
nand U581 (N_581,In_205,In_78);
xor U582 (N_582,In_959,In_1446);
nand U583 (N_583,In_2,In_1410);
or U584 (N_584,In_1401,In_323);
and U585 (N_585,In_1248,In_98);
xor U586 (N_586,In_242,In_938);
or U587 (N_587,In_408,In_1472);
and U588 (N_588,In_806,In_872);
nor U589 (N_589,In_315,In_1193);
nand U590 (N_590,In_897,In_1196);
nor U591 (N_591,In_250,In_727);
nor U592 (N_592,In_81,In_209);
nand U593 (N_593,In_192,In_821);
nand U594 (N_594,In_221,In_1328);
nor U595 (N_595,In_142,In_496);
or U596 (N_596,In_862,In_1307);
nand U597 (N_597,In_208,In_533);
nor U598 (N_598,In_516,In_1032);
and U599 (N_599,In_515,In_838);
and U600 (N_600,In_1239,In_707);
nand U601 (N_601,In_251,In_642);
nor U602 (N_602,In_724,In_649);
and U603 (N_603,In_1198,In_803);
and U604 (N_604,In_717,In_819);
or U605 (N_605,In_318,In_1397);
and U606 (N_606,In_118,In_1026);
and U607 (N_607,In_836,In_559);
nand U608 (N_608,In_1135,In_341);
nand U609 (N_609,In_704,In_531);
nand U610 (N_610,In_983,In_933);
nor U611 (N_611,In_1114,In_818);
and U612 (N_612,In_1279,In_479);
xor U613 (N_613,In_439,In_73);
nand U614 (N_614,In_1020,In_616);
or U615 (N_615,In_345,In_1469);
nand U616 (N_616,In_968,In_720);
and U617 (N_617,In_1261,In_1225);
or U618 (N_618,In_470,In_1141);
nor U619 (N_619,In_1120,In_1476);
nor U620 (N_620,In_695,In_526);
xnor U621 (N_621,In_1324,In_1001);
nor U622 (N_622,In_325,In_565);
nand U623 (N_623,In_1121,In_1251);
or U624 (N_624,In_220,In_499);
and U625 (N_625,In_743,In_1106);
or U626 (N_626,In_1227,In_448);
nor U627 (N_627,In_412,In_511);
xor U628 (N_628,In_1204,In_676);
nor U629 (N_629,In_9,In_944);
or U630 (N_630,In_777,In_772);
or U631 (N_631,In_899,In_796);
xnor U632 (N_632,In_1158,In_980);
or U633 (N_633,In_802,In_333);
nand U634 (N_634,In_238,In_400);
nor U635 (N_635,In_1331,In_472);
and U636 (N_636,In_1423,In_1145);
nor U637 (N_637,In_200,In_845);
nor U638 (N_638,In_20,In_541);
and U639 (N_639,In_760,In_87);
or U640 (N_640,In_509,In_1474);
nand U641 (N_641,In_1011,In_1483);
nor U642 (N_642,In_425,In_525);
or U643 (N_643,In_1102,In_1124);
nor U644 (N_644,In_721,In_1060);
nand U645 (N_645,In_143,In_288);
nand U646 (N_646,In_1271,In_166);
or U647 (N_647,In_1396,In_88);
and U648 (N_648,In_787,In_963);
or U649 (N_649,In_1179,In_357);
or U650 (N_650,In_577,In_1495);
or U651 (N_651,In_122,In_1338);
and U652 (N_652,In_1143,In_157);
or U653 (N_653,In_133,In_1433);
and U654 (N_654,In_273,In_769);
nor U655 (N_655,In_733,In_599);
nand U656 (N_656,In_1003,In_60);
or U657 (N_657,In_110,In_571);
nor U658 (N_658,In_1078,In_1325);
or U659 (N_659,In_1136,In_1084);
and U660 (N_660,In_1309,In_494);
and U661 (N_661,In_212,In_1125);
or U662 (N_662,In_604,In_582);
nor U663 (N_663,In_429,In_27);
or U664 (N_664,In_1089,In_906);
and U665 (N_665,In_860,In_501);
nand U666 (N_666,In_1421,In_278);
nor U667 (N_667,In_939,In_708);
and U668 (N_668,In_277,In_977);
nor U669 (N_669,In_455,In_886);
nor U670 (N_670,In_465,In_666);
nor U671 (N_671,In_1167,In_292);
or U672 (N_672,In_735,In_303);
nand U673 (N_673,In_1101,In_376);
or U674 (N_674,In_1459,In_1117);
nor U675 (N_675,In_985,In_900);
and U676 (N_676,In_824,In_741);
and U677 (N_677,In_216,In_545);
or U678 (N_678,In_1390,In_89);
and U679 (N_679,In_445,In_1155);
nand U680 (N_680,In_1486,In_952);
and U681 (N_681,In_1165,In_569);
nand U682 (N_682,In_926,In_788);
nor U683 (N_683,In_1051,In_1096);
or U684 (N_684,In_669,In_764);
nor U685 (N_685,In_94,In_1093);
or U686 (N_686,In_1361,In_54);
nand U687 (N_687,In_966,In_188);
xor U688 (N_688,In_646,In_927);
or U689 (N_689,In_956,In_103);
or U690 (N_690,In_336,In_334);
or U691 (N_691,In_1332,In_1313);
or U692 (N_692,In_758,In_1237);
nor U693 (N_693,In_113,In_626);
nand U694 (N_694,In_1284,In_841);
nand U695 (N_695,In_1166,In_159);
nor U696 (N_696,In_39,In_890);
nor U697 (N_697,In_181,In_1375);
or U698 (N_698,In_685,In_1180);
nand U699 (N_699,In_847,In_1485);
or U700 (N_700,In_898,In_227);
and U701 (N_701,In_1097,In_1122);
and U702 (N_702,In_1425,In_128);
nor U703 (N_703,In_1036,In_95);
or U704 (N_704,In_280,In_1326);
or U705 (N_705,In_510,In_348);
or U706 (N_706,In_560,In_1458);
and U707 (N_707,In_1149,In_654);
nor U708 (N_708,In_964,In_149);
nand U709 (N_709,In_252,In_1137);
or U710 (N_710,In_1416,In_96);
nor U711 (N_711,In_126,In_1028);
nand U712 (N_712,In_1054,In_363);
and U713 (N_713,In_922,In_49);
nand U714 (N_714,In_147,In_317);
nor U715 (N_715,In_1371,In_861);
nand U716 (N_716,In_822,In_923);
and U717 (N_717,In_969,In_908);
and U718 (N_718,In_179,In_680);
or U719 (N_719,In_949,In_1132);
and U720 (N_720,In_540,In_1215);
nand U721 (N_721,In_233,In_1062);
nor U722 (N_722,In_21,In_1113);
and U723 (N_723,In_937,In_364);
nand U724 (N_724,In_840,In_1098);
and U725 (N_725,In_353,In_738);
nand U726 (N_726,In_1354,In_289);
nor U727 (N_727,In_1038,In_449);
and U728 (N_728,In_486,In_256);
or U729 (N_729,In_1342,In_1202);
nand U730 (N_730,In_132,In_884);
nor U731 (N_731,In_684,In_41);
nand U732 (N_732,In_1236,In_682);
nand U733 (N_733,In_0,In_572);
and U734 (N_734,In_644,In_613);
nor U735 (N_735,In_61,In_546);
nand U736 (N_736,In_1270,In_1048);
nand U737 (N_737,In_396,In_1426);
nand U738 (N_738,In_659,In_1187);
or U739 (N_739,In_1112,In_170);
and U740 (N_740,In_370,In_296);
or U741 (N_741,In_413,In_151);
or U742 (N_742,In_1213,In_1083);
or U743 (N_743,In_732,In_595);
nand U744 (N_744,In_1258,In_253);
and U745 (N_745,In_1388,In_1039);
nand U746 (N_746,In_957,In_422);
nor U747 (N_747,In_1386,In_770);
nor U748 (N_748,In_1025,In_382);
or U749 (N_749,In_881,In_262);
nand U750 (N_750,In_1069,In_1456);
nand U751 (N_751,In_1191,In_1221);
nand U752 (N_752,In_294,In_1018);
and U753 (N_753,In_455,In_1114);
nor U754 (N_754,In_734,In_483);
nand U755 (N_755,In_810,In_456);
nor U756 (N_756,In_1122,In_1476);
and U757 (N_757,In_1213,In_664);
or U758 (N_758,In_826,In_122);
or U759 (N_759,In_273,In_1074);
nand U760 (N_760,In_513,In_1075);
nand U761 (N_761,In_172,In_10);
or U762 (N_762,In_920,In_168);
or U763 (N_763,In_1176,In_383);
and U764 (N_764,In_936,In_222);
or U765 (N_765,In_1174,In_1294);
nor U766 (N_766,In_429,In_462);
and U767 (N_767,In_1409,In_787);
nand U768 (N_768,In_573,In_734);
xnor U769 (N_769,In_1077,In_1110);
nor U770 (N_770,In_617,In_1467);
or U771 (N_771,In_1220,In_1321);
or U772 (N_772,In_713,In_1116);
nor U773 (N_773,In_120,In_94);
nand U774 (N_774,In_1447,In_980);
and U775 (N_775,In_1148,In_1139);
nand U776 (N_776,In_1255,In_636);
nand U777 (N_777,In_1050,In_464);
or U778 (N_778,In_948,In_618);
or U779 (N_779,In_1218,In_155);
or U780 (N_780,In_1215,In_1348);
nand U781 (N_781,In_1268,In_646);
nand U782 (N_782,In_627,In_332);
nor U783 (N_783,In_1277,In_537);
nor U784 (N_784,In_438,In_322);
and U785 (N_785,In_294,In_266);
or U786 (N_786,In_949,In_832);
and U787 (N_787,In_1160,In_407);
nand U788 (N_788,In_946,In_763);
nor U789 (N_789,In_1406,In_1226);
nor U790 (N_790,In_857,In_335);
nand U791 (N_791,In_908,In_1104);
nor U792 (N_792,In_577,In_171);
and U793 (N_793,In_870,In_934);
or U794 (N_794,In_439,In_1180);
or U795 (N_795,In_1432,In_851);
nand U796 (N_796,In_1383,In_1223);
nor U797 (N_797,In_622,In_547);
or U798 (N_798,In_1158,In_546);
and U799 (N_799,In_768,In_1252);
or U800 (N_800,In_776,In_107);
and U801 (N_801,In_1353,In_135);
or U802 (N_802,In_1360,In_618);
and U803 (N_803,In_861,In_1009);
nand U804 (N_804,In_1483,In_49);
or U805 (N_805,In_1039,In_669);
nand U806 (N_806,In_483,In_290);
and U807 (N_807,In_365,In_1195);
or U808 (N_808,In_721,In_756);
or U809 (N_809,In_411,In_465);
nor U810 (N_810,In_966,In_221);
and U811 (N_811,In_490,In_416);
nor U812 (N_812,In_1357,In_1425);
nor U813 (N_813,In_8,In_904);
nand U814 (N_814,In_612,In_844);
nor U815 (N_815,In_690,In_995);
nand U816 (N_816,In_162,In_111);
and U817 (N_817,In_282,In_181);
nand U818 (N_818,In_1413,In_669);
and U819 (N_819,In_232,In_565);
or U820 (N_820,In_937,In_366);
or U821 (N_821,In_1023,In_197);
and U822 (N_822,In_334,In_1193);
nor U823 (N_823,In_76,In_1069);
and U824 (N_824,In_945,In_559);
nand U825 (N_825,In_360,In_964);
and U826 (N_826,In_236,In_90);
nor U827 (N_827,In_226,In_713);
nor U828 (N_828,In_137,In_1211);
and U829 (N_829,In_1117,In_1401);
and U830 (N_830,In_1140,In_626);
nand U831 (N_831,In_651,In_187);
nand U832 (N_832,In_1459,In_958);
nor U833 (N_833,In_1193,In_464);
nor U834 (N_834,In_1308,In_1432);
nand U835 (N_835,In_307,In_1316);
nor U836 (N_836,In_422,In_1476);
nor U837 (N_837,In_691,In_584);
or U838 (N_838,In_402,In_1040);
or U839 (N_839,In_646,In_483);
and U840 (N_840,In_713,In_994);
xor U841 (N_841,In_549,In_831);
and U842 (N_842,In_290,In_892);
nor U843 (N_843,In_79,In_603);
or U844 (N_844,In_297,In_118);
nor U845 (N_845,In_114,In_339);
and U846 (N_846,In_1161,In_1378);
or U847 (N_847,In_593,In_868);
nand U848 (N_848,In_541,In_310);
and U849 (N_849,In_1374,In_18);
nor U850 (N_850,In_1122,In_991);
or U851 (N_851,In_805,In_245);
and U852 (N_852,In_588,In_155);
or U853 (N_853,In_797,In_1115);
and U854 (N_854,In_1268,In_1320);
nand U855 (N_855,In_670,In_424);
nor U856 (N_856,In_499,In_265);
and U857 (N_857,In_916,In_1421);
nor U858 (N_858,In_66,In_641);
nor U859 (N_859,In_1037,In_174);
or U860 (N_860,In_758,In_216);
and U861 (N_861,In_427,In_1062);
and U862 (N_862,In_830,In_902);
nand U863 (N_863,In_725,In_717);
nand U864 (N_864,In_1191,In_1382);
nand U865 (N_865,In_835,In_988);
nand U866 (N_866,In_1055,In_329);
xor U867 (N_867,In_571,In_18);
nor U868 (N_868,In_1230,In_827);
or U869 (N_869,In_788,In_1482);
nand U870 (N_870,In_640,In_131);
nor U871 (N_871,In_586,In_330);
nor U872 (N_872,In_1490,In_314);
or U873 (N_873,In_728,In_885);
xor U874 (N_874,In_621,In_591);
and U875 (N_875,In_190,In_1313);
or U876 (N_876,In_101,In_1161);
and U877 (N_877,In_185,In_204);
and U878 (N_878,In_484,In_344);
xnor U879 (N_879,In_656,In_351);
and U880 (N_880,In_1003,In_1060);
and U881 (N_881,In_797,In_1280);
nor U882 (N_882,In_1208,In_1165);
and U883 (N_883,In_1349,In_1169);
nor U884 (N_884,In_209,In_383);
or U885 (N_885,In_802,In_239);
and U886 (N_886,In_1372,In_421);
nand U887 (N_887,In_1443,In_525);
nand U888 (N_888,In_529,In_1492);
or U889 (N_889,In_516,In_292);
xor U890 (N_890,In_451,In_5);
or U891 (N_891,In_1407,In_271);
nand U892 (N_892,In_936,In_512);
nor U893 (N_893,In_925,In_420);
and U894 (N_894,In_350,In_628);
nand U895 (N_895,In_266,In_1345);
nand U896 (N_896,In_1426,In_1391);
and U897 (N_897,In_1091,In_1080);
xor U898 (N_898,In_909,In_50);
nand U899 (N_899,In_60,In_1377);
xor U900 (N_900,In_932,In_1299);
or U901 (N_901,In_489,In_713);
nand U902 (N_902,In_376,In_648);
and U903 (N_903,In_358,In_68);
and U904 (N_904,In_442,In_503);
nor U905 (N_905,In_317,In_762);
or U906 (N_906,In_1236,In_786);
or U907 (N_907,In_678,In_942);
or U908 (N_908,In_1176,In_338);
nand U909 (N_909,In_511,In_902);
and U910 (N_910,In_1401,In_883);
nor U911 (N_911,In_434,In_1340);
and U912 (N_912,In_1434,In_488);
and U913 (N_913,In_224,In_1495);
nand U914 (N_914,In_674,In_718);
nor U915 (N_915,In_1404,In_1135);
nand U916 (N_916,In_1368,In_417);
and U917 (N_917,In_1364,In_1486);
and U918 (N_918,In_5,In_654);
or U919 (N_919,In_190,In_1259);
or U920 (N_920,In_241,In_881);
or U921 (N_921,In_1254,In_96);
or U922 (N_922,In_897,In_828);
or U923 (N_923,In_237,In_595);
or U924 (N_924,In_1076,In_213);
nand U925 (N_925,In_847,In_295);
nand U926 (N_926,In_1450,In_809);
and U927 (N_927,In_673,In_741);
xor U928 (N_928,In_1442,In_1046);
nor U929 (N_929,In_208,In_850);
or U930 (N_930,In_273,In_768);
xor U931 (N_931,In_1176,In_1428);
nor U932 (N_932,In_52,In_1439);
xor U933 (N_933,In_1096,In_1335);
nand U934 (N_934,In_1038,In_682);
nand U935 (N_935,In_1376,In_108);
or U936 (N_936,In_1056,In_366);
nand U937 (N_937,In_1105,In_1388);
and U938 (N_938,In_1481,In_1006);
nor U939 (N_939,In_1421,In_743);
or U940 (N_940,In_190,In_733);
and U941 (N_941,In_1279,In_1149);
nor U942 (N_942,In_1311,In_1135);
nor U943 (N_943,In_304,In_1279);
nand U944 (N_944,In_1085,In_458);
nor U945 (N_945,In_478,In_400);
or U946 (N_946,In_892,In_487);
nor U947 (N_947,In_1460,In_104);
and U948 (N_948,In_1238,In_826);
and U949 (N_949,In_1059,In_1262);
nand U950 (N_950,In_829,In_823);
nand U951 (N_951,In_227,In_62);
nand U952 (N_952,In_571,In_1445);
nand U953 (N_953,In_1389,In_910);
nor U954 (N_954,In_85,In_141);
nor U955 (N_955,In_434,In_9);
and U956 (N_956,In_799,In_194);
and U957 (N_957,In_723,In_1182);
or U958 (N_958,In_108,In_1496);
and U959 (N_959,In_943,In_1029);
or U960 (N_960,In_514,In_767);
or U961 (N_961,In_911,In_319);
nand U962 (N_962,In_1305,In_772);
nor U963 (N_963,In_27,In_861);
nor U964 (N_964,In_24,In_1455);
nand U965 (N_965,In_1119,In_568);
and U966 (N_966,In_737,In_987);
or U967 (N_967,In_1289,In_776);
nand U968 (N_968,In_228,In_166);
and U969 (N_969,In_441,In_244);
and U970 (N_970,In_986,In_265);
nand U971 (N_971,In_2,In_627);
nor U972 (N_972,In_1044,In_216);
and U973 (N_973,In_1491,In_938);
nand U974 (N_974,In_527,In_1075);
nand U975 (N_975,In_955,In_1261);
or U976 (N_976,In_1311,In_1375);
and U977 (N_977,In_346,In_419);
or U978 (N_978,In_977,In_267);
nand U979 (N_979,In_742,In_655);
and U980 (N_980,In_289,In_438);
or U981 (N_981,In_1365,In_153);
nand U982 (N_982,In_177,In_1301);
nor U983 (N_983,In_398,In_1063);
or U984 (N_984,In_86,In_337);
nor U985 (N_985,In_407,In_816);
nor U986 (N_986,In_800,In_1202);
and U987 (N_987,In_1259,In_44);
nand U988 (N_988,In_986,In_1018);
or U989 (N_989,In_1155,In_414);
and U990 (N_990,In_523,In_411);
or U991 (N_991,In_1209,In_576);
or U992 (N_992,In_957,In_31);
nor U993 (N_993,In_1484,In_493);
or U994 (N_994,In_991,In_1395);
nor U995 (N_995,In_1087,In_885);
or U996 (N_996,In_871,In_1220);
nand U997 (N_997,In_997,In_994);
and U998 (N_998,In_896,In_138);
nor U999 (N_999,In_1023,In_945);
nor U1000 (N_1000,In_659,In_908);
or U1001 (N_1001,In_120,In_828);
or U1002 (N_1002,In_330,In_460);
or U1003 (N_1003,In_534,In_102);
nand U1004 (N_1004,In_1105,In_416);
and U1005 (N_1005,In_682,In_376);
nand U1006 (N_1006,In_1007,In_674);
nand U1007 (N_1007,In_304,In_985);
and U1008 (N_1008,In_1492,In_258);
nor U1009 (N_1009,In_1459,In_31);
nor U1010 (N_1010,In_1480,In_682);
nand U1011 (N_1011,In_381,In_690);
nand U1012 (N_1012,In_239,In_1494);
and U1013 (N_1013,In_185,In_32);
nand U1014 (N_1014,In_1159,In_392);
nor U1015 (N_1015,In_1221,In_233);
and U1016 (N_1016,In_385,In_350);
nor U1017 (N_1017,In_785,In_528);
nor U1018 (N_1018,In_1049,In_328);
nor U1019 (N_1019,In_1372,In_759);
and U1020 (N_1020,In_1496,In_1070);
or U1021 (N_1021,In_1040,In_1200);
or U1022 (N_1022,In_1467,In_791);
nand U1023 (N_1023,In_1213,In_291);
nand U1024 (N_1024,In_948,In_1005);
nor U1025 (N_1025,In_645,In_1140);
or U1026 (N_1026,In_461,In_118);
xnor U1027 (N_1027,In_1414,In_47);
xnor U1028 (N_1028,In_1166,In_96);
or U1029 (N_1029,In_626,In_1216);
nand U1030 (N_1030,In_138,In_321);
nand U1031 (N_1031,In_5,In_467);
xor U1032 (N_1032,In_138,In_1400);
nor U1033 (N_1033,In_164,In_42);
or U1034 (N_1034,In_425,In_1431);
or U1035 (N_1035,In_359,In_945);
nand U1036 (N_1036,In_174,In_883);
and U1037 (N_1037,In_301,In_1436);
and U1038 (N_1038,In_374,In_1131);
and U1039 (N_1039,In_92,In_1435);
or U1040 (N_1040,In_759,In_1365);
nor U1041 (N_1041,In_109,In_566);
nand U1042 (N_1042,In_769,In_1291);
or U1043 (N_1043,In_150,In_1058);
or U1044 (N_1044,In_1365,In_717);
or U1045 (N_1045,In_618,In_1239);
or U1046 (N_1046,In_85,In_150);
and U1047 (N_1047,In_1372,In_1339);
nor U1048 (N_1048,In_132,In_252);
and U1049 (N_1049,In_760,In_126);
or U1050 (N_1050,In_459,In_1263);
nand U1051 (N_1051,In_469,In_1268);
nor U1052 (N_1052,In_693,In_605);
nor U1053 (N_1053,In_355,In_420);
and U1054 (N_1054,In_1085,In_733);
nor U1055 (N_1055,In_1439,In_1248);
nor U1056 (N_1056,In_652,In_557);
or U1057 (N_1057,In_572,In_199);
and U1058 (N_1058,In_1134,In_1012);
and U1059 (N_1059,In_285,In_79);
nand U1060 (N_1060,In_452,In_591);
nand U1061 (N_1061,In_1499,In_710);
and U1062 (N_1062,In_1038,In_107);
or U1063 (N_1063,In_955,In_1149);
and U1064 (N_1064,In_707,In_449);
nand U1065 (N_1065,In_367,In_510);
nand U1066 (N_1066,In_322,In_754);
or U1067 (N_1067,In_1168,In_1129);
nand U1068 (N_1068,In_807,In_1249);
nor U1069 (N_1069,In_919,In_787);
nand U1070 (N_1070,In_6,In_11);
or U1071 (N_1071,In_714,In_268);
or U1072 (N_1072,In_416,In_258);
or U1073 (N_1073,In_1190,In_1421);
or U1074 (N_1074,In_1108,In_1220);
nand U1075 (N_1075,In_379,In_555);
or U1076 (N_1076,In_425,In_547);
nor U1077 (N_1077,In_2,In_1160);
or U1078 (N_1078,In_187,In_1322);
nand U1079 (N_1079,In_1062,In_1112);
nand U1080 (N_1080,In_1339,In_436);
and U1081 (N_1081,In_417,In_972);
and U1082 (N_1082,In_354,In_1111);
and U1083 (N_1083,In_270,In_937);
or U1084 (N_1084,In_1217,In_202);
and U1085 (N_1085,In_562,In_1276);
xor U1086 (N_1086,In_15,In_1453);
or U1087 (N_1087,In_228,In_762);
and U1088 (N_1088,In_567,In_576);
nand U1089 (N_1089,In_234,In_85);
nor U1090 (N_1090,In_1236,In_1018);
and U1091 (N_1091,In_981,In_1432);
xor U1092 (N_1092,In_88,In_405);
xor U1093 (N_1093,In_1271,In_1400);
nand U1094 (N_1094,In_230,In_298);
or U1095 (N_1095,In_618,In_224);
and U1096 (N_1096,In_100,In_392);
and U1097 (N_1097,In_274,In_610);
or U1098 (N_1098,In_1365,In_511);
or U1099 (N_1099,In_1349,In_1382);
nor U1100 (N_1100,In_823,In_17);
nand U1101 (N_1101,In_1435,In_399);
nand U1102 (N_1102,In_534,In_676);
nand U1103 (N_1103,In_1251,In_469);
nor U1104 (N_1104,In_458,In_980);
nand U1105 (N_1105,In_479,In_458);
and U1106 (N_1106,In_18,In_467);
nand U1107 (N_1107,In_161,In_546);
and U1108 (N_1108,In_1081,In_1453);
nor U1109 (N_1109,In_573,In_1166);
xor U1110 (N_1110,In_501,In_450);
or U1111 (N_1111,In_1389,In_1163);
and U1112 (N_1112,In_447,In_218);
nand U1113 (N_1113,In_615,In_1317);
and U1114 (N_1114,In_6,In_545);
xor U1115 (N_1115,In_36,In_1197);
nor U1116 (N_1116,In_394,In_1407);
or U1117 (N_1117,In_274,In_1245);
nor U1118 (N_1118,In_722,In_31);
nand U1119 (N_1119,In_682,In_397);
and U1120 (N_1120,In_428,In_189);
nand U1121 (N_1121,In_852,In_939);
and U1122 (N_1122,In_353,In_1427);
nand U1123 (N_1123,In_1301,In_317);
nand U1124 (N_1124,In_1379,In_486);
and U1125 (N_1125,In_1032,In_830);
and U1126 (N_1126,In_616,In_297);
nand U1127 (N_1127,In_1207,In_721);
and U1128 (N_1128,In_844,In_1311);
nand U1129 (N_1129,In_1325,In_1123);
or U1130 (N_1130,In_493,In_549);
and U1131 (N_1131,In_1344,In_198);
or U1132 (N_1132,In_891,In_1335);
or U1133 (N_1133,In_791,In_1133);
nor U1134 (N_1134,In_223,In_83);
or U1135 (N_1135,In_802,In_1106);
nand U1136 (N_1136,In_1484,In_1422);
nand U1137 (N_1137,In_369,In_1461);
or U1138 (N_1138,In_1218,In_80);
or U1139 (N_1139,In_341,In_307);
and U1140 (N_1140,In_916,In_177);
or U1141 (N_1141,In_1460,In_532);
or U1142 (N_1142,In_1465,In_348);
nor U1143 (N_1143,In_1412,In_36);
nor U1144 (N_1144,In_1052,In_238);
or U1145 (N_1145,In_796,In_1032);
and U1146 (N_1146,In_992,In_1117);
and U1147 (N_1147,In_731,In_1472);
or U1148 (N_1148,In_1062,In_995);
nand U1149 (N_1149,In_1194,In_1424);
nor U1150 (N_1150,In_16,In_408);
nor U1151 (N_1151,In_519,In_1359);
and U1152 (N_1152,In_113,In_734);
nand U1153 (N_1153,In_221,In_428);
and U1154 (N_1154,In_1393,In_758);
nor U1155 (N_1155,In_1067,In_284);
nor U1156 (N_1156,In_1320,In_570);
nand U1157 (N_1157,In_403,In_1440);
nor U1158 (N_1158,In_448,In_939);
or U1159 (N_1159,In_62,In_1007);
nand U1160 (N_1160,In_1462,In_88);
nor U1161 (N_1161,In_841,In_863);
or U1162 (N_1162,In_256,In_1164);
nand U1163 (N_1163,In_1298,In_448);
nand U1164 (N_1164,In_1213,In_533);
or U1165 (N_1165,In_834,In_30);
nand U1166 (N_1166,In_229,In_827);
or U1167 (N_1167,In_1273,In_1387);
nor U1168 (N_1168,In_261,In_729);
and U1169 (N_1169,In_887,In_849);
nand U1170 (N_1170,In_51,In_635);
or U1171 (N_1171,In_998,In_1199);
or U1172 (N_1172,In_373,In_418);
and U1173 (N_1173,In_298,In_851);
or U1174 (N_1174,In_1487,In_1004);
and U1175 (N_1175,In_1156,In_235);
or U1176 (N_1176,In_966,In_428);
nand U1177 (N_1177,In_1334,In_1447);
or U1178 (N_1178,In_309,In_400);
nor U1179 (N_1179,In_480,In_430);
nor U1180 (N_1180,In_1120,In_1419);
and U1181 (N_1181,In_354,In_366);
or U1182 (N_1182,In_679,In_827);
or U1183 (N_1183,In_743,In_249);
nor U1184 (N_1184,In_17,In_970);
nand U1185 (N_1185,In_987,In_1334);
and U1186 (N_1186,In_1229,In_765);
nand U1187 (N_1187,In_66,In_1220);
and U1188 (N_1188,In_1465,In_1357);
or U1189 (N_1189,In_919,In_402);
nand U1190 (N_1190,In_790,In_1126);
and U1191 (N_1191,In_1343,In_137);
or U1192 (N_1192,In_625,In_580);
nand U1193 (N_1193,In_1249,In_435);
or U1194 (N_1194,In_44,In_76);
nor U1195 (N_1195,In_1258,In_531);
nand U1196 (N_1196,In_591,In_269);
nand U1197 (N_1197,In_447,In_69);
nor U1198 (N_1198,In_1491,In_176);
nand U1199 (N_1199,In_839,In_782);
or U1200 (N_1200,In_312,In_644);
nor U1201 (N_1201,In_1439,In_293);
and U1202 (N_1202,In_954,In_6);
nand U1203 (N_1203,In_1367,In_1064);
nor U1204 (N_1204,In_405,In_1361);
nor U1205 (N_1205,In_432,In_1305);
nand U1206 (N_1206,In_1274,In_819);
nor U1207 (N_1207,In_243,In_675);
nor U1208 (N_1208,In_498,In_20);
or U1209 (N_1209,In_1164,In_199);
and U1210 (N_1210,In_469,In_1055);
or U1211 (N_1211,In_291,In_260);
or U1212 (N_1212,In_383,In_329);
and U1213 (N_1213,In_1412,In_604);
nand U1214 (N_1214,In_1345,In_1250);
nor U1215 (N_1215,In_606,In_817);
and U1216 (N_1216,In_1295,In_932);
or U1217 (N_1217,In_1306,In_1167);
and U1218 (N_1218,In_197,In_243);
and U1219 (N_1219,In_1071,In_246);
nor U1220 (N_1220,In_684,In_1266);
nand U1221 (N_1221,In_783,In_1494);
and U1222 (N_1222,In_1328,In_1340);
and U1223 (N_1223,In_732,In_880);
nor U1224 (N_1224,In_625,In_29);
or U1225 (N_1225,In_1400,In_596);
nand U1226 (N_1226,In_621,In_1367);
nor U1227 (N_1227,In_1149,In_702);
or U1228 (N_1228,In_14,In_498);
xnor U1229 (N_1229,In_100,In_229);
nand U1230 (N_1230,In_865,In_197);
and U1231 (N_1231,In_644,In_1190);
nand U1232 (N_1232,In_958,In_1344);
nor U1233 (N_1233,In_404,In_546);
nor U1234 (N_1234,In_6,In_144);
nand U1235 (N_1235,In_148,In_1003);
nand U1236 (N_1236,In_1004,In_164);
and U1237 (N_1237,In_532,In_811);
or U1238 (N_1238,In_1078,In_252);
nor U1239 (N_1239,In_652,In_801);
or U1240 (N_1240,In_150,In_442);
and U1241 (N_1241,In_1405,In_1142);
nand U1242 (N_1242,In_589,In_106);
or U1243 (N_1243,In_643,In_1093);
nand U1244 (N_1244,In_754,In_1117);
nand U1245 (N_1245,In_1121,In_1044);
and U1246 (N_1246,In_1361,In_278);
and U1247 (N_1247,In_1218,In_1461);
nor U1248 (N_1248,In_1450,In_151);
and U1249 (N_1249,In_226,In_820);
nand U1250 (N_1250,In_805,In_138);
nor U1251 (N_1251,In_1258,In_1218);
nand U1252 (N_1252,In_892,In_1062);
nor U1253 (N_1253,In_579,In_197);
nor U1254 (N_1254,In_1027,In_175);
nand U1255 (N_1255,In_499,In_152);
or U1256 (N_1256,In_193,In_1477);
or U1257 (N_1257,In_989,In_13);
xor U1258 (N_1258,In_1066,In_788);
and U1259 (N_1259,In_1411,In_821);
and U1260 (N_1260,In_926,In_163);
or U1261 (N_1261,In_591,In_896);
nand U1262 (N_1262,In_1081,In_1036);
nor U1263 (N_1263,In_2,In_10);
or U1264 (N_1264,In_993,In_162);
xor U1265 (N_1265,In_1250,In_1307);
or U1266 (N_1266,In_1114,In_1154);
nand U1267 (N_1267,In_546,In_1087);
nor U1268 (N_1268,In_732,In_247);
nor U1269 (N_1269,In_103,In_1479);
or U1270 (N_1270,In_482,In_278);
nand U1271 (N_1271,In_305,In_1075);
and U1272 (N_1272,In_111,In_925);
or U1273 (N_1273,In_942,In_130);
or U1274 (N_1274,In_1215,In_1033);
and U1275 (N_1275,In_721,In_2);
nor U1276 (N_1276,In_703,In_1240);
or U1277 (N_1277,In_616,In_1046);
and U1278 (N_1278,In_1495,In_1219);
or U1279 (N_1279,In_1016,In_125);
or U1280 (N_1280,In_1298,In_761);
nand U1281 (N_1281,In_586,In_166);
nand U1282 (N_1282,In_564,In_314);
and U1283 (N_1283,In_348,In_63);
and U1284 (N_1284,In_112,In_1087);
and U1285 (N_1285,In_516,In_473);
or U1286 (N_1286,In_220,In_793);
and U1287 (N_1287,In_1322,In_907);
or U1288 (N_1288,In_440,In_808);
and U1289 (N_1289,In_773,In_974);
or U1290 (N_1290,In_395,In_973);
or U1291 (N_1291,In_322,In_1189);
xor U1292 (N_1292,In_313,In_839);
or U1293 (N_1293,In_1331,In_1049);
and U1294 (N_1294,In_930,In_489);
and U1295 (N_1295,In_765,In_278);
nor U1296 (N_1296,In_154,In_72);
nand U1297 (N_1297,In_1008,In_35);
and U1298 (N_1298,In_962,In_466);
or U1299 (N_1299,In_219,In_725);
and U1300 (N_1300,In_1301,In_631);
and U1301 (N_1301,In_150,In_701);
and U1302 (N_1302,In_302,In_580);
nor U1303 (N_1303,In_566,In_622);
nand U1304 (N_1304,In_1187,In_861);
nand U1305 (N_1305,In_839,In_1086);
xnor U1306 (N_1306,In_737,In_991);
nor U1307 (N_1307,In_1044,In_842);
nand U1308 (N_1308,In_772,In_1090);
nand U1309 (N_1309,In_105,In_752);
and U1310 (N_1310,In_788,In_1088);
nand U1311 (N_1311,In_1379,In_1153);
or U1312 (N_1312,In_553,In_1062);
and U1313 (N_1313,In_1210,In_349);
or U1314 (N_1314,In_579,In_1109);
and U1315 (N_1315,In_351,In_203);
and U1316 (N_1316,In_522,In_589);
nor U1317 (N_1317,In_1252,In_988);
and U1318 (N_1318,In_1247,In_862);
and U1319 (N_1319,In_959,In_1163);
and U1320 (N_1320,In_1300,In_1397);
or U1321 (N_1321,In_396,In_703);
nor U1322 (N_1322,In_1476,In_1258);
nand U1323 (N_1323,In_1411,In_673);
nor U1324 (N_1324,In_1311,In_207);
or U1325 (N_1325,In_1376,In_1102);
nor U1326 (N_1326,In_1055,In_1484);
or U1327 (N_1327,In_943,In_1040);
and U1328 (N_1328,In_598,In_1415);
nor U1329 (N_1329,In_951,In_1207);
and U1330 (N_1330,In_257,In_1345);
nand U1331 (N_1331,In_881,In_1470);
or U1332 (N_1332,In_1057,In_409);
or U1333 (N_1333,In_18,In_960);
or U1334 (N_1334,In_974,In_853);
and U1335 (N_1335,In_454,In_1436);
nand U1336 (N_1336,In_1351,In_201);
and U1337 (N_1337,In_72,In_1410);
nor U1338 (N_1338,In_457,In_1016);
or U1339 (N_1339,In_931,In_1152);
xnor U1340 (N_1340,In_59,In_1232);
nor U1341 (N_1341,In_335,In_48);
nand U1342 (N_1342,In_272,In_759);
and U1343 (N_1343,In_1349,In_1376);
nor U1344 (N_1344,In_1077,In_17);
nand U1345 (N_1345,In_889,In_1234);
nand U1346 (N_1346,In_1227,In_613);
nand U1347 (N_1347,In_388,In_618);
and U1348 (N_1348,In_1409,In_1041);
or U1349 (N_1349,In_190,In_918);
or U1350 (N_1350,In_797,In_460);
nand U1351 (N_1351,In_507,In_451);
xnor U1352 (N_1352,In_927,In_327);
nand U1353 (N_1353,In_1444,In_1453);
and U1354 (N_1354,In_553,In_1232);
nand U1355 (N_1355,In_927,In_401);
or U1356 (N_1356,In_1436,In_445);
or U1357 (N_1357,In_162,In_786);
and U1358 (N_1358,In_415,In_71);
nand U1359 (N_1359,In_419,In_1452);
and U1360 (N_1360,In_486,In_1283);
nor U1361 (N_1361,In_278,In_185);
nand U1362 (N_1362,In_1467,In_610);
nand U1363 (N_1363,In_649,In_1461);
and U1364 (N_1364,In_827,In_238);
nand U1365 (N_1365,In_900,In_965);
nand U1366 (N_1366,In_903,In_407);
or U1367 (N_1367,In_493,In_989);
nand U1368 (N_1368,In_473,In_288);
nand U1369 (N_1369,In_1482,In_1125);
or U1370 (N_1370,In_49,In_1252);
or U1371 (N_1371,In_932,In_751);
nand U1372 (N_1372,In_837,In_389);
and U1373 (N_1373,In_942,In_116);
and U1374 (N_1374,In_960,In_673);
and U1375 (N_1375,In_1490,In_641);
or U1376 (N_1376,In_442,In_224);
and U1377 (N_1377,In_1423,In_173);
and U1378 (N_1378,In_1314,In_129);
nor U1379 (N_1379,In_1358,In_155);
nor U1380 (N_1380,In_834,In_1087);
nor U1381 (N_1381,In_94,In_634);
and U1382 (N_1382,In_175,In_970);
or U1383 (N_1383,In_17,In_683);
nor U1384 (N_1384,In_115,In_1265);
and U1385 (N_1385,In_1239,In_20);
nand U1386 (N_1386,In_827,In_1331);
or U1387 (N_1387,In_1095,In_950);
nand U1388 (N_1388,In_230,In_955);
nor U1389 (N_1389,In_495,In_294);
and U1390 (N_1390,In_520,In_477);
or U1391 (N_1391,In_518,In_1496);
nand U1392 (N_1392,In_750,In_361);
or U1393 (N_1393,In_464,In_1427);
and U1394 (N_1394,In_181,In_1249);
nor U1395 (N_1395,In_1036,In_1104);
xnor U1396 (N_1396,In_885,In_1157);
nand U1397 (N_1397,In_499,In_868);
or U1398 (N_1398,In_89,In_62);
and U1399 (N_1399,In_229,In_829);
or U1400 (N_1400,In_1451,In_606);
nor U1401 (N_1401,In_1078,In_1463);
nand U1402 (N_1402,In_1043,In_909);
nor U1403 (N_1403,In_1494,In_78);
and U1404 (N_1404,In_783,In_964);
nand U1405 (N_1405,In_449,In_75);
or U1406 (N_1406,In_185,In_578);
nand U1407 (N_1407,In_199,In_721);
or U1408 (N_1408,In_1261,In_741);
nor U1409 (N_1409,In_588,In_318);
nor U1410 (N_1410,In_169,In_804);
and U1411 (N_1411,In_1044,In_999);
or U1412 (N_1412,In_1178,In_971);
or U1413 (N_1413,In_158,In_1036);
nand U1414 (N_1414,In_158,In_1164);
nor U1415 (N_1415,In_511,In_892);
or U1416 (N_1416,In_727,In_712);
and U1417 (N_1417,In_1102,In_526);
and U1418 (N_1418,In_394,In_328);
nor U1419 (N_1419,In_899,In_251);
nor U1420 (N_1420,In_1122,In_649);
nor U1421 (N_1421,In_92,In_401);
or U1422 (N_1422,In_277,In_680);
or U1423 (N_1423,In_979,In_492);
or U1424 (N_1424,In_515,In_1456);
nand U1425 (N_1425,In_471,In_74);
nor U1426 (N_1426,In_101,In_1242);
nor U1427 (N_1427,In_1268,In_1322);
nor U1428 (N_1428,In_1117,In_1349);
nand U1429 (N_1429,In_161,In_1016);
nand U1430 (N_1430,In_917,In_56);
nor U1431 (N_1431,In_344,In_1008);
nand U1432 (N_1432,In_1255,In_1494);
and U1433 (N_1433,In_1352,In_1285);
and U1434 (N_1434,In_588,In_786);
nand U1435 (N_1435,In_581,In_766);
and U1436 (N_1436,In_630,In_182);
nor U1437 (N_1437,In_174,In_902);
nand U1438 (N_1438,In_1090,In_847);
nand U1439 (N_1439,In_111,In_285);
nand U1440 (N_1440,In_273,In_808);
or U1441 (N_1441,In_1148,In_880);
nor U1442 (N_1442,In_295,In_1001);
and U1443 (N_1443,In_598,In_1474);
or U1444 (N_1444,In_1238,In_79);
nand U1445 (N_1445,In_804,In_172);
and U1446 (N_1446,In_41,In_1235);
and U1447 (N_1447,In_1346,In_1368);
or U1448 (N_1448,In_40,In_551);
and U1449 (N_1449,In_959,In_1352);
nand U1450 (N_1450,In_1114,In_105);
nor U1451 (N_1451,In_389,In_1123);
nand U1452 (N_1452,In_854,In_331);
or U1453 (N_1453,In_602,In_1301);
nand U1454 (N_1454,In_1223,In_1100);
nor U1455 (N_1455,In_71,In_863);
and U1456 (N_1456,In_841,In_984);
or U1457 (N_1457,In_560,In_738);
xnor U1458 (N_1458,In_165,In_302);
nand U1459 (N_1459,In_401,In_1258);
or U1460 (N_1460,In_468,In_712);
or U1461 (N_1461,In_699,In_142);
or U1462 (N_1462,In_1180,In_1411);
nor U1463 (N_1463,In_485,In_468);
nand U1464 (N_1464,In_1172,In_1117);
nand U1465 (N_1465,In_1192,In_63);
nor U1466 (N_1466,In_359,In_874);
and U1467 (N_1467,In_88,In_104);
or U1468 (N_1468,In_203,In_553);
nor U1469 (N_1469,In_691,In_292);
or U1470 (N_1470,In_1465,In_1290);
nor U1471 (N_1471,In_202,In_481);
nor U1472 (N_1472,In_201,In_613);
and U1473 (N_1473,In_697,In_208);
and U1474 (N_1474,In_1330,In_57);
or U1475 (N_1475,In_783,In_1137);
nor U1476 (N_1476,In_406,In_221);
or U1477 (N_1477,In_1212,In_1141);
nor U1478 (N_1478,In_709,In_1331);
or U1479 (N_1479,In_1488,In_941);
xor U1480 (N_1480,In_416,In_1024);
nand U1481 (N_1481,In_1031,In_1058);
nand U1482 (N_1482,In_442,In_549);
and U1483 (N_1483,In_315,In_1460);
and U1484 (N_1484,In_512,In_924);
and U1485 (N_1485,In_288,In_527);
nand U1486 (N_1486,In_1291,In_1431);
or U1487 (N_1487,In_1216,In_1460);
and U1488 (N_1488,In_361,In_588);
or U1489 (N_1489,In_593,In_1420);
or U1490 (N_1490,In_596,In_1186);
and U1491 (N_1491,In_1326,In_288);
and U1492 (N_1492,In_876,In_131);
nor U1493 (N_1493,In_627,In_74);
nand U1494 (N_1494,In_544,In_956);
nor U1495 (N_1495,In_487,In_39);
nand U1496 (N_1496,In_800,In_1140);
or U1497 (N_1497,In_1105,In_1232);
xor U1498 (N_1498,In_408,In_545);
nor U1499 (N_1499,In_1046,In_1236);
or U1500 (N_1500,In_1,In_606);
or U1501 (N_1501,In_336,In_886);
and U1502 (N_1502,In_957,In_1084);
or U1503 (N_1503,In_970,In_531);
nor U1504 (N_1504,In_1004,In_868);
nor U1505 (N_1505,In_980,In_21);
nand U1506 (N_1506,In_355,In_874);
and U1507 (N_1507,In_1020,In_756);
or U1508 (N_1508,In_481,In_217);
xor U1509 (N_1509,In_375,In_1155);
and U1510 (N_1510,In_1176,In_478);
or U1511 (N_1511,In_187,In_598);
nor U1512 (N_1512,In_872,In_598);
or U1513 (N_1513,In_799,In_523);
and U1514 (N_1514,In_27,In_521);
and U1515 (N_1515,In_577,In_93);
nand U1516 (N_1516,In_169,In_952);
nand U1517 (N_1517,In_1380,In_1353);
and U1518 (N_1518,In_281,In_527);
nand U1519 (N_1519,In_1136,In_1450);
xor U1520 (N_1520,In_314,In_844);
nor U1521 (N_1521,In_1454,In_621);
or U1522 (N_1522,In_50,In_16);
nand U1523 (N_1523,In_1050,In_218);
or U1524 (N_1524,In_406,In_52);
or U1525 (N_1525,In_806,In_668);
nand U1526 (N_1526,In_1029,In_1437);
nand U1527 (N_1527,In_1288,In_1403);
nand U1528 (N_1528,In_557,In_302);
nor U1529 (N_1529,In_1147,In_905);
nor U1530 (N_1530,In_933,In_535);
nand U1531 (N_1531,In_414,In_738);
and U1532 (N_1532,In_1027,In_1351);
nand U1533 (N_1533,In_979,In_762);
or U1534 (N_1534,In_801,In_197);
and U1535 (N_1535,In_651,In_917);
nor U1536 (N_1536,In_671,In_33);
or U1537 (N_1537,In_358,In_1387);
nand U1538 (N_1538,In_1365,In_1263);
and U1539 (N_1539,In_567,In_464);
nand U1540 (N_1540,In_1100,In_410);
nor U1541 (N_1541,In_426,In_222);
or U1542 (N_1542,In_616,In_331);
xor U1543 (N_1543,In_111,In_290);
nand U1544 (N_1544,In_856,In_827);
and U1545 (N_1545,In_601,In_866);
nor U1546 (N_1546,In_760,In_1057);
nand U1547 (N_1547,In_693,In_788);
and U1548 (N_1548,In_1337,In_858);
nand U1549 (N_1549,In_1355,In_830);
nand U1550 (N_1550,In_851,In_238);
or U1551 (N_1551,In_191,In_200);
and U1552 (N_1552,In_777,In_956);
or U1553 (N_1553,In_1162,In_1368);
nor U1554 (N_1554,In_293,In_532);
and U1555 (N_1555,In_1472,In_204);
and U1556 (N_1556,In_595,In_20);
and U1557 (N_1557,In_564,In_1401);
nor U1558 (N_1558,In_1386,In_1345);
or U1559 (N_1559,In_1339,In_1491);
or U1560 (N_1560,In_1056,In_939);
nand U1561 (N_1561,In_658,In_197);
nor U1562 (N_1562,In_1054,In_838);
and U1563 (N_1563,In_819,In_768);
and U1564 (N_1564,In_907,In_155);
nand U1565 (N_1565,In_1411,In_179);
and U1566 (N_1566,In_567,In_179);
nor U1567 (N_1567,In_1321,In_434);
or U1568 (N_1568,In_379,In_561);
nor U1569 (N_1569,In_1102,In_1392);
nor U1570 (N_1570,In_1129,In_64);
nor U1571 (N_1571,In_594,In_1141);
nand U1572 (N_1572,In_463,In_1087);
nor U1573 (N_1573,In_243,In_12);
nand U1574 (N_1574,In_703,In_968);
nor U1575 (N_1575,In_1063,In_703);
nand U1576 (N_1576,In_233,In_872);
nand U1577 (N_1577,In_1310,In_1452);
nand U1578 (N_1578,In_297,In_964);
and U1579 (N_1579,In_235,In_215);
nand U1580 (N_1580,In_899,In_1344);
and U1581 (N_1581,In_253,In_396);
and U1582 (N_1582,In_64,In_791);
nor U1583 (N_1583,In_1142,In_1182);
nand U1584 (N_1584,In_605,In_1334);
and U1585 (N_1585,In_1439,In_1344);
and U1586 (N_1586,In_739,In_1369);
xnor U1587 (N_1587,In_726,In_1141);
or U1588 (N_1588,In_1404,In_862);
nand U1589 (N_1589,In_1133,In_70);
or U1590 (N_1590,In_671,In_904);
nand U1591 (N_1591,In_472,In_969);
nor U1592 (N_1592,In_458,In_1178);
nor U1593 (N_1593,In_626,In_460);
and U1594 (N_1594,In_1193,In_1472);
or U1595 (N_1595,In_320,In_1442);
and U1596 (N_1596,In_1316,In_401);
or U1597 (N_1597,In_1138,In_1272);
nor U1598 (N_1598,In_519,In_1346);
and U1599 (N_1599,In_771,In_810);
and U1600 (N_1600,In_799,In_1073);
xor U1601 (N_1601,In_141,In_545);
nor U1602 (N_1602,In_736,In_451);
or U1603 (N_1603,In_409,In_505);
or U1604 (N_1604,In_1254,In_1333);
or U1605 (N_1605,In_46,In_70);
and U1606 (N_1606,In_320,In_934);
or U1607 (N_1607,In_853,In_615);
nor U1608 (N_1608,In_897,In_10);
nand U1609 (N_1609,In_607,In_818);
and U1610 (N_1610,In_555,In_531);
or U1611 (N_1611,In_1454,In_904);
nor U1612 (N_1612,In_793,In_296);
nor U1613 (N_1613,In_1010,In_971);
nor U1614 (N_1614,In_672,In_12);
nand U1615 (N_1615,In_945,In_914);
and U1616 (N_1616,In_586,In_66);
nor U1617 (N_1617,In_426,In_1144);
nor U1618 (N_1618,In_1172,In_192);
nor U1619 (N_1619,In_630,In_914);
or U1620 (N_1620,In_546,In_1286);
and U1621 (N_1621,In_1380,In_1068);
nor U1622 (N_1622,In_777,In_917);
and U1623 (N_1623,In_368,In_1042);
nor U1624 (N_1624,In_596,In_211);
nor U1625 (N_1625,In_1272,In_1253);
nand U1626 (N_1626,In_230,In_810);
nand U1627 (N_1627,In_409,In_395);
nand U1628 (N_1628,In_827,In_316);
or U1629 (N_1629,In_1084,In_1433);
or U1630 (N_1630,In_931,In_1131);
or U1631 (N_1631,In_363,In_93);
or U1632 (N_1632,In_434,In_1269);
and U1633 (N_1633,In_328,In_714);
nand U1634 (N_1634,In_64,In_626);
nand U1635 (N_1635,In_295,In_772);
or U1636 (N_1636,In_1175,In_802);
nor U1637 (N_1637,In_361,In_941);
nand U1638 (N_1638,In_377,In_393);
or U1639 (N_1639,In_773,In_424);
nand U1640 (N_1640,In_1178,In_1114);
or U1641 (N_1641,In_11,In_1276);
nand U1642 (N_1642,In_1067,In_685);
or U1643 (N_1643,In_601,In_584);
nor U1644 (N_1644,In_740,In_1356);
nor U1645 (N_1645,In_1210,In_1347);
and U1646 (N_1646,In_1259,In_735);
nand U1647 (N_1647,In_982,In_1406);
and U1648 (N_1648,In_1359,In_175);
or U1649 (N_1649,In_363,In_868);
nor U1650 (N_1650,In_28,In_1131);
and U1651 (N_1651,In_1240,In_63);
or U1652 (N_1652,In_869,In_374);
nand U1653 (N_1653,In_788,In_296);
nor U1654 (N_1654,In_47,In_1195);
and U1655 (N_1655,In_174,In_776);
nand U1656 (N_1656,In_678,In_667);
xor U1657 (N_1657,In_1200,In_964);
or U1658 (N_1658,In_1053,In_345);
and U1659 (N_1659,In_568,In_553);
nor U1660 (N_1660,In_791,In_342);
nand U1661 (N_1661,In_628,In_428);
nand U1662 (N_1662,In_1427,In_254);
nor U1663 (N_1663,In_1274,In_1466);
nand U1664 (N_1664,In_1484,In_1161);
nor U1665 (N_1665,In_1233,In_900);
and U1666 (N_1666,In_1395,In_56);
xor U1667 (N_1667,In_1488,In_561);
nand U1668 (N_1668,In_878,In_1137);
and U1669 (N_1669,In_418,In_1061);
nor U1670 (N_1670,In_543,In_1380);
or U1671 (N_1671,In_1036,In_1206);
or U1672 (N_1672,In_127,In_96);
nor U1673 (N_1673,In_164,In_377);
or U1674 (N_1674,In_87,In_738);
and U1675 (N_1675,In_1211,In_176);
nor U1676 (N_1676,In_1080,In_593);
nand U1677 (N_1677,In_694,In_715);
or U1678 (N_1678,In_578,In_1210);
nand U1679 (N_1679,In_1305,In_991);
nor U1680 (N_1680,In_828,In_1273);
or U1681 (N_1681,In_281,In_1314);
nor U1682 (N_1682,In_922,In_712);
nor U1683 (N_1683,In_928,In_94);
nor U1684 (N_1684,In_664,In_599);
nand U1685 (N_1685,In_1002,In_1254);
xnor U1686 (N_1686,In_1096,In_369);
nor U1687 (N_1687,In_82,In_393);
and U1688 (N_1688,In_1255,In_573);
and U1689 (N_1689,In_1310,In_850);
nor U1690 (N_1690,In_638,In_861);
nand U1691 (N_1691,In_1080,In_881);
and U1692 (N_1692,In_1238,In_52);
or U1693 (N_1693,In_1224,In_236);
or U1694 (N_1694,In_1474,In_851);
nor U1695 (N_1695,In_548,In_1309);
and U1696 (N_1696,In_229,In_1077);
and U1697 (N_1697,In_1093,In_1393);
and U1698 (N_1698,In_483,In_1371);
or U1699 (N_1699,In_1350,In_515);
or U1700 (N_1700,In_1297,In_755);
nand U1701 (N_1701,In_792,In_764);
and U1702 (N_1702,In_1229,In_815);
nor U1703 (N_1703,In_465,In_12);
nand U1704 (N_1704,In_182,In_94);
nor U1705 (N_1705,In_369,In_1033);
or U1706 (N_1706,In_1002,In_735);
nor U1707 (N_1707,In_322,In_805);
or U1708 (N_1708,In_1250,In_757);
nor U1709 (N_1709,In_763,In_511);
or U1710 (N_1710,In_855,In_1452);
nor U1711 (N_1711,In_423,In_1284);
or U1712 (N_1712,In_362,In_187);
or U1713 (N_1713,In_1353,In_1028);
nand U1714 (N_1714,In_423,In_1069);
or U1715 (N_1715,In_245,In_1276);
nand U1716 (N_1716,In_482,In_103);
nand U1717 (N_1717,In_396,In_912);
nor U1718 (N_1718,In_712,In_602);
nand U1719 (N_1719,In_1296,In_58);
or U1720 (N_1720,In_211,In_814);
nand U1721 (N_1721,In_94,In_880);
or U1722 (N_1722,In_707,In_1324);
nor U1723 (N_1723,In_939,In_1270);
nand U1724 (N_1724,In_386,In_837);
and U1725 (N_1725,In_731,In_640);
or U1726 (N_1726,In_964,In_867);
nor U1727 (N_1727,In_965,In_69);
and U1728 (N_1728,In_1249,In_1264);
nand U1729 (N_1729,In_938,In_870);
or U1730 (N_1730,In_944,In_176);
nor U1731 (N_1731,In_628,In_688);
nand U1732 (N_1732,In_529,In_481);
xor U1733 (N_1733,In_393,In_467);
nand U1734 (N_1734,In_421,In_1414);
nand U1735 (N_1735,In_1389,In_1397);
and U1736 (N_1736,In_1200,In_1133);
nor U1737 (N_1737,In_29,In_647);
nor U1738 (N_1738,In_1109,In_151);
and U1739 (N_1739,In_865,In_679);
or U1740 (N_1740,In_1377,In_1437);
and U1741 (N_1741,In_722,In_343);
or U1742 (N_1742,In_1047,In_1064);
nand U1743 (N_1743,In_670,In_930);
nand U1744 (N_1744,In_626,In_637);
or U1745 (N_1745,In_1390,In_267);
and U1746 (N_1746,In_1155,In_755);
and U1747 (N_1747,In_996,In_459);
and U1748 (N_1748,In_794,In_837);
nor U1749 (N_1749,In_682,In_621);
nand U1750 (N_1750,In_545,In_1044);
or U1751 (N_1751,In_809,In_1129);
and U1752 (N_1752,In_750,In_893);
nor U1753 (N_1753,In_1378,In_1060);
nand U1754 (N_1754,In_214,In_850);
nor U1755 (N_1755,In_1486,In_1122);
or U1756 (N_1756,In_1104,In_540);
and U1757 (N_1757,In_1026,In_165);
nand U1758 (N_1758,In_1006,In_530);
nor U1759 (N_1759,In_860,In_906);
nand U1760 (N_1760,In_1229,In_676);
or U1761 (N_1761,In_122,In_37);
nand U1762 (N_1762,In_168,In_506);
or U1763 (N_1763,In_1466,In_314);
nand U1764 (N_1764,In_989,In_1187);
or U1765 (N_1765,In_1178,In_153);
nor U1766 (N_1766,In_606,In_244);
nand U1767 (N_1767,In_855,In_849);
nand U1768 (N_1768,In_1172,In_471);
nor U1769 (N_1769,In_1079,In_381);
nor U1770 (N_1770,In_779,In_1016);
and U1771 (N_1771,In_619,In_877);
or U1772 (N_1772,In_314,In_1236);
nor U1773 (N_1773,In_939,In_908);
or U1774 (N_1774,In_639,In_58);
nor U1775 (N_1775,In_313,In_1003);
nor U1776 (N_1776,In_1419,In_1144);
nor U1777 (N_1777,In_1080,In_112);
nand U1778 (N_1778,In_325,In_826);
nor U1779 (N_1779,In_1316,In_1425);
nand U1780 (N_1780,In_851,In_414);
xor U1781 (N_1781,In_1063,In_696);
nor U1782 (N_1782,In_220,In_111);
nand U1783 (N_1783,In_1171,In_143);
nor U1784 (N_1784,In_1485,In_852);
nand U1785 (N_1785,In_1054,In_47);
or U1786 (N_1786,In_153,In_467);
xnor U1787 (N_1787,In_1113,In_862);
and U1788 (N_1788,In_1371,In_1386);
nor U1789 (N_1789,In_1070,In_885);
xor U1790 (N_1790,In_356,In_1030);
nand U1791 (N_1791,In_137,In_685);
nor U1792 (N_1792,In_1155,In_197);
or U1793 (N_1793,In_906,In_920);
nor U1794 (N_1794,In_485,In_1260);
and U1795 (N_1795,In_562,In_1101);
nand U1796 (N_1796,In_718,In_1276);
and U1797 (N_1797,In_968,In_1111);
and U1798 (N_1798,In_140,In_656);
nor U1799 (N_1799,In_659,In_1487);
nor U1800 (N_1800,In_1468,In_698);
nand U1801 (N_1801,In_17,In_159);
nand U1802 (N_1802,In_954,In_709);
nor U1803 (N_1803,In_1204,In_726);
nand U1804 (N_1804,In_1289,In_586);
nand U1805 (N_1805,In_1231,In_739);
nor U1806 (N_1806,In_939,In_1376);
nand U1807 (N_1807,In_113,In_356);
nor U1808 (N_1808,In_81,In_30);
and U1809 (N_1809,In_1003,In_822);
nor U1810 (N_1810,In_738,In_1472);
or U1811 (N_1811,In_567,In_490);
nor U1812 (N_1812,In_195,In_1284);
nand U1813 (N_1813,In_412,In_708);
nand U1814 (N_1814,In_659,In_1068);
or U1815 (N_1815,In_1062,In_507);
and U1816 (N_1816,In_389,In_758);
nor U1817 (N_1817,In_1481,In_1247);
and U1818 (N_1818,In_61,In_344);
and U1819 (N_1819,In_472,In_203);
and U1820 (N_1820,In_825,In_807);
nor U1821 (N_1821,In_985,In_842);
and U1822 (N_1822,In_796,In_535);
or U1823 (N_1823,In_333,In_1488);
or U1824 (N_1824,In_190,In_1303);
nor U1825 (N_1825,In_460,In_1439);
and U1826 (N_1826,In_1087,In_147);
and U1827 (N_1827,In_1095,In_503);
nor U1828 (N_1828,In_1236,In_1275);
or U1829 (N_1829,In_451,In_79);
nor U1830 (N_1830,In_1169,In_845);
or U1831 (N_1831,In_538,In_44);
and U1832 (N_1832,In_738,In_583);
nor U1833 (N_1833,In_84,In_628);
nor U1834 (N_1834,In_1109,In_752);
nor U1835 (N_1835,In_1103,In_1212);
or U1836 (N_1836,In_383,In_668);
and U1837 (N_1837,In_1114,In_1462);
or U1838 (N_1838,In_419,In_1201);
and U1839 (N_1839,In_723,In_618);
nand U1840 (N_1840,In_648,In_1030);
nand U1841 (N_1841,In_1338,In_608);
nand U1842 (N_1842,In_619,In_581);
and U1843 (N_1843,In_711,In_308);
nor U1844 (N_1844,In_951,In_778);
nand U1845 (N_1845,In_1480,In_771);
and U1846 (N_1846,In_1410,In_1183);
nand U1847 (N_1847,In_886,In_580);
nand U1848 (N_1848,In_181,In_1325);
and U1849 (N_1849,In_870,In_851);
or U1850 (N_1850,In_571,In_1281);
and U1851 (N_1851,In_1360,In_253);
or U1852 (N_1852,In_381,In_1256);
and U1853 (N_1853,In_250,In_780);
or U1854 (N_1854,In_1107,In_1472);
and U1855 (N_1855,In_1432,In_459);
or U1856 (N_1856,In_1150,In_1466);
or U1857 (N_1857,In_44,In_872);
nor U1858 (N_1858,In_40,In_685);
nor U1859 (N_1859,In_616,In_334);
nand U1860 (N_1860,In_1497,In_939);
and U1861 (N_1861,In_1056,In_812);
or U1862 (N_1862,In_1362,In_123);
or U1863 (N_1863,In_31,In_1011);
or U1864 (N_1864,In_541,In_1027);
or U1865 (N_1865,In_442,In_748);
or U1866 (N_1866,In_190,In_1290);
nand U1867 (N_1867,In_105,In_1499);
or U1868 (N_1868,In_374,In_341);
nor U1869 (N_1869,In_1406,In_599);
nand U1870 (N_1870,In_831,In_78);
nor U1871 (N_1871,In_634,In_156);
or U1872 (N_1872,In_1163,In_1056);
or U1873 (N_1873,In_440,In_788);
and U1874 (N_1874,In_427,In_726);
nand U1875 (N_1875,In_235,In_483);
nand U1876 (N_1876,In_1167,In_1453);
and U1877 (N_1877,In_333,In_886);
nor U1878 (N_1878,In_1367,In_665);
nand U1879 (N_1879,In_930,In_1406);
nand U1880 (N_1880,In_1343,In_2);
nor U1881 (N_1881,In_745,In_451);
nand U1882 (N_1882,In_1384,In_964);
and U1883 (N_1883,In_769,In_30);
nand U1884 (N_1884,In_1063,In_1304);
nand U1885 (N_1885,In_1169,In_289);
or U1886 (N_1886,In_763,In_620);
nand U1887 (N_1887,In_572,In_70);
nor U1888 (N_1888,In_404,In_1498);
nor U1889 (N_1889,In_1305,In_1405);
and U1890 (N_1890,In_345,In_1064);
and U1891 (N_1891,In_646,In_1327);
nor U1892 (N_1892,In_906,In_1271);
and U1893 (N_1893,In_1387,In_1137);
and U1894 (N_1894,In_1466,In_986);
and U1895 (N_1895,In_1446,In_972);
nand U1896 (N_1896,In_319,In_1482);
nand U1897 (N_1897,In_214,In_273);
or U1898 (N_1898,In_524,In_1187);
nor U1899 (N_1899,In_309,In_384);
nor U1900 (N_1900,In_1011,In_591);
or U1901 (N_1901,In_338,In_552);
and U1902 (N_1902,In_879,In_30);
xnor U1903 (N_1903,In_1286,In_584);
and U1904 (N_1904,In_633,In_1156);
or U1905 (N_1905,In_1279,In_324);
nand U1906 (N_1906,In_1448,In_1115);
nor U1907 (N_1907,In_825,In_1195);
nand U1908 (N_1908,In_171,In_127);
and U1909 (N_1909,In_809,In_587);
nor U1910 (N_1910,In_1417,In_1362);
nor U1911 (N_1911,In_1237,In_232);
and U1912 (N_1912,In_334,In_517);
or U1913 (N_1913,In_426,In_692);
or U1914 (N_1914,In_714,In_506);
or U1915 (N_1915,In_244,In_895);
and U1916 (N_1916,In_1186,In_974);
and U1917 (N_1917,In_804,In_500);
and U1918 (N_1918,In_89,In_1153);
nand U1919 (N_1919,In_435,In_75);
or U1920 (N_1920,In_1037,In_0);
or U1921 (N_1921,In_287,In_1296);
or U1922 (N_1922,In_658,In_313);
and U1923 (N_1923,In_1062,In_699);
nand U1924 (N_1924,In_774,In_1133);
and U1925 (N_1925,In_616,In_409);
or U1926 (N_1926,In_1355,In_1446);
xnor U1927 (N_1927,In_1229,In_710);
or U1928 (N_1928,In_247,In_132);
nand U1929 (N_1929,In_511,In_750);
and U1930 (N_1930,In_437,In_378);
nand U1931 (N_1931,In_411,In_412);
nand U1932 (N_1932,In_1203,In_1279);
nand U1933 (N_1933,In_1278,In_382);
nand U1934 (N_1934,In_688,In_88);
or U1935 (N_1935,In_129,In_1156);
or U1936 (N_1936,In_185,In_591);
nor U1937 (N_1937,In_984,In_968);
nand U1938 (N_1938,In_1053,In_1499);
nand U1939 (N_1939,In_1416,In_1335);
nand U1940 (N_1940,In_709,In_1095);
and U1941 (N_1941,In_1199,In_852);
and U1942 (N_1942,In_239,In_854);
and U1943 (N_1943,In_426,In_1319);
nor U1944 (N_1944,In_843,In_673);
nand U1945 (N_1945,In_740,In_1337);
or U1946 (N_1946,In_641,In_1283);
and U1947 (N_1947,In_891,In_1309);
and U1948 (N_1948,In_480,In_203);
nand U1949 (N_1949,In_246,In_976);
or U1950 (N_1950,In_1454,In_746);
or U1951 (N_1951,In_247,In_351);
and U1952 (N_1952,In_375,In_402);
or U1953 (N_1953,In_690,In_1419);
or U1954 (N_1954,In_315,In_625);
nor U1955 (N_1955,In_1485,In_578);
nand U1956 (N_1956,In_1294,In_1078);
and U1957 (N_1957,In_537,In_585);
nor U1958 (N_1958,In_1204,In_542);
or U1959 (N_1959,In_1120,In_469);
and U1960 (N_1960,In_1390,In_1268);
and U1961 (N_1961,In_635,In_1282);
nand U1962 (N_1962,In_361,In_1122);
or U1963 (N_1963,In_1308,In_564);
or U1964 (N_1964,In_1413,In_345);
nand U1965 (N_1965,In_984,In_34);
and U1966 (N_1966,In_1111,In_430);
nor U1967 (N_1967,In_569,In_676);
nand U1968 (N_1968,In_998,In_328);
nand U1969 (N_1969,In_1208,In_8);
nand U1970 (N_1970,In_478,In_865);
and U1971 (N_1971,In_1090,In_673);
nand U1972 (N_1972,In_1080,In_906);
nand U1973 (N_1973,In_304,In_13);
nand U1974 (N_1974,In_252,In_1314);
or U1975 (N_1975,In_371,In_1347);
nand U1976 (N_1976,In_1273,In_1109);
and U1977 (N_1977,In_630,In_725);
nor U1978 (N_1978,In_1068,In_42);
nand U1979 (N_1979,In_423,In_1202);
nand U1980 (N_1980,In_818,In_943);
xor U1981 (N_1981,In_903,In_792);
nand U1982 (N_1982,In_1162,In_1057);
nand U1983 (N_1983,In_1098,In_1227);
and U1984 (N_1984,In_771,In_385);
or U1985 (N_1985,In_820,In_522);
nor U1986 (N_1986,In_1088,In_1114);
or U1987 (N_1987,In_681,In_479);
and U1988 (N_1988,In_558,In_1419);
nand U1989 (N_1989,In_263,In_374);
xor U1990 (N_1990,In_1458,In_1360);
and U1991 (N_1991,In_42,In_60);
nand U1992 (N_1992,In_736,In_473);
nand U1993 (N_1993,In_324,In_1468);
and U1994 (N_1994,In_438,In_1480);
nand U1995 (N_1995,In_1184,In_979);
nand U1996 (N_1996,In_349,In_10);
or U1997 (N_1997,In_1381,In_1070);
nand U1998 (N_1998,In_1227,In_721);
nand U1999 (N_1999,In_763,In_1165);
and U2000 (N_2000,In_453,In_157);
and U2001 (N_2001,In_1437,In_112);
nand U2002 (N_2002,In_865,In_876);
or U2003 (N_2003,In_569,In_1451);
and U2004 (N_2004,In_882,In_1247);
nor U2005 (N_2005,In_57,In_1377);
and U2006 (N_2006,In_634,In_597);
nand U2007 (N_2007,In_322,In_508);
or U2008 (N_2008,In_395,In_183);
nor U2009 (N_2009,In_1287,In_385);
nand U2010 (N_2010,In_605,In_547);
nor U2011 (N_2011,In_1122,In_1008);
and U2012 (N_2012,In_280,In_313);
xnor U2013 (N_2013,In_1254,In_231);
or U2014 (N_2014,In_525,In_1215);
nand U2015 (N_2015,In_1109,In_949);
nand U2016 (N_2016,In_840,In_1038);
and U2017 (N_2017,In_458,In_538);
and U2018 (N_2018,In_281,In_9);
xor U2019 (N_2019,In_1131,In_543);
and U2020 (N_2020,In_320,In_560);
xnor U2021 (N_2021,In_1089,In_7);
nor U2022 (N_2022,In_799,In_1488);
nor U2023 (N_2023,In_306,In_1458);
or U2024 (N_2024,In_119,In_531);
or U2025 (N_2025,In_542,In_1390);
nor U2026 (N_2026,In_1099,In_271);
or U2027 (N_2027,In_430,In_265);
nor U2028 (N_2028,In_4,In_167);
or U2029 (N_2029,In_1291,In_818);
and U2030 (N_2030,In_1301,In_138);
nand U2031 (N_2031,In_866,In_1383);
nor U2032 (N_2032,In_101,In_1375);
and U2033 (N_2033,In_1481,In_1449);
nor U2034 (N_2034,In_474,In_123);
or U2035 (N_2035,In_358,In_1085);
or U2036 (N_2036,In_42,In_874);
nand U2037 (N_2037,In_1389,In_593);
xor U2038 (N_2038,In_1422,In_1483);
nor U2039 (N_2039,In_34,In_442);
nand U2040 (N_2040,In_1408,In_250);
nand U2041 (N_2041,In_620,In_163);
nand U2042 (N_2042,In_8,In_688);
nor U2043 (N_2043,In_460,In_299);
or U2044 (N_2044,In_45,In_427);
and U2045 (N_2045,In_1115,In_1330);
or U2046 (N_2046,In_1422,In_519);
nand U2047 (N_2047,In_682,In_250);
and U2048 (N_2048,In_1479,In_452);
or U2049 (N_2049,In_1466,In_573);
nand U2050 (N_2050,In_804,In_1185);
and U2051 (N_2051,In_1168,In_1376);
nor U2052 (N_2052,In_594,In_587);
nor U2053 (N_2053,In_644,In_1213);
and U2054 (N_2054,In_320,In_283);
nor U2055 (N_2055,In_54,In_1223);
nor U2056 (N_2056,In_1137,In_1395);
nor U2057 (N_2057,In_958,In_1466);
or U2058 (N_2058,In_120,In_1460);
nor U2059 (N_2059,In_98,In_846);
and U2060 (N_2060,In_705,In_933);
nand U2061 (N_2061,In_335,In_674);
nor U2062 (N_2062,In_104,In_1212);
or U2063 (N_2063,In_214,In_720);
or U2064 (N_2064,In_429,In_994);
nor U2065 (N_2065,In_124,In_787);
nand U2066 (N_2066,In_74,In_92);
or U2067 (N_2067,In_430,In_1059);
and U2068 (N_2068,In_169,In_1398);
nor U2069 (N_2069,In_1345,In_928);
and U2070 (N_2070,In_814,In_342);
or U2071 (N_2071,In_1152,In_114);
and U2072 (N_2072,In_164,In_97);
nor U2073 (N_2073,In_564,In_1341);
or U2074 (N_2074,In_506,In_692);
or U2075 (N_2075,In_1456,In_524);
and U2076 (N_2076,In_673,In_29);
nor U2077 (N_2077,In_426,In_99);
nor U2078 (N_2078,In_919,In_62);
and U2079 (N_2079,In_732,In_399);
xor U2080 (N_2080,In_1474,In_50);
and U2081 (N_2081,In_971,In_1375);
or U2082 (N_2082,In_641,In_141);
nand U2083 (N_2083,In_1238,In_101);
or U2084 (N_2084,In_690,In_1151);
xnor U2085 (N_2085,In_1308,In_323);
nand U2086 (N_2086,In_1063,In_932);
nor U2087 (N_2087,In_1482,In_245);
nand U2088 (N_2088,In_926,In_1011);
nor U2089 (N_2089,In_967,In_1199);
and U2090 (N_2090,In_494,In_928);
nand U2091 (N_2091,In_1192,In_1290);
or U2092 (N_2092,In_570,In_708);
nor U2093 (N_2093,In_204,In_1457);
or U2094 (N_2094,In_1247,In_201);
and U2095 (N_2095,In_628,In_700);
and U2096 (N_2096,In_678,In_1470);
or U2097 (N_2097,In_887,In_988);
nor U2098 (N_2098,In_132,In_566);
and U2099 (N_2099,In_720,In_283);
or U2100 (N_2100,In_85,In_815);
nor U2101 (N_2101,In_109,In_1133);
nand U2102 (N_2102,In_695,In_1162);
or U2103 (N_2103,In_1006,In_512);
xor U2104 (N_2104,In_942,In_1293);
nor U2105 (N_2105,In_1116,In_74);
nand U2106 (N_2106,In_1104,In_164);
and U2107 (N_2107,In_823,In_118);
and U2108 (N_2108,In_10,In_728);
nor U2109 (N_2109,In_752,In_928);
or U2110 (N_2110,In_1105,In_649);
nand U2111 (N_2111,In_449,In_316);
nor U2112 (N_2112,In_176,In_885);
or U2113 (N_2113,In_51,In_770);
or U2114 (N_2114,In_1310,In_1448);
and U2115 (N_2115,In_1303,In_1220);
and U2116 (N_2116,In_314,In_571);
and U2117 (N_2117,In_638,In_482);
or U2118 (N_2118,In_1094,In_1196);
nand U2119 (N_2119,In_878,In_264);
nand U2120 (N_2120,In_1208,In_1142);
xnor U2121 (N_2121,In_1312,In_203);
nor U2122 (N_2122,In_446,In_672);
nor U2123 (N_2123,In_942,In_213);
nor U2124 (N_2124,In_1481,In_543);
or U2125 (N_2125,In_220,In_913);
nand U2126 (N_2126,In_270,In_434);
or U2127 (N_2127,In_1122,In_120);
nor U2128 (N_2128,In_1403,In_753);
nor U2129 (N_2129,In_317,In_1298);
or U2130 (N_2130,In_1261,In_798);
and U2131 (N_2131,In_432,In_2);
and U2132 (N_2132,In_838,In_330);
nand U2133 (N_2133,In_401,In_777);
or U2134 (N_2134,In_1426,In_526);
nor U2135 (N_2135,In_1068,In_687);
nor U2136 (N_2136,In_1320,In_613);
nand U2137 (N_2137,In_462,In_391);
or U2138 (N_2138,In_802,In_1058);
or U2139 (N_2139,In_1365,In_342);
or U2140 (N_2140,In_1381,In_1094);
nor U2141 (N_2141,In_1363,In_1019);
or U2142 (N_2142,In_716,In_1003);
and U2143 (N_2143,In_34,In_650);
or U2144 (N_2144,In_1481,In_557);
nand U2145 (N_2145,In_742,In_1351);
and U2146 (N_2146,In_291,In_1272);
nor U2147 (N_2147,In_1060,In_755);
nor U2148 (N_2148,In_511,In_924);
and U2149 (N_2149,In_541,In_350);
nand U2150 (N_2150,In_803,In_39);
or U2151 (N_2151,In_56,In_1383);
and U2152 (N_2152,In_1024,In_1139);
or U2153 (N_2153,In_1391,In_1289);
and U2154 (N_2154,In_1024,In_732);
nand U2155 (N_2155,In_1182,In_1150);
or U2156 (N_2156,In_927,In_435);
and U2157 (N_2157,In_1434,In_389);
nand U2158 (N_2158,In_278,In_831);
and U2159 (N_2159,In_170,In_1193);
nor U2160 (N_2160,In_584,In_411);
and U2161 (N_2161,In_1452,In_832);
nand U2162 (N_2162,In_93,In_825);
and U2163 (N_2163,In_43,In_1342);
and U2164 (N_2164,In_1299,In_649);
nor U2165 (N_2165,In_739,In_1141);
and U2166 (N_2166,In_185,In_137);
nor U2167 (N_2167,In_1414,In_520);
nor U2168 (N_2168,In_226,In_1464);
nor U2169 (N_2169,In_783,In_61);
nand U2170 (N_2170,In_282,In_242);
xnor U2171 (N_2171,In_1335,In_1439);
and U2172 (N_2172,In_1284,In_811);
or U2173 (N_2173,In_749,In_942);
or U2174 (N_2174,In_959,In_1447);
nor U2175 (N_2175,In_1126,In_1288);
nor U2176 (N_2176,In_574,In_555);
nand U2177 (N_2177,In_203,In_234);
nand U2178 (N_2178,In_920,In_521);
and U2179 (N_2179,In_220,In_69);
or U2180 (N_2180,In_9,In_32);
or U2181 (N_2181,In_1246,In_1102);
or U2182 (N_2182,In_230,In_1221);
nand U2183 (N_2183,In_1447,In_250);
or U2184 (N_2184,In_67,In_44);
or U2185 (N_2185,In_804,In_1038);
and U2186 (N_2186,In_312,In_1184);
nand U2187 (N_2187,In_719,In_195);
and U2188 (N_2188,In_135,In_1164);
nand U2189 (N_2189,In_1449,In_888);
and U2190 (N_2190,In_747,In_207);
nor U2191 (N_2191,In_444,In_767);
or U2192 (N_2192,In_1484,In_475);
or U2193 (N_2193,In_1293,In_546);
nor U2194 (N_2194,In_1148,In_585);
and U2195 (N_2195,In_1312,In_275);
nand U2196 (N_2196,In_98,In_1413);
nand U2197 (N_2197,In_935,In_1478);
nor U2198 (N_2198,In_510,In_1199);
nand U2199 (N_2199,In_1090,In_1414);
or U2200 (N_2200,In_487,In_1317);
nor U2201 (N_2201,In_752,In_1173);
and U2202 (N_2202,In_804,In_1377);
nor U2203 (N_2203,In_1289,In_687);
or U2204 (N_2204,In_151,In_565);
and U2205 (N_2205,In_1427,In_563);
or U2206 (N_2206,In_735,In_759);
nand U2207 (N_2207,In_1299,In_808);
and U2208 (N_2208,In_1138,In_19);
nand U2209 (N_2209,In_1484,In_1240);
and U2210 (N_2210,In_779,In_144);
and U2211 (N_2211,In_607,In_697);
nand U2212 (N_2212,In_977,In_931);
nor U2213 (N_2213,In_918,In_670);
or U2214 (N_2214,In_700,In_890);
nor U2215 (N_2215,In_1377,In_1106);
nor U2216 (N_2216,In_568,In_952);
nor U2217 (N_2217,In_1391,In_574);
and U2218 (N_2218,In_840,In_695);
nor U2219 (N_2219,In_1395,In_836);
nor U2220 (N_2220,In_1326,In_286);
or U2221 (N_2221,In_1202,In_305);
nor U2222 (N_2222,In_103,In_912);
nand U2223 (N_2223,In_577,In_1055);
nand U2224 (N_2224,In_93,In_1046);
or U2225 (N_2225,In_1444,In_197);
nor U2226 (N_2226,In_515,In_539);
or U2227 (N_2227,In_1290,In_1004);
and U2228 (N_2228,In_1478,In_494);
and U2229 (N_2229,In_1161,In_1085);
nand U2230 (N_2230,In_863,In_877);
nor U2231 (N_2231,In_458,In_697);
or U2232 (N_2232,In_436,In_611);
nand U2233 (N_2233,In_65,In_345);
or U2234 (N_2234,In_1278,In_1269);
and U2235 (N_2235,In_49,In_1072);
nor U2236 (N_2236,In_832,In_842);
or U2237 (N_2237,In_788,In_158);
nor U2238 (N_2238,In_690,In_910);
xor U2239 (N_2239,In_424,In_1102);
or U2240 (N_2240,In_836,In_926);
nand U2241 (N_2241,In_1475,In_165);
nor U2242 (N_2242,In_669,In_1116);
nand U2243 (N_2243,In_25,In_1419);
nand U2244 (N_2244,In_104,In_528);
nor U2245 (N_2245,In_324,In_1041);
nand U2246 (N_2246,In_322,In_669);
nor U2247 (N_2247,In_292,In_525);
or U2248 (N_2248,In_194,In_281);
nor U2249 (N_2249,In_890,In_1025);
nand U2250 (N_2250,In_796,In_939);
and U2251 (N_2251,In_1107,In_1292);
nor U2252 (N_2252,In_36,In_1293);
and U2253 (N_2253,In_456,In_889);
nor U2254 (N_2254,In_704,In_1265);
or U2255 (N_2255,In_126,In_608);
nand U2256 (N_2256,In_1011,In_531);
nor U2257 (N_2257,In_335,In_1433);
or U2258 (N_2258,In_790,In_695);
or U2259 (N_2259,In_533,In_1367);
and U2260 (N_2260,In_806,In_1169);
and U2261 (N_2261,In_1344,In_764);
or U2262 (N_2262,In_1111,In_50);
nor U2263 (N_2263,In_140,In_554);
or U2264 (N_2264,In_227,In_835);
xor U2265 (N_2265,In_1349,In_618);
or U2266 (N_2266,In_152,In_752);
and U2267 (N_2267,In_1266,In_1045);
nand U2268 (N_2268,In_257,In_933);
and U2269 (N_2269,In_237,In_1075);
and U2270 (N_2270,In_7,In_51);
or U2271 (N_2271,In_592,In_1405);
nand U2272 (N_2272,In_302,In_630);
or U2273 (N_2273,In_1262,In_472);
nor U2274 (N_2274,In_1472,In_100);
or U2275 (N_2275,In_1033,In_1057);
nor U2276 (N_2276,In_531,In_553);
and U2277 (N_2277,In_1238,In_951);
nor U2278 (N_2278,In_1287,In_762);
and U2279 (N_2279,In_717,In_821);
nor U2280 (N_2280,In_265,In_275);
or U2281 (N_2281,In_1117,In_1196);
nand U2282 (N_2282,In_1027,In_1438);
or U2283 (N_2283,In_418,In_339);
xor U2284 (N_2284,In_1292,In_539);
nor U2285 (N_2285,In_257,In_436);
and U2286 (N_2286,In_763,In_1432);
nor U2287 (N_2287,In_339,In_877);
nor U2288 (N_2288,In_366,In_1259);
or U2289 (N_2289,In_370,In_83);
nor U2290 (N_2290,In_260,In_154);
nor U2291 (N_2291,In_241,In_1344);
and U2292 (N_2292,In_297,In_157);
nor U2293 (N_2293,In_1060,In_217);
and U2294 (N_2294,In_1400,In_669);
and U2295 (N_2295,In_583,In_505);
or U2296 (N_2296,In_1340,In_133);
nand U2297 (N_2297,In_382,In_1277);
nand U2298 (N_2298,In_910,In_1399);
nor U2299 (N_2299,In_1369,In_974);
and U2300 (N_2300,In_412,In_1389);
nor U2301 (N_2301,In_1156,In_676);
or U2302 (N_2302,In_142,In_793);
or U2303 (N_2303,In_485,In_601);
and U2304 (N_2304,In_340,In_573);
nand U2305 (N_2305,In_1022,In_628);
xor U2306 (N_2306,In_319,In_917);
nor U2307 (N_2307,In_460,In_368);
nor U2308 (N_2308,In_139,In_61);
nor U2309 (N_2309,In_1018,In_1211);
or U2310 (N_2310,In_653,In_560);
or U2311 (N_2311,In_1432,In_479);
and U2312 (N_2312,In_120,In_1165);
nor U2313 (N_2313,In_69,In_1076);
and U2314 (N_2314,In_1176,In_137);
or U2315 (N_2315,In_796,In_307);
nor U2316 (N_2316,In_68,In_715);
xnor U2317 (N_2317,In_745,In_1322);
nor U2318 (N_2318,In_238,In_320);
or U2319 (N_2319,In_94,In_1377);
nand U2320 (N_2320,In_1228,In_284);
nor U2321 (N_2321,In_1468,In_369);
nor U2322 (N_2322,In_99,In_318);
nor U2323 (N_2323,In_150,In_1218);
nand U2324 (N_2324,In_259,In_855);
or U2325 (N_2325,In_115,In_583);
nor U2326 (N_2326,In_247,In_839);
and U2327 (N_2327,In_81,In_793);
nor U2328 (N_2328,In_778,In_177);
nor U2329 (N_2329,In_407,In_1240);
nand U2330 (N_2330,In_1445,In_521);
nand U2331 (N_2331,In_308,In_888);
and U2332 (N_2332,In_688,In_395);
and U2333 (N_2333,In_492,In_341);
and U2334 (N_2334,In_148,In_326);
or U2335 (N_2335,In_779,In_113);
nor U2336 (N_2336,In_756,In_83);
or U2337 (N_2337,In_1186,In_414);
nor U2338 (N_2338,In_1155,In_836);
and U2339 (N_2339,In_1352,In_877);
nor U2340 (N_2340,In_983,In_979);
or U2341 (N_2341,In_1174,In_664);
or U2342 (N_2342,In_403,In_20);
xor U2343 (N_2343,In_1371,In_907);
nor U2344 (N_2344,In_1439,In_1429);
nor U2345 (N_2345,In_423,In_153);
nand U2346 (N_2346,In_976,In_1150);
or U2347 (N_2347,In_1032,In_421);
or U2348 (N_2348,In_1455,In_1387);
nand U2349 (N_2349,In_1370,In_1008);
nand U2350 (N_2350,In_1308,In_1150);
and U2351 (N_2351,In_1284,In_685);
nand U2352 (N_2352,In_1083,In_1304);
nor U2353 (N_2353,In_427,In_287);
nand U2354 (N_2354,In_420,In_879);
and U2355 (N_2355,In_982,In_1148);
or U2356 (N_2356,In_1375,In_358);
nand U2357 (N_2357,In_966,In_200);
and U2358 (N_2358,In_978,In_664);
and U2359 (N_2359,In_789,In_643);
nor U2360 (N_2360,In_1316,In_1131);
and U2361 (N_2361,In_700,In_438);
nor U2362 (N_2362,In_410,In_295);
nand U2363 (N_2363,In_804,In_54);
or U2364 (N_2364,In_890,In_788);
nand U2365 (N_2365,In_110,In_43);
and U2366 (N_2366,In_51,In_662);
nor U2367 (N_2367,In_1173,In_223);
and U2368 (N_2368,In_715,In_975);
or U2369 (N_2369,In_1249,In_164);
and U2370 (N_2370,In_704,In_241);
or U2371 (N_2371,In_712,In_496);
or U2372 (N_2372,In_608,In_535);
nor U2373 (N_2373,In_339,In_18);
xor U2374 (N_2374,In_1465,In_484);
nor U2375 (N_2375,In_173,In_86);
nand U2376 (N_2376,In_745,In_757);
and U2377 (N_2377,In_908,In_18);
and U2378 (N_2378,In_1084,In_1368);
nor U2379 (N_2379,In_459,In_860);
or U2380 (N_2380,In_231,In_175);
or U2381 (N_2381,In_1079,In_788);
nor U2382 (N_2382,In_849,In_667);
nand U2383 (N_2383,In_642,In_1499);
and U2384 (N_2384,In_1067,In_120);
nor U2385 (N_2385,In_951,In_1222);
or U2386 (N_2386,In_1031,In_573);
nand U2387 (N_2387,In_1253,In_305);
nor U2388 (N_2388,In_1271,In_1036);
and U2389 (N_2389,In_36,In_865);
and U2390 (N_2390,In_1142,In_53);
nor U2391 (N_2391,In_704,In_1008);
or U2392 (N_2392,In_1066,In_304);
or U2393 (N_2393,In_243,In_1353);
nor U2394 (N_2394,In_151,In_979);
and U2395 (N_2395,In_488,In_680);
or U2396 (N_2396,In_141,In_1115);
and U2397 (N_2397,In_763,In_728);
and U2398 (N_2398,In_335,In_1280);
nand U2399 (N_2399,In_1304,In_710);
nor U2400 (N_2400,In_1046,In_1037);
nand U2401 (N_2401,In_1117,In_1171);
nand U2402 (N_2402,In_903,In_726);
or U2403 (N_2403,In_343,In_1278);
nand U2404 (N_2404,In_1073,In_968);
nand U2405 (N_2405,In_1424,In_268);
or U2406 (N_2406,In_1140,In_1396);
or U2407 (N_2407,In_470,In_1172);
nor U2408 (N_2408,In_113,In_1207);
or U2409 (N_2409,In_1454,In_1416);
or U2410 (N_2410,In_460,In_713);
or U2411 (N_2411,In_1175,In_1019);
nand U2412 (N_2412,In_17,In_1015);
nor U2413 (N_2413,In_1388,In_932);
and U2414 (N_2414,In_194,In_824);
nor U2415 (N_2415,In_1095,In_600);
nor U2416 (N_2416,In_836,In_1055);
xnor U2417 (N_2417,In_734,In_1070);
and U2418 (N_2418,In_1319,In_1216);
nand U2419 (N_2419,In_1170,In_906);
nor U2420 (N_2420,In_1257,In_141);
nor U2421 (N_2421,In_770,In_764);
or U2422 (N_2422,In_312,In_125);
and U2423 (N_2423,In_909,In_53);
nor U2424 (N_2424,In_1196,In_823);
and U2425 (N_2425,In_876,In_1443);
and U2426 (N_2426,In_823,In_375);
and U2427 (N_2427,In_751,In_435);
nor U2428 (N_2428,In_446,In_62);
and U2429 (N_2429,In_603,In_1030);
and U2430 (N_2430,In_252,In_461);
and U2431 (N_2431,In_714,In_838);
or U2432 (N_2432,In_1208,In_1432);
and U2433 (N_2433,In_1375,In_1084);
and U2434 (N_2434,In_774,In_587);
nor U2435 (N_2435,In_1261,In_1113);
nor U2436 (N_2436,In_169,In_74);
nand U2437 (N_2437,In_495,In_989);
or U2438 (N_2438,In_1065,In_1061);
nand U2439 (N_2439,In_615,In_641);
nor U2440 (N_2440,In_1195,In_1057);
and U2441 (N_2441,In_385,In_843);
and U2442 (N_2442,In_1013,In_1294);
and U2443 (N_2443,In_862,In_680);
nand U2444 (N_2444,In_523,In_1300);
or U2445 (N_2445,In_140,In_1465);
nor U2446 (N_2446,In_121,In_1357);
nand U2447 (N_2447,In_438,In_1266);
nor U2448 (N_2448,In_1140,In_914);
or U2449 (N_2449,In_301,In_676);
nand U2450 (N_2450,In_924,In_845);
or U2451 (N_2451,In_1256,In_757);
nor U2452 (N_2452,In_1065,In_1233);
and U2453 (N_2453,In_1395,In_1068);
and U2454 (N_2454,In_1384,In_486);
or U2455 (N_2455,In_358,In_1200);
or U2456 (N_2456,In_1326,In_199);
nand U2457 (N_2457,In_723,In_825);
or U2458 (N_2458,In_721,In_456);
nand U2459 (N_2459,In_425,In_371);
nor U2460 (N_2460,In_483,In_1464);
nand U2461 (N_2461,In_1114,In_887);
nor U2462 (N_2462,In_629,In_648);
nor U2463 (N_2463,In_1303,In_1063);
or U2464 (N_2464,In_1166,In_1244);
or U2465 (N_2465,In_452,In_1461);
nor U2466 (N_2466,In_450,In_919);
nand U2467 (N_2467,In_879,In_516);
nand U2468 (N_2468,In_165,In_759);
and U2469 (N_2469,In_470,In_1070);
nor U2470 (N_2470,In_288,In_807);
nand U2471 (N_2471,In_1437,In_1353);
nand U2472 (N_2472,In_413,In_343);
nor U2473 (N_2473,In_248,In_1462);
nand U2474 (N_2474,In_416,In_343);
or U2475 (N_2475,In_862,In_185);
nor U2476 (N_2476,In_1054,In_823);
nand U2477 (N_2477,In_435,In_257);
xor U2478 (N_2478,In_1476,In_1018);
nor U2479 (N_2479,In_464,In_124);
or U2480 (N_2480,In_234,In_847);
or U2481 (N_2481,In_311,In_437);
and U2482 (N_2482,In_708,In_1297);
nand U2483 (N_2483,In_1415,In_630);
nand U2484 (N_2484,In_1190,In_1288);
nand U2485 (N_2485,In_871,In_1180);
or U2486 (N_2486,In_783,In_985);
and U2487 (N_2487,In_1374,In_1155);
nand U2488 (N_2488,In_256,In_638);
nand U2489 (N_2489,In_1424,In_412);
nand U2490 (N_2490,In_775,In_526);
or U2491 (N_2491,In_1354,In_347);
and U2492 (N_2492,In_1437,In_1045);
and U2493 (N_2493,In_1297,In_270);
or U2494 (N_2494,In_1427,In_1263);
and U2495 (N_2495,In_368,In_1270);
or U2496 (N_2496,In_395,In_370);
or U2497 (N_2497,In_1261,In_479);
nor U2498 (N_2498,In_662,In_1459);
xnor U2499 (N_2499,In_152,In_890);
or U2500 (N_2500,In_690,In_1041);
and U2501 (N_2501,In_483,In_486);
or U2502 (N_2502,In_459,In_1248);
or U2503 (N_2503,In_173,In_501);
or U2504 (N_2504,In_1390,In_885);
or U2505 (N_2505,In_686,In_350);
and U2506 (N_2506,In_509,In_565);
nor U2507 (N_2507,In_1385,In_147);
nand U2508 (N_2508,In_290,In_496);
or U2509 (N_2509,In_112,In_843);
nand U2510 (N_2510,In_1355,In_239);
or U2511 (N_2511,In_1315,In_522);
or U2512 (N_2512,In_296,In_360);
or U2513 (N_2513,In_1029,In_800);
or U2514 (N_2514,In_74,In_646);
and U2515 (N_2515,In_688,In_15);
nand U2516 (N_2516,In_1403,In_137);
and U2517 (N_2517,In_315,In_1104);
or U2518 (N_2518,In_1459,In_67);
or U2519 (N_2519,In_1204,In_1477);
and U2520 (N_2520,In_418,In_849);
and U2521 (N_2521,In_858,In_47);
or U2522 (N_2522,In_226,In_851);
or U2523 (N_2523,In_761,In_1060);
and U2524 (N_2524,In_141,In_1330);
xor U2525 (N_2525,In_1364,In_402);
and U2526 (N_2526,In_307,In_1278);
nor U2527 (N_2527,In_40,In_1077);
and U2528 (N_2528,In_872,In_738);
and U2529 (N_2529,In_1335,In_1176);
or U2530 (N_2530,In_168,In_529);
and U2531 (N_2531,In_1349,In_1397);
and U2532 (N_2532,In_1312,In_1199);
and U2533 (N_2533,In_1074,In_1130);
nand U2534 (N_2534,In_644,In_948);
or U2535 (N_2535,In_395,In_157);
nor U2536 (N_2536,In_1023,In_1293);
nor U2537 (N_2537,In_1253,In_998);
nor U2538 (N_2538,In_264,In_1366);
or U2539 (N_2539,In_637,In_406);
nand U2540 (N_2540,In_1452,In_449);
nor U2541 (N_2541,In_685,In_1173);
and U2542 (N_2542,In_651,In_739);
or U2543 (N_2543,In_843,In_1076);
and U2544 (N_2544,In_1063,In_348);
or U2545 (N_2545,In_887,In_1027);
nor U2546 (N_2546,In_735,In_1028);
or U2547 (N_2547,In_53,In_488);
nor U2548 (N_2548,In_995,In_85);
and U2549 (N_2549,In_33,In_1069);
nor U2550 (N_2550,In_1254,In_519);
nor U2551 (N_2551,In_957,In_1077);
and U2552 (N_2552,In_1026,In_1377);
or U2553 (N_2553,In_1288,In_598);
nor U2554 (N_2554,In_1135,In_1238);
nand U2555 (N_2555,In_53,In_583);
nand U2556 (N_2556,In_170,In_1328);
or U2557 (N_2557,In_1033,In_801);
nand U2558 (N_2558,In_170,In_516);
or U2559 (N_2559,In_897,In_1332);
nor U2560 (N_2560,In_507,In_1221);
or U2561 (N_2561,In_77,In_243);
nand U2562 (N_2562,In_1417,In_895);
or U2563 (N_2563,In_394,In_840);
or U2564 (N_2564,In_797,In_481);
nor U2565 (N_2565,In_1403,In_578);
nand U2566 (N_2566,In_1054,In_1435);
and U2567 (N_2567,In_270,In_223);
nor U2568 (N_2568,In_604,In_705);
or U2569 (N_2569,In_993,In_340);
or U2570 (N_2570,In_518,In_329);
nand U2571 (N_2571,In_13,In_382);
nor U2572 (N_2572,In_1291,In_760);
and U2573 (N_2573,In_1060,In_33);
and U2574 (N_2574,In_1446,In_479);
or U2575 (N_2575,In_1389,In_283);
or U2576 (N_2576,In_1008,In_404);
nand U2577 (N_2577,In_1175,In_22);
and U2578 (N_2578,In_158,In_403);
and U2579 (N_2579,In_895,In_1319);
and U2580 (N_2580,In_1277,In_737);
nand U2581 (N_2581,In_745,In_836);
nor U2582 (N_2582,In_480,In_1022);
and U2583 (N_2583,In_314,In_198);
or U2584 (N_2584,In_202,In_514);
nand U2585 (N_2585,In_1110,In_484);
nor U2586 (N_2586,In_1011,In_1004);
or U2587 (N_2587,In_33,In_1024);
nand U2588 (N_2588,In_353,In_115);
and U2589 (N_2589,In_1457,In_1335);
or U2590 (N_2590,In_720,In_1118);
nor U2591 (N_2591,In_458,In_1014);
or U2592 (N_2592,In_1476,In_1339);
nand U2593 (N_2593,In_412,In_57);
or U2594 (N_2594,In_793,In_281);
or U2595 (N_2595,In_582,In_371);
and U2596 (N_2596,In_78,In_297);
and U2597 (N_2597,In_1298,In_800);
and U2598 (N_2598,In_589,In_10);
or U2599 (N_2599,In_1136,In_740);
or U2600 (N_2600,In_787,In_1284);
nor U2601 (N_2601,In_1384,In_35);
nor U2602 (N_2602,In_79,In_1324);
xor U2603 (N_2603,In_557,In_466);
nor U2604 (N_2604,In_262,In_31);
nand U2605 (N_2605,In_339,In_1148);
or U2606 (N_2606,In_375,In_920);
nand U2607 (N_2607,In_41,In_686);
nand U2608 (N_2608,In_247,In_973);
and U2609 (N_2609,In_471,In_599);
nand U2610 (N_2610,In_225,In_1188);
and U2611 (N_2611,In_47,In_718);
or U2612 (N_2612,In_296,In_310);
and U2613 (N_2613,In_689,In_1173);
nor U2614 (N_2614,In_12,In_1054);
nor U2615 (N_2615,In_1368,In_529);
nor U2616 (N_2616,In_754,In_328);
nand U2617 (N_2617,In_103,In_217);
or U2618 (N_2618,In_505,In_1444);
and U2619 (N_2619,In_1345,In_659);
or U2620 (N_2620,In_3,In_1074);
nor U2621 (N_2621,In_681,In_227);
and U2622 (N_2622,In_353,In_572);
or U2623 (N_2623,In_602,In_445);
nor U2624 (N_2624,In_293,In_1046);
and U2625 (N_2625,In_561,In_446);
or U2626 (N_2626,In_1324,In_1238);
nor U2627 (N_2627,In_1246,In_4);
nand U2628 (N_2628,In_1150,In_196);
or U2629 (N_2629,In_886,In_694);
nor U2630 (N_2630,In_81,In_516);
or U2631 (N_2631,In_1180,In_247);
and U2632 (N_2632,In_785,In_985);
nand U2633 (N_2633,In_1029,In_1030);
nand U2634 (N_2634,In_708,In_618);
or U2635 (N_2635,In_1325,In_989);
or U2636 (N_2636,In_959,In_746);
and U2637 (N_2637,In_435,In_678);
and U2638 (N_2638,In_280,In_1000);
nand U2639 (N_2639,In_65,In_553);
or U2640 (N_2640,In_1240,In_770);
or U2641 (N_2641,In_805,In_851);
nand U2642 (N_2642,In_866,In_593);
and U2643 (N_2643,In_1316,In_1269);
and U2644 (N_2644,In_397,In_309);
xor U2645 (N_2645,In_245,In_933);
or U2646 (N_2646,In_895,In_703);
xor U2647 (N_2647,In_803,In_1005);
and U2648 (N_2648,In_375,In_1250);
and U2649 (N_2649,In_1070,In_822);
and U2650 (N_2650,In_1170,In_683);
nor U2651 (N_2651,In_884,In_1453);
nor U2652 (N_2652,In_109,In_827);
or U2653 (N_2653,In_541,In_1381);
nor U2654 (N_2654,In_1155,In_1050);
nand U2655 (N_2655,In_644,In_165);
nand U2656 (N_2656,In_799,In_79);
nand U2657 (N_2657,In_433,In_1084);
or U2658 (N_2658,In_1099,In_1467);
or U2659 (N_2659,In_357,In_245);
or U2660 (N_2660,In_728,In_653);
and U2661 (N_2661,In_1219,In_266);
and U2662 (N_2662,In_891,In_548);
or U2663 (N_2663,In_1076,In_403);
xnor U2664 (N_2664,In_1279,In_847);
nor U2665 (N_2665,In_1078,In_1412);
or U2666 (N_2666,In_446,In_848);
nor U2667 (N_2667,In_1146,In_1076);
or U2668 (N_2668,In_698,In_293);
nand U2669 (N_2669,In_1147,In_903);
nand U2670 (N_2670,In_1073,In_55);
or U2671 (N_2671,In_416,In_840);
and U2672 (N_2672,In_1162,In_557);
and U2673 (N_2673,In_405,In_564);
nand U2674 (N_2674,In_241,In_1111);
nand U2675 (N_2675,In_1028,In_462);
nand U2676 (N_2676,In_1041,In_921);
nand U2677 (N_2677,In_172,In_953);
nor U2678 (N_2678,In_317,In_951);
nor U2679 (N_2679,In_55,In_538);
nand U2680 (N_2680,In_788,In_1041);
or U2681 (N_2681,In_484,In_980);
and U2682 (N_2682,In_926,In_212);
or U2683 (N_2683,In_976,In_995);
and U2684 (N_2684,In_39,In_166);
and U2685 (N_2685,In_858,In_1065);
and U2686 (N_2686,In_465,In_564);
nand U2687 (N_2687,In_1496,In_609);
and U2688 (N_2688,In_1498,In_131);
and U2689 (N_2689,In_201,In_730);
and U2690 (N_2690,In_245,In_99);
and U2691 (N_2691,In_985,In_695);
nand U2692 (N_2692,In_844,In_1144);
nor U2693 (N_2693,In_807,In_372);
nand U2694 (N_2694,In_285,In_354);
and U2695 (N_2695,In_315,In_186);
and U2696 (N_2696,In_1346,In_972);
or U2697 (N_2697,In_96,In_1373);
or U2698 (N_2698,In_106,In_165);
and U2699 (N_2699,In_755,In_528);
nor U2700 (N_2700,In_360,In_48);
and U2701 (N_2701,In_1388,In_1395);
nor U2702 (N_2702,In_1005,In_1382);
nand U2703 (N_2703,In_1436,In_493);
nor U2704 (N_2704,In_316,In_734);
and U2705 (N_2705,In_1219,In_1251);
nor U2706 (N_2706,In_648,In_540);
or U2707 (N_2707,In_100,In_693);
and U2708 (N_2708,In_976,In_483);
nor U2709 (N_2709,In_372,In_1362);
or U2710 (N_2710,In_1361,In_625);
nand U2711 (N_2711,In_619,In_1222);
and U2712 (N_2712,In_1184,In_198);
nand U2713 (N_2713,In_340,In_1218);
nand U2714 (N_2714,In_405,In_239);
nor U2715 (N_2715,In_895,In_690);
nand U2716 (N_2716,In_142,In_1375);
and U2717 (N_2717,In_320,In_1291);
nand U2718 (N_2718,In_149,In_1465);
or U2719 (N_2719,In_944,In_386);
nand U2720 (N_2720,In_424,In_1474);
or U2721 (N_2721,In_670,In_1296);
or U2722 (N_2722,In_1237,In_1309);
or U2723 (N_2723,In_742,In_1288);
or U2724 (N_2724,In_907,In_403);
and U2725 (N_2725,In_741,In_193);
or U2726 (N_2726,In_0,In_667);
or U2727 (N_2727,In_1334,In_769);
nand U2728 (N_2728,In_827,In_1134);
and U2729 (N_2729,In_85,In_1440);
and U2730 (N_2730,In_737,In_465);
nand U2731 (N_2731,In_296,In_455);
xor U2732 (N_2732,In_1414,In_665);
nand U2733 (N_2733,In_1472,In_523);
nand U2734 (N_2734,In_318,In_1269);
or U2735 (N_2735,In_1286,In_633);
and U2736 (N_2736,In_1181,In_1307);
nor U2737 (N_2737,In_1244,In_170);
nor U2738 (N_2738,In_1407,In_166);
nand U2739 (N_2739,In_994,In_1429);
and U2740 (N_2740,In_1108,In_1186);
or U2741 (N_2741,In_1109,In_70);
and U2742 (N_2742,In_715,In_980);
or U2743 (N_2743,In_1452,In_79);
or U2744 (N_2744,In_1046,In_1476);
nor U2745 (N_2745,In_671,In_1246);
nand U2746 (N_2746,In_211,In_1480);
nand U2747 (N_2747,In_1429,In_207);
xnor U2748 (N_2748,In_313,In_1398);
or U2749 (N_2749,In_1276,In_573);
or U2750 (N_2750,In_375,In_866);
and U2751 (N_2751,In_330,In_21);
and U2752 (N_2752,In_388,In_1280);
nor U2753 (N_2753,In_353,In_212);
and U2754 (N_2754,In_286,In_1372);
or U2755 (N_2755,In_188,In_590);
or U2756 (N_2756,In_622,In_894);
nor U2757 (N_2757,In_259,In_758);
and U2758 (N_2758,In_1132,In_835);
nor U2759 (N_2759,In_788,In_533);
and U2760 (N_2760,In_694,In_483);
nor U2761 (N_2761,In_368,In_1087);
nor U2762 (N_2762,In_314,In_381);
nand U2763 (N_2763,In_1284,In_218);
nor U2764 (N_2764,In_999,In_1314);
and U2765 (N_2765,In_160,In_672);
and U2766 (N_2766,In_1429,In_384);
and U2767 (N_2767,In_1100,In_281);
and U2768 (N_2768,In_1053,In_28);
nand U2769 (N_2769,In_1209,In_1121);
or U2770 (N_2770,In_421,In_515);
and U2771 (N_2771,In_699,In_1033);
and U2772 (N_2772,In_964,In_694);
nand U2773 (N_2773,In_384,In_49);
nor U2774 (N_2774,In_1267,In_906);
nand U2775 (N_2775,In_1267,In_33);
nand U2776 (N_2776,In_231,In_539);
and U2777 (N_2777,In_539,In_818);
or U2778 (N_2778,In_739,In_89);
nor U2779 (N_2779,In_1422,In_972);
nand U2780 (N_2780,In_112,In_1224);
nand U2781 (N_2781,In_1320,In_1236);
and U2782 (N_2782,In_1299,In_1308);
and U2783 (N_2783,In_424,In_60);
nor U2784 (N_2784,In_1198,In_370);
and U2785 (N_2785,In_85,In_744);
and U2786 (N_2786,In_946,In_185);
nor U2787 (N_2787,In_198,In_1014);
nor U2788 (N_2788,In_720,In_1424);
and U2789 (N_2789,In_1032,In_573);
or U2790 (N_2790,In_1463,In_308);
or U2791 (N_2791,In_492,In_801);
or U2792 (N_2792,In_1283,In_244);
nor U2793 (N_2793,In_703,In_1318);
and U2794 (N_2794,In_1386,In_1095);
nor U2795 (N_2795,In_927,In_157);
or U2796 (N_2796,In_879,In_825);
nor U2797 (N_2797,In_635,In_432);
and U2798 (N_2798,In_855,In_1284);
nand U2799 (N_2799,In_694,In_837);
xor U2800 (N_2800,In_820,In_646);
or U2801 (N_2801,In_196,In_1017);
nor U2802 (N_2802,In_1266,In_335);
nor U2803 (N_2803,In_1114,In_369);
nor U2804 (N_2804,In_1402,In_588);
nand U2805 (N_2805,In_848,In_1148);
and U2806 (N_2806,In_119,In_1285);
and U2807 (N_2807,In_146,In_382);
or U2808 (N_2808,In_452,In_754);
or U2809 (N_2809,In_463,In_255);
nor U2810 (N_2810,In_176,In_906);
xnor U2811 (N_2811,In_644,In_326);
nor U2812 (N_2812,In_799,In_181);
nand U2813 (N_2813,In_1457,In_514);
nand U2814 (N_2814,In_886,In_337);
or U2815 (N_2815,In_964,In_1410);
nor U2816 (N_2816,In_215,In_35);
and U2817 (N_2817,In_872,In_785);
nand U2818 (N_2818,In_1454,In_112);
or U2819 (N_2819,In_735,In_336);
nand U2820 (N_2820,In_874,In_211);
and U2821 (N_2821,In_208,In_1355);
or U2822 (N_2822,In_1483,In_233);
or U2823 (N_2823,In_939,In_381);
nor U2824 (N_2824,In_414,In_1436);
and U2825 (N_2825,In_436,In_512);
nand U2826 (N_2826,In_818,In_1357);
nor U2827 (N_2827,In_796,In_85);
and U2828 (N_2828,In_1358,In_752);
nor U2829 (N_2829,In_1193,In_1033);
xor U2830 (N_2830,In_1239,In_445);
and U2831 (N_2831,In_433,In_43);
nand U2832 (N_2832,In_1112,In_338);
nand U2833 (N_2833,In_1177,In_32);
or U2834 (N_2834,In_574,In_148);
or U2835 (N_2835,In_117,In_792);
nand U2836 (N_2836,In_1316,In_562);
nor U2837 (N_2837,In_868,In_1262);
nand U2838 (N_2838,In_924,In_556);
nor U2839 (N_2839,In_850,In_1447);
nand U2840 (N_2840,In_62,In_1116);
or U2841 (N_2841,In_712,In_500);
or U2842 (N_2842,In_330,In_931);
and U2843 (N_2843,In_377,In_277);
nand U2844 (N_2844,In_91,In_1135);
nor U2845 (N_2845,In_474,In_263);
nor U2846 (N_2846,In_976,In_1098);
xnor U2847 (N_2847,In_646,In_810);
nor U2848 (N_2848,In_1054,In_455);
nand U2849 (N_2849,In_141,In_80);
nand U2850 (N_2850,In_778,In_419);
or U2851 (N_2851,In_1180,In_655);
nand U2852 (N_2852,In_1227,In_676);
nor U2853 (N_2853,In_707,In_453);
nand U2854 (N_2854,In_1099,In_1092);
nand U2855 (N_2855,In_1310,In_738);
nand U2856 (N_2856,In_742,In_555);
or U2857 (N_2857,In_383,In_59);
or U2858 (N_2858,In_130,In_829);
nor U2859 (N_2859,In_484,In_532);
nor U2860 (N_2860,In_1380,In_894);
or U2861 (N_2861,In_325,In_1090);
nand U2862 (N_2862,In_1255,In_534);
nand U2863 (N_2863,In_910,In_538);
nand U2864 (N_2864,In_1396,In_294);
nor U2865 (N_2865,In_1144,In_301);
nand U2866 (N_2866,In_261,In_1229);
nand U2867 (N_2867,In_1420,In_1030);
or U2868 (N_2868,In_12,In_390);
nor U2869 (N_2869,In_654,In_207);
nor U2870 (N_2870,In_342,In_521);
nor U2871 (N_2871,In_356,In_429);
and U2872 (N_2872,In_932,In_155);
nand U2873 (N_2873,In_918,In_216);
or U2874 (N_2874,In_153,In_1237);
and U2875 (N_2875,In_1039,In_853);
nor U2876 (N_2876,In_597,In_229);
nand U2877 (N_2877,In_813,In_1358);
nor U2878 (N_2878,In_614,In_1332);
nor U2879 (N_2879,In_1447,In_260);
or U2880 (N_2880,In_612,In_359);
and U2881 (N_2881,In_848,In_887);
and U2882 (N_2882,In_698,In_301);
nand U2883 (N_2883,In_1072,In_174);
nand U2884 (N_2884,In_558,In_530);
and U2885 (N_2885,In_322,In_1442);
nand U2886 (N_2886,In_1294,In_240);
or U2887 (N_2887,In_425,In_1357);
nand U2888 (N_2888,In_1298,In_364);
or U2889 (N_2889,In_614,In_1319);
nor U2890 (N_2890,In_706,In_257);
nand U2891 (N_2891,In_379,In_1071);
and U2892 (N_2892,In_1155,In_1107);
nor U2893 (N_2893,In_212,In_1229);
nand U2894 (N_2894,In_901,In_306);
nor U2895 (N_2895,In_772,In_146);
nor U2896 (N_2896,In_563,In_40);
nand U2897 (N_2897,In_97,In_1419);
or U2898 (N_2898,In_1112,In_211);
nand U2899 (N_2899,In_1205,In_450);
or U2900 (N_2900,In_1461,In_1323);
or U2901 (N_2901,In_1400,In_1173);
and U2902 (N_2902,In_194,In_1052);
xor U2903 (N_2903,In_1426,In_613);
nand U2904 (N_2904,In_282,In_1209);
nand U2905 (N_2905,In_782,In_713);
or U2906 (N_2906,In_1084,In_1202);
and U2907 (N_2907,In_1164,In_1049);
nor U2908 (N_2908,In_972,In_156);
nor U2909 (N_2909,In_863,In_251);
and U2910 (N_2910,In_1456,In_629);
nand U2911 (N_2911,In_1181,In_1483);
and U2912 (N_2912,In_1466,In_641);
and U2913 (N_2913,In_841,In_1247);
nand U2914 (N_2914,In_976,In_806);
and U2915 (N_2915,In_471,In_733);
and U2916 (N_2916,In_974,In_79);
nor U2917 (N_2917,In_801,In_732);
nor U2918 (N_2918,In_1324,In_31);
nand U2919 (N_2919,In_598,In_1308);
nand U2920 (N_2920,In_143,In_959);
nand U2921 (N_2921,In_449,In_630);
and U2922 (N_2922,In_1073,In_594);
nand U2923 (N_2923,In_301,In_639);
and U2924 (N_2924,In_1432,In_381);
or U2925 (N_2925,In_1135,In_1155);
nand U2926 (N_2926,In_1124,In_770);
and U2927 (N_2927,In_680,In_67);
or U2928 (N_2928,In_1339,In_832);
nor U2929 (N_2929,In_419,In_1371);
nand U2930 (N_2930,In_1301,In_230);
nand U2931 (N_2931,In_462,In_450);
nor U2932 (N_2932,In_165,In_950);
nand U2933 (N_2933,In_1186,In_580);
and U2934 (N_2934,In_791,In_456);
nor U2935 (N_2935,In_1467,In_281);
and U2936 (N_2936,In_1347,In_694);
or U2937 (N_2937,In_37,In_1078);
and U2938 (N_2938,In_1277,In_201);
or U2939 (N_2939,In_451,In_1453);
and U2940 (N_2940,In_935,In_672);
or U2941 (N_2941,In_1020,In_273);
or U2942 (N_2942,In_384,In_192);
nand U2943 (N_2943,In_705,In_378);
nor U2944 (N_2944,In_740,In_1129);
nor U2945 (N_2945,In_656,In_162);
nand U2946 (N_2946,In_48,In_121);
nor U2947 (N_2947,In_5,In_951);
nor U2948 (N_2948,In_723,In_828);
and U2949 (N_2949,In_81,In_186);
and U2950 (N_2950,In_474,In_724);
nand U2951 (N_2951,In_1495,In_581);
nor U2952 (N_2952,In_1491,In_113);
nor U2953 (N_2953,In_170,In_979);
nand U2954 (N_2954,In_586,In_155);
xor U2955 (N_2955,In_270,In_1078);
nor U2956 (N_2956,In_1075,In_1282);
and U2957 (N_2957,In_549,In_172);
nor U2958 (N_2958,In_264,In_863);
nand U2959 (N_2959,In_1446,In_15);
or U2960 (N_2960,In_1321,In_1070);
nand U2961 (N_2961,In_316,In_517);
and U2962 (N_2962,In_502,In_473);
or U2963 (N_2963,In_1274,In_531);
and U2964 (N_2964,In_1042,In_1153);
or U2965 (N_2965,In_75,In_650);
and U2966 (N_2966,In_1347,In_1268);
nor U2967 (N_2967,In_930,In_125);
nor U2968 (N_2968,In_864,In_765);
and U2969 (N_2969,In_1131,In_1433);
nand U2970 (N_2970,In_580,In_1172);
xnor U2971 (N_2971,In_303,In_228);
or U2972 (N_2972,In_247,In_1315);
or U2973 (N_2973,In_1260,In_201);
nand U2974 (N_2974,In_447,In_893);
nand U2975 (N_2975,In_959,In_216);
or U2976 (N_2976,In_374,In_813);
nand U2977 (N_2977,In_877,In_1198);
nand U2978 (N_2978,In_193,In_1359);
or U2979 (N_2979,In_1475,In_975);
or U2980 (N_2980,In_454,In_362);
or U2981 (N_2981,In_705,In_501);
nand U2982 (N_2982,In_977,In_1011);
xnor U2983 (N_2983,In_549,In_833);
and U2984 (N_2984,In_232,In_1357);
nand U2985 (N_2985,In_1307,In_1315);
xor U2986 (N_2986,In_343,In_697);
and U2987 (N_2987,In_23,In_85);
nand U2988 (N_2988,In_1459,In_1098);
or U2989 (N_2989,In_477,In_588);
and U2990 (N_2990,In_629,In_679);
and U2991 (N_2991,In_914,In_111);
nand U2992 (N_2992,In_969,In_552);
nand U2993 (N_2993,In_383,In_302);
nor U2994 (N_2994,In_175,In_372);
nor U2995 (N_2995,In_874,In_1155);
or U2996 (N_2996,In_808,In_1151);
nand U2997 (N_2997,In_1022,In_1023);
nand U2998 (N_2998,In_54,In_1244);
and U2999 (N_2999,In_1491,In_809);
nand U3000 (N_3000,N_372,N_2192);
and U3001 (N_3001,N_2466,N_2439);
nor U3002 (N_3002,N_684,N_1782);
nand U3003 (N_3003,N_336,N_2414);
nand U3004 (N_3004,N_1497,N_1536);
nand U3005 (N_3005,N_1893,N_2313);
nand U3006 (N_3006,N_2462,N_2868);
and U3007 (N_3007,N_491,N_854);
and U3008 (N_3008,N_979,N_2693);
or U3009 (N_3009,N_999,N_663);
nor U3010 (N_3010,N_642,N_2833);
or U3011 (N_3011,N_2514,N_1472);
nand U3012 (N_3012,N_437,N_1896);
and U3013 (N_3013,N_247,N_244);
nand U3014 (N_3014,N_992,N_260);
nand U3015 (N_3015,N_623,N_1729);
and U3016 (N_3016,N_697,N_1609);
nand U3017 (N_3017,N_781,N_2948);
nand U3018 (N_3018,N_2130,N_1561);
or U3019 (N_3019,N_2206,N_2870);
or U3020 (N_3020,N_172,N_2594);
nor U3021 (N_3021,N_1097,N_1725);
nand U3022 (N_3022,N_2639,N_267);
and U3023 (N_3023,N_1200,N_2068);
and U3024 (N_3024,N_1899,N_1891);
nand U3025 (N_3025,N_2178,N_780);
or U3026 (N_3026,N_421,N_231);
nor U3027 (N_3027,N_2698,N_2054);
and U3028 (N_3028,N_1921,N_707);
nor U3029 (N_3029,N_2658,N_713);
and U3030 (N_3030,N_2747,N_2685);
nor U3031 (N_3031,N_1713,N_2898);
and U3032 (N_3032,N_811,N_1836);
and U3033 (N_3033,N_10,N_986);
or U3034 (N_3034,N_1979,N_2857);
and U3035 (N_3035,N_925,N_718);
and U3036 (N_3036,N_2989,N_2910);
and U3037 (N_3037,N_755,N_1201);
xor U3038 (N_3038,N_541,N_2542);
nand U3039 (N_3039,N_1682,N_1249);
or U3040 (N_3040,N_419,N_2449);
and U3041 (N_3041,N_2999,N_2271);
nand U3042 (N_3042,N_56,N_2617);
and U3043 (N_3043,N_2456,N_2064);
or U3044 (N_3044,N_1614,N_1586);
nor U3045 (N_3045,N_535,N_1428);
and U3046 (N_3046,N_2880,N_2166);
nand U3047 (N_3047,N_1294,N_629);
nor U3048 (N_3048,N_2330,N_1569);
nor U3049 (N_3049,N_1911,N_392);
nand U3050 (N_3050,N_2032,N_2173);
nor U3051 (N_3051,N_2279,N_2382);
nand U3052 (N_3052,N_277,N_2866);
and U3053 (N_3053,N_433,N_1761);
nor U3054 (N_3054,N_996,N_2583);
nor U3055 (N_3055,N_2849,N_168);
or U3056 (N_3056,N_1997,N_2308);
and U3057 (N_3057,N_1041,N_1388);
and U3058 (N_3058,N_1494,N_2713);
or U3059 (N_3059,N_1898,N_2426);
xnor U3060 (N_3060,N_2520,N_2453);
or U3061 (N_3061,N_11,N_2306);
xor U3062 (N_3062,N_2077,N_1033);
or U3063 (N_3063,N_1545,N_1463);
or U3064 (N_3064,N_2180,N_1150);
nand U3065 (N_3065,N_2268,N_2315);
nor U3066 (N_3066,N_2018,N_2042);
and U3067 (N_3067,N_1177,N_1853);
nor U3068 (N_3068,N_2679,N_1110);
or U3069 (N_3069,N_2204,N_2103);
nand U3070 (N_3070,N_1863,N_2415);
or U3071 (N_3071,N_2067,N_2988);
nor U3072 (N_3072,N_1931,N_685);
or U3073 (N_3073,N_1877,N_2794);
nor U3074 (N_3074,N_373,N_2319);
nor U3075 (N_3075,N_332,N_468);
nor U3076 (N_3076,N_2863,N_2758);
or U3077 (N_3077,N_2263,N_2247);
or U3078 (N_3078,N_1669,N_2288);
nor U3079 (N_3079,N_1302,N_98);
nand U3080 (N_3080,N_1115,N_1289);
nand U3081 (N_3081,N_611,N_2629);
nor U3082 (N_3082,N_211,N_1990);
or U3083 (N_3083,N_1337,N_601);
and U3084 (N_3084,N_758,N_2580);
nand U3085 (N_3085,N_1651,N_2187);
nand U3086 (N_3086,N_1399,N_2641);
or U3087 (N_3087,N_632,N_99);
nand U3088 (N_3088,N_2145,N_737);
or U3089 (N_3089,N_1356,N_2797);
or U3090 (N_3090,N_1544,N_2702);
or U3091 (N_3091,N_1269,N_1687);
nand U3092 (N_3092,N_112,N_2371);
or U3093 (N_3093,N_2655,N_1319);
nor U3094 (N_3094,N_1955,N_8);
nand U3095 (N_3095,N_1724,N_2266);
and U3096 (N_3096,N_167,N_575);
nand U3097 (N_3097,N_1112,N_1897);
nand U3098 (N_3098,N_1883,N_1610);
nor U3099 (N_3099,N_2927,N_1776);
and U3100 (N_3100,N_2841,N_1625);
nand U3101 (N_3101,N_2984,N_2222);
nand U3102 (N_3102,N_2390,N_2095);
nand U3103 (N_3103,N_215,N_2671);
nand U3104 (N_3104,N_1787,N_1040);
or U3105 (N_3105,N_2590,N_1263);
nand U3106 (N_3106,N_2132,N_2888);
and U3107 (N_3107,N_1973,N_711);
nor U3108 (N_3108,N_1262,N_2516);
nor U3109 (N_3109,N_916,N_953);
and U3110 (N_3110,N_2460,N_994);
nand U3111 (N_3111,N_2924,N_1322);
and U3112 (N_3112,N_2640,N_627);
nor U3113 (N_3113,N_1312,N_683);
nand U3114 (N_3114,N_2485,N_1556);
nand U3115 (N_3115,N_538,N_599);
and U3116 (N_3116,N_2316,N_886);
nor U3117 (N_3117,N_101,N_843);
and U3118 (N_3118,N_2684,N_2527);
and U3119 (N_3119,N_263,N_525);
and U3120 (N_3120,N_1437,N_816);
nand U3121 (N_3121,N_2047,N_2842);
and U3122 (N_3122,N_92,N_184);
nand U3123 (N_3123,N_2404,N_2269);
nand U3124 (N_3124,N_1274,N_2930);
nor U3125 (N_3125,N_2473,N_258);
nor U3126 (N_3126,N_1620,N_1500);
and U3127 (N_3127,N_1382,N_2048);
and U3128 (N_3128,N_760,N_2987);
or U3129 (N_3129,N_2962,N_118);
nand U3130 (N_3130,N_1922,N_1491);
nor U3131 (N_3131,N_2447,N_2537);
or U3132 (N_3132,N_1080,N_785);
and U3133 (N_3133,N_411,N_865);
nand U3134 (N_3134,N_475,N_156);
or U3135 (N_3135,N_1368,N_1416);
nor U3136 (N_3136,N_1422,N_770);
nor U3137 (N_3137,N_578,N_2109);
and U3138 (N_3138,N_300,N_233);
or U3139 (N_3139,N_2899,N_763);
or U3140 (N_3140,N_793,N_1583);
nor U3141 (N_3141,N_2376,N_2710);
nor U3142 (N_3142,N_1241,N_2219);
or U3143 (N_3143,N_797,N_688);
or U3144 (N_3144,N_226,N_1275);
or U3145 (N_3145,N_504,N_456);
nor U3146 (N_3146,N_2270,N_2091);
xor U3147 (N_3147,N_577,N_1732);
nand U3148 (N_3148,N_2723,N_2153);
nand U3149 (N_3149,N_1044,N_2181);
nand U3150 (N_3150,N_828,N_2920);
nor U3151 (N_3151,N_1601,N_2043);
nor U3152 (N_3152,N_308,N_2718);
and U3153 (N_3153,N_1783,N_1435);
and U3154 (N_3154,N_815,N_894);
nand U3155 (N_3155,N_2726,N_102);
or U3156 (N_3156,N_1128,N_956);
nor U3157 (N_3157,N_2167,N_1876);
and U3158 (N_3158,N_1498,N_1690);
and U3159 (N_3159,N_1006,N_1693);
or U3160 (N_3160,N_1704,N_2776);
or U3161 (N_3161,N_2163,N_867);
nand U3162 (N_3162,N_2258,N_1756);
nand U3163 (N_3163,N_1144,N_2400);
nand U3164 (N_3164,N_1096,N_2618);
nand U3165 (N_3165,N_667,N_2364);
nand U3166 (N_3166,N_939,N_178);
and U3167 (N_3167,N_1377,N_1509);
xor U3168 (N_3168,N_1092,N_1767);
nand U3169 (N_3169,N_930,N_1471);
or U3170 (N_3170,N_1451,N_2585);
or U3171 (N_3171,N_1467,N_495);
nand U3172 (N_3172,N_2416,N_1082);
or U3173 (N_3173,N_526,N_633);
nand U3174 (N_3174,N_7,N_2809);
or U3175 (N_3175,N_2242,N_249);
and U3176 (N_3176,N_1532,N_2100);
and U3177 (N_3177,N_669,N_379);
and U3178 (N_3178,N_1234,N_428);
xor U3179 (N_3179,N_1228,N_2309);
and U3180 (N_3180,N_1306,N_1659);
nand U3181 (N_3181,N_2628,N_424);
nor U3182 (N_3182,N_2484,N_2452);
nor U3183 (N_3183,N_2804,N_1236);
or U3184 (N_3184,N_1197,N_2276);
or U3185 (N_3185,N_1167,N_16);
nand U3186 (N_3186,N_228,N_870);
and U3187 (N_3187,N_1159,N_851);
nand U3188 (N_3188,N_62,N_1606);
nand U3189 (N_3189,N_144,N_682);
and U3190 (N_3190,N_443,N_808);
nand U3191 (N_3191,N_2738,N_2946);
nor U3192 (N_3192,N_1304,N_1022);
nand U3193 (N_3193,N_2234,N_2184);
and U3194 (N_3194,N_321,N_941);
nor U3195 (N_3195,N_1255,N_501);
and U3196 (N_3196,N_1492,N_2424);
nor U3197 (N_3197,N_2409,N_33);
and U3198 (N_3198,N_1213,N_1176);
or U3199 (N_3199,N_1061,N_2335);
nor U3200 (N_3200,N_1345,N_1443);
nand U3201 (N_3201,N_1420,N_1157);
nor U3202 (N_3202,N_2207,N_1615);
nor U3203 (N_3203,N_351,N_2521);
nor U3204 (N_3204,N_1487,N_27);
nand U3205 (N_3205,N_967,N_1285);
and U3206 (N_3206,N_1266,N_192);
or U3207 (N_3207,N_1519,N_2372);
nand U3208 (N_3208,N_426,N_1702);
or U3209 (N_3209,N_910,N_1951);
or U3210 (N_3210,N_1215,N_2593);
nand U3211 (N_3211,N_2096,N_1632);
nor U3212 (N_3212,N_1242,N_2929);
or U3213 (N_3213,N_1709,N_1282);
or U3214 (N_3214,N_847,N_639);
nor U3215 (N_3215,N_1064,N_1980);
nor U3216 (N_3216,N_46,N_2186);
and U3217 (N_3217,N_1715,N_2046);
xor U3218 (N_3218,N_777,N_1804);
or U3219 (N_3219,N_2651,N_2122);
nand U3220 (N_3220,N_230,N_1387);
or U3221 (N_3221,N_2119,N_2255);
and U3222 (N_3222,N_1649,N_1160);
or U3223 (N_3223,N_0,N_1111);
and U3224 (N_3224,N_1790,N_944);
xor U3225 (N_3225,N_2800,N_1999);
nand U3226 (N_3226,N_554,N_1245);
or U3227 (N_3227,N_963,N_2076);
nor U3228 (N_3228,N_2027,N_521);
or U3229 (N_3229,N_948,N_1404);
or U3230 (N_3230,N_1698,N_418);
nor U3231 (N_3231,N_1385,N_1101);
and U3232 (N_3232,N_761,N_119);
nor U3233 (N_3233,N_1888,N_2872);
nand U3234 (N_3234,N_2297,N_1460);
or U3235 (N_3235,N_2025,N_1063);
nand U3236 (N_3236,N_1260,N_2762);
and U3237 (N_3237,N_626,N_2835);
nand U3238 (N_3238,N_2867,N_269);
or U3239 (N_3239,N_1462,N_2189);
and U3240 (N_3240,N_1,N_1524);
or U3241 (N_3241,N_756,N_561);
nor U3242 (N_3242,N_951,N_1009);
nand U3243 (N_3243,N_1954,N_224);
or U3244 (N_3244,N_732,N_991);
nand U3245 (N_3245,N_841,N_1407);
nand U3246 (N_3246,N_2914,N_2890);
xnor U3247 (N_3247,N_940,N_2026);
nand U3248 (N_3248,N_1220,N_743);
nor U3249 (N_3249,N_2230,N_1515);
nor U3250 (N_3250,N_1208,N_447);
and U3251 (N_3251,N_1359,N_2137);
nor U3252 (N_3252,N_2483,N_616);
nand U3253 (N_3253,N_548,N_2503);
nor U3254 (N_3254,N_1288,N_845);
nand U3255 (N_3255,N_1461,N_774);
nand U3256 (N_3256,N_2136,N_1842);
nand U3257 (N_3257,N_2820,N_296);
nand U3258 (N_3258,N_2464,N_844);
nor U3259 (N_3259,N_1786,N_1528);
nor U3260 (N_3260,N_137,N_2879);
and U3261 (N_3261,N_976,N_1254);
and U3262 (N_3262,N_2495,N_23);
or U3263 (N_3263,N_568,N_1038);
nor U3264 (N_3264,N_176,N_1346);
and U3265 (N_3265,N_1301,N_1759);
or U3266 (N_3266,N_2413,N_720);
and U3267 (N_3267,N_2344,N_239);
nor U3268 (N_3268,N_1588,N_2195);
nand U3269 (N_3269,N_2338,N_1607);
nand U3270 (N_3270,N_610,N_2208);
and U3271 (N_3271,N_2701,N_2293);
xor U3272 (N_3272,N_1358,N_2896);
or U3273 (N_3273,N_2650,N_2683);
nor U3274 (N_3274,N_729,N_1278);
or U3275 (N_3275,N_814,N_650);
nand U3276 (N_3276,N_2862,N_1626);
nand U3277 (N_3277,N_2821,N_2445);
and U3278 (N_3278,N_2506,N_2353);
nand U3279 (N_3279,N_849,N_2913);
nor U3280 (N_3280,N_839,N_2957);
nand U3281 (N_3281,N_2668,N_345);
or U3282 (N_3282,N_2039,N_513);
and U3283 (N_3283,N_2351,N_1848);
nand U3284 (N_3284,N_1172,N_476);
or U3285 (N_3285,N_1296,N_1415);
nand U3286 (N_3286,N_1578,N_2455);
and U3287 (N_3287,N_138,N_298);
nand U3288 (N_3288,N_1361,N_1957);
nor U3289 (N_3289,N_2408,N_2691);
or U3290 (N_3290,N_2644,N_1585);
or U3291 (N_3291,N_2533,N_1143);
and U3292 (N_3292,N_1264,N_1037);
or U3293 (N_3293,N_1726,N_2450);
nand U3294 (N_3294,N_246,N_407);
and U3295 (N_3295,N_2791,N_2795);
nor U3296 (N_3296,N_1689,N_909);
and U3297 (N_3297,N_649,N_2979);
and U3298 (N_3298,N_1117,N_708);
and U3299 (N_3299,N_2487,N_1452);
nor U3300 (N_3300,N_1093,N_2596);
nand U3301 (N_3301,N_427,N_2501);
or U3302 (N_3302,N_2154,N_2363);
nand U3303 (N_3303,N_1637,N_183);
or U3304 (N_3304,N_9,N_2201);
nor U3305 (N_3305,N_378,N_1994);
and U3306 (N_3306,N_2556,N_2009);
or U3307 (N_3307,N_1811,N_2725);
and U3308 (N_3308,N_133,N_2576);
and U3309 (N_3309,N_1231,N_2134);
and U3310 (N_3310,N_2689,N_1364);
nand U3311 (N_3311,N_1950,N_1243);
nand U3312 (N_3312,N_2401,N_596);
or U3313 (N_3313,N_2475,N_2970);
nor U3314 (N_3314,N_545,N_1819);
xor U3315 (N_3315,N_716,N_1224);
nor U3316 (N_3316,N_125,N_326);
nand U3317 (N_3317,N_749,N_1905);
or U3318 (N_3318,N_47,N_1675);
nor U3319 (N_3319,N_2435,N_462);
nor U3320 (N_3320,N_1179,N_735);
or U3321 (N_3321,N_423,N_2298);
nand U3322 (N_3322,N_1923,N_1555);
nor U3323 (N_3323,N_2528,N_132);
and U3324 (N_3324,N_2417,N_93);
or U3325 (N_3325,N_904,N_603);
nand U3326 (N_3326,N_2228,N_2433);
nor U3327 (N_3327,N_129,N_279);
or U3328 (N_3328,N_127,N_547);
nor U3329 (N_3329,N_2170,N_2547);
and U3330 (N_3330,N_64,N_352);
and U3331 (N_3331,N_1229,N_2003);
or U3332 (N_3332,N_343,N_164);
nor U3333 (N_3333,N_2532,N_2015);
nand U3334 (N_3334,N_1360,N_2785);
or U3335 (N_3335,N_728,N_982);
nand U3336 (N_3336,N_2493,N_350);
nand U3337 (N_3337,N_1777,N_1571);
nand U3338 (N_3338,N_2748,N_924);
nand U3339 (N_3339,N_2570,N_2865);
nor U3340 (N_3340,N_1855,N_2564);
xnor U3341 (N_3341,N_202,N_725);
and U3342 (N_3342,N_74,N_2394);
nand U3343 (N_3343,N_2055,N_161);
and U3344 (N_3344,N_1192,N_2006);
nor U3345 (N_3345,N_1822,N_2775);
nor U3346 (N_3346,N_2421,N_151);
nand U3347 (N_3347,N_82,N_439);
and U3348 (N_3348,N_645,N_2034);
nand U3349 (N_3349,N_2118,N_747);
nand U3350 (N_3350,N_460,N_1155);
or U3351 (N_3351,N_2648,N_2294);
and U3352 (N_3352,N_36,N_2446);
nand U3353 (N_3353,N_1843,N_1089);
nand U3354 (N_3354,N_2824,N_1791);
nor U3355 (N_3355,N_259,N_15);
nand U3356 (N_3356,N_1478,N_1132);
and U3357 (N_3357,N_2074,N_409);
nor U3358 (N_3358,N_1495,N_2620);
and U3359 (N_3359,N_1330,N_2735);
or U3360 (N_3360,N_191,N_1147);
and U3361 (N_3361,N_1316,N_2711);
nand U3362 (N_3362,N_1365,N_1070);
nand U3363 (N_3363,N_552,N_319);
nand U3364 (N_3364,N_1605,N_383);
nand U3365 (N_3365,N_1629,N_1701);
or U3366 (N_3366,N_2746,N_2759);
or U3367 (N_3367,N_617,N_2138);
xor U3368 (N_3368,N_1014,N_2660);
nor U3369 (N_3369,N_134,N_1792);
nor U3370 (N_3370,N_1173,N_374);
nor U3371 (N_3371,N_2325,N_805);
nand U3372 (N_3372,N_2002,N_1481);
nor U3373 (N_3373,N_2322,N_2341);
nand U3374 (N_3374,N_965,N_2816);
nor U3375 (N_3375,N_1801,N_2429);
and U3376 (N_3376,N_975,N_1785);
or U3377 (N_3377,N_2481,N_1042);
nand U3378 (N_3378,N_2810,N_2811);
nor U3379 (N_3379,N_1328,N_265);
and U3380 (N_3380,N_717,N_17);
and U3381 (N_3381,N_1741,N_2087);
or U3382 (N_3382,N_1740,N_2161);
nand U3383 (N_3383,N_2158,N_2472);
nand U3384 (N_3384,N_486,N_218);
nand U3385 (N_3385,N_254,N_802);
nor U3386 (N_3386,N_977,N_1712);
and U3387 (N_3387,N_2912,N_1284);
nor U3388 (N_3388,N_1329,N_1570);
or U3389 (N_3389,N_2014,N_1652);
nand U3390 (N_3390,N_1720,N_1942);
or U3391 (N_3391,N_171,N_1589);
or U3392 (N_3392,N_1849,N_2995);
nor U3393 (N_3393,N_1017,N_906);
or U3394 (N_3394,N_2839,N_21);
xnor U3395 (N_3395,N_2454,N_914);
and U3396 (N_3396,N_821,N_973);
and U3397 (N_3397,N_806,N_2788);
and U3398 (N_3398,N_2147,N_474);
and U3399 (N_3399,N_2699,N_182);
xor U3400 (N_3400,N_397,N_51);
and U3401 (N_3401,N_386,N_543);
and U3402 (N_3402,N_1279,N_2348);
or U3403 (N_3403,N_1403,N_358);
nor U3404 (N_3404,N_822,N_1317);
or U3405 (N_3405,N_1182,N_1579);
xor U3406 (N_3406,N_2587,N_1318);
nand U3407 (N_3407,N_166,N_188);
nand U3408 (N_3408,N_2541,N_30);
and U3409 (N_3409,N_2958,N_1806);
nand U3410 (N_3410,N_2732,N_2536);
and U3411 (N_3411,N_1930,N_284);
or U3412 (N_3412,N_937,N_2675);
nor U3413 (N_3413,N_2635,N_1178);
nand U3414 (N_3414,N_1004,N_2235);
and U3415 (N_3415,N_377,N_2772);
or U3416 (N_3416,N_2961,N_465);
or U3417 (N_3417,N_1723,N_67);
or U3418 (N_3418,N_219,N_1617);
nand U3419 (N_3419,N_1065,N_1459);
nor U3420 (N_3420,N_2966,N_2061);
nand U3421 (N_3421,N_2465,N_1225);
nor U3422 (N_3422,N_995,N_301);
and U3423 (N_3423,N_2793,N_2743);
nand U3424 (N_3424,N_809,N_1861);
and U3425 (N_3425,N_60,N_2632);
nor U3426 (N_3426,N_1141,N_2071);
and U3427 (N_3427,N_938,N_194);
nand U3428 (N_3428,N_1493,N_564);
nor U3429 (N_3429,N_121,N_922);
nand U3430 (N_3430,N_208,N_387);
nand U3431 (N_3431,N_291,N_339);
and U3432 (N_3432,N_207,N_1214);
nor U3433 (N_3433,N_511,N_1352);
nor U3434 (N_3434,N_1880,N_285);
nand U3435 (N_3435,N_1120,N_955);
nor U3436 (N_3436,N_1780,N_371);
nor U3437 (N_3437,N_1036,N_2673);
nor U3438 (N_3438,N_2767,N_2406);
or U3439 (N_3439,N_1369,N_533);
nor U3440 (N_3440,N_1184,N_1015);
and U3441 (N_3441,N_1107,N_1012);
and U3442 (N_3442,N_1933,N_1985);
nor U3443 (N_3443,N_466,N_1755);
nand U3444 (N_3444,N_103,N_1575);
and U3445 (N_3445,N_823,N_1773);
nor U3446 (N_3446,N_158,N_562);
nor U3447 (N_3447,N_949,N_709);
nor U3448 (N_3448,N_1217,N_305);
nor U3449 (N_3449,N_1142,N_2203);
nor U3450 (N_3450,N_1530,N_573);
nand U3451 (N_3451,N_1291,N_1809);
nand U3452 (N_3452,N_2,N_2120);
and U3453 (N_3453,N_450,N_2320);
nand U3454 (N_3454,N_1261,N_592);
xor U3455 (N_3455,N_2670,N_2146);
or U3456 (N_3456,N_1476,N_302);
nor U3457 (N_3457,N_2942,N_367);
or U3458 (N_3458,N_2612,N_2717);
and U3459 (N_3459,N_327,N_677);
and U3460 (N_3460,N_341,N_205);
nand U3461 (N_3461,N_1251,N_1916);
nor U3462 (N_3462,N_96,N_1152);
or U3463 (N_3463,N_2686,N_1331);
nand U3464 (N_3464,N_1554,N_2245);
or U3465 (N_3465,N_2169,N_1517);
and U3466 (N_3466,N_2214,N_40);
or U3467 (N_3467,N_69,N_2592);
nor U3468 (N_3468,N_1003,N_2994);
and U3469 (N_3469,N_606,N_2864);
and U3470 (N_3470,N_2000,N_227);
nand U3471 (N_3471,N_506,N_106);
nand U3472 (N_3472,N_1829,N_1936);
or U3473 (N_3473,N_1841,N_2549);
nor U3474 (N_3474,N_2678,N_1533);
and U3475 (N_3475,N_2148,N_1297);
nand U3476 (N_3476,N_2507,N_344);
nor U3477 (N_3477,N_214,N_2359);
nand U3478 (N_3478,N_510,N_492);
or U3479 (N_3479,N_1349,N_123);
and U3480 (N_3480,N_2282,N_1490);
xnor U3481 (N_3481,N_2274,N_2967);
nor U3482 (N_3482,N_985,N_342);
nand U3483 (N_3483,N_2405,N_2807);
nand U3484 (N_3484,N_2937,N_790);
and U3485 (N_3485,N_275,N_2990);
nor U3486 (N_3486,N_1456,N_2769);
nand U3487 (N_3487,N_2381,N_1864);
nor U3488 (N_3488,N_1338,N_2964);
nor U3489 (N_3489,N_340,N_1870);
nor U3490 (N_3490,N_1026,N_2437);
nand U3491 (N_3491,N_2126,N_1223);
or U3492 (N_3492,N_2223,N_2229);
and U3493 (N_3493,N_800,N_702);
or U3494 (N_3494,N_2403,N_2347);
and U3495 (N_3495,N_2524,N_1639);
or U3496 (N_3496,N_2358,N_1433);
and U3497 (N_3497,N_789,N_2871);
or U3498 (N_3498,N_856,N_2349);
and U3499 (N_3499,N_1397,N_1194);
and U3500 (N_3500,N_1926,N_2724);
or U3501 (N_3501,N_2669,N_2892);
nand U3502 (N_3502,N_2287,N_2264);
nand U3503 (N_3503,N_1692,N_1350);
and U3504 (N_3504,N_416,N_576);
or U3505 (N_3505,N_2645,N_1882);
or U3506 (N_3506,N_585,N_557);
nand U3507 (N_3507,N_117,N_2215);
and U3508 (N_3508,N_2730,N_1386);
or U3509 (N_3509,N_79,N_1910);
or U3510 (N_3510,N_1449,N_622);
xnor U3511 (N_3511,N_1315,N_604);
nand U3512 (N_3512,N_594,N_2088);
or U3513 (N_3513,N_641,N_1354);
and U3514 (N_3514,N_2496,N_2277);
nand U3515 (N_3515,N_820,N_2248);
or U3516 (N_3516,N_2550,N_1246);
and U3517 (N_3517,N_323,N_2324);
or U3518 (N_3518,N_1781,N_2665);
nand U3519 (N_3519,N_784,N_2001);
nor U3520 (N_3520,N_1644,N_1440);
or U3521 (N_3521,N_2940,N_1455);
nor U3522 (N_3522,N_614,N_2057);
or U3523 (N_3523,N_1623,N_2336);
nor U3524 (N_3524,N_1314,N_1100);
and U3525 (N_3525,N_1442,N_966);
nor U3526 (N_3526,N_908,N_1518);
nor U3527 (N_3527,N_514,N_2923);
or U3528 (N_3528,N_2012,N_2687);
nor U3529 (N_3529,N_274,N_542);
nor U3530 (N_3530,N_61,N_1052);
or U3531 (N_3531,N_1043,N_1744);
xnor U3532 (N_3532,N_1839,N_42);
nor U3533 (N_3533,N_2886,N_1788);
or U3534 (N_3534,N_1280,N_2396);
and U3535 (N_3535,N_1090,N_2438);
and U3536 (N_3536,N_1753,N_1634);
and U3537 (N_3537,N_307,N_640);
and U3538 (N_3538,N_2051,N_395);
nor U3539 (N_3539,N_1591,N_2373);
nand U3540 (N_3540,N_2834,N_1130);
and U3541 (N_3541,N_1303,N_186);
and U3542 (N_3542,N_2106,N_890);
nand U3543 (N_3543,N_560,N_1380);
nor U3544 (N_3544,N_282,N_457);
or U3545 (N_3545,N_2591,N_512);
nand U3546 (N_3546,N_1488,N_318);
or U3547 (N_3547,N_401,N_236);
and U3548 (N_3548,N_2060,N_2572);
nand U3549 (N_3549,N_2915,N_530);
nand U3550 (N_3550,N_2884,N_2720);
nor U3551 (N_3551,N_2090,N_2656);
or U3552 (N_3552,N_1411,N_2448);
nand U3553 (N_3553,N_1593,N_892);
nand U3554 (N_3554,N_2385,N_1616);
and U3555 (N_3555,N_1865,N_584);
nand U3556 (N_3556,N_741,N_2918);
or U3557 (N_3557,N_448,N_1430);
or U3558 (N_3558,N_2712,N_2604);
nor U3559 (N_3559,N_2070,N_116);
and U3560 (N_3560,N_177,N_2257);
nor U3561 (N_3561,N_1859,N_32);
or U3562 (N_3562,N_497,N_2124);
nor U3563 (N_3563,N_1068,N_459);
or U3564 (N_3564,N_76,N_2011);
and U3565 (N_3565,N_2739,N_2023);
or U3566 (N_3566,N_2789,N_2992);
or U3567 (N_3567,N_2598,N_1479);
nor U3568 (N_3568,N_1975,N_245);
and U3569 (N_3569,N_83,N_1728);
nand U3570 (N_3570,N_1307,N_1457);
nor U3571 (N_3571,N_1486,N_310);
nand U3572 (N_3572,N_242,N_687);
or U3573 (N_3573,N_896,N_567);
nor U3574 (N_3574,N_2694,N_571);
or U3575 (N_3575,N_324,N_1599);
and U3576 (N_3576,N_255,N_1808);
and U3577 (N_3577,N_2577,N_2943);
or U3578 (N_3578,N_1233,N_2489);
and U3579 (N_3579,N_1645,N_2017);
or U3580 (N_3580,N_1595,N_110);
nand U3581 (N_3581,N_636,N_2069);
nor U3582 (N_3582,N_2036,N_2093);
and U3583 (N_3583,N_1230,N_2224);
or U3584 (N_3584,N_78,N_1655);
nand U3585 (N_3585,N_2383,N_2151);
and U3586 (N_3586,N_2281,N_470);
nor U3587 (N_3587,N_2243,N_313);
nand U3588 (N_3588,N_1531,N_2649);
or U3589 (N_3589,N_2250,N_316);
nand U3590 (N_3590,N_740,N_881);
nor U3591 (N_3591,N_115,N_2150);
nor U3592 (N_3592,N_1600,N_2608);
or U3593 (N_3593,N_2210,N_1371);
or U3594 (N_3594,N_1127,N_1055);
or U3595 (N_3595,N_2741,N_974);
nand U3596 (N_3596,N_1323,N_1608);
nor U3597 (N_3597,N_2143,N_1348);
or U3598 (N_3598,N_1271,N_722);
nand U3599 (N_3599,N_2252,N_2399);
xnor U3600 (N_3600,N_648,N_1633);
and U3601 (N_3601,N_1894,N_727);
nor U3602 (N_3602,N_502,N_1572);
or U3603 (N_3603,N_2078,N_1256);
and U3604 (N_3604,N_898,N_2661);
and U3605 (N_3605,N_1534,N_1965);
or U3606 (N_3606,N_299,N_834);
or U3607 (N_3607,N_1768,N_2333);
xor U3608 (N_3608,N_2110,N_1886);
and U3609 (N_3609,N_883,N_1219);
or U3610 (N_3610,N_1384,N_2367);
and U3611 (N_3611,N_612,N_1636);
nand U3612 (N_3612,N_704,N_55);
nor U3613 (N_3613,N_1874,N_425);
and U3614 (N_3614,N_1679,N_2904);
or U3615 (N_3615,N_835,N_2246);
nand U3616 (N_3616,N_689,N_2688);
or U3617 (N_3617,N_1083,N_195);
nand U3618 (N_3618,N_723,N_2798);
nand U3619 (N_3619,N_2786,N_782);
nand U3620 (N_3620,N_665,N_2318);
or U3621 (N_3621,N_1087,N_317);
or U3622 (N_3622,N_2831,N_2254);
or U3623 (N_3623,N_1059,N_2615);
and U3624 (N_3624,N_1913,N_444);
nor U3625 (N_3625,N_936,N_810);
and U3626 (N_3626,N_1941,N_2362);
nor U3627 (N_3627,N_1559,N_2790);
and U3628 (N_3628,N_320,N_791);
and U3629 (N_3629,N_2568,N_1867);
nor U3630 (N_3630,N_1453,N_2261);
nand U3631 (N_3631,N_2273,N_1618);
nor U3632 (N_3632,N_1362,N_2005);
and U3633 (N_3633,N_767,N_2272);
or U3634 (N_3634,N_2941,N_2621);
nand U3635 (N_3635,N_2211,N_921);
and U3636 (N_3636,N_403,N_1820);
and U3637 (N_3637,N_1114,N_1963);
or U3638 (N_3638,N_2016,N_2624);
nand U3639 (N_3639,N_672,N_2356);
or U3640 (N_3640,N_2545,N_402);
nand U3641 (N_3641,N_1681,N_1574);
nor U3642 (N_3642,N_1206,N_1011);
and U3643 (N_3643,N_1991,N_2700);
or U3644 (N_3644,N_2386,N_1417);
nand U3645 (N_3645,N_29,N_488);
nand U3646 (N_3646,N_333,N_754);
or U3647 (N_3647,N_2766,N_2895);
xnor U3648 (N_3648,N_1775,N_961);
nand U3649 (N_3649,N_998,N_666);
and U3650 (N_3650,N_2412,N_2030);
or U3651 (N_3651,N_394,N_1205);
xnor U3652 (N_3652,N_2468,N_1094);
and U3653 (N_3653,N_1547,N_349);
nor U3654 (N_3654,N_1821,N_290);
nand U3655 (N_3655,N_2565,N_2963);
and U3656 (N_3656,N_1441,N_2832);
nand U3657 (N_3657,N_2312,N_1624);
nor U3658 (N_3658,N_803,N_926);
nand U3659 (N_3659,N_2737,N_113);
or U3660 (N_3660,N_1934,N_1857);
or U3661 (N_3661,N_1548,N_157);
nand U3662 (N_3662,N_2664,N_905);
nor U3663 (N_3663,N_2551,N_952);
and U3664 (N_3664,N_1981,N_1538);
or U3665 (N_3665,N_1714,N_2610);
nor U3666 (N_3666,N_1427,N_1642);
or U3667 (N_3667,N_338,N_1845);
nor U3668 (N_3668,N_2781,N_496);
and U3669 (N_3669,N_884,N_1253);
and U3670 (N_3670,N_836,N_1680);
nand U3671 (N_3671,N_1660,N_2112);
or U3672 (N_3672,N_2019,N_2082);
or U3673 (N_3673,N_2114,N_1171);
or U3674 (N_3674,N_1398,N_278);
nand U3675 (N_3675,N_2721,N_84);
nor U3676 (N_3676,N_489,N_2909);
and U3677 (N_3677,N_619,N_1151);
or U3678 (N_3678,N_1852,N_1496);
or U3679 (N_3679,N_694,N_2740);
nand U3680 (N_3680,N_1077,N_1858);
nand U3681 (N_3681,N_1204,N_2331);
and U3682 (N_3682,N_1031,N_990);
nand U3683 (N_3683,N_1914,N_48);
and U3684 (N_3684,N_796,N_1631);
and U3685 (N_3685,N_580,N_565);
xnor U3686 (N_3686,N_876,N_314);
nor U3687 (N_3687,N_1366,N_2052);
nor U3688 (N_3688,N_2262,N_621);
and U3689 (N_3689,N_2897,N_1267);
nand U3690 (N_3690,N_2213,N_2600);
or U3691 (N_3691,N_589,N_2860);
nor U3692 (N_3692,N_1071,N_59);
or U3693 (N_3693,N_2075,N_838);
nor U3694 (N_3694,N_2848,N_376);
nand U3695 (N_3695,N_2152,N_1683);
and U3696 (N_3696,N_2733,N_2558);
and U3697 (N_3697,N_712,N_833);
nor U3698 (N_3698,N_2802,N_1736);
and U3699 (N_3699,N_772,N_52);
and U3700 (N_3700,N_1832,N_1106);
or U3701 (N_3701,N_2323,N_1125);
or U3702 (N_3702,N_44,N_2066);
and U3703 (N_3703,N_1529,N_1439);
or U3704 (N_3704,N_868,N_1272);
nand U3705 (N_3705,N_216,N_558);
nor U3706 (N_3706,N_1025,N_1210);
nand U3707 (N_3707,N_2975,N_1222);
or U3708 (N_3708,N_605,N_671);
or U3709 (N_3709,N_1581,N_2554);
or U3710 (N_3710,N_2823,N_885);
or U3711 (N_3711,N_270,N_1067);
or U3712 (N_3712,N_2332,N_1102);
nor U3713 (N_3713,N_436,N_273);
nor U3714 (N_3714,N_294,N_72);
nand U3715 (N_3715,N_644,N_2007);
nand U3716 (N_3716,N_1408,N_2513);
xnor U3717 (N_3717,N_507,N_2954);
or U3718 (N_3718,N_1860,N_87);
and U3719 (N_3719,N_2236,N_2960);
or U3720 (N_3720,N_2657,N_863);
or U3721 (N_3721,N_1945,N_500);
or U3722 (N_3722,N_2729,N_2708);
and U3723 (N_3723,N_1772,N_1469);
xnor U3724 (N_3724,N_389,N_220);
and U3725 (N_3725,N_2259,N_613);
nor U3726 (N_3726,N_77,N_901);
nor U3727 (N_3727,N_1032,N_2080);
nand U3728 (N_3728,N_1750,N_1019);
or U3729 (N_3729,N_1676,N_1851);
xnor U3730 (N_3730,N_1543,N_2567);
or U3731 (N_3731,N_935,N_1149);
nand U3732 (N_3732,N_818,N_1504);
and U3733 (N_3733,N_2305,N_866);
or U3734 (N_3734,N_2716,N_2826);
or U3735 (N_3735,N_2681,N_670);
nand U3736 (N_3736,N_2326,N_1996);
nor U3737 (N_3737,N_390,N_1900);
xnor U3738 (N_3738,N_1190,N_1162);
nor U3739 (N_3739,N_1730,N_1485);
nor U3740 (N_3740,N_2499,N_22);
and U3741 (N_3741,N_2337,N_739);
or U3742 (N_3742,N_70,N_705);
nor U3743 (N_3743,N_600,N_1321);
or U3744 (N_3744,N_1622,N_520);
nor U3745 (N_3745,N_1342,N_2378);
nor U3746 (N_3746,N_2117,N_857);
nand U3747 (N_3747,N_591,N_1946);
and U3748 (N_3748,N_2492,N_551);
nor U3749 (N_3749,N_962,N_1976);
or U3750 (N_3750,N_2284,N_2217);
or U3751 (N_3751,N_1295,N_730);
nand U3752 (N_3752,N_2602,N_2840);
and U3753 (N_3753,N_1627,N_1719);
or U3754 (N_3754,N_370,N_1630);
and U3755 (N_3755,N_28,N_2407);
nor U3756 (N_3756,N_574,N_2470);
nand U3757 (N_3757,N_5,N_104);
nand U3758 (N_3758,N_1050,N_2168);
or U3759 (N_3759,N_1300,N_209);
or U3760 (N_3760,N_2062,N_1763);
nand U3761 (N_3761,N_1161,N_240);
and U3762 (N_3762,N_1558,N_1995);
or U3763 (N_3763,N_1868,N_1124);
and U3764 (N_3764,N_2467,N_2197);
or U3765 (N_3765,N_1468,N_2300);
nor U3766 (N_3766,N_950,N_2285);
and U3767 (N_3767,N_1540,N_2428);
nand U3768 (N_3768,N_1292,N_1743);
nor U3769 (N_3769,N_1961,N_2703);
nand U3770 (N_3770,N_1587,N_1847);
nand U3771 (N_3771,N_2159,N_1392);
and U3772 (N_3772,N_907,N_1562);
or U3773 (N_3773,N_787,N_253);
and U3774 (N_3774,N_1138,N_2763);
and U3775 (N_3775,N_2822,N_2637);
nand U3776 (N_3776,N_2079,N_2578);
or U3777 (N_3777,N_417,N_1830);
or U3778 (N_3778,N_2976,N_1351);
and U3779 (N_3779,N_2508,N_1584);
xnor U3780 (N_3780,N_1446,N_2212);
or U3781 (N_3781,N_2727,N_2350);
xnor U3782 (N_3782,N_1754,N_2936);
and U3783 (N_3783,N_969,N_2969);
xor U3784 (N_3784,N_2198,N_2444);
or U3785 (N_3785,N_108,N_726);
or U3786 (N_3786,N_1119,N_1673);
nand U3787 (N_3787,N_1598,N_2441);
nand U3788 (N_3788,N_508,N_1716);
nor U3789 (N_3789,N_1166,N_234);
or U3790 (N_3790,N_590,N_131);
nand U3791 (N_3791,N_1146,N_2502);
nand U3792 (N_3792,N_1747,N_1871);
xnor U3793 (N_3793,N_1465,N_1060);
nor U3794 (N_3794,N_2286,N_2707);
or U3795 (N_3795,N_742,N_430);
nor U3796 (N_3796,N_1188,N_2965);
or U3797 (N_3797,N_2402,N_1552);
nand U3798 (N_3798,N_2374,N_1244);
and U3799 (N_3799,N_2171,N_2827);
nand U3800 (N_3800,N_1978,N_1156);
nand U3801 (N_3801,N_1470,N_256);
and U3802 (N_3802,N_452,N_2073);
and U3803 (N_3803,N_1542,N_2647);
and U3804 (N_3804,N_1641,N_615);
and U3805 (N_3805,N_2497,N_850);
or U3806 (N_3806,N_2973,N_2156);
nor U3807 (N_3807,N_2770,N_366);
nand U3808 (N_3808,N_653,N_819);
nor U3809 (N_3809,N_2606,N_1817);
nor U3810 (N_3810,N_1862,N_1298);
nand U3811 (N_3811,N_2692,N_2233);
nor U3812 (N_3812,N_2216,N_1932);
and U3813 (N_3813,N_68,N_1909);
and U3814 (N_3814,N_569,N_795);
or U3815 (N_3815,N_1334,N_393);
and U3816 (N_3816,N_786,N_2538);
nor U3817 (N_3817,N_2586,N_928);
nand U3818 (N_3818,N_1273,N_2289);
nand U3819 (N_3819,N_1769,N_37);
or U3820 (N_3820,N_2425,N_1749);
and U3821 (N_3821,N_2498,N_2951);
and U3822 (N_3822,N_2050,N_765);
nand U3823 (N_3823,N_1539,N_812);
nor U3824 (N_3824,N_38,N_1854);
nor U3825 (N_3825,N_2561,N_1752);
nand U3826 (N_3826,N_1814,N_2360);
and U3827 (N_3827,N_24,N_2696);
or U3828 (N_3828,N_2477,N_1088);
or U3829 (N_3829,N_1959,N_162);
or U3830 (N_3830,N_2165,N_2662);
and U3831 (N_3831,N_607,N_1103);
and U3832 (N_3832,N_1590,N_1066);
nand U3833 (N_3833,N_1409,N_276);
and U3834 (N_3834,N_1180,N_1174);
and U3835 (N_3835,N_446,N_3);
and U3836 (N_3836,N_2837,N_1925);
nand U3837 (N_3837,N_2622,N_618);
or U3838 (N_3838,N_2010,N_2205);
nand U3839 (N_3839,N_165,N_2291);
and U3840 (N_3840,N_524,N_2099);
and U3841 (N_3841,N_1553,N_2307);
nand U3842 (N_3842,N_73,N_2045);
or U3843 (N_3843,N_1027,N_1475);
or U3844 (N_3844,N_2044,N_1657);
xor U3845 (N_3845,N_2361,N_1573);
nor U3846 (N_3846,N_658,N_1774);
and U3847 (N_3847,N_1799,N_2634);
or U3848 (N_3848,N_2546,N_1968);
or U3849 (N_3849,N_2474,N_2905);
nand U3850 (N_3850,N_1834,N_369);
nor U3851 (N_3851,N_1974,N_2133);
nor U3852 (N_3852,N_2579,N_173);
or U3853 (N_3853,N_485,N_2125);
nand U3854 (N_3854,N_900,N_2267);
nor U3855 (N_3855,N_2933,N_155);
nand U3856 (N_3856,N_2575,N_595);
nand U3857 (N_3857,N_1844,N_1643);
xor U3858 (N_3858,N_570,N_1535);
or U3859 (N_3859,N_1878,N_920);
or U3860 (N_3860,N_325,N_523);
or U3861 (N_3861,N_1121,N_624);
nor U3862 (N_3862,N_2525,N_2921);
nand U3863 (N_3863,N_1432,N_1045);
nor U3864 (N_3864,N_295,N_435);
nor U3865 (N_3865,N_2968,N_1104);
or U3866 (N_3866,N_1734,N_458);
xnor U3867 (N_3867,N_375,N_947);
or U3868 (N_3868,N_25,N_2185);
and U3869 (N_3869,N_1145,N_1708);
or U3870 (N_3870,N_943,N_2771);
and U3871 (N_3871,N_2237,N_1447);
nor U3872 (N_3872,N_2935,N_2127);
or U3873 (N_3873,N_2311,N_813);
or U3874 (N_3874,N_2784,N_2423);
nand U3875 (N_3875,N_960,N_2135);
and U3876 (N_3876,N_1480,N_26);
nand U3877 (N_3877,N_41,N_363);
and U3878 (N_3878,N_1193,N_505);
nand U3879 (N_3879,N_837,N_2265);
nand U3880 (N_3880,N_2911,N_1816);
or U3881 (N_3881,N_579,N_2626);
or U3882 (N_3882,N_1506,N_2218);
nor U3883 (N_3883,N_1333,N_1473);
or U3884 (N_3884,N_2705,N_1688);
nor U3885 (N_3885,N_1029,N_2164);
and U3886 (N_3886,N_213,N_1454);
nor U3887 (N_3887,N_2571,N_412);
and U3888 (N_3888,N_2697,N_1232);
and U3889 (N_3889,N_2129,N_1268);
nor U3890 (N_3890,N_2815,N_1423);
or U3891 (N_3891,N_628,N_2955);
and U3892 (N_3892,N_2858,N_414);
nor U3893 (N_3893,N_18,N_794);
or U3894 (N_3894,N_2916,N_53);
nand U3895 (N_3895,N_2369,N_2985);
or U3896 (N_3896,N_2856,N_1560);
nor U3897 (N_3897,N_2183,N_1802);
or U3898 (N_3898,N_1341,N_286);
and U3899 (N_3899,N_2751,N_1766);
or U3900 (N_3900,N_381,N_2366);
or U3901 (N_3901,N_848,N_2812);
or U3902 (N_3902,N_238,N_1290);
or U3903 (N_3903,N_807,N_1270);
or U3904 (N_3904,N_1347,N_2859);
and U3905 (N_3905,N_1393,N_65);
nand U3906 (N_3906,N_2715,N_360);
nand U3907 (N_3907,N_1937,N_550);
nand U3908 (N_3908,N_1056,N_2633);
nand U3909 (N_3909,N_306,N_498);
nor U3910 (N_3910,N_1313,N_2534);
or U3911 (N_3911,N_2625,N_2768);
nor U3912 (N_3912,N_1311,N_478);
and U3913 (N_3913,N_2419,N_2540);
nand U3914 (N_3914,N_2486,N_731);
nand U3915 (N_3915,N_2033,N_553);
xnor U3916 (N_3916,N_532,N_2232);
and U3917 (N_3917,N_2038,N_2877);
and U3918 (N_3918,N_2175,N_503);
and U3919 (N_3919,N_2340,N_1489);
nand U3920 (N_3920,N_1276,N_66);
or U3921 (N_3921,N_1944,N_2825);
or U3922 (N_3922,N_120,N_1073);
or U3923 (N_3923,N_2398,N_957);
nor U3924 (N_3924,N_145,N_1135);
and U3925 (N_3925,N_1153,N_1650);
nor U3926 (N_3926,N_410,N_1154);
nand U3927 (N_3927,N_1765,N_1694);
and U3928 (N_3928,N_1653,N_1988);
nor U3929 (N_3929,N_679,N_1638);
nor U3930 (N_3930,N_2505,N_2959);
or U3931 (N_3931,N_405,N_2597);
and U3932 (N_3932,N_2607,N_2240);
or U3933 (N_3933,N_354,N_1363);
and U3934 (N_3934,N_1126,N_1952);
nand U3935 (N_3935,N_1706,N_100);
or U3936 (N_3936,N_1131,N_2663);
nand U3937 (N_3937,N_748,N_2049);
and U3938 (N_3938,N_2339,N_1218);
or U3939 (N_3939,N_2855,N_396);
nor U3940 (N_3940,N_1158,N_1105);
and U3941 (N_3941,N_2092,N_1434);
nor U3942 (N_3942,N_181,N_2458);
or U3943 (N_3943,N_1293,N_329);
or U3944 (N_3944,N_2630,N_1902);
or U3945 (N_3945,N_660,N_2116);
or U3946 (N_3946,N_1746,N_2646);
nor U3947 (N_3947,N_2996,N_509);
nand U3948 (N_3948,N_1076,N_903);
and U3949 (N_3949,N_2535,N_348);
nand U3950 (N_3950,N_1237,N_2295);
nor U3951 (N_3951,N_34,N_724);
nand U3952 (N_3952,N_1081,N_2928);
nor U3953 (N_3953,N_2149,N_2354);
or U3954 (N_3954,N_652,N_455);
nor U3955 (N_3955,N_357,N_243);
nand U3956 (N_3956,N_637,N_1810);
or U3957 (N_3957,N_1075,N_1049);
nor U3958 (N_3958,N_1550,N_2131);
or U3959 (N_3959,N_2845,N_2938);
nor U3960 (N_3960,N_440,N_1464);
and U3961 (N_3961,N_690,N_775);
nor U3962 (N_3962,N_634,N_1718);
nor U3963 (N_3963,N_80,N_1710);
nor U3964 (N_3964,N_1523,N_283);
and U3965 (N_3965,N_1596,N_361);
nor U3966 (N_3966,N_2874,N_987);
and U3967 (N_3967,N_1879,N_2638);
and U3968 (N_3968,N_130,N_1873);
nand U3969 (N_3969,N_1257,N_2993);
or U3970 (N_3970,N_773,N_2084);
and U3971 (N_3971,N_964,N_331);
nand U3972 (N_3972,N_983,N_1695);
or U3973 (N_3973,N_432,N_746);
nor U3974 (N_3974,N_1320,N_472);
or U3975 (N_3975,N_1970,N_2631);
or U3976 (N_3976,N_1969,N_2543);
or U3977 (N_3977,N_2491,N_1611);
or U3978 (N_3978,N_398,N_95);
xnor U3979 (N_3979,N_50,N_893);
nand U3980 (N_3980,N_1748,N_1418);
nand U3981 (N_3981,N_635,N_170);
or U3982 (N_3982,N_1482,N_2846);
or U3983 (N_3983,N_1010,N_1445);
and U3984 (N_3984,N_6,N_2883);
and U3985 (N_3985,N_1389,N_2107);
and U3986 (N_3986,N_146,N_1001);
nand U3987 (N_3987,N_656,N_1426);
nand U3988 (N_3988,N_1514,N_879);
nand U3989 (N_3989,N_149,N_1665);
and U3990 (N_3990,N_281,N_1108);
and U3991 (N_3991,N_2764,N_139);
and U3992 (N_3992,N_676,N_2843);
nor U3993 (N_3993,N_1477,N_2907);
or U3994 (N_3994,N_461,N_1429);
and U3995 (N_3995,N_1248,N_289);
nand U3996 (N_3996,N_1940,N_768);
and U3997 (N_3997,N_1379,N_2544);
xor U3998 (N_3998,N_1484,N_878);
or U3999 (N_3999,N_1196,N_2482);
nand U4000 (N_4000,N_1760,N_2539);
nor U4001 (N_4001,N_933,N_347);
and U4002 (N_4002,N_2345,N_2557);
nand U4003 (N_4003,N_877,N_516);
nor U4004 (N_4004,N_1972,N_678);
nand U4005 (N_4005,N_14,N_2518);
nor U4006 (N_4006,N_2202,N_1139);
or U4007 (N_4007,N_2379,N_1510);
or U4008 (N_4008,N_1895,N_2783);
nand U4009 (N_4009,N_422,N_262);
nor U4010 (N_4010,N_63,N_2900);
and U4011 (N_4011,N_257,N_1030);
and U4012 (N_4012,N_2588,N_1209);
nand U4013 (N_4013,N_2653,N_293);
nand U4014 (N_4014,N_481,N_1919);
nand U4015 (N_4015,N_1181,N_1109);
nand U4016 (N_4016,N_388,N_1327);
or U4017 (N_4017,N_2244,N_1502);
xor U4018 (N_4018,N_1797,N_1958);
and U4019 (N_4019,N_2053,N_873);
or U4020 (N_4020,N_1265,N_880);
or U4021 (N_4021,N_1567,N_2850);
and U4022 (N_4022,N_2728,N_2056);
nor U4023 (N_4023,N_1410,N_1928);
or U4024 (N_4024,N_1866,N_2803);
and U4025 (N_4025,N_1400,N_1887);
nor U4026 (N_4026,N_2020,N_1198);
nor U4027 (N_4027,N_978,N_152);
nand U4028 (N_4028,N_544,N_1696);
and U4029 (N_4029,N_1000,N_1287);
and U4030 (N_4030,N_1137,N_1982);
nor U4031 (N_4031,N_1235,N_206);
nand U4032 (N_4032,N_1424,N_1856);
or U4033 (N_4033,N_1668,N_126);
nor U4034 (N_4034,N_1837,N_2599);
and U4035 (N_4035,N_2829,N_315);
nand U4036 (N_4036,N_2299,N_1207);
nand U4037 (N_4037,N_1168,N_2752);
nor U4038 (N_4038,N_1058,N_2805);
and U4039 (N_4039,N_1671,N_2256);
nor U4040 (N_4040,N_861,N_515);
or U4041 (N_4041,N_954,N_97);
or U4042 (N_4042,N_1123,N_529);
nor U4043 (N_4043,N_1023,N_2226);
nand U4044 (N_4044,N_1987,N_875);
or U4045 (N_4045,N_89,N_1635);
and U4046 (N_4046,N_1960,N_537);
nor U4047 (N_4047,N_1099,N_2199);
and U4048 (N_4048,N_2510,N_902);
or U4049 (N_4049,N_2667,N_1252);
and U4050 (N_4050,N_1953,N_248);
nor U4051 (N_4051,N_368,N_1016);
and U4052 (N_4052,N_1165,N_413);
nand U4053 (N_4053,N_309,N_199);
and U4054 (N_4054,N_1967,N_582);
or U4055 (N_4055,N_2719,N_631);
xor U4056 (N_4056,N_1336,N_1935);
nor U4057 (N_4057,N_1007,N_1202);
nand U4058 (N_4058,N_464,N_2479);
or U4059 (N_4059,N_958,N_1458);
xor U4060 (N_4060,N_1722,N_1013);
or U4061 (N_4061,N_2814,N_2377);
xor U4062 (N_4062,N_1685,N_1129);
nand U4063 (N_4063,N_882,N_1904);
and U4064 (N_4064,N_1727,N_94);
nand U4065 (N_4065,N_2947,N_400);
or U4066 (N_4066,N_473,N_659);
or U4067 (N_4067,N_654,N_1920);
nand U4068 (N_4068,N_2643,N_431);
or U4069 (N_4069,N_2411,N_111);
nor U4070 (N_4070,N_2440,N_1762);
nor U4071 (N_4071,N_912,N_2901);
nor U4072 (N_4072,N_2278,N_19);
nor U4073 (N_4073,N_1947,N_204);
or U4074 (N_4074,N_1658,N_1711);
or U4075 (N_4075,N_647,N_2779);
or U4076 (N_4076,N_1784,N_1344);
or U4077 (N_4077,N_1034,N_587);
and U4078 (N_4078,N_1133,N_696);
and U4079 (N_4079,N_2241,N_2393);
nor U4080 (N_4080,N_2552,N_45);
or U4081 (N_4081,N_1283,N_2457);
and U4082 (N_4082,N_2392,N_2548);
nor U4083 (N_4083,N_1375,N_2595);
nand U4084 (N_4084,N_2365,N_753);
and U4085 (N_4085,N_2024,N_776);
nand U4086 (N_4086,N_2659,N_266);
or U4087 (N_4087,N_1024,N_2722);
nor U4088 (N_4088,N_2847,N_1827);
nand U4089 (N_4089,N_2040,N_1374);
or U4090 (N_4090,N_2562,N_2680);
or U4091 (N_4091,N_1881,N_429);
or U4092 (N_4092,N_2983,N_159);
and U4093 (N_4093,N_2526,N_442);
and U4094 (N_4094,N_2238,N_752);
nor U4095 (N_4095,N_2885,N_1929);
nor U4096 (N_4096,N_2609,N_2089);
or U4097 (N_4097,N_1604,N_539);
and U4098 (N_4098,N_2108,N_1021);
or U4099 (N_4099,N_1885,N_1551);
nor U4100 (N_4100,N_1824,N_798);
nor U4101 (N_4101,N_714,N_241);
nor U4102 (N_4102,N_91,N_945);
and U4103 (N_4103,N_2851,N_54);
and U4104 (N_4104,N_620,N_699);
nand U4105 (N_4105,N_2749,N_1705);
nand U4106 (N_4106,N_2742,N_304);
and U4107 (N_4107,N_2917,N_913);
nand U4108 (N_4108,N_1503,N_1815);
nor U4109 (N_4109,N_2157,N_2352);
and U4110 (N_4110,N_2614,N_1884);
or U4111 (N_4111,N_583,N_1949);
nand U4112 (N_4112,N_2388,N_1324);
or U4113 (N_4113,N_1850,N_1373);
and U4114 (N_4114,N_2488,N_646);
and U4115 (N_4115,N_783,N_2801);
nand U4116 (N_4116,N_2553,N_1678);
and U4117 (N_4117,N_31,N_2792);
nand U4118 (N_4118,N_1697,N_2346);
and U4119 (N_4119,N_559,N_691);
and U4120 (N_4120,N_471,N_2654);
or U4121 (N_4121,N_1047,N_988);
nand U4122 (N_4122,N_2515,N_929);
nand U4123 (N_4123,N_1053,N_2111);
nand U4124 (N_4124,N_1654,N_2098);
nand U4125 (N_4125,N_1140,N_2695);
or U4126 (N_4126,N_2225,N_2574);
nand U4127 (N_4127,N_1226,N_2155);
nor U4128 (N_4128,N_225,N_855);
and U4129 (N_4129,N_700,N_2008);
and U4130 (N_4130,N_1406,N_1414);
and U4131 (N_4131,N_546,N_2375);
or U4132 (N_4132,N_2314,N_989);
or U4133 (N_4133,N_334,N_1020);
or U4134 (N_4134,N_420,N_1250);
and U4135 (N_4135,N_1907,N_2191);
nor U4136 (N_4136,N_2887,N_2844);
nand U4137 (N_4137,N_2603,N_1187);
or U4138 (N_4138,N_1738,N_1666);
nor U4139 (N_4139,N_2573,N_1956);
or U4140 (N_4140,N_1136,N_1908);
and U4141 (N_4141,N_1191,N_1648);
nor U4142 (N_4142,N_1833,N_2436);
nand U4143 (N_4143,N_88,N_1677);
nand U4144 (N_4144,N_2926,N_2873);
or U4145 (N_4145,N_135,N_1989);
or U4146 (N_4146,N_2317,N_250);
or U4147 (N_4147,N_872,N_1005);
nand U4148 (N_4148,N_2063,N_887);
and U4149 (N_4149,N_2522,N_1597);
nor U4150 (N_4150,N_2290,N_563);
nand U4151 (N_4151,N_105,N_1378);
or U4152 (N_4152,N_1084,N_2494);
nor U4153 (N_4153,N_625,N_2559);
nand U4154 (N_4154,N_2853,N_1674);
nor U4155 (N_4155,N_2756,N_1085);
nand U4156 (N_4156,N_408,N_846);
or U4157 (N_4157,N_2744,N_1568);
nand U4158 (N_4158,N_251,N_2260);
nor U4159 (N_4159,N_2736,N_2037);
and U4160 (N_4160,N_655,N_2945);
nor U4161 (N_4161,N_764,N_661);
nand U4162 (N_4162,N_2517,N_597);
nor U4163 (N_4163,N_2301,N_942);
nor U4164 (N_4164,N_968,N_2623);
or U4165 (N_4165,N_1203,N_1474);
nor U4166 (N_4166,N_142,N_1594);
and U4167 (N_4167,N_1686,N_4);
nor U4168 (N_4168,N_1511,N_2903);
or U4169 (N_4169,N_1603,N_2636);
nand U4170 (N_4170,N_971,N_451);
nand U4171 (N_4171,N_2998,N_1240);
nor U4172 (N_4172,N_2476,N_237);
nand U4173 (N_4173,N_1619,N_2690);
and U4174 (N_4174,N_58,N_1122);
and U4175 (N_4175,N_824,N_35);
and U4176 (N_4176,N_927,N_2881);
nand U4177 (N_4177,N_441,N_1875);
nor U4178 (N_4178,N_193,N_1332);
or U4179 (N_4179,N_984,N_1943);
or U4180 (N_4180,N_75,N_517);
xor U4181 (N_4181,N_2451,N_190);
nand U4182 (N_4182,N_2777,N_2420);
nor U4183 (N_4183,N_1546,N_1621);
or U4184 (N_4184,N_1258,N_536);
and U4185 (N_4185,N_695,N_1733);
nor U4186 (N_4186,N_1116,N_1370);
nor U4187 (N_4187,N_2174,N_122);
nand U4188 (N_4188,N_1281,N_2329);
nand U4189 (N_4189,N_1742,N_2387);
or U4190 (N_4190,N_2031,N_1818);
or U4191 (N_4191,N_1662,N_235);
or U4192 (N_4192,N_404,N_2908);
and U4193 (N_4193,N_673,N_2982);
nor U4194 (N_4194,N_2384,N_1745);
and U4195 (N_4195,N_664,N_899);
nand U4196 (N_4196,N_454,N_449);
and U4197 (N_4197,N_827,N_2529);
or U4198 (N_4198,N_2627,N_2179);
or U4199 (N_4199,N_2519,N_1565);
nor U4200 (N_4200,N_2509,N_2581);
nor U4201 (N_4201,N_566,N_1069);
and U4202 (N_4202,N_2321,N_2757);
nor U4203 (N_4203,N_303,N_197);
and U4204 (N_4204,N_630,N_212);
or U4205 (N_4205,N_2141,N_2500);
and U4206 (N_4206,N_1466,N_2370);
nand U4207 (N_4207,N_1798,N_1175);
or U4208 (N_4208,N_415,N_817);
nor U4209 (N_4209,N_2085,N_2176);
nand U4210 (N_4210,N_2162,N_721);
nor U4211 (N_4211,N_445,N_522);
nand U4212 (N_4212,N_2977,N_2105);
and U4213 (N_4213,N_1566,N_825);
nor U4214 (N_4214,N_2511,N_71);
and U4215 (N_4215,N_2227,N_385);
xnor U4216 (N_4216,N_494,N_2303);
or U4217 (N_4217,N_2469,N_490);
nor U4218 (N_4218,N_271,N_322);
nand U4219 (N_4219,N_2932,N_499);
and U4220 (N_4220,N_2220,N_769);
and U4221 (N_4221,N_2978,N_1794);
and U4222 (N_4222,N_406,N_292);
and U4223 (N_4223,N_1079,N_2058);
nand U4224 (N_4224,N_931,N_1091);
nor U4225 (N_4225,N_549,N_1395);
or U4226 (N_4226,N_2397,N_2986);
and U4227 (N_4227,N_766,N_483);
xnor U4228 (N_4228,N_762,N_335);
and U4229 (N_4229,N_715,N_869);
or U4230 (N_4230,N_2128,N_2714);
nor U4231 (N_4231,N_2882,N_1499);
and U4232 (N_4232,N_1367,N_2731);
or U4233 (N_4233,N_1527,N_1372);
or U4234 (N_4234,N_384,N_2523);
or U4235 (N_4235,N_1672,N_1305);
or U4236 (N_4236,N_2619,N_175);
nand U4237 (N_4237,N_2755,N_2925);
nand U4238 (N_4238,N_203,N_2889);
nand U4239 (N_4239,N_1739,N_2934);
nor U4240 (N_4240,N_2704,N_1381);
nand U4241 (N_4241,N_2283,N_261);
nor U4242 (N_4242,N_2796,N_12);
nand U4243 (N_4243,N_1793,N_391);
or U4244 (N_4244,N_2121,N_2869);
and U4245 (N_4245,N_1889,N_154);
nor U4246 (N_4246,N_2613,N_2875);
xor U4247 (N_4247,N_1086,N_1018);
nand U4248 (N_4248,N_1835,N_840);
nor U4249 (N_4249,N_196,N_2139);
or U4250 (N_4250,N_2774,N_1915);
or U4251 (N_4251,N_2140,N_852);
nand U4252 (N_4252,N_1872,N_39);
xnor U4253 (N_4253,N_757,N_1148);
nor U4254 (N_4254,N_2028,N_1918);
nand U4255 (N_4255,N_2782,N_2209);
nor U4256 (N_4256,N_1448,N_1512);
nand U4257 (N_4257,N_2022,N_1051);
or U4258 (N_4258,N_1823,N_1737);
nand U4259 (N_4259,N_734,N_1984);
nand U4260 (N_4260,N_706,N_2342);
xnor U4261 (N_4261,N_738,N_1221);
and U4262 (N_4262,N_1516,N_826);
and U4263 (N_4263,N_359,N_581);
nor U4264 (N_4264,N_2878,N_467);
nand U4265 (N_4265,N_710,N_540);
nand U4266 (N_4266,N_1938,N_1062);
or U4267 (N_4267,N_586,N_853);
or U4268 (N_4268,N_2555,N_1831);
and U4269 (N_4269,N_1505,N_871);
nor U4270 (N_4270,N_1164,N_1717);
xor U4271 (N_4271,N_364,N_1118);
nand U4272 (N_4272,N_1612,N_382);
or U4273 (N_4273,N_353,N_114);
and U4274 (N_4274,N_1247,N_2115);
xor U4275 (N_4275,N_692,N_804);
nor U4276 (N_4276,N_1431,N_2461);
or U4277 (N_4277,N_2709,N_2980);
nor U4278 (N_4278,N_1795,N_651);
and U4279 (N_4279,N_2442,N_859);
and U4280 (N_4280,N_934,N_2004);
nor U4281 (N_4281,N_778,N_482);
and U4282 (N_4282,N_1299,N_993);
and U4283 (N_4283,N_2512,N_1425);
or U4284 (N_4284,N_919,N_2430);
and U4285 (N_4285,N_1355,N_399);
nor U4286 (N_4286,N_733,N_1277);
nor U4287 (N_4287,N_2193,N_703);
or U4288 (N_4288,N_745,N_362);
and U4289 (N_4289,N_643,N_2296);
and U4290 (N_4290,N_1039,N_1035);
and U4291 (N_4291,N_2480,N_2991);
or U4292 (N_4292,N_2891,N_2778);
or U4293 (N_4293,N_932,N_2478);
or U4294 (N_4294,N_2327,N_2081);
nand U4295 (N_4295,N_2569,N_2950);
or U4296 (N_4296,N_829,N_2459);
and U4297 (N_4297,N_751,N_1522);
or U4298 (N_4298,N_1828,N_1663);
or U4299 (N_4299,N_2083,N_2589);
nand U4300 (N_4300,N_759,N_469);
nand U4301 (N_4301,N_148,N_2894);
and U4302 (N_4302,N_1906,N_1646);
or U4303 (N_4303,N_479,N_1383);
nor U4304 (N_4304,N_1286,N_657);
and U4305 (N_4305,N_1576,N_842);
and U4306 (N_4306,N_2059,N_2422);
and U4307 (N_4307,N_1707,N_858);
and U4308 (N_4308,N_2674,N_2672);
and U4309 (N_4309,N_864,N_1939);
nand U4310 (N_4310,N_1757,N_1340);
nand U4311 (N_4311,N_1656,N_946);
nor U4312 (N_4312,N_20,N_2677);
nand U4313 (N_4313,N_330,N_1846);
nand U4314 (N_4314,N_1869,N_1800);
nor U4315 (N_4315,N_2944,N_2253);
and U4316 (N_4316,N_2041,N_232);
nand U4317 (N_4317,N_1072,N_531);
nand U4318 (N_4318,N_1326,N_917);
nand U4319 (N_4319,N_434,N_484);
xnor U4320 (N_4320,N_2806,N_2434);
xor U4321 (N_4321,N_185,N_268);
nor U4322 (N_4322,N_555,N_918);
and U4323 (N_4323,N_2808,N_1582);
nor U4324 (N_4324,N_2836,N_609);
nand U4325 (N_4325,N_2601,N_2838);
or U4326 (N_4326,N_179,N_1735);
and U4327 (N_4327,N_2605,N_2123);
or U4328 (N_4328,N_2819,N_1513);
nor U4329 (N_4329,N_2304,N_1840);
and U4330 (N_4330,N_229,N_2761);
nor U4331 (N_4331,N_602,N_1661);
or U4332 (N_4332,N_200,N_771);
nand U4333 (N_4333,N_701,N_674);
and U4334 (N_4334,N_1966,N_2395);
nor U4335 (N_4335,N_2765,N_1216);
or U4336 (N_4336,N_888,N_1357);
or U4337 (N_4337,N_527,N_889);
or U4338 (N_4338,N_2094,N_143);
xnor U4339 (N_4339,N_1667,N_280);
nand U4340 (N_4340,N_1912,N_163);
or U4341 (N_4341,N_1983,N_2652);
nor U4342 (N_4342,N_2971,N_668);
xor U4343 (N_4343,N_2666,N_1335);
or U4344 (N_4344,N_174,N_2560);
or U4345 (N_4345,N_2642,N_1211);
nor U4346 (N_4346,N_2563,N_830);
nand U4347 (N_4347,N_2102,N_2432);
nand U4348 (N_4348,N_311,N_1520);
nor U4349 (N_4349,N_2231,N_638);
and U4350 (N_4350,N_1390,N_1438);
and U4351 (N_4351,N_2813,N_686);
and U4352 (N_4352,N_2086,N_556);
or U4353 (N_4353,N_1227,N_2343);
nand U4354 (N_4354,N_1002,N_1564);
nand U4355 (N_4355,N_2328,N_2611);
and U4356 (N_4356,N_2582,N_1376);
and U4357 (N_4357,N_1537,N_1046);
nand U4358 (N_4358,N_487,N_2368);
nor U4359 (N_4359,N_1444,N_480);
and U4360 (N_4360,N_2104,N_337);
nand U4361 (N_4361,N_2021,N_2876);
nor U4362 (N_4362,N_1770,N_136);
nor U4363 (N_4363,N_1992,N_2799);
or U4364 (N_4364,N_2787,N_2753);
nor U4365 (N_4365,N_1095,N_1339);
or U4366 (N_4366,N_1751,N_970);
and U4367 (N_4367,N_1838,N_518);
nand U4368 (N_4368,N_2196,N_160);
and U4369 (N_4369,N_493,N_1993);
nand U4370 (N_4370,N_140,N_264);
and U4371 (N_4371,N_2817,N_346);
or U4372 (N_4372,N_2531,N_593);
nand U4373 (N_4373,N_1183,N_2906);
and U4374 (N_4374,N_2160,N_1964);
and U4375 (N_4375,N_1986,N_1977);
nand U4376 (N_4376,N_2194,N_1700);
xnor U4377 (N_4377,N_2200,N_2922);
and U4378 (N_4378,N_2182,N_189);
and U4379 (N_4379,N_150,N_1892);
or U4380 (N_4380,N_792,N_2431);
or U4381 (N_4381,N_1789,N_297);
or U4382 (N_4382,N_43,N_187);
nand U4383 (N_4383,N_736,N_1212);
or U4384 (N_4384,N_1691,N_1647);
and U4385 (N_4385,N_1054,N_2418);
nor U4386 (N_4386,N_2931,N_1008);
nor U4387 (N_4387,N_1803,N_2113);
nand U4388 (N_4388,N_217,N_1098);
nand U4389 (N_4389,N_1640,N_1195);
nor U4390 (N_4390,N_2190,N_1309);
or U4391 (N_4391,N_2750,N_681);
nor U4392 (N_4392,N_2310,N_2389);
or U4393 (N_4393,N_2754,N_832);
or U4394 (N_4394,N_719,N_972);
nand U4395 (N_4395,N_2490,N_355);
nor U4396 (N_4396,N_2952,N_356);
nor U4397 (N_4397,N_287,N_1134);
nor U4398 (N_4398,N_608,N_1308);
nor U4399 (N_4399,N_1948,N_2355);
or U4400 (N_4400,N_2029,N_222);
nor U4401 (N_4401,N_2072,N_1412);
nor U4402 (N_4402,N_1507,N_2760);
nand U4403 (N_4403,N_2177,N_1199);
or U4404 (N_4404,N_2893,N_109);
and U4405 (N_4405,N_1421,N_1664);
nand U4406 (N_4406,N_1703,N_1343);
nand U4407 (N_4407,N_693,N_1541);
nand U4408 (N_4408,N_2773,N_1450);
nand U4409 (N_4409,N_1185,N_1325);
and U4410 (N_4410,N_153,N_2939);
or U4411 (N_4411,N_1779,N_1419);
or U4412 (N_4412,N_2616,N_2380);
and U4413 (N_4413,N_2302,N_1074);
or U4414 (N_4414,N_1962,N_895);
or U4415 (N_4415,N_2097,N_1169);
nor U4416 (N_4416,N_128,N_1436);
or U4417 (N_4417,N_1483,N_141);
and U4418 (N_4418,N_572,N_223);
nor U4419 (N_4419,N_2251,N_1917);
or U4420 (N_4420,N_1699,N_744);
nand U4421 (N_4421,N_180,N_1563);
nor U4422 (N_4422,N_1580,N_147);
and U4423 (N_4423,N_2334,N_1508);
nor U4424 (N_4424,N_1731,N_169);
and U4425 (N_4425,N_862,N_1998);
nand U4426 (N_4426,N_799,N_2035);
and U4427 (N_4427,N_2427,N_2280);
and U4428 (N_4428,N_2972,N_288);
xor U4429 (N_4429,N_2682,N_272);
nor U4430 (N_4430,N_662,N_2443);
nor U4431 (N_4431,N_2249,N_891);
and U4432 (N_4432,N_1721,N_2981);
and U4433 (N_4433,N_923,N_2828);
nor U4434 (N_4434,N_1927,N_2997);
and U4435 (N_4435,N_2172,N_1670);
nor U4436 (N_4436,N_312,N_788);
nor U4437 (N_4437,N_1758,N_2852);
nor U4438 (N_4438,N_1310,N_1771);
and U4439 (N_4439,N_2956,N_1796);
and U4440 (N_4440,N_1592,N_675);
or U4441 (N_4441,N_252,N_2861);
or U4442 (N_4442,N_1764,N_1396);
nand U4443 (N_4443,N_1259,N_2830);
or U4444 (N_4444,N_1521,N_1353);
nor U4445 (N_4445,N_1078,N_1826);
nor U4446 (N_4446,N_1413,N_981);
nand U4447 (N_4447,N_2471,N_210);
nor U4448 (N_4448,N_2854,N_107);
nand U4449 (N_4449,N_1189,N_1048);
nor U4450 (N_4450,N_2391,N_2188);
nand U4451 (N_4451,N_2530,N_201);
xnor U4452 (N_4452,N_85,N_588);
nor U4453 (N_4453,N_1613,N_1170);
or U4454 (N_4454,N_911,N_750);
nand U4455 (N_4455,N_2221,N_1526);
nor U4456 (N_4456,N_2818,N_1924);
and U4457 (N_4457,N_1549,N_1028);
or U4458 (N_4458,N_598,N_463);
nor U4459 (N_4459,N_365,N_528);
and U4460 (N_4460,N_1391,N_534);
and U4461 (N_4461,N_57,N_1402);
and U4462 (N_4462,N_1813,N_1394);
nand U4463 (N_4463,N_2566,N_519);
or U4464 (N_4464,N_1812,N_86);
or U4465 (N_4465,N_2292,N_380);
and U4466 (N_4466,N_959,N_1903);
nor U4467 (N_4467,N_1890,N_2584);
or U4468 (N_4468,N_2101,N_698);
nor U4469 (N_4469,N_2974,N_831);
xor U4470 (N_4470,N_2504,N_1238);
and U4471 (N_4471,N_2953,N_1405);
and U4472 (N_4472,N_1971,N_897);
and U4473 (N_4473,N_2949,N_2745);
or U4474 (N_4474,N_2144,N_221);
nor U4475 (N_4475,N_477,N_997);
or U4476 (N_4476,N_124,N_1807);
or U4477 (N_4477,N_860,N_13);
or U4478 (N_4478,N_1163,N_2410);
or U4479 (N_4479,N_779,N_874);
or U4480 (N_4480,N_198,N_2463);
nor U4481 (N_4481,N_2065,N_90);
xnor U4482 (N_4482,N_2919,N_2676);
or U4483 (N_4483,N_1778,N_1113);
nand U4484 (N_4484,N_2013,N_1557);
nor U4485 (N_4485,N_2902,N_1602);
or U4486 (N_4486,N_801,N_81);
nor U4487 (N_4487,N_2275,N_1805);
nor U4488 (N_4488,N_1684,N_2780);
nor U4489 (N_4489,N_2706,N_453);
and U4490 (N_4490,N_680,N_1401);
or U4491 (N_4491,N_2734,N_2142);
and U4492 (N_4492,N_2357,N_1525);
and U4493 (N_4493,N_328,N_438);
or U4494 (N_4494,N_1239,N_1501);
nand U4495 (N_4495,N_1628,N_915);
nor U4496 (N_4496,N_1577,N_2239);
nor U4497 (N_4497,N_49,N_980);
nand U4498 (N_4498,N_1901,N_1825);
and U4499 (N_4499,N_1186,N_1057);
and U4500 (N_4500,N_1598,N_2437);
or U4501 (N_4501,N_139,N_2696);
nand U4502 (N_4502,N_1709,N_1359);
and U4503 (N_4503,N_2605,N_2107);
nand U4504 (N_4504,N_86,N_2409);
nand U4505 (N_4505,N_1722,N_1826);
or U4506 (N_4506,N_2899,N_656);
nor U4507 (N_4507,N_654,N_1708);
nor U4508 (N_4508,N_2224,N_2515);
or U4509 (N_4509,N_1472,N_2022);
nand U4510 (N_4510,N_513,N_168);
nor U4511 (N_4511,N_1824,N_2330);
nand U4512 (N_4512,N_174,N_2050);
nor U4513 (N_4513,N_1634,N_861);
or U4514 (N_4514,N_340,N_616);
and U4515 (N_4515,N_2699,N_1628);
nor U4516 (N_4516,N_29,N_943);
and U4517 (N_4517,N_1947,N_578);
xnor U4518 (N_4518,N_2152,N_1854);
nand U4519 (N_4519,N_1386,N_1366);
nand U4520 (N_4520,N_2361,N_2706);
nand U4521 (N_4521,N_2216,N_861);
nor U4522 (N_4522,N_1255,N_1725);
and U4523 (N_4523,N_1120,N_39);
nor U4524 (N_4524,N_2069,N_1082);
and U4525 (N_4525,N_975,N_849);
and U4526 (N_4526,N_358,N_2757);
and U4527 (N_4527,N_2266,N_2701);
nor U4528 (N_4528,N_948,N_1135);
nor U4529 (N_4529,N_1984,N_1300);
nor U4530 (N_4530,N_2248,N_1551);
xor U4531 (N_4531,N_2247,N_796);
and U4532 (N_4532,N_1444,N_2870);
or U4533 (N_4533,N_392,N_1515);
or U4534 (N_4534,N_2501,N_289);
and U4535 (N_4535,N_2932,N_2745);
and U4536 (N_4536,N_1941,N_1094);
or U4537 (N_4537,N_1993,N_446);
nand U4538 (N_4538,N_697,N_26);
or U4539 (N_4539,N_1642,N_1562);
nor U4540 (N_4540,N_2954,N_175);
nor U4541 (N_4541,N_2918,N_1664);
and U4542 (N_4542,N_2839,N_225);
and U4543 (N_4543,N_2389,N_1637);
nor U4544 (N_4544,N_93,N_2832);
nor U4545 (N_4545,N_2850,N_2765);
or U4546 (N_4546,N_251,N_2186);
and U4547 (N_4547,N_1728,N_2675);
nor U4548 (N_4548,N_1028,N_889);
nand U4549 (N_4549,N_197,N_1279);
and U4550 (N_4550,N_902,N_923);
nand U4551 (N_4551,N_225,N_1610);
nor U4552 (N_4552,N_1010,N_397);
nand U4553 (N_4553,N_1249,N_2421);
nor U4554 (N_4554,N_752,N_2462);
nor U4555 (N_4555,N_2493,N_332);
nand U4556 (N_4556,N_2695,N_709);
nand U4557 (N_4557,N_271,N_925);
nand U4558 (N_4558,N_1683,N_2582);
nor U4559 (N_4559,N_1199,N_625);
nor U4560 (N_4560,N_826,N_1257);
and U4561 (N_4561,N_2732,N_2906);
and U4562 (N_4562,N_1692,N_1563);
and U4563 (N_4563,N_2840,N_620);
and U4564 (N_4564,N_1074,N_1043);
or U4565 (N_4565,N_894,N_49);
and U4566 (N_4566,N_476,N_2982);
nor U4567 (N_4567,N_1054,N_965);
nor U4568 (N_4568,N_1638,N_2592);
and U4569 (N_4569,N_2517,N_2279);
and U4570 (N_4570,N_1173,N_1174);
nor U4571 (N_4571,N_1594,N_2817);
or U4572 (N_4572,N_1516,N_2476);
or U4573 (N_4573,N_1787,N_1336);
nand U4574 (N_4574,N_207,N_1175);
nor U4575 (N_4575,N_99,N_1283);
xor U4576 (N_4576,N_1906,N_1468);
or U4577 (N_4577,N_1635,N_114);
or U4578 (N_4578,N_1792,N_2845);
nand U4579 (N_4579,N_2725,N_2188);
and U4580 (N_4580,N_2814,N_2109);
nand U4581 (N_4581,N_1596,N_2040);
or U4582 (N_4582,N_2412,N_1166);
nand U4583 (N_4583,N_2749,N_2365);
nor U4584 (N_4584,N_2435,N_2324);
and U4585 (N_4585,N_518,N_863);
nor U4586 (N_4586,N_2497,N_2908);
or U4587 (N_4587,N_2424,N_1697);
nand U4588 (N_4588,N_2622,N_2638);
and U4589 (N_4589,N_114,N_1920);
nor U4590 (N_4590,N_2108,N_1029);
or U4591 (N_4591,N_960,N_1236);
or U4592 (N_4592,N_1826,N_944);
and U4593 (N_4593,N_2475,N_2371);
or U4594 (N_4594,N_1521,N_1920);
nand U4595 (N_4595,N_1846,N_1948);
xor U4596 (N_4596,N_1112,N_216);
nor U4597 (N_4597,N_876,N_1980);
nor U4598 (N_4598,N_1641,N_267);
nor U4599 (N_4599,N_1124,N_924);
nor U4600 (N_4600,N_505,N_2171);
and U4601 (N_4601,N_2454,N_1998);
and U4602 (N_4602,N_2360,N_68);
and U4603 (N_4603,N_1079,N_2187);
nand U4604 (N_4604,N_448,N_1066);
or U4605 (N_4605,N_335,N_2085);
or U4606 (N_4606,N_1906,N_2731);
or U4607 (N_4607,N_233,N_1817);
or U4608 (N_4608,N_1597,N_2429);
nand U4609 (N_4609,N_2496,N_1087);
nor U4610 (N_4610,N_2831,N_2153);
nand U4611 (N_4611,N_1745,N_748);
nor U4612 (N_4612,N_646,N_2768);
or U4613 (N_4613,N_1253,N_466);
or U4614 (N_4614,N_2498,N_366);
or U4615 (N_4615,N_1361,N_1241);
and U4616 (N_4616,N_33,N_2045);
or U4617 (N_4617,N_2794,N_1141);
and U4618 (N_4618,N_2941,N_2642);
and U4619 (N_4619,N_650,N_2120);
and U4620 (N_4620,N_1496,N_2135);
nand U4621 (N_4621,N_2128,N_2475);
nand U4622 (N_4622,N_1436,N_2986);
and U4623 (N_4623,N_1363,N_1911);
nand U4624 (N_4624,N_2427,N_1119);
xnor U4625 (N_4625,N_2331,N_2233);
nor U4626 (N_4626,N_2206,N_1666);
or U4627 (N_4627,N_2139,N_1738);
or U4628 (N_4628,N_1905,N_1694);
and U4629 (N_4629,N_2891,N_2906);
nor U4630 (N_4630,N_395,N_1548);
or U4631 (N_4631,N_968,N_672);
nand U4632 (N_4632,N_2843,N_412);
nor U4633 (N_4633,N_1878,N_2406);
or U4634 (N_4634,N_346,N_1629);
nor U4635 (N_4635,N_2895,N_2070);
and U4636 (N_4636,N_132,N_1404);
xnor U4637 (N_4637,N_2552,N_2589);
nor U4638 (N_4638,N_2906,N_791);
and U4639 (N_4639,N_822,N_1910);
nor U4640 (N_4640,N_2953,N_1135);
and U4641 (N_4641,N_99,N_2009);
and U4642 (N_4642,N_124,N_900);
and U4643 (N_4643,N_917,N_806);
or U4644 (N_4644,N_1436,N_2097);
and U4645 (N_4645,N_1516,N_1908);
or U4646 (N_4646,N_1082,N_1361);
nand U4647 (N_4647,N_1110,N_767);
nor U4648 (N_4648,N_2998,N_1573);
or U4649 (N_4649,N_510,N_1757);
or U4650 (N_4650,N_1833,N_1719);
and U4651 (N_4651,N_700,N_1692);
nand U4652 (N_4652,N_194,N_2359);
or U4653 (N_4653,N_2777,N_1971);
nor U4654 (N_4654,N_955,N_775);
and U4655 (N_4655,N_688,N_237);
and U4656 (N_4656,N_1208,N_2959);
nor U4657 (N_4657,N_2159,N_724);
nand U4658 (N_4658,N_2605,N_628);
nand U4659 (N_4659,N_65,N_299);
and U4660 (N_4660,N_1447,N_417);
and U4661 (N_4661,N_1960,N_521);
nor U4662 (N_4662,N_2882,N_2962);
nor U4663 (N_4663,N_2420,N_1464);
or U4664 (N_4664,N_2299,N_2088);
and U4665 (N_4665,N_425,N_2651);
and U4666 (N_4666,N_2259,N_2011);
and U4667 (N_4667,N_1608,N_246);
nand U4668 (N_4668,N_2645,N_228);
and U4669 (N_4669,N_590,N_1286);
and U4670 (N_4670,N_2243,N_2626);
or U4671 (N_4671,N_190,N_2845);
xnor U4672 (N_4672,N_353,N_1154);
and U4673 (N_4673,N_741,N_1177);
or U4674 (N_4674,N_174,N_391);
or U4675 (N_4675,N_304,N_2465);
and U4676 (N_4676,N_1157,N_1423);
nor U4677 (N_4677,N_930,N_2069);
nor U4678 (N_4678,N_1124,N_2519);
nand U4679 (N_4679,N_2783,N_1727);
nand U4680 (N_4680,N_2494,N_2302);
nor U4681 (N_4681,N_1964,N_1283);
or U4682 (N_4682,N_1977,N_1257);
nor U4683 (N_4683,N_928,N_1317);
nor U4684 (N_4684,N_318,N_1205);
or U4685 (N_4685,N_214,N_773);
or U4686 (N_4686,N_2329,N_1949);
and U4687 (N_4687,N_1145,N_744);
nand U4688 (N_4688,N_2592,N_1873);
and U4689 (N_4689,N_784,N_1775);
and U4690 (N_4690,N_2463,N_1484);
xnor U4691 (N_4691,N_363,N_2760);
nor U4692 (N_4692,N_2244,N_1131);
and U4693 (N_4693,N_1801,N_2192);
or U4694 (N_4694,N_1744,N_2198);
or U4695 (N_4695,N_2153,N_608);
xnor U4696 (N_4696,N_285,N_1602);
nor U4697 (N_4697,N_1305,N_98);
nand U4698 (N_4698,N_1175,N_777);
nor U4699 (N_4699,N_199,N_1132);
and U4700 (N_4700,N_1144,N_1299);
or U4701 (N_4701,N_253,N_326);
xor U4702 (N_4702,N_592,N_2197);
and U4703 (N_4703,N_2057,N_2023);
nor U4704 (N_4704,N_398,N_1369);
nor U4705 (N_4705,N_2384,N_2440);
and U4706 (N_4706,N_13,N_2847);
or U4707 (N_4707,N_1715,N_872);
or U4708 (N_4708,N_2444,N_2541);
and U4709 (N_4709,N_1362,N_1858);
and U4710 (N_4710,N_2801,N_789);
nor U4711 (N_4711,N_680,N_2449);
or U4712 (N_4712,N_2025,N_1402);
or U4713 (N_4713,N_25,N_1455);
nand U4714 (N_4714,N_1644,N_1807);
and U4715 (N_4715,N_2565,N_2384);
nand U4716 (N_4716,N_1796,N_194);
or U4717 (N_4717,N_1166,N_1485);
nand U4718 (N_4718,N_2833,N_533);
and U4719 (N_4719,N_2448,N_2097);
nand U4720 (N_4720,N_831,N_2093);
and U4721 (N_4721,N_2742,N_2901);
or U4722 (N_4722,N_1839,N_2361);
or U4723 (N_4723,N_1825,N_996);
and U4724 (N_4724,N_2111,N_1391);
nand U4725 (N_4725,N_1840,N_688);
or U4726 (N_4726,N_999,N_758);
or U4727 (N_4727,N_1753,N_2687);
or U4728 (N_4728,N_557,N_2390);
nor U4729 (N_4729,N_1275,N_664);
nand U4730 (N_4730,N_2679,N_1133);
nor U4731 (N_4731,N_298,N_2079);
nor U4732 (N_4732,N_1064,N_2822);
xnor U4733 (N_4733,N_1566,N_2003);
nor U4734 (N_4734,N_2711,N_1770);
nand U4735 (N_4735,N_2287,N_1184);
and U4736 (N_4736,N_2546,N_2184);
nand U4737 (N_4737,N_673,N_2683);
and U4738 (N_4738,N_1870,N_1315);
nand U4739 (N_4739,N_2589,N_1649);
nand U4740 (N_4740,N_50,N_2953);
nor U4741 (N_4741,N_1064,N_754);
nor U4742 (N_4742,N_2489,N_1201);
nor U4743 (N_4743,N_1574,N_2595);
nor U4744 (N_4744,N_2065,N_1905);
nor U4745 (N_4745,N_1667,N_2602);
or U4746 (N_4746,N_2026,N_2258);
or U4747 (N_4747,N_2751,N_389);
and U4748 (N_4748,N_2593,N_540);
and U4749 (N_4749,N_1709,N_1625);
xnor U4750 (N_4750,N_1055,N_748);
or U4751 (N_4751,N_1344,N_1316);
nor U4752 (N_4752,N_1276,N_121);
nor U4753 (N_4753,N_1493,N_534);
nand U4754 (N_4754,N_1552,N_1709);
nor U4755 (N_4755,N_1426,N_2935);
nor U4756 (N_4756,N_1810,N_1295);
or U4757 (N_4757,N_1883,N_1220);
nor U4758 (N_4758,N_1045,N_1641);
nand U4759 (N_4759,N_1991,N_878);
nand U4760 (N_4760,N_1034,N_698);
nor U4761 (N_4761,N_367,N_1357);
and U4762 (N_4762,N_1448,N_1679);
nand U4763 (N_4763,N_2894,N_2705);
nand U4764 (N_4764,N_1039,N_2834);
and U4765 (N_4765,N_1529,N_2088);
nor U4766 (N_4766,N_1049,N_772);
nand U4767 (N_4767,N_2059,N_2225);
or U4768 (N_4768,N_1479,N_2646);
and U4769 (N_4769,N_2542,N_2086);
nand U4770 (N_4770,N_2214,N_1257);
or U4771 (N_4771,N_1861,N_2773);
or U4772 (N_4772,N_2403,N_2120);
and U4773 (N_4773,N_481,N_443);
or U4774 (N_4774,N_1548,N_2887);
nand U4775 (N_4775,N_1520,N_1699);
and U4776 (N_4776,N_882,N_1167);
nor U4777 (N_4777,N_387,N_79);
and U4778 (N_4778,N_1504,N_1143);
nand U4779 (N_4779,N_2582,N_2789);
nand U4780 (N_4780,N_1876,N_2781);
and U4781 (N_4781,N_377,N_598);
and U4782 (N_4782,N_2662,N_1748);
or U4783 (N_4783,N_739,N_2937);
nor U4784 (N_4784,N_2399,N_839);
nor U4785 (N_4785,N_723,N_1411);
xor U4786 (N_4786,N_715,N_1957);
and U4787 (N_4787,N_2004,N_1300);
nand U4788 (N_4788,N_1520,N_2474);
or U4789 (N_4789,N_2768,N_1786);
nor U4790 (N_4790,N_1641,N_1193);
and U4791 (N_4791,N_2433,N_2793);
or U4792 (N_4792,N_275,N_884);
and U4793 (N_4793,N_625,N_10);
nand U4794 (N_4794,N_1033,N_39);
nor U4795 (N_4795,N_1395,N_2558);
or U4796 (N_4796,N_2941,N_920);
or U4797 (N_4797,N_2390,N_1699);
or U4798 (N_4798,N_2901,N_2306);
and U4799 (N_4799,N_2232,N_2713);
nand U4800 (N_4800,N_930,N_2852);
nand U4801 (N_4801,N_737,N_2593);
nand U4802 (N_4802,N_679,N_1319);
nand U4803 (N_4803,N_2640,N_1599);
nand U4804 (N_4804,N_610,N_1925);
and U4805 (N_4805,N_488,N_487);
or U4806 (N_4806,N_2284,N_1594);
or U4807 (N_4807,N_380,N_1954);
or U4808 (N_4808,N_2627,N_1382);
nor U4809 (N_4809,N_1002,N_1550);
xnor U4810 (N_4810,N_854,N_2540);
nor U4811 (N_4811,N_87,N_575);
and U4812 (N_4812,N_532,N_1333);
nor U4813 (N_4813,N_476,N_1320);
nor U4814 (N_4814,N_331,N_385);
nand U4815 (N_4815,N_2802,N_1953);
and U4816 (N_4816,N_1514,N_17);
and U4817 (N_4817,N_1182,N_1994);
nor U4818 (N_4818,N_2480,N_1660);
and U4819 (N_4819,N_2903,N_521);
nand U4820 (N_4820,N_2305,N_1511);
and U4821 (N_4821,N_2007,N_2383);
xor U4822 (N_4822,N_476,N_99);
nand U4823 (N_4823,N_466,N_730);
nor U4824 (N_4824,N_2836,N_2060);
nand U4825 (N_4825,N_750,N_2500);
nor U4826 (N_4826,N_1903,N_2015);
xor U4827 (N_4827,N_2198,N_1265);
nor U4828 (N_4828,N_2536,N_1871);
or U4829 (N_4829,N_1935,N_799);
nor U4830 (N_4830,N_1213,N_347);
and U4831 (N_4831,N_462,N_537);
and U4832 (N_4832,N_1661,N_1311);
and U4833 (N_4833,N_2901,N_102);
and U4834 (N_4834,N_2022,N_1591);
nand U4835 (N_4835,N_1188,N_1029);
or U4836 (N_4836,N_1719,N_1220);
or U4837 (N_4837,N_1970,N_2664);
or U4838 (N_4838,N_2170,N_1564);
nand U4839 (N_4839,N_907,N_1798);
or U4840 (N_4840,N_1953,N_2405);
and U4841 (N_4841,N_2698,N_163);
and U4842 (N_4842,N_834,N_1674);
xnor U4843 (N_4843,N_2712,N_1415);
or U4844 (N_4844,N_2706,N_2315);
or U4845 (N_4845,N_1894,N_179);
nand U4846 (N_4846,N_1280,N_388);
or U4847 (N_4847,N_2566,N_1764);
and U4848 (N_4848,N_161,N_2829);
nand U4849 (N_4849,N_2803,N_1875);
nor U4850 (N_4850,N_2528,N_1262);
and U4851 (N_4851,N_1078,N_557);
nand U4852 (N_4852,N_2285,N_848);
nand U4853 (N_4853,N_1893,N_1513);
nor U4854 (N_4854,N_2077,N_10);
and U4855 (N_4855,N_2839,N_100);
xor U4856 (N_4856,N_2334,N_1384);
and U4857 (N_4857,N_2215,N_2881);
nor U4858 (N_4858,N_2320,N_1453);
or U4859 (N_4859,N_2850,N_2021);
and U4860 (N_4860,N_818,N_2268);
or U4861 (N_4861,N_2744,N_1628);
nor U4862 (N_4862,N_2179,N_2597);
or U4863 (N_4863,N_952,N_2189);
nor U4864 (N_4864,N_263,N_1684);
or U4865 (N_4865,N_901,N_2886);
xnor U4866 (N_4866,N_2610,N_382);
nor U4867 (N_4867,N_1454,N_711);
nand U4868 (N_4868,N_1331,N_2746);
or U4869 (N_4869,N_2281,N_2235);
and U4870 (N_4870,N_1614,N_2879);
or U4871 (N_4871,N_1224,N_221);
nor U4872 (N_4872,N_2904,N_1712);
or U4873 (N_4873,N_2586,N_318);
and U4874 (N_4874,N_1544,N_1340);
or U4875 (N_4875,N_1652,N_1057);
or U4876 (N_4876,N_2561,N_2727);
nor U4877 (N_4877,N_1248,N_249);
nor U4878 (N_4878,N_1315,N_856);
and U4879 (N_4879,N_24,N_1362);
nand U4880 (N_4880,N_675,N_2944);
nor U4881 (N_4881,N_237,N_776);
and U4882 (N_4882,N_1125,N_289);
and U4883 (N_4883,N_2333,N_2738);
and U4884 (N_4884,N_821,N_1802);
nor U4885 (N_4885,N_2691,N_1057);
nand U4886 (N_4886,N_335,N_2901);
or U4887 (N_4887,N_2308,N_1520);
or U4888 (N_4888,N_2427,N_1616);
nand U4889 (N_4889,N_1387,N_1903);
nor U4890 (N_4890,N_1817,N_1376);
and U4891 (N_4891,N_1970,N_2243);
or U4892 (N_4892,N_1432,N_2600);
nand U4893 (N_4893,N_2820,N_1587);
or U4894 (N_4894,N_2327,N_293);
or U4895 (N_4895,N_1111,N_1456);
or U4896 (N_4896,N_580,N_2090);
and U4897 (N_4897,N_1231,N_1013);
nand U4898 (N_4898,N_1987,N_1330);
or U4899 (N_4899,N_2329,N_2778);
and U4900 (N_4900,N_781,N_1824);
nor U4901 (N_4901,N_1081,N_2115);
and U4902 (N_4902,N_2861,N_434);
and U4903 (N_4903,N_1292,N_2728);
or U4904 (N_4904,N_1031,N_1665);
nand U4905 (N_4905,N_1791,N_2421);
or U4906 (N_4906,N_1888,N_1609);
or U4907 (N_4907,N_1068,N_628);
or U4908 (N_4908,N_1200,N_35);
or U4909 (N_4909,N_194,N_975);
or U4910 (N_4910,N_1601,N_1524);
and U4911 (N_4911,N_2350,N_2935);
and U4912 (N_4912,N_697,N_201);
nand U4913 (N_4913,N_1729,N_1127);
nand U4914 (N_4914,N_127,N_1856);
nand U4915 (N_4915,N_840,N_1702);
or U4916 (N_4916,N_855,N_1060);
nand U4917 (N_4917,N_1629,N_1808);
and U4918 (N_4918,N_1877,N_2841);
or U4919 (N_4919,N_1241,N_2867);
nand U4920 (N_4920,N_84,N_2286);
nor U4921 (N_4921,N_452,N_906);
and U4922 (N_4922,N_517,N_816);
or U4923 (N_4923,N_1862,N_1311);
nand U4924 (N_4924,N_2256,N_1250);
or U4925 (N_4925,N_2997,N_687);
nand U4926 (N_4926,N_2797,N_2349);
nand U4927 (N_4927,N_301,N_2046);
nand U4928 (N_4928,N_1700,N_1423);
nand U4929 (N_4929,N_2957,N_1534);
nor U4930 (N_4930,N_2082,N_1230);
nor U4931 (N_4931,N_2491,N_1145);
or U4932 (N_4932,N_2827,N_2363);
and U4933 (N_4933,N_2432,N_331);
and U4934 (N_4934,N_1575,N_743);
nor U4935 (N_4935,N_2358,N_2335);
or U4936 (N_4936,N_213,N_1142);
nand U4937 (N_4937,N_199,N_2459);
nand U4938 (N_4938,N_1772,N_548);
or U4939 (N_4939,N_2692,N_1055);
or U4940 (N_4940,N_394,N_1023);
and U4941 (N_4941,N_806,N_2562);
nand U4942 (N_4942,N_1275,N_2886);
nor U4943 (N_4943,N_943,N_2359);
nand U4944 (N_4944,N_1015,N_2280);
nor U4945 (N_4945,N_578,N_288);
or U4946 (N_4946,N_2889,N_2976);
or U4947 (N_4947,N_2641,N_1867);
or U4948 (N_4948,N_1532,N_271);
or U4949 (N_4949,N_1602,N_782);
nor U4950 (N_4950,N_2638,N_1399);
nor U4951 (N_4951,N_2919,N_1711);
or U4952 (N_4952,N_1020,N_2334);
nor U4953 (N_4953,N_2933,N_2948);
nor U4954 (N_4954,N_1472,N_1811);
or U4955 (N_4955,N_2636,N_2431);
xnor U4956 (N_4956,N_2596,N_1261);
nor U4957 (N_4957,N_348,N_2734);
nor U4958 (N_4958,N_540,N_2049);
and U4959 (N_4959,N_1186,N_1899);
or U4960 (N_4960,N_1067,N_2878);
and U4961 (N_4961,N_1557,N_1965);
or U4962 (N_4962,N_928,N_1706);
or U4963 (N_4963,N_961,N_632);
and U4964 (N_4964,N_2551,N_144);
nand U4965 (N_4965,N_263,N_1244);
and U4966 (N_4966,N_1603,N_1183);
or U4967 (N_4967,N_26,N_2818);
nor U4968 (N_4968,N_1663,N_1156);
nor U4969 (N_4969,N_2542,N_2309);
and U4970 (N_4970,N_2193,N_1463);
nand U4971 (N_4971,N_1224,N_567);
nor U4972 (N_4972,N_666,N_2005);
nand U4973 (N_4973,N_1931,N_767);
nor U4974 (N_4974,N_2920,N_2224);
and U4975 (N_4975,N_273,N_1028);
nand U4976 (N_4976,N_1607,N_472);
or U4977 (N_4977,N_513,N_438);
or U4978 (N_4978,N_2053,N_551);
nor U4979 (N_4979,N_209,N_1986);
and U4980 (N_4980,N_2723,N_1187);
nand U4981 (N_4981,N_222,N_1224);
nand U4982 (N_4982,N_2058,N_2427);
nand U4983 (N_4983,N_1103,N_1601);
nand U4984 (N_4984,N_1352,N_921);
nand U4985 (N_4985,N_1224,N_1384);
nor U4986 (N_4986,N_2150,N_2616);
nor U4987 (N_4987,N_912,N_889);
and U4988 (N_4988,N_380,N_2527);
xnor U4989 (N_4989,N_793,N_1390);
xnor U4990 (N_4990,N_2053,N_1905);
nor U4991 (N_4991,N_606,N_1374);
nor U4992 (N_4992,N_2656,N_2511);
and U4993 (N_4993,N_2083,N_615);
nor U4994 (N_4994,N_1138,N_2951);
nor U4995 (N_4995,N_1869,N_255);
and U4996 (N_4996,N_353,N_585);
xnor U4997 (N_4997,N_2736,N_1917);
and U4998 (N_4998,N_2316,N_340);
and U4999 (N_4999,N_1472,N_606);
nand U5000 (N_5000,N_1288,N_2465);
nor U5001 (N_5001,N_1195,N_1679);
and U5002 (N_5002,N_520,N_1669);
and U5003 (N_5003,N_309,N_709);
and U5004 (N_5004,N_2045,N_1322);
and U5005 (N_5005,N_1165,N_267);
nand U5006 (N_5006,N_2096,N_1112);
nand U5007 (N_5007,N_826,N_1741);
and U5008 (N_5008,N_494,N_2186);
nor U5009 (N_5009,N_2811,N_585);
or U5010 (N_5010,N_865,N_591);
nand U5011 (N_5011,N_1341,N_322);
nor U5012 (N_5012,N_176,N_2083);
xor U5013 (N_5013,N_204,N_2203);
or U5014 (N_5014,N_1449,N_1632);
and U5015 (N_5015,N_896,N_35);
and U5016 (N_5016,N_2053,N_2182);
nor U5017 (N_5017,N_1666,N_734);
or U5018 (N_5018,N_2792,N_265);
and U5019 (N_5019,N_2590,N_2455);
or U5020 (N_5020,N_2538,N_1088);
and U5021 (N_5021,N_620,N_174);
or U5022 (N_5022,N_1811,N_504);
nand U5023 (N_5023,N_2210,N_98);
or U5024 (N_5024,N_2412,N_532);
nor U5025 (N_5025,N_1768,N_1264);
and U5026 (N_5026,N_193,N_2264);
nand U5027 (N_5027,N_2979,N_2512);
nor U5028 (N_5028,N_54,N_2278);
and U5029 (N_5029,N_890,N_277);
nand U5030 (N_5030,N_1112,N_1868);
or U5031 (N_5031,N_2656,N_551);
and U5032 (N_5032,N_2960,N_1692);
or U5033 (N_5033,N_2967,N_1543);
nor U5034 (N_5034,N_1127,N_1784);
nor U5035 (N_5035,N_2555,N_1711);
nor U5036 (N_5036,N_476,N_1593);
nand U5037 (N_5037,N_2458,N_928);
and U5038 (N_5038,N_627,N_2397);
and U5039 (N_5039,N_2557,N_1946);
nand U5040 (N_5040,N_2566,N_2986);
xor U5041 (N_5041,N_674,N_2226);
and U5042 (N_5042,N_1661,N_2729);
and U5043 (N_5043,N_2370,N_864);
or U5044 (N_5044,N_1270,N_260);
nor U5045 (N_5045,N_54,N_2928);
nand U5046 (N_5046,N_828,N_2266);
nand U5047 (N_5047,N_341,N_2002);
nand U5048 (N_5048,N_2261,N_987);
nor U5049 (N_5049,N_2526,N_1361);
or U5050 (N_5050,N_2734,N_1605);
nor U5051 (N_5051,N_2332,N_1033);
nand U5052 (N_5052,N_13,N_684);
xnor U5053 (N_5053,N_2330,N_2849);
and U5054 (N_5054,N_525,N_1054);
nor U5055 (N_5055,N_1453,N_204);
and U5056 (N_5056,N_2133,N_498);
and U5057 (N_5057,N_365,N_672);
and U5058 (N_5058,N_676,N_1843);
or U5059 (N_5059,N_2529,N_1686);
and U5060 (N_5060,N_1370,N_1807);
and U5061 (N_5061,N_534,N_2693);
or U5062 (N_5062,N_2300,N_271);
and U5063 (N_5063,N_45,N_2257);
nor U5064 (N_5064,N_807,N_225);
or U5065 (N_5065,N_745,N_1276);
and U5066 (N_5066,N_2501,N_536);
or U5067 (N_5067,N_2312,N_2482);
or U5068 (N_5068,N_1434,N_2609);
and U5069 (N_5069,N_763,N_1985);
nor U5070 (N_5070,N_2795,N_993);
or U5071 (N_5071,N_1800,N_2903);
nand U5072 (N_5072,N_1145,N_1838);
nor U5073 (N_5073,N_800,N_2811);
nor U5074 (N_5074,N_2734,N_102);
xnor U5075 (N_5075,N_2067,N_1289);
and U5076 (N_5076,N_1940,N_1677);
nand U5077 (N_5077,N_2629,N_2855);
and U5078 (N_5078,N_238,N_2126);
xor U5079 (N_5079,N_2393,N_2026);
or U5080 (N_5080,N_2286,N_2606);
nand U5081 (N_5081,N_136,N_1648);
nor U5082 (N_5082,N_1451,N_2716);
nor U5083 (N_5083,N_2532,N_1976);
nand U5084 (N_5084,N_384,N_300);
nand U5085 (N_5085,N_841,N_1693);
nand U5086 (N_5086,N_1888,N_1759);
nor U5087 (N_5087,N_562,N_1009);
nor U5088 (N_5088,N_1233,N_617);
or U5089 (N_5089,N_1722,N_1464);
and U5090 (N_5090,N_2256,N_988);
or U5091 (N_5091,N_1546,N_1644);
or U5092 (N_5092,N_1433,N_2890);
and U5093 (N_5093,N_2903,N_1470);
or U5094 (N_5094,N_2726,N_1203);
and U5095 (N_5095,N_559,N_924);
and U5096 (N_5096,N_349,N_2176);
or U5097 (N_5097,N_581,N_1664);
or U5098 (N_5098,N_720,N_462);
nor U5099 (N_5099,N_658,N_34);
nand U5100 (N_5100,N_1763,N_1733);
or U5101 (N_5101,N_1322,N_1783);
or U5102 (N_5102,N_1984,N_2110);
nor U5103 (N_5103,N_2028,N_259);
or U5104 (N_5104,N_1012,N_963);
nand U5105 (N_5105,N_2470,N_2140);
nand U5106 (N_5106,N_2999,N_2164);
or U5107 (N_5107,N_2193,N_2266);
and U5108 (N_5108,N_2519,N_815);
nand U5109 (N_5109,N_453,N_1610);
nor U5110 (N_5110,N_545,N_1753);
nand U5111 (N_5111,N_1598,N_1976);
nand U5112 (N_5112,N_1481,N_2111);
nor U5113 (N_5113,N_197,N_709);
and U5114 (N_5114,N_1324,N_93);
and U5115 (N_5115,N_409,N_1928);
nor U5116 (N_5116,N_2373,N_1852);
nand U5117 (N_5117,N_2292,N_1727);
nand U5118 (N_5118,N_2295,N_315);
and U5119 (N_5119,N_1010,N_2687);
nand U5120 (N_5120,N_2924,N_803);
nor U5121 (N_5121,N_2054,N_2763);
nor U5122 (N_5122,N_447,N_1370);
nor U5123 (N_5123,N_1801,N_398);
xor U5124 (N_5124,N_1595,N_2465);
or U5125 (N_5125,N_135,N_686);
or U5126 (N_5126,N_2906,N_724);
nand U5127 (N_5127,N_1080,N_1670);
or U5128 (N_5128,N_641,N_1359);
nand U5129 (N_5129,N_1000,N_1652);
nor U5130 (N_5130,N_979,N_1823);
xor U5131 (N_5131,N_2083,N_2336);
nand U5132 (N_5132,N_2129,N_2003);
nand U5133 (N_5133,N_2829,N_145);
and U5134 (N_5134,N_2050,N_1282);
or U5135 (N_5135,N_1735,N_654);
or U5136 (N_5136,N_1366,N_2703);
nand U5137 (N_5137,N_2102,N_792);
and U5138 (N_5138,N_2747,N_2072);
nor U5139 (N_5139,N_2563,N_2084);
and U5140 (N_5140,N_2340,N_2366);
and U5141 (N_5141,N_2745,N_1470);
nand U5142 (N_5142,N_2328,N_710);
nand U5143 (N_5143,N_2776,N_2902);
nand U5144 (N_5144,N_2556,N_2542);
or U5145 (N_5145,N_229,N_448);
nor U5146 (N_5146,N_1596,N_1245);
and U5147 (N_5147,N_1694,N_1725);
and U5148 (N_5148,N_275,N_281);
or U5149 (N_5149,N_2501,N_1378);
nor U5150 (N_5150,N_2036,N_1689);
and U5151 (N_5151,N_2480,N_123);
nor U5152 (N_5152,N_1757,N_1397);
or U5153 (N_5153,N_688,N_1480);
nand U5154 (N_5154,N_869,N_2380);
or U5155 (N_5155,N_802,N_704);
nor U5156 (N_5156,N_256,N_2478);
and U5157 (N_5157,N_2408,N_113);
or U5158 (N_5158,N_2490,N_1923);
and U5159 (N_5159,N_2755,N_931);
nor U5160 (N_5160,N_1204,N_1540);
or U5161 (N_5161,N_511,N_2116);
and U5162 (N_5162,N_2140,N_544);
or U5163 (N_5163,N_219,N_1823);
nor U5164 (N_5164,N_2814,N_1619);
and U5165 (N_5165,N_131,N_1253);
and U5166 (N_5166,N_1196,N_2735);
nand U5167 (N_5167,N_1771,N_2335);
xnor U5168 (N_5168,N_2790,N_2658);
and U5169 (N_5169,N_2642,N_2892);
and U5170 (N_5170,N_2664,N_859);
or U5171 (N_5171,N_2460,N_1253);
xnor U5172 (N_5172,N_2398,N_2582);
or U5173 (N_5173,N_734,N_1486);
nand U5174 (N_5174,N_2249,N_1005);
nand U5175 (N_5175,N_456,N_1519);
nor U5176 (N_5176,N_2635,N_2869);
nand U5177 (N_5177,N_798,N_2449);
and U5178 (N_5178,N_1409,N_2175);
xor U5179 (N_5179,N_929,N_109);
and U5180 (N_5180,N_1484,N_2994);
and U5181 (N_5181,N_1726,N_207);
nand U5182 (N_5182,N_976,N_231);
and U5183 (N_5183,N_1650,N_1375);
nand U5184 (N_5184,N_2160,N_4);
xor U5185 (N_5185,N_741,N_981);
nand U5186 (N_5186,N_1778,N_1317);
and U5187 (N_5187,N_2128,N_217);
nand U5188 (N_5188,N_613,N_1591);
nand U5189 (N_5189,N_2494,N_672);
nor U5190 (N_5190,N_654,N_2099);
and U5191 (N_5191,N_2752,N_808);
and U5192 (N_5192,N_935,N_1455);
and U5193 (N_5193,N_1877,N_2724);
nand U5194 (N_5194,N_1903,N_68);
or U5195 (N_5195,N_320,N_2589);
nor U5196 (N_5196,N_2977,N_2531);
nand U5197 (N_5197,N_2293,N_399);
nor U5198 (N_5198,N_2058,N_1820);
or U5199 (N_5199,N_2899,N_272);
nand U5200 (N_5200,N_1168,N_313);
or U5201 (N_5201,N_1728,N_850);
and U5202 (N_5202,N_1909,N_1644);
nand U5203 (N_5203,N_2573,N_2290);
nor U5204 (N_5204,N_2593,N_2735);
and U5205 (N_5205,N_396,N_2698);
nand U5206 (N_5206,N_1917,N_2381);
and U5207 (N_5207,N_1361,N_1768);
nor U5208 (N_5208,N_1106,N_1451);
or U5209 (N_5209,N_1463,N_2552);
and U5210 (N_5210,N_256,N_561);
nand U5211 (N_5211,N_904,N_154);
and U5212 (N_5212,N_1717,N_1144);
nand U5213 (N_5213,N_2048,N_2771);
nand U5214 (N_5214,N_2296,N_377);
nand U5215 (N_5215,N_2503,N_949);
nand U5216 (N_5216,N_1656,N_739);
or U5217 (N_5217,N_2379,N_2112);
nand U5218 (N_5218,N_2293,N_556);
and U5219 (N_5219,N_2007,N_1246);
or U5220 (N_5220,N_1042,N_641);
and U5221 (N_5221,N_1282,N_2548);
nor U5222 (N_5222,N_2008,N_1703);
or U5223 (N_5223,N_2878,N_587);
nand U5224 (N_5224,N_1871,N_2483);
nand U5225 (N_5225,N_2618,N_2960);
and U5226 (N_5226,N_2524,N_2214);
nor U5227 (N_5227,N_55,N_597);
and U5228 (N_5228,N_2772,N_1604);
nand U5229 (N_5229,N_410,N_2645);
nand U5230 (N_5230,N_326,N_1398);
or U5231 (N_5231,N_225,N_2659);
or U5232 (N_5232,N_466,N_575);
xor U5233 (N_5233,N_84,N_2983);
nor U5234 (N_5234,N_1957,N_1278);
nand U5235 (N_5235,N_1750,N_640);
nor U5236 (N_5236,N_1816,N_2279);
or U5237 (N_5237,N_1239,N_771);
xor U5238 (N_5238,N_2470,N_1502);
and U5239 (N_5239,N_2494,N_529);
and U5240 (N_5240,N_1028,N_2220);
nand U5241 (N_5241,N_1392,N_667);
and U5242 (N_5242,N_930,N_1422);
or U5243 (N_5243,N_1972,N_2352);
xnor U5244 (N_5244,N_1170,N_1182);
nand U5245 (N_5245,N_2911,N_2892);
and U5246 (N_5246,N_2673,N_251);
nand U5247 (N_5247,N_594,N_2517);
xnor U5248 (N_5248,N_523,N_1136);
nand U5249 (N_5249,N_963,N_889);
xor U5250 (N_5250,N_2274,N_2216);
or U5251 (N_5251,N_2918,N_1119);
nand U5252 (N_5252,N_770,N_2228);
and U5253 (N_5253,N_935,N_141);
nor U5254 (N_5254,N_2274,N_509);
nand U5255 (N_5255,N_356,N_1727);
and U5256 (N_5256,N_2087,N_2548);
nand U5257 (N_5257,N_372,N_878);
or U5258 (N_5258,N_1161,N_2545);
and U5259 (N_5259,N_1845,N_963);
and U5260 (N_5260,N_2395,N_1922);
or U5261 (N_5261,N_1472,N_2992);
and U5262 (N_5262,N_1336,N_2181);
and U5263 (N_5263,N_2525,N_2303);
or U5264 (N_5264,N_379,N_2979);
or U5265 (N_5265,N_2254,N_87);
nor U5266 (N_5266,N_2001,N_2403);
nand U5267 (N_5267,N_727,N_2468);
or U5268 (N_5268,N_1835,N_105);
and U5269 (N_5269,N_2134,N_2296);
or U5270 (N_5270,N_225,N_2153);
nor U5271 (N_5271,N_111,N_590);
nand U5272 (N_5272,N_790,N_2087);
nor U5273 (N_5273,N_1055,N_437);
or U5274 (N_5274,N_2730,N_1733);
nand U5275 (N_5275,N_2281,N_1035);
or U5276 (N_5276,N_2081,N_325);
xor U5277 (N_5277,N_2204,N_2254);
nor U5278 (N_5278,N_2276,N_1570);
and U5279 (N_5279,N_2117,N_1402);
nor U5280 (N_5280,N_632,N_1765);
nand U5281 (N_5281,N_899,N_2326);
and U5282 (N_5282,N_1262,N_1968);
and U5283 (N_5283,N_1190,N_990);
and U5284 (N_5284,N_1125,N_1755);
nand U5285 (N_5285,N_2062,N_1777);
nand U5286 (N_5286,N_2023,N_574);
and U5287 (N_5287,N_1668,N_2405);
nor U5288 (N_5288,N_261,N_361);
or U5289 (N_5289,N_1703,N_2543);
and U5290 (N_5290,N_1889,N_2597);
nor U5291 (N_5291,N_925,N_1655);
or U5292 (N_5292,N_1234,N_682);
nor U5293 (N_5293,N_1731,N_2247);
or U5294 (N_5294,N_585,N_1727);
nand U5295 (N_5295,N_1772,N_984);
nor U5296 (N_5296,N_458,N_1428);
nand U5297 (N_5297,N_630,N_294);
and U5298 (N_5298,N_42,N_1518);
nand U5299 (N_5299,N_2593,N_0);
or U5300 (N_5300,N_885,N_1401);
or U5301 (N_5301,N_1053,N_2666);
or U5302 (N_5302,N_1340,N_1620);
nor U5303 (N_5303,N_736,N_54);
nor U5304 (N_5304,N_2400,N_1280);
nand U5305 (N_5305,N_1555,N_1297);
or U5306 (N_5306,N_216,N_1138);
nand U5307 (N_5307,N_354,N_195);
or U5308 (N_5308,N_2186,N_1508);
nand U5309 (N_5309,N_2184,N_2017);
and U5310 (N_5310,N_2274,N_2440);
nor U5311 (N_5311,N_2139,N_284);
nor U5312 (N_5312,N_719,N_12);
nor U5313 (N_5313,N_669,N_833);
xor U5314 (N_5314,N_2550,N_2238);
and U5315 (N_5315,N_40,N_646);
or U5316 (N_5316,N_2587,N_959);
nor U5317 (N_5317,N_2622,N_2434);
or U5318 (N_5318,N_327,N_1321);
nand U5319 (N_5319,N_873,N_1557);
or U5320 (N_5320,N_2647,N_2098);
or U5321 (N_5321,N_2037,N_2529);
nand U5322 (N_5322,N_2915,N_2743);
nand U5323 (N_5323,N_1538,N_760);
and U5324 (N_5324,N_2105,N_2067);
and U5325 (N_5325,N_1606,N_936);
or U5326 (N_5326,N_2035,N_2891);
nand U5327 (N_5327,N_872,N_1221);
or U5328 (N_5328,N_1881,N_338);
nor U5329 (N_5329,N_398,N_1022);
nor U5330 (N_5330,N_2192,N_2124);
or U5331 (N_5331,N_821,N_1520);
nand U5332 (N_5332,N_1470,N_1884);
or U5333 (N_5333,N_2661,N_1307);
or U5334 (N_5334,N_1587,N_119);
xor U5335 (N_5335,N_2078,N_154);
and U5336 (N_5336,N_2274,N_2979);
xnor U5337 (N_5337,N_706,N_915);
and U5338 (N_5338,N_2281,N_789);
nand U5339 (N_5339,N_1029,N_1160);
and U5340 (N_5340,N_2434,N_1007);
nor U5341 (N_5341,N_1333,N_2492);
nor U5342 (N_5342,N_2550,N_2666);
nor U5343 (N_5343,N_2330,N_89);
or U5344 (N_5344,N_2319,N_2998);
or U5345 (N_5345,N_1257,N_247);
nor U5346 (N_5346,N_669,N_2020);
nand U5347 (N_5347,N_1600,N_2859);
nor U5348 (N_5348,N_152,N_1767);
nor U5349 (N_5349,N_1499,N_2119);
and U5350 (N_5350,N_989,N_665);
nor U5351 (N_5351,N_2850,N_614);
nand U5352 (N_5352,N_2056,N_2468);
nor U5353 (N_5353,N_2356,N_2349);
nor U5354 (N_5354,N_1166,N_2837);
nand U5355 (N_5355,N_1178,N_725);
nor U5356 (N_5356,N_104,N_2767);
or U5357 (N_5357,N_2615,N_33);
or U5358 (N_5358,N_534,N_2773);
and U5359 (N_5359,N_551,N_1106);
nor U5360 (N_5360,N_1152,N_197);
and U5361 (N_5361,N_377,N_2836);
or U5362 (N_5362,N_2141,N_1064);
and U5363 (N_5363,N_1304,N_1362);
or U5364 (N_5364,N_2763,N_946);
nand U5365 (N_5365,N_344,N_268);
or U5366 (N_5366,N_1571,N_2330);
or U5367 (N_5367,N_61,N_996);
or U5368 (N_5368,N_466,N_2466);
nand U5369 (N_5369,N_577,N_864);
nor U5370 (N_5370,N_1163,N_2312);
and U5371 (N_5371,N_1256,N_2437);
nand U5372 (N_5372,N_1280,N_979);
nor U5373 (N_5373,N_1737,N_217);
or U5374 (N_5374,N_938,N_2272);
nor U5375 (N_5375,N_127,N_2328);
and U5376 (N_5376,N_2362,N_2470);
and U5377 (N_5377,N_776,N_612);
nand U5378 (N_5378,N_123,N_244);
nand U5379 (N_5379,N_1321,N_2047);
or U5380 (N_5380,N_2339,N_741);
and U5381 (N_5381,N_2127,N_1171);
or U5382 (N_5382,N_991,N_2726);
nand U5383 (N_5383,N_459,N_157);
and U5384 (N_5384,N_1810,N_1008);
nand U5385 (N_5385,N_2059,N_707);
nor U5386 (N_5386,N_1475,N_789);
and U5387 (N_5387,N_1866,N_600);
or U5388 (N_5388,N_2789,N_2364);
nand U5389 (N_5389,N_300,N_1367);
or U5390 (N_5390,N_964,N_2111);
nor U5391 (N_5391,N_2613,N_2374);
nor U5392 (N_5392,N_259,N_1075);
or U5393 (N_5393,N_2393,N_1155);
or U5394 (N_5394,N_2882,N_1557);
and U5395 (N_5395,N_2759,N_2916);
and U5396 (N_5396,N_704,N_31);
nor U5397 (N_5397,N_612,N_899);
or U5398 (N_5398,N_2268,N_156);
and U5399 (N_5399,N_1303,N_1872);
xnor U5400 (N_5400,N_667,N_2034);
and U5401 (N_5401,N_177,N_384);
and U5402 (N_5402,N_1570,N_2166);
or U5403 (N_5403,N_893,N_1047);
nand U5404 (N_5404,N_1429,N_756);
or U5405 (N_5405,N_1491,N_1227);
or U5406 (N_5406,N_1091,N_2153);
nor U5407 (N_5407,N_1973,N_1431);
and U5408 (N_5408,N_990,N_2462);
nor U5409 (N_5409,N_2087,N_34);
and U5410 (N_5410,N_856,N_2903);
nor U5411 (N_5411,N_992,N_247);
nor U5412 (N_5412,N_440,N_2017);
nor U5413 (N_5413,N_104,N_469);
nor U5414 (N_5414,N_218,N_491);
nand U5415 (N_5415,N_2310,N_1339);
and U5416 (N_5416,N_2630,N_146);
nor U5417 (N_5417,N_170,N_2584);
or U5418 (N_5418,N_2231,N_2426);
or U5419 (N_5419,N_2645,N_350);
or U5420 (N_5420,N_1361,N_816);
or U5421 (N_5421,N_2186,N_1224);
nand U5422 (N_5422,N_1901,N_994);
nand U5423 (N_5423,N_2110,N_699);
nor U5424 (N_5424,N_945,N_1604);
nor U5425 (N_5425,N_714,N_1517);
nor U5426 (N_5426,N_276,N_1262);
nor U5427 (N_5427,N_2718,N_2627);
nor U5428 (N_5428,N_1337,N_708);
nor U5429 (N_5429,N_2352,N_879);
nor U5430 (N_5430,N_315,N_623);
nand U5431 (N_5431,N_415,N_2260);
or U5432 (N_5432,N_1526,N_2404);
nor U5433 (N_5433,N_1335,N_477);
or U5434 (N_5434,N_1721,N_603);
nand U5435 (N_5435,N_1299,N_276);
nor U5436 (N_5436,N_355,N_1365);
and U5437 (N_5437,N_1102,N_1679);
or U5438 (N_5438,N_1198,N_2264);
and U5439 (N_5439,N_2777,N_1657);
nor U5440 (N_5440,N_481,N_1090);
nand U5441 (N_5441,N_1102,N_1090);
or U5442 (N_5442,N_131,N_2790);
or U5443 (N_5443,N_1452,N_1861);
nor U5444 (N_5444,N_2187,N_234);
nor U5445 (N_5445,N_1422,N_1348);
xnor U5446 (N_5446,N_2315,N_148);
nand U5447 (N_5447,N_2504,N_581);
nor U5448 (N_5448,N_2066,N_2507);
nor U5449 (N_5449,N_2007,N_2695);
nand U5450 (N_5450,N_2799,N_2947);
nand U5451 (N_5451,N_549,N_872);
nor U5452 (N_5452,N_2239,N_2039);
nor U5453 (N_5453,N_402,N_1107);
and U5454 (N_5454,N_2159,N_1308);
and U5455 (N_5455,N_1399,N_143);
nand U5456 (N_5456,N_707,N_2687);
and U5457 (N_5457,N_815,N_1770);
or U5458 (N_5458,N_659,N_2314);
or U5459 (N_5459,N_2753,N_2621);
nor U5460 (N_5460,N_17,N_2973);
and U5461 (N_5461,N_1451,N_826);
and U5462 (N_5462,N_238,N_667);
nor U5463 (N_5463,N_913,N_714);
nand U5464 (N_5464,N_1118,N_847);
or U5465 (N_5465,N_923,N_2717);
or U5466 (N_5466,N_1751,N_323);
xnor U5467 (N_5467,N_255,N_2861);
nor U5468 (N_5468,N_2515,N_2971);
or U5469 (N_5469,N_1755,N_1079);
or U5470 (N_5470,N_2301,N_1511);
nand U5471 (N_5471,N_1220,N_2520);
and U5472 (N_5472,N_661,N_1075);
nand U5473 (N_5473,N_2586,N_115);
or U5474 (N_5474,N_825,N_1590);
and U5475 (N_5475,N_2765,N_1996);
and U5476 (N_5476,N_2606,N_2132);
nor U5477 (N_5477,N_391,N_934);
or U5478 (N_5478,N_314,N_1240);
nand U5479 (N_5479,N_1486,N_1150);
nor U5480 (N_5480,N_256,N_1959);
nor U5481 (N_5481,N_2150,N_2679);
nor U5482 (N_5482,N_660,N_604);
and U5483 (N_5483,N_1255,N_67);
and U5484 (N_5484,N_450,N_1946);
or U5485 (N_5485,N_2690,N_1286);
and U5486 (N_5486,N_4,N_2231);
and U5487 (N_5487,N_2032,N_2025);
and U5488 (N_5488,N_1244,N_2828);
and U5489 (N_5489,N_2782,N_2178);
and U5490 (N_5490,N_2508,N_2784);
nand U5491 (N_5491,N_2404,N_2904);
xor U5492 (N_5492,N_322,N_1050);
or U5493 (N_5493,N_2213,N_2349);
and U5494 (N_5494,N_30,N_972);
and U5495 (N_5495,N_191,N_1178);
and U5496 (N_5496,N_1778,N_1640);
nand U5497 (N_5497,N_596,N_2197);
nor U5498 (N_5498,N_376,N_1413);
or U5499 (N_5499,N_2373,N_1511);
nand U5500 (N_5500,N_1543,N_2449);
and U5501 (N_5501,N_1903,N_1140);
or U5502 (N_5502,N_1228,N_804);
or U5503 (N_5503,N_1903,N_1828);
and U5504 (N_5504,N_2610,N_2229);
or U5505 (N_5505,N_784,N_1553);
and U5506 (N_5506,N_814,N_2192);
nand U5507 (N_5507,N_1452,N_1115);
nand U5508 (N_5508,N_413,N_1867);
or U5509 (N_5509,N_2669,N_891);
and U5510 (N_5510,N_1927,N_1304);
nand U5511 (N_5511,N_2293,N_2234);
nor U5512 (N_5512,N_2757,N_2133);
nor U5513 (N_5513,N_779,N_785);
and U5514 (N_5514,N_1250,N_2764);
or U5515 (N_5515,N_2271,N_1134);
or U5516 (N_5516,N_978,N_2484);
or U5517 (N_5517,N_2108,N_1559);
nor U5518 (N_5518,N_2614,N_2084);
or U5519 (N_5519,N_924,N_1447);
xnor U5520 (N_5520,N_1853,N_2400);
and U5521 (N_5521,N_2503,N_255);
xor U5522 (N_5522,N_517,N_85);
or U5523 (N_5523,N_2138,N_2840);
nand U5524 (N_5524,N_321,N_832);
nor U5525 (N_5525,N_2488,N_19);
nor U5526 (N_5526,N_2548,N_1337);
and U5527 (N_5527,N_649,N_1579);
nor U5528 (N_5528,N_2385,N_504);
or U5529 (N_5529,N_560,N_1428);
or U5530 (N_5530,N_1335,N_2726);
nor U5531 (N_5531,N_1809,N_914);
and U5532 (N_5532,N_2981,N_5);
and U5533 (N_5533,N_1391,N_1780);
nand U5534 (N_5534,N_2178,N_1787);
and U5535 (N_5535,N_496,N_2633);
and U5536 (N_5536,N_2467,N_396);
xor U5537 (N_5537,N_2141,N_601);
nand U5538 (N_5538,N_2834,N_79);
or U5539 (N_5539,N_1791,N_2475);
nor U5540 (N_5540,N_915,N_2611);
nor U5541 (N_5541,N_375,N_755);
nor U5542 (N_5542,N_503,N_1404);
and U5543 (N_5543,N_165,N_725);
and U5544 (N_5544,N_1983,N_1542);
nand U5545 (N_5545,N_255,N_2767);
or U5546 (N_5546,N_2987,N_1719);
nor U5547 (N_5547,N_1826,N_748);
or U5548 (N_5548,N_1602,N_2699);
nor U5549 (N_5549,N_1960,N_2734);
or U5550 (N_5550,N_535,N_2151);
nand U5551 (N_5551,N_2196,N_1589);
and U5552 (N_5552,N_795,N_2945);
nand U5553 (N_5553,N_2994,N_1758);
nor U5554 (N_5554,N_2997,N_818);
or U5555 (N_5555,N_2726,N_900);
or U5556 (N_5556,N_2023,N_1455);
or U5557 (N_5557,N_500,N_676);
nand U5558 (N_5558,N_1322,N_2914);
and U5559 (N_5559,N_2345,N_1013);
nand U5560 (N_5560,N_2361,N_2232);
nand U5561 (N_5561,N_526,N_337);
nor U5562 (N_5562,N_2352,N_432);
or U5563 (N_5563,N_280,N_499);
nand U5564 (N_5564,N_847,N_1019);
and U5565 (N_5565,N_2858,N_1644);
and U5566 (N_5566,N_1923,N_504);
nor U5567 (N_5567,N_1449,N_656);
nor U5568 (N_5568,N_396,N_1503);
or U5569 (N_5569,N_203,N_634);
or U5570 (N_5570,N_1719,N_2264);
or U5571 (N_5571,N_2604,N_858);
nand U5572 (N_5572,N_1854,N_1815);
and U5573 (N_5573,N_2516,N_165);
nand U5574 (N_5574,N_1257,N_1205);
and U5575 (N_5575,N_1498,N_1496);
nor U5576 (N_5576,N_2606,N_2519);
nor U5577 (N_5577,N_1925,N_898);
nand U5578 (N_5578,N_1086,N_1400);
or U5579 (N_5579,N_644,N_2116);
nand U5580 (N_5580,N_1092,N_2819);
nand U5581 (N_5581,N_2655,N_2450);
nand U5582 (N_5582,N_1091,N_879);
or U5583 (N_5583,N_1806,N_375);
and U5584 (N_5584,N_2237,N_2228);
nand U5585 (N_5585,N_2551,N_1940);
or U5586 (N_5586,N_621,N_1486);
and U5587 (N_5587,N_2763,N_1853);
or U5588 (N_5588,N_922,N_2978);
or U5589 (N_5589,N_571,N_1779);
nand U5590 (N_5590,N_2305,N_6);
nand U5591 (N_5591,N_1477,N_561);
or U5592 (N_5592,N_880,N_253);
nand U5593 (N_5593,N_786,N_1270);
and U5594 (N_5594,N_1715,N_141);
nand U5595 (N_5595,N_2729,N_1096);
or U5596 (N_5596,N_2542,N_1064);
nor U5597 (N_5597,N_1795,N_1681);
and U5598 (N_5598,N_2812,N_2453);
nor U5599 (N_5599,N_2228,N_180);
or U5600 (N_5600,N_1399,N_1449);
and U5601 (N_5601,N_1553,N_1752);
nor U5602 (N_5602,N_286,N_1260);
nor U5603 (N_5603,N_1116,N_1286);
nand U5604 (N_5604,N_142,N_1250);
nor U5605 (N_5605,N_1333,N_2660);
and U5606 (N_5606,N_433,N_813);
and U5607 (N_5607,N_2423,N_1598);
and U5608 (N_5608,N_367,N_1524);
nand U5609 (N_5609,N_121,N_2693);
nand U5610 (N_5610,N_1080,N_2762);
and U5611 (N_5611,N_1204,N_2281);
and U5612 (N_5612,N_2114,N_2041);
or U5613 (N_5613,N_1360,N_1323);
or U5614 (N_5614,N_2379,N_2591);
nor U5615 (N_5615,N_1619,N_44);
and U5616 (N_5616,N_2367,N_1051);
nor U5617 (N_5617,N_2117,N_513);
and U5618 (N_5618,N_616,N_970);
and U5619 (N_5619,N_728,N_1698);
or U5620 (N_5620,N_1730,N_179);
nor U5621 (N_5621,N_1965,N_646);
nor U5622 (N_5622,N_1242,N_1381);
and U5623 (N_5623,N_2909,N_2821);
nor U5624 (N_5624,N_2651,N_2773);
or U5625 (N_5625,N_1647,N_1628);
and U5626 (N_5626,N_2379,N_102);
nand U5627 (N_5627,N_1013,N_125);
and U5628 (N_5628,N_1331,N_73);
and U5629 (N_5629,N_1209,N_988);
and U5630 (N_5630,N_762,N_2394);
or U5631 (N_5631,N_892,N_165);
and U5632 (N_5632,N_673,N_1217);
nor U5633 (N_5633,N_694,N_463);
nor U5634 (N_5634,N_911,N_1319);
xnor U5635 (N_5635,N_1768,N_1626);
nand U5636 (N_5636,N_216,N_1364);
nand U5637 (N_5637,N_15,N_1116);
or U5638 (N_5638,N_2628,N_2337);
and U5639 (N_5639,N_796,N_2289);
nand U5640 (N_5640,N_771,N_284);
or U5641 (N_5641,N_705,N_2847);
or U5642 (N_5642,N_1013,N_2671);
or U5643 (N_5643,N_2981,N_2644);
or U5644 (N_5644,N_258,N_1441);
or U5645 (N_5645,N_1545,N_2083);
or U5646 (N_5646,N_678,N_1171);
or U5647 (N_5647,N_847,N_1446);
nor U5648 (N_5648,N_1514,N_2898);
nor U5649 (N_5649,N_1516,N_527);
and U5650 (N_5650,N_2774,N_995);
and U5651 (N_5651,N_1953,N_1926);
nand U5652 (N_5652,N_990,N_1694);
nand U5653 (N_5653,N_602,N_823);
nor U5654 (N_5654,N_820,N_277);
nor U5655 (N_5655,N_1060,N_232);
or U5656 (N_5656,N_2634,N_1060);
and U5657 (N_5657,N_2517,N_1635);
and U5658 (N_5658,N_2532,N_309);
nand U5659 (N_5659,N_2983,N_121);
and U5660 (N_5660,N_264,N_820);
and U5661 (N_5661,N_2109,N_2911);
nor U5662 (N_5662,N_2831,N_1904);
nand U5663 (N_5663,N_1038,N_413);
nor U5664 (N_5664,N_1005,N_1491);
nor U5665 (N_5665,N_1527,N_2453);
or U5666 (N_5666,N_2608,N_2995);
nor U5667 (N_5667,N_1416,N_542);
and U5668 (N_5668,N_2813,N_2075);
or U5669 (N_5669,N_3,N_2666);
nand U5670 (N_5670,N_821,N_281);
nor U5671 (N_5671,N_1727,N_1730);
and U5672 (N_5672,N_1103,N_1597);
and U5673 (N_5673,N_2730,N_1447);
xnor U5674 (N_5674,N_2039,N_2626);
nor U5675 (N_5675,N_823,N_312);
nand U5676 (N_5676,N_2429,N_2924);
nand U5677 (N_5677,N_715,N_2375);
nand U5678 (N_5678,N_1417,N_2229);
nand U5679 (N_5679,N_2508,N_2732);
nand U5680 (N_5680,N_1280,N_1685);
nor U5681 (N_5681,N_613,N_2385);
or U5682 (N_5682,N_621,N_2839);
and U5683 (N_5683,N_950,N_2619);
or U5684 (N_5684,N_955,N_639);
nand U5685 (N_5685,N_839,N_993);
or U5686 (N_5686,N_2563,N_2777);
or U5687 (N_5687,N_2236,N_1955);
and U5688 (N_5688,N_233,N_867);
nor U5689 (N_5689,N_1604,N_1150);
nor U5690 (N_5690,N_747,N_2704);
nand U5691 (N_5691,N_1575,N_2511);
nand U5692 (N_5692,N_966,N_2927);
or U5693 (N_5693,N_1090,N_239);
or U5694 (N_5694,N_654,N_1485);
and U5695 (N_5695,N_2350,N_2212);
nand U5696 (N_5696,N_2297,N_190);
nand U5697 (N_5697,N_2003,N_64);
nand U5698 (N_5698,N_570,N_1105);
and U5699 (N_5699,N_1649,N_1629);
and U5700 (N_5700,N_577,N_1806);
nor U5701 (N_5701,N_195,N_470);
or U5702 (N_5702,N_1371,N_2357);
or U5703 (N_5703,N_2660,N_1671);
and U5704 (N_5704,N_1047,N_1396);
or U5705 (N_5705,N_1417,N_1094);
nand U5706 (N_5706,N_1331,N_2721);
nor U5707 (N_5707,N_389,N_898);
nand U5708 (N_5708,N_2448,N_1956);
and U5709 (N_5709,N_2292,N_1468);
and U5710 (N_5710,N_1579,N_2516);
or U5711 (N_5711,N_339,N_2565);
nor U5712 (N_5712,N_6,N_1142);
nand U5713 (N_5713,N_2190,N_16);
and U5714 (N_5714,N_1312,N_2972);
nand U5715 (N_5715,N_1942,N_2943);
or U5716 (N_5716,N_569,N_2132);
or U5717 (N_5717,N_32,N_1792);
nand U5718 (N_5718,N_396,N_483);
and U5719 (N_5719,N_2248,N_374);
and U5720 (N_5720,N_2352,N_1138);
nor U5721 (N_5721,N_347,N_112);
nand U5722 (N_5722,N_2047,N_2173);
nor U5723 (N_5723,N_2516,N_2230);
and U5724 (N_5724,N_1676,N_1599);
and U5725 (N_5725,N_1285,N_2906);
nor U5726 (N_5726,N_2129,N_1669);
nand U5727 (N_5727,N_854,N_1367);
nand U5728 (N_5728,N_2872,N_2129);
xor U5729 (N_5729,N_749,N_2188);
or U5730 (N_5730,N_1253,N_2968);
nor U5731 (N_5731,N_2535,N_2530);
and U5732 (N_5732,N_2258,N_1714);
or U5733 (N_5733,N_1772,N_1833);
and U5734 (N_5734,N_788,N_1019);
and U5735 (N_5735,N_2358,N_1595);
nor U5736 (N_5736,N_2608,N_2434);
nand U5737 (N_5737,N_2827,N_96);
nand U5738 (N_5738,N_1530,N_386);
nand U5739 (N_5739,N_485,N_1408);
nor U5740 (N_5740,N_426,N_353);
or U5741 (N_5741,N_588,N_723);
or U5742 (N_5742,N_2302,N_1298);
and U5743 (N_5743,N_26,N_2755);
nor U5744 (N_5744,N_679,N_1852);
and U5745 (N_5745,N_506,N_939);
or U5746 (N_5746,N_1540,N_215);
nand U5747 (N_5747,N_859,N_1629);
or U5748 (N_5748,N_1107,N_2162);
nand U5749 (N_5749,N_1855,N_1899);
or U5750 (N_5750,N_919,N_2758);
or U5751 (N_5751,N_630,N_580);
nand U5752 (N_5752,N_2259,N_1277);
nor U5753 (N_5753,N_245,N_243);
nor U5754 (N_5754,N_1108,N_2506);
or U5755 (N_5755,N_212,N_1107);
nand U5756 (N_5756,N_2364,N_1328);
nor U5757 (N_5757,N_1225,N_2390);
nand U5758 (N_5758,N_485,N_1009);
or U5759 (N_5759,N_98,N_166);
and U5760 (N_5760,N_2496,N_863);
nor U5761 (N_5761,N_704,N_590);
nand U5762 (N_5762,N_2234,N_2926);
nand U5763 (N_5763,N_2269,N_2889);
and U5764 (N_5764,N_622,N_1897);
nor U5765 (N_5765,N_1436,N_2882);
nor U5766 (N_5766,N_2592,N_809);
and U5767 (N_5767,N_2174,N_1939);
and U5768 (N_5768,N_2095,N_53);
nand U5769 (N_5769,N_1059,N_953);
and U5770 (N_5770,N_216,N_937);
or U5771 (N_5771,N_997,N_1901);
nand U5772 (N_5772,N_2526,N_2724);
nor U5773 (N_5773,N_1480,N_2457);
xor U5774 (N_5774,N_2848,N_78);
nor U5775 (N_5775,N_409,N_2554);
nand U5776 (N_5776,N_1245,N_278);
nor U5777 (N_5777,N_1957,N_891);
and U5778 (N_5778,N_148,N_2720);
and U5779 (N_5779,N_2010,N_1007);
nand U5780 (N_5780,N_368,N_2241);
nand U5781 (N_5781,N_62,N_2823);
nor U5782 (N_5782,N_2349,N_299);
and U5783 (N_5783,N_424,N_930);
and U5784 (N_5784,N_999,N_1205);
nor U5785 (N_5785,N_908,N_1241);
nand U5786 (N_5786,N_348,N_178);
nand U5787 (N_5787,N_2859,N_1120);
and U5788 (N_5788,N_527,N_1072);
nor U5789 (N_5789,N_2676,N_175);
nand U5790 (N_5790,N_2881,N_2214);
xnor U5791 (N_5791,N_2780,N_147);
or U5792 (N_5792,N_1688,N_2487);
and U5793 (N_5793,N_1763,N_273);
or U5794 (N_5794,N_1037,N_1176);
nand U5795 (N_5795,N_301,N_1562);
nand U5796 (N_5796,N_2370,N_2884);
nor U5797 (N_5797,N_1779,N_1560);
or U5798 (N_5798,N_2483,N_1525);
xnor U5799 (N_5799,N_2771,N_265);
xor U5800 (N_5800,N_1164,N_973);
or U5801 (N_5801,N_635,N_1925);
or U5802 (N_5802,N_1820,N_561);
and U5803 (N_5803,N_278,N_84);
or U5804 (N_5804,N_2273,N_2188);
or U5805 (N_5805,N_1300,N_1355);
or U5806 (N_5806,N_2907,N_118);
or U5807 (N_5807,N_806,N_1917);
and U5808 (N_5808,N_2379,N_1813);
and U5809 (N_5809,N_2598,N_2376);
nand U5810 (N_5810,N_126,N_1762);
and U5811 (N_5811,N_1674,N_2267);
or U5812 (N_5812,N_1615,N_1635);
nand U5813 (N_5813,N_2992,N_2759);
or U5814 (N_5814,N_2667,N_712);
and U5815 (N_5815,N_1977,N_1328);
or U5816 (N_5816,N_2300,N_2551);
and U5817 (N_5817,N_539,N_2139);
nor U5818 (N_5818,N_1965,N_108);
nor U5819 (N_5819,N_1968,N_1052);
or U5820 (N_5820,N_2912,N_2147);
nor U5821 (N_5821,N_11,N_1161);
and U5822 (N_5822,N_2864,N_2441);
and U5823 (N_5823,N_866,N_1914);
and U5824 (N_5824,N_1370,N_1513);
and U5825 (N_5825,N_682,N_926);
or U5826 (N_5826,N_637,N_1165);
nor U5827 (N_5827,N_1676,N_463);
nor U5828 (N_5828,N_586,N_132);
xor U5829 (N_5829,N_1330,N_48);
nor U5830 (N_5830,N_1985,N_2483);
or U5831 (N_5831,N_550,N_1725);
or U5832 (N_5832,N_2962,N_2478);
nand U5833 (N_5833,N_2263,N_2833);
or U5834 (N_5834,N_1989,N_215);
nand U5835 (N_5835,N_2358,N_2122);
or U5836 (N_5836,N_1797,N_938);
nor U5837 (N_5837,N_92,N_2066);
or U5838 (N_5838,N_2448,N_2149);
and U5839 (N_5839,N_729,N_1979);
and U5840 (N_5840,N_713,N_1817);
nor U5841 (N_5841,N_2589,N_1618);
and U5842 (N_5842,N_1316,N_2034);
nor U5843 (N_5843,N_471,N_645);
nor U5844 (N_5844,N_1077,N_2279);
nor U5845 (N_5845,N_88,N_2015);
and U5846 (N_5846,N_2102,N_2115);
nor U5847 (N_5847,N_748,N_1331);
or U5848 (N_5848,N_1469,N_957);
or U5849 (N_5849,N_787,N_1000);
nor U5850 (N_5850,N_1889,N_1782);
and U5851 (N_5851,N_992,N_1758);
nand U5852 (N_5852,N_331,N_2479);
or U5853 (N_5853,N_50,N_279);
nor U5854 (N_5854,N_276,N_403);
nand U5855 (N_5855,N_427,N_895);
and U5856 (N_5856,N_1354,N_2091);
nand U5857 (N_5857,N_1775,N_2756);
xnor U5858 (N_5858,N_591,N_1904);
and U5859 (N_5859,N_2540,N_1478);
nor U5860 (N_5860,N_1952,N_1304);
nor U5861 (N_5861,N_2711,N_1239);
and U5862 (N_5862,N_375,N_87);
nand U5863 (N_5863,N_2006,N_847);
or U5864 (N_5864,N_1095,N_2037);
and U5865 (N_5865,N_2176,N_1167);
nor U5866 (N_5866,N_1297,N_2206);
nor U5867 (N_5867,N_622,N_2620);
and U5868 (N_5868,N_461,N_81);
or U5869 (N_5869,N_1614,N_891);
nand U5870 (N_5870,N_2716,N_1988);
or U5871 (N_5871,N_2529,N_2586);
nor U5872 (N_5872,N_1546,N_773);
nor U5873 (N_5873,N_1262,N_1324);
and U5874 (N_5874,N_54,N_909);
nor U5875 (N_5875,N_848,N_981);
and U5876 (N_5876,N_1201,N_2098);
nand U5877 (N_5877,N_1352,N_1488);
nor U5878 (N_5878,N_1595,N_700);
nand U5879 (N_5879,N_1205,N_2804);
nand U5880 (N_5880,N_71,N_355);
nand U5881 (N_5881,N_2547,N_1716);
or U5882 (N_5882,N_1887,N_1078);
nor U5883 (N_5883,N_1253,N_1854);
nor U5884 (N_5884,N_732,N_108);
nand U5885 (N_5885,N_859,N_139);
xnor U5886 (N_5886,N_1087,N_1019);
nand U5887 (N_5887,N_986,N_2559);
and U5888 (N_5888,N_935,N_287);
nor U5889 (N_5889,N_2821,N_1798);
and U5890 (N_5890,N_2192,N_2733);
or U5891 (N_5891,N_1175,N_2373);
nor U5892 (N_5892,N_904,N_1806);
nand U5893 (N_5893,N_1921,N_976);
nand U5894 (N_5894,N_2760,N_1940);
and U5895 (N_5895,N_2434,N_2187);
nor U5896 (N_5896,N_685,N_2843);
nor U5897 (N_5897,N_303,N_2037);
or U5898 (N_5898,N_2145,N_2790);
and U5899 (N_5899,N_2387,N_2688);
nor U5900 (N_5900,N_362,N_1660);
or U5901 (N_5901,N_2177,N_1631);
or U5902 (N_5902,N_352,N_1913);
and U5903 (N_5903,N_2104,N_929);
or U5904 (N_5904,N_236,N_2930);
nand U5905 (N_5905,N_323,N_2314);
or U5906 (N_5906,N_2980,N_562);
and U5907 (N_5907,N_2296,N_1188);
and U5908 (N_5908,N_2576,N_2245);
nand U5909 (N_5909,N_1943,N_2371);
or U5910 (N_5910,N_2200,N_2086);
nand U5911 (N_5911,N_28,N_2562);
nor U5912 (N_5912,N_388,N_1725);
nor U5913 (N_5913,N_2331,N_2290);
or U5914 (N_5914,N_1013,N_248);
nor U5915 (N_5915,N_1748,N_960);
nand U5916 (N_5916,N_436,N_2222);
nor U5917 (N_5917,N_1624,N_72);
and U5918 (N_5918,N_2387,N_1036);
nand U5919 (N_5919,N_675,N_1556);
nand U5920 (N_5920,N_867,N_2473);
or U5921 (N_5921,N_1831,N_2154);
nor U5922 (N_5922,N_1434,N_1404);
xor U5923 (N_5923,N_36,N_486);
xor U5924 (N_5924,N_1698,N_995);
nor U5925 (N_5925,N_2863,N_2839);
or U5926 (N_5926,N_2055,N_349);
nand U5927 (N_5927,N_1175,N_1482);
xnor U5928 (N_5928,N_2326,N_485);
and U5929 (N_5929,N_2505,N_2486);
nor U5930 (N_5930,N_369,N_846);
or U5931 (N_5931,N_450,N_1181);
and U5932 (N_5932,N_1952,N_567);
nor U5933 (N_5933,N_2180,N_2757);
nand U5934 (N_5934,N_732,N_2836);
nor U5935 (N_5935,N_896,N_136);
and U5936 (N_5936,N_474,N_74);
nor U5937 (N_5937,N_300,N_1402);
and U5938 (N_5938,N_2269,N_2159);
and U5939 (N_5939,N_2498,N_895);
nor U5940 (N_5940,N_717,N_852);
nor U5941 (N_5941,N_739,N_889);
nor U5942 (N_5942,N_2167,N_251);
and U5943 (N_5943,N_2163,N_1837);
nor U5944 (N_5944,N_2396,N_2046);
or U5945 (N_5945,N_35,N_238);
nand U5946 (N_5946,N_891,N_1324);
nand U5947 (N_5947,N_2511,N_2005);
or U5948 (N_5948,N_1381,N_1096);
nor U5949 (N_5949,N_61,N_2507);
nor U5950 (N_5950,N_1603,N_2680);
nand U5951 (N_5951,N_290,N_674);
nand U5952 (N_5952,N_954,N_2316);
nor U5953 (N_5953,N_884,N_76);
nand U5954 (N_5954,N_855,N_2003);
nor U5955 (N_5955,N_2585,N_1109);
and U5956 (N_5956,N_524,N_1150);
nand U5957 (N_5957,N_1483,N_1363);
nor U5958 (N_5958,N_2802,N_1448);
nor U5959 (N_5959,N_1220,N_2189);
and U5960 (N_5960,N_1797,N_2607);
or U5961 (N_5961,N_2721,N_2751);
or U5962 (N_5962,N_2111,N_957);
nand U5963 (N_5963,N_2927,N_1072);
or U5964 (N_5964,N_2980,N_1126);
and U5965 (N_5965,N_2443,N_1726);
and U5966 (N_5966,N_1706,N_1551);
or U5967 (N_5967,N_2395,N_775);
nor U5968 (N_5968,N_586,N_1539);
and U5969 (N_5969,N_893,N_396);
or U5970 (N_5970,N_654,N_2031);
or U5971 (N_5971,N_316,N_1015);
and U5972 (N_5972,N_1719,N_2611);
nor U5973 (N_5973,N_2913,N_1625);
or U5974 (N_5974,N_1353,N_2532);
or U5975 (N_5975,N_163,N_1548);
nand U5976 (N_5976,N_1332,N_2591);
and U5977 (N_5977,N_1039,N_2037);
and U5978 (N_5978,N_2833,N_2534);
xor U5979 (N_5979,N_1995,N_2749);
nand U5980 (N_5980,N_728,N_635);
nand U5981 (N_5981,N_178,N_968);
or U5982 (N_5982,N_1725,N_1031);
or U5983 (N_5983,N_2151,N_1605);
and U5984 (N_5984,N_882,N_1577);
nor U5985 (N_5985,N_1852,N_2757);
and U5986 (N_5986,N_1891,N_1490);
or U5987 (N_5987,N_393,N_1508);
nor U5988 (N_5988,N_797,N_706);
and U5989 (N_5989,N_2943,N_1915);
or U5990 (N_5990,N_92,N_1615);
nand U5991 (N_5991,N_2596,N_2156);
xnor U5992 (N_5992,N_618,N_2155);
and U5993 (N_5993,N_1235,N_1156);
nand U5994 (N_5994,N_2317,N_1249);
nand U5995 (N_5995,N_1452,N_80);
and U5996 (N_5996,N_232,N_1175);
nand U5997 (N_5997,N_436,N_2264);
and U5998 (N_5998,N_2114,N_93);
nand U5999 (N_5999,N_1407,N_466);
or U6000 (N_6000,N_5605,N_5272);
or U6001 (N_6001,N_3886,N_3083);
nand U6002 (N_6002,N_4014,N_3281);
nor U6003 (N_6003,N_3158,N_5607);
and U6004 (N_6004,N_3800,N_5449);
or U6005 (N_6005,N_4740,N_5353);
and U6006 (N_6006,N_5107,N_4353);
nor U6007 (N_6007,N_4366,N_3374);
and U6008 (N_6008,N_5046,N_4526);
nor U6009 (N_6009,N_4576,N_3557);
nand U6010 (N_6010,N_3108,N_5079);
nand U6011 (N_6011,N_4351,N_3353);
and U6012 (N_6012,N_5524,N_4896);
nor U6013 (N_6013,N_4993,N_3975);
nor U6014 (N_6014,N_5385,N_3348);
or U6015 (N_6015,N_4385,N_3872);
nand U6016 (N_6016,N_4204,N_4399);
or U6017 (N_6017,N_3604,N_4037);
nand U6018 (N_6018,N_5369,N_3571);
or U6019 (N_6019,N_3031,N_4857);
nand U6020 (N_6020,N_3069,N_3330);
and U6021 (N_6021,N_3350,N_4965);
and U6022 (N_6022,N_5039,N_5878);
or U6023 (N_6023,N_3465,N_3251);
nor U6024 (N_6024,N_5440,N_4061);
nand U6025 (N_6025,N_3779,N_5806);
nor U6026 (N_6026,N_3665,N_4550);
nand U6027 (N_6027,N_5137,N_3971);
nor U6028 (N_6028,N_5451,N_4003);
nor U6029 (N_6029,N_3494,N_3169);
and U6030 (N_6030,N_5196,N_3153);
and U6031 (N_6031,N_4442,N_4391);
xnor U6032 (N_6032,N_3848,N_4678);
nand U6033 (N_6033,N_3984,N_3220);
and U6034 (N_6034,N_3061,N_3492);
or U6035 (N_6035,N_5366,N_3462);
nor U6036 (N_6036,N_5742,N_5185);
or U6037 (N_6037,N_5638,N_4540);
xnor U6038 (N_6038,N_3898,N_5627);
nor U6039 (N_6039,N_5651,N_3004);
nand U6040 (N_6040,N_5811,N_3088);
or U6041 (N_6041,N_5916,N_5781);
or U6042 (N_6042,N_4105,N_4631);
nand U6043 (N_6043,N_4541,N_5795);
nand U6044 (N_6044,N_4790,N_3005);
or U6045 (N_6045,N_4510,N_3894);
and U6046 (N_6046,N_5175,N_5677);
nand U6047 (N_6047,N_4024,N_4575);
and U6048 (N_6048,N_4245,N_4131);
nand U6049 (N_6049,N_3122,N_4788);
or U6050 (N_6050,N_4411,N_3424);
or U6051 (N_6051,N_4592,N_3545);
or U6052 (N_6052,N_3786,N_3246);
or U6053 (N_6053,N_4444,N_4318);
nand U6054 (N_6054,N_3086,N_3548);
xor U6055 (N_6055,N_5427,N_4546);
nand U6056 (N_6056,N_4607,N_3946);
or U6057 (N_6057,N_5955,N_4109);
nand U6058 (N_6058,N_4641,N_4943);
and U6059 (N_6059,N_5303,N_4899);
or U6060 (N_6060,N_4213,N_4590);
and U6061 (N_6061,N_3039,N_3645);
nand U6062 (N_6062,N_3318,N_3321);
nor U6063 (N_6063,N_5410,N_4012);
nand U6064 (N_6064,N_3751,N_3923);
nor U6065 (N_6065,N_3202,N_5585);
nor U6066 (N_6066,N_5267,N_4230);
nor U6067 (N_6067,N_3904,N_5249);
xnor U6068 (N_6068,N_4143,N_4598);
and U6069 (N_6069,N_3412,N_5172);
nand U6070 (N_6070,N_3680,N_5764);
or U6071 (N_6071,N_5662,N_3369);
nand U6072 (N_6072,N_3835,N_4202);
or U6073 (N_6073,N_3326,N_5756);
nand U6074 (N_6074,N_3160,N_3688);
or U6075 (N_6075,N_3407,N_3147);
nand U6076 (N_6076,N_3953,N_4949);
and U6077 (N_6077,N_5074,N_4916);
nand U6078 (N_6078,N_5115,N_5981);
and U6079 (N_6079,N_4505,N_5056);
nand U6080 (N_6080,N_4936,N_3782);
nor U6081 (N_6081,N_4897,N_5459);
or U6082 (N_6082,N_5120,N_5329);
or U6083 (N_6083,N_3903,N_4272);
nor U6084 (N_6084,N_3881,N_4404);
xnor U6085 (N_6085,N_4597,N_5094);
and U6086 (N_6086,N_3466,N_3634);
and U6087 (N_6087,N_3217,N_5332);
nand U6088 (N_6088,N_5821,N_5346);
nor U6089 (N_6089,N_4359,N_5494);
and U6090 (N_6090,N_4049,N_4218);
or U6091 (N_6091,N_4725,N_5921);
nand U6092 (N_6092,N_4201,N_4043);
or U6093 (N_6093,N_5340,N_5684);
nor U6094 (N_6094,N_5579,N_4729);
nand U6095 (N_6095,N_4470,N_5118);
and U6096 (N_6096,N_3935,N_3385);
xor U6097 (N_6097,N_5264,N_3780);
xnor U6098 (N_6098,N_4847,N_4853);
or U6099 (N_6099,N_4950,N_3105);
and U6100 (N_6100,N_5371,N_4026);
xnor U6101 (N_6101,N_4461,N_4246);
nand U6102 (N_6102,N_4700,N_5370);
nand U6103 (N_6103,N_3519,N_4591);
or U6104 (N_6104,N_5481,N_4117);
nand U6105 (N_6105,N_5802,N_5723);
and U6106 (N_6106,N_3674,N_3499);
nor U6107 (N_6107,N_3416,N_4080);
nor U6108 (N_6108,N_5626,N_3832);
nor U6109 (N_6109,N_3197,N_5113);
nor U6110 (N_6110,N_5296,N_3533);
xnor U6111 (N_6111,N_4651,N_4255);
and U6112 (N_6112,N_3829,N_3491);
nor U6113 (N_6113,N_3698,N_3440);
nor U6114 (N_6114,N_5472,N_5152);
or U6115 (N_6115,N_4119,N_3066);
nand U6116 (N_6116,N_4009,N_5500);
nor U6117 (N_6117,N_3743,N_4179);
nor U6118 (N_6118,N_5206,N_5289);
or U6119 (N_6119,N_5349,N_4984);
or U6120 (N_6120,N_4138,N_3672);
and U6121 (N_6121,N_5038,N_5636);
or U6122 (N_6122,N_3482,N_4711);
or U6123 (N_6123,N_3431,N_3776);
nand U6124 (N_6124,N_3945,N_4284);
and U6125 (N_6125,N_5474,N_3297);
nand U6126 (N_6126,N_4969,N_3697);
and U6127 (N_6127,N_4091,N_5401);
nand U6128 (N_6128,N_5694,N_4452);
and U6129 (N_6129,N_5194,N_3589);
or U6130 (N_6130,N_3359,N_3397);
and U6131 (N_6131,N_5142,N_5344);
xor U6132 (N_6132,N_4587,N_5754);
and U6133 (N_6133,N_4483,N_5839);
and U6134 (N_6134,N_3419,N_5750);
nor U6135 (N_6135,N_5455,N_5442);
or U6136 (N_6136,N_3370,N_5300);
xor U6137 (N_6137,N_5621,N_3728);
nand U6138 (N_6138,N_5693,N_3826);
or U6139 (N_6139,N_4384,N_4823);
nand U6140 (N_6140,N_4212,N_3902);
nand U6141 (N_6141,N_3418,N_5940);
nor U6142 (N_6142,N_5884,N_5661);
and U6143 (N_6143,N_3346,N_3542);
nand U6144 (N_6144,N_5531,N_3806);
nor U6145 (N_6145,N_5925,N_5260);
and U6146 (N_6146,N_4277,N_4660);
nand U6147 (N_6147,N_5796,N_3855);
nor U6148 (N_6148,N_4044,N_4970);
nand U6149 (N_6149,N_4333,N_5555);
nor U6150 (N_6150,N_4456,N_4234);
and U6151 (N_6151,N_5944,N_4369);
nand U6152 (N_6152,N_4240,N_4273);
nand U6153 (N_6153,N_5527,N_5520);
nor U6154 (N_6154,N_5514,N_3067);
or U6155 (N_6155,N_3243,N_5497);
and U6156 (N_6156,N_4098,N_3534);
nor U6157 (N_6157,N_5648,N_5470);
or U6158 (N_6158,N_3444,N_5829);
nand U6159 (N_6159,N_3304,N_3613);
nand U6160 (N_6160,N_3390,N_3831);
or U6161 (N_6161,N_5019,N_3130);
xor U6162 (N_6162,N_4635,N_4382);
nor U6163 (N_6163,N_5012,N_4567);
nor U6164 (N_6164,N_5013,N_4599);
or U6165 (N_6165,N_5911,N_5571);
nor U6166 (N_6166,N_4948,N_3183);
nand U6167 (N_6167,N_5215,N_3659);
and U6168 (N_6168,N_5178,N_3159);
nand U6169 (N_6169,N_5269,N_5667);
nor U6170 (N_6170,N_5951,N_5904);
xnor U6171 (N_6171,N_4642,N_3964);
or U6172 (N_6172,N_3576,N_3460);
xor U6173 (N_6173,N_5515,N_3819);
and U6174 (N_6174,N_4545,N_4945);
and U6175 (N_6175,N_5771,N_4862);
nor U6176 (N_6176,N_4926,N_3033);
nor U6177 (N_6177,N_5256,N_5328);
nand U6178 (N_6178,N_5659,N_3085);
or U6179 (N_6179,N_4543,N_5225);
and U6180 (N_6180,N_4895,N_4454);
nand U6181 (N_6181,N_3023,N_4270);
or U6182 (N_6182,N_4403,N_4961);
or U6183 (N_6183,N_4187,N_3034);
and U6184 (N_6184,N_5982,N_3907);
nand U6185 (N_6185,N_4754,N_3739);
or U6186 (N_6186,N_3549,N_5564);
nor U6187 (N_6187,N_5772,N_5299);
or U6188 (N_6188,N_4923,N_4900);
or U6189 (N_6189,N_5584,N_5241);
nor U6190 (N_6190,N_5570,N_5156);
nand U6191 (N_6191,N_3137,N_5054);
and U6192 (N_6192,N_5526,N_5498);
nor U6193 (N_6193,N_4983,N_3750);
or U6194 (N_6194,N_5546,N_3495);
nor U6195 (N_6195,N_4652,N_4077);
and U6196 (N_6196,N_4718,N_5861);
nand U6197 (N_6197,N_3653,N_5587);
or U6198 (N_6198,N_3524,N_4289);
and U6199 (N_6199,N_4643,N_4428);
nand U6200 (N_6200,N_3675,N_3591);
nor U6201 (N_6201,N_3203,N_5236);
nor U6202 (N_6202,N_3165,N_3386);
and U6203 (N_6203,N_5624,N_5834);
or U6204 (N_6204,N_4458,N_4374);
or U6205 (N_6205,N_3300,N_5832);
or U6206 (N_6206,N_3565,N_3252);
or U6207 (N_6207,N_4523,N_3154);
or U6208 (N_6208,N_4209,N_5434);
or U6209 (N_6209,N_3741,N_4615);
nand U6210 (N_6210,N_5288,N_5489);
or U6211 (N_6211,N_4683,N_3025);
nor U6212 (N_6212,N_4102,N_4023);
nand U6213 (N_6213,N_4028,N_5209);
or U6214 (N_6214,N_5454,N_4267);
or U6215 (N_6215,N_4311,N_4247);
or U6216 (N_6216,N_3996,N_3999);
nand U6217 (N_6217,N_4140,N_3809);
xor U6218 (N_6218,N_4379,N_3535);
nand U6219 (N_6219,N_4219,N_3011);
nor U6220 (N_6220,N_3422,N_5704);
or U6221 (N_6221,N_5024,N_5250);
nand U6222 (N_6222,N_5210,N_5511);
nor U6223 (N_6223,N_3291,N_5422);
nand U6224 (N_6224,N_3009,N_3262);
nor U6225 (N_6225,N_5941,N_3423);
nand U6226 (N_6226,N_5809,N_5485);
nand U6227 (N_6227,N_4464,N_5907);
and U6228 (N_6228,N_5167,N_4947);
and U6229 (N_6229,N_4530,N_4763);
nor U6230 (N_6230,N_3354,N_5827);
nor U6231 (N_6231,N_4820,N_5943);
or U6232 (N_6232,N_5510,N_5186);
and U6233 (N_6233,N_5402,N_5559);
or U6234 (N_6234,N_5622,N_5998);
nand U6235 (N_6235,N_5613,N_5864);
nand U6236 (N_6236,N_3897,N_3815);
nand U6237 (N_6237,N_3884,N_5432);
nor U6238 (N_6238,N_3598,N_4256);
nor U6239 (N_6239,N_4376,N_5453);
nand U6240 (N_6240,N_3581,N_5599);
and U6241 (N_6241,N_3406,N_3471);
and U6242 (N_6242,N_4180,N_4063);
and U6243 (N_6243,N_5352,N_4223);
xnor U6244 (N_6244,N_5357,N_3379);
xnor U6245 (N_6245,N_3400,N_4345);
nand U6246 (N_6246,N_3569,N_4739);
and U6247 (N_6247,N_5810,N_3112);
and U6248 (N_6248,N_3226,N_5934);
nand U6249 (N_6249,N_5135,N_3630);
nand U6250 (N_6250,N_5297,N_3433);
xor U6251 (N_6251,N_5676,N_4364);
or U6252 (N_6252,N_4360,N_5244);
and U6253 (N_6253,N_5088,N_4322);
xnor U6254 (N_6254,N_3028,N_3849);
nor U6255 (N_6255,N_4835,N_3455);
and U6256 (N_6256,N_5950,N_4441);
nor U6257 (N_6257,N_3794,N_4685);
or U6258 (N_6258,N_3677,N_4735);
and U6259 (N_6259,N_4697,N_3237);
or U6260 (N_6260,N_4482,N_4446);
or U6261 (N_6261,N_3081,N_5116);
or U6262 (N_6262,N_3518,N_5538);
or U6263 (N_6263,N_5100,N_5695);
xor U6264 (N_6264,N_4626,N_5128);
nor U6265 (N_6265,N_3955,N_3839);
or U6266 (N_6266,N_5174,N_3525);
nor U6267 (N_6267,N_4922,N_5252);
and U6268 (N_6268,N_3956,N_4988);
or U6269 (N_6269,N_4327,N_3991);
nor U6270 (N_6270,N_5713,N_3489);
nand U6271 (N_6271,N_5799,N_3432);
and U6272 (N_6272,N_3893,N_3757);
nor U6273 (N_6273,N_4000,N_5032);
nand U6274 (N_6274,N_5224,N_3944);
nor U6275 (N_6275,N_3436,N_4815);
or U6276 (N_6276,N_5376,N_4166);
nor U6277 (N_6277,N_5708,N_3684);
or U6278 (N_6278,N_4604,N_5285);
nor U6279 (N_6279,N_3487,N_4455);
and U6280 (N_6280,N_4930,N_3836);
nand U6281 (N_6281,N_4509,N_5807);
nand U6282 (N_6282,N_3622,N_4648);
nor U6283 (N_6283,N_4216,N_5231);
nand U6284 (N_6284,N_5488,N_3452);
nor U6285 (N_6285,N_4554,N_5658);
or U6286 (N_6286,N_5203,N_4981);
nor U6287 (N_6287,N_3788,N_4146);
nand U6288 (N_6288,N_3820,N_5302);
nor U6289 (N_6289,N_5964,N_4181);
nand U6290 (N_6290,N_4083,N_5978);
nand U6291 (N_6291,N_3584,N_5602);
or U6292 (N_6292,N_4705,N_5325);
nor U6293 (N_6293,N_5486,N_3954);
and U6294 (N_6294,N_3283,N_4402);
and U6295 (N_6295,N_5390,N_5327);
nand U6296 (N_6296,N_3103,N_3201);
nor U6297 (N_6297,N_3026,N_3555);
nand U6298 (N_6298,N_5961,N_3967);
or U6299 (N_6299,N_3498,N_4137);
and U6300 (N_6300,N_4108,N_4486);
and U6301 (N_6301,N_5738,N_5894);
nor U6302 (N_6302,N_4424,N_3529);
nor U6303 (N_6303,N_5159,N_4795);
nor U6304 (N_6304,N_3381,N_4197);
xnor U6305 (N_6305,N_3276,N_5595);
and U6306 (N_6306,N_3152,N_5592);
nor U6307 (N_6307,N_4367,N_3875);
and U6308 (N_6308,N_4335,N_5912);
nor U6309 (N_6309,N_5614,N_3612);
or U6310 (N_6310,N_3871,N_5673);
nor U6311 (N_6311,N_4120,N_4148);
and U6312 (N_6312,N_4445,N_4925);
or U6313 (N_6313,N_3631,N_4356);
nand U6314 (N_6314,N_3446,N_4858);
and U6315 (N_6315,N_4462,N_5093);
nor U6316 (N_6316,N_5542,N_5221);
nor U6317 (N_6317,N_3842,N_3857);
or U6318 (N_6318,N_3678,N_3241);
nand U6319 (N_6319,N_5248,N_3171);
and U6320 (N_6320,N_3439,N_4429);
or U6321 (N_6321,N_5041,N_5026);
nand U6322 (N_6322,N_3959,N_4142);
and U6323 (N_6323,N_3585,N_3707);
and U6324 (N_6324,N_3408,N_5229);
and U6325 (N_6325,N_3219,N_5766);
nor U6326 (N_6326,N_4565,N_4286);
and U6327 (N_6327,N_4671,N_3254);
nor U6328 (N_6328,N_5703,N_4594);
nor U6329 (N_6329,N_4830,N_4103);
or U6330 (N_6330,N_3587,N_3179);
or U6331 (N_6331,N_3900,N_3415);
or U6332 (N_6332,N_5166,N_3080);
nand U6333 (N_6333,N_4808,N_5130);
or U6334 (N_6334,N_4324,N_4944);
nor U6335 (N_6335,N_4624,N_5308);
nor U6336 (N_6336,N_3943,N_4440);
nor U6337 (N_6337,N_4357,N_3822);
and U6338 (N_6338,N_5919,N_4346);
or U6339 (N_6339,N_4997,N_3784);
nor U6340 (N_6340,N_3213,N_3483);
nand U6341 (N_6341,N_3552,N_5569);
and U6342 (N_6342,N_5989,N_5845);
nand U6343 (N_6343,N_4466,N_5805);
nand U6344 (N_6344,N_4583,N_3573);
xor U6345 (N_6345,N_5675,N_4924);
and U6346 (N_6346,N_3764,N_5242);
or U6347 (N_6347,N_5833,N_5007);
and U6348 (N_6348,N_5927,N_4872);
and U6349 (N_6349,N_3572,N_3168);
and U6350 (N_6350,N_4413,N_4839);
or U6351 (N_6351,N_5815,N_3995);
nand U6352 (N_6352,N_3352,N_5755);
nor U6353 (N_6353,N_3141,N_4793);
and U6354 (N_6354,N_4749,N_3940);
nor U6355 (N_6355,N_4251,N_5158);
and U6356 (N_6356,N_3742,N_5326);
nor U6357 (N_6357,N_4977,N_5915);
and U6358 (N_6358,N_4779,N_4076);
nor U6359 (N_6359,N_5523,N_5318);
and U6360 (N_6360,N_3629,N_5027);
nand U6361 (N_6361,N_4147,N_5949);
or U6362 (N_6362,N_4007,N_5014);
or U6363 (N_6363,N_4536,N_3577);
and U6364 (N_6364,N_3072,N_5005);
nand U6365 (N_6365,N_3843,N_3970);
and U6366 (N_6366,N_3323,N_4165);
or U6367 (N_6367,N_4688,N_3854);
nand U6368 (N_6368,N_3609,N_3207);
and U6369 (N_6369,N_4877,N_4016);
nor U6370 (N_6370,N_4757,N_3076);
nand U6371 (N_6371,N_4701,N_4295);
and U6372 (N_6372,N_5280,N_3889);
nor U6373 (N_6373,N_3926,N_4172);
or U6374 (N_6374,N_4057,N_3858);
nand U6375 (N_6375,N_5565,N_4906);
nand U6376 (N_6376,N_4661,N_4618);
and U6377 (N_6377,N_5067,N_3803);
and U6378 (N_6378,N_5952,N_3063);
or U6379 (N_6379,N_5887,N_5709);
or U6380 (N_6380,N_5593,N_3914);
nor U6381 (N_6381,N_3002,N_4194);
and U6382 (N_6382,N_3867,N_3176);
or U6383 (N_6383,N_4531,N_5899);
and U6384 (N_6384,N_3515,N_4401);
nor U6385 (N_6385,N_4229,N_3376);
nor U6386 (N_6386,N_5149,N_5572);
and U6387 (N_6387,N_5926,N_3445);
nand U6388 (N_6388,N_5954,N_5856);
nand U6389 (N_6389,N_4625,N_4752);
and U6390 (N_6390,N_3461,N_5640);
and U6391 (N_6391,N_5023,N_3502);
nor U6392 (N_6392,N_5540,N_4864);
and U6393 (N_6393,N_3759,N_5501);
nand U6394 (N_6394,N_3801,N_5133);
and U6395 (N_6395,N_5482,N_3664);
nor U6396 (N_6396,N_4696,N_5478);
nand U6397 (N_6397,N_5307,N_3711);
xor U6398 (N_6398,N_5011,N_5534);
or U6399 (N_6399,N_5965,N_5388);
and U6400 (N_6400,N_4848,N_5247);
nor U6401 (N_6401,N_4075,N_3522);
and U6402 (N_6402,N_3365,N_3856);
nor U6403 (N_6403,N_4804,N_5315);
and U6404 (N_6404,N_3544,N_5403);
nand U6405 (N_6405,N_4796,N_3100);
and U6406 (N_6406,N_5271,N_3934);
and U6407 (N_6407,N_4114,N_5428);
and U6408 (N_6408,N_5789,N_3018);
or U6409 (N_6409,N_4233,N_5936);
and U6410 (N_6410,N_4350,N_5153);
and U6411 (N_6411,N_3218,N_4745);
or U6412 (N_6412,N_5596,N_4476);
nor U6413 (N_6413,N_4030,N_5657);
nor U6414 (N_6414,N_4975,N_5028);
xnor U6415 (N_6415,N_4099,N_5903);
or U6416 (N_6416,N_5140,N_4349);
nor U6417 (N_6417,N_3942,N_4659);
nand U6418 (N_6418,N_5890,N_3050);
nor U6419 (N_6419,N_5452,N_3172);
and U6420 (N_6420,N_4959,N_5310);
nor U6421 (N_6421,N_3235,N_3356);
xor U6422 (N_6422,N_3766,N_4776);
or U6423 (N_6423,N_4017,N_5182);
and U6424 (N_6424,N_3641,N_3977);
nand U6425 (N_6425,N_5974,N_4585);
or U6426 (N_6426,N_4822,N_3273);
nand U6427 (N_6427,N_3312,N_3216);
nand U6428 (N_6428,N_4673,N_4859);
or U6429 (N_6429,N_5373,N_3570);
or U6430 (N_6430,N_3199,N_4275);
and U6431 (N_6431,N_5518,N_3700);
or U6432 (N_6432,N_3380,N_5847);
nor U6433 (N_6433,N_4400,N_5652);
nor U6434 (N_6434,N_3421,N_3827);
and U6435 (N_6435,N_3267,N_5102);
nand U6436 (N_6436,N_3378,N_4654);
nor U6437 (N_6437,N_4886,N_4071);
nor U6438 (N_6438,N_5211,N_5457);
nand U6439 (N_6439,N_4901,N_5858);
nand U6440 (N_6440,N_5034,N_4759);
and U6441 (N_6441,N_4963,N_4515);
or U6442 (N_6442,N_3094,N_5380);
and U6443 (N_6443,N_3689,N_4321);
or U6444 (N_6444,N_4791,N_5558);
nor U6445 (N_6445,N_4538,N_3363);
nor U6446 (N_6446,N_4723,N_5483);
nand U6447 (N_6447,N_4005,N_5022);
nor U6448 (N_6448,N_5687,N_5042);
and U6449 (N_6449,N_5767,N_5008);
nand U6450 (N_6450,N_3719,N_4773);
nand U6451 (N_6451,N_3920,N_5761);
nand U6452 (N_6452,N_5139,N_4459);
nand U6453 (N_6453,N_4573,N_5816);
or U6454 (N_6454,N_4314,N_3905);
xor U6455 (N_6455,N_5258,N_3212);
nor U6456 (N_6456,N_5099,N_4789);
nor U6457 (N_6457,N_5150,N_4999);
and U6458 (N_6458,N_3607,N_3327);
nor U6459 (N_6459,N_5291,N_5001);
nor U6460 (N_6460,N_5702,N_3256);
or U6461 (N_6461,N_3047,N_4315);
nor U6462 (N_6462,N_4477,N_4371);
nand U6463 (N_6463,N_3562,N_4134);
or U6464 (N_6464,N_3919,N_5319);
or U6465 (N_6465,N_4570,N_3939);
and U6466 (N_6466,N_5286,N_3825);
and U6467 (N_6467,N_4046,N_5568);
nor U6468 (N_6468,N_5902,N_5108);
nor U6469 (N_6469,N_4894,N_3608);
or U6470 (N_6470,N_4337,N_5716);
nor U6471 (N_6471,N_5790,N_5970);
nor U6472 (N_6472,N_4638,N_3345);
nand U6473 (N_6473,N_4451,N_5293);
or U6474 (N_6474,N_3334,N_4406);
or U6475 (N_6475,N_4110,N_5469);
nor U6476 (N_6476,N_4876,N_5335);
and U6477 (N_6477,N_5183,N_5404);
and U6478 (N_6478,N_5591,N_5456);
and U6479 (N_6479,N_4269,N_4145);
nand U6480 (N_6480,N_4447,N_5825);
nor U6481 (N_6481,N_3937,N_3029);
or U6482 (N_6482,N_4062,N_4582);
and U6483 (N_6483,N_3038,N_4670);
nand U6484 (N_6484,N_5874,N_5461);
and U6485 (N_6485,N_4562,N_5618);
nor U6486 (N_6486,N_5393,N_5737);
and U6487 (N_6487,N_4807,N_3490);
nand U6488 (N_6488,N_5313,N_3847);
and U6489 (N_6489,N_5730,N_3733);
nor U6490 (N_6490,N_4302,N_3024);
nor U6491 (N_6491,N_5844,N_5548);
and U6492 (N_6492,N_5680,N_4529);
or U6493 (N_6493,N_3113,N_4574);
xor U6494 (N_6494,N_4086,N_5777);
or U6495 (N_6495,N_4614,N_3985);
and U6496 (N_6496,N_4130,N_4308);
nor U6497 (N_6497,N_4232,N_3770);
xor U6498 (N_6498,N_5836,N_3837);
and U6499 (N_6499,N_5862,N_3274);
and U6500 (N_6500,N_5803,N_5932);
or U6501 (N_6501,N_4714,N_3073);
nor U6502 (N_6502,N_4060,N_3249);
nand U6503 (N_6503,N_4387,N_4448);
nor U6504 (N_6504,N_3974,N_4978);
or U6505 (N_6505,N_4047,N_4511);
or U6506 (N_6506,N_5634,N_4632);
nand U6507 (N_6507,N_3866,N_5262);
nor U6508 (N_6508,N_5068,N_4265);
nand U6509 (N_6509,N_4433,N_5117);
and U6510 (N_6510,N_5914,N_4837);
and U6511 (N_6511,N_5946,N_3650);
nand U6512 (N_6512,N_3679,N_4496);
nand U6513 (N_6513,N_3245,N_5619);
xor U6514 (N_6514,N_4693,N_5240);
and U6515 (N_6515,N_5732,N_4123);
or U6516 (N_6516,N_5097,N_5064);
nand U6517 (N_6517,N_4668,N_3833);
xnor U6518 (N_6518,N_5924,N_3288);
and U6519 (N_6519,N_3505,N_4548);
nor U6520 (N_6520,N_4199,N_3104);
and U6521 (N_6521,N_3718,N_4514);
nand U6522 (N_6522,N_4812,N_3738);
nand U6523 (N_6523,N_4398,N_3778);
and U6524 (N_6524,N_5261,N_5119);
or U6525 (N_6525,N_4902,N_4935);
and U6526 (N_6526,N_4084,N_4301);
and U6527 (N_6527,N_5098,N_4549);
or U6528 (N_6528,N_4533,N_4694);
or U6529 (N_6529,N_4328,N_5398);
nand U6530 (N_6530,N_5070,N_5047);
nand U6531 (N_6531,N_4608,N_3131);
or U6532 (N_6532,N_3789,N_4809);
or U6533 (N_6533,N_5562,N_3402);
xor U6534 (N_6534,N_5104,N_5784);
or U6535 (N_6535,N_4260,N_4794);
and U6536 (N_6536,N_5905,N_3450);
nor U6537 (N_6537,N_5933,N_5207);
or U6538 (N_6538,N_4726,N_4339);
nand U6539 (N_6539,N_4845,N_3810);
nor U6540 (N_6540,N_5824,N_5991);
or U6541 (N_6541,N_3399,N_3232);
and U6542 (N_6542,N_3392,N_5808);
or U6543 (N_6543,N_4602,N_5298);
nand U6544 (N_6544,N_5187,N_3215);
and U6545 (N_6545,N_3253,N_4572);
nor U6546 (N_6546,N_4031,N_3309);
nand U6547 (N_6547,N_3196,N_3375);
nor U6548 (N_6548,N_4681,N_4506);
nor U6549 (N_6549,N_3351,N_3222);
nor U6550 (N_6550,N_4962,N_4487);
nor U6551 (N_6551,N_3804,N_4792);
or U6552 (N_6552,N_4512,N_4422);
and U6553 (N_6553,N_5746,N_4824);
or U6554 (N_6554,N_5748,N_4954);
nor U6555 (N_6555,N_3632,N_5567);
or U6556 (N_6556,N_4589,N_5669);
and U6557 (N_6557,N_4898,N_4474);
or U6558 (N_6558,N_3567,N_3454);
and U6559 (N_6559,N_5381,N_3795);
nand U6560 (N_6560,N_4653,N_4383);
and U6561 (N_6561,N_4699,N_5220);
and U6562 (N_6562,N_4908,N_3877);
nand U6563 (N_6563,N_4891,N_3062);
xor U6564 (N_6564,N_5420,N_4785);
and U6565 (N_6565,N_5556,N_4481);
nor U6566 (N_6566,N_4929,N_5201);
nand U6567 (N_6567,N_5817,N_5900);
nor U6568 (N_6568,N_5223,N_4816);
nor U6569 (N_6569,N_3853,N_5739);
or U6570 (N_6570,N_4933,N_4666);
nor U6571 (N_6571,N_5179,N_4497);
or U6572 (N_6572,N_3606,N_3434);
nand U6573 (N_6573,N_4866,N_4136);
nor U6574 (N_6574,N_3458,N_3187);
or U6575 (N_6575,N_5164,N_3910);
nand U6576 (N_6576,N_3485,N_3371);
nor U6577 (N_6577,N_5421,N_4527);
and U6578 (N_6578,N_4905,N_5377);
nand U6579 (N_6579,N_4425,N_3756);
nand U6580 (N_6580,N_5445,N_5063);
nor U6581 (N_6581,N_3911,N_5686);
nor U6582 (N_6582,N_4431,N_3895);
nor U6583 (N_6583,N_5697,N_3145);
and U6584 (N_6584,N_5061,N_3355);
nor U6585 (N_6585,N_5101,N_4449);
and U6586 (N_6586,N_5125,N_3150);
and U6587 (N_6587,N_3367,N_4831);
and U6588 (N_6588,N_3775,N_3277);
and U6589 (N_6589,N_5945,N_3090);
nor U6590 (N_6590,N_3056,N_4293);
or U6591 (N_6591,N_3990,N_4827);
and U6592 (N_6592,N_5642,N_4534);
or U6593 (N_6593,N_5405,N_3547);
and U6594 (N_6594,N_5439,N_3662);
nand U6595 (N_6595,N_5109,N_4706);
or U6596 (N_6596,N_4798,N_5553);
or U6597 (N_6597,N_3174,N_4222);
or U6598 (N_6598,N_5893,N_3929);
or U6599 (N_6599,N_5090,N_5292);
nand U6600 (N_6600,N_3538,N_3242);
nor U6601 (N_6601,N_5132,N_3978);
or U6602 (N_6602,N_5051,N_3229);
or U6603 (N_6603,N_5823,N_4094);
nor U6604 (N_6604,N_5055,N_4081);
nand U6605 (N_6605,N_3349,N_5496);
or U6606 (N_6606,N_5509,N_4904);
nand U6607 (N_6607,N_5988,N_5502);
nand U6608 (N_6608,N_5972,N_3404);
nand U6609 (N_6609,N_3435,N_4586);
nor U6610 (N_6610,N_3225,N_4079);
nand U6611 (N_6611,N_5043,N_3124);
nor U6612 (N_6612,N_3624,N_4152);
nor U6613 (N_6613,N_5342,N_5753);
nand U6614 (N_6614,N_4674,N_5386);
nor U6615 (N_6615,N_3726,N_5958);
nand U6616 (N_6616,N_4774,N_4940);
and U6617 (N_6617,N_4095,N_5347);
or U6618 (N_6618,N_3194,N_4174);
and U6619 (N_6619,N_4702,N_3762);
or U6620 (N_6620,N_4765,N_5707);
nor U6621 (N_6621,N_4680,N_4722);
nor U6622 (N_6622,N_4432,N_3000);
or U6623 (N_6623,N_3714,N_4288);
nand U6624 (N_6624,N_3221,N_3611);
nor U6625 (N_6625,N_4348,N_4377);
nand U6626 (N_6626,N_5060,N_5681);
nor U6627 (N_6627,N_3101,N_4832);
or U6628 (N_6628,N_5173,N_5506);
or U6629 (N_6629,N_4252,N_4861);
nand U6630 (N_6630,N_4127,N_3908);
or U6631 (N_6631,N_5020,N_4629);
nor U6632 (N_6632,N_5528,N_4596);
or U6633 (N_6633,N_4786,N_4262);
xor U6634 (N_6634,N_4524,N_5867);
nor U6635 (N_6635,N_3469,N_5979);
or U6636 (N_6636,N_5654,N_3189);
nor U6637 (N_6637,N_4956,N_4679);
and U6638 (N_6638,N_4151,N_3595);
or U6639 (N_6639,N_4883,N_5399);
nor U6640 (N_6640,N_4101,N_5625);
or U6641 (N_6641,N_3696,N_3891);
nand U6642 (N_6642,N_5822,N_5069);
and U6643 (N_6643,N_3517,N_4814);
nand U6644 (N_6644,N_4716,N_3467);
nor U6645 (N_6645,N_5891,N_5612);
or U6646 (N_6646,N_5641,N_5254);
nand U6647 (N_6647,N_4810,N_4479);
or U6648 (N_6648,N_5923,N_5610);
and U6649 (N_6649,N_5414,N_4412);
nand U6650 (N_6650,N_5760,N_4153);
and U6651 (N_6651,N_4728,N_3405);
nand U6652 (N_6652,N_3532,N_4860);
xor U6653 (N_6653,N_4994,N_5278);
nor U6654 (N_6654,N_3055,N_5917);
and U6655 (N_6655,N_3746,N_4185);
nor U6656 (N_6656,N_3049,N_5598);
or U6657 (N_6657,N_5015,N_3874);
nor U6658 (N_6658,N_3702,N_5204);
nand U6659 (N_6659,N_3030,N_4236);
or U6660 (N_6660,N_5199,N_5239);
nand U6661 (N_6661,N_5848,N_5080);
and U6662 (N_6662,N_4919,N_3087);
nor U6663 (N_6663,N_5180,N_4717);
nor U6664 (N_6664,N_4771,N_3093);
nor U6665 (N_6665,N_5688,N_3883);
or U6666 (N_6666,N_4982,N_4747);
or U6667 (N_6667,N_4336,N_5078);
nor U6668 (N_6668,N_5463,N_3343);
nand U6669 (N_6669,N_5287,N_3824);
or U6670 (N_6670,N_5892,N_4525);
nor U6671 (N_6671,N_5604,N_4601);
and U6672 (N_6672,N_5871,N_4427);
nor U6673 (N_6673,N_5356,N_3817);
or U6674 (N_6674,N_4027,N_3773);
xnor U6675 (N_6675,N_3239,N_4719);
and U6676 (N_6676,N_5889,N_5725);
or U6677 (N_6677,N_4106,N_4090);
nor U6678 (N_6678,N_5645,N_3736);
nand U6679 (N_6679,N_3761,N_5851);
xnor U6680 (N_6680,N_4188,N_4215);
or U6681 (N_6681,N_5383,N_5536);
and U6682 (N_6682,N_4974,N_4453);
nand U6683 (N_6683,N_5082,N_3307);
nand U6684 (N_6684,N_5769,N_4516);
nand U6685 (N_6685,N_4319,N_4996);
or U6686 (N_6686,N_3329,N_3296);
and U6687 (N_6687,N_4182,N_3396);
nand U6688 (N_6688,N_5877,N_3084);
nand U6689 (N_6689,N_3470,N_3270);
nand U6690 (N_6690,N_5505,N_4358);
and U6691 (N_6691,N_4287,N_4584);
nor U6692 (N_6692,N_4426,N_4312);
or U6693 (N_6693,N_4734,N_4968);
and U6694 (N_6694,N_5301,N_5105);
nor U6695 (N_6695,N_5551,N_5849);
and U6696 (N_6696,N_5413,N_5854);
and U6697 (N_6697,N_5859,N_5646);
nand U6698 (N_6698,N_3694,N_3302);
nor U6699 (N_6699,N_4677,N_4239);
or U6700 (N_6700,N_5050,N_4912);
nand U6701 (N_6701,N_3823,N_4537);
and U6702 (N_6702,N_3708,N_3036);
nor U6703 (N_6703,N_5519,N_5025);
nand U6704 (N_6704,N_4168,N_3504);
nand U6705 (N_6705,N_4778,N_3428);
and U6706 (N_6706,N_3337,N_4892);
or U6707 (N_6707,N_3155,N_5729);
nand U6708 (N_6708,N_3811,N_5216);
nand U6709 (N_6709,N_4294,N_3298);
or U6710 (N_6710,N_3706,N_4494);
or U6711 (N_6711,N_3228,N_4813);
nor U6712 (N_6712,N_4619,N_3957);
or U6713 (N_6713,N_5986,N_5717);
nand U6714 (N_6714,N_5479,N_4190);
and U6715 (N_6715,N_3372,N_3701);
nor U6716 (N_6716,N_3899,N_3754);
nand U6717 (N_6717,N_3042,N_5812);
nand U6718 (N_6718,N_4609,N_4292);
or U6719 (N_6719,N_5751,N_4687);
and U6720 (N_6720,N_4029,N_3870);
and U6721 (N_6721,N_5081,N_4244);
nand U6722 (N_6722,N_4662,N_3593);
or U6723 (N_6723,N_4874,N_3933);
or U6724 (N_6724,N_4183,N_5237);
nor U6725 (N_6725,N_5444,N_3496);
or U6726 (N_6726,N_4310,N_3639);
nand U6727 (N_6727,N_5106,N_3414);
nor U6728 (N_6728,N_4196,N_4551);
nor U6729 (N_6729,N_3868,N_4817);
and U6730 (N_6730,N_5276,N_5906);
or U6731 (N_6731,N_5712,N_5685);
nor U6732 (N_6732,N_5138,N_3206);
xor U6733 (N_6733,N_3941,N_3841);
and U6734 (N_6734,N_5417,N_5533);
and U6735 (N_6735,N_4909,N_4686);
nand U6736 (N_6736,N_3873,N_3308);
nand U6737 (N_6737,N_3068,N_5692);
or U6738 (N_6738,N_5490,N_5181);
and U6739 (N_6739,N_3361,N_4274);
nor U6740 (N_6740,N_4220,N_5791);
and U6741 (N_6741,N_5257,N_3161);
and U6742 (N_6742,N_5606,N_4838);
and U6743 (N_6743,N_4002,N_4354);
nand U6744 (N_6744,N_5843,N_4564);
and U6745 (N_6745,N_4317,N_5378);
or U6746 (N_6746,N_5305,N_4157);
or U6747 (N_6747,N_3772,N_3962);
and U6748 (N_6748,N_3133,N_5363);
nor U6749 (N_6749,N_5886,N_4710);
nand U6750 (N_6750,N_5710,N_3191);
or U6751 (N_6751,N_4087,N_5666);
and U6752 (N_6752,N_5151,N_5163);
nor U6753 (N_6753,N_4439,N_5814);
nor U6754 (N_6754,N_5617,N_4787);
and U6755 (N_6755,N_4560,N_3879);
nor U6756 (N_6756,N_5424,N_5243);
and U6757 (N_6757,N_4542,N_5205);
nor U6758 (N_6758,N_5492,N_5009);
or U6759 (N_6759,N_4663,N_3054);
and U6760 (N_6760,N_4051,N_5541);
or U6761 (N_6761,N_3703,N_3117);
xnor U6762 (N_6762,N_4689,N_5045);
nor U6763 (N_6763,N_4365,N_5749);
or U6764 (N_6764,N_4058,N_3438);
or U6765 (N_6765,N_5169,N_4885);
nand U6766 (N_6766,N_3389,N_3447);
nor U6767 (N_6767,N_4299,N_5547);
nand U6768 (N_6768,N_5029,N_5581);
nand U6769 (N_6769,N_5495,N_4113);
and U6770 (N_6770,N_3682,N_4703);
nor U6771 (N_6771,N_4160,N_5529);
nor U6772 (N_6772,N_3457,N_5395);
xnor U6773 (N_6773,N_3119,N_5425);
nor U6774 (N_6774,N_3388,N_5030);
nand U6775 (N_6775,N_3845,N_3134);
or U6776 (N_6776,N_3695,N_3115);
and U6777 (N_6777,N_3240,N_4911);
and U6778 (N_6778,N_4122,N_5084);
xnor U6779 (N_6779,N_5391,N_4563);
nand U6780 (N_6780,N_3052,N_4547);
and U6781 (N_6781,N_5462,N_3566);
or U6782 (N_6782,N_3559,N_3661);
nand U6783 (N_6783,N_4568,N_5230);
nor U6784 (N_6784,N_3723,N_4501);
and U6785 (N_6785,N_4036,N_5111);
nand U6786 (N_6786,N_5901,N_4522);
nand U6787 (N_6787,N_3834,N_3493);
nand U6788 (N_6788,N_3715,N_3921);
or U6789 (N_6789,N_4767,N_4467);
nor U6790 (N_6790,N_4208,N_5499);
and U6791 (N_6791,N_4676,N_5997);
or U6792 (N_6792,N_4450,N_5129);
xor U6793 (N_6793,N_4721,N_3089);
and U6794 (N_6794,N_3790,N_5522);
xor U6795 (N_6795,N_4928,N_5477);
or U6796 (N_6796,N_3448,N_3503);
and U6797 (N_6797,N_3184,N_3997);
or U6798 (N_6798,N_5213,N_4227);
nand U6799 (N_6799,N_4006,N_3802);
or U6800 (N_6800,N_3384,N_3537);
and U6801 (N_6801,N_5460,N_5736);
and U6802 (N_6802,N_4715,N_3136);
and U6803 (N_6803,N_4297,N_3335);
and U6804 (N_6804,N_3655,N_4732);
nand U6805 (N_6805,N_5465,N_3521);
nor U6806 (N_6806,N_3007,N_5162);
nand U6807 (N_6807,N_5544,N_5842);
nor U6808 (N_6808,N_4015,N_4748);
nor U6809 (N_6809,N_5017,N_4634);
nand U6810 (N_6810,N_3224,N_4772);
nand U6811 (N_6811,N_4851,N_3864);
and U6812 (N_6812,N_4805,N_3705);
and U6813 (N_6813,N_4304,N_3744);
or U6814 (N_6814,N_3961,N_3127);
nor U6815 (N_6815,N_4580,N_5217);
nand U6816 (N_6816,N_5870,N_5740);
nand U6817 (N_6817,N_3647,N_5883);
or U6818 (N_6818,N_4664,N_3601);
or U6819 (N_6819,N_3317,N_3513);
nand U6820 (N_6820,N_3580,N_5345);
nor U6821 (N_6821,N_3814,N_4393);
nor U6822 (N_6822,N_4844,N_4434);
nand U6823 (N_6823,N_4231,N_5637);
nand U6824 (N_6824,N_3430,N_5372);
and U6825 (N_6825,N_4177,N_4893);
nor U6826 (N_6826,N_5035,N_4309);
nor U6827 (N_6827,N_5752,N_4841);
and U6828 (N_6828,N_5157,N_3003);
nor U6829 (N_6829,N_5306,N_3887);
nand U6830 (N_6830,N_5696,N_4672);
xnor U6831 (N_6831,N_5146,N_5689);
nor U6832 (N_6832,N_3099,N_3401);
nand U6833 (N_6833,N_3464,N_5114);
nand U6834 (N_6834,N_4163,N_3478);
and U6835 (N_6835,N_4976,N_3771);
or U6836 (N_6836,N_4639,N_3132);
nand U6837 (N_6837,N_3182,N_3821);
nor U6838 (N_6838,N_3146,N_4628);
or U6839 (N_6839,N_3109,N_3516);
and U6840 (N_6840,N_3320,N_4979);
nor U6841 (N_6841,N_3223,N_3074);
nor U6842 (N_6842,N_5663,N_4821);
nor U6843 (N_6843,N_5031,N_3306);
nor U6844 (N_6844,N_5826,N_3960);
nor U6845 (N_6845,N_3156,N_3468);
nor U6846 (N_6846,N_4407,N_3511);
nand U6847 (N_6847,N_5480,N_5517);
nor U6848 (N_6848,N_5913,N_4880);
nand U6849 (N_6849,N_5037,N_4937);
nor U6850 (N_6850,N_3869,N_3777);
nand U6851 (N_6851,N_5999,N_5411);
or U6852 (N_6852,N_4995,N_3753);
or U6853 (N_6853,N_4254,N_4363);
nand U6854 (N_6854,N_4990,N_5350);
or U6855 (N_6855,N_4133,N_3994);
nor U6856 (N_6856,N_5700,N_4285);
and U6857 (N_6857,N_3812,N_3627);
and U6858 (N_6858,N_5577,N_3721);
or U6859 (N_6859,N_3983,N_5683);
and U6860 (N_6860,N_4667,N_5284);
nor U6861 (N_6861,N_4556,N_5010);
and U6862 (N_6862,N_5597,N_3284);
nand U6863 (N_6863,N_5792,N_3387);
and U6864 (N_6864,N_5574,N_3913);
and U6865 (N_6865,N_4096,N_5537);
nor U6866 (N_6866,N_3808,N_4558);
or U6867 (N_6867,N_3667,N_5880);
and U6868 (N_6868,N_4303,N_4155);
or U6869 (N_6869,N_3106,N_4173);
xor U6870 (N_6870,N_5255,N_3043);
nor U6871 (N_6871,N_5672,N_4720);
or U6872 (N_6872,N_5699,N_3303);
nand U6873 (N_6873,N_4819,N_3669);
and U6874 (N_6874,N_3799,N_4242);
and U6875 (N_6875,N_3748,N_3558);
nand U6876 (N_6876,N_5468,N_3107);
or U6877 (N_6877,N_5277,N_3097);
and U6878 (N_6878,N_4225,N_4865);
nand U6879 (N_6879,N_3623,N_5788);
or U6880 (N_6880,N_5379,N_3366);
and U6881 (N_6881,N_3021,N_5876);
or U6882 (N_6882,N_3070,N_4887);
nor U6883 (N_6883,N_5578,N_4186);
or U6884 (N_6884,N_5134,N_3463);
and U6885 (N_6885,N_3319,N_4603);
or U6886 (N_6886,N_4842,N_5368);
nor U6887 (N_6887,N_4769,N_4078);
and U6888 (N_6888,N_5953,N_3749);
or U6889 (N_6889,N_5690,N_3745);
and U6890 (N_6890,N_4647,N_5218);
and U6891 (N_6891,N_3932,N_5628);
nor U6892 (N_6892,N_3979,N_5801);
nand U6893 (N_6893,N_5512,N_3965);
or U6894 (N_6894,N_5155,N_5840);
and U6895 (N_6895,N_5644,N_3071);
and U6896 (N_6896,N_3144,N_3948);
and U6897 (N_6897,N_5273,N_4727);
xor U6898 (N_6898,N_3594,N_4491);
nor U6899 (N_6899,N_3484,N_3077);
nand U6900 (N_6900,N_3735,N_5714);
and U6901 (N_6901,N_3347,N_3118);
nor U6902 (N_6902,N_5813,N_3579);
nor U6903 (N_6903,N_4665,N_3666);
nor U6904 (N_6904,N_3691,N_4504);
nand U6905 (N_6905,N_4972,N_5360);
xor U6906 (N_6906,N_3725,N_5195);
or U6907 (N_6907,N_5176,N_5762);
or U6908 (N_6908,N_5124,N_4559);
or U6909 (N_6909,N_4801,N_5566);
or U6910 (N_6910,N_5348,N_5554);
or U6911 (N_6911,N_3643,N_4761);
and U6912 (N_6912,N_3992,N_4868);
nand U6913 (N_6913,N_5358,N_3266);
or U6914 (N_6914,N_4918,N_3791);
nor U6915 (N_6915,N_5334,N_5226);
and U6916 (N_6916,N_3163,N_3765);
nand U6917 (N_6917,N_3966,N_3712);
nand U6918 (N_6918,N_5706,N_3096);
nor U6919 (N_6919,N_4158,N_4650);
xor U6920 (N_6920,N_5336,N_4169);
or U6921 (N_6921,N_4637,N_3362);
and U6922 (N_6922,N_5909,N_4544);
xnor U6923 (N_6923,N_5331,N_3963);
nor U6924 (N_6924,N_3596,N_3687);
nor U6925 (N_6925,N_5400,N_5535);
or U6926 (N_6926,N_4126,N_5364);
nand U6927 (N_6927,N_3188,N_5283);
nand U6928 (N_6928,N_4764,N_3648);
nand U6929 (N_6929,N_3451,N_4684);
nand U6930 (N_6930,N_4217,N_4566);
and U6931 (N_6931,N_5580,N_3017);
or U6932 (N_6932,N_4226,N_3514);
xor U6933 (N_6933,N_4203,N_5866);
nand U6934 (N_6934,N_3015,N_3110);
or U6935 (N_6935,N_5994,N_3583);
nand U6936 (N_6936,N_5122,N_3620);
and U6937 (N_6937,N_3394,N_4198);
or U6938 (N_6938,N_4658,N_5525);
and U6939 (N_6939,N_5875,N_5323);
nor U6940 (N_6940,N_5971,N_5670);
nor U6941 (N_6941,N_5160,N_3805);
or U6942 (N_6942,N_4264,N_3878);
nor U6943 (N_6943,N_4072,N_4927);
nand U6944 (N_6944,N_3618,N_4176);
nor U6945 (N_6945,N_5731,N_3091);
or U6946 (N_6946,N_3531,N_5219);
xor U6947 (N_6947,N_4951,N_4485);
nor U6948 (N_6948,N_3763,N_5200);
or U6949 (N_6949,N_5021,N_3506);
or U6950 (N_6950,N_3747,N_5561);
or U6951 (N_6951,N_4991,N_3980);
xor U6952 (N_6952,N_5092,N_3673);
and U6953 (N_6953,N_5423,N_3474);
or U6954 (N_6954,N_5793,N_4942);
nand U6955 (N_6955,N_4054,N_3259);
and U6956 (N_6956,N_5629,N_3373);
or U6957 (N_6957,N_3481,N_4088);
nand U6958 (N_6958,N_3512,N_3227);
and U6959 (N_6959,N_5320,N_3325);
nor U6960 (N_6960,N_5782,N_5768);
or U6961 (N_6961,N_3644,N_3210);
or U6962 (N_6962,N_3637,N_5198);
or U6963 (N_6963,N_5096,N_4342);
nand U6964 (N_6964,N_5189,N_3315);
and U6965 (N_6965,N_3523,N_4595);
nand U6966 (N_6966,N_3449,N_4224);
or U6967 (N_6967,N_4704,N_3477);
and U6968 (N_6968,N_4781,N_5086);
or U6969 (N_6969,N_3403,N_4192);
nand U6970 (N_6970,N_3078,N_4035);
and U6971 (N_6971,N_5359,N_3553);
or U6972 (N_6972,N_4171,N_3798);
and U6973 (N_6973,N_4397,N_4852);
and U6974 (N_6974,N_3238,N_4191);
nor U6975 (N_6975,N_4281,N_3704);
nor U6976 (N_6976,N_3204,N_3285);
nand U6977 (N_6977,N_5316,N_5431);
nor U6978 (N_6978,N_4139,N_4228);
nand U6979 (N_6979,N_4780,N_5550);
or U6980 (N_6980,N_3368,N_3014);
and U6981 (N_6981,N_5615,N_4682);
or U6982 (N_6982,N_4320,N_5763);
and U6983 (N_6983,N_3479,N_5608);
or U6984 (N_6984,N_3027,N_3657);
nor U6985 (N_6985,N_3818,N_5048);
nand U6986 (N_6986,N_3610,N_4755);
and U6987 (N_6987,N_3065,N_5881);
and U6988 (N_6988,N_5733,N_4124);
nand U6989 (N_6989,N_5743,N_3475);
nand U6990 (N_6990,N_3417,N_3128);
and U6991 (N_6991,N_4381,N_4833);
nand U6992 (N_6992,N_4355,N_3987);
nand U6993 (N_6993,N_3880,N_3286);
or U6994 (N_6994,N_5337,N_4724);
or U6995 (N_6995,N_3079,N_3724);
nor U6996 (N_6996,N_4971,N_5635);
and U6997 (N_6997,N_5908,N_4128);
nor U6998 (N_6998,N_4064,N_5611);
and U6999 (N_6999,N_5190,N_4713);
and U7000 (N_7000,N_3890,N_5245);
or U7001 (N_7001,N_5052,N_5820);
or U7002 (N_7002,N_4042,N_5476);
nor U7003 (N_7003,N_5148,N_4141);
nand U7004 (N_7004,N_5387,N_3045);
nor U7005 (N_7005,N_4736,N_4953);
and U7006 (N_7006,N_5126,N_4890);
or U7007 (N_7007,N_5966,N_3727);
nand U7008 (N_7008,N_3969,N_3716);
nor U7009 (N_7009,N_5263,N_5208);
nand U7010 (N_7010,N_5392,N_5234);
nor U7011 (N_7011,N_3268,N_5759);
and U7012 (N_7012,N_5508,N_5968);
xnor U7013 (N_7013,N_4243,N_5314);
or U7014 (N_7014,N_4826,N_3257);
xnor U7015 (N_7015,N_5266,N_5765);
or U7016 (N_7016,N_3316,N_4253);
nor U7017 (N_7017,N_5192,N_5656);
nand U7018 (N_7018,N_5552,N_5852);
or U7019 (N_7019,N_3530,N_4867);
nor U7020 (N_7020,N_4283,N_5623);
nor U7021 (N_7021,N_5016,N_4802);
nor U7022 (N_7022,N_4489,N_5942);
or U7023 (N_7023,N_4316,N_4987);
nand U7024 (N_7024,N_4870,N_5956);
or U7025 (N_7025,N_3922,N_4008);
or U7026 (N_7026,N_4205,N_5794);
nor U7027 (N_7027,N_4498,N_3357);
nand U7028 (N_7028,N_4430,N_3528);
nor U7029 (N_7029,N_5869,N_4018);
or U7030 (N_7030,N_3064,N_5312);
nor U7031 (N_7031,N_4115,N_3617);
nor U7032 (N_7032,N_4465,N_5583);
or U7033 (N_7033,N_5123,N_5441);
and U7034 (N_7034,N_4175,N_4089);
nand U7035 (N_7035,N_3507,N_5000);
and U7036 (N_7036,N_4600,N_3663);
nor U7037 (N_7037,N_5679,N_5193);
or U7038 (N_7038,N_3993,N_4235);
and U7039 (N_7039,N_3931,N_4675);
or U7040 (N_7040,N_4473,N_4695);
nand U7041 (N_7041,N_3722,N_3459);
or U7042 (N_7042,N_3035,N_3260);
nor U7043 (N_7043,N_3774,N_5491);
and U7044 (N_7044,N_4557,N_4210);
or U7045 (N_7045,N_5724,N_4623);
nand U7046 (N_7046,N_4296,N_3048);
and U7047 (N_7047,N_5603,N_4743);
or U7048 (N_7048,N_3950,N_5426);
or U7049 (N_7049,N_4756,N_4834);
nand U7050 (N_7050,N_5757,N_4121);
and U7051 (N_7051,N_5977,N_4952);
nor U7052 (N_7052,N_5212,N_3230);
and U7053 (N_7053,N_3195,N_4211);
nand U7054 (N_7054,N_3139,N_4352);
nand U7055 (N_7055,N_4263,N_5317);
or U7056 (N_7056,N_5233,N_5671);
or U7057 (N_7057,N_5747,N_4368);
nor U7058 (N_7058,N_4612,N_4657);
nand U7059 (N_7059,N_5018,N_4960);
or U7060 (N_7060,N_3614,N_4611);
or U7061 (N_7061,N_4766,N_3692);
or U7062 (N_7062,N_3111,N_4836);
or U7063 (N_7063,N_4581,N_5418);
nand U7064 (N_7064,N_4758,N_5783);
and U7065 (N_7065,N_3391,N_4931);
nor U7066 (N_7066,N_4162,N_4074);
and U7067 (N_7067,N_5653,N_4050);
nand U7068 (N_7068,N_5361,N_4640);
nand U7069 (N_7069,N_3590,N_5721);
nor U7070 (N_7070,N_5466,N_3338);
nor U7071 (N_7071,N_3998,N_3968);
nand U7072 (N_7072,N_3234,N_4471);
nor U7073 (N_7073,N_5835,N_4032);
and U7074 (N_7074,N_5549,N_5590);
nand U7075 (N_7075,N_4958,N_5779);
nor U7076 (N_7076,N_4170,N_4414);
nor U7077 (N_7077,N_3830,N_4132);
nor U7078 (N_7078,N_5253,N_4107);
or U7079 (N_7079,N_3173,N_4326);
or U7080 (N_7080,N_3755,N_4806);
nand U7081 (N_7081,N_3828,N_5238);
and U7082 (N_7082,N_3554,N_4394);
nand U7083 (N_7083,N_4370,N_4135);
or U7084 (N_7084,N_5643,N_5429);
or U7085 (N_7085,N_5447,N_5057);
or U7086 (N_7086,N_3787,N_4846);
or U7087 (N_7087,N_4313,N_5321);
nor U7088 (N_7088,N_3292,N_4873);
and U7089 (N_7089,N_4004,N_4503);
nand U7090 (N_7090,N_4052,N_3658);
or U7091 (N_7091,N_4421,N_4669);
and U7092 (N_7092,N_5655,N_5521);
or U7093 (N_7093,N_4617,N_4437);
nand U7094 (N_7094,N_4478,N_3936);
nor U7095 (N_7095,N_3564,N_5232);
nand U7096 (N_7096,N_4164,N_3295);
nand U7097 (N_7097,N_5493,N_3876);
nor U7098 (N_7098,N_4266,N_4323);
xor U7099 (N_7099,N_3322,N_3114);
nor U7100 (N_7100,N_3001,N_3151);
and U7101 (N_7101,N_4116,N_5475);
or U7102 (N_7102,N_4998,N_5059);
nor U7103 (N_7103,N_4343,N_3180);
xnor U7104 (N_7104,N_3269,N_3543);
and U7105 (N_7105,N_3536,N_5705);
nor U7106 (N_7106,N_4104,N_5711);
and U7107 (N_7107,N_3717,N_5774);
nand U7108 (N_7108,N_4097,N_5467);
nor U7109 (N_7109,N_5131,N_5165);
nand U7110 (N_7110,N_4329,N_3851);
or U7111 (N_7111,N_3500,N_5033);
and U7112 (N_7112,N_5575,N_3642);
nor U7113 (N_7113,N_4150,N_4380);
xnor U7114 (N_7114,N_3807,N_4443);
or U7115 (N_7115,N_4300,N_4472);
nor U7116 (N_7116,N_3540,N_5620);
and U7117 (N_7117,N_5539,N_4118);
nand U7118 (N_7118,N_3588,N_5973);
nand U7119 (N_7119,N_5633,N_4799);
and U7120 (N_7120,N_4941,N_3621);
or U7121 (N_7121,N_4698,N_3476);
or U7122 (N_7122,N_3592,N_5144);
or U7123 (N_7123,N_3178,N_4875);
xnor U7124 (N_7124,N_3233,N_4068);
and U7125 (N_7125,N_3986,N_5235);
and U7126 (N_7126,N_3699,N_5770);
and U7127 (N_7127,N_4850,N_4784);
nand U7128 (N_7128,N_4518,N_3411);
nor U7129 (N_7129,N_3636,N_4340);
or U7130 (N_7130,N_5831,N_3393);
or U7131 (N_7131,N_4409,N_5975);
or U7132 (N_7132,N_5897,N_4001);
or U7133 (N_7133,N_5650,N_3918);
and U7134 (N_7134,N_5691,N_3205);
nor U7135 (N_7135,N_4555,N_5563);
or U7136 (N_7136,N_5103,N_4207);
nor U7137 (N_7137,N_5898,N_5228);
and U7138 (N_7138,N_3314,N_5601);
or U7139 (N_7139,N_4338,N_5865);
or U7140 (N_7140,N_4373,N_4056);
nor U7141 (N_7141,N_5396,N_4738);
and U7142 (N_7142,N_3729,N_3901);
or U7143 (N_7143,N_4964,N_4144);
or U7144 (N_7144,N_4552,N_4741);
nand U7145 (N_7145,N_5664,N_4372);
or U7146 (N_7146,N_5698,N_4605);
and U7147 (N_7147,N_4125,N_4730);
nand U7148 (N_7148,N_5882,N_4620);
or U7149 (N_7149,N_3947,N_4913);
or U7150 (N_7150,N_3383,N_3646);
nor U7151 (N_7151,N_3258,N_4206);
or U7152 (N_7152,N_3783,N_3760);
nand U7153 (N_7153,N_4038,N_5804);
and U7154 (N_7154,N_3792,N_3731);
nor U7155 (N_7155,N_3265,N_3892);
nand U7156 (N_7156,N_3289,N_3443);
xor U7157 (N_7157,N_3785,N_5415);
nor U7158 (N_7158,N_3040,N_4707);
or U7159 (N_7159,N_4633,N_5076);
or U7160 (N_7160,N_3275,N_3863);
nand U7161 (N_7161,N_3976,N_5780);
or U7162 (N_7162,N_3116,N_5775);
and U7163 (N_7163,N_3649,N_4571);
or U7164 (N_7164,N_5630,N_5773);
nor U7165 (N_7165,N_3186,N_3927);
nand U7166 (N_7166,N_3602,N_5259);
nand U7167 (N_7167,N_3181,N_3425);
nor U7168 (N_7168,N_3852,N_4392);
or U7169 (N_7169,N_3768,N_4973);
or U7170 (N_7170,N_5154,N_3336);
or U7171 (N_7171,N_4843,N_4100);
or U7172 (N_7172,N_4645,N_3209);
nor U7173 (N_7173,N_5513,N_4492);
or U7174 (N_7174,N_3164,N_3915);
and U7175 (N_7175,N_4708,N_4878);
nand U7176 (N_7176,N_5141,N_3020);
nand U7177 (N_7177,N_5419,N_3175);
and U7178 (N_7178,N_3619,N_4416);
nand U7179 (N_7179,N_4250,N_5960);
nor U7180 (N_7180,N_5557,N_3539);
nand U7181 (N_7181,N_4513,N_4709);
or U7182 (N_7182,N_4539,N_3437);
or U7183 (N_7183,N_4914,N_4622);
nand U7184 (N_7184,N_5311,N_5969);
nand U7185 (N_7185,N_5136,N_4856);
nor U7186 (N_7186,N_4305,N_4731);
and U7187 (N_7187,N_4613,N_4055);
nand U7188 (N_7188,N_4577,N_4517);
or U7189 (N_7189,N_3324,N_3058);
nand U7190 (N_7190,N_4578,N_4268);
or U7191 (N_7191,N_5959,N_5860);
nand U7192 (N_7192,N_5800,N_5274);
nor U7193 (N_7193,N_4649,N_4418);
and U7194 (N_7194,N_4502,N_4248);
or U7195 (N_7195,N_3364,N_4484);
or U7196 (N_7196,N_5294,N_4750);
and U7197 (N_7197,N_3796,N_4818);
nand U7198 (N_7198,N_3906,N_5002);
xnor U7199 (N_7199,N_5722,N_5734);
xor U7200 (N_7200,N_3248,N_5171);
nand U7201 (N_7201,N_3924,N_5545);
or U7202 (N_7202,N_5962,N_3013);
and U7203 (N_7203,N_3982,N_4347);
nor U7204 (N_7204,N_4630,N_3640);
nand U7205 (N_7205,N_3409,N_4193);
and U7206 (N_7206,N_5735,N_3190);
nand U7207 (N_7207,N_4457,N_3167);
or U7208 (N_7208,N_4396,N_4746);
nor U7209 (N_7209,N_4325,N_3037);
nor U7210 (N_7210,N_3473,N_3720);
and U7211 (N_7211,N_5091,N_3041);
or U7212 (N_7212,N_3429,N_3200);
nor U7213 (N_7213,N_5367,N_3556);
nand U7214 (N_7214,N_4423,N_5343);
or U7215 (N_7215,N_3121,N_3272);
or U7216 (N_7216,N_5270,N_3019);
nor U7217 (N_7217,N_3293,N_3671);
xor U7218 (N_7218,N_5066,N_3082);
or U7219 (N_7219,N_3192,N_3551);
nor U7220 (N_7220,N_3693,N_5745);
nor U7221 (N_7221,N_4907,N_4828);
nand U7222 (N_7222,N_5963,N_4034);
nor U7223 (N_7223,N_4241,N_3280);
nor U7224 (N_7224,N_4184,N_3398);
nand U7225 (N_7225,N_3126,N_3341);
and U7226 (N_7226,N_3615,N_4249);
nor U7227 (N_7227,N_3769,N_4655);
nor U7228 (N_7228,N_5718,N_3909);
nor U7229 (N_7229,N_5279,N_5374);
and U7230 (N_7230,N_3654,N_5668);
nor U7231 (N_7231,N_4438,N_4800);
or U7232 (N_7232,N_3988,N_3651);
and U7233 (N_7233,N_3888,N_4344);
nand U7234 (N_7234,N_3046,N_3342);
and U7235 (N_7235,N_4692,N_3413);
nand U7236 (N_7236,N_3157,N_4520);
and U7237 (N_7237,N_4469,N_3676);
nor U7238 (N_7238,N_4261,N_4829);
and U7239 (N_7239,N_5450,N_5576);
nor U7240 (N_7240,N_4992,N_3059);
nor U7241 (N_7241,N_3550,N_4825);
nor U7242 (N_7242,N_5435,N_5935);
nor U7243 (N_7243,N_3917,N_3605);
xnor U7244 (N_7244,N_3426,N_5786);
nand U7245 (N_7245,N_5295,N_5351);
nor U7246 (N_7246,N_4013,N_5484);
nor U7247 (N_7247,N_3301,N_5837);
nor U7248 (N_7248,N_3299,N_3143);
nor U7249 (N_7249,N_3734,N_3938);
and U7250 (N_7250,N_4782,N_4610);
or U7251 (N_7251,N_3022,N_5660);
nor U7252 (N_7252,N_3509,N_4733);
and U7253 (N_7253,N_5863,N_5616);
or U7254 (N_7254,N_4768,N_3958);
or U7255 (N_7255,N_4395,N_5487);
xor U7256 (N_7256,N_3793,N_3510);
and U7257 (N_7257,N_3008,N_3850);
or U7258 (N_7258,N_4762,N_3427);
or U7259 (N_7259,N_3840,N_5062);
nor U7260 (N_7260,N_3683,N_5741);
or U7261 (N_7261,N_3060,N_3140);
nor U7262 (N_7262,N_3767,N_5448);
and U7263 (N_7263,N_3816,N_5918);
or U7264 (N_7264,N_3247,N_5407);
nand U7265 (N_7265,N_4507,N_5885);
or U7266 (N_7266,N_3797,N_3250);
and U7267 (N_7267,N_3638,N_5309);
or U7268 (N_7268,N_3972,N_4436);
or U7269 (N_7269,N_5397,N_5720);
and U7270 (N_7270,N_4280,N_3737);
nand U7271 (N_7271,N_5828,N_4033);
nor U7272 (N_7272,N_4712,N_5758);
or U7273 (N_7273,N_3125,N_4934);
nor U7274 (N_7274,N_4279,N_4903);
nor U7275 (N_7275,N_3730,N_4488);
or U7276 (N_7276,N_5947,N_3279);
nand U7277 (N_7277,N_4388,N_5072);
or U7278 (N_7278,N_5177,N_3255);
nor U7279 (N_7279,N_3095,N_5006);
or U7280 (N_7280,N_5987,N_5168);
nand U7281 (N_7281,N_4189,N_3012);
xor U7282 (N_7282,N_5394,N_4985);
nand U7283 (N_7283,N_3006,N_5639);
nor U7284 (N_7284,N_3546,N_3508);
xnor U7285 (N_7285,N_4378,N_5983);
or U7286 (N_7286,N_3713,N_3358);
nand U7287 (N_7287,N_5586,N_5674);
or U7288 (N_7288,N_4777,N_5701);
nand U7289 (N_7289,N_5188,N_3973);
or U7290 (N_7290,N_4039,N_4881);
and U7291 (N_7291,N_5719,N_4073);
and U7292 (N_7292,N_5003,N_5145);
xnor U7293 (N_7293,N_4957,N_4307);
nand U7294 (N_7294,N_3305,N_5990);
or U7295 (N_7295,N_4849,N_4361);
or U7296 (N_7296,N_4070,N_3264);
nand U7297 (N_7297,N_5112,N_4069);
and U7298 (N_7298,N_3603,N_4435);
nor U7299 (N_7299,N_5127,N_5049);
and U7300 (N_7300,N_3928,N_3313);
nand U7301 (N_7301,N_5855,N_3670);
nor U7302 (N_7302,N_4744,N_4111);
or U7303 (N_7303,N_5437,N_3010);
and U7304 (N_7304,N_5324,N_3497);
or U7305 (N_7305,N_4258,N_5085);
and U7306 (N_7306,N_5647,N_4938);
nand U7307 (N_7307,N_4156,N_5985);
and U7308 (N_7308,N_3652,N_5227);
or U7309 (N_7309,N_4362,N_5976);
nand U7310 (N_7310,N_3271,N_3860);
nand U7311 (N_7311,N_3282,N_4621);
or U7312 (N_7312,N_4463,N_3563);
xnor U7313 (N_7313,N_5530,N_5471);
or U7314 (N_7314,N_4811,N_4691);
nor U7315 (N_7315,N_5744,N_5928);
and U7316 (N_7316,N_5888,N_5281);
and U7317 (N_7317,N_5993,N_3211);
or U7318 (N_7318,N_3925,N_5438);
nand U7319 (N_7319,N_4375,N_5446);
nand U7320 (N_7320,N_4290,N_4408);
nor U7321 (N_7321,N_4636,N_4917);
and U7322 (N_7322,N_5362,N_4085);
nor U7323 (N_7323,N_3526,N_5053);
nand U7324 (N_7324,N_4690,N_4410);
nand U7325 (N_7325,N_3633,N_4067);
nor U7326 (N_7326,N_5560,N_4646);
nand U7327 (N_7327,N_5930,N_5304);
xnor U7328 (N_7328,N_4237,N_4797);
nor U7329 (N_7329,N_3882,N_4282);
or U7330 (N_7330,N_5967,N_3075);
and U7331 (N_7331,N_5202,N_4021);
and U7332 (N_7332,N_3148,N_4500);
nand U7333 (N_7333,N_4855,N_3453);
nor U7334 (N_7334,N_5330,N_3294);
or U7335 (N_7335,N_5632,N_5532);
nor U7336 (N_7336,N_5246,N_4490);
nor U7337 (N_7337,N_3656,N_4332);
and U7338 (N_7338,N_5600,N_5458);
xor U7339 (N_7339,N_5594,N_3597);
nand U7340 (N_7340,N_4214,N_5073);
nor U7341 (N_7341,N_4154,N_5609);
nor U7342 (N_7342,N_3865,N_4480);
and U7343 (N_7343,N_5896,N_5338);
nand U7344 (N_7344,N_4066,N_3311);
and U7345 (N_7345,N_3752,N_5044);
or U7346 (N_7346,N_4386,N_4129);
and U7347 (N_7347,N_3930,N_3098);
nor U7348 (N_7348,N_4059,N_3410);
and U7349 (N_7349,N_4010,N_5879);
and U7350 (N_7350,N_5095,N_5170);
xnor U7351 (N_7351,N_4871,N_4022);
and U7352 (N_7352,N_4405,N_3912);
nand U7353 (N_7353,N_3166,N_3740);
nor U7354 (N_7354,N_3129,N_4967);
or U7355 (N_7355,N_5543,N_3838);
or U7356 (N_7356,N_5433,N_4840);
and U7357 (N_7357,N_5375,N_4775);
nor U7358 (N_7358,N_4495,N_4753);
or U7359 (N_7359,N_3102,N_3781);
xnor U7360 (N_7360,N_5995,N_3846);
and U7361 (N_7361,N_5121,N_5726);
nor U7362 (N_7362,N_4092,N_5275);
nand U7363 (N_7363,N_3681,N_3635);
nor U7364 (N_7364,N_4869,N_5573);
or U7365 (N_7365,N_5939,N_3758);
xor U7366 (N_7366,N_3599,N_4221);
nor U7367 (N_7367,N_3578,N_3332);
or U7368 (N_7368,N_5354,N_4306);
or U7369 (N_7369,N_5776,N_5516);
nor U7370 (N_7370,N_5339,N_5416);
nand U7371 (N_7371,N_4879,N_5920);
or U7372 (N_7372,N_5984,N_5929);
nor U7373 (N_7373,N_3690,N_5268);
nand U7374 (N_7374,N_3709,N_3339);
or U7375 (N_7375,N_5322,N_4065);
or U7376 (N_7376,N_4535,N_5191);
nand U7377 (N_7377,N_5957,N_5077);
nor U7378 (N_7378,N_4521,N_4737);
or U7379 (N_7379,N_5184,N_4616);
or U7380 (N_7380,N_3520,N_3310);
and U7381 (N_7381,N_5071,N_4946);
nor U7382 (N_7382,N_5222,N_4257);
or U7383 (N_7383,N_4863,N_4644);
nand U7384 (N_7384,N_5147,N_4167);
and U7385 (N_7385,N_5365,N_3885);
or U7386 (N_7386,N_3135,N_5992);
or U7387 (N_7387,N_5161,N_4420);
nand U7388 (N_7388,N_5412,N_4298);
and U7389 (N_7389,N_3600,N_4278);
nand U7390 (N_7390,N_5841,N_3193);
or U7391 (N_7391,N_4920,N_5996);
or U7392 (N_7392,N_3686,N_3057);
or U7393 (N_7393,N_3456,N_5389);
or U7394 (N_7394,N_4579,N_5853);
nand U7395 (N_7395,N_5948,N_3244);
and U7396 (N_7396,N_3340,N_5582);
or U7397 (N_7397,N_4161,N_4627);
nand U7398 (N_7398,N_3032,N_3016);
or U7399 (N_7399,N_4330,N_5409);
or U7400 (N_7400,N_3044,N_4334);
or U7401 (N_7401,N_3149,N_4760);
or U7402 (N_7402,N_5682,N_5143);
or U7403 (N_7403,N_4291,N_4803);
nand U7404 (N_7404,N_5873,N_5678);
and U7405 (N_7405,N_5430,N_5850);
xor U7406 (N_7406,N_4415,N_3441);
nand U7407 (N_7407,N_4932,N_3660);
or U7408 (N_7408,N_4331,N_3142);
or U7409 (N_7409,N_3527,N_5819);
and U7410 (N_7410,N_5787,N_5785);
and U7411 (N_7411,N_5382,N_3278);
and U7412 (N_7412,N_4915,N_3092);
nor U7413 (N_7413,N_5089,N_4200);
nor U7414 (N_7414,N_5036,N_3162);
nor U7415 (N_7415,N_3120,N_3916);
nor U7416 (N_7416,N_4889,N_5282);
or U7417 (N_7417,N_5665,N_4178);
nor U7418 (N_7418,N_5464,N_5290);
nor U7419 (N_7419,N_5436,N_3951);
nand U7420 (N_7420,N_5087,N_4390);
and U7421 (N_7421,N_4493,N_5931);
nor U7422 (N_7422,N_5058,N_4389);
or U7423 (N_7423,N_3586,N_4751);
or U7424 (N_7424,N_3261,N_4011);
nor U7425 (N_7425,N_5727,N_5251);
nor U7426 (N_7426,N_3231,N_3989);
nand U7427 (N_7427,N_5846,N_3952);
nor U7428 (N_7428,N_3668,N_4082);
or U7429 (N_7429,N_5355,N_5040);
and U7430 (N_7430,N_4588,N_3051);
nor U7431 (N_7431,N_4417,N_4783);
nand U7432 (N_7432,N_5197,N_5922);
nand U7433 (N_7433,N_4093,N_3710);
nand U7434 (N_7434,N_3859,N_4025);
or U7435 (N_7435,N_5083,N_3472);
nor U7436 (N_7436,N_3198,N_4419);
nor U7437 (N_7437,N_3420,N_4966);
or U7438 (N_7438,N_5406,N_4238);
or U7439 (N_7439,N_3480,N_4989);
and U7440 (N_7440,N_4519,N_4048);
nor U7441 (N_7441,N_5507,N_3053);
xor U7442 (N_7442,N_3844,N_3382);
nand U7443 (N_7443,N_4888,N_4656);
or U7444 (N_7444,N_3442,N_4045);
nand U7445 (N_7445,N_3360,N_4939);
nor U7446 (N_7446,N_5408,N_4508);
nor U7447 (N_7447,N_5503,N_3501);
or U7448 (N_7448,N_5473,N_4532);
nor U7449 (N_7449,N_5341,N_4149);
nand U7450 (N_7450,N_4593,N_4195);
nand U7451 (N_7451,N_4019,N_5715);
nor U7452 (N_7452,N_4468,N_4040);
or U7453 (N_7453,N_5649,N_5588);
nor U7454 (N_7454,N_4475,N_4259);
and U7455 (N_7455,N_3560,N_5910);
or U7456 (N_7456,N_5443,N_3395);
or U7457 (N_7457,N_4882,N_5631);
and U7458 (N_7458,N_5778,N_3949);
and U7459 (N_7459,N_4041,N_3170);
nand U7460 (N_7460,N_5384,N_3123);
and U7461 (N_7461,N_5857,N_3185);
and U7462 (N_7462,N_5937,N_3616);
and U7463 (N_7463,N_5980,N_5838);
or U7464 (N_7464,N_5589,N_4770);
and U7465 (N_7465,N_5818,N_4955);
nor U7466 (N_7466,N_4921,N_5065);
nand U7467 (N_7467,N_5797,N_3138);
nand U7468 (N_7468,N_4053,N_4499);
nor U7469 (N_7469,N_4980,N_3333);
nor U7470 (N_7470,N_4606,N_3626);
nor U7471 (N_7471,N_3861,N_4884);
nand U7472 (N_7472,N_3328,N_3582);
nand U7473 (N_7473,N_4553,N_3561);
nand U7474 (N_7474,N_3541,N_4528);
nor U7475 (N_7475,N_3732,N_5214);
and U7476 (N_7476,N_3575,N_3208);
and U7477 (N_7477,N_5895,N_5728);
nand U7478 (N_7478,N_4854,N_3862);
or U7479 (N_7479,N_4986,N_5504);
nand U7480 (N_7480,N_5798,N_4341);
and U7481 (N_7481,N_3214,N_3625);
nor U7482 (N_7482,N_3331,N_5938);
and U7483 (N_7483,N_3981,N_5868);
and U7484 (N_7484,N_4460,N_3287);
nor U7485 (N_7485,N_3628,N_5110);
nand U7486 (N_7486,N_3290,N_3685);
or U7487 (N_7487,N_5004,N_3377);
and U7488 (N_7488,N_4112,N_3486);
and U7489 (N_7489,N_3177,N_4276);
or U7490 (N_7490,N_4569,N_3236);
and U7491 (N_7491,N_3568,N_5075);
and U7492 (N_7492,N_4742,N_3896);
nor U7493 (N_7493,N_5872,N_3813);
or U7494 (N_7494,N_3488,N_5265);
and U7495 (N_7495,N_4910,N_4561);
nand U7496 (N_7496,N_3263,N_4271);
and U7497 (N_7497,N_4159,N_5830);
and U7498 (N_7498,N_3574,N_4020);
nand U7499 (N_7499,N_5333,N_3344);
and U7500 (N_7500,N_4217,N_4336);
and U7501 (N_7501,N_4605,N_4303);
nor U7502 (N_7502,N_4875,N_3269);
or U7503 (N_7503,N_5232,N_3881);
nand U7504 (N_7504,N_3706,N_3877);
and U7505 (N_7505,N_4441,N_5684);
nand U7506 (N_7506,N_4111,N_5008);
nand U7507 (N_7507,N_4256,N_3182);
or U7508 (N_7508,N_5972,N_3163);
and U7509 (N_7509,N_3261,N_5976);
nand U7510 (N_7510,N_4443,N_4864);
nand U7511 (N_7511,N_5446,N_4608);
or U7512 (N_7512,N_5596,N_4258);
nor U7513 (N_7513,N_3977,N_5545);
or U7514 (N_7514,N_3696,N_3133);
nand U7515 (N_7515,N_5972,N_5674);
nand U7516 (N_7516,N_3253,N_3958);
nand U7517 (N_7517,N_4459,N_4260);
and U7518 (N_7518,N_5542,N_4430);
and U7519 (N_7519,N_4648,N_4891);
nor U7520 (N_7520,N_5175,N_5322);
nand U7521 (N_7521,N_5691,N_3514);
or U7522 (N_7522,N_5042,N_3750);
nand U7523 (N_7523,N_5277,N_4655);
nand U7524 (N_7524,N_3689,N_4426);
nand U7525 (N_7525,N_5651,N_4663);
nand U7526 (N_7526,N_5320,N_4803);
nor U7527 (N_7527,N_4203,N_3372);
and U7528 (N_7528,N_4036,N_3341);
nand U7529 (N_7529,N_4552,N_5959);
and U7530 (N_7530,N_3688,N_4363);
or U7531 (N_7531,N_4510,N_3887);
nor U7532 (N_7532,N_5804,N_3123);
nand U7533 (N_7533,N_5191,N_4241);
nor U7534 (N_7534,N_5204,N_3325);
and U7535 (N_7535,N_4666,N_4927);
nor U7536 (N_7536,N_4924,N_4940);
and U7537 (N_7537,N_5209,N_4617);
nor U7538 (N_7538,N_3942,N_4714);
nor U7539 (N_7539,N_5287,N_4188);
nand U7540 (N_7540,N_5180,N_3178);
and U7541 (N_7541,N_4584,N_4033);
nor U7542 (N_7542,N_4615,N_3119);
or U7543 (N_7543,N_4450,N_3352);
and U7544 (N_7544,N_3976,N_3454);
nand U7545 (N_7545,N_4262,N_5313);
nand U7546 (N_7546,N_4913,N_4011);
and U7547 (N_7547,N_3787,N_5054);
nor U7548 (N_7548,N_4526,N_4098);
or U7549 (N_7549,N_5241,N_5164);
nor U7550 (N_7550,N_3647,N_5334);
and U7551 (N_7551,N_5060,N_4951);
and U7552 (N_7552,N_3638,N_4643);
and U7553 (N_7553,N_3900,N_3450);
nor U7554 (N_7554,N_5719,N_3651);
and U7555 (N_7555,N_5049,N_3751);
nor U7556 (N_7556,N_3540,N_3112);
and U7557 (N_7557,N_5382,N_3618);
nand U7558 (N_7558,N_5950,N_5670);
and U7559 (N_7559,N_3575,N_3535);
nand U7560 (N_7560,N_5037,N_3466);
or U7561 (N_7561,N_5314,N_4334);
or U7562 (N_7562,N_4539,N_5836);
nor U7563 (N_7563,N_3776,N_3766);
nor U7564 (N_7564,N_5215,N_4838);
or U7565 (N_7565,N_3532,N_5236);
nor U7566 (N_7566,N_5599,N_4412);
or U7567 (N_7567,N_4421,N_5252);
nand U7568 (N_7568,N_4104,N_4516);
nor U7569 (N_7569,N_5592,N_5595);
nand U7570 (N_7570,N_3361,N_3895);
nor U7571 (N_7571,N_3008,N_3282);
and U7572 (N_7572,N_5929,N_5558);
xnor U7573 (N_7573,N_3008,N_4724);
and U7574 (N_7574,N_5108,N_5182);
or U7575 (N_7575,N_3777,N_4331);
nor U7576 (N_7576,N_5612,N_4427);
and U7577 (N_7577,N_5817,N_5963);
or U7578 (N_7578,N_4711,N_5391);
or U7579 (N_7579,N_5922,N_4150);
and U7580 (N_7580,N_4744,N_4896);
nand U7581 (N_7581,N_4734,N_3689);
nand U7582 (N_7582,N_3982,N_5799);
nand U7583 (N_7583,N_5656,N_3367);
nor U7584 (N_7584,N_4437,N_5020);
nor U7585 (N_7585,N_5133,N_4494);
and U7586 (N_7586,N_4554,N_5880);
or U7587 (N_7587,N_4454,N_3657);
or U7588 (N_7588,N_5706,N_5761);
or U7589 (N_7589,N_5648,N_4123);
or U7590 (N_7590,N_4612,N_5012);
nor U7591 (N_7591,N_3837,N_4123);
or U7592 (N_7592,N_5583,N_3566);
and U7593 (N_7593,N_3860,N_5986);
nand U7594 (N_7594,N_4879,N_5466);
nor U7595 (N_7595,N_4462,N_4772);
xnor U7596 (N_7596,N_3792,N_4795);
or U7597 (N_7597,N_4826,N_3886);
or U7598 (N_7598,N_4196,N_5228);
and U7599 (N_7599,N_5062,N_5545);
nor U7600 (N_7600,N_3909,N_5822);
nand U7601 (N_7601,N_5655,N_4022);
or U7602 (N_7602,N_3473,N_3858);
and U7603 (N_7603,N_4138,N_5007);
and U7604 (N_7604,N_4378,N_4447);
or U7605 (N_7605,N_4994,N_4762);
and U7606 (N_7606,N_3028,N_5813);
nand U7607 (N_7607,N_3972,N_4596);
or U7608 (N_7608,N_3484,N_4440);
nor U7609 (N_7609,N_4448,N_5948);
nand U7610 (N_7610,N_3074,N_3721);
nor U7611 (N_7611,N_3263,N_4613);
or U7612 (N_7612,N_3145,N_3707);
and U7613 (N_7613,N_3957,N_5964);
nor U7614 (N_7614,N_4270,N_4018);
xnor U7615 (N_7615,N_3344,N_5673);
or U7616 (N_7616,N_3009,N_5105);
nor U7617 (N_7617,N_3255,N_4181);
nor U7618 (N_7618,N_5912,N_3146);
nor U7619 (N_7619,N_5943,N_5888);
nand U7620 (N_7620,N_5141,N_3239);
nor U7621 (N_7621,N_5079,N_3939);
nor U7622 (N_7622,N_5679,N_5384);
or U7623 (N_7623,N_4218,N_5278);
or U7624 (N_7624,N_5800,N_5460);
or U7625 (N_7625,N_4942,N_4749);
or U7626 (N_7626,N_4999,N_3395);
nand U7627 (N_7627,N_4787,N_3606);
nand U7628 (N_7628,N_4310,N_4976);
nor U7629 (N_7629,N_3487,N_3535);
nand U7630 (N_7630,N_3958,N_5389);
and U7631 (N_7631,N_4204,N_4791);
and U7632 (N_7632,N_3075,N_3562);
and U7633 (N_7633,N_3384,N_5070);
or U7634 (N_7634,N_3710,N_3461);
and U7635 (N_7635,N_4845,N_5327);
nor U7636 (N_7636,N_4863,N_4056);
nor U7637 (N_7637,N_5525,N_5997);
nor U7638 (N_7638,N_5318,N_4302);
or U7639 (N_7639,N_4275,N_4498);
nand U7640 (N_7640,N_3319,N_5443);
and U7641 (N_7641,N_4862,N_3734);
xnor U7642 (N_7642,N_4352,N_3203);
nand U7643 (N_7643,N_3546,N_5941);
nor U7644 (N_7644,N_5028,N_3824);
nor U7645 (N_7645,N_3737,N_5747);
or U7646 (N_7646,N_5130,N_3971);
nand U7647 (N_7647,N_4225,N_4344);
nor U7648 (N_7648,N_3773,N_4362);
and U7649 (N_7649,N_3552,N_5066);
nand U7650 (N_7650,N_4357,N_4510);
and U7651 (N_7651,N_4037,N_5571);
nor U7652 (N_7652,N_4930,N_5014);
and U7653 (N_7653,N_4786,N_4842);
nor U7654 (N_7654,N_3817,N_5980);
nand U7655 (N_7655,N_5177,N_5900);
or U7656 (N_7656,N_5731,N_3125);
and U7657 (N_7657,N_3129,N_4310);
nor U7658 (N_7658,N_4339,N_3669);
and U7659 (N_7659,N_3838,N_4471);
nand U7660 (N_7660,N_5329,N_5595);
nand U7661 (N_7661,N_3618,N_4675);
nand U7662 (N_7662,N_3039,N_5660);
or U7663 (N_7663,N_5617,N_5781);
and U7664 (N_7664,N_4977,N_5568);
or U7665 (N_7665,N_5863,N_4489);
nand U7666 (N_7666,N_3276,N_3313);
nand U7667 (N_7667,N_5705,N_5782);
and U7668 (N_7668,N_4848,N_3271);
or U7669 (N_7669,N_4113,N_5493);
nand U7670 (N_7670,N_4365,N_3195);
or U7671 (N_7671,N_3684,N_3141);
nand U7672 (N_7672,N_3964,N_3065);
or U7673 (N_7673,N_3886,N_3555);
nor U7674 (N_7674,N_3644,N_5036);
nor U7675 (N_7675,N_5674,N_4732);
nor U7676 (N_7676,N_4534,N_5906);
or U7677 (N_7677,N_3089,N_3020);
or U7678 (N_7678,N_4715,N_3706);
nor U7679 (N_7679,N_4926,N_3212);
nand U7680 (N_7680,N_5301,N_4343);
and U7681 (N_7681,N_3648,N_4653);
or U7682 (N_7682,N_5669,N_4686);
nand U7683 (N_7683,N_3731,N_3448);
or U7684 (N_7684,N_4289,N_4072);
nor U7685 (N_7685,N_5305,N_3412);
and U7686 (N_7686,N_5892,N_3459);
xnor U7687 (N_7687,N_4446,N_5441);
or U7688 (N_7688,N_5370,N_4778);
nor U7689 (N_7689,N_5831,N_3747);
xor U7690 (N_7690,N_3168,N_4048);
and U7691 (N_7691,N_3408,N_4468);
or U7692 (N_7692,N_5059,N_5408);
or U7693 (N_7693,N_3267,N_4431);
and U7694 (N_7694,N_5974,N_5559);
nand U7695 (N_7695,N_5746,N_5483);
nand U7696 (N_7696,N_5345,N_5727);
and U7697 (N_7697,N_3097,N_5063);
or U7698 (N_7698,N_4119,N_3372);
or U7699 (N_7699,N_3070,N_4562);
nand U7700 (N_7700,N_5598,N_4055);
and U7701 (N_7701,N_5514,N_4369);
and U7702 (N_7702,N_3064,N_5206);
or U7703 (N_7703,N_3431,N_5853);
nor U7704 (N_7704,N_5867,N_4124);
nor U7705 (N_7705,N_3259,N_4224);
and U7706 (N_7706,N_5989,N_5943);
or U7707 (N_7707,N_4387,N_5310);
and U7708 (N_7708,N_5110,N_4588);
and U7709 (N_7709,N_4205,N_5704);
nand U7710 (N_7710,N_4560,N_5340);
or U7711 (N_7711,N_5412,N_3128);
nor U7712 (N_7712,N_4770,N_4050);
or U7713 (N_7713,N_4592,N_3731);
or U7714 (N_7714,N_3990,N_3603);
nand U7715 (N_7715,N_4748,N_3772);
nand U7716 (N_7716,N_4755,N_5193);
nor U7717 (N_7717,N_4042,N_5890);
or U7718 (N_7718,N_3643,N_3401);
nor U7719 (N_7719,N_4971,N_5661);
or U7720 (N_7720,N_4874,N_5516);
nor U7721 (N_7721,N_3232,N_5785);
or U7722 (N_7722,N_3048,N_5603);
and U7723 (N_7723,N_3121,N_5534);
nor U7724 (N_7724,N_5193,N_3857);
nand U7725 (N_7725,N_5411,N_4975);
and U7726 (N_7726,N_3009,N_5821);
or U7727 (N_7727,N_5945,N_5260);
nand U7728 (N_7728,N_3739,N_5762);
nor U7729 (N_7729,N_4827,N_3900);
nor U7730 (N_7730,N_4966,N_4679);
nor U7731 (N_7731,N_5447,N_4394);
or U7732 (N_7732,N_4842,N_5737);
or U7733 (N_7733,N_4973,N_4501);
xor U7734 (N_7734,N_5263,N_4032);
or U7735 (N_7735,N_5365,N_5377);
and U7736 (N_7736,N_4509,N_3596);
and U7737 (N_7737,N_4196,N_3204);
nand U7738 (N_7738,N_5748,N_3510);
nand U7739 (N_7739,N_5591,N_3309);
nand U7740 (N_7740,N_4196,N_5166);
xor U7741 (N_7741,N_5042,N_3470);
or U7742 (N_7742,N_5446,N_3328);
nand U7743 (N_7743,N_5302,N_3368);
and U7744 (N_7744,N_5624,N_5379);
nor U7745 (N_7745,N_5773,N_3472);
nand U7746 (N_7746,N_4369,N_4493);
nand U7747 (N_7747,N_4247,N_4240);
and U7748 (N_7748,N_4442,N_5903);
and U7749 (N_7749,N_3579,N_4989);
nor U7750 (N_7750,N_3988,N_3098);
nor U7751 (N_7751,N_4705,N_4164);
and U7752 (N_7752,N_5132,N_4119);
and U7753 (N_7753,N_3249,N_4798);
or U7754 (N_7754,N_5515,N_5344);
nand U7755 (N_7755,N_3769,N_5441);
nor U7756 (N_7756,N_5365,N_5934);
or U7757 (N_7757,N_5672,N_5599);
or U7758 (N_7758,N_3581,N_3012);
or U7759 (N_7759,N_5716,N_4668);
nor U7760 (N_7760,N_3459,N_4964);
nand U7761 (N_7761,N_5190,N_5361);
or U7762 (N_7762,N_5196,N_3201);
and U7763 (N_7763,N_5975,N_3612);
nor U7764 (N_7764,N_3561,N_5402);
and U7765 (N_7765,N_4931,N_4291);
or U7766 (N_7766,N_3495,N_4142);
nand U7767 (N_7767,N_3463,N_3669);
and U7768 (N_7768,N_4697,N_5055);
nand U7769 (N_7769,N_3791,N_5054);
nand U7770 (N_7770,N_5211,N_5650);
nand U7771 (N_7771,N_4838,N_5782);
or U7772 (N_7772,N_3863,N_3257);
nor U7773 (N_7773,N_3349,N_5376);
and U7774 (N_7774,N_4195,N_5986);
nor U7775 (N_7775,N_4526,N_3121);
and U7776 (N_7776,N_4628,N_4277);
nand U7777 (N_7777,N_4423,N_4244);
and U7778 (N_7778,N_5841,N_4673);
nand U7779 (N_7779,N_3165,N_5054);
nor U7780 (N_7780,N_4254,N_5973);
or U7781 (N_7781,N_5981,N_3700);
or U7782 (N_7782,N_3754,N_3234);
nand U7783 (N_7783,N_3231,N_3715);
nand U7784 (N_7784,N_3462,N_3047);
nor U7785 (N_7785,N_4738,N_3147);
nand U7786 (N_7786,N_5064,N_5288);
nor U7787 (N_7787,N_4502,N_3044);
nand U7788 (N_7788,N_5448,N_3911);
or U7789 (N_7789,N_3435,N_3959);
xor U7790 (N_7790,N_5839,N_3440);
and U7791 (N_7791,N_5725,N_4244);
nand U7792 (N_7792,N_3588,N_5390);
and U7793 (N_7793,N_4300,N_4653);
nand U7794 (N_7794,N_3564,N_5196);
nand U7795 (N_7795,N_4128,N_4239);
and U7796 (N_7796,N_4278,N_3993);
and U7797 (N_7797,N_3831,N_3416);
nor U7798 (N_7798,N_4913,N_5495);
or U7799 (N_7799,N_4524,N_3186);
xnor U7800 (N_7800,N_4021,N_5191);
nor U7801 (N_7801,N_3507,N_4315);
and U7802 (N_7802,N_5575,N_3999);
nand U7803 (N_7803,N_4105,N_3365);
and U7804 (N_7804,N_5560,N_4284);
and U7805 (N_7805,N_3495,N_3056);
nor U7806 (N_7806,N_4898,N_3854);
or U7807 (N_7807,N_4444,N_4645);
and U7808 (N_7808,N_4916,N_3442);
or U7809 (N_7809,N_5646,N_3614);
nor U7810 (N_7810,N_4707,N_4833);
nor U7811 (N_7811,N_4676,N_5352);
and U7812 (N_7812,N_5895,N_3591);
nor U7813 (N_7813,N_3137,N_5085);
or U7814 (N_7814,N_4165,N_3186);
or U7815 (N_7815,N_4126,N_3282);
or U7816 (N_7816,N_4874,N_3734);
and U7817 (N_7817,N_4960,N_4325);
nor U7818 (N_7818,N_3928,N_5337);
nand U7819 (N_7819,N_3541,N_5044);
nor U7820 (N_7820,N_3583,N_3461);
or U7821 (N_7821,N_5334,N_4145);
xor U7822 (N_7822,N_3500,N_4924);
and U7823 (N_7823,N_5045,N_5879);
and U7824 (N_7824,N_4857,N_5829);
and U7825 (N_7825,N_4004,N_3937);
nand U7826 (N_7826,N_3746,N_4985);
nor U7827 (N_7827,N_4388,N_3562);
nor U7828 (N_7828,N_5047,N_4855);
nor U7829 (N_7829,N_4691,N_5781);
or U7830 (N_7830,N_4462,N_3024);
nor U7831 (N_7831,N_4197,N_3417);
or U7832 (N_7832,N_5919,N_3836);
and U7833 (N_7833,N_3220,N_4351);
nand U7834 (N_7834,N_4264,N_3992);
or U7835 (N_7835,N_5206,N_4277);
nand U7836 (N_7836,N_3686,N_3883);
nor U7837 (N_7837,N_4650,N_5799);
nand U7838 (N_7838,N_4345,N_4457);
nor U7839 (N_7839,N_5459,N_4270);
and U7840 (N_7840,N_4962,N_4778);
nand U7841 (N_7841,N_4286,N_3619);
or U7842 (N_7842,N_4200,N_4062);
or U7843 (N_7843,N_5205,N_3405);
and U7844 (N_7844,N_5442,N_4890);
xor U7845 (N_7845,N_4496,N_3412);
nor U7846 (N_7846,N_4650,N_5131);
or U7847 (N_7847,N_4361,N_3964);
nand U7848 (N_7848,N_4074,N_4674);
nand U7849 (N_7849,N_4268,N_4706);
nor U7850 (N_7850,N_5226,N_3687);
nor U7851 (N_7851,N_5380,N_5749);
nor U7852 (N_7852,N_4053,N_5442);
nor U7853 (N_7853,N_3479,N_3638);
or U7854 (N_7854,N_4681,N_3720);
nand U7855 (N_7855,N_3858,N_5497);
and U7856 (N_7856,N_3274,N_5551);
nor U7857 (N_7857,N_5521,N_3536);
nor U7858 (N_7858,N_4326,N_5544);
or U7859 (N_7859,N_3418,N_4460);
or U7860 (N_7860,N_4003,N_4200);
and U7861 (N_7861,N_4107,N_3255);
nor U7862 (N_7862,N_5305,N_5256);
nand U7863 (N_7863,N_5974,N_3102);
or U7864 (N_7864,N_3850,N_4331);
or U7865 (N_7865,N_5332,N_4451);
and U7866 (N_7866,N_5330,N_3265);
nand U7867 (N_7867,N_3999,N_3799);
and U7868 (N_7868,N_5882,N_4776);
or U7869 (N_7869,N_5669,N_4770);
and U7870 (N_7870,N_5463,N_4657);
and U7871 (N_7871,N_3783,N_3273);
nand U7872 (N_7872,N_5856,N_3314);
or U7873 (N_7873,N_5748,N_5994);
nor U7874 (N_7874,N_3720,N_5303);
or U7875 (N_7875,N_3676,N_4930);
nand U7876 (N_7876,N_4714,N_3144);
nand U7877 (N_7877,N_3413,N_3805);
nor U7878 (N_7878,N_3496,N_5134);
nor U7879 (N_7879,N_4822,N_3508);
nor U7880 (N_7880,N_5390,N_3303);
and U7881 (N_7881,N_5607,N_4780);
xnor U7882 (N_7882,N_4171,N_5375);
or U7883 (N_7883,N_4596,N_3030);
and U7884 (N_7884,N_5860,N_4119);
nand U7885 (N_7885,N_4615,N_4408);
and U7886 (N_7886,N_3135,N_5000);
nand U7887 (N_7887,N_5397,N_3172);
or U7888 (N_7888,N_5369,N_4958);
nand U7889 (N_7889,N_4518,N_3041);
nor U7890 (N_7890,N_4993,N_5012);
nor U7891 (N_7891,N_4711,N_4543);
and U7892 (N_7892,N_5505,N_5626);
or U7893 (N_7893,N_4444,N_5342);
or U7894 (N_7894,N_4899,N_5175);
nand U7895 (N_7895,N_4312,N_4481);
nand U7896 (N_7896,N_3095,N_3309);
nand U7897 (N_7897,N_3555,N_4980);
or U7898 (N_7898,N_4787,N_3944);
nor U7899 (N_7899,N_4952,N_5548);
nand U7900 (N_7900,N_3566,N_5914);
or U7901 (N_7901,N_4794,N_5023);
and U7902 (N_7902,N_4937,N_3678);
or U7903 (N_7903,N_4130,N_4843);
nor U7904 (N_7904,N_5679,N_3602);
nand U7905 (N_7905,N_5718,N_3574);
nand U7906 (N_7906,N_5955,N_4819);
or U7907 (N_7907,N_4095,N_5130);
nand U7908 (N_7908,N_5728,N_3934);
nor U7909 (N_7909,N_5500,N_3662);
or U7910 (N_7910,N_3053,N_4857);
xnor U7911 (N_7911,N_3582,N_5951);
nor U7912 (N_7912,N_5263,N_3290);
or U7913 (N_7913,N_4376,N_5839);
or U7914 (N_7914,N_4553,N_4673);
xor U7915 (N_7915,N_4537,N_4951);
and U7916 (N_7916,N_3145,N_4196);
nand U7917 (N_7917,N_4392,N_4830);
or U7918 (N_7918,N_3664,N_4734);
nand U7919 (N_7919,N_3000,N_3494);
or U7920 (N_7920,N_3026,N_4144);
nor U7921 (N_7921,N_5391,N_4089);
nand U7922 (N_7922,N_4254,N_3687);
or U7923 (N_7923,N_3583,N_5701);
nor U7924 (N_7924,N_3281,N_3702);
and U7925 (N_7925,N_3440,N_4351);
nand U7926 (N_7926,N_3593,N_3590);
or U7927 (N_7927,N_5774,N_4472);
and U7928 (N_7928,N_4722,N_4475);
nand U7929 (N_7929,N_3099,N_4848);
nor U7930 (N_7930,N_5248,N_4246);
nand U7931 (N_7931,N_4006,N_3008);
xnor U7932 (N_7932,N_3892,N_4097);
nor U7933 (N_7933,N_5564,N_3126);
nand U7934 (N_7934,N_4002,N_5570);
or U7935 (N_7935,N_3217,N_3847);
or U7936 (N_7936,N_5396,N_4238);
nor U7937 (N_7937,N_3518,N_3713);
and U7938 (N_7938,N_3756,N_5533);
or U7939 (N_7939,N_4648,N_3158);
nand U7940 (N_7940,N_4984,N_5687);
nor U7941 (N_7941,N_5935,N_5619);
or U7942 (N_7942,N_3851,N_3423);
nor U7943 (N_7943,N_5422,N_3706);
or U7944 (N_7944,N_3478,N_4152);
and U7945 (N_7945,N_3234,N_5832);
or U7946 (N_7946,N_3181,N_4164);
xnor U7947 (N_7947,N_3613,N_3734);
nor U7948 (N_7948,N_5579,N_4474);
nor U7949 (N_7949,N_3320,N_4708);
or U7950 (N_7950,N_5071,N_3419);
and U7951 (N_7951,N_3489,N_3978);
or U7952 (N_7952,N_4284,N_4574);
nand U7953 (N_7953,N_5374,N_5510);
nand U7954 (N_7954,N_4301,N_3832);
or U7955 (N_7955,N_4492,N_5614);
xor U7956 (N_7956,N_3581,N_5063);
or U7957 (N_7957,N_4564,N_5934);
nor U7958 (N_7958,N_5482,N_5685);
or U7959 (N_7959,N_4187,N_3439);
and U7960 (N_7960,N_3553,N_5310);
nor U7961 (N_7961,N_4650,N_4687);
or U7962 (N_7962,N_4986,N_5123);
nand U7963 (N_7963,N_5775,N_4709);
nor U7964 (N_7964,N_5522,N_3615);
nand U7965 (N_7965,N_4959,N_3076);
nand U7966 (N_7966,N_5621,N_5840);
or U7967 (N_7967,N_5114,N_5842);
nor U7968 (N_7968,N_4780,N_4617);
nand U7969 (N_7969,N_5014,N_4571);
nand U7970 (N_7970,N_5726,N_3730);
or U7971 (N_7971,N_5816,N_3359);
or U7972 (N_7972,N_4440,N_5013);
or U7973 (N_7973,N_3347,N_3737);
nand U7974 (N_7974,N_3362,N_4894);
or U7975 (N_7975,N_4825,N_5358);
or U7976 (N_7976,N_4947,N_4262);
and U7977 (N_7977,N_4819,N_3415);
nand U7978 (N_7978,N_5609,N_4697);
nand U7979 (N_7979,N_5153,N_4499);
and U7980 (N_7980,N_4922,N_3131);
nor U7981 (N_7981,N_5460,N_5967);
or U7982 (N_7982,N_3762,N_4098);
nand U7983 (N_7983,N_5619,N_4191);
and U7984 (N_7984,N_3112,N_5143);
or U7985 (N_7985,N_4262,N_5365);
or U7986 (N_7986,N_5518,N_5131);
nand U7987 (N_7987,N_4684,N_4353);
and U7988 (N_7988,N_3834,N_5917);
or U7989 (N_7989,N_5403,N_3927);
nand U7990 (N_7990,N_5182,N_3291);
nor U7991 (N_7991,N_3503,N_3376);
nand U7992 (N_7992,N_4325,N_4269);
nand U7993 (N_7993,N_3676,N_3868);
and U7994 (N_7994,N_5940,N_4759);
nand U7995 (N_7995,N_5920,N_5439);
nor U7996 (N_7996,N_5525,N_3520);
and U7997 (N_7997,N_4362,N_3316);
and U7998 (N_7998,N_4462,N_3184);
nand U7999 (N_7999,N_3797,N_4089);
and U8000 (N_8000,N_3286,N_3588);
nor U8001 (N_8001,N_5662,N_4285);
nand U8002 (N_8002,N_4570,N_4995);
nand U8003 (N_8003,N_3857,N_3225);
or U8004 (N_8004,N_4839,N_5321);
nor U8005 (N_8005,N_4806,N_4617);
nand U8006 (N_8006,N_5329,N_5245);
or U8007 (N_8007,N_3546,N_4717);
and U8008 (N_8008,N_4973,N_4060);
or U8009 (N_8009,N_5576,N_3812);
nor U8010 (N_8010,N_5522,N_3614);
nand U8011 (N_8011,N_5379,N_3511);
nand U8012 (N_8012,N_3482,N_4407);
and U8013 (N_8013,N_4781,N_3068);
nor U8014 (N_8014,N_5686,N_4638);
nand U8015 (N_8015,N_3889,N_5531);
and U8016 (N_8016,N_4762,N_4071);
or U8017 (N_8017,N_5667,N_5718);
nor U8018 (N_8018,N_4061,N_4606);
nor U8019 (N_8019,N_3724,N_4190);
or U8020 (N_8020,N_4939,N_4360);
nand U8021 (N_8021,N_5553,N_3267);
or U8022 (N_8022,N_3564,N_4289);
and U8023 (N_8023,N_3400,N_3717);
nand U8024 (N_8024,N_4887,N_3976);
nand U8025 (N_8025,N_4932,N_4778);
and U8026 (N_8026,N_5912,N_3577);
nand U8027 (N_8027,N_5506,N_4659);
and U8028 (N_8028,N_5939,N_5113);
and U8029 (N_8029,N_4008,N_4063);
xor U8030 (N_8030,N_3691,N_5128);
nand U8031 (N_8031,N_3630,N_3006);
or U8032 (N_8032,N_3322,N_5783);
nand U8033 (N_8033,N_5742,N_4730);
nor U8034 (N_8034,N_5753,N_4762);
and U8035 (N_8035,N_3791,N_5565);
nor U8036 (N_8036,N_3370,N_5468);
nor U8037 (N_8037,N_5814,N_4035);
and U8038 (N_8038,N_3153,N_5379);
nand U8039 (N_8039,N_4919,N_5103);
nand U8040 (N_8040,N_5956,N_3610);
or U8041 (N_8041,N_3133,N_4807);
and U8042 (N_8042,N_5639,N_4749);
or U8043 (N_8043,N_3750,N_4663);
or U8044 (N_8044,N_3384,N_4018);
and U8045 (N_8045,N_4490,N_5371);
or U8046 (N_8046,N_4199,N_5248);
nor U8047 (N_8047,N_3947,N_3291);
or U8048 (N_8048,N_5811,N_3678);
nand U8049 (N_8049,N_5748,N_4487);
nand U8050 (N_8050,N_4496,N_3279);
xor U8051 (N_8051,N_3812,N_5273);
nor U8052 (N_8052,N_3495,N_4683);
or U8053 (N_8053,N_3103,N_5548);
nand U8054 (N_8054,N_3585,N_3898);
and U8055 (N_8055,N_4410,N_4370);
nand U8056 (N_8056,N_4151,N_4261);
or U8057 (N_8057,N_4550,N_3839);
nand U8058 (N_8058,N_5683,N_3334);
and U8059 (N_8059,N_4749,N_5524);
nand U8060 (N_8060,N_4709,N_4411);
or U8061 (N_8061,N_3946,N_5677);
and U8062 (N_8062,N_5951,N_5704);
nand U8063 (N_8063,N_3592,N_5750);
nor U8064 (N_8064,N_3934,N_5762);
nor U8065 (N_8065,N_4346,N_5971);
and U8066 (N_8066,N_5367,N_3846);
and U8067 (N_8067,N_5965,N_5239);
or U8068 (N_8068,N_3794,N_4155);
nor U8069 (N_8069,N_3054,N_3357);
nor U8070 (N_8070,N_5403,N_4308);
nand U8071 (N_8071,N_4223,N_3526);
nor U8072 (N_8072,N_5915,N_5791);
and U8073 (N_8073,N_3791,N_5862);
and U8074 (N_8074,N_4280,N_4889);
and U8075 (N_8075,N_4243,N_4524);
xor U8076 (N_8076,N_5411,N_4739);
and U8077 (N_8077,N_5702,N_4143);
and U8078 (N_8078,N_3235,N_4512);
nor U8079 (N_8079,N_4710,N_3813);
and U8080 (N_8080,N_3564,N_5518);
and U8081 (N_8081,N_4163,N_5785);
nand U8082 (N_8082,N_5589,N_4309);
and U8083 (N_8083,N_3560,N_3608);
nand U8084 (N_8084,N_4381,N_3201);
nand U8085 (N_8085,N_4022,N_5054);
or U8086 (N_8086,N_3794,N_4769);
xnor U8087 (N_8087,N_3529,N_4829);
nand U8088 (N_8088,N_5204,N_5570);
xnor U8089 (N_8089,N_4800,N_4842);
or U8090 (N_8090,N_5032,N_5886);
and U8091 (N_8091,N_3471,N_5809);
nand U8092 (N_8092,N_4010,N_5994);
and U8093 (N_8093,N_5420,N_5001);
and U8094 (N_8094,N_3618,N_4252);
and U8095 (N_8095,N_5655,N_3920);
or U8096 (N_8096,N_4709,N_3834);
xnor U8097 (N_8097,N_4437,N_3943);
nand U8098 (N_8098,N_5210,N_3729);
or U8099 (N_8099,N_3417,N_5709);
nand U8100 (N_8100,N_5703,N_4394);
or U8101 (N_8101,N_4278,N_3943);
nor U8102 (N_8102,N_5347,N_3126);
and U8103 (N_8103,N_5456,N_5505);
nor U8104 (N_8104,N_3669,N_5596);
and U8105 (N_8105,N_4699,N_5127);
or U8106 (N_8106,N_5996,N_5670);
nand U8107 (N_8107,N_3386,N_4869);
nand U8108 (N_8108,N_5974,N_5776);
or U8109 (N_8109,N_3989,N_5367);
and U8110 (N_8110,N_3608,N_5899);
nand U8111 (N_8111,N_5627,N_3097);
nand U8112 (N_8112,N_5391,N_3848);
and U8113 (N_8113,N_5306,N_3272);
and U8114 (N_8114,N_5550,N_4680);
or U8115 (N_8115,N_5224,N_4397);
or U8116 (N_8116,N_3183,N_5734);
nor U8117 (N_8117,N_4581,N_4033);
and U8118 (N_8118,N_4661,N_3973);
and U8119 (N_8119,N_5438,N_3777);
or U8120 (N_8120,N_3455,N_3389);
nor U8121 (N_8121,N_5618,N_3034);
nor U8122 (N_8122,N_4974,N_4122);
nor U8123 (N_8123,N_3295,N_3426);
and U8124 (N_8124,N_5665,N_5224);
xor U8125 (N_8125,N_3529,N_5929);
and U8126 (N_8126,N_3583,N_5015);
and U8127 (N_8127,N_5953,N_5777);
or U8128 (N_8128,N_5745,N_5132);
and U8129 (N_8129,N_3438,N_4993);
or U8130 (N_8130,N_5788,N_5798);
and U8131 (N_8131,N_5748,N_4411);
and U8132 (N_8132,N_3432,N_3291);
and U8133 (N_8133,N_4293,N_4942);
xnor U8134 (N_8134,N_3920,N_5024);
nand U8135 (N_8135,N_3153,N_4652);
nor U8136 (N_8136,N_5884,N_5083);
nor U8137 (N_8137,N_5165,N_3005);
nand U8138 (N_8138,N_5341,N_3329);
or U8139 (N_8139,N_4932,N_4928);
and U8140 (N_8140,N_5926,N_3913);
nand U8141 (N_8141,N_4424,N_5176);
and U8142 (N_8142,N_4908,N_5207);
nor U8143 (N_8143,N_5113,N_3661);
and U8144 (N_8144,N_3177,N_5641);
nor U8145 (N_8145,N_4697,N_3859);
or U8146 (N_8146,N_5558,N_3520);
and U8147 (N_8147,N_3203,N_4161);
nand U8148 (N_8148,N_3922,N_5932);
nand U8149 (N_8149,N_4843,N_4288);
and U8150 (N_8150,N_3095,N_3740);
and U8151 (N_8151,N_3243,N_3204);
and U8152 (N_8152,N_3221,N_4009);
xnor U8153 (N_8153,N_4867,N_4922);
nor U8154 (N_8154,N_5283,N_3977);
nand U8155 (N_8155,N_3004,N_3003);
or U8156 (N_8156,N_3102,N_3503);
or U8157 (N_8157,N_4899,N_3596);
nor U8158 (N_8158,N_5714,N_5144);
or U8159 (N_8159,N_5916,N_4218);
nor U8160 (N_8160,N_5954,N_5284);
xor U8161 (N_8161,N_3199,N_4620);
and U8162 (N_8162,N_3181,N_4446);
nor U8163 (N_8163,N_3833,N_3261);
nand U8164 (N_8164,N_5377,N_5459);
nand U8165 (N_8165,N_5461,N_3807);
nor U8166 (N_8166,N_5048,N_4429);
and U8167 (N_8167,N_4062,N_4087);
and U8168 (N_8168,N_3431,N_3850);
nand U8169 (N_8169,N_5867,N_5662);
nor U8170 (N_8170,N_5022,N_5029);
and U8171 (N_8171,N_5505,N_3045);
nand U8172 (N_8172,N_5710,N_4678);
or U8173 (N_8173,N_3282,N_4890);
or U8174 (N_8174,N_5183,N_4234);
or U8175 (N_8175,N_4865,N_3159);
and U8176 (N_8176,N_3094,N_4236);
or U8177 (N_8177,N_4782,N_4650);
xnor U8178 (N_8178,N_4646,N_3924);
nand U8179 (N_8179,N_5803,N_5743);
nor U8180 (N_8180,N_5712,N_4672);
nor U8181 (N_8181,N_4112,N_5831);
or U8182 (N_8182,N_3834,N_5713);
and U8183 (N_8183,N_3498,N_4249);
or U8184 (N_8184,N_5576,N_4068);
nor U8185 (N_8185,N_4320,N_3450);
and U8186 (N_8186,N_5531,N_4130);
nand U8187 (N_8187,N_4404,N_5881);
or U8188 (N_8188,N_5389,N_5111);
and U8189 (N_8189,N_4124,N_4718);
nand U8190 (N_8190,N_4551,N_3884);
or U8191 (N_8191,N_4423,N_5272);
nand U8192 (N_8192,N_5183,N_5664);
nand U8193 (N_8193,N_4910,N_4680);
or U8194 (N_8194,N_3197,N_5124);
and U8195 (N_8195,N_4591,N_4555);
and U8196 (N_8196,N_4345,N_4871);
nand U8197 (N_8197,N_3541,N_5931);
or U8198 (N_8198,N_5465,N_3045);
and U8199 (N_8199,N_3983,N_4811);
nor U8200 (N_8200,N_5628,N_3869);
nor U8201 (N_8201,N_3837,N_5010);
and U8202 (N_8202,N_3886,N_4667);
or U8203 (N_8203,N_3369,N_4838);
or U8204 (N_8204,N_3149,N_4488);
nand U8205 (N_8205,N_3649,N_3362);
and U8206 (N_8206,N_5136,N_5535);
or U8207 (N_8207,N_5868,N_3671);
nor U8208 (N_8208,N_5464,N_4081);
or U8209 (N_8209,N_3458,N_3681);
nand U8210 (N_8210,N_5384,N_3263);
nand U8211 (N_8211,N_5913,N_5530);
and U8212 (N_8212,N_4883,N_3576);
nor U8213 (N_8213,N_4659,N_4041);
and U8214 (N_8214,N_4311,N_5809);
nand U8215 (N_8215,N_3212,N_3961);
or U8216 (N_8216,N_3292,N_5064);
nor U8217 (N_8217,N_4860,N_5301);
nor U8218 (N_8218,N_4617,N_5152);
or U8219 (N_8219,N_3511,N_5264);
and U8220 (N_8220,N_3811,N_4987);
or U8221 (N_8221,N_3451,N_4887);
nor U8222 (N_8222,N_4348,N_5564);
nor U8223 (N_8223,N_4119,N_4802);
nand U8224 (N_8224,N_4294,N_5300);
or U8225 (N_8225,N_5362,N_5922);
or U8226 (N_8226,N_3775,N_5930);
and U8227 (N_8227,N_5997,N_5623);
nand U8228 (N_8228,N_3833,N_4949);
nor U8229 (N_8229,N_3358,N_3192);
nor U8230 (N_8230,N_3814,N_4232);
or U8231 (N_8231,N_3754,N_5693);
nand U8232 (N_8232,N_4591,N_4723);
nor U8233 (N_8233,N_4161,N_5314);
and U8234 (N_8234,N_4421,N_5732);
and U8235 (N_8235,N_4316,N_5323);
or U8236 (N_8236,N_3687,N_3738);
nor U8237 (N_8237,N_4804,N_4147);
xnor U8238 (N_8238,N_5483,N_3883);
nor U8239 (N_8239,N_4917,N_3798);
nor U8240 (N_8240,N_5974,N_5210);
nand U8241 (N_8241,N_5288,N_5323);
nor U8242 (N_8242,N_4843,N_3897);
and U8243 (N_8243,N_4141,N_5079);
nand U8244 (N_8244,N_3278,N_4798);
nor U8245 (N_8245,N_3704,N_3731);
nand U8246 (N_8246,N_5899,N_5075);
and U8247 (N_8247,N_3875,N_5679);
nand U8248 (N_8248,N_4225,N_4591);
or U8249 (N_8249,N_3774,N_3221);
nor U8250 (N_8250,N_4176,N_3489);
nor U8251 (N_8251,N_4735,N_3517);
or U8252 (N_8252,N_3138,N_4378);
nand U8253 (N_8253,N_5128,N_4994);
nor U8254 (N_8254,N_5746,N_3568);
nand U8255 (N_8255,N_5802,N_5096);
or U8256 (N_8256,N_4347,N_3929);
nor U8257 (N_8257,N_5097,N_4600);
nor U8258 (N_8258,N_3237,N_3299);
or U8259 (N_8259,N_5869,N_3635);
and U8260 (N_8260,N_5006,N_5009);
nand U8261 (N_8261,N_5989,N_4155);
or U8262 (N_8262,N_5661,N_3188);
or U8263 (N_8263,N_4978,N_4510);
nand U8264 (N_8264,N_3084,N_3832);
and U8265 (N_8265,N_5035,N_3350);
and U8266 (N_8266,N_5578,N_5958);
nand U8267 (N_8267,N_5215,N_5305);
nor U8268 (N_8268,N_5801,N_3946);
nand U8269 (N_8269,N_5265,N_4309);
and U8270 (N_8270,N_3450,N_3980);
nor U8271 (N_8271,N_5325,N_3993);
and U8272 (N_8272,N_3264,N_3245);
or U8273 (N_8273,N_3930,N_3245);
and U8274 (N_8274,N_4664,N_4761);
nor U8275 (N_8275,N_3927,N_4529);
and U8276 (N_8276,N_5464,N_3783);
nor U8277 (N_8277,N_3615,N_4416);
nor U8278 (N_8278,N_3979,N_5933);
and U8279 (N_8279,N_3695,N_3186);
nand U8280 (N_8280,N_5527,N_3441);
and U8281 (N_8281,N_5352,N_3360);
or U8282 (N_8282,N_5356,N_5663);
and U8283 (N_8283,N_5469,N_5287);
and U8284 (N_8284,N_4943,N_3016);
or U8285 (N_8285,N_5355,N_4808);
and U8286 (N_8286,N_4683,N_3721);
and U8287 (N_8287,N_5850,N_5299);
nor U8288 (N_8288,N_4131,N_4834);
xnor U8289 (N_8289,N_3643,N_4961);
or U8290 (N_8290,N_5394,N_4459);
nor U8291 (N_8291,N_3870,N_3269);
or U8292 (N_8292,N_4750,N_3333);
and U8293 (N_8293,N_4392,N_4287);
or U8294 (N_8294,N_3123,N_5762);
nand U8295 (N_8295,N_5625,N_4377);
and U8296 (N_8296,N_3186,N_3871);
and U8297 (N_8297,N_5439,N_5714);
xnor U8298 (N_8298,N_5950,N_5997);
nor U8299 (N_8299,N_3223,N_3961);
nand U8300 (N_8300,N_5307,N_3999);
and U8301 (N_8301,N_4913,N_3256);
or U8302 (N_8302,N_5293,N_4122);
nand U8303 (N_8303,N_4067,N_5590);
and U8304 (N_8304,N_4993,N_4695);
nand U8305 (N_8305,N_4678,N_4397);
nand U8306 (N_8306,N_4920,N_3236);
nor U8307 (N_8307,N_5040,N_5506);
or U8308 (N_8308,N_4947,N_3989);
nor U8309 (N_8309,N_5469,N_3093);
or U8310 (N_8310,N_4998,N_4600);
nand U8311 (N_8311,N_4420,N_5724);
nand U8312 (N_8312,N_3889,N_3471);
and U8313 (N_8313,N_4368,N_3563);
or U8314 (N_8314,N_3334,N_4497);
and U8315 (N_8315,N_4338,N_5777);
nand U8316 (N_8316,N_3523,N_3270);
nand U8317 (N_8317,N_3708,N_5533);
nor U8318 (N_8318,N_5539,N_4063);
or U8319 (N_8319,N_3242,N_3978);
and U8320 (N_8320,N_5050,N_4433);
nand U8321 (N_8321,N_5409,N_4907);
or U8322 (N_8322,N_5756,N_3640);
and U8323 (N_8323,N_4931,N_5734);
nor U8324 (N_8324,N_5918,N_5229);
nand U8325 (N_8325,N_5546,N_5009);
nand U8326 (N_8326,N_4990,N_5041);
or U8327 (N_8327,N_4831,N_3053);
or U8328 (N_8328,N_3767,N_3339);
or U8329 (N_8329,N_4328,N_4396);
and U8330 (N_8330,N_4111,N_5801);
or U8331 (N_8331,N_4086,N_3609);
nand U8332 (N_8332,N_5696,N_4366);
or U8333 (N_8333,N_5281,N_4224);
and U8334 (N_8334,N_3989,N_4466);
nor U8335 (N_8335,N_4345,N_4226);
and U8336 (N_8336,N_4082,N_5465);
nand U8337 (N_8337,N_5172,N_3005);
or U8338 (N_8338,N_3594,N_4673);
and U8339 (N_8339,N_4768,N_3581);
and U8340 (N_8340,N_4780,N_3421);
and U8341 (N_8341,N_3638,N_3658);
or U8342 (N_8342,N_5336,N_3207);
nand U8343 (N_8343,N_3567,N_4497);
nor U8344 (N_8344,N_3612,N_5418);
nand U8345 (N_8345,N_4639,N_5082);
or U8346 (N_8346,N_3839,N_5931);
nor U8347 (N_8347,N_5560,N_5318);
nor U8348 (N_8348,N_3578,N_3023);
nand U8349 (N_8349,N_3778,N_3994);
or U8350 (N_8350,N_3065,N_4792);
or U8351 (N_8351,N_4803,N_5512);
and U8352 (N_8352,N_5980,N_4206);
or U8353 (N_8353,N_4436,N_5960);
nor U8354 (N_8354,N_5477,N_4369);
nor U8355 (N_8355,N_4906,N_4230);
nor U8356 (N_8356,N_5164,N_4378);
and U8357 (N_8357,N_4600,N_3853);
or U8358 (N_8358,N_4891,N_5273);
nand U8359 (N_8359,N_3486,N_4497);
nor U8360 (N_8360,N_4194,N_3540);
nor U8361 (N_8361,N_3991,N_4417);
nand U8362 (N_8362,N_5851,N_5810);
nand U8363 (N_8363,N_5971,N_3331);
nand U8364 (N_8364,N_3338,N_4456);
or U8365 (N_8365,N_3305,N_5433);
nor U8366 (N_8366,N_4138,N_3105);
nand U8367 (N_8367,N_5989,N_3333);
and U8368 (N_8368,N_3001,N_5947);
nand U8369 (N_8369,N_4908,N_5280);
nand U8370 (N_8370,N_4761,N_5403);
and U8371 (N_8371,N_3862,N_3832);
nor U8372 (N_8372,N_5318,N_5870);
or U8373 (N_8373,N_3690,N_4029);
nand U8374 (N_8374,N_5074,N_4599);
nand U8375 (N_8375,N_4548,N_3117);
nand U8376 (N_8376,N_3218,N_5655);
or U8377 (N_8377,N_3151,N_3236);
or U8378 (N_8378,N_5251,N_5675);
and U8379 (N_8379,N_4225,N_3095);
nor U8380 (N_8380,N_5418,N_3844);
nor U8381 (N_8381,N_5427,N_4131);
and U8382 (N_8382,N_4093,N_3520);
and U8383 (N_8383,N_5208,N_4154);
and U8384 (N_8384,N_5533,N_5674);
nand U8385 (N_8385,N_4105,N_4407);
or U8386 (N_8386,N_5387,N_3495);
and U8387 (N_8387,N_5228,N_5549);
and U8388 (N_8388,N_5565,N_3780);
nand U8389 (N_8389,N_5844,N_3658);
nand U8390 (N_8390,N_4411,N_5749);
xnor U8391 (N_8391,N_4067,N_4646);
nand U8392 (N_8392,N_4673,N_5025);
and U8393 (N_8393,N_3481,N_5476);
or U8394 (N_8394,N_3382,N_4375);
xor U8395 (N_8395,N_5065,N_3438);
and U8396 (N_8396,N_3012,N_5864);
and U8397 (N_8397,N_5674,N_3100);
nor U8398 (N_8398,N_3227,N_4216);
or U8399 (N_8399,N_3269,N_4461);
nor U8400 (N_8400,N_4315,N_5498);
nand U8401 (N_8401,N_4386,N_5993);
or U8402 (N_8402,N_3125,N_4922);
nand U8403 (N_8403,N_3537,N_4047);
or U8404 (N_8404,N_4615,N_3349);
nand U8405 (N_8405,N_3377,N_5488);
nand U8406 (N_8406,N_3774,N_5062);
nor U8407 (N_8407,N_5136,N_3069);
and U8408 (N_8408,N_3723,N_3611);
nor U8409 (N_8409,N_3591,N_4947);
nand U8410 (N_8410,N_5639,N_3377);
nor U8411 (N_8411,N_3881,N_5086);
or U8412 (N_8412,N_5430,N_5759);
and U8413 (N_8413,N_5550,N_4603);
or U8414 (N_8414,N_5705,N_4070);
nand U8415 (N_8415,N_4390,N_5766);
or U8416 (N_8416,N_5784,N_4187);
nand U8417 (N_8417,N_4350,N_3009);
or U8418 (N_8418,N_4114,N_4514);
nand U8419 (N_8419,N_4279,N_4574);
and U8420 (N_8420,N_4141,N_4408);
or U8421 (N_8421,N_4519,N_4788);
and U8422 (N_8422,N_5150,N_5338);
nor U8423 (N_8423,N_4674,N_5524);
or U8424 (N_8424,N_3541,N_3816);
or U8425 (N_8425,N_4629,N_4566);
nor U8426 (N_8426,N_3213,N_3789);
or U8427 (N_8427,N_4724,N_5788);
nor U8428 (N_8428,N_3099,N_4422);
nand U8429 (N_8429,N_3624,N_3967);
nand U8430 (N_8430,N_4304,N_5005);
or U8431 (N_8431,N_4509,N_5683);
and U8432 (N_8432,N_4113,N_4117);
nor U8433 (N_8433,N_3732,N_5218);
and U8434 (N_8434,N_4124,N_3291);
and U8435 (N_8435,N_3077,N_3118);
or U8436 (N_8436,N_4411,N_4058);
nand U8437 (N_8437,N_3529,N_5595);
nor U8438 (N_8438,N_5446,N_4869);
or U8439 (N_8439,N_3629,N_3436);
and U8440 (N_8440,N_3566,N_4177);
and U8441 (N_8441,N_4476,N_4337);
nor U8442 (N_8442,N_3842,N_4882);
nor U8443 (N_8443,N_5368,N_5390);
or U8444 (N_8444,N_3113,N_5545);
nor U8445 (N_8445,N_5169,N_3164);
nand U8446 (N_8446,N_5086,N_3527);
and U8447 (N_8447,N_4950,N_5043);
nand U8448 (N_8448,N_4348,N_3090);
nor U8449 (N_8449,N_5699,N_3144);
nand U8450 (N_8450,N_3098,N_3200);
nor U8451 (N_8451,N_4780,N_5065);
and U8452 (N_8452,N_3289,N_3404);
or U8453 (N_8453,N_4775,N_3864);
nand U8454 (N_8454,N_3969,N_4157);
nand U8455 (N_8455,N_4490,N_4028);
nor U8456 (N_8456,N_4720,N_4795);
or U8457 (N_8457,N_5782,N_3748);
nor U8458 (N_8458,N_3360,N_3860);
and U8459 (N_8459,N_3175,N_3452);
or U8460 (N_8460,N_3178,N_5477);
or U8461 (N_8461,N_4013,N_4532);
and U8462 (N_8462,N_4456,N_4334);
or U8463 (N_8463,N_5825,N_5904);
nand U8464 (N_8464,N_5221,N_3950);
or U8465 (N_8465,N_4907,N_3799);
nor U8466 (N_8466,N_3283,N_4187);
nor U8467 (N_8467,N_3708,N_4364);
or U8468 (N_8468,N_5054,N_5418);
and U8469 (N_8469,N_4243,N_4583);
and U8470 (N_8470,N_3988,N_5224);
or U8471 (N_8471,N_5180,N_5794);
or U8472 (N_8472,N_3058,N_3563);
or U8473 (N_8473,N_5775,N_5466);
nand U8474 (N_8474,N_4653,N_4948);
or U8475 (N_8475,N_5940,N_3259);
and U8476 (N_8476,N_3636,N_5596);
and U8477 (N_8477,N_4675,N_5745);
and U8478 (N_8478,N_3549,N_4586);
nand U8479 (N_8479,N_5597,N_5332);
or U8480 (N_8480,N_4984,N_3911);
and U8481 (N_8481,N_5008,N_4731);
and U8482 (N_8482,N_5932,N_4929);
nor U8483 (N_8483,N_5540,N_4275);
or U8484 (N_8484,N_4688,N_4478);
and U8485 (N_8485,N_3835,N_3840);
nand U8486 (N_8486,N_3526,N_4997);
nand U8487 (N_8487,N_3894,N_3178);
or U8488 (N_8488,N_5256,N_4913);
or U8489 (N_8489,N_5305,N_3501);
or U8490 (N_8490,N_4057,N_4616);
nand U8491 (N_8491,N_5121,N_4594);
nor U8492 (N_8492,N_4086,N_5389);
or U8493 (N_8493,N_4873,N_4012);
or U8494 (N_8494,N_3657,N_4059);
nor U8495 (N_8495,N_5339,N_5217);
nand U8496 (N_8496,N_4281,N_4977);
and U8497 (N_8497,N_4124,N_4332);
nand U8498 (N_8498,N_3594,N_3761);
nand U8499 (N_8499,N_5528,N_4496);
or U8500 (N_8500,N_4703,N_5159);
or U8501 (N_8501,N_4808,N_3996);
or U8502 (N_8502,N_3794,N_3433);
and U8503 (N_8503,N_4370,N_3330);
nand U8504 (N_8504,N_5339,N_5525);
xor U8505 (N_8505,N_4685,N_4698);
nor U8506 (N_8506,N_3425,N_5491);
nand U8507 (N_8507,N_4526,N_3878);
and U8508 (N_8508,N_3026,N_3691);
nor U8509 (N_8509,N_3656,N_3172);
and U8510 (N_8510,N_3479,N_3084);
nor U8511 (N_8511,N_5854,N_4397);
or U8512 (N_8512,N_5354,N_5625);
or U8513 (N_8513,N_5987,N_3126);
and U8514 (N_8514,N_5402,N_5463);
xor U8515 (N_8515,N_4977,N_4430);
nand U8516 (N_8516,N_4917,N_3928);
xor U8517 (N_8517,N_4426,N_5129);
or U8518 (N_8518,N_5219,N_3465);
and U8519 (N_8519,N_3249,N_4232);
nand U8520 (N_8520,N_5156,N_4176);
nand U8521 (N_8521,N_3097,N_5588);
nand U8522 (N_8522,N_3227,N_3110);
nor U8523 (N_8523,N_5223,N_3428);
or U8524 (N_8524,N_5456,N_3232);
or U8525 (N_8525,N_4347,N_5927);
and U8526 (N_8526,N_5644,N_4340);
or U8527 (N_8527,N_4122,N_5327);
xor U8528 (N_8528,N_5818,N_5469);
and U8529 (N_8529,N_5958,N_4259);
and U8530 (N_8530,N_4926,N_3270);
or U8531 (N_8531,N_3827,N_4297);
nor U8532 (N_8532,N_4527,N_4684);
or U8533 (N_8533,N_3091,N_3906);
or U8534 (N_8534,N_5341,N_5235);
nor U8535 (N_8535,N_3881,N_3331);
nand U8536 (N_8536,N_5566,N_5072);
nand U8537 (N_8537,N_4963,N_4373);
nand U8538 (N_8538,N_5127,N_5309);
and U8539 (N_8539,N_3070,N_4860);
nand U8540 (N_8540,N_3154,N_3947);
or U8541 (N_8541,N_3868,N_4327);
nor U8542 (N_8542,N_3653,N_5637);
nor U8543 (N_8543,N_4297,N_5699);
and U8544 (N_8544,N_4527,N_5290);
and U8545 (N_8545,N_4427,N_4367);
nor U8546 (N_8546,N_5452,N_5278);
and U8547 (N_8547,N_5463,N_3690);
or U8548 (N_8548,N_4442,N_5409);
and U8549 (N_8549,N_5206,N_3172);
nand U8550 (N_8550,N_5045,N_3105);
nor U8551 (N_8551,N_5656,N_3678);
nand U8552 (N_8552,N_3831,N_3232);
or U8553 (N_8553,N_4836,N_4671);
nand U8554 (N_8554,N_4554,N_3315);
nand U8555 (N_8555,N_5102,N_4957);
or U8556 (N_8556,N_3865,N_5825);
and U8557 (N_8557,N_3287,N_5244);
nand U8558 (N_8558,N_4904,N_5887);
or U8559 (N_8559,N_4568,N_5810);
nor U8560 (N_8560,N_4120,N_3929);
nor U8561 (N_8561,N_5418,N_5101);
nor U8562 (N_8562,N_5448,N_3002);
nand U8563 (N_8563,N_3441,N_4071);
or U8564 (N_8564,N_5925,N_5542);
and U8565 (N_8565,N_4102,N_4210);
or U8566 (N_8566,N_4569,N_4552);
and U8567 (N_8567,N_5883,N_4033);
or U8568 (N_8568,N_5392,N_4189);
nor U8569 (N_8569,N_4910,N_5265);
and U8570 (N_8570,N_4982,N_3752);
and U8571 (N_8571,N_5394,N_5009);
nand U8572 (N_8572,N_4956,N_4982);
nand U8573 (N_8573,N_4884,N_4608);
nand U8574 (N_8574,N_4450,N_5975);
nor U8575 (N_8575,N_3689,N_4199);
nor U8576 (N_8576,N_5611,N_3958);
nor U8577 (N_8577,N_4228,N_3115);
or U8578 (N_8578,N_5438,N_4432);
or U8579 (N_8579,N_5445,N_5577);
and U8580 (N_8580,N_3741,N_4276);
and U8581 (N_8581,N_5834,N_3413);
and U8582 (N_8582,N_3456,N_4242);
and U8583 (N_8583,N_4385,N_3087);
and U8584 (N_8584,N_4132,N_4068);
or U8585 (N_8585,N_5030,N_4580);
or U8586 (N_8586,N_4209,N_3519);
and U8587 (N_8587,N_3222,N_4326);
or U8588 (N_8588,N_3871,N_5972);
xor U8589 (N_8589,N_4678,N_4138);
and U8590 (N_8590,N_4268,N_3810);
nor U8591 (N_8591,N_3977,N_3533);
nor U8592 (N_8592,N_5726,N_5908);
nand U8593 (N_8593,N_5739,N_4545);
nor U8594 (N_8594,N_3514,N_3154);
and U8595 (N_8595,N_4672,N_5619);
nand U8596 (N_8596,N_4913,N_3853);
nor U8597 (N_8597,N_5919,N_5360);
nor U8598 (N_8598,N_3851,N_4379);
nand U8599 (N_8599,N_5968,N_4141);
nor U8600 (N_8600,N_3090,N_5013);
nand U8601 (N_8601,N_4700,N_4110);
or U8602 (N_8602,N_5539,N_5290);
or U8603 (N_8603,N_3280,N_5619);
and U8604 (N_8604,N_5594,N_5307);
or U8605 (N_8605,N_4494,N_5565);
nor U8606 (N_8606,N_4660,N_5631);
or U8607 (N_8607,N_3521,N_4278);
nand U8608 (N_8608,N_4368,N_3439);
and U8609 (N_8609,N_4276,N_3107);
nand U8610 (N_8610,N_3757,N_4407);
nand U8611 (N_8611,N_4519,N_3791);
or U8612 (N_8612,N_3795,N_3063);
or U8613 (N_8613,N_5797,N_5465);
nor U8614 (N_8614,N_4775,N_4437);
or U8615 (N_8615,N_5498,N_4503);
or U8616 (N_8616,N_3990,N_4372);
nand U8617 (N_8617,N_5824,N_5904);
or U8618 (N_8618,N_3412,N_3131);
and U8619 (N_8619,N_5307,N_3185);
nand U8620 (N_8620,N_3171,N_3464);
nor U8621 (N_8621,N_4543,N_4382);
or U8622 (N_8622,N_5139,N_3521);
or U8623 (N_8623,N_4048,N_4531);
and U8624 (N_8624,N_3873,N_4505);
or U8625 (N_8625,N_4970,N_5010);
nand U8626 (N_8626,N_5845,N_5564);
nor U8627 (N_8627,N_3855,N_3626);
and U8628 (N_8628,N_5799,N_4932);
nor U8629 (N_8629,N_4772,N_4282);
nand U8630 (N_8630,N_3393,N_3704);
and U8631 (N_8631,N_4112,N_4684);
nor U8632 (N_8632,N_3250,N_3164);
nand U8633 (N_8633,N_4585,N_5477);
nor U8634 (N_8634,N_3520,N_4984);
nand U8635 (N_8635,N_4107,N_5573);
nor U8636 (N_8636,N_3162,N_3501);
nand U8637 (N_8637,N_5252,N_4103);
nand U8638 (N_8638,N_3981,N_3765);
nor U8639 (N_8639,N_5577,N_3023);
and U8640 (N_8640,N_3150,N_3233);
nor U8641 (N_8641,N_5901,N_5386);
and U8642 (N_8642,N_3748,N_3552);
nand U8643 (N_8643,N_5361,N_5806);
and U8644 (N_8644,N_3647,N_4902);
or U8645 (N_8645,N_5298,N_4241);
and U8646 (N_8646,N_4139,N_4012);
nand U8647 (N_8647,N_4331,N_3081);
nand U8648 (N_8648,N_3482,N_5320);
and U8649 (N_8649,N_3777,N_5105);
nor U8650 (N_8650,N_4278,N_3319);
and U8651 (N_8651,N_5435,N_4808);
nand U8652 (N_8652,N_5288,N_5384);
and U8653 (N_8653,N_4515,N_5604);
nand U8654 (N_8654,N_3811,N_5844);
nor U8655 (N_8655,N_3189,N_4182);
and U8656 (N_8656,N_4033,N_5945);
or U8657 (N_8657,N_4430,N_5892);
or U8658 (N_8658,N_5270,N_3448);
nor U8659 (N_8659,N_3683,N_3711);
or U8660 (N_8660,N_5609,N_4248);
nand U8661 (N_8661,N_4822,N_4159);
xor U8662 (N_8662,N_5972,N_3268);
nand U8663 (N_8663,N_3588,N_5871);
xor U8664 (N_8664,N_3102,N_4761);
or U8665 (N_8665,N_5193,N_5781);
nand U8666 (N_8666,N_3926,N_5709);
and U8667 (N_8667,N_3153,N_3312);
nor U8668 (N_8668,N_4700,N_4620);
or U8669 (N_8669,N_4638,N_5424);
or U8670 (N_8670,N_4077,N_4099);
nor U8671 (N_8671,N_5351,N_5310);
nand U8672 (N_8672,N_4551,N_3065);
or U8673 (N_8673,N_3808,N_3691);
nand U8674 (N_8674,N_4498,N_5582);
nor U8675 (N_8675,N_3157,N_4801);
nor U8676 (N_8676,N_5235,N_3716);
nand U8677 (N_8677,N_3957,N_4609);
nor U8678 (N_8678,N_4322,N_5728);
and U8679 (N_8679,N_4112,N_3832);
nand U8680 (N_8680,N_4320,N_5348);
nand U8681 (N_8681,N_5568,N_4058);
nor U8682 (N_8682,N_5114,N_5346);
nand U8683 (N_8683,N_3025,N_3189);
and U8684 (N_8684,N_3802,N_3316);
nor U8685 (N_8685,N_4996,N_5368);
or U8686 (N_8686,N_4605,N_3500);
xor U8687 (N_8687,N_3612,N_5844);
or U8688 (N_8688,N_5550,N_4458);
nand U8689 (N_8689,N_4443,N_5743);
or U8690 (N_8690,N_5397,N_5822);
nand U8691 (N_8691,N_5135,N_4083);
and U8692 (N_8692,N_5754,N_5711);
nand U8693 (N_8693,N_4778,N_3231);
and U8694 (N_8694,N_4407,N_5139);
and U8695 (N_8695,N_3318,N_3537);
nand U8696 (N_8696,N_5723,N_3583);
nor U8697 (N_8697,N_5826,N_5928);
nor U8698 (N_8698,N_5435,N_5104);
or U8699 (N_8699,N_4846,N_5173);
nor U8700 (N_8700,N_4725,N_5794);
nand U8701 (N_8701,N_5023,N_3580);
and U8702 (N_8702,N_5780,N_4119);
nor U8703 (N_8703,N_5512,N_3969);
or U8704 (N_8704,N_3567,N_5078);
and U8705 (N_8705,N_4193,N_4442);
and U8706 (N_8706,N_3951,N_3032);
and U8707 (N_8707,N_3623,N_5441);
nand U8708 (N_8708,N_3649,N_5422);
or U8709 (N_8709,N_3058,N_5183);
nand U8710 (N_8710,N_5410,N_3637);
and U8711 (N_8711,N_3423,N_3021);
and U8712 (N_8712,N_4342,N_4979);
nand U8713 (N_8713,N_5380,N_4696);
nand U8714 (N_8714,N_4321,N_3844);
or U8715 (N_8715,N_3883,N_5404);
nor U8716 (N_8716,N_5567,N_4561);
or U8717 (N_8717,N_4803,N_5472);
xnor U8718 (N_8718,N_3237,N_4910);
nor U8719 (N_8719,N_4708,N_3406);
and U8720 (N_8720,N_5320,N_5302);
and U8721 (N_8721,N_3645,N_4310);
and U8722 (N_8722,N_5510,N_5698);
nor U8723 (N_8723,N_5893,N_3808);
nor U8724 (N_8724,N_3693,N_5779);
or U8725 (N_8725,N_3241,N_3736);
nand U8726 (N_8726,N_4574,N_3817);
nor U8727 (N_8727,N_3779,N_5292);
or U8728 (N_8728,N_5847,N_3781);
or U8729 (N_8729,N_4739,N_4475);
nand U8730 (N_8730,N_3285,N_4994);
or U8731 (N_8731,N_5915,N_3256);
and U8732 (N_8732,N_4628,N_3677);
or U8733 (N_8733,N_3479,N_5009);
and U8734 (N_8734,N_3448,N_5132);
nand U8735 (N_8735,N_4129,N_5246);
nand U8736 (N_8736,N_3012,N_4837);
and U8737 (N_8737,N_4999,N_4315);
or U8738 (N_8738,N_3149,N_3774);
nor U8739 (N_8739,N_5941,N_4432);
or U8740 (N_8740,N_4786,N_3336);
nand U8741 (N_8741,N_5982,N_4486);
nor U8742 (N_8742,N_4724,N_3698);
nand U8743 (N_8743,N_5513,N_3607);
nand U8744 (N_8744,N_4539,N_3984);
or U8745 (N_8745,N_3917,N_3203);
or U8746 (N_8746,N_5933,N_4519);
or U8747 (N_8747,N_5812,N_5717);
nand U8748 (N_8748,N_5750,N_3429);
nand U8749 (N_8749,N_3970,N_5661);
and U8750 (N_8750,N_5582,N_4063);
nand U8751 (N_8751,N_5457,N_3711);
or U8752 (N_8752,N_3388,N_3367);
and U8753 (N_8753,N_4124,N_3360);
and U8754 (N_8754,N_5097,N_4609);
nand U8755 (N_8755,N_4178,N_3383);
xor U8756 (N_8756,N_5463,N_3202);
nand U8757 (N_8757,N_5863,N_4861);
and U8758 (N_8758,N_3646,N_5265);
and U8759 (N_8759,N_4469,N_3712);
nand U8760 (N_8760,N_3408,N_4846);
nand U8761 (N_8761,N_4664,N_3410);
nor U8762 (N_8762,N_5924,N_5969);
nor U8763 (N_8763,N_5698,N_5125);
or U8764 (N_8764,N_3767,N_4417);
and U8765 (N_8765,N_5885,N_3895);
nor U8766 (N_8766,N_3767,N_4869);
or U8767 (N_8767,N_3404,N_3435);
nand U8768 (N_8768,N_3339,N_4189);
and U8769 (N_8769,N_5902,N_3580);
nor U8770 (N_8770,N_4714,N_3833);
nand U8771 (N_8771,N_5575,N_3771);
nand U8772 (N_8772,N_5522,N_3684);
nand U8773 (N_8773,N_5095,N_5807);
or U8774 (N_8774,N_4176,N_5848);
nor U8775 (N_8775,N_4373,N_4478);
or U8776 (N_8776,N_4096,N_4613);
or U8777 (N_8777,N_5267,N_3668);
nor U8778 (N_8778,N_4425,N_3499);
nor U8779 (N_8779,N_4653,N_4544);
nand U8780 (N_8780,N_5277,N_5071);
nor U8781 (N_8781,N_5143,N_5478);
nand U8782 (N_8782,N_5820,N_5748);
nand U8783 (N_8783,N_5131,N_5564);
and U8784 (N_8784,N_5488,N_4536);
nand U8785 (N_8785,N_5236,N_3168);
and U8786 (N_8786,N_3130,N_4120);
nor U8787 (N_8787,N_3801,N_4202);
and U8788 (N_8788,N_3351,N_4822);
nor U8789 (N_8789,N_5828,N_5203);
or U8790 (N_8790,N_5759,N_5644);
and U8791 (N_8791,N_4689,N_5818);
and U8792 (N_8792,N_5020,N_5357);
or U8793 (N_8793,N_3097,N_4470);
xnor U8794 (N_8794,N_5038,N_5290);
xor U8795 (N_8795,N_3428,N_3532);
nand U8796 (N_8796,N_5937,N_5797);
and U8797 (N_8797,N_5021,N_3779);
or U8798 (N_8798,N_3343,N_5925);
nor U8799 (N_8799,N_3283,N_3188);
and U8800 (N_8800,N_3074,N_5054);
nor U8801 (N_8801,N_5761,N_3453);
and U8802 (N_8802,N_3653,N_3560);
nor U8803 (N_8803,N_5403,N_3631);
and U8804 (N_8804,N_5927,N_5935);
and U8805 (N_8805,N_5581,N_3334);
or U8806 (N_8806,N_5815,N_3318);
and U8807 (N_8807,N_5673,N_5949);
or U8808 (N_8808,N_3412,N_5240);
nand U8809 (N_8809,N_4740,N_5062);
and U8810 (N_8810,N_3006,N_5082);
and U8811 (N_8811,N_3271,N_4910);
or U8812 (N_8812,N_3803,N_4676);
nand U8813 (N_8813,N_3606,N_5209);
nor U8814 (N_8814,N_5681,N_4984);
xor U8815 (N_8815,N_4142,N_5982);
nand U8816 (N_8816,N_5033,N_4221);
and U8817 (N_8817,N_5421,N_4021);
and U8818 (N_8818,N_5585,N_4311);
and U8819 (N_8819,N_4651,N_4785);
or U8820 (N_8820,N_4532,N_4351);
nor U8821 (N_8821,N_4863,N_4988);
or U8822 (N_8822,N_3091,N_4029);
and U8823 (N_8823,N_4886,N_4824);
nor U8824 (N_8824,N_5698,N_4809);
nand U8825 (N_8825,N_5806,N_3724);
nor U8826 (N_8826,N_4458,N_5599);
and U8827 (N_8827,N_3799,N_5079);
nand U8828 (N_8828,N_4772,N_4399);
xor U8829 (N_8829,N_3551,N_4701);
or U8830 (N_8830,N_4594,N_5270);
nand U8831 (N_8831,N_4253,N_5343);
nor U8832 (N_8832,N_5335,N_3138);
xnor U8833 (N_8833,N_3056,N_3566);
and U8834 (N_8834,N_5891,N_5002);
nor U8835 (N_8835,N_4370,N_4034);
or U8836 (N_8836,N_3983,N_3090);
or U8837 (N_8837,N_5222,N_5712);
or U8838 (N_8838,N_5340,N_4093);
and U8839 (N_8839,N_3293,N_5633);
nor U8840 (N_8840,N_4576,N_3132);
nand U8841 (N_8841,N_4388,N_5186);
and U8842 (N_8842,N_3961,N_4422);
nand U8843 (N_8843,N_3009,N_4952);
and U8844 (N_8844,N_5750,N_3227);
and U8845 (N_8845,N_4358,N_5231);
nor U8846 (N_8846,N_4282,N_3231);
or U8847 (N_8847,N_4031,N_5424);
and U8848 (N_8848,N_3657,N_4885);
or U8849 (N_8849,N_5479,N_3710);
and U8850 (N_8850,N_4349,N_3752);
nor U8851 (N_8851,N_4444,N_5233);
nor U8852 (N_8852,N_3375,N_5937);
or U8853 (N_8853,N_5212,N_4617);
nand U8854 (N_8854,N_3929,N_3330);
nor U8855 (N_8855,N_5216,N_4725);
nor U8856 (N_8856,N_4427,N_4202);
nand U8857 (N_8857,N_3246,N_5255);
and U8858 (N_8858,N_5238,N_5766);
nor U8859 (N_8859,N_3965,N_4592);
and U8860 (N_8860,N_4998,N_4046);
or U8861 (N_8861,N_4814,N_4435);
nor U8862 (N_8862,N_4018,N_5436);
or U8863 (N_8863,N_4747,N_5528);
and U8864 (N_8864,N_4875,N_4171);
and U8865 (N_8865,N_3045,N_3497);
or U8866 (N_8866,N_5866,N_3981);
and U8867 (N_8867,N_5328,N_3523);
and U8868 (N_8868,N_5631,N_5755);
and U8869 (N_8869,N_4133,N_3850);
or U8870 (N_8870,N_5227,N_5675);
or U8871 (N_8871,N_4239,N_5220);
and U8872 (N_8872,N_5520,N_3477);
nor U8873 (N_8873,N_4154,N_5196);
nand U8874 (N_8874,N_4179,N_5782);
and U8875 (N_8875,N_4625,N_3926);
nor U8876 (N_8876,N_5058,N_4279);
nand U8877 (N_8877,N_4324,N_5677);
or U8878 (N_8878,N_4293,N_3569);
nand U8879 (N_8879,N_5649,N_3069);
nor U8880 (N_8880,N_3406,N_4126);
nor U8881 (N_8881,N_4595,N_3427);
or U8882 (N_8882,N_3771,N_5009);
and U8883 (N_8883,N_4234,N_4895);
nand U8884 (N_8884,N_5375,N_5717);
nor U8885 (N_8885,N_4412,N_4212);
and U8886 (N_8886,N_5852,N_4645);
nand U8887 (N_8887,N_4074,N_4260);
or U8888 (N_8888,N_5613,N_4998);
and U8889 (N_8889,N_3691,N_5502);
or U8890 (N_8890,N_4613,N_3208);
nand U8891 (N_8891,N_3261,N_4107);
or U8892 (N_8892,N_3109,N_4403);
nor U8893 (N_8893,N_4476,N_4227);
or U8894 (N_8894,N_4273,N_5703);
or U8895 (N_8895,N_4575,N_5711);
or U8896 (N_8896,N_5212,N_4414);
nor U8897 (N_8897,N_3629,N_4052);
nor U8898 (N_8898,N_4911,N_4448);
nor U8899 (N_8899,N_4041,N_4902);
or U8900 (N_8900,N_5587,N_5135);
or U8901 (N_8901,N_5377,N_4811);
nand U8902 (N_8902,N_3134,N_3439);
nor U8903 (N_8903,N_4257,N_5926);
and U8904 (N_8904,N_3043,N_3002);
nor U8905 (N_8905,N_3774,N_5250);
and U8906 (N_8906,N_5784,N_3128);
nor U8907 (N_8907,N_5038,N_3006);
nand U8908 (N_8908,N_5325,N_5449);
nor U8909 (N_8909,N_3503,N_5530);
nor U8910 (N_8910,N_4010,N_5231);
and U8911 (N_8911,N_5208,N_5088);
nor U8912 (N_8912,N_5569,N_5778);
and U8913 (N_8913,N_3302,N_4743);
and U8914 (N_8914,N_3024,N_5946);
nor U8915 (N_8915,N_4136,N_5833);
nand U8916 (N_8916,N_4762,N_4486);
nand U8917 (N_8917,N_3757,N_4132);
nand U8918 (N_8918,N_5002,N_3729);
nor U8919 (N_8919,N_4800,N_4210);
and U8920 (N_8920,N_3477,N_3229);
and U8921 (N_8921,N_3576,N_3262);
and U8922 (N_8922,N_3204,N_4499);
and U8923 (N_8923,N_5774,N_5507);
nor U8924 (N_8924,N_5567,N_4031);
or U8925 (N_8925,N_5543,N_4489);
nand U8926 (N_8926,N_3497,N_3553);
nand U8927 (N_8927,N_3281,N_3620);
or U8928 (N_8928,N_3994,N_4397);
nor U8929 (N_8929,N_3114,N_5624);
nor U8930 (N_8930,N_3142,N_3446);
xor U8931 (N_8931,N_4168,N_4050);
nor U8932 (N_8932,N_3944,N_4615);
nand U8933 (N_8933,N_3485,N_4740);
or U8934 (N_8934,N_3849,N_5566);
nor U8935 (N_8935,N_5199,N_4390);
nand U8936 (N_8936,N_5476,N_3475);
and U8937 (N_8937,N_5945,N_5150);
xnor U8938 (N_8938,N_3890,N_4063);
nand U8939 (N_8939,N_4667,N_5240);
or U8940 (N_8940,N_5950,N_4077);
or U8941 (N_8941,N_4843,N_4832);
xnor U8942 (N_8942,N_5466,N_4704);
and U8943 (N_8943,N_5787,N_3040);
nand U8944 (N_8944,N_3704,N_3750);
or U8945 (N_8945,N_4698,N_3664);
and U8946 (N_8946,N_5612,N_3344);
or U8947 (N_8947,N_4885,N_5401);
or U8948 (N_8948,N_5392,N_5817);
and U8949 (N_8949,N_4918,N_5670);
nand U8950 (N_8950,N_4340,N_5920);
nor U8951 (N_8951,N_3530,N_5351);
nor U8952 (N_8952,N_5790,N_3315);
and U8953 (N_8953,N_3861,N_4107);
and U8954 (N_8954,N_3264,N_4636);
nand U8955 (N_8955,N_5408,N_3327);
nor U8956 (N_8956,N_5763,N_3976);
nor U8957 (N_8957,N_4796,N_5562);
and U8958 (N_8958,N_3010,N_5571);
nor U8959 (N_8959,N_3651,N_4152);
or U8960 (N_8960,N_4659,N_5706);
nand U8961 (N_8961,N_5542,N_4135);
and U8962 (N_8962,N_5659,N_5925);
or U8963 (N_8963,N_4202,N_5270);
nor U8964 (N_8964,N_5799,N_4035);
and U8965 (N_8965,N_5529,N_5383);
nor U8966 (N_8966,N_5498,N_5591);
and U8967 (N_8967,N_4737,N_5374);
nor U8968 (N_8968,N_5675,N_3673);
nand U8969 (N_8969,N_5260,N_5983);
nor U8970 (N_8970,N_4056,N_5060);
and U8971 (N_8971,N_4359,N_3955);
nor U8972 (N_8972,N_5503,N_4103);
and U8973 (N_8973,N_4022,N_3631);
or U8974 (N_8974,N_3764,N_4642);
nor U8975 (N_8975,N_4474,N_5447);
nor U8976 (N_8976,N_3009,N_4493);
and U8977 (N_8977,N_3353,N_4684);
or U8978 (N_8978,N_4470,N_3959);
nor U8979 (N_8979,N_3144,N_3979);
or U8980 (N_8980,N_5988,N_4881);
or U8981 (N_8981,N_3254,N_4036);
nand U8982 (N_8982,N_4846,N_3089);
and U8983 (N_8983,N_3624,N_5294);
or U8984 (N_8984,N_5909,N_4283);
and U8985 (N_8985,N_5845,N_5036);
nor U8986 (N_8986,N_5933,N_4520);
nand U8987 (N_8987,N_4547,N_4222);
nor U8988 (N_8988,N_4162,N_3812);
nor U8989 (N_8989,N_3885,N_4570);
and U8990 (N_8990,N_3215,N_5502);
nand U8991 (N_8991,N_5545,N_3049);
and U8992 (N_8992,N_3192,N_3890);
or U8993 (N_8993,N_5246,N_4428);
nor U8994 (N_8994,N_3456,N_4127);
nand U8995 (N_8995,N_4927,N_5730);
nand U8996 (N_8996,N_5940,N_3159);
xor U8997 (N_8997,N_5301,N_5623);
nand U8998 (N_8998,N_3771,N_4362);
nor U8999 (N_8999,N_4501,N_4529);
xnor U9000 (N_9000,N_6712,N_7333);
or U9001 (N_9001,N_7266,N_7024);
or U9002 (N_9002,N_8022,N_7530);
nor U9003 (N_9003,N_7281,N_8011);
or U9004 (N_9004,N_8860,N_8788);
nand U9005 (N_9005,N_7257,N_8965);
or U9006 (N_9006,N_6899,N_7450);
nor U9007 (N_9007,N_6403,N_8659);
and U9008 (N_9008,N_6308,N_7105);
and U9009 (N_9009,N_8255,N_7693);
nand U9010 (N_9010,N_8419,N_7354);
and U9011 (N_9011,N_8998,N_6323);
or U9012 (N_9012,N_7498,N_8677);
nor U9013 (N_9013,N_6816,N_6410);
nand U9014 (N_9014,N_6602,N_6087);
and U9015 (N_9015,N_6979,N_8603);
or U9016 (N_9016,N_8383,N_8322);
or U9017 (N_9017,N_8171,N_6779);
xnor U9018 (N_9018,N_6359,N_8729);
and U9019 (N_9019,N_6691,N_6495);
nor U9020 (N_9020,N_8735,N_7873);
nand U9021 (N_9021,N_8911,N_6548);
or U9022 (N_9022,N_6862,N_6438);
and U9023 (N_9023,N_8177,N_8543);
and U9024 (N_9024,N_7004,N_6633);
and U9025 (N_9025,N_7397,N_6027);
and U9026 (N_9026,N_6915,N_7437);
and U9027 (N_9027,N_6958,N_6268);
nand U9028 (N_9028,N_8232,N_6757);
nand U9029 (N_9029,N_8651,N_6888);
nand U9030 (N_9030,N_7468,N_7310);
and U9031 (N_9031,N_6156,N_8639);
or U9032 (N_9032,N_6075,N_7378);
nand U9033 (N_9033,N_7395,N_6569);
nand U9034 (N_9034,N_7211,N_6695);
nand U9035 (N_9035,N_7252,N_7444);
nand U9036 (N_9036,N_6292,N_6188);
or U9037 (N_9037,N_8721,N_7718);
and U9038 (N_9038,N_7603,N_6611);
nand U9039 (N_9039,N_7454,N_8319);
nand U9040 (N_9040,N_7825,N_8823);
or U9041 (N_9041,N_7910,N_7001);
or U9042 (N_9042,N_8618,N_8036);
nand U9043 (N_9043,N_6190,N_7569);
nand U9044 (N_9044,N_6989,N_8400);
nor U9045 (N_9045,N_7883,N_8790);
or U9046 (N_9046,N_8738,N_8945);
nor U9047 (N_9047,N_7092,N_6825);
nand U9048 (N_9048,N_6728,N_7697);
nor U9049 (N_9049,N_7962,N_8754);
nand U9050 (N_9050,N_7694,N_7106);
and U9051 (N_9051,N_8562,N_8575);
nor U9052 (N_9052,N_6701,N_6982);
nand U9053 (N_9053,N_7533,N_8699);
or U9054 (N_9054,N_6697,N_6251);
and U9055 (N_9055,N_6226,N_6029);
and U9056 (N_9056,N_7710,N_7654);
or U9057 (N_9057,N_6497,N_8500);
nor U9058 (N_9058,N_8139,N_7089);
or U9059 (N_9059,N_8850,N_7937);
and U9060 (N_9060,N_8637,N_8154);
nand U9061 (N_9061,N_6956,N_7897);
or U9062 (N_9062,N_8898,N_7506);
nand U9063 (N_9063,N_7088,N_8986);
or U9064 (N_9064,N_7431,N_8170);
and U9065 (N_9065,N_8100,N_7941);
nor U9066 (N_9066,N_8143,N_6318);
and U9067 (N_9067,N_8789,N_8498);
or U9068 (N_9068,N_7278,N_8877);
nand U9069 (N_9069,N_6651,N_6022);
nand U9070 (N_9070,N_8441,N_7866);
nor U9071 (N_9071,N_8774,N_8309);
nand U9072 (N_9072,N_6386,N_6930);
nand U9073 (N_9073,N_8270,N_7615);
nand U9074 (N_9074,N_6872,N_8303);
nand U9075 (N_9075,N_6142,N_6686);
nand U9076 (N_9076,N_7069,N_6132);
and U9077 (N_9077,N_6504,N_6940);
nor U9078 (N_9078,N_6452,N_6471);
nand U9079 (N_9079,N_7125,N_6809);
nor U9080 (N_9080,N_6833,N_6258);
or U9081 (N_9081,N_6923,N_8094);
nand U9082 (N_9082,N_7110,N_8041);
or U9083 (N_9083,N_7008,N_6551);
and U9084 (N_9084,N_6484,N_7610);
nor U9085 (N_9085,N_8121,N_8365);
nand U9086 (N_9086,N_6222,N_7302);
or U9087 (N_9087,N_8919,N_6916);
and U9088 (N_9088,N_6131,N_6017);
nor U9089 (N_9089,N_7400,N_8035);
and U9090 (N_9090,N_7308,N_8403);
and U9091 (N_9091,N_6562,N_8669);
nor U9092 (N_9092,N_8028,N_8631);
and U9093 (N_9093,N_7597,N_8452);
nor U9094 (N_9094,N_7413,N_7970);
nor U9095 (N_9095,N_6482,N_7619);
or U9096 (N_9096,N_8222,N_7653);
nand U9097 (N_9097,N_8952,N_7967);
or U9098 (N_9098,N_6453,N_8890);
nand U9099 (N_9099,N_6593,N_6669);
nand U9100 (N_9100,N_7746,N_6086);
nand U9101 (N_9101,N_6882,N_6441);
and U9102 (N_9102,N_6466,N_8101);
and U9103 (N_9103,N_8853,N_6641);
and U9104 (N_9104,N_6741,N_6626);
or U9105 (N_9105,N_8996,N_7396);
or U9106 (N_9106,N_7276,N_8082);
or U9107 (N_9107,N_7629,N_8897);
nand U9108 (N_9108,N_7785,N_6890);
or U9109 (N_9109,N_8787,N_8000);
nor U9110 (N_9110,N_6874,N_7340);
or U9111 (N_9111,N_6970,N_6309);
nand U9112 (N_9112,N_6010,N_7770);
nand U9113 (N_9113,N_6286,N_7129);
and U9114 (N_9114,N_7799,N_8475);
nor U9115 (N_9115,N_8152,N_8535);
or U9116 (N_9116,N_7461,N_8885);
or U9117 (N_9117,N_7227,N_7581);
nand U9118 (N_9118,N_8081,N_7440);
nor U9119 (N_9119,N_7784,N_7856);
and U9120 (N_9120,N_8662,N_7280);
and U9121 (N_9121,N_8807,N_6205);
nand U9122 (N_9122,N_7441,N_7501);
and U9123 (N_9123,N_8524,N_8974);
and U9124 (N_9124,N_8624,N_6181);
and U9125 (N_9125,N_7151,N_7261);
and U9126 (N_9126,N_6578,N_8185);
nand U9127 (N_9127,N_7933,N_6692);
or U9128 (N_9128,N_8769,N_8192);
nand U9129 (N_9129,N_7052,N_7073);
xor U9130 (N_9130,N_6588,N_7368);
or U9131 (N_9131,N_8463,N_8399);
nand U9132 (N_9132,N_6853,N_7868);
or U9133 (N_9133,N_6330,N_7251);
nand U9134 (N_9134,N_7657,N_6366);
nand U9135 (N_9135,N_8156,N_6931);
and U9136 (N_9136,N_6362,N_6854);
and U9137 (N_9137,N_8153,N_6442);
nor U9138 (N_9138,N_6841,N_8380);
and U9139 (N_9139,N_8886,N_6472);
or U9140 (N_9140,N_6408,N_7604);
and U9141 (N_9141,N_7067,N_7234);
and U9142 (N_9142,N_7406,N_6901);
or U9143 (N_9143,N_8375,N_7231);
or U9144 (N_9144,N_7021,N_6861);
nor U9145 (N_9145,N_7594,N_8636);
xor U9146 (N_9146,N_8578,N_7344);
nor U9147 (N_9147,N_6850,N_7741);
or U9148 (N_9148,N_7453,N_7375);
nor U9149 (N_9149,N_8984,N_7828);
or U9150 (N_9150,N_8893,N_7595);
or U9151 (N_9151,N_6015,N_8717);
and U9152 (N_9152,N_6744,N_8931);
nor U9153 (N_9153,N_6341,N_6594);
nand U9154 (N_9154,N_7078,N_7372);
nand U9155 (N_9155,N_7179,N_6476);
xor U9156 (N_9156,N_8961,N_8382);
and U9157 (N_9157,N_6020,N_8751);
and U9158 (N_9158,N_6846,N_7640);
nand U9159 (N_9159,N_8838,N_6467);
nand U9160 (N_9160,N_7051,N_7751);
or U9161 (N_9161,N_6420,N_6404);
nor U9162 (N_9162,N_6334,N_7842);
nand U9163 (N_9163,N_7079,N_8800);
nand U9164 (N_9164,N_6040,N_6939);
nor U9165 (N_9165,N_8756,N_6628);
nor U9166 (N_9166,N_6148,N_8078);
nand U9167 (N_9167,N_6987,N_8001);
and U9168 (N_9168,N_6058,N_8158);
or U9169 (N_9169,N_8155,N_7117);
or U9170 (N_9170,N_6619,N_6450);
and U9171 (N_9171,N_6306,N_7470);
and U9172 (N_9172,N_8835,N_6090);
nor U9173 (N_9173,N_8806,N_8138);
or U9174 (N_9174,N_7643,N_6274);
xnor U9175 (N_9175,N_6567,N_7200);
and U9176 (N_9176,N_7817,N_8874);
nor U9177 (N_9177,N_6380,N_7309);
and U9178 (N_9178,N_8221,N_8727);
and U9179 (N_9179,N_7291,N_8615);
and U9180 (N_9180,N_8709,N_6771);
nand U9181 (N_9181,N_6895,N_7865);
nor U9182 (N_9182,N_6470,N_7509);
nand U9183 (N_9183,N_6212,N_6689);
and U9184 (N_9184,N_6083,N_6097);
and U9185 (N_9185,N_6655,N_6926);
nor U9186 (N_9186,N_7191,N_7293);
and U9187 (N_9187,N_8980,N_7432);
and U9188 (N_9188,N_6179,N_7745);
nand U9189 (N_9189,N_7561,N_8124);
nand U9190 (N_9190,N_7793,N_7656);
nand U9191 (N_9191,N_7322,N_7666);
nand U9192 (N_9192,N_7072,N_8406);
nor U9193 (N_9193,N_8167,N_6517);
nand U9194 (N_9194,N_6117,N_7325);
and U9195 (N_9195,N_8541,N_7859);
nor U9196 (N_9196,N_7153,N_6592);
nor U9197 (N_9197,N_8266,N_8292);
and U9198 (N_9198,N_6737,N_8679);
and U9199 (N_9199,N_7382,N_6049);
nor U9200 (N_9200,N_8157,N_8061);
xor U9201 (N_9201,N_8570,N_8982);
nor U9202 (N_9202,N_7305,N_6917);
or U9203 (N_9203,N_7819,N_7235);
nor U9204 (N_9204,N_7788,N_7102);
nand U9205 (N_9205,N_6963,N_8581);
nand U9206 (N_9206,N_6041,N_8103);
xnor U9207 (N_9207,N_8329,N_8917);
or U9208 (N_9208,N_7459,N_6640);
xor U9209 (N_9209,N_8294,N_7210);
and U9210 (N_9210,N_6394,N_7535);
or U9211 (N_9211,N_6024,N_8630);
nand U9212 (N_9212,N_8083,N_8644);
nor U9213 (N_9213,N_6465,N_7659);
or U9214 (N_9214,N_8687,N_8076);
xnor U9215 (N_9215,N_6234,N_7928);
nor U9216 (N_9216,N_7849,N_8596);
and U9217 (N_9217,N_7848,N_8063);
nand U9218 (N_9218,N_6598,N_8247);
nor U9219 (N_9219,N_6167,N_7734);
nand U9220 (N_9220,N_8533,N_8102);
or U9221 (N_9221,N_6896,N_7850);
nand U9222 (N_9222,N_6540,N_8418);
and U9223 (N_9223,N_7899,N_8527);
or U9224 (N_9224,N_8275,N_6823);
or U9225 (N_9225,N_7513,N_7651);
nor U9226 (N_9226,N_7748,N_8528);
and U9227 (N_9227,N_8310,N_6604);
or U9228 (N_9228,N_8655,N_8796);
nor U9229 (N_9229,N_7776,N_8069);
or U9230 (N_9230,N_7685,N_8490);
or U9231 (N_9231,N_6413,N_6787);
xor U9232 (N_9232,N_6925,N_6373);
nor U9233 (N_9233,N_7399,N_7242);
or U9234 (N_9234,N_6698,N_6337);
nor U9235 (N_9235,N_7735,N_6834);
and U9236 (N_9236,N_8362,N_8750);
nand U9237 (N_9237,N_7076,N_6676);
and U9238 (N_9238,N_7335,N_8914);
and U9239 (N_9239,N_7992,N_6199);
nor U9240 (N_9240,N_8220,N_8424);
and U9241 (N_9241,N_8136,N_8048);
or U9242 (N_9242,N_8391,N_7987);
and U9243 (N_9243,N_6705,N_7913);
nand U9244 (N_9244,N_7930,N_7548);
or U9245 (N_9245,N_8812,N_8600);
or U9246 (N_9246,N_7475,N_7598);
or U9247 (N_9247,N_6770,N_7057);
and U9248 (N_9248,N_8511,N_6550);
nand U9249 (N_9249,N_6262,N_7923);
nor U9250 (N_9250,N_8647,N_7159);
and U9251 (N_9251,N_7605,N_7524);
nor U9252 (N_9252,N_7875,N_6388);
nand U9253 (N_9253,N_8314,N_6125);
and U9254 (N_9254,N_6894,N_6508);
nand U9255 (N_9255,N_6168,N_8161);
and U9256 (N_9256,N_6719,N_8002);
and U9257 (N_9257,N_8127,N_8859);
or U9258 (N_9258,N_7119,N_7912);
nand U9259 (N_9259,N_8110,N_8300);
and U9260 (N_9260,N_7932,N_6510);
nand U9261 (N_9261,N_6563,N_6751);
or U9262 (N_9262,N_6295,N_7763);
or U9263 (N_9263,N_6171,N_8340);
nor U9264 (N_9264,N_7938,N_6233);
xor U9265 (N_9265,N_6101,N_8026);
nor U9266 (N_9266,N_7502,N_8708);
xnor U9267 (N_9267,N_6019,N_8445);
and U9268 (N_9268,N_7846,N_6216);
and U9269 (N_9269,N_6773,N_7542);
or U9270 (N_9270,N_6758,N_6433);
or U9271 (N_9271,N_7661,N_6736);
nor U9272 (N_9272,N_8281,N_7225);
or U9273 (N_9273,N_8967,N_7256);
nor U9274 (N_9274,N_6445,N_6525);
and U9275 (N_9275,N_8009,N_7360);
nor U9276 (N_9276,N_7632,N_7152);
or U9277 (N_9277,N_6514,N_6146);
or U9278 (N_9278,N_6391,N_8684);
nand U9279 (N_9279,N_6228,N_6727);
or U9280 (N_9280,N_7177,N_7262);
nor U9281 (N_9281,N_6990,N_7889);
and U9282 (N_9282,N_7414,N_7445);
nor U9283 (N_9283,N_8461,N_6332);
nand U9284 (N_9284,N_8989,N_7424);
or U9285 (N_9285,N_6129,N_8620);
nor U9286 (N_9286,N_6107,N_6710);
and U9287 (N_9287,N_6724,N_7772);
and U9288 (N_9288,N_7725,N_8010);
and U9289 (N_9289,N_7096,N_7279);
nor U9290 (N_9290,N_7924,N_7165);
nor U9291 (N_9291,N_7044,N_8905);
and U9292 (N_9292,N_8262,N_7046);
or U9293 (N_9293,N_7835,N_6952);
nand U9294 (N_9294,N_7267,N_6050);
nand U9295 (N_9295,N_8964,N_6473);
and U9296 (N_9296,N_7915,N_6449);
or U9297 (N_9297,N_7170,N_8466);
nor U9298 (N_9298,N_8146,N_7155);
nor U9299 (N_9299,N_6532,N_8782);
nand U9300 (N_9300,N_7220,N_6071);
and U9301 (N_9301,N_6672,N_8568);
and U9302 (N_9302,N_7085,N_8480);
and U9303 (N_9303,N_7701,N_6423);
nand U9304 (N_9304,N_8323,N_6650);
nand U9305 (N_9305,N_7197,N_8759);
xor U9306 (N_9306,N_6080,N_6706);
nand U9307 (N_9307,N_6509,N_8887);
nand U9308 (N_9308,N_7587,N_6906);
nand U9309 (N_9309,N_7668,N_6743);
or U9310 (N_9310,N_8326,N_7224);
and U9311 (N_9311,N_7209,N_8748);
or U9312 (N_9312,N_7931,N_7381);
and U9313 (N_9313,N_8566,N_7321);
nand U9314 (N_9314,N_8390,N_8858);
nand U9315 (N_9315,N_8492,N_8333);
or U9316 (N_9316,N_6824,N_8560);
and U9317 (N_9317,N_7936,N_6671);
or U9318 (N_9318,N_6516,N_8515);
nor U9319 (N_9319,N_7295,N_8271);
nand U9320 (N_9320,N_7775,N_6443);
nor U9321 (N_9321,N_7499,N_8957);
nor U9322 (N_9322,N_8920,N_7313);
xnor U9323 (N_9323,N_8357,N_6335);
nand U9324 (N_9324,N_7664,N_6063);
or U9325 (N_9325,N_7645,N_8050);
nand U9326 (N_9326,N_6774,N_7973);
or U9327 (N_9327,N_7390,N_6105);
or U9328 (N_9328,N_8531,N_8546);
nor U9329 (N_9329,N_7346,N_7503);
and U9330 (N_9330,N_6867,N_7149);
and U9331 (N_9331,N_8246,N_8619);
or U9332 (N_9332,N_6369,N_6880);
and U9333 (N_9333,N_6485,N_6791);
and U9334 (N_9334,N_6478,N_6827);
nor U9335 (N_9335,N_7099,N_6848);
and U9336 (N_9336,N_7374,N_8785);
or U9337 (N_9337,N_8707,N_8868);
or U9338 (N_9338,N_6991,N_7221);
and U9339 (N_9339,N_6648,N_6372);
nor U9340 (N_9340,N_7929,N_8387);
nor U9341 (N_9341,N_7827,N_7755);
nand U9342 (N_9342,N_7623,N_7168);
nor U9343 (N_9343,N_8473,N_7794);
nor U9344 (N_9344,N_6828,N_8767);
nand U9345 (N_9345,N_8491,N_8719);
nand U9346 (N_9346,N_7226,N_6822);
nor U9347 (N_9347,N_8203,N_7841);
and U9348 (N_9348,N_6056,N_6618);
or U9349 (N_9349,N_7583,N_6847);
and U9350 (N_9350,N_7202,N_6155);
and U9351 (N_9351,N_6902,N_8829);
or U9352 (N_9352,N_7655,N_7056);
and U9353 (N_9353,N_6252,N_7528);
or U9354 (N_9354,N_8057,N_8373);
nand U9355 (N_9355,N_8554,N_8224);
and U9356 (N_9356,N_8386,N_8163);
or U9357 (N_9357,N_7109,N_6570);
or U9358 (N_9358,N_6191,N_8025);
xnor U9359 (N_9359,N_7000,N_8683);
and U9360 (N_9360,N_6273,N_7030);
and U9361 (N_9361,N_7860,N_7781);
nor U9362 (N_9362,N_6708,N_7438);
and U9363 (N_9363,N_8693,N_6186);
nand U9364 (N_9364,N_6536,N_8297);
nor U9365 (N_9365,N_7917,N_8346);
nor U9366 (N_9366,N_8369,N_6422);
nand U9367 (N_9367,N_6333,N_8066);
xnor U9368 (N_9368,N_6440,N_8062);
nand U9369 (N_9369,N_7166,N_7675);
and U9370 (N_9370,N_6948,N_6585);
nor U9371 (N_9371,N_8027,N_6519);
and U9372 (N_9372,N_8106,N_7779);
nor U9373 (N_9373,N_8488,N_7876);
and U9374 (N_9374,N_6102,N_6277);
or U9375 (N_9375,N_7443,N_7403);
nor U9376 (N_9376,N_7270,N_8431);
nor U9377 (N_9377,N_8927,N_6079);
and U9378 (N_9378,N_6474,N_6907);
nor U9379 (N_9379,N_7804,N_7285);
nor U9380 (N_9380,N_8182,N_7641);
nand U9381 (N_9381,N_6831,N_7916);
or U9382 (N_9382,N_6634,N_7199);
nor U9383 (N_9383,N_7233,N_8432);
and U9384 (N_9384,N_7189,N_6392);
nand U9385 (N_9385,N_7803,N_8287);
nand U9386 (N_9386,N_8839,N_8617);
or U9387 (N_9387,N_6203,N_6196);
nor U9388 (N_9388,N_7306,N_7742);
and U9389 (N_9389,N_7379,N_7562);
nand U9390 (N_9390,N_6808,N_7350);
nor U9391 (N_9391,N_7362,N_8526);
nor U9392 (N_9392,N_8414,N_6756);
or U9393 (N_9393,N_7780,N_8409);
nand U9394 (N_9394,N_8706,N_6638);
nand U9395 (N_9395,N_8962,N_8530);
nand U9396 (N_9396,N_8983,N_8460);
and U9397 (N_9397,N_7521,N_8694);
xor U9398 (N_9398,N_7269,N_8450);
or U9399 (N_9399,N_6621,N_8234);
nor U9400 (N_9400,N_8878,N_8016);
and U9401 (N_9401,N_6430,N_6389);
nand U9402 (N_9402,N_7128,N_8656);
nor U9403 (N_9403,N_8777,N_8194);
nand U9404 (N_9404,N_7728,N_8744);
nand U9405 (N_9405,N_6393,N_8770);
nor U9406 (N_9406,N_8064,N_8206);
nor U9407 (N_9407,N_8781,N_6182);
or U9408 (N_9408,N_7287,N_6266);
and U9409 (N_9409,N_7778,N_6008);
and U9410 (N_9410,N_7223,N_8700);
nor U9411 (N_9411,N_8739,N_8430);
or U9412 (N_9412,N_6169,N_8755);
xor U9413 (N_9413,N_8941,N_8653);
or U9414 (N_9414,N_8621,N_8623);
and U9415 (N_9415,N_7175,N_7023);
nor U9416 (N_9416,N_8160,N_7731);
nor U9417 (N_9417,N_7909,N_8724);
or U9418 (N_9418,N_8892,N_8834);
nand U9419 (N_9419,N_7014,N_7357);
and U9420 (N_9420,N_6028,N_7749);
or U9421 (N_9421,N_7434,N_8325);
and U9422 (N_9422,N_8273,N_6835);
nand U9423 (N_9423,N_6067,N_8280);
and U9424 (N_9424,N_6564,N_7971);
nor U9425 (N_9425,N_8184,N_6546);
nor U9426 (N_9426,N_7744,N_8891);
or U9427 (N_9427,N_6488,N_7886);
nor U9428 (N_9428,N_8261,N_8863);
or U9429 (N_9429,N_6754,N_8256);
nor U9430 (N_9430,N_7602,N_7371);
nand U9431 (N_9431,N_7187,N_7810);
nand U9432 (N_9432,N_6084,N_7144);
nor U9433 (N_9433,N_6193,N_6717);
nor U9434 (N_9434,N_8005,N_8689);
or U9435 (N_9435,N_8702,N_6615);
nor U9436 (N_9436,N_6764,N_7891);
and U9437 (N_9437,N_7384,N_6576);
nor U9438 (N_9438,N_7721,N_7264);
and U9439 (N_9439,N_7205,N_8195);
nor U9440 (N_9440,N_7764,N_8416);
or U9441 (N_9441,N_8197,N_6047);
nand U9442 (N_9442,N_8944,N_7045);
nor U9443 (N_9443,N_7173,N_8147);
and U9444 (N_9444,N_7487,N_7663);
or U9445 (N_9445,N_7042,N_6929);
nand U9446 (N_9446,N_8376,N_6180);
or U9447 (N_9447,N_8137,N_6348);
nand U9448 (N_9448,N_6137,N_6629);
or U9449 (N_9449,N_7364,N_8259);
or U9450 (N_9450,N_7950,N_7050);
nor U9451 (N_9451,N_6675,N_6884);
nand U9452 (N_9452,N_8842,N_7060);
nand U9453 (N_9453,N_7567,N_8494);
and U9454 (N_9454,N_7797,N_8402);
and U9455 (N_9455,N_8169,N_8657);
nor U9456 (N_9456,N_7547,N_8046);
or U9457 (N_9457,N_8540,N_7787);
nand U9458 (N_9458,N_8095,N_7284);
nand U9459 (N_9459,N_8730,N_6257);
nand U9460 (N_9460,N_8720,N_6803);
nand U9461 (N_9461,N_7366,N_8589);
xnor U9462 (N_9462,N_8675,N_8556);
or U9463 (N_9463,N_7719,N_6799);
nand U9464 (N_9464,N_7563,N_6030);
or U9465 (N_9465,N_8698,N_6863);
or U9466 (N_9466,N_8606,N_8301);
nand U9467 (N_9467,N_7132,N_6819);
or U9468 (N_9468,N_8946,N_7123);
and U9469 (N_9469,N_6673,N_8004);
nor U9470 (N_9470,N_6043,N_7141);
nor U9471 (N_9471,N_6918,N_6328);
or U9472 (N_9472,N_8470,N_7792);
nor U9473 (N_9473,N_6042,N_8202);
or U9474 (N_9474,N_8910,N_8595);
and U9475 (N_9475,N_8397,N_6682);
or U9476 (N_9476,N_8336,N_8704);
or U9477 (N_9477,N_8140,N_8553);
nor U9478 (N_9478,N_8318,N_7771);
or U9479 (N_9479,N_6238,N_7537);
nor U9480 (N_9480,N_8368,N_6535);
nand U9481 (N_9481,N_7204,N_6002);
and U9482 (N_9482,N_8040,N_6133);
and U9483 (N_9483,N_7774,N_7131);
and U9484 (N_9484,N_8934,N_7895);
nor U9485 (N_9485,N_7178,N_6074);
nor U9486 (N_9486,N_8133,N_7591);
nor U9487 (N_9487,N_7887,N_7237);
or U9488 (N_9488,N_8634,N_8105);
and U9489 (N_9489,N_6275,N_6945);
or U9490 (N_9490,N_8469,N_6734);
and U9491 (N_9491,N_8997,N_6885);
or U9492 (N_9492,N_6730,N_8239);
nand U9493 (N_9493,N_6905,N_7695);
nor U9494 (N_9494,N_8966,N_8253);
and U9495 (N_9495,N_7523,N_7122);
and U9496 (N_9496,N_6781,N_7512);
nor U9497 (N_9497,N_7240,N_7670);
nand U9498 (N_9498,N_7831,N_6997);
nor U9499 (N_9499,N_6396,N_7113);
nand U9500 (N_9500,N_7037,N_8417);
nor U9501 (N_9501,N_7999,N_7036);
nand U9502 (N_9502,N_6177,N_6685);
nor U9503 (N_9503,N_8956,N_8901);
nand U9504 (N_9504,N_8695,N_6387);
nor U9505 (N_9505,N_6579,N_6479);
nor U9506 (N_9506,N_7249,N_6908);
xor U9507 (N_9507,N_6868,N_7473);
nor U9508 (N_9508,N_6243,N_6166);
nor U9509 (N_9509,N_6696,N_6976);
nor U9510 (N_9510,N_7935,N_6006);
nand U9511 (N_9511,N_7738,N_8018);
xor U9512 (N_9512,N_6946,N_7737);
and U9513 (N_9513,N_6613,N_7157);
or U9514 (N_9514,N_6807,N_6897);
nor U9515 (N_9515,N_6973,N_8685);
nor U9516 (N_9516,N_7762,N_6812);
nor U9517 (N_9517,N_6051,N_8285);
or U9518 (N_9518,N_8268,N_8557);
nor U9519 (N_9519,N_8395,N_6953);
nor U9520 (N_9520,N_7075,N_8958);
nand U9521 (N_9521,N_7786,N_8625);
or U9522 (N_9522,N_8742,N_6921);
or U9523 (N_9523,N_6250,N_6220);
nand U9524 (N_9524,N_6539,N_6378);
nor U9525 (N_9525,N_8830,N_8216);
nor U9526 (N_9526,N_7054,N_6670);
or U9527 (N_9527,N_6608,N_8977);
and U9528 (N_9528,N_8217,N_7593);
and U9529 (N_9529,N_8179,N_8384);
or U9530 (N_9530,N_8894,N_8960);
and U9531 (N_9531,N_8479,N_6725);
and U9532 (N_9532,N_8355,N_8434);
nand U9533 (N_9533,N_8225,N_7053);
and U9534 (N_9534,N_6405,N_7981);
and U9535 (N_9535,N_8506,N_6584);
and U9536 (N_9536,N_8539,N_6280);
nand U9537 (N_9537,N_8343,N_8950);
and U9538 (N_9538,N_7495,N_6254);
or U9539 (N_9539,N_8579,N_8658);
nor U9540 (N_9540,N_8274,N_8725);
or U9541 (N_9541,N_7894,N_6871);
and U9542 (N_9542,N_7588,N_6236);
or U9543 (N_9543,N_6646,N_6784);
nand U9544 (N_9544,N_8663,N_7671);
nand U9545 (N_9545,N_6983,N_8747);
xnor U9546 (N_9546,N_6313,N_7550);
or U9547 (N_9547,N_7405,N_8313);
nand U9548 (N_9548,N_8542,N_6418);
nand U9549 (N_9549,N_6127,N_6211);
nand U9550 (N_9550,N_8521,N_7943);
nand U9551 (N_9551,N_6339,N_6733);
and U9552 (N_9552,N_6738,N_7709);
nand U9553 (N_9553,N_6070,N_6195);
nand U9554 (N_9554,N_6095,N_6599);
or U9555 (N_9555,N_6283,N_6590);
nand U9556 (N_9556,N_6653,N_6780);
nand U9557 (N_9557,N_6270,N_7964);
nand U9558 (N_9558,N_7118,N_7465);
or U9559 (N_9559,N_8587,N_7606);
or U9560 (N_9560,N_8257,N_6390);
nand U9561 (N_9561,N_8736,N_8715);
nand U9562 (N_9562,N_6623,N_8489);
or U9563 (N_9563,N_8923,N_6005);
xnor U9564 (N_9564,N_6501,N_8096);
nand U9565 (N_9565,N_8181,N_8145);
nor U9566 (N_9566,N_7011,N_8586);
nor U9567 (N_9567,N_7985,N_6627);
xor U9568 (N_9568,N_8734,N_8218);
nand U9569 (N_9569,N_7833,N_6582);
nor U9570 (N_9570,N_7616,N_8054);
nor U9571 (N_9571,N_6112,N_6011);
nand U9572 (N_9572,N_7975,N_8827);
nand U9573 (N_9573,N_6175,N_6398);
and U9574 (N_9574,N_8236,N_6986);
nand U9575 (N_9575,N_8840,N_7691);
or U9576 (N_9576,N_7904,N_6235);
or U9577 (N_9577,N_8565,N_8569);
or U9578 (N_9578,N_6575,N_8613);
nand U9579 (N_9579,N_8398,N_6740);
or U9580 (N_9580,N_7980,N_8786);
and U9581 (N_9581,N_6340,N_7682);
and U9582 (N_9582,N_8519,N_7194);
and U9583 (N_9583,N_6464,N_6702);
and U9584 (N_9584,N_6797,N_8649);
or U9585 (N_9585,N_6239,N_7976);
and U9586 (N_9586,N_6096,N_6844);
or U9587 (N_9587,N_6364,N_7133);
nand U9588 (N_9588,N_8544,N_8446);
nand U9589 (N_9589,N_6126,N_8033);
nor U9590 (N_9590,N_7680,N_6116);
nand U9591 (N_9591,N_7253,N_7622);
and U9592 (N_9592,N_6496,N_8353);
nor U9593 (N_9593,N_6693,N_7408);
nor U9594 (N_9594,N_7161,N_8849);
xnor U9595 (N_9595,N_6984,N_6596);
nand U9596 (N_9596,N_8678,N_8168);
or U9597 (N_9597,N_6134,N_6259);
nand U9598 (N_9598,N_6855,N_8696);
and U9599 (N_9599,N_6487,N_8464);
nor U9600 (N_9600,N_6568,N_8741);
and U9601 (N_9601,N_7290,N_7193);
nor U9602 (N_9602,N_6269,N_6382);
and U9603 (N_9603,N_6574,N_8128);
or U9604 (N_9604,N_7185,N_8737);
nor U9605 (N_9605,N_7908,N_7997);
nand U9606 (N_9606,N_7988,N_7843);
and U9607 (N_9607,N_8210,N_6992);
and U9608 (N_9608,N_6377,N_7126);
and U9609 (N_9609,N_8073,N_6612);
and U9610 (N_9610,N_7956,N_8626);
nand U9611 (N_9611,N_7517,N_7672);
nand U9612 (N_9612,N_8315,N_6928);
and U9613 (N_9613,N_7061,N_6399);
nor U9614 (N_9614,N_7582,N_6310);
nand U9615 (N_9615,N_7186,N_6491);
or U9616 (N_9616,N_7496,N_7529);
nor U9617 (N_9617,N_7714,N_7034);
and U9618 (N_9618,N_8458,N_7015);
and U9619 (N_9619,N_7590,N_8244);
or U9620 (N_9620,N_8091,N_6531);
nor U9621 (N_9621,N_7690,N_6062);
nand U9622 (N_9622,N_8045,N_8472);
and U9623 (N_9623,N_8199,N_7312);
nor U9624 (N_9624,N_7058,N_6350);
nor U9625 (N_9625,N_8862,N_6045);
and U9626 (N_9626,N_6542,N_7990);
nand U9627 (N_9627,N_7882,N_6012);
nor U9628 (N_9628,N_7301,N_7028);
or U9629 (N_9629,N_7519,N_8921);
nand U9630 (N_9630,N_6499,N_8797);
and U9631 (N_9631,N_6643,N_8111);
and U9632 (N_9632,N_7934,N_6829);
or U9633 (N_9633,N_6647,N_7016);
nand U9634 (N_9634,N_6707,N_8439);
or U9635 (N_9635,N_8571,N_7064);
and U9636 (N_9636,N_6750,N_8049);
nor U9637 (N_9637,N_7739,N_6761);
nor U9638 (N_9638,N_8308,N_6104);
or U9639 (N_9639,N_6678,N_8588);
or U9640 (N_9640,N_6139,N_7049);
or U9641 (N_9641,N_6721,N_7767);
or U9642 (N_9642,N_8633,N_8743);
and U9643 (N_9643,N_8389,N_6320);
nor U9644 (N_9644,N_8003,N_7790);
nor U9645 (N_9645,N_8971,N_6072);
xnor U9646 (N_9646,N_6432,N_6140);
nor U9647 (N_9647,N_6289,N_7995);
nor U9648 (N_9648,N_8364,N_7947);
and U9649 (N_9649,N_7631,N_8334);
or U9650 (N_9650,N_7822,N_6614);
xor U9651 (N_9651,N_7481,N_7867);
and U9652 (N_9652,N_7699,N_6343);
nand U9653 (N_9653,N_7715,N_7518);
nor U9654 (N_9654,N_7458,N_7353);
nand U9655 (N_9655,N_8349,N_8360);
nand U9656 (N_9656,N_6149,N_7336);
and U9657 (N_9657,N_6739,N_6515);
or U9658 (N_9658,N_7412,N_8229);
nand U9659 (N_9659,N_6775,N_6662);
and U9660 (N_9660,N_7365,N_7871);
or U9661 (N_9661,N_6778,N_8345);
or U9662 (N_9662,N_6316,N_7207);
nor U9663 (N_9663,N_7857,N_7723);
nand U9664 (N_9664,N_7658,N_8879);
nand U9665 (N_9665,N_7679,N_8713);
or U9666 (N_9666,N_7634,N_7704);
or U9667 (N_9667,N_6726,N_7195);
and U9668 (N_9668,N_7979,N_8267);
nand U9669 (N_9669,N_6204,N_7116);
and U9670 (N_9670,N_8451,N_6007);
or U9671 (N_9671,N_8404,N_8538);
xor U9672 (N_9672,N_6431,N_8692);
and U9673 (N_9673,N_6713,N_6609);
and U9674 (N_9674,N_7316,N_8454);
nor U9675 (N_9675,N_6407,N_8443);
nand U9676 (N_9676,N_7662,N_7229);
nand U9677 (N_9677,N_6559,N_7352);
nand U9678 (N_9678,N_7472,N_8801);
nor U9679 (N_9679,N_7949,N_8943);
and U9680 (N_9680,N_6356,N_7389);
nor U9681 (N_9681,N_8607,N_6700);
nand U9682 (N_9682,N_8248,N_6845);
or U9683 (N_9683,N_7637,N_8745);
and U9684 (N_9684,N_6964,N_8723);
nor U9685 (N_9685,N_7698,N_6114);
and U9686 (N_9686,N_6138,N_8493);
xor U9687 (N_9687,N_8561,N_7376);
nand U9688 (N_9688,N_8065,N_8778);
nor U9689 (N_9689,N_8071,N_7953);
and U9690 (N_9690,N_7250,N_8444);
and U9691 (N_9691,N_7646,N_6066);
nand U9692 (N_9692,N_6709,N_6498);
nor U9693 (N_9693,N_8407,N_7417);
or U9694 (N_9694,N_7314,N_7983);
nand U9695 (N_9695,N_8808,N_6189);
or U9696 (N_9696,N_6255,N_7243);
and U9697 (N_9697,N_8228,N_7888);
or U9698 (N_9698,N_8420,N_7222);
or U9699 (N_9699,N_6486,N_7600);
or U9700 (N_9700,N_8299,N_6246);
nand U9701 (N_9701,N_8109,N_6637);
nand U9702 (N_9702,N_7244,N_8471);
xor U9703 (N_9703,N_6253,N_6753);
nor U9704 (N_9704,N_8632,N_7359);
nand U9705 (N_9705,N_6617,N_6397);
and U9706 (N_9706,N_7753,N_6794);
and U9707 (N_9707,N_8779,N_7573);
nand U9708 (N_9708,N_7836,N_6694);
and U9709 (N_9709,N_6384,N_7022);
or U9710 (N_9710,N_8924,N_6981);
nand U9711 (N_9711,N_8366,N_8503);
or U9712 (N_9712,N_7171,N_8970);
and U9713 (N_9713,N_6060,N_6098);
nor U9714 (N_9714,N_8344,N_8254);
or U9715 (N_9715,N_8131,N_7407);
nand U9716 (N_9716,N_8661,N_7216);
nand U9717 (N_9717,N_8367,N_8576);
or U9718 (N_9718,N_7480,N_8436);
or U9719 (N_9719,N_8311,N_6645);
and U9720 (N_9720,N_8317,N_8135);
nor U9721 (N_9721,N_8551,N_6795);
nand U9722 (N_9722,N_8250,N_8995);
or U9723 (N_9723,N_8495,N_6860);
or U9724 (N_9724,N_8245,N_6124);
nand U9725 (N_9725,N_7246,N_7339);
nand U9726 (N_9726,N_6383,N_8975);
nor U9727 (N_9727,N_7585,N_7627);
nor U9728 (N_9728,N_7556,N_8332);
or U9729 (N_9729,N_7169,N_6157);
nand U9730 (N_9730,N_8815,N_7678);
nand U9731 (N_9731,N_7013,N_6152);
nand U9732 (N_9732,N_6505,N_7579);
and U9733 (N_9733,N_7277,N_8908);
nand U9734 (N_9734,N_6038,N_6287);
and U9735 (N_9735,N_6891,N_6256);
nand U9736 (N_9736,N_8552,N_7265);
nor U9737 (N_9737,N_6924,N_7198);
or U9738 (N_9738,N_6247,N_8178);
nand U9739 (N_9739,N_6814,N_8939);
nand U9740 (N_9740,N_7494,N_8496);
nor U9741 (N_9741,N_8129,N_8822);
nor U9742 (N_9742,N_8938,N_8305);
nand U9743 (N_9743,N_6164,N_7713);
nor U9744 (N_9744,N_7188,N_7968);
or U9745 (N_9745,N_8209,N_7217);
nand U9746 (N_9746,N_7415,N_6601);
and U9747 (N_9747,N_6630,N_7884);
or U9748 (N_9748,N_8688,N_8012);
or U9749 (N_9749,N_8680,N_6788);
nor U9750 (N_9750,N_8523,N_6961);
nor U9751 (N_9751,N_7839,N_8085);
nand U9752 (N_9752,N_8775,N_6457);
or U9753 (N_9753,N_6998,N_6119);
and U9754 (N_9754,N_7791,N_8705);
or U9755 (N_9755,N_6943,N_8447);
nand U9756 (N_9756,N_6914,N_8930);
or U9757 (N_9757,N_8673,N_6037);
or U9758 (N_9758,N_8594,N_8487);
or U9759 (N_9759,N_7944,N_6968);
and U9760 (N_9760,N_8093,N_7012);
nor U9761 (N_9761,N_7740,N_7525);
nand U9762 (N_9762,N_8327,N_8214);
and U9763 (N_9763,N_7761,N_8510);
or U9764 (N_9764,N_6217,N_7272);
nand U9765 (N_9765,N_8902,N_7107);
and U9766 (N_9766,N_8701,N_8126);
and U9767 (N_9767,N_7752,N_7717);
or U9768 (N_9768,N_6089,N_6883);
nor U9769 (N_9769,N_6344,N_8855);
and U9770 (N_9770,N_8585,N_7477);
nor U9771 (N_9771,N_7743,N_8117);
nor U9772 (N_9772,N_6589,N_7271);
and U9773 (N_9773,N_6209,N_8211);
nor U9774 (N_9774,N_8144,N_7019);
nor U9775 (N_9775,N_7342,N_6526);
and U9776 (N_9776,N_7268,N_8819);
nand U9777 (N_9777,N_8514,N_7215);
and U9778 (N_9778,N_6554,N_8857);
and U9779 (N_9779,N_6249,N_6454);
xnor U9780 (N_9780,N_7946,N_6512);
or U9781 (N_9781,N_6938,N_7555);
xnor U9782 (N_9782,N_6716,N_7736);
or U9783 (N_9783,N_8803,N_8200);
or U9784 (N_9784,N_8113,N_7070);
xor U9785 (N_9785,N_6061,N_7954);
nor U9786 (N_9786,N_7427,N_8335);
and U9787 (N_9787,N_6321,N_8753);
nand U9788 (N_9788,N_8752,N_6544);
or U9789 (N_9789,N_7847,N_6336);
nor U9790 (N_9790,N_6120,N_8252);
nor U9791 (N_9791,N_6857,N_8584);
nand U9792 (N_9792,N_6460,N_8502);
nor U9793 (N_9793,N_6684,N_7994);
or U9794 (N_9794,N_7660,N_7766);
nand U9795 (N_9795,N_6881,N_6798);
or U9796 (N_9796,N_8712,N_8972);
nand U9797 (N_9797,N_8437,N_7665);
xnor U9798 (N_9798,N_8532,N_6185);
nand U9799 (N_9799,N_8865,N_7906);
or U9800 (N_9800,N_7463,N_8242);
xor U9801 (N_9801,N_8122,N_8670);
or U9802 (N_9802,N_7274,N_8312);
and U9803 (N_9803,N_7808,N_7838);
and U9804 (N_9804,N_7522,N_7167);
and U9805 (N_9805,N_7789,N_6207);
or U9806 (N_9806,N_8534,N_7254);
and U9807 (N_9807,N_8485,N_8077);
and U9808 (N_9808,N_8872,N_8370);
nor U9809 (N_9809,N_8969,N_8286);
or U9810 (N_9810,N_8764,N_7607);
nor U9811 (N_9811,N_6789,N_6910);
nand U9812 (N_9812,N_8599,N_8328);
and U9813 (N_9813,N_8371,N_7108);
nand U9814 (N_9814,N_8086,N_8190);
or U9815 (N_9815,N_6000,N_7478);
and U9816 (N_9816,N_8339,N_8051);
and U9817 (N_9817,N_8037,N_8762);
xor U9818 (N_9818,N_7570,N_8728);
and U9819 (N_9819,N_7489,N_6747);
or U9820 (N_9820,N_7317,N_7777);
nand U9821 (N_9821,N_6527,N_8176);
and U9822 (N_9822,N_6108,N_7416);
and U9823 (N_9823,N_7881,N_8929);
nor U9824 (N_9824,N_6044,N_6376);
or U9825 (N_9825,N_7121,N_7162);
or U9826 (N_9826,N_8968,N_8173);
nor U9827 (N_9827,N_7476,N_8622);
nor U9828 (N_9828,N_6543,N_7586);
nor U9829 (N_9829,N_6714,N_7464);
nand U9830 (N_9830,N_8529,N_7644);
xnor U9831 (N_9831,N_6301,N_7398);
nor U9832 (N_9832,N_7258,N_6806);
and U9833 (N_9833,N_6631,N_7558);
and U9834 (N_9834,N_6033,N_8112);
nand U9835 (N_9835,N_7630,N_8610);
nand U9836 (N_9836,N_7300,N_8053);
and U9837 (N_9837,N_8092,N_7039);
and U9838 (N_9838,N_7411,N_6208);
nor U9839 (N_9839,N_6796,N_6877);
xor U9840 (N_9840,N_7902,N_7307);
nor U9841 (N_9841,N_6265,N_8425);
or U9842 (N_9842,N_7673,N_8015);
or U9843 (N_9843,N_8422,N_6290);
or U9844 (N_9844,N_8665,N_7041);
xor U9845 (N_9845,N_7900,N_7238);
or U9846 (N_9846,N_7040,N_7832);
nor U9847 (N_9847,N_8141,N_7722);
nand U9848 (N_9848,N_7802,N_6288);
nor U9849 (N_9849,N_6036,N_8627);
or U9850 (N_9850,N_7756,N_6415);
or U9851 (N_9851,N_6760,N_7601);
nor U9852 (N_9852,N_7142,N_6875);
nor U9853 (N_9853,N_7457,N_7724);
nor U9854 (N_9854,N_7520,N_6401);
nor U9855 (N_9855,N_6839,N_7633);
nand U9856 (N_9856,N_8802,N_8130);
nor U9857 (N_9857,N_6023,N_7388);
and U9858 (N_9858,N_7683,N_8572);
or U9859 (N_9859,N_6583,N_7304);
or U9860 (N_9860,N_6800,N_6425);
nand U9861 (N_9861,N_8710,N_7462);
or U9862 (N_9862,N_8522,N_8059);
or U9863 (N_9863,N_6811,N_8501);
nand U9864 (N_9864,N_8408,N_6837);
and U9865 (N_9865,N_7921,N_8278);
nor U9866 (N_9866,N_8558,N_8833);
nor U9867 (N_9867,N_6858,N_6974);
nor U9868 (N_9868,N_8591,N_6113);
nand U9869 (N_9869,N_8377,N_6573);
and U9870 (N_9870,N_8044,N_6225);
and U9871 (N_9871,N_8468,N_7135);
and U9872 (N_9872,N_7958,N_7806);
nor U9873 (N_9873,N_8201,N_8356);
nor U9874 (N_9874,N_6426,N_8504);
nor U9875 (N_9875,N_6115,N_8084);
nand U9876 (N_9876,N_7154,N_7647);
or U9877 (N_9877,N_6690,N_8848);
or U9878 (N_9878,N_8426,N_8150);
or U9879 (N_9879,N_6511,N_8321);
and U9880 (N_9880,N_6859,N_7319);
or U9881 (N_9881,N_7206,N_7283);
or U9882 (N_9882,N_6305,N_6913);
nor U9883 (N_9883,N_7720,N_7705);
or U9884 (N_9884,N_7286,N_6688);
nand U9885 (N_9885,N_6507,N_6912);
nor U9886 (N_9886,N_6272,N_8075);
nand U9887 (N_9887,N_7773,N_6151);
nand U9888 (N_9888,N_8226,N_7551);
or U9889 (N_9889,N_8654,N_7241);
nor U9890 (N_9890,N_6842,N_8580);
nor U9891 (N_9891,N_7486,N_7747);
nor U9892 (N_9892,N_7689,N_8013);
and U9893 (N_9893,N_6136,N_7363);
and U9894 (N_9894,N_6533,N_6777);
xor U9895 (N_9895,N_6103,N_6985);
and U9896 (N_9896,N_8949,N_6264);
or U9897 (N_9897,N_8107,N_8711);
nand U9898 (N_9898,N_6625,N_6163);
or U9899 (N_9899,N_7393,N_6322);
or U9900 (N_9900,N_7263,N_7686);
and U9901 (N_9901,N_7425,N_6052);
nor U9902 (N_9902,N_8338,N_7820);
or U9903 (N_9903,N_7112,N_6765);
nand U9904 (N_9904,N_8574,N_6851);
and U9905 (N_9905,N_7898,N_6624);
and U9906 (N_9906,N_8478,N_7294);
nor U9907 (N_9907,N_7874,N_8372);
nand U9908 (N_9908,N_6864,N_8864);
or U9909 (N_9909,N_8304,N_8352);
nand U9910 (N_9910,N_6537,N_7989);
or U9911 (N_9911,N_7095,N_7328);
nand U9912 (N_9912,N_8985,N_8861);
and U9913 (N_9913,N_7572,N_7514);
or U9914 (N_9914,N_7331,N_6427);
and U9915 (N_9915,N_7580,N_6248);
and U9916 (N_9916,N_6159,N_8060);
and U9917 (N_9917,N_6419,N_8047);
or U9918 (N_9918,N_6031,N_6766);
nor U9919 (N_9919,N_6429,N_7150);
or U9920 (N_9920,N_7965,N_7903);
nor U9921 (N_9921,N_8058,N_8771);
and U9922 (N_9922,N_7103,N_7114);
and U9923 (N_9923,N_8148,N_7059);
and U9924 (N_9924,N_6951,N_7347);
nand U9925 (N_9925,N_7885,N_8302);
and U9926 (N_9926,N_6681,N_7297);
or U9927 (N_9927,N_6230,N_8401);
and U9928 (N_9928,N_8279,N_6009);
or U9929 (N_9929,N_6534,N_6715);
nand U9930 (N_9930,N_8283,N_8187);
and U9931 (N_9931,N_7538,N_8805);
and U9932 (N_9932,N_6772,N_7006);
and U9933 (N_9933,N_8766,N_8359);
nor U9934 (N_9934,N_7553,N_7667);
nor U9935 (N_9935,N_7007,N_8429);
nand U9936 (N_9936,N_7732,N_8240);
or U9937 (N_9937,N_6571,N_7318);
and U9938 (N_9938,N_8841,N_6055);
nand U9939 (N_9939,N_6980,N_7652);
and U9940 (N_9940,N_6329,N_7608);
nor U9941 (N_9941,N_7323,N_6100);
nand U9942 (N_9942,N_7526,N_8411);
or U9943 (N_9943,N_6954,N_6215);
and U9944 (N_9944,N_7620,N_7460);
nand U9945 (N_9945,N_8899,N_8381);
nor U9946 (N_9946,N_8149,N_8337);
or U9947 (N_9947,N_7181,N_8188);
or U9948 (N_9948,N_7201,N_7212);
and U9949 (N_9949,N_7164,N_6959);
or U9950 (N_9950,N_6654,N_7729);
or U9951 (N_9951,N_6001,N_6170);
and U9952 (N_9952,N_8165,N_7565);
nand U9953 (N_9953,N_8818,N_8088);
nand U9954 (N_9954,N_8032,N_7681);
nand U9955 (N_9955,N_6245,N_6161);
nor U9956 (N_9956,N_6870,N_7282);
nor U9957 (N_9957,N_6720,N_8650);
and U9958 (N_9958,N_6150,N_6683);
or U9959 (N_9959,N_7901,N_6581);
and U9960 (N_9960,N_6370,N_8955);
or U9961 (N_9961,N_7578,N_6975);
and U9962 (N_9962,N_7957,N_6657);
or U9963 (N_9963,N_8851,N_7248);
nand U9964 (N_9964,N_6547,N_6972);
or U9965 (N_9965,N_6718,N_6663);
nor U9966 (N_9966,N_7419,N_7872);
nand U9967 (N_9967,N_8017,N_6307);
and U9968 (N_9968,N_7289,N_8881);
nand U9969 (N_9969,N_8484,N_7020);
nand U9970 (N_9970,N_8196,N_6606);
nand U9971 (N_9971,N_8198,N_8664);
nand U9972 (N_9972,N_8641,N_6091);
nand U9973 (N_9973,N_8976,N_6162);
and U9974 (N_9974,N_8602,N_7446);
nor U9975 (N_9975,N_7527,N_6852);
and U9976 (N_9976,N_7974,N_7176);
and U9977 (N_9977,N_7467,N_8341);
and U9978 (N_9978,N_8854,N_8342);
and U9979 (N_9979,N_7435,N_6732);
or U9980 (N_9980,N_6558,N_6300);
and U9981 (N_9981,N_7035,N_6130);
nor U9982 (N_9982,N_8763,N_8746);
or U9983 (N_9983,N_6406,N_6904);
or U9984 (N_9984,N_8525,N_6603);
and U9985 (N_9985,N_7260,N_7373);
or U9986 (N_9986,N_7184,N_7824);
nand U9987 (N_9987,N_8249,N_8123);
or U9988 (N_9988,N_7942,N_7584);
xnor U9989 (N_9989,N_6231,N_6173);
nor U9990 (N_9990,N_6046,N_6538);
nand U9991 (N_9991,N_7493,N_8907);
nand U9992 (N_9992,N_7471,N_6996);
nand U9993 (N_9993,N_8718,N_6421);
or U9994 (N_9994,N_6224,N_8260);
or U9995 (N_9995,N_6605,N_8640);
and U9996 (N_9996,N_7358,N_7077);
nand U9997 (N_9997,N_7676,N_6820);
nand U9998 (N_9998,N_8564,N_7959);
xnor U9999 (N_9999,N_8813,N_8090);
or U10000 (N_10000,N_8440,N_7549);
or U10001 (N_10001,N_8795,N_7148);
or U10002 (N_10002,N_7315,N_6767);
and U10003 (N_10003,N_6552,N_7174);
and U10004 (N_10004,N_7410,N_7837);
or U10005 (N_10005,N_8608,N_6949);
nor U10006 (N_10006,N_6658,N_6069);
nor U10007 (N_10007,N_6094,N_6666);
and U10008 (N_10008,N_6687,N_8691);
nand U10009 (N_10009,N_7557,N_7047);
nor U10010 (N_10010,N_7758,N_6381);
nand U10011 (N_10011,N_7324,N_8477);
or U10012 (N_10012,N_7090,N_6886);
or U10013 (N_10013,N_6500,N_6832);
and U10014 (N_10014,N_7420,N_6659);
nor U10015 (N_10015,N_7492,N_6093);
nor U10016 (N_10016,N_7559,N_6319);
or U10017 (N_10017,N_6414,N_6294);
nand U10018 (N_10018,N_7137,N_8916);
nand U10019 (N_10019,N_8410,N_7003);
nand U10020 (N_10020,N_6342,N_8825);
nand U10021 (N_10021,N_6898,N_6154);
and U10022 (N_10022,N_8951,N_6580);
xor U10023 (N_10023,N_6644,N_6545);
and U10024 (N_10024,N_7479,N_6197);
nor U10025 (N_10025,N_6933,N_7048);
nand U10026 (N_10026,N_8731,N_7628);
or U10027 (N_10027,N_6291,N_8189);
nand U10028 (N_10028,N_8765,N_7355);
nor U10029 (N_10029,N_8089,N_8241);
nand U10030 (N_10030,N_6999,N_7649);
nand U10031 (N_10031,N_7609,N_6490);
or U10032 (N_10032,N_7320,N_8114);
or U10033 (N_10033,N_7456,N_8159);
nand U10034 (N_10034,N_7348,N_8509);
and U10035 (N_10035,N_6560,N_7708);
nor U10036 (N_10036,N_6919,N_6099);
or U10037 (N_10037,N_7091,N_8172);
nand U10038 (N_10038,N_7993,N_7351);
or U10039 (N_10039,N_8243,N_8846);
xnor U10040 (N_10040,N_8947,N_6944);
nand U10041 (N_10041,N_8582,N_6065);
and U10042 (N_10042,N_8505,N_6271);
or U10043 (N_10043,N_8213,N_6360);
or U10044 (N_10044,N_6660,N_7712);
nand U10045 (N_10045,N_6966,N_6993);
nor U10046 (N_10046,N_8428,N_6417);
or U10047 (N_10047,N_7960,N_6843);
nor U10048 (N_10048,N_7120,N_6458);
nand U10049 (N_10049,N_6444,N_8296);
nand U10050 (N_10050,N_8716,N_8031);
nor U10051 (N_10051,N_7978,N_6357);
nand U10052 (N_10052,N_8922,N_8347);
nor U10053 (N_10053,N_6434,N_7104);
and U10054 (N_10054,N_6456,N_7982);
nor U10055 (N_10055,N_7733,N_6524);
nor U10056 (N_10056,N_8517,N_8690);
and U10057 (N_10057,N_6311,N_6804);
and U10058 (N_10058,N_8433,N_8856);
nand U10059 (N_10059,N_6160,N_8378);
or U10060 (N_10060,N_8798,N_8055);
nand U10061 (N_10061,N_7560,N_7688);
or U10062 (N_10062,N_6053,N_7566);
and U10063 (N_10063,N_6371,N_8474);
or U10064 (N_10064,N_6437,N_6889);
or U10065 (N_10065,N_8108,N_8583);
or U10066 (N_10066,N_7858,N_8667);
or U10067 (N_10067,N_7638,N_7299);
nor U10068 (N_10068,N_6762,N_8733);
and U10069 (N_10069,N_6586,N_8918);
nor U10070 (N_10070,N_8421,N_7098);
and U10071 (N_10071,N_6346,N_6489);
nor U10072 (N_10072,N_6085,N_7991);
nor U10073 (N_10073,N_8021,N_7853);
nor U10074 (N_10074,N_6481,N_6572);
or U10075 (N_10075,N_7341,N_6703);
nand U10076 (N_10076,N_7484,N_7922);
nor U10077 (N_10077,N_7031,N_7613);
or U10078 (N_10078,N_7356,N_6462);
nor U10079 (N_10079,N_6128,N_6942);
or U10080 (N_10080,N_8455,N_8547);
and U10081 (N_10081,N_6354,N_6557);
or U10082 (N_10082,N_6978,N_7236);
nand U10083 (N_10083,N_6639,N_8265);
and U10084 (N_10084,N_7370,N_7329);
or U10085 (N_10085,N_8483,N_6616);
nand U10086 (N_10086,N_8573,N_6110);
xnor U10087 (N_10087,N_6746,N_7765);
or U10088 (N_10088,N_8869,N_8697);
nand U10089 (N_10089,N_7273,N_6866);
and U10090 (N_10090,N_8331,N_6665);
and U10091 (N_10091,N_7303,N_7966);
and U10092 (N_10092,N_6679,N_8412);
nand U10093 (N_10093,N_6494,N_7855);
or U10094 (N_10094,N_8643,N_7490);
nand U10095 (N_10095,N_6849,N_7816);
or U10096 (N_10096,N_6600,N_6242);
nor U10097 (N_10097,N_8836,N_8883);
or U10098 (N_10098,N_8933,N_6282);
or U10099 (N_10099,N_7914,N_6267);
nand U10100 (N_10100,N_8212,N_7716);
nor U10101 (N_10101,N_7083,N_8992);
and U10102 (N_10102,N_6610,N_8722);
nor U10103 (N_10103,N_8794,N_7027);
nor U10104 (N_10104,N_6299,N_6039);
nand U10105 (N_10105,N_8388,N_8598);
nand U10106 (N_10106,N_8672,N_7455);
or U10107 (N_10107,N_8520,N_6206);
nor U10108 (N_10108,N_8882,N_7409);
nand U10109 (N_10109,N_6025,N_7288);
nand U10110 (N_10110,N_6218,N_7801);
nand U10111 (N_10111,N_6521,N_7626);
and U10112 (N_10112,N_8132,N_6184);
or U10113 (N_10113,N_8973,N_7796);
or U10114 (N_10114,N_6988,N_7068);
nand U10115 (N_10115,N_6059,N_6395);
or U10116 (N_10116,N_8537,N_8449);
nand U10117 (N_10117,N_6977,N_7592);
nand U10118 (N_10118,N_7880,N_7436);
or U10119 (N_10119,N_7469,N_7636);
and U10120 (N_10120,N_8456,N_8396);
and U10121 (N_10121,N_8508,N_7896);
or U10122 (N_10122,N_6793,N_6068);
nor U10123 (N_10123,N_7343,N_6261);
and U10124 (N_10124,N_8120,N_8563);
xor U10125 (N_10125,N_6722,N_7190);
or U10126 (N_10126,N_6566,N_6661);
and U10127 (N_10127,N_6805,N_8457);
nand U10128 (N_10128,N_6597,N_6123);
nand U10129 (N_10129,N_7554,N_7918);
and U10130 (N_10130,N_7877,N_7998);
or U10131 (N_10131,N_7863,N_6374);
nor U10132 (N_10132,N_8183,N_7311);
nand U10133 (N_10133,N_7066,N_6296);
or U10134 (N_10134,N_6202,N_6118);
or U10135 (N_10135,N_8019,N_8363);
or U10136 (N_10136,N_7183,N_6461);
nor U10137 (N_10137,N_8671,N_8928);
and U10138 (N_10138,N_8904,N_7807);
and U10139 (N_10139,N_8832,N_6492);
and U10140 (N_10140,N_7730,N_8896);
and U10141 (N_10141,N_6109,N_6742);
or U10142 (N_10142,N_6802,N_6735);
nand U10143 (N_10143,N_8115,N_6878);
nor U10144 (N_10144,N_6810,N_6503);
nor U10145 (N_10145,N_6416,N_6776);
or U10146 (N_10146,N_6111,N_7029);
nor U10147 (N_10147,N_8810,N_6210);
nand U10148 (N_10148,N_7101,N_6950);
nand U10149 (N_10149,N_6187,N_7497);
or U10150 (N_10150,N_7577,N_7130);
or U10151 (N_10151,N_6749,N_6297);
and U10152 (N_10152,N_6830,N_7172);
xnor U10153 (N_10153,N_8453,N_7124);
nand U10154 (N_10154,N_7969,N_7541);
nand U10155 (N_10155,N_8809,N_6284);
nor U10156 (N_10156,N_6016,N_6363);
nand U10157 (N_10157,N_6677,N_8306);
and U10158 (N_10158,N_7367,N_7952);
nor U10159 (N_10159,N_6281,N_8438);
or U10160 (N_10160,N_6729,N_7147);
or U10161 (N_10161,N_8820,N_7466);
nand U10162 (N_10162,N_8852,N_8978);
nor U10163 (N_10163,N_6365,N_6936);
xor U10164 (N_10164,N_6911,N_8413);
nand U10165 (N_10165,N_6409,N_6276);
xor U10166 (N_10166,N_6176,N_7447);
nor U10167 (N_10167,N_6178,N_6607);
and U10168 (N_10168,N_8298,N_6424);
or U10169 (N_10169,N_6455,N_7018);
and U10170 (N_10170,N_8007,N_8350);
or U10171 (N_10171,N_7488,N_8948);
and U10172 (N_10172,N_8358,N_8732);
nand U10173 (N_10173,N_6375,N_8925);
or U10174 (N_10174,N_7180,N_7614);
and U10175 (N_10175,N_6355,N_8845);
nand U10176 (N_10176,N_7208,N_6385);
nand U10177 (N_10177,N_7385,N_8042);
nand U10178 (N_10178,N_8394,N_7951);
and U10179 (N_10179,N_7821,N_6447);
and U10180 (N_10180,N_7642,N_7539);
or U10181 (N_10181,N_8497,N_6549);
or U10182 (N_10182,N_8290,N_8932);
or U10183 (N_10183,N_6763,N_7574);
nor U10184 (N_10184,N_8116,N_7404);
or U10185 (N_10185,N_6219,N_6865);
and U10186 (N_10186,N_7203,N_8590);
and U10187 (N_10187,N_7977,N_7612);
or U10188 (N_10188,N_7650,N_7387);
and U10189 (N_10189,N_8593,N_8427);
or U10190 (N_10190,N_7760,N_7239);
or U10191 (N_10191,N_8180,N_6971);
and U10192 (N_10192,N_7800,N_8024);
or U10193 (N_10193,N_7009,N_6260);
xnor U10194 (N_10194,N_6237,N_7296);
nand U10195 (N_10195,N_8592,N_8616);
or U10196 (N_10196,N_8043,N_8324);
nand U10197 (N_10197,N_7361,N_8142);
nand U10198 (N_10198,N_7648,N_8817);
nor U10199 (N_10199,N_6026,N_8215);
nor U10200 (N_10200,N_7515,N_8550);
and U10201 (N_10201,N_6565,N_8284);
nand U10202 (N_10202,N_8219,N_6223);
nor U10203 (N_10203,N_8816,N_8954);
and U10204 (N_10204,N_7684,N_7635);
and U10205 (N_10205,N_7696,N_7421);
nor U10206 (N_10206,N_7576,N_6003);
and U10207 (N_10207,N_8507,N_6955);
nor U10208 (N_10208,N_7097,N_8909);
and U10209 (N_10209,N_6900,N_6934);
nor U10210 (N_10210,N_8330,N_8871);
and U10211 (N_10211,N_7086,N_6475);
or U10212 (N_10212,N_8104,N_6723);
xor U10213 (N_10213,N_8629,N_6347);
and U10214 (N_10214,N_8423,N_8953);
and U10215 (N_10215,N_8486,N_7854);
nor U10216 (N_10216,N_7702,N_7759);
and U10217 (N_10217,N_7805,N_6200);
nand U10218 (N_10218,N_8605,N_7532);
nor U10219 (N_10219,N_7852,N_7428);
nor U10220 (N_10220,N_8393,N_6147);
or U10221 (N_10221,N_8768,N_6304);
nand U10222 (N_10222,N_8295,N_8513);
nand U10223 (N_10223,N_8068,N_6361);
or U10224 (N_10224,N_6317,N_7818);
nor U10225 (N_10225,N_8681,N_8811);
nand U10226 (N_10226,N_8125,N_7625);
and U10227 (N_10227,N_7005,N_7862);
or U10228 (N_10228,N_7677,N_7955);
nor U10229 (N_10229,N_8884,N_7893);
nor U10230 (N_10230,N_7139,N_7426);
nor U10231 (N_10231,N_6144,N_7394);
and U10232 (N_10232,N_7025,N_6879);
or U10233 (N_10233,N_7984,N_8442);
nor U10234 (N_10234,N_8269,N_6048);
nand U10235 (N_10235,N_7879,N_7380);
or U10236 (N_10236,N_7508,N_6635);
and U10237 (N_10237,N_7809,N_6887);
nand U10238 (N_10238,N_7449,N_8666);
nor U10239 (N_10239,N_7448,N_6032);
nand U10240 (N_10240,N_7383,N_8070);
nand U10241 (N_10241,N_6229,N_7292);
and U10242 (N_10242,N_6263,N_7504);
and U10243 (N_10243,N_8204,N_6523);
nand U10244 (N_10244,N_8783,N_6448);
nor U10245 (N_10245,N_7377,N_6106);
nand U10246 (N_10246,N_8512,N_7483);
nand U10247 (N_10247,N_6541,N_8448);
and U10248 (N_10248,N_6962,N_7531);
and U10249 (N_10249,N_6632,N_7062);
or U10250 (N_10250,N_8348,N_8889);
and U10251 (N_10251,N_6748,N_6468);
and U10252 (N_10252,N_8320,N_8761);
or U10253 (N_10253,N_6352,N_7706);
and U10254 (N_10254,N_7826,N_6088);
and U10255 (N_10255,N_7146,N_8703);
nor U10256 (N_10256,N_7500,N_8555);
or U10257 (N_10257,N_8821,N_6021);
and U10258 (N_10258,N_6278,N_6194);
and U10259 (N_10259,N_8351,N_7002);
or U10260 (N_10260,N_6922,N_8837);
and U10261 (N_10261,N_6556,N_7798);
nand U10262 (N_10262,N_8119,N_6838);
nand U10263 (N_10263,N_6518,N_8994);
nor U10264 (N_10264,N_6555,N_7055);
and U10265 (N_10265,N_7919,N_7511);
and U10266 (N_10266,N_8991,N_8847);
or U10267 (N_10267,N_8614,N_7892);
nand U10268 (N_10268,N_8876,N_6214);
nor U10269 (N_10269,N_6324,N_6769);
and U10270 (N_10270,N_6459,N_8166);
and U10271 (N_10271,N_8604,N_6668);
and U10272 (N_10272,N_6680,N_6135);
nor U10273 (N_10273,N_8231,N_6873);
xnor U10274 (N_10274,N_8264,N_6801);
nor U10275 (N_10275,N_8936,N_8674);
or U10276 (N_10276,N_6073,N_6325);
nor U10277 (N_10277,N_6768,N_7540);
and U10278 (N_10278,N_6477,N_6221);
nand U10279 (N_10279,N_8814,N_8870);
nand U10280 (N_10280,N_7143,N_8193);
and U10281 (N_10281,N_6241,N_7510);
nor U10282 (N_10282,N_7218,N_8935);
nand U10283 (N_10283,N_7442,N_7082);
and U10284 (N_10284,N_6818,N_7063);
or U10285 (N_10285,N_6969,N_7543);
and U10286 (N_10286,N_6314,N_8080);
nand U10287 (N_10287,N_6620,N_8638);
nor U10288 (N_10288,N_7245,N_8682);
nor U10289 (N_10289,N_8828,N_8415);
nor U10290 (N_10290,N_6122,N_6892);
nand U10291 (N_10291,N_6711,N_8668);
nor U10292 (N_10292,N_7337,N_6411);
or U10293 (N_10293,N_7536,N_8067);
or U10294 (N_10294,N_8354,N_6145);
and U10295 (N_10295,N_8462,N_8999);
and U10296 (N_10296,N_7115,N_7158);
nor U10297 (N_10297,N_7386,N_8039);
nor U10298 (N_10298,N_7575,N_6076);
and U10299 (N_10299,N_6174,N_8758);
nor U10300 (N_10300,N_6667,N_8374);
and U10301 (N_10301,N_8087,N_8230);
nor U10302 (N_10302,N_6158,N_8915);
nand U10303 (N_10303,N_8186,N_7334);
or U10304 (N_10304,N_8612,N_7213);
and U10305 (N_10305,N_8993,N_7948);
or U10306 (N_10306,N_7100,N_8780);
nor U10307 (N_10307,N_7996,N_6367);
or U10308 (N_10308,N_8867,N_6244);
nand U10309 (N_10309,N_6893,N_6506);
or U10310 (N_10310,N_7127,N_8008);
nor U10311 (N_10311,N_7451,N_7878);
nor U10312 (N_10312,N_6078,N_6577);
and U10313 (N_10313,N_8645,N_7065);
and U10314 (N_10314,N_7429,N_8880);
and U10315 (N_10315,N_7703,N_8559);
or U10316 (N_10316,N_7830,N_8784);
or U10317 (N_10317,N_6699,N_6752);
nor U10318 (N_10318,N_7754,N_6642);
and U10319 (N_10319,N_8263,N_6439);
or U10320 (N_10320,N_7228,N_6927);
nor U10321 (N_10321,N_6995,N_8895);
and U10322 (N_10322,N_6240,N_7093);
and U10323 (N_10323,N_7768,N_8981);
or U10324 (N_10324,N_7750,N_8937);
xnor U10325 (N_10325,N_6004,N_6435);
nor U10326 (N_10326,N_7145,N_6121);
or U10327 (N_10327,N_7332,N_6821);
nor U10328 (N_10328,N_6402,N_6446);
or U10329 (N_10329,N_8029,N_6480);
nor U10330 (N_10330,N_8272,N_6279);
or U10331 (N_10331,N_6745,N_8990);
nor U10332 (N_10332,N_8888,N_6759);
nand U10333 (N_10333,N_7247,N_6553);
nand U10334 (N_10334,N_6412,N_7214);
nand U10335 (N_10335,N_8959,N_8006);
and U10336 (N_10336,N_7138,N_7621);
or U10337 (N_10337,N_7452,N_6856);
and U10338 (N_10338,N_6674,N_8963);
xor U10339 (N_10339,N_7433,N_7134);
nand U10340 (N_10340,N_7156,N_7925);
or U10341 (N_10341,N_7617,N_6876);
nand U10342 (N_10342,N_8499,N_7823);
or U10343 (N_10343,N_8258,N_8749);
nor U10344 (N_10344,N_6463,N_6081);
nand U10345 (N_10345,N_6869,N_6817);
and U10346 (N_10346,N_8237,N_6018);
and U10347 (N_10347,N_8208,N_8293);
nand U10348 (N_10348,N_6285,N_8175);
nor U10349 (N_10349,N_8379,N_8174);
nand U10350 (N_10350,N_6172,N_8205);
nand U10351 (N_10351,N_7402,N_7870);
xnor U10352 (N_10352,N_8979,N_6153);
or U10353 (N_10353,N_8518,N_7707);
and U10354 (N_10354,N_6529,N_8799);
or U10355 (N_10355,N_8648,N_8726);
and U10356 (N_10356,N_7963,N_6649);
nor U10357 (N_10357,N_7813,N_8549);
and U10358 (N_10358,N_8207,N_6813);
or U10359 (N_10359,N_7726,N_6013);
nand U10360 (N_10360,N_6326,N_7516);
nor U10361 (N_10361,N_6338,N_7546);
nor U10362 (N_10362,N_7571,N_6014);
nor U10363 (N_10363,N_7840,N_6790);
nand U10364 (N_10364,N_7422,N_6755);
xnor U10365 (N_10365,N_7851,N_8034);
or U10366 (N_10366,N_7259,N_6379);
nor U10367 (N_10367,N_6782,N_8906);
or U10368 (N_10368,N_8238,N_7033);
or U10369 (N_10369,N_7687,N_7692);
nor U10370 (N_10370,N_7232,N_8476);
or U10371 (N_10371,N_8646,N_8118);
nand U10372 (N_10372,N_6092,N_7330);
nand U10373 (N_10373,N_6587,N_6792);
and U10374 (N_10374,N_8760,N_8757);
and U10375 (N_10375,N_6836,N_6345);
and U10376 (N_10376,N_7611,N_8481);
or U10377 (N_10377,N_8942,N_7552);
nand U10378 (N_10378,N_6298,N_6656);
and U10379 (N_10379,N_8056,N_6353);
nor U10380 (N_10380,N_6227,N_8804);
nor U10381 (N_10381,N_7026,N_6783);
and U10382 (N_10382,N_6183,N_6636);
nand U10383 (N_10383,N_6704,N_7326);
and U10384 (N_10384,N_7160,N_8233);
and U10385 (N_10385,N_8903,N_7907);
nor U10386 (N_10386,N_8482,N_8913);
or U10387 (N_10387,N_8567,N_8074);
or U10388 (N_10388,N_8772,N_7255);
nand U10389 (N_10389,N_7275,N_6082);
nand U10390 (N_10390,N_8714,N_8023);
or U10391 (N_10391,N_7230,N_7589);
and U10392 (N_10392,N_6349,N_8776);
or U10393 (N_10393,N_7624,N_8072);
or U10394 (N_10394,N_8467,N_8628);
and U10395 (N_10395,N_6331,N_6428);
and U10396 (N_10396,N_6994,N_8052);
nor U10397 (N_10397,N_6937,N_6358);
nand U10398 (N_10398,N_7961,N_8545);
and U10399 (N_10399,N_7545,N_7815);
and U10400 (N_10400,N_8824,N_7418);
nor U10401 (N_10401,N_8831,N_8660);
nor U10402 (N_10402,N_8316,N_6201);
or U10403 (N_10403,N_7811,N_7905);
nand U10404 (N_10404,N_6591,N_7564);
xor U10405 (N_10405,N_7507,N_6960);
or U10406 (N_10406,N_8988,N_6213);
and U10407 (N_10407,N_8099,N_8652);
and U10408 (N_10408,N_6493,N_8392);
and U10409 (N_10409,N_7534,N_6165);
or U10410 (N_10410,N_7192,N_7327);
nand U10411 (N_10411,N_8792,N_7795);
or U10412 (N_10412,N_6530,N_8235);
or U10413 (N_10413,N_6351,N_7639);
nand U10414 (N_10414,N_6057,N_7017);
xor U10415 (N_10415,N_7338,N_7986);
or U10416 (N_10416,N_6513,N_8151);
or U10417 (N_10417,N_8686,N_7727);
xnor U10418 (N_10418,N_8548,N_8601);
nor U10419 (N_10419,N_7369,N_8609);
nor U10420 (N_10420,N_8740,N_8030);
nand U10421 (N_10421,N_7474,N_6664);
and U10422 (N_10422,N_8516,N_7081);
nor U10423 (N_10423,N_7094,N_6368);
nand U10424 (N_10424,N_7599,N_8251);
xor U10425 (N_10425,N_6840,N_7140);
nor U10426 (N_10426,N_6967,N_6826);
and U10427 (N_10427,N_8676,N_6731);
xnor U10428 (N_10428,N_7163,N_7430);
nand U10429 (N_10429,N_8385,N_8926);
nor U10430 (N_10430,N_6785,N_7423);
nand U10431 (N_10431,N_6064,N_8227);
or U10432 (N_10432,N_8164,N_8459);
or U10433 (N_10433,N_6957,N_7345);
nor U10434 (N_10434,N_7219,N_8577);
and U10435 (N_10435,N_8844,N_6303);
and U10436 (N_10436,N_7439,N_8079);
and U10437 (N_10437,N_8288,N_7136);
and U10438 (N_10438,N_7491,N_6965);
or U10439 (N_10439,N_8465,N_7544);
or U10440 (N_10440,N_7401,N_8162);
xor U10441 (N_10441,N_6232,N_7700);
and U10442 (N_10442,N_6400,N_7568);
nor U10443 (N_10443,N_6909,N_8361);
nor U10444 (N_10444,N_7864,N_8611);
nor U10445 (N_10445,N_8038,N_6652);
and U10446 (N_10446,N_8097,N_8098);
and U10447 (N_10447,N_6903,N_7669);
nand U10448 (N_10448,N_8291,N_7814);
or U10449 (N_10449,N_7812,N_8791);
or U10450 (N_10450,N_6451,N_6947);
xor U10451 (N_10451,N_6327,N_8020);
nor U10452 (N_10452,N_7927,N_6941);
nand U10453 (N_10453,N_7349,N_6483);
and U10454 (N_10454,N_8134,N_7829);
nand U10455 (N_10455,N_7757,N_7111);
nor U10456 (N_10456,N_7392,N_8405);
and U10457 (N_10457,N_6054,N_6815);
and U10458 (N_10458,N_6932,N_8866);
and U10459 (N_10459,N_6312,N_7945);
nand U10460 (N_10460,N_7972,N_7939);
and U10461 (N_10461,N_6436,N_7010);
or U10462 (N_10462,N_8014,N_7074);
nor U10463 (N_10463,N_7043,N_7482);
nor U10464 (N_10464,N_6502,N_8536);
nor U10465 (N_10465,N_6528,N_8773);
nand U10466 (N_10466,N_8191,N_6034);
or U10467 (N_10467,N_7618,N_7087);
and U10468 (N_10468,N_6143,N_8843);
nand U10469 (N_10469,N_6035,N_8277);
nor U10470 (N_10470,N_7861,N_7769);
nand U10471 (N_10471,N_6522,N_7845);
nor U10472 (N_10472,N_6561,N_7071);
nor U10473 (N_10473,N_7782,N_7485);
nor U10474 (N_10474,N_6077,N_6920);
and U10475 (N_10475,N_6935,N_8793);
or U10476 (N_10476,N_8900,N_7911);
nand U10477 (N_10477,N_7196,N_7038);
xor U10478 (N_10478,N_8223,N_8642);
or U10479 (N_10479,N_7084,N_7869);
nor U10480 (N_10480,N_7391,N_6315);
or U10481 (N_10481,N_7182,N_7596);
or U10482 (N_10482,N_7783,N_7032);
or U10483 (N_10483,N_8873,N_6293);
xor U10484 (N_10484,N_6786,N_6595);
nor U10485 (N_10485,N_8307,N_7920);
nand U10486 (N_10486,N_8912,N_8276);
and U10487 (N_10487,N_6520,N_7505);
and U10488 (N_10488,N_6141,N_8597);
and U10489 (N_10489,N_8435,N_7844);
nand U10490 (N_10490,N_8289,N_7834);
xor U10491 (N_10491,N_6302,N_8940);
and U10492 (N_10492,N_8826,N_7940);
nand U10493 (N_10493,N_8635,N_7711);
nand U10494 (N_10494,N_8282,N_7080);
nor U10495 (N_10495,N_8875,N_6192);
nor U10496 (N_10496,N_8987,N_7298);
nor U10497 (N_10497,N_7926,N_6622);
nand U10498 (N_10498,N_7890,N_6198);
nand U10499 (N_10499,N_6469,N_7674);
and U10500 (N_10500,N_7923,N_7071);
nand U10501 (N_10501,N_6785,N_6482);
and U10502 (N_10502,N_8176,N_6470);
nand U10503 (N_10503,N_8061,N_6279);
nand U10504 (N_10504,N_7783,N_8220);
and U10505 (N_10505,N_7148,N_8430);
nand U10506 (N_10506,N_8686,N_8465);
or U10507 (N_10507,N_8395,N_7480);
and U10508 (N_10508,N_8040,N_6552);
or U10509 (N_10509,N_8785,N_6932);
nor U10510 (N_10510,N_8696,N_6151);
xor U10511 (N_10511,N_7103,N_7206);
nand U10512 (N_10512,N_8530,N_8057);
nor U10513 (N_10513,N_6550,N_6502);
or U10514 (N_10514,N_8522,N_8108);
or U10515 (N_10515,N_6745,N_8856);
or U10516 (N_10516,N_7746,N_7476);
nor U10517 (N_10517,N_8213,N_6162);
nor U10518 (N_10518,N_8139,N_8904);
or U10519 (N_10519,N_6918,N_8394);
nand U10520 (N_10520,N_6213,N_6361);
nand U10521 (N_10521,N_8832,N_7035);
nor U10522 (N_10522,N_6040,N_7114);
or U10523 (N_10523,N_7437,N_7802);
nor U10524 (N_10524,N_8916,N_7232);
nand U10525 (N_10525,N_6967,N_8122);
xnor U10526 (N_10526,N_8207,N_6215);
or U10527 (N_10527,N_8019,N_7201);
and U10528 (N_10528,N_7899,N_8469);
or U10529 (N_10529,N_8574,N_7202);
nor U10530 (N_10530,N_7995,N_7918);
nor U10531 (N_10531,N_8401,N_8056);
nand U10532 (N_10532,N_6643,N_6744);
nand U10533 (N_10533,N_6886,N_6461);
and U10534 (N_10534,N_6742,N_6091);
nor U10535 (N_10535,N_8916,N_8000);
or U10536 (N_10536,N_7250,N_7567);
or U10537 (N_10537,N_6626,N_6917);
and U10538 (N_10538,N_8059,N_6817);
and U10539 (N_10539,N_7174,N_6774);
nand U10540 (N_10540,N_6584,N_7738);
nand U10541 (N_10541,N_6490,N_6093);
and U10542 (N_10542,N_6675,N_8836);
nand U10543 (N_10543,N_8695,N_6052);
nor U10544 (N_10544,N_7296,N_6251);
or U10545 (N_10545,N_8476,N_7632);
and U10546 (N_10546,N_6692,N_8613);
nand U10547 (N_10547,N_7777,N_8304);
and U10548 (N_10548,N_7575,N_8712);
nor U10549 (N_10549,N_8471,N_7476);
and U10550 (N_10550,N_8352,N_7045);
or U10551 (N_10551,N_6712,N_6889);
nand U10552 (N_10552,N_8867,N_6087);
and U10553 (N_10553,N_7716,N_8556);
and U10554 (N_10554,N_7690,N_7723);
and U10555 (N_10555,N_6669,N_6856);
nand U10556 (N_10556,N_7250,N_7115);
or U10557 (N_10557,N_8527,N_6517);
or U10558 (N_10558,N_7340,N_8007);
nor U10559 (N_10559,N_6027,N_8445);
nor U10560 (N_10560,N_8850,N_8743);
nand U10561 (N_10561,N_8108,N_7762);
and U10562 (N_10562,N_8867,N_8510);
nand U10563 (N_10563,N_7638,N_8872);
and U10564 (N_10564,N_7303,N_6168);
or U10565 (N_10565,N_8676,N_6751);
and U10566 (N_10566,N_6987,N_6428);
and U10567 (N_10567,N_8161,N_8276);
nor U10568 (N_10568,N_6863,N_6641);
or U10569 (N_10569,N_6825,N_8699);
nor U10570 (N_10570,N_8934,N_6583);
nor U10571 (N_10571,N_6981,N_8460);
or U10572 (N_10572,N_6489,N_6217);
nand U10573 (N_10573,N_8896,N_6373);
nor U10574 (N_10574,N_8136,N_7855);
nor U10575 (N_10575,N_6459,N_6208);
and U10576 (N_10576,N_7774,N_7061);
nand U10577 (N_10577,N_6814,N_7060);
or U10578 (N_10578,N_8308,N_7319);
nand U10579 (N_10579,N_6650,N_6065);
xor U10580 (N_10580,N_8470,N_6739);
nand U10581 (N_10581,N_7682,N_8766);
and U10582 (N_10582,N_8914,N_6016);
and U10583 (N_10583,N_6473,N_8096);
nor U10584 (N_10584,N_8023,N_8197);
xor U10585 (N_10585,N_6025,N_7354);
or U10586 (N_10586,N_6700,N_8777);
and U10587 (N_10587,N_6015,N_7684);
nand U10588 (N_10588,N_6688,N_8299);
nand U10589 (N_10589,N_8653,N_8752);
nor U10590 (N_10590,N_7909,N_6925);
nand U10591 (N_10591,N_7596,N_8353);
or U10592 (N_10592,N_8010,N_7447);
or U10593 (N_10593,N_8884,N_6815);
or U10594 (N_10594,N_8690,N_7210);
nor U10595 (N_10595,N_7316,N_8323);
nor U10596 (N_10596,N_6943,N_8475);
and U10597 (N_10597,N_7528,N_6761);
and U10598 (N_10598,N_8937,N_8191);
xor U10599 (N_10599,N_7388,N_7400);
nand U10600 (N_10600,N_6171,N_8705);
nor U10601 (N_10601,N_7593,N_7290);
or U10602 (N_10602,N_8040,N_6611);
or U10603 (N_10603,N_8440,N_7228);
nor U10604 (N_10604,N_8213,N_7675);
or U10605 (N_10605,N_7371,N_8711);
nand U10606 (N_10606,N_6215,N_7866);
nand U10607 (N_10607,N_6940,N_7438);
or U10608 (N_10608,N_6881,N_6102);
nor U10609 (N_10609,N_6821,N_6398);
and U10610 (N_10610,N_8692,N_6152);
nor U10611 (N_10611,N_7642,N_8443);
nor U10612 (N_10612,N_6015,N_6653);
nor U10613 (N_10613,N_7983,N_8093);
nand U10614 (N_10614,N_7563,N_6494);
or U10615 (N_10615,N_6007,N_8580);
nor U10616 (N_10616,N_8352,N_8108);
and U10617 (N_10617,N_8577,N_7187);
and U10618 (N_10618,N_7935,N_6159);
xnor U10619 (N_10619,N_8593,N_7457);
nand U10620 (N_10620,N_8782,N_6342);
nor U10621 (N_10621,N_8623,N_8785);
nor U10622 (N_10622,N_6672,N_8074);
nor U10623 (N_10623,N_7453,N_8336);
nor U10624 (N_10624,N_8733,N_6775);
nand U10625 (N_10625,N_8746,N_7849);
or U10626 (N_10626,N_7486,N_8934);
xor U10627 (N_10627,N_6110,N_8132);
nand U10628 (N_10628,N_6136,N_7108);
and U10629 (N_10629,N_7444,N_6737);
and U10630 (N_10630,N_8100,N_8826);
or U10631 (N_10631,N_8194,N_6204);
and U10632 (N_10632,N_6614,N_8845);
and U10633 (N_10633,N_7133,N_7176);
or U10634 (N_10634,N_8622,N_8005);
nand U10635 (N_10635,N_6579,N_6182);
or U10636 (N_10636,N_7077,N_8857);
and U10637 (N_10637,N_6225,N_6556);
and U10638 (N_10638,N_6963,N_6789);
nand U10639 (N_10639,N_7657,N_8183);
nor U10640 (N_10640,N_6888,N_7740);
or U10641 (N_10641,N_7912,N_6398);
nand U10642 (N_10642,N_8581,N_7834);
and U10643 (N_10643,N_7986,N_6266);
or U10644 (N_10644,N_6709,N_8810);
nand U10645 (N_10645,N_6954,N_8777);
or U10646 (N_10646,N_6482,N_7103);
nand U10647 (N_10647,N_7698,N_7177);
nand U10648 (N_10648,N_8878,N_8903);
or U10649 (N_10649,N_8541,N_6765);
or U10650 (N_10650,N_7200,N_6651);
nor U10651 (N_10651,N_6975,N_6816);
and U10652 (N_10652,N_6890,N_6837);
or U10653 (N_10653,N_7102,N_7849);
and U10654 (N_10654,N_7380,N_8384);
or U10655 (N_10655,N_8926,N_7911);
or U10656 (N_10656,N_7803,N_6360);
nor U10657 (N_10657,N_6463,N_8319);
nor U10658 (N_10658,N_6328,N_7176);
nand U10659 (N_10659,N_6749,N_7327);
or U10660 (N_10660,N_8458,N_7782);
nand U10661 (N_10661,N_8485,N_8597);
and U10662 (N_10662,N_7586,N_8884);
or U10663 (N_10663,N_8497,N_6419);
nand U10664 (N_10664,N_6414,N_8477);
nor U10665 (N_10665,N_8260,N_6854);
or U10666 (N_10666,N_6374,N_6667);
and U10667 (N_10667,N_8620,N_7177);
or U10668 (N_10668,N_7578,N_8917);
nor U10669 (N_10669,N_6869,N_6902);
nor U10670 (N_10670,N_6876,N_7533);
and U10671 (N_10671,N_7197,N_8901);
nand U10672 (N_10672,N_6218,N_6883);
nor U10673 (N_10673,N_8769,N_7010);
and U10674 (N_10674,N_6934,N_6300);
or U10675 (N_10675,N_7672,N_7642);
and U10676 (N_10676,N_7474,N_6152);
nor U10677 (N_10677,N_8545,N_6053);
and U10678 (N_10678,N_6378,N_7219);
and U10679 (N_10679,N_7069,N_7946);
or U10680 (N_10680,N_7772,N_6406);
nor U10681 (N_10681,N_7363,N_7063);
or U10682 (N_10682,N_7066,N_6938);
nand U10683 (N_10683,N_6538,N_8563);
nor U10684 (N_10684,N_8947,N_8388);
nor U10685 (N_10685,N_8335,N_7468);
and U10686 (N_10686,N_7678,N_6746);
and U10687 (N_10687,N_7524,N_7789);
nor U10688 (N_10688,N_7538,N_6065);
or U10689 (N_10689,N_6406,N_8570);
and U10690 (N_10690,N_7561,N_6468);
nand U10691 (N_10691,N_6569,N_7817);
or U10692 (N_10692,N_8615,N_6966);
nor U10693 (N_10693,N_6411,N_7202);
nand U10694 (N_10694,N_7574,N_6035);
nand U10695 (N_10695,N_8454,N_8609);
nand U10696 (N_10696,N_7427,N_7978);
nor U10697 (N_10697,N_7562,N_6187);
nor U10698 (N_10698,N_8086,N_7231);
or U10699 (N_10699,N_7883,N_6964);
nor U10700 (N_10700,N_8713,N_6668);
nand U10701 (N_10701,N_8155,N_6522);
nand U10702 (N_10702,N_8695,N_6135);
nand U10703 (N_10703,N_7956,N_7753);
and U10704 (N_10704,N_8781,N_8276);
and U10705 (N_10705,N_8648,N_8677);
and U10706 (N_10706,N_6577,N_6375);
nand U10707 (N_10707,N_7002,N_8130);
nor U10708 (N_10708,N_8594,N_8981);
nor U10709 (N_10709,N_6022,N_6950);
or U10710 (N_10710,N_8842,N_6874);
or U10711 (N_10711,N_7264,N_8916);
and U10712 (N_10712,N_6932,N_6265);
nor U10713 (N_10713,N_7565,N_6005);
nand U10714 (N_10714,N_6310,N_8853);
nand U10715 (N_10715,N_7217,N_7554);
and U10716 (N_10716,N_8512,N_7959);
or U10717 (N_10717,N_7321,N_7983);
or U10718 (N_10718,N_8665,N_8832);
nand U10719 (N_10719,N_7653,N_6373);
and U10720 (N_10720,N_6069,N_6611);
nor U10721 (N_10721,N_6913,N_7633);
nor U10722 (N_10722,N_7351,N_8198);
nand U10723 (N_10723,N_7891,N_7465);
nor U10724 (N_10724,N_8873,N_8980);
nor U10725 (N_10725,N_8706,N_7197);
and U10726 (N_10726,N_8001,N_7265);
nor U10727 (N_10727,N_6559,N_8809);
or U10728 (N_10728,N_6213,N_8952);
and U10729 (N_10729,N_7122,N_7170);
nor U10730 (N_10730,N_8052,N_8764);
nor U10731 (N_10731,N_6320,N_7098);
or U10732 (N_10732,N_6599,N_6075);
or U10733 (N_10733,N_6779,N_8840);
nand U10734 (N_10734,N_6018,N_7021);
or U10735 (N_10735,N_7662,N_6343);
or U10736 (N_10736,N_8871,N_7055);
and U10737 (N_10737,N_7297,N_8051);
or U10738 (N_10738,N_6252,N_8604);
or U10739 (N_10739,N_8002,N_7997);
nand U10740 (N_10740,N_7078,N_6705);
or U10741 (N_10741,N_7827,N_8634);
or U10742 (N_10742,N_8445,N_8924);
nand U10743 (N_10743,N_8626,N_6611);
or U10744 (N_10744,N_8462,N_8891);
nor U10745 (N_10745,N_8812,N_6081);
or U10746 (N_10746,N_7968,N_7800);
or U10747 (N_10747,N_7076,N_6053);
and U10748 (N_10748,N_8518,N_6209);
and U10749 (N_10749,N_6875,N_7376);
or U10750 (N_10750,N_8125,N_7182);
nand U10751 (N_10751,N_8787,N_6403);
xor U10752 (N_10752,N_6342,N_6140);
or U10753 (N_10753,N_7685,N_8238);
and U10754 (N_10754,N_7076,N_8493);
nand U10755 (N_10755,N_6104,N_6049);
nor U10756 (N_10756,N_6935,N_6650);
or U10757 (N_10757,N_6710,N_8353);
nor U10758 (N_10758,N_8425,N_6521);
or U10759 (N_10759,N_7969,N_6541);
or U10760 (N_10760,N_7150,N_7257);
and U10761 (N_10761,N_7964,N_6219);
or U10762 (N_10762,N_8529,N_6164);
and U10763 (N_10763,N_6184,N_7481);
or U10764 (N_10764,N_8962,N_8705);
nor U10765 (N_10765,N_6932,N_7233);
nand U10766 (N_10766,N_7499,N_8547);
nor U10767 (N_10767,N_6353,N_8921);
nand U10768 (N_10768,N_8120,N_6465);
nand U10769 (N_10769,N_7320,N_8692);
xnor U10770 (N_10770,N_6686,N_8583);
nor U10771 (N_10771,N_7439,N_6364);
or U10772 (N_10772,N_6948,N_8348);
or U10773 (N_10773,N_7265,N_8360);
nor U10774 (N_10774,N_8904,N_8574);
nor U10775 (N_10775,N_7967,N_7995);
nor U10776 (N_10776,N_8450,N_8036);
and U10777 (N_10777,N_8587,N_7174);
nor U10778 (N_10778,N_6017,N_8813);
and U10779 (N_10779,N_6851,N_6754);
xor U10780 (N_10780,N_8971,N_8549);
nor U10781 (N_10781,N_7391,N_7547);
and U10782 (N_10782,N_6588,N_8368);
nand U10783 (N_10783,N_6269,N_8482);
and U10784 (N_10784,N_8297,N_6337);
or U10785 (N_10785,N_8191,N_6563);
nand U10786 (N_10786,N_7328,N_7675);
or U10787 (N_10787,N_7495,N_7015);
or U10788 (N_10788,N_7314,N_7018);
nand U10789 (N_10789,N_6802,N_6221);
and U10790 (N_10790,N_8865,N_8051);
nand U10791 (N_10791,N_8051,N_6217);
nor U10792 (N_10792,N_7314,N_8641);
and U10793 (N_10793,N_8419,N_6162);
nor U10794 (N_10794,N_6772,N_8591);
and U10795 (N_10795,N_8533,N_7448);
nand U10796 (N_10796,N_7606,N_8490);
or U10797 (N_10797,N_6387,N_7605);
nand U10798 (N_10798,N_6989,N_8049);
nor U10799 (N_10799,N_7999,N_7695);
nor U10800 (N_10800,N_7983,N_7904);
and U10801 (N_10801,N_8586,N_6163);
or U10802 (N_10802,N_6341,N_8080);
or U10803 (N_10803,N_8260,N_7116);
or U10804 (N_10804,N_7985,N_6575);
nor U10805 (N_10805,N_6250,N_8737);
and U10806 (N_10806,N_7166,N_7328);
or U10807 (N_10807,N_7593,N_7051);
or U10808 (N_10808,N_7115,N_8385);
xor U10809 (N_10809,N_7029,N_7701);
nor U10810 (N_10810,N_6377,N_8004);
nor U10811 (N_10811,N_7018,N_7764);
xor U10812 (N_10812,N_6745,N_7406);
nand U10813 (N_10813,N_8694,N_8893);
nor U10814 (N_10814,N_7867,N_6534);
and U10815 (N_10815,N_6701,N_8714);
nor U10816 (N_10816,N_8345,N_8967);
nand U10817 (N_10817,N_7400,N_7047);
and U10818 (N_10818,N_6170,N_7829);
nor U10819 (N_10819,N_8143,N_8447);
or U10820 (N_10820,N_7865,N_6928);
or U10821 (N_10821,N_6534,N_6773);
nor U10822 (N_10822,N_7255,N_7522);
nor U10823 (N_10823,N_8901,N_6075);
and U10824 (N_10824,N_6853,N_8554);
nand U10825 (N_10825,N_8619,N_7191);
nand U10826 (N_10826,N_8090,N_6709);
nor U10827 (N_10827,N_6058,N_8188);
nor U10828 (N_10828,N_8679,N_8524);
or U10829 (N_10829,N_8544,N_7065);
and U10830 (N_10830,N_8924,N_8717);
or U10831 (N_10831,N_6223,N_8143);
nand U10832 (N_10832,N_7237,N_8137);
nor U10833 (N_10833,N_7550,N_6550);
and U10834 (N_10834,N_6856,N_6582);
nor U10835 (N_10835,N_6932,N_6621);
or U10836 (N_10836,N_6237,N_6977);
and U10837 (N_10837,N_7662,N_7684);
and U10838 (N_10838,N_6146,N_7074);
or U10839 (N_10839,N_7906,N_6230);
and U10840 (N_10840,N_8521,N_7495);
nor U10841 (N_10841,N_6967,N_7311);
nor U10842 (N_10842,N_7953,N_7091);
and U10843 (N_10843,N_8918,N_6391);
and U10844 (N_10844,N_6430,N_7125);
nor U10845 (N_10845,N_6946,N_8910);
or U10846 (N_10846,N_8805,N_6189);
or U10847 (N_10847,N_6141,N_6159);
and U10848 (N_10848,N_8200,N_7968);
nor U10849 (N_10849,N_6625,N_7394);
nor U10850 (N_10850,N_6766,N_7478);
nand U10851 (N_10851,N_7700,N_8774);
and U10852 (N_10852,N_8064,N_8022);
nor U10853 (N_10853,N_7534,N_7873);
nor U10854 (N_10854,N_6740,N_8315);
or U10855 (N_10855,N_7768,N_6367);
or U10856 (N_10856,N_8943,N_6752);
or U10857 (N_10857,N_7744,N_6937);
or U10858 (N_10858,N_8068,N_8168);
or U10859 (N_10859,N_8543,N_6253);
and U10860 (N_10860,N_7661,N_7433);
and U10861 (N_10861,N_7282,N_7860);
nor U10862 (N_10862,N_6380,N_7757);
nand U10863 (N_10863,N_8685,N_8047);
and U10864 (N_10864,N_7891,N_7112);
nand U10865 (N_10865,N_8515,N_7363);
nor U10866 (N_10866,N_7924,N_8336);
or U10867 (N_10867,N_7237,N_6260);
nor U10868 (N_10868,N_7597,N_6101);
nand U10869 (N_10869,N_8288,N_7798);
and U10870 (N_10870,N_7331,N_7809);
and U10871 (N_10871,N_6433,N_7309);
nor U10872 (N_10872,N_8442,N_7102);
nor U10873 (N_10873,N_8263,N_6671);
nand U10874 (N_10874,N_8221,N_7765);
or U10875 (N_10875,N_6179,N_7526);
nor U10876 (N_10876,N_6867,N_7048);
nand U10877 (N_10877,N_7348,N_6397);
nor U10878 (N_10878,N_8577,N_8739);
nand U10879 (N_10879,N_8949,N_6534);
nor U10880 (N_10880,N_7839,N_7038);
or U10881 (N_10881,N_7786,N_7379);
nand U10882 (N_10882,N_7329,N_8952);
nor U10883 (N_10883,N_8260,N_8932);
and U10884 (N_10884,N_8702,N_6745);
nand U10885 (N_10885,N_6613,N_7451);
and U10886 (N_10886,N_7717,N_6972);
and U10887 (N_10887,N_6518,N_8909);
or U10888 (N_10888,N_8885,N_6381);
nand U10889 (N_10889,N_6422,N_8519);
nor U10890 (N_10890,N_8448,N_8669);
and U10891 (N_10891,N_8503,N_6255);
nor U10892 (N_10892,N_8907,N_7142);
or U10893 (N_10893,N_8893,N_8355);
nor U10894 (N_10894,N_6836,N_7462);
or U10895 (N_10895,N_6909,N_7248);
or U10896 (N_10896,N_8206,N_6043);
or U10897 (N_10897,N_7867,N_8715);
and U10898 (N_10898,N_8513,N_7112);
and U10899 (N_10899,N_8414,N_8254);
nand U10900 (N_10900,N_6425,N_8404);
xnor U10901 (N_10901,N_6919,N_6251);
nand U10902 (N_10902,N_7154,N_8965);
nand U10903 (N_10903,N_6778,N_7360);
and U10904 (N_10904,N_7436,N_7388);
or U10905 (N_10905,N_8841,N_7053);
nor U10906 (N_10906,N_7422,N_6026);
and U10907 (N_10907,N_7046,N_7148);
and U10908 (N_10908,N_7797,N_6615);
nand U10909 (N_10909,N_7690,N_8267);
and U10910 (N_10910,N_8749,N_8773);
and U10911 (N_10911,N_7235,N_8781);
and U10912 (N_10912,N_6461,N_8232);
or U10913 (N_10913,N_6979,N_7869);
or U10914 (N_10914,N_7541,N_6436);
nand U10915 (N_10915,N_6420,N_7412);
and U10916 (N_10916,N_7303,N_6937);
or U10917 (N_10917,N_6262,N_8225);
nand U10918 (N_10918,N_8108,N_6474);
and U10919 (N_10919,N_6403,N_6621);
and U10920 (N_10920,N_6678,N_8758);
and U10921 (N_10921,N_6668,N_8477);
or U10922 (N_10922,N_8629,N_8656);
or U10923 (N_10923,N_6983,N_6516);
nor U10924 (N_10924,N_8838,N_6863);
and U10925 (N_10925,N_6211,N_6701);
or U10926 (N_10926,N_7848,N_7054);
nor U10927 (N_10927,N_7593,N_7950);
nand U10928 (N_10928,N_7941,N_7662);
or U10929 (N_10929,N_8553,N_8033);
and U10930 (N_10930,N_8447,N_7777);
nand U10931 (N_10931,N_8673,N_8011);
nand U10932 (N_10932,N_6972,N_6573);
nand U10933 (N_10933,N_8689,N_7155);
nor U10934 (N_10934,N_8682,N_8758);
nand U10935 (N_10935,N_7652,N_6649);
and U10936 (N_10936,N_7094,N_6057);
nor U10937 (N_10937,N_7306,N_6194);
and U10938 (N_10938,N_7115,N_7134);
and U10939 (N_10939,N_6472,N_7012);
and U10940 (N_10940,N_7157,N_6897);
or U10941 (N_10941,N_7147,N_8002);
nand U10942 (N_10942,N_6879,N_6048);
or U10943 (N_10943,N_7163,N_6324);
and U10944 (N_10944,N_6106,N_8181);
and U10945 (N_10945,N_7597,N_6332);
nand U10946 (N_10946,N_7356,N_7755);
and U10947 (N_10947,N_8329,N_7138);
nand U10948 (N_10948,N_6097,N_8889);
and U10949 (N_10949,N_7653,N_6504);
nor U10950 (N_10950,N_8297,N_8622);
nand U10951 (N_10951,N_8039,N_7530);
nor U10952 (N_10952,N_6564,N_7457);
and U10953 (N_10953,N_8464,N_8135);
nor U10954 (N_10954,N_7255,N_6519);
or U10955 (N_10955,N_7340,N_7480);
nor U10956 (N_10956,N_6152,N_6787);
and U10957 (N_10957,N_8558,N_6967);
nand U10958 (N_10958,N_6289,N_7010);
nand U10959 (N_10959,N_7242,N_6114);
or U10960 (N_10960,N_6747,N_7478);
and U10961 (N_10961,N_8157,N_7405);
xnor U10962 (N_10962,N_6943,N_8196);
nor U10963 (N_10963,N_7785,N_8479);
and U10964 (N_10964,N_8441,N_8674);
or U10965 (N_10965,N_7877,N_6277);
xor U10966 (N_10966,N_6548,N_6198);
or U10967 (N_10967,N_7414,N_7162);
and U10968 (N_10968,N_6015,N_6586);
nand U10969 (N_10969,N_6801,N_6293);
nand U10970 (N_10970,N_7086,N_6240);
or U10971 (N_10971,N_6915,N_8225);
or U10972 (N_10972,N_6887,N_7142);
and U10973 (N_10973,N_7050,N_8703);
nor U10974 (N_10974,N_7433,N_7759);
and U10975 (N_10975,N_6165,N_7864);
nand U10976 (N_10976,N_7835,N_7462);
or U10977 (N_10977,N_6204,N_8309);
or U10978 (N_10978,N_6991,N_7292);
nor U10979 (N_10979,N_6288,N_8580);
and U10980 (N_10980,N_6167,N_7313);
nand U10981 (N_10981,N_8449,N_7715);
and U10982 (N_10982,N_6983,N_6979);
or U10983 (N_10983,N_7001,N_7334);
or U10984 (N_10984,N_7798,N_6757);
or U10985 (N_10985,N_6586,N_8407);
and U10986 (N_10986,N_7578,N_7845);
or U10987 (N_10987,N_7649,N_8729);
nand U10988 (N_10988,N_6992,N_8112);
or U10989 (N_10989,N_8624,N_6741);
or U10990 (N_10990,N_6532,N_7582);
or U10991 (N_10991,N_7754,N_6014);
or U10992 (N_10992,N_6420,N_7948);
and U10993 (N_10993,N_6525,N_6573);
and U10994 (N_10994,N_8110,N_7893);
nor U10995 (N_10995,N_6526,N_8931);
nor U10996 (N_10996,N_7896,N_8000);
nand U10997 (N_10997,N_8552,N_6005);
nor U10998 (N_10998,N_7127,N_8786);
or U10999 (N_10999,N_7750,N_7007);
or U11000 (N_11000,N_7815,N_7891);
nand U11001 (N_11001,N_8427,N_6310);
nand U11002 (N_11002,N_6164,N_7101);
and U11003 (N_11003,N_7750,N_6673);
nor U11004 (N_11004,N_6650,N_8342);
nand U11005 (N_11005,N_8351,N_6606);
and U11006 (N_11006,N_8572,N_7658);
and U11007 (N_11007,N_7254,N_8339);
nand U11008 (N_11008,N_7108,N_7518);
nand U11009 (N_11009,N_7575,N_8738);
nand U11010 (N_11010,N_7891,N_7228);
and U11011 (N_11011,N_6071,N_8769);
or U11012 (N_11012,N_8436,N_7741);
nand U11013 (N_11013,N_6959,N_8152);
or U11014 (N_11014,N_8955,N_7444);
nand U11015 (N_11015,N_6870,N_6435);
nand U11016 (N_11016,N_8847,N_6110);
xor U11017 (N_11017,N_7159,N_6988);
or U11018 (N_11018,N_7979,N_7288);
nand U11019 (N_11019,N_8166,N_7167);
nor U11020 (N_11020,N_7928,N_8644);
or U11021 (N_11021,N_8779,N_7181);
and U11022 (N_11022,N_8474,N_6844);
and U11023 (N_11023,N_8300,N_7222);
nand U11024 (N_11024,N_7818,N_6736);
nand U11025 (N_11025,N_7669,N_7023);
or U11026 (N_11026,N_7857,N_6842);
or U11027 (N_11027,N_8992,N_6014);
nor U11028 (N_11028,N_7944,N_6570);
or U11029 (N_11029,N_8055,N_8987);
nor U11030 (N_11030,N_7142,N_6690);
nand U11031 (N_11031,N_7959,N_7926);
or U11032 (N_11032,N_7868,N_6179);
nand U11033 (N_11033,N_7608,N_6869);
or U11034 (N_11034,N_6573,N_8260);
nand U11035 (N_11035,N_7421,N_7648);
nand U11036 (N_11036,N_7244,N_6815);
or U11037 (N_11037,N_8436,N_6942);
or U11038 (N_11038,N_8342,N_7918);
nand U11039 (N_11039,N_8662,N_6687);
nand U11040 (N_11040,N_7984,N_7184);
or U11041 (N_11041,N_8993,N_7679);
nor U11042 (N_11042,N_6074,N_7216);
nor U11043 (N_11043,N_8389,N_6502);
nand U11044 (N_11044,N_7805,N_8970);
or U11045 (N_11045,N_8523,N_7657);
or U11046 (N_11046,N_8798,N_6636);
and U11047 (N_11047,N_8762,N_7234);
nor U11048 (N_11048,N_8860,N_6195);
nor U11049 (N_11049,N_7395,N_8581);
nor U11050 (N_11050,N_8989,N_8336);
nor U11051 (N_11051,N_8665,N_6073);
nand U11052 (N_11052,N_8444,N_6256);
and U11053 (N_11053,N_7363,N_8289);
nor U11054 (N_11054,N_6970,N_6312);
or U11055 (N_11055,N_7947,N_6115);
or U11056 (N_11056,N_6780,N_8568);
or U11057 (N_11057,N_7300,N_8567);
and U11058 (N_11058,N_7956,N_6810);
nor U11059 (N_11059,N_7954,N_7280);
and U11060 (N_11060,N_8867,N_6309);
nand U11061 (N_11061,N_8969,N_7551);
or U11062 (N_11062,N_6948,N_6077);
or U11063 (N_11063,N_8498,N_7401);
or U11064 (N_11064,N_8686,N_8340);
xor U11065 (N_11065,N_8827,N_6082);
or U11066 (N_11066,N_8281,N_8546);
nand U11067 (N_11067,N_7552,N_8071);
xor U11068 (N_11068,N_7134,N_6868);
and U11069 (N_11069,N_6746,N_6408);
and U11070 (N_11070,N_8313,N_7502);
and U11071 (N_11071,N_8380,N_6397);
nand U11072 (N_11072,N_6199,N_8955);
nand U11073 (N_11073,N_6881,N_7810);
nand U11074 (N_11074,N_7997,N_7252);
or U11075 (N_11075,N_7999,N_7749);
nand U11076 (N_11076,N_7527,N_6947);
and U11077 (N_11077,N_8625,N_8421);
and U11078 (N_11078,N_8677,N_8878);
nand U11079 (N_11079,N_8509,N_6890);
nor U11080 (N_11080,N_7665,N_7308);
and U11081 (N_11081,N_6314,N_8462);
nor U11082 (N_11082,N_6790,N_6594);
nor U11083 (N_11083,N_6233,N_6242);
nand U11084 (N_11084,N_8028,N_8442);
nor U11085 (N_11085,N_6844,N_8723);
and U11086 (N_11086,N_8963,N_7612);
nand U11087 (N_11087,N_7773,N_8232);
nand U11088 (N_11088,N_7318,N_7497);
nand U11089 (N_11089,N_6705,N_7418);
and U11090 (N_11090,N_7612,N_6419);
nor U11091 (N_11091,N_7833,N_8486);
or U11092 (N_11092,N_7432,N_8092);
nor U11093 (N_11093,N_6411,N_7297);
nand U11094 (N_11094,N_7901,N_6212);
nor U11095 (N_11095,N_6276,N_8362);
nor U11096 (N_11096,N_8861,N_6631);
and U11097 (N_11097,N_8836,N_6169);
or U11098 (N_11098,N_7346,N_7839);
and U11099 (N_11099,N_6757,N_6642);
or U11100 (N_11100,N_7635,N_8321);
and U11101 (N_11101,N_7560,N_7353);
nand U11102 (N_11102,N_7962,N_8721);
nor U11103 (N_11103,N_6567,N_7642);
and U11104 (N_11104,N_8570,N_8550);
or U11105 (N_11105,N_7597,N_7243);
nor U11106 (N_11106,N_7735,N_8447);
nor U11107 (N_11107,N_6238,N_7409);
and U11108 (N_11108,N_8960,N_8603);
nor U11109 (N_11109,N_6821,N_7948);
nand U11110 (N_11110,N_6090,N_6741);
nor U11111 (N_11111,N_6106,N_7245);
or U11112 (N_11112,N_6533,N_8005);
nor U11113 (N_11113,N_7982,N_7585);
nand U11114 (N_11114,N_7155,N_6052);
nor U11115 (N_11115,N_6680,N_6370);
and U11116 (N_11116,N_6182,N_6503);
nand U11117 (N_11117,N_8605,N_7684);
or U11118 (N_11118,N_8869,N_8214);
xnor U11119 (N_11119,N_7962,N_8525);
nor U11120 (N_11120,N_7939,N_6746);
and U11121 (N_11121,N_7079,N_8436);
nor U11122 (N_11122,N_7294,N_7349);
nor U11123 (N_11123,N_6269,N_7757);
nor U11124 (N_11124,N_6531,N_8542);
nand U11125 (N_11125,N_7492,N_6307);
nor U11126 (N_11126,N_6496,N_7462);
or U11127 (N_11127,N_6409,N_6195);
nand U11128 (N_11128,N_6873,N_6234);
and U11129 (N_11129,N_8474,N_8805);
nor U11130 (N_11130,N_8272,N_6136);
nor U11131 (N_11131,N_6774,N_7340);
nand U11132 (N_11132,N_7337,N_6407);
or U11133 (N_11133,N_6962,N_8046);
nor U11134 (N_11134,N_6600,N_8784);
or U11135 (N_11135,N_7842,N_6696);
nand U11136 (N_11136,N_8697,N_8506);
and U11137 (N_11137,N_8332,N_7546);
and U11138 (N_11138,N_7859,N_8656);
nor U11139 (N_11139,N_8710,N_8828);
and U11140 (N_11140,N_7468,N_7732);
nor U11141 (N_11141,N_6356,N_8370);
and U11142 (N_11142,N_8136,N_7443);
nor U11143 (N_11143,N_7189,N_7425);
nor U11144 (N_11144,N_8927,N_7886);
nor U11145 (N_11145,N_8565,N_6598);
and U11146 (N_11146,N_7368,N_8340);
and U11147 (N_11147,N_6418,N_8124);
nand U11148 (N_11148,N_8007,N_8105);
and U11149 (N_11149,N_8427,N_6457);
nand U11150 (N_11150,N_8764,N_6367);
or U11151 (N_11151,N_7787,N_6956);
or U11152 (N_11152,N_6502,N_7706);
nor U11153 (N_11153,N_7826,N_6871);
nor U11154 (N_11154,N_7025,N_6206);
nor U11155 (N_11155,N_7518,N_7186);
and U11156 (N_11156,N_7966,N_7875);
nor U11157 (N_11157,N_6553,N_8764);
and U11158 (N_11158,N_6484,N_6688);
nand U11159 (N_11159,N_7320,N_8240);
nand U11160 (N_11160,N_7206,N_8518);
or U11161 (N_11161,N_8475,N_6715);
xnor U11162 (N_11162,N_6280,N_6268);
nand U11163 (N_11163,N_8769,N_6227);
nand U11164 (N_11164,N_7957,N_7610);
nor U11165 (N_11165,N_6151,N_6930);
and U11166 (N_11166,N_8201,N_7868);
xnor U11167 (N_11167,N_7725,N_8887);
xnor U11168 (N_11168,N_6975,N_6984);
nand U11169 (N_11169,N_6798,N_7831);
xnor U11170 (N_11170,N_7454,N_8237);
and U11171 (N_11171,N_8712,N_7464);
nand U11172 (N_11172,N_8476,N_8806);
nand U11173 (N_11173,N_8141,N_7059);
nor U11174 (N_11174,N_7673,N_8022);
nand U11175 (N_11175,N_7222,N_6726);
or U11176 (N_11176,N_8086,N_8328);
nor U11177 (N_11177,N_8877,N_6589);
nor U11178 (N_11178,N_7727,N_6737);
or U11179 (N_11179,N_7900,N_8307);
or U11180 (N_11180,N_6169,N_8161);
nor U11181 (N_11181,N_7862,N_6268);
nor U11182 (N_11182,N_7232,N_8443);
nand U11183 (N_11183,N_6083,N_6397);
nor U11184 (N_11184,N_8565,N_6414);
nand U11185 (N_11185,N_6277,N_6274);
or U11186 (N_11186,N_6051,N_6551);
or U11187 (N_11187,N_6572,N_6636);
or U11188 (N_11188,N_7458,N_7026);
or U11189 (N_11189,N_8789,N_8496);
or U11190 (N_11190,N_6416,N_7014);
nand U11191 (N_11191,N_6808,N_8653);
and U11192 (N_11192,N_6830,N_7813);
nor U11193 (N_11193,N_6921,N_6765);
nand U11194 (N_11194,N_7772,N_6941);
xor U11195 (N_11195,N_8001,N_8496);
nor U11196 (N_11196,N_7052,N_6547);
nor U11197 (N_11197,N_7769,N_6164);
nor U11198 (N_11198,N_6476,N_8207);
or U11199 (N_11199,N_6371,N_8801);
nor U11200 (N_11200,N_7824,N_7436);
and U11201 (N_11201,N_7346,N_6664);
or U11202 (N_11202,N_8643,N_8413);
nand U11203 (N_11203,N_6036,N_6293);
nand U11204 (N_11204,N_7221,N_7700);
nand U11205 (N_11205,N_6149,N_7998);
nor U11206 (N_11206,N_7408,N_7417);
nor U11207 (N_11207,N_6182,N_6029);
nand U11208 (N_11208,N_6277,N_6979);
or U11209 (N_11209,N_7466,N_8777);
nand U11210 (N_11210,N_8589,N_8706);
and U11211 (N_11211,N_6006,N_6770);
and U11212 (N_11212,N_6522,N_7791);
or U11213 (N_11213,N_7528,N_7734);
or U11214 (N_11214,N_8728,N_6654);
nor U11215 (N_11215,N_6781,N_7950);
and U11216 (N_11216,N_8793,N_8352);
nor U11217 (N_11217,N_8774,N_7731);
nor U11218 (N_11218,N_6274,N_8626);
nand U11219 (N_11219,N_7496,N_6126);
nor U11220 (N_11220,N_8325,N_6810);
nand U11221 (N_11221,N_6756,N_6481);
nor U11222 (N_11222,N_8176,N_8550);
nor U11223 (N_11223,N_7532,N_7261);
nand U11224 (N_11224,N_6815,N_8111);
and U11225 (N_11225,N_7976,N_7374);
and U11226 (N_11226,N_6949,N_6140);
or U11227 (N_11227,N_6794,N_7012);
or U11228 (N_11228,N_6081,N_8828);
and U11229 (N_11229,N_6347,N_7414);
nand U11230 (N_11230,N_8968,N_7525);
nor U11231 (N_11231,N_8810,N_8156);
and U11232 (N_11232,N_6033,N_7167);
or U11233 (N_11233,N_7229,N_6679);
nor U11234 (N_11234,N_6122,N_6682);
nand U11235 (N_11235,N_7790,N_7252);
and U11236 (N_11236,N_6451,N_8045);
and U11237 (N_11237,N_7686,N_6078);
nand U11238 (N_11238,N_7269,N_6176);
and U11239 (N_11239,N_7049,N_7140);
nand U11240 (N_11240,N_8914,N_6582);
and U11241 (N_11241,N_8509,N_6012);
nand U11242 (N_11242,N_7007,N_6030);
nand U11243 (N_11243,N_7184,N_6695);
nor U11244 (N_11244,N_8010,N_8936);
nor U11245 (N_11245,N_6068,N_7439);
nor U11246 (N_11246,N_8106,N_8740);
and U11247 (N_11247,N_8710,N_8667);
and U11248 (N_11248,N_6958,N_6978);
and U11249 (N_11249,N_7927,N_7434);
and U11250 (N_11250,N_6709,N_7155);
nor U11251 (N_11251,N_6529,N_7264);
nor U11252 (N_11252,N_7884,N_6707);
nor U11253 (N_11253,N_7784,N_6132);
nand U11254 (N_11254,N_6456,N_6275);
and U11255 (N_11255,N_7072,N_8133);
nand U11256 (N_11256,N_6617,N_8354);
nand U11257 (N_11257,N_8326,N_7132);
and U11258 (N_11258,N_7520,N_7521);
or U11259 (N_11259,N_8055,N_8585);
nor U11260 (N_11260,N_6049,N_7377);
and U11261 (N_11261,N_7404,N_6429);
or U11262 (N_11262,N_8134,N_7206);
and U11263 (N_11263,N_8869,N_6525);
and U11264 (N_11264,N_8643,N_6954);
nand U11265 (N_11265,N_6548,N_6388);
nand U11266 (N_11266,N_7912,N_7422);
nand U11267 (N_11267,N_7586,N_6885);
nor U11268 (N_11268,N_7482,N_6477);
and U11269 (N_11269,N_7286,N_7100);
nor U11270 (N_11270,N_7314,N_6349);
and U11271 (N_11271,N_8319,N_7218);
and U11272 (N_11272,N_8098,N_7404);
and U11273 (N_11273,N_6160,N_6185);
nand U11274 (N_11274,N_6975,N_6620);
or U11275 (N_11275,N_6360,N_8852);
and U11276 (N_11276,N_6861,N_8050);
or U11277 (N_11277,N_6247,N_6788);
nand U11278 (N_11278,N_8795,N_8770);
and U11279 (N_11279,N_7813,N_6788);
and U11280 (N_11280,N_6818,N_7717);
nand U11281 (N_11281,N_7004,N_8870);
nor U11282 (N_11282,N_7549,N_6650);
xnor U11283 (N_11283,N_8182,N_8195);
nor U11284 (N_11284,N_6199,N_8835);
nor U11285 (N_11285,N_6989,N_8974);
nand U11286 (N_11286,N_6270,N_8815);
nand U11287 (N_11287,N_8562,N_6120);
and U11288 (N_11288,N_6110,N_8503);
nand U11289 (N_11289,N_6446,N_6252);
and U11290 (N_11290,N_7928,N_8752);
nor U11291 (N_11291,N_7833,N_7582);
nor U11292 (N_11292,N_6857,N_6550);
and U11293 (N_11293,N_6685,N_7536);
nor U11294 (N_11294,N_8507,N_6300);
and U11295 (N_11295,N_6894,N_8400);
nand U11296 (N_11296,N_7042,N_6314);
and U11297 (N_11297,N_6317,N_6786);
or U11298 (N_11298,N_7374,N_6863);
nor U11299 (N_11299,N_6944,N_7392);
and U11300 (N_11300,N_6913,N_7205);
nor U11301 (N_11301,N_7263,N_6626);
nor U11302 (N_11302,N_8751,N_7363);
nor U11303 (N_11303,N_7935,N_6665);
nor U11304 (N_11304,N_8268,N_7041);
nor U11305 (N_11305,N_8957,N_7675);
xnor U11306 (N_11306,N_7864,N_6934);
or U11307 (N_11307,N_7599,N_6950);
nor U11308 (N_11308,N_6054,N_7333);
nand U11309 (N_11309,N_6534,N_7694);
nor U11310 (N_11310,N_6070,N_6116);
or U11311 (N_11311,N_7786,N_8601);
nor U11312 (N_11312,N_7510,N_7500);
nor U11313 (N_11313,N_8074,N_8760);
nand U11314 (N_11314,N_7812,N_8149);
or U11315 (N_11315,N_8492,N_6940);
and U11316 (N_11316,N_8206,N_7691);
nor U11317 (N_11317,N_8773,N_6478);
and U11318 (N_11318,N_7394,N_8674);
and U11319 (N_11319,N_6752,N_7257);
and U11320 (N_11320,N_6533,N_7533);
nor U11321 (N_11321,N_7048,N_7856);
nor U11322 (N_11322,N_6035,N_7403);
or U11323 (N_11323,N_7462,N_6431);
nor U11324 (N_11324,N_8278,N_6043);
or U11325 (N_11325,N_7742,N_8277);
nand U11326 (N_11326,N_6788,N_7477);
nand U11327 (N_11327,N_8950,N_8172);
nand U11328 (N_11328,N_8106,N_8652);
nand U11329 (N_11329,N_6681,N_6403);
or U11330 (N_11330,N_8172,N_6244);
nor U11331 (N_11331,N_8465,N_8038);
nor U11332 (N_11332,N_8158,N_8433);
and U11333 (N_11333,N_8568,N_8191);
nand U11334 (N_11334,N_8062,N_6116);
and U11335 (N_11335,N_7775,N_7288);
nand U11336 (N_11336,N_7593,N_6794);
or U11337 (N_11337,N_7779,N_6167);
or U11338 (N_11338,N_6421,N_6252);
nor U11339 (N_11339,N_8680,N_7490);
and U11340 (N_11340,N_8232,N_6448);
and U11341 (N_11341,N_6167,N_7272);
nor U11342 (N_11342,N_7275,N_6878);
nand U11343 (N_11343,N_7731,N_7667);
nor U11344 (N_11344,N_6338,N_6439);
nor U11345 (N_11345,N_8299,N_8064);
or U11346 (N_11346,N_8269,N_7137);
or U11347 (N_11347,N_8716,N_7833);
nor U11348 (N_11348,N_6304,N_7903);
or U11349 (N_11349,N_8539,N_8001);
or U11350 (N_11350,N_8264,N_6422);
or U11351 (N_11351,N_6490,N_6578);
nor U11352 (N_11352,N_6801,N_6498);
and U11353 (N_11353,N_7894,N_8789);
or U11354 (N_11354,N_7145,N_6344);
or U11355 (N_11355,N_7234,N_8274);
nand U11356 (N_11356,N_8821,N_7028);
and U11357 (N_11357,N_8812,N_7994);
and U11358 (N_11358,N_7912,N_7655);
nor U11359 (N_11359,N_7290,N_7371);
nand U11360 (N_11360,N_7401,N_6486);
nand U11361 (N_11361,N_8376,N_7473);
nand U11362 (N_11362,N_8544,N_6773);
nor U11363 (N_11363,N_8450,N_7511);
and U11364 (N_11364,N_7879,N_6918);
or U11365 (N_11365,N_6205,N_8283);
nor U11366 (N_11366,N_8844,N_7093);
and U11367 (N_11367,N_7287,N_8005);
or U11368 (N_11368,N_6027,N_7975);
and U11369 (N_11369,N_7912,N_8650);
nand U11370 (N_11370,N_6122,N_6115);
nand U11371 (N_11371,N_7379,N_7254);
nor U11372 (N_11372,N_6270,N_8781);
nor U11373 (N_11373,N_8644,N_6254);
and U11374 (N_11374,N_8242,N_8300);
nor U11375 (N_11375,N_6873,N_7071);
nor U11376 (N_11376,N_7710,N_8605);
and U11377 (N_11377,N_6217,N_8650);
nor U11378 (N_11378,N_7186,N_6959);
or U11379 (N_11379,N_6154,N_8933);
or U11380 (N_11380,N_7575,N_8355);
nor U11381 (N_11381,N_7202,N_7798);
nor U11382 (N_11382,N_7622,N_6015);
or U11383 (N_11383,N_8811,N_8096);
xnor U11384 (N_11384,N_7643,N_8712);
and U11385 (N_11385,N_6366,N_7832);
and U11386 (N_11386,N_7363,N_8924);
nand U11387 (N_11387,N_6660,N_6617);
nor U11388 (N_11388,N_8715,N_6800);
or U11389 (N_11389,N_8689,N_8066);
and U11390 (N_11390,N_7690,N_6486);
nor U11391 (N_11391,N_6575,N_6629);
nand U11392 (N_11392,N_7317,N_6954);
nand U11393 (N_11393,N_8281,N_6519);
and U11394 (N_11394,N_8035,N_6540);
and U11395 (N_11395,N_8543,N_7693);
and U11396 (N_11396,N_8677,N_6558);
nand U11397 (N_11397,N_6651,N_8231);
nor U11398 (N_11398,N_7789,N_6334);
or U11399 (N_11399,N_6017,N_8726);
nor U11400 (N_11400,N_8419,N_7582);
and U11401 (N_11401,N_7894,N_7030);
nand U11402 (N_11402,N_8578,N_8930);
and U11403 (N_11403,N_6534,N_8871);
and U11404 (N_11404,N_7375,N_6491);
or U11405 (N_11405,N_6816,N_6012);
and U11406 (N_11406,N_6172,N_8146);
or U11407 (N_11407,N_7218,N_7179);
nor U11408 (N_11408,N_7602,N_8057);
nand U11409 (N_11409,N_7777,N_6173);
or U11410 (N_11410,N_8551,N_8780);
nand U11411 (N_11411,N_7212,N_7253);
nor U11412 (N_11412,N_7035,N_7486);
and U11413 (N_11413,N_7207,N_8192);
or U11414 (N_11414,N_6371,N_6034);
nand U11415 (N_11415,N_6347,N_8011);
or U11416 (N_11416,N_6155,N_6118);
and U11417 (N_11417,N_7399,N_6119);
and U11418 (N_11418,N_7571,N_8260);
and U11419 (N_11419,N_7607,N_6261);
xnor U11420 (N_11420,N_8953,N_7924);
and U11421 (N_11421,N_6272,N_7942);
nand U11422 (N_11422,N_6137,N_8513);
and U11423 (N_11423,N_6085,N_6060);
xor U11424 (N_11424,N_8010,N_6958);
or U11425 (N_11425,N_6677,N_8447);
nor U11426 (N_11426,N_8775,N_6686);
and U11427 (N_11427,N_6591,N_6814);
nor U11428 (N_11428,N_6418,N_7578);
nor U11429 (N_11429,N_7569,N_7942);
nand U11430 (N_11430,N_7743,N_7160);
and U11431 (N_11431,N_7780,N_6657);
nor U11432 (N_11432,N_6175,N_8543);
nor U11433 (N_11433,N_8150,N_7419);
and U11434 (N_11434,N_8688,N_6087);
and U11435 (N_11435,N_6605,N_6288);
nand U11436 (N_11436,N_8845,N_6517);
or U11437 (N_11437,N_7644,N_8249);
and U11438 (N_11438,N_7491,N_7951);
and U11439 (N_11439,N_8966,N_7000);
nor U11440 (N_11440,N_6053,N_7271);
nor U11441 (N_11441,N_6420,N_7543);
nor U11442 (N_11442,N_7894,N_7915);
and U11443 (N_11443,N_6340,N_6918);
nand U11444 (N_11444,N_8179,N_8003);
or U11445 (N_11445,N_8947,N_8566);
or U11446 (N_11446,N_6118,N_6336);
and U11447 (N_11447,N_8570,N_7764);
nor U11448 (N_11448,N_6828,N_7011);
nor U11449 (N_11449,N_8298,N_6682);
or U11450 (N_11450,N_7160,N_7325);
nand U11451 (N_11451,N_8034,N_7135);
nor U11452 (N_11452,N_6394,N_7946);
or U11453 (N_11453,N_7753,N_8348);
nand U11454 (N_11454,N_8281,N_6820);
nor U11455 (N_11455,N_6523,N_8313);
nand U11456 (N_11456,N_6263,N_6227);
and U11457 (N_11457,N_7552,N_7569);
xor U11458 (N_11458,N_8202,N_8591);
xor U11459 (N_11459,N_8202,N_8872);
or U11460 (N_11460,N_8886,N_8475);
nand U11461 (N_11461,N_8633,N_7282);
nor U11462 (N_11462,N_6027,N_6539);
and U11463 (N_11463,N_7337,N_7730);
or U11464 (N_11464,N_6576,N_7684);
nand U11465 (N_11465,N_8364,N_7601);
and U11466 (N_11466,N_6792,N_8203);
nor U11467 (N_11467,N_6003,N_7779);
or U11468 (N_11468,N_6679,N_8184);
or U11469 (N_11469,N_8121,N_8411);
and U11470 (N_11470,N_7618,N_8831);
nor U11471 (N_11471,N_7296,N_7392);
or U11472 (N_11472,N_8982,N_8877);
and U11473 (N_11473,N_8683,N_6420);
xnor U11474 (N_11474,N_7964,N_6714);
nand U11475 (N_11475,N_8334,N_7002);
xor U11476 (N_11476,N_6176,N_6904);
and U11477 (N_11477,N_8767,N_8685);
or U11478 (N_11478,N_7299,N_8039);
and U11479 (N_11479,N_7429,N_8268);
nor U11480 (N_11480,N_8367,N_7155);
and U11481 (N_11481,N_6736,N_8923);
nor U11482 (N_11482,N_7008,N_8547);
nand U11483 (N_11483,N_7876,N_8793);
and U11484 (N_11484,N_6677,N_6203);
nand U11485 (N_11485,N_7520,N_6190);
nand U11486 (N_11486,N_8988,N_8777);
nor U11487 (N_11487,N_6385,N_8325);
nor U11488 (N_11488,N_6528,N_7929);
nand U11489 (N_11489,N_6803,N_6125);
nand U11490 (N_11490,N_6593,N_8142);
nor U11491 (N_11491,N_6380,N_8384);
nor U11492 (N_11492,N_8384,N_7437);
nand U11493 (N_11493,N_6722,N_7797);
or U11494 (N_11494,N_8579,N_6825);
or U11495 (N_11495,N_7810,N_6815);
nand U11496 (N_11496,N_6980,N_6525);
nand U11497 (N_11497,N_7896,N_6543);
or U11498 (N_11498,N_8761,N_8548);
and U11499 (N_11499,N_7128,N_6384);
nand U11500 (N_11500,N_6945,N_6880);
nor U11501 (N_11501,N_8194,N_6086);
nand U11502 (N_11502,N_7936,N_7510);
nor U11503 (N_11503,N_7850,N_7185);
nor U11504 (N_11504,N_6694,N_7810);
and U11505 (N_11505,N_7943,N_7597);
nand U11506 (N_11506,N_6735,N_6402);
nor U11507 (N_11507,N_8483,N_8345);
and U11508 (N_11508,N_6841,N_8261);
or U11509 (N_11509,N_7107,N_8493);
or U11510 (N_11510,N_8131,N_7302);
and U11511 (N_11511,N_7746,N_8129);
or U11512 (N_11512,N_6926,N_7460);
and U11513 (N_11513,N_7408,N_7342);
nor U11514 (N_11514,N_7875,N_6836);
or U11515 (N_11515,N_6762,N_6646);
nor U11516 (N_11516,N_8213,N_8796);
or U11517 (N_11517,N_8577,N_6896);
nand U11518 (N_11518,N_7286,N_8595);
or U11519 (N_11519,N_6314,N_7311);
or U11520 (N_11520,N_8239,N_8551);
and U11521 (N_11521,N_6465,N_7391);
nor U11522 (N_11522,N_7305,N_6854);
nor U11523 (N_11523,N_8767,N_6332);
or U11524 (N_11524,N_6443,N_6566);
and U11525 (N_11525,N_7887,N_8412);
nand U11526 (N_11526,N_7824,N_7134);
nand U11527 (N_11527,N_8380,N_8059);
nor U11528 (N_11528,N_7132,N_7011);
or U11529 (N_11529,N_6339,N_6808);
and U11530 (N_11530,N_8023,N_8919);
nor U11531 (N_11531,N_7068,N_8610);
and U11532 (N_11532,N_6049,N_6858);
nand U11533 (N_11533,N_7737,N_7228);
nor U11534 (N_11534,N_8301,N_7665);
nand U11535 (N_11535,N_6800,N_6606);
and U11536 (N_11536,N_6985,N_8052);
nor U11537 (N_11537,N_6377,N_6096);
and U11538 (N_11538,N_7811,N_7013);
and U11539 (N_11539,N_6677,N_7304);
and U11540 (N_11540,N_7586,N_6402);
nand U11541 (N_11541,N_7663,N_7829);
nor U11542 (N_11542,N_6261,N_6790);
nand U11543 (N_11543,N_7441,N_8248);
or U11544 (N_11544,N_8702,N_6333);
and U11545 (N_11545,N_8074,N_6901);
nor U11546 (N_11546,N_6818,N_6113);
nor U11547 (N_11547,N_6238,N_7565);
and U11548 (N_11548,N_6429,N_6338);
nand U11549 (N_11549,N_6427,N_6716);
nand U11550 (N_11550,N_8229,N_7953);
nor U11551 (N_11551,N_6990,N_7880);
or U11552 (N_11552,N_8720,N_7038);
nor U11553 (N_11553,N_8877,N_8500);
nor U11554 (N_11554,N_7503,N_7251);
nand U11555 (N_11555,N_7818,N_6820);
or U11556 (N_11556,N_6009,N_7997);
nor U11557 (N_11557,N_6490,N_7336);
nor U11558 (N_11558,N_6321,N_8419);
nand U11559 (N_11559,N_6017,N_7099);
nand U11560 (N_11560,N_7875,N_6336);
nor U11561 (N_11561,N_8411,N_7683);
nor U11562 (N_11562,N_7306,N_8199);
or U11563 (N_11563,N_8598,N_6678);
nand U11564 (N_11564,N_6504,N_7667);
nor U11565 (N_11565,N_8280,N_6316);
nor U11566 (N_11566,N_8194,N_6232);
or U11567 (N_11567,N_8072,N_7619);
nand U11568 (N_11568,N_7723,N_7825);
xnor U11569 (N_11569,N_8730,N_8303);
nand U11570 (N_11570,N_8522,N_7638);
nand U11571 (N_11571,N_6618,N_6101);
nand U11572 (N_11572,N_7551,N_7839);
and U11573 (N_11573,N_8875,N_7331);
nand U11574 (N_11574,N_7339,N_8282);
nor U11575 (N_11575,N_6730,N_7643);
nand U11576 (N_11576,N_8540,N_8023);
or U11577 (N_11577,N_8875,N_8078);
nand U11578 (N_11578,N_8460,N_8828);
nand U11579 (N_11579,N_8245,N_7562);
or U11580 (N_11580,N_6518,N_6967);
or U11581 (N_11581,N_8566,N_7753);
and U11582 (N_11582,N_6186,N_7882);
and U11583 (N_11583,N_8384,N_6983);
and U11584 (N_11584,N_7922,N_7940);
nor U11585 (N_11585,N_6163,N_6490);
or U11586 (N_11586,N_7357,N_6951);
and U11587 (N_11587,N_7963,N_6693);
and U11588 (N_11588,N_7415,N_8579);
or U11589 (N_11589,N_6058,N_6570);
nand U11590 (N_11590,N_6223,N_7180);
nand U11591 (N_11591,N_6900,N_7462);
nor U11592 (N_11592,N_8574,N_8298);
or U11593 (N_11593,N_8904,N_6208);
nor U11594 (N_11594,N_8278,N_6791);
nand U11595 (N_11595,N_8251,N_7688);
nand U11596 (N_11596,N_7251,N_6705);
nand U11597 (N_11597,N_8552,N_6603);
and U11598 (N_11598,N_7343,N_8454);
nor U11599 (N_11599,N_8588,N_6873);
or U11600 (N_11600,N_7636,N_8822);
nor U11601 (N_11601,N_8527,N_8600);
and U11602 (N_11602,N_8379,N_8736);
nand U11603 (N_11603,N_8204,N_8010);
nand U11604 (N_11604,N_7248,N_7397);
or U11605 (N_11605,N_7807,N_8737);
nor U11606 (N_11606,N_7199,N_6929);
nand U11607 (N_11607,N_7059,N_7012);
nor U11608 (N_11608,N_6174,N_8415);
nor U11609 (N_11609,N_8588,N_7730);
and U11610 (N_11610,N_8626,N_7742);
nor U11611 (N_11611,N_8654,N_6815);
nand U11612 (N_11612,N_6711,N_7297);
or U11613 (N_11613,N_8298,N_6830);
nand U11614 (N_11614,N_8416,N_6141);
or U11615 (N_11615,N_8786,N_7099);
and U11616 (N_11616,N_7608,N_7778);
and U11617 (N_11617,N_7963,N_7285);
and U11618 (N_11618,N_8661,N_8752);
or U11619 (N_11619,N_6920,N_8612);
nor U11620 (N_11620,N_8015,N_6251);
xnor U11621 (N_11621,N_7748,N_6163);
or U11622 (N_11622,N_6771,N_7085);
nand U11623 (N_11623,N_8033,N_8942);
xor U11624 (N_11624,N_8738,N_6777);
nor U11625 (N_11625,N_8538,N_8768);
or U11626 (N_11626,N_6959,N_8411);
and U11627 (N_11627,N_6639,N_6585);
nor U11628 (N_11628,N_8703,N_7111);
and U11629 (N_11629,N_6156,N_6625);
or U11630 (N_11630,N_6571,N_6126);
nor U11631 (N_11631,N_7950,N_7723);
nand U11632 (N_11632,N_7721,N_8861);
or U11633 (N_11633,N_6168,N_6833);
nor U11634 (N_11634,N_8119,N_7705);
nand U11635 (N_11635,N_7178,N_6746);
xor U11636 (N_11636,N_7685,N_7326);
nand U11637 (N_11637,N_6047,N_7359);
nand U11638 (N_11638,N_7367,N_8594);
nor U11639 (N_11639,N_6125,N_8104);
nor U11640 (N_11640,N_8594,N_7776);
or U11641 (N_11641,N_8675,N_8833);
xnor U11642 (N_11642,N_8449,N_7466);
or U11643 (N_11643,N_6119,N_7931);
nand U11644 (N_11644,N_6266,N_7312);
and U11645 (N_11645,N_6571,N_7582);
and U11646 (N_11646,N_6235,N_6199);
nand U11647 (N_11647,N_7342,N_8761);
or U11648 (N_11648,N_8858,N_6440);
nand U11649 (N_11649,N_7438,N_6688);
and U11650 (N_11650,N_8810,N_6823);
nor U11651 (N_11651,N_6816,N_7536);
nand U11652 (N_11652,N_8828,N_7515);
and U11653 (N_11653,N_6136,N_7382);
nand U11654 (N_11654,N_6984,N_7647);
or U11655 (N_11655,N_6739,N_8043);
nor U11656 (N_11656,N_7201,N_6542);
and U11657 (N_11657,N_6256,N_7687);
or U11658 (N_11658,N_7066,N_7326);
nand U11659 (N_11659,N_8704,N_7420);
and U11660 (N_11660,N_6947,N_6838);
or U11661 (N_11661,N_8118,N_6390);
or U11662 (N_11662,N_8128,N_6116);
or U11663 (N_11663,N_7611,N_8931);
or U11664 (N_11664,N_8803,N_8494);
nand U11665 (N_11665,N_8173,N_8418);
or U11666 (N_11666,N_7508,N_7586);
nor U11667 (N_11667,N_8626,N_7924);
nor U11668 (N_11668,N_8885,N_8706);
nor U11669 (N_11669,N_8952,N_6235);
nand U11670 (N_11670,N_7262,N_7729);
nor U11671 (N_11671,N_6167,N_6284);
nor U11672 (N_11672,N_8288,N_6614);
xor U11673 (N_11673,N_6130,N_8949);
nand U11674 (N_11674,N_7652,N_8068);
nor U11675 (N_11675,N_6433,N_8033);
and U11676 (N_11676,N_6033,N_8704);
or U11677 (N_11677,N_8020,N_7344);
or U11678 (N_11678,N_8772,N_6453);
xnor U11679 (N_11679,N_6167,N_6918);
nand U11680 (N_11680,N_7500,N_7073);
nor U11681 (N_11681,N_7251,N_7600);
and U11682 (N_11682,N_6184,N_8181);
nand U11683 (N_11683,N_6835,N_6108);
nor U11684 (N_11684,N_6529,N_6328);
nand U11685 (N_11685,N_7879,N_7808);
or U11686 (N_11686,N_8951,N_7488);
nand U11687 (N_11687,N_8469,N_8605);
nor U11688 (N_11688,N_7291,N_8928);
nand U11689 (N_11689,N_7507,N_6686);
nor U11690 (N_11690,N_7301,N_7005);
or U11691 (N_11691,N_7409,N_8466);
and U11692 (N_11692,N_7180,N_8327);
and U11693 (N_11693,N_8362,N_8830);
or U11694 (N_11694,N_8539,N_6833);
xor U11695 (N_11695,N_6092,N_7994);
nor U11696 (N_11696,N_8123,N_7514);
and U11697 (N_11697,N_7277,N_8287);
or U11698 (N_11698,N_7109,N_8869);
nand U11699 (N_11699,N_6211,N_8086);
nand U11700 (N_11700,N_7168,N_6754);
and U11701 (N_11701,N_6183,N_8065);
or U11702 (N_11702,N_7665,N_7443);
nor U11703 (N_11703,N_7905,N_7673);
and U11704 (N_11704,N_7818,N_8260);
nand U11705 (N_11705,N_8886,N_7113);
and U11706 (N_11706,N_7575,N_7901);
and U11707 (N_11707,N_8195,N_7232);
nand U11708 (N_11708,N_8499,N_7525);
nand U11709 (N_11709,N_7072,N_8267);
nand U11710 (N_11710,N_7289,N_6740);
nand U11711 (N_11711,N_7563,N_7383);
and U11712 (N_11712,N_7382,N_6183);
and U11713 (N_11713,N_8807,N_8779);
nor U11714 (N_11714,N_6385,N_7562);
nand U11715 (N_11715,N_6148,N_6128);
nor U11716 (N_11716,N_8941,N_8542);
nand U11717 (N_11717,N_6645,N_6082);
nor U11718 (N_11718,N_7491,N_7780);
or U11719 (N_11719,N_6402,N_7451);
or U11720 (N_11720,N_8965,N_6413);
nand U11721 (N_11721,N_7138,N_8395);
nand U11722 (N_11722,N_7507,N_7338);
and U11723 (N_11723,N_7066,N_7406);
nand U11724 (N_11724,N_6029,N_7816);
nor U11725 (N_11725,N_6762,N_7530);
or U11726 (N_11726,N_7292,N_6665);
or U11727 (N_11727,N_8523,N_7964);
or U11728 (N_11728,N_6342,N_6960);
nor U11729 (N_11729,N_6559,N_8892);
nand U11730 (N_11730,N_8269,N_7777);
and U11731 (N_11731,N_6319,N_7823);
and U11732 (N_11732,N_6200,N_8020);
or U11733 (N_11733,N_8734,N_7750);
xnor U11734 (N_11734,N_8059,N_6154);
or U11735 (N_11735,N_8539,N_6576);
and U11736 (N_11736,N_8415,N_7635);
nor U11737 (N_11737,N_8989,N_7692);
or U11738 (N_11738,N_7197,N_8540);
xor U11739 (N_11739,N_8638,N_7829);
nand U11740 (N_11740,N_6363,N_6213);
nor U11741 (N_11741,N_7213,N_8368);
or U11742 (N_11742,N_7650,N_7731);
nor U11743 (N_11743,N_8492,N_7067);
nand U11744 (N_11744,N_6034,N_8112);
or U11745 (N_11745,N_7839,N_7007);
and U11746 (N_11746,N_8562,N_8999);
nor U11747 (N_11747,N_7032,N_8673);
or U11748 (N_11748,N_7283,N_6604);
and U11749 (N_11749,N_8680,N_8441);
or U11750 (N_11750,N_6726,N_8910);
nand U11751 (N_11751,N_8973,N_6753);
nand U11752 (N_11752,N_8323,N_7200);
or U11753 (N_11753,N_8139,N_6579);
nand U11754 (N_11754,N_7422,N_6851);
and U11755 (N_11755,N_7823,N_6250);
or U11756 (N_11756,N_7448,N_8576);
nand U11757 (N_11757,N_8518,N_8859);
and U11758 (N_11758,N_6931,N_6125);
and U11759 (N_11759,N_6693,N_8305);
nand U11760 (N_11760,N_8403,N_8879);
nand U11761 (N_11761,N_6539,N_7279);
and U11762 (N_11762,N_8484,N_8273);
nor U11763 (N_11763,N_8540,N_8368);
and U11764 (N_11764,N_6466,N_7013);
and U11765 (N_11765,N_8261,N_6645);
and U11766 (N_11766,N_8991,N_6556);
or U11767 (N_11767,N_8936,N_7007);
or U11768 (N_11768,N_6640,N_8801);
nor U11769 (N_11769,N_8137,N_7793);
xnor U11770 (N_11770,N_8489,N_8533);
nor U11771 (N_11771,N_8407,N_8178);
or U11772 (N_11772,N_7813,N_7720);
and U11773 (N_11773,N_6288,N_8572);
and U11774 (N_11774,N_8810,N_8510);
nor U11775 (N_11775,N_7542,N_8547);
nand U11776 (N_11776,N_7687,N_8009);
nor U11777 (N_11777,N_7772,N_7868);
nor U11778 (N_11778,N_6694,N_6507);
or U11779 (N_11779,N_7390,N_8626);
or U11780 (N_11780,N_8019,N_7429);
and U11781 (N_11781,N_7045,N_6386);
and U11782 (N_11782,N_8465,N_6009);
nand U11783 (N_11783,N_7415,N_6076);
and U11784 (N_11784,N_7546,N_6164);
or U11785 (N_11785,N_7610,N_7105);
nand U11786 (N_11786,N_7821,N_7508);
and U11787 (N_11787,N_6240,N_7765);
nand U11788 (N_11788,N_8349,N_6664);
and U11789 (N_11789,N_8990,N_8525);
nor U11790 (N_11790,N_8649,N_7376);
or U11791 (N_11791,N_8604,N_8567);
and U11792 (N_11792,N_7705,N_6923);
nand U11793 (N_11793,N_6565,N_6816);
nand U11794 (N_11794,N_7618,N_6390);
nand U11795 (N_11795,N_7133,N_8534);
and U11796 (N_11796,N_6220,N_7119);
nor U11797 (N_11797,N_7471,N_7974);
nand U11798 (N_11798,N_7545,N_8887);
and U11799 (N_11799,N_7817,N_6650);
nand U11800 (N_11800,N_7772,N_6843);
or U11801 (N_11801,N_7076,N_6167);
nand U11802 (N_11802,N_6040,N_6266);
nand U11803 (N_11803,N_6231,N_7335);
and U11804 (N_11804,N_8823,N_8187);
or U11805 (N_11805,N_6319,N_8021);
nor U11806 (N_11806,N_7418,N_8326);
nor U11807 (N_11807,N_7743,N_6000);
and U11808 (N_11808,N_6208,N_6185);
and U11809 (N_11809,N_8982,N_6264);
and U11810 (N_11810,N_8596,N_7146);
xnor U11811 (N_11811,N_6667,N_6685);
or U11812 (N_11812,N_8318,N_7847);
and U11813 (N_11813,N_7907,N_8708);
or U11814 (N_11814,N_8134,N_6110);
nand U11815 (N_11815,N_7758,N_8651);
nand U11816 (N_11816,N_6758,N_6782);
nor U11817 (N_11817,N_8819,N_8362);
nor U11818 (N_11818,N_6824,N_7776);
and U11819 (N_11819,N_6591,N_7036);
nor U11820 (N_11820,N_8142,N_6343);
and U11821 (N_11821,N_6194,N_7798);
nand U11822 (N_11822,N_8894,N_8961);
or U11823 (N_11823,N_8965,N_6021);
xor U11824 (N_11824,N_8760,N_7324);
and U11825 (N_11825,N_7891,N_7476);
nor U11826 (N_11826,N_8286,N_7878);
nor U11827 (N_11827,N_7121,N_7234);
nand U11828 (N_11828,N_6723,N_6417);
or U11829 (N_11829,N_8936,N_8656);
nor U11830 (N_11830,N_7941,N_7989);
and U11831 (N_11831,N_8684,N_7973);
nand U11832 (N_11832,N_7588,N_8961);
nand U11833 (N_11833,N_6900,N_7865);
or U11834 (N_11834,N_6129,N_7364);
nand U11835 (N_11835,N_6660,N_6443);
nor U11836 (N_11836,N_8800,N_8609);
nor U11837 (N_11837,N_6022,N_7816);
or U11838 (N_11838,N_6324,N_7321);
nor U11839 (N_11839,N_8801,N_8661);
nand U11840 (N_11840,N_8289,N_7517);
or U11841 (N_11841,N_6733,N_7949);
nand U11842 (N_11842,N_8760,N_8595);
nand U11843 (N_11843,N_7277,N_6722);
nand U11844 (N_11844,N_6258,N_6645);
nor U11845 (N_11845,N_6293,N_6937);
nand U11846 (N_11846,N_6211,N_6373);
or U11847 (N_11847,N_8897,N_8312);
nand U11848 (N_11848,N_7059,N_7517);
and U11849 (N_11849,N_8727,N_6973);
and U11850 (N_11850,N_8397,N_6765);
nor U11851 (N_11851,N_8088,N_6391);
or U11852 (N_11852,N_7802,N_7394);
or U11853 (N_11853,N_8042,N_7690);
nand U11854 (N_11854,N_6217,N_6834);
and U11855 (N_11855,N_8742,N_7205);
and U11856 (N_11856,N_7295,N_7689);
xnor U11857 (N_11857,N_8819,N_6617);
or U11858 (N_11858,N_8650,N_8504);
and U11859 (N_11859,N_7667,N_8322);
or U11860 (N_11860,N_8372,N_7832);
or U11861 (N_11861,N_6168,N_7762);
and U11862 (N_11862,N_7363,N_7446);
or U11863 (N_11863,N_7097,N_7016);
xor U11864 (N_11864,N_6295,N_7299);
nand U11865 (N_11865,N_6404,N_7165);
nor U11866 (N_11866,N_8170,N_7815);
and U11867 (N_11867,N_7297,N_7905);
nor U11868 (N_11868,N_7355,N_8742);
or U11869 (N_11869,N_7678,N_6054);
or U11870 (N_11870,N_7780,N_7795);
nand U11871 (N_11871,N_6623,N_6129);
or U11872 (N_11872,N_6508,N_8398);
or U11873 (N_11873,N_7453,N_6828);
nor U11874 (N_11874,N_7697,N_8244);
nor U11875 (N_11875,N_6272,N_8089);
and U11876 (N_11876,N_6740,N_8012);
nand U11877 (N_11877,N_8360,N_7223);
or U11878 (N_11878,N_6643,N_7552);
nor U11879 (N_11879,N_8975,N_7421);
and U11880 (N_11880,N_6234,N_6400);
nand U11881 (N_11881,N_7544,N_8887);
or U11882 (N_11882,N_7854,N_8434);
or U11883 (N_11883,N_8574,N_8064);
and U11884 (N_11884,N_8772,N_6861);
or U11885 (N_11885,N_6264,N_7435);
nand U11886 (N_11886,N_7241,N_6953);
nand U11887 (N_11887,N_7509,N_7801);
nand U11888 (N_11888,N_6422,N_8620);
nand U11889 (N_11889,N_6079,N_6714);
nand U11890 (N_11890,N_8908,N_8468);
nand U11891 (N_11891,N_6096,N_6996);
nand U11892 (N_11892,N_7185,N_8961);
or U11893 (N_11893,N_6039,N_7591);
and U11894 (N_11894,N_6174,N_8401);
nor U11895 (N_11895,N_8988,N_6496);
nor U11896 (N_11896,N_6646,N_7975);
or U11897 (N_11897,N_7611,N_6513);
or U11898 (N_11898,N_8857,N_6369);
and U11899 (N_11899,N_8225,N_6946);
or U11900 (N_11900,N_7827,N_7995);
or U11901 (N_11901,N_8066,N_8579);
nand U11902 (N_11902,N_8187,N_6343);
nor U11903 (N_11903,N_6982,N_7183);
and U11904 (N_11904,N_8297,N_7485);
and U11905 (N_11905,N_8729,N_6812);
nor U11906 (N_11906,N_6136,N_8433);
and U11907 (N_11907,N_7680,N_6272);
and U11908 (N_11908,N_6824,N_8062);
and U11909 (N_11909,N_6833,N_6651);
and U11910 (N_11910,N_7740,N_8644);
nor U11911 (N_11911,N_8694,N_6909);
xnor U11912 (N_11912,N_8199,N_7853);
or U11913 (N_11913,N_8868,N_6419);
or U11914 (N_11914,N_8024,N_8063);
and U11915 (N_11915,N_6131,N_6465);
nor U11916 (N_11916,N_8118,N_8627);
or U11917 (N_11917,N_8754,N_6784);
or U11918 (N_11918,N_7205,N_7088);
or U11919 (N_11919,N_7003,N_8924);
nand U11920 (N_11920,N_8027,N_7223);
and U11921 (N_11921,N_8925,N_7976);
or U11922 (N_11922,N_7790,N_8745);
nor U11923 (N_11923,N_6240,N_7699);
nor U11924 (N_11924,N_6631,N_7574);
and U11925 (N_11925,N_6628,N_7048);
and U11926 (N_11926,N_7102,N_8245);
and U11927 (N_11927,N_6879,N_6405);
or U11928 (N_11928,N_6977,N_6456);
and U11929 (N_11929,N_7722,N_7975);
or U11930 (N_11930,N_8706,N_6017);
nand U11931 (N_11931,N_8884,N_8008);
nor U11932 (N_11932,N_8103,N_7394);
nor U11933 (N_11933,N_6388,N_6719);
and U11934 (N_11934,N_8269,N_7606);
nand U11935 (N_11935,N_7024,N_6917);
or U11936 (N_11936,N_8399,N_6945);
xnor U11937 (N_11937,N_8101,N_8226);
and U11938 (N_11938,N_6592,N_7569);
or U11939 (N_11939,N_7522,N_7006);
xor U11940 (N_11940,N_8043,N_7773);
nor U11941 (N_11941,N_7999,N_8135);
and U11942 (N_11942,N_7224,N_7054);
nor U11943 (N_11943,N_6875,N_7827);
and U11944 (N_11944,N_6927,N_7378);
nor U11945 (N_11945,N_6098,N_8184);
nor U11946 (N_11946,N_6479,N_7677);
or U11947 (N_11947,N_7260,N_8351);
and U11948 (N_11948,N_7503,N_8443);
and U11949 (N_11949,N_6599,N_8742);
or U11950 (N_11950,N_7032,N_8375);
nand U11951 (N_11951,N_6242,N_6430);
nand U11952 (N_11952,N_6109,N_8698);
nand U11953 (N_11953,N_7192,N_8099);
nand U11954 (N_11954,N_7183,N_7271);
nor U11955 (N_11955,N_7764,N_8207);
nand U11956 (N_11956,N_6034,N_6153);
and U11957 (N_11957,N_6186,N_8608);
nor U11958 (N_11958,N_7502,N_6270);
nor U11959 (N_11959,N_6019,N_8162);
or U11960 (N_11960,N_8450,N_7964);
or U11961 (N_11961,N_6895,N_8044);
and U11962 (N_11962,N_6802,N_8740);
or U11963 (N_11963,N_7152,N_8568);
nor U11964 (N_11964,N_7594,N_7856);
nand U11965 (N_11965,N_6817,N_8865);
and U11966 (N_11966,N_7529,N_6069);
or U11967 (N_11967,N_8650,N_7913);
and U11968 (N_11968,N_7743,N_6597);
nand U11969 (N_11969,N_7920,N_8788);
or U11970 (N_11970,N_8400,N_7955);
and U11971 (N_11971,N_7080,N_7371);
nor U11972 (N_11972,N_7349,N_8488);
or U11973 (N_11973,N_7976,N_8959);
nand U11974 (N_11974,N_7210,N_8380);
nor U11975 (N_11975,N_7341,N_8670);
nor U11976 (N_11976,N_8685,N_8543);
nand U11977 (N_11977,N_6008,N_6074);
nand U11978 (N_11978,N_8957,N_6517);
and U11979 (N_11979,N_8250,N_6435);
or U11980 (N_11980,N_8289,N_6392);
nor U11981 (N_11981,N_6247,N_7250);
nand U11982 (N_11982,N_6103,N_6863);
or U11983 (N_11983,N_7117,N_6928);
xnor U11984 (N_11984,N_7824,N_7259);
or U11985 (N_11985,N_6369,N_8287);
or U11986 (N_11986,N_7521,N_7875);
nand U11987 (N_11987,N_8075,N_7344);
nor U11988 (N_11988,N_7051,N_6602);
and U11989 (N_11989,N_6808,N_6103);
nand U11990 (N_11990,N_6218,N_7581);
and U11991 (N_11991,N_6479,N_7676);
or U11992 (N_11992,N_8075,N_7116);
and U11993 (N_11993,N_6898,N_8708);
or U11994 (N_11994,N_8930,N_6118);
or U11995 (N_11995,N_6010,N_6054);
and U11996 (N_11996,N_7719,N_8418);
nand U11997 (N_11997,N_8498,N_8120);
nand U11998 (N_11998,N_8254,N_7121);
or U11999 (N_11999,N_6695,N_8620);
nor U12000 (N_12000,N_10896,N_10623);
xor U12001 (N_12001,N_11487,N_10968);
or U12002 (N_12002,N_11334,N_9004);
nor U12003 (N_12003,N_10009,N_10384);
nand U12004 (N_12004,N_10396,N_9402);
nor U12005 (N_12005,N_11572,N_9432);
and U12006 (N_12006,N_11836,N_10912);
and U12007 (N_12007,N_11100,N_10350);
nand U12008 (N_12008,N_11856,N_11648);
xnor U12009 (N_12009,N_9870,N_10681);
or U12010 (N_12010,N_11419,N_11767);
or U12011 (N_12011,N_9816,N_9046);
nand U12012 (N_12012,N_10054,N_9990);
nand U12013 (N_12013,N_9273,N_10921);
nor U12014 (N_12014,N_11886,N_11101);
or U12015 (N_12015,N_9584,N_10686);
nor U12016 (N_12016,N_10892,N_9940);
or U12017 (N_12017,N_10819,N_11337);
nor U12018 (N_12018,N_9221,N_10514);
or U12019 (N_12019,N_10366,N_10327);
xor U12020 (N_12020,N_10421,N_10598);
nor U12021 (N_12021,N_9802,N_9744);
nand U12022 (N_12022,N_11874,N_10763);
and U12023 (N_12023,N_11335,N_11561);
nor U12024 (N_12024,N_9857,N_10390);
and U12025 (N_12025,N_11560,N_9727);
nand U12026 (N_12026,N_10594,N_10742);
nor U12027 (N_12027,N_9934,N_11197);
nor U12028 (N_12028,N_10096,N_11175);
or U12029 (N_12029,N_11557,N_10687);
nor U12030 (N_12030,N_9406,N_11440);
xor U12031 (N_12031,N_10380,N_11319);
or U12032 (N_12032,N_11899,N_10236);
nor U12033 (N_12033,N_10443,N_10342);
and U12034 (N_12034,N_10472,N_11852);
nand U12035 (N_12035,N_10886,N_10745);
nand U12036 (N_12036,N_11643,N_10126);
and U12037 (N_12037,N_11609,N_10647);
or U12038 (N_12038,N_9707,N_9070);
nor U12039 (N_12039,N_10949,N_9813);
nand U12040 (N_12040,N_9886,N_10489);
nor U12041 (N_12041,N_11592,N_10531);
and U12042 (N_12042,N_9709,N_11739);
and U12043 (N_12043,N_9010,N_10964);
or U12044 (N_12044,N_10442,N_10908);
or U12045 (N_12045,N_11356,N_11107);
or U12046 (N_12046,N_10279,N_9248);
or U12047 (N_12047,N_10125,N_9664);
nor U12048 (N_12048,N_10178,N_10501);
and U12049 (N_12049,N_9423,N_9941);
nor U12050 (N_12050,N_10631,N_9349);
or U12051 (N_12051,N_10170,N_11841);
and U12052 (N_12052,N_11503,N_10382);
nand U12053 (N_12053,N_10294,N_9550);
nand U12054 (N_12054,N_10065,N_9906);
and U12055 (N_12055,N_10665,N_11033);
nor U12056 (N_12056,N_10171,N_9877);
nor U12057 (N_12057,N_11127,N_11629);
or U12058 (N_12058,N_10369,N_10247);
or U12059 (N_12059,N_11584,N_11153);
and U12060 (N_12060,N_9387,N_11928);
nand U12061 (N_12061,N_11243,N_11695);
and U12062 (N_12062,N_11099,N_10099);
nand U12063 (N_12063,N_9102,N_11714);
nand U12064 (N_12064,N_9189,N_10420);
nor U12065 (N_12065,N_11908,N_10910);
nand U12066 (N_12066,N_9170,N_10441);
nor U12067 (N_12067,N_10930,N_10156);
nand U12068 (N_12068,N_9195,N_9056);
nand U12069 (N_12069,N_11800,N_9413);
nand U12070 (N_12070,N_9723,N_9117);
xnor U12071 (N_12071,N_9401,N_9355);
nand U12072 (N_12072,N_11895,N_11855);
nand U12073 (N_12073,N_10504,N_10363);
or U12074 (N_12074,N_9122,N_10761);
nor U12075 (N_12075,N_9521,N_10856);
nor U12076 (N_12076,N_9607,N_10884);
and U12077 (N_12077,N_9927,N_11376);
and U12078 (N_12078,N_9210,N_9784);
nor U12079 (N_12079,N_10608,N_11486);
and U12080 (N_12080,N_11192,N_9568);
or U12081 (N_12081,N_10164,N_9683);
or U12082 (N_12082,N_9446,N_9951);
nand U12083 (N_12083,N_9515,N_9205);
or U12084 (N_12084,N_9147,N_11513);
and U12085 (N_12085,N_9471,N_11881);
nor U12086 (N_12086,N_9220,N_9800);
nand U12087 (N_12087,N_10121,N_11047);
or U12088 (N_12088,N_11461,N_9576);
xnor U12089 (N_12089,N_11581,N_11422);
nor U12090 (N_12090,N_11317,N_11273);
nor U12091 (N_12091,N_9352,N_10597);
and U12092 (N_12092,N_9632,N_9790);
or U12093 (N_12093,N_11787,N_11129);
nand U12094 (N_12094,N_10796,N_10337);
nor U12095 (N_12095,N_11237,N_9234);
nand U12096 (N_12096,N_9995,N_10020);
or U12097 (N_12097,N_11046,N_10061);
and U12098 (N_12098,N_11193,N_9315);
nand U12099 (N_12099,N_11857,N_10640);
or U12100 (N_12100,N_11601,N_10264);
and U12101 (N_12101,N_10655,N_10852);
and U12102 (N_12102,N_10979,N_11362);
xnor U12103 (N_12103,N_10301,N_11270);
nand U12104 (N_12104,N_11141,N_10188);
and U12105 (N_12105,N_10496,N_11843);
nor U12106 (N_12106,N_10223,N_9980);
nor U12107 (N_12107,N_9998,N_10593);
nand U12108 (N_12108,N_9326,N_10580);
or U12109 (N_12109,N_11035,N_9517);
or U12110 (N_12110,N_9575,N_11331);
or U12111 (N_12111,N_9144,N_9611);
nor U12112 (N_12112,N_10603,N_9811);
and U12113 (N_12113,N_10016,N_9883);
or U12114 (N_12114,N_9682,N_11671);
nand U12115 (N_12115,N_10941,N_10971);
xnor U12116 (N_12116,N_10833,N_9809);
and U12117 (N_12117,N_11730,N_10877);
or U12118 (N_12118,N_9215,N_11490);
or U12119 (N_12119,N_9781,N_9474);
nor U12120 (N_12120,N_9845,N_9725);
xor U12121 (N_12121,N_9614,N_10660);
or U12122 (N_12122,N_11533,N_11640);
nand U12123 (N_12123,N_10999,N_11736);
nor U12124 (N_12124,N_9093,N_11201);
nand U12125 (N_12125,N_9443,N_10516);
and U12126 (N_12126,N_9898,N_10544);
nand U12127 (N_12127,N_10333,N_10142);
and U12128 (N_12128,N_9097,N_10173);
and U12129 (N_12129,N_9871,N_11240);
and U12130 (N_12130,N_11016,N_11027);
nand U12131 (N_12131,N_9271,N_10253);
or U12132 (N_12132,N_10585,N_9492);
or U12133 (N_12133,N_11447,N_10144);
or U12134 (N_12134,N_9291,N_9452);
nand U12135 (N_12135,N_10642,N_9211);
or U12136 (N_12136,N_9403,N_9253);
nand U12137 (N_12137,N_9282,N_10860);
or U12138 (N_12138,N_10521,N_10050);
nor U12139 (N_12139,N_10936,N_9854);
nand U12140 (N_12140,N_10809,N_11302);
and U12141 (N_12141,N_11512,N_11316);
or U12142 (N_12142,N_10602,N_10071);
nor U12143 (N_12143,N_11116,N_9645);
or U12144 (N_12144,N_11931,N_11187);
nand U12145 (N_12145,N_10703,N_11683);
nand U12146 (N_12146,N_10210,N_11795);
nand U12147 (N_12147,N_9184,N_11920);
nor U12148 (N_12148,N_9982,N_10181);
nor U12149 (N_12149,N_9101,N_9742);
or U12150 (N_12150,N_11410,N_9848);
and U12151 (N_12151,N_9174,N_10952);
and U12152 (N_12152,N_11936,N_10619);
or U12153 (N_12153,N_9063,N_11670);
nand U12154 (N_12154,N_9157,N_11799);
nor U12155 (N_12155,N_10175,N_11733);
and U12156 (N_12156,N_9141,N_9656);
nor U12157 (N_12157,N_11152,N_10747);
nor U12158 (N_12158,N_11975,N_9755);
and U12159 (N_12159,N_11235,N_10548);
and U12160 (N_12160,N_9098,N_9180);
nor U12161 (N_12161,N_11021,N_10041);
nor U12162 (N_12162,N_10756,N_9372);
or U12163 (N_12163,N_10826,N_10627);
or U12164 (N_12164,N_11682,N_11217);
and U12165 (N_12165,N_11250,N_9735);
nor U12166 (N_12166,N_10300,N_9922);
nor U12167 (N_12167,N_9267,N_10755);
and U12168 (N_12168,N_9398,N_10101);
nor U12169 (N_12169,N_9503,N_10733);
and U12170 (N_12170,N_9137,N_9060);
or U12171 (N_12171,N_11300,N_11357);
nor U12172 (N_12172,N_9701,N_11173);
or U12173 (N_12173,N_9260,N_11970);
or U12174 (N_12174,N_10292,N_9684);
nand U12175 (N_12175,N_9539,N_9670);
nand U12176 (N_12176,N_10015,N_9936);
nor U12177 (N_12177,N_9767,N_10974);
nand U12178 (N_12178,N_10083,N_10078);
and U12179 (N_12179,N_10572,N_9868);
and U12180 (N_12180,N_9777,N_11114);
or U12181 (N_12181,N_9047,N_10255);
and U12182 (N_12182,N_10351,N_11451);
and U12183 (N_12183,N_10538,N_9397);
nor U12184 (N_12184,N_9564,N_10958);
and U12185 (N_12185,N_11408,N_9694);
and U12186 (N_12186,N_9208,N_9703);
or U12187 (N_12187,N_9495,N_11806);
or U12188 (N_12188,N_9400,N_11900);
nand U12189 (N_12189,N_10866,N_9597);
and U12190 (N_12190,N_9009,N_11721);
nand U12191 (N_12191,N_11511,N_11504);
and U12192 (N_12192,N_10764,N_9776);
xnor U12193 (N_12193,N_10996,N_10663);
or U12194 (N_12194,N_10618,N_10639);
or U12195 (N_12195,N_9178,N_10717);
or U12196 (N_12196,N_11722,N_11922);
and U12197 (N_12197,N_11759,N_10330);
and U12198 (N_12198,N_11232,N_9194);
nand U12199 (N_12199,N_9407,N_11760);
and U12200 (N_12200,N_10124,N_11359);
nor U12201 (N_12201,N_10452,N_10191);
xor U12202 (N_12202,N_9015,N_9792);
or U12203 (N_12203,N_9064,N_10295);
nand U12204 (N_12204,N_11271,N_11200);
or U12205 (N_12205,N_9499,N_10708);
or U12206 (N_12206,N_10069,N_11876);
nand U12207 (N_12207,N_11860,N_10671);
or U12208 (N_12208,N_10937,N_10743);
or U12209 (N_12209,N_11977,N_11929);
and U12210 (N_12210,N_11915,N_10482);
nor U12211 (N_12211,N_9510,N_10832);
nor U12212 (N_12212,N_9788,N_10878);
and U12213 (N_12213,N_9615,N_11205);
and U12214 (N_12214,N_11870,N_10495);
and U12215 (N_12215,N_10837,N_10468);
nand U12216 (N_12216,N_9625,N_9241);
nand U12217 (N_12217,N_9544,N_10803);
nand U12218 (N_12218,N_9609,N_11530);
xor U12219 (N_12219,N_11594,N_10929);
nand U12220 (N_12220,N_10407,N_9223);
nand U12221 (N_12221,N_10997,N_10129);
nor U12222 (N_12222,N_10824,N_11402);
or U12223 (N_12223,N_11780,N_11961);
or U12224 (N_12224,N_11123,N_9095);
or U12225 (N_12225,N_9172,N_10356);
nor U12226 (N_12226,N_9022,N_11496);
nor U12227 (N_12227,N_9573,N_9970);
nor U12228 (N_12228,N_10477,N_11219);
nand U12229 (N_12229,N_9890,N_11040);
or U12230 (N_12230,N_11838,N_9572);
nand U12231 (N_12231,N_11934,N_9774);
and U12232 (N_12232,N_11276,N_11091);
nand U12233 (N_12233,N_9496,N_11311);
nand U12234 (N_12234,N_9066,N_9043);
and U12235 (N_12235,N_11108,N_9738);
or U12236 (N_12236,N_9786,N_10036);
and U12237 (N_12237,N_10527,N_10274);
nor U12238 (N_12238,N_9294,N_11207);
nor U12239 (N_12239,N_9014,N_9981);
and U12240 (N_12240,N_10726,N_9337);
or U12241 (N_12241,N_10995,N_11326);
and U12242 (N_12242,N_11269,N_10749);
xnor U12243 (N_12243,N_9266,N_11313);
nor U12244 (N_12244,N_10409,N_9479);
or U12245 (N_12245,N_10141,N_10638);
and U12246 (N_12246,N_9239,N_9449);
and U12247 (N_12247,N_11966,N_10123);
or U12248 (N_12248,N_10862,N_11738);
or U12249 (N_12249,N_10307,N_9287);
nand U12250 (N_12250,N_10524,N_10272);
nor U12251 (N_12251,N_10375,N_9866);
nand U12252 (N_12252,N_11549,N_9276);
nand U12253 (N_12253,N_10143,N_11679);
or U12254 (N_12254,N_10791,N_9975);
nor U12255 (N_12255,N_10221,N_11524);
or U12256 (N_12256,N_11927,N_11517);
nor U12257 (N_12257,N_9916,N_10578);
and U12258 (N_12258,N_11887,N_10925);
or U12259 (N_12259,N_10656,N_11343);
and U12260 (N_12260,N_11167,N_11850);
or U12261 (N_12261,N_9080,N_11073);
and U12262 (N_12262,N_11399,N_11652);
nor U12263 (N_12263,N_11083,N_9290);
nor U12264 (N_12264,N_9460,N_11994);
nand U12265 (N_12265,N_11398,N_11568);
and U12266 (N_12266,N_11778,N_9750);
or U12267 (N_12267,N_11784,N_11480);
or U12268 (N_12268,N_10177,N_11412);
nand U12269 (N_12269,N_11206,N_11186);
or U12270 (N_12270,N_9263,N_10336);
and U12271 (N_12271,N_9347,N_9518);
or U12272 (N_12272,N_9123,N_10880);
nor U12273 (N_12273,N_10725,N_11770);
nand U12274 (N_12274,N_10739,N_10182);
or U12275 (N_12275,N_11805,N_10648);
nand U12276 (N_12276,N_9148,N_9605);
nand U12277 (N_12277,N_11158,N_9236);
or U12278 (N_12278,N_10817,N_11550);
or U12279 (N_12279,N_11904,N_10969);
or U12280 (N_12280,N_9209,N_9278);
nand U12281 (N_12281,N_9894,N_10984);
nand U12282 (N_12282,N_11665,N_11891);
and U12283 (N_12283,N_11545,N_10471);
and U12284 (N_12284,N_10372,N_9391);
and U12285 (N_12285,N_9847,N_10683);
nor U12286 (N_12286,N_11942,N_10368);
nor U12287 (N_12287,N_10397,N_11605);
nor U12288 (N_12288,N_11325,N_10289);
nor U12289 (N_12289,N_9646,N_9595);
nand U12290 (N_12290,N_11840,N_11905);
nor U12291 (N_12291,N_9902,N_11124);
and U12292 (N_12292,N_9453,N_11148);
nor U12293 (N_12293,N_10435,N_10208);
and U12294 (N_12294,N_9280,N_11074);
or U12295 (N_12295,N_10026,N_9578);
nand U12296 (N_12296,N_9021,N_9803);
and U12297 (N_12297,N_9907,N_10373);
nor U12298 (N_12298,N_10954,N_9011);
nand U12299 (N_12299,N_11468,N_11688);
or U12300 (N_12300,N_9306,N_11514);
xnor U12301 (N_12301,N_9556,N_10304);
nand U12302 (N_12302,N_10576,N_10857);
nand U12303 (N_12303,N_11731,N_9024);
or U12304 (N_12304,N_11969,N_10712);
and U12305 (N_12305,N_11898,N_11241);
or U12306 (N_12306,N_10486,N_9500);
nor U12307 (N_12307,N_9965,N_9341);
nand U12308 (N_12308,N_9904,N_11725);
and U12309 (N_12309,N_11383,N_11157);
and U12310 (N_12310,N_10159,N_11639);
and U12311 (N_12311,N_11110,N_10270);
nor U12312 (N_12312,N_9366,N_9244);
nor U12313 (N_12313,N_11754,N_11715);
and U12314 (N_12314,N_11813,N_9062);
nor U12315 (N_12315,N_11195,N_10163);
nor U12316 (N_12316,N_10894,N_9476);
nand U12317 (N_12317,N_11510,N_11819);
and U12318 (N_12318,N_9143,N_11950);
and U12319 (N_12319,N_10560,N_10515);
nand U12320 (N_12320,N_9431,N_10268);
or U12321 (N_12321,N_11828,N_11830);
or U12322 (N_12322,N_9509,N_11793);
or U12323 (N_12323,N_10775,N_11010);
nand U12324 (N_12324,N_10714,N_11833);
and U12325 (N_12325,N_10469,N_10924);
or U12326 (N_12326,N_11626,N_10861);
and U12327 (N_12327,N_9218,N_11491);
xnor U12328 (N_12328,N_11299,N_11143);
nor U12329 (N_12329,N_10034,N_11582);
nand U12330 (N_12330,N_11687,N_11242);
and U12331 (N_12331,N_11776,N_11464);
nand U12332 (N_12332,N_11102,N_9841);
or U12333 (N_12333,N_11538,N_9963);
and U12334 (N_12334,N_10447,N_11467);
nor U12335 (N_12335,N_9569,N_11038);
nand U12336 (N_12336,N_10014,N_11354);
nand U12337 (N_12337,N_11740,N_9115);
nand U12338 (N_12338,N_11603,N_9462);
nor U12339 (N_12339,N_11689,N_10115);
or U12340 (N_12340,N_9613,N_11749);
nand U12341 (N_12341,N_11015,N_11477);
nor U12342 (N_12342,N_11937,N_11223);
nor U12343 (N_12343,N_11735,N_10260);
nor U12344 (N_12344,N_9171,N_11863);
nor U12345 (N_12345,N_9749,N_10012);
and U12346 (N_12346,N_11763,N_9103);
nor U12347 (N_12347,N_11052,N_10398);
or U12348 (N_12348,N_11796,N_9959);
nand U12349 (N_12349,N_9654,N_9514);
and U12350 (N_12350,N_10564,N_9549);
or U12351 (N_12351,N_10781,N_10296);
or U12352 (N_12352,N_11846,N_9183);
nand U12353 (N_12353,N_10475,N_9869);
nor U12354 (N_12354,N_11726,N_10508);
nand U12355 (N_12355,N_9311,N_9477);
nand U12356 (N_12356,N_9344,N_11750);
and U12357 (N_12357,N_10573,N_10762);
nand U12358 (N_12358,N_9835,N_10137);
or U12359 (N_12359,N_9444,N_9938);
and U12360 (N_12360,N_9418,N_9393);
nand U12361 (N_12361,N_9833,N_9801);
and U12362 (N_12362,N_9363,N_10613);
nor U12363 (N_12363,N_10068,N_11498);
xnor U12364 (N_12364,N_11161,N_11065);
and U12365 (N_12365,N_11154,N_10644);
nor U12366 (N_12366,N_11439,N_10821);
and U12367 (N_12367,N_9036,N_10519);
or U12368 (N_12368,N_9298,N_9677);
and U12369 (N_12369,N_10520,N_9931);
or U12370 (N_12370,N_9256,N_9169);
nor U12371 (N_12371,N_9765,N_11347);
or U12372 (N_12372,N_10339,N_11087);
and U12373 (N_12373,N_11281,N_10040);
and U12374 (N_12374,N_10353,N_10157);
nand U12375 (N_12375,N_9222,N_10694);
nand U12376 (N_12376,N_9483,N_11132);
or U12377 (N_12377,N_11711,N_10919);
nor U12378 (N_12378,N_9913,N_9330);
xor U12379 (N_12379,N_9561,N_10523);
and U12380 (N_12380,N_9988,N_11309);
and U12381 (N_12381,N_11400,N_11867);
or U12382 (N_12382,N_9269,N_11675);
xnor U12383 (N_12383,N_11879,N_9130);
nand U12384 (N_12384,N_10591,N_10891);
nand U12385 (N_12385,N_9016,N_11086);
and U12386 (N_12386,N_11667,N_9292);
nand U12387 (N_12387,N_10771,N_9506);
nor U12388 (N_12388,N_10875,N_9384);
and U12389 (N_12389,N_10847,N_11164);
nor U12390 (N_12390,N_11017,N_9771);
or U12391 (N_12391,N_9649,N_11792);
or U12392 (N_12392,N_10556,N_9810);
or U12393 (N_12393,N_11983,N_10211);
nand U12394 (N_12394,N_11989,N_10321);
nand U12395 (N_12395,N_11231,N_11284);
or U12396 (N_12396,N_10415,N_9971);
nand U12397 (N_12397,N_11142,N_10645);
nor U12398 (N_12398,N_10830,N_9643);
or U12399 (N_12399,N_10309,N_10674);
nor U12400 (N_12400,N_11475,N_11213);
or U12401 (N_12401,N_10865,N_9381);
nand U12402 (N_12402,N_9695,N_10579);
or U12403 (N_12403,N_10478,N_10535);
nand U12404 (N_12404,N_11960,N_10432);
and U12405 (N_12405,N_11310,N_10285);
nand U12406 (N_12406,N_9603,N_11072);
nor U12407 (N_12407,N_9702,N_9919);
xor U12408 (N_12408,N_9405,N_11471);
nand U12409 (N_12409,N_10414,N_10252);
or U12410 (N_12410,N_11542,N_11563);
nand U12411 (N_12411,N_11368,N_9120);
or U12412 (N_12412,N_10165,N_11914);
xor U12413 (N_12413,N_11972,N_11764);
nor U12414 (N_12414,N_10231,N_10804);
or U12415 (N_12415,N_11394,N_10042);
and U12416 (N_12416,N_10206,N_10058);
or U12417 (N_12417,N_10731,N_10565);
nor U12418 (N_12418,N_10960,N_9528);
nor U12419 (N_12419,N_11162,N_9668);
xnor U12420 (N_12420,N_10750,N_10760);
nor U12421 (N_12421,N_10198,N_10909);
or U12422 (N_12422,N_11616,N_9125);
or U12423 (N_12423,N_10951,N_10777);
nand U12424 (N_12424,N_10690,N_9068);
nor U12425 (N_12425,N_11199,N_9259);
or U12426 (N_12426,N_9834,N_11495);
or U12427 (N_12427,N_10596,N_11214);
nor U12428 (N_12428,N_9823,N_9301);
and U12429 (N_12429,N_9849,N_10013);
nor U12430 (N_12430,N_9574,N_11808);
or U12431 (N_12431,N_11979,N_11460);
and U12432 (N_12432,N_11117,N_9438);
or U12433 (N_12433,N_11058,N_11527);
nor U12434 (N_12434,N_10753,N_9339);
and U12435 (N_12435,N_9224,N_10533);
nor U12436 (N_12436,N_9756,N_9012);
and U12437 (N_12437,N_11168,N_11098);
nor U12438 (N_12438,N_10149,N_10217);
nand U12439 (N_12439,N_11505,N_10055);
or U12440 (N_12440,N_10216,N_10147);
nor U12441 (N_12441,N_11777,N_9524);
nand U12442 (N_12442,N_10870,N_10453);
xnor U12443 (N_12443,N_11336,N_11022);
xnor U12444 (N_12444,N_10248,N_11554);
nor U12445 (N_12445,N_10479,N_11734);
and U12446 (N_12446,N_10732,N_11179);
or U12447 (N_12447,N_11203,N_11441);
nand U12448 (N_12448,N_10766,N_11834);
or U12449 (N_12449,N_10662,N_9893);
nor U12450 (N_12450,N_11432,N_10389);
and U12451 (N_12451,N_11121,N_9262);
or U12452 (N_12452,N_10340,N_9053);
or U12453 (N_12453,N_9875,N_9176);
or U12454 (N_12454,N_10679,N_10239);
nand U12455 (N_12455,N_9075,N_10668);
nand U12456 (N_12456,N_9454,N_11463);
nand U12457 (N_12457,N_11188,N_11658);
nand U12458 (N_12458,N_9754,N_10800);
or U12459 (N_12459,N_10583,N_11246);
nand U12460 (N_12460,N_11272,N_10953);
nor U12461 (N_12461,N_11637,N_11096);
or U12462 (N_12462,N_9592,N_9678);
or U12463 (N_12463,N_11973,N_10172);
nor U12464 (N_12464,N_9693,N_9567);
and U12465 (N_12465,N_11570,N_9589);
nor U12466 (N_12466,N_9559,N_10823);
and U12467 (N_12467,N_9031,N_9563);
nand U12468 (N_12468,N_10035,N_11133);
nand U12469 (N_12469,N_10428,N_10305);
nand U12470 (N_12470,N_9037,N_11562);
or U12471 (N_12471,N_11955,N_9129);
and U12472 (N_12472,N_9861,N_10916);
nand U12473 (N_12473,N_10155,N_11350);
and U12474 (N_12474,N_9554,N_10493);
nor U12475 (N_12475,N_10972,N_9994);
nand U12476 (N_12476,N_11699,N_11516);
or U12477 (N_12477,N_11662,N_11364);
and U12478 (N_12478,N_11621,N_10704);
and U12479 (N_12479,N_11267,N_10431);
nor U12480 (N_12480,N_9579,N_11174);
or U12481 (N_12481,N_11919,N_11000);
nand U12482 (N_12482,N_10798,N_11897);
nand U12483 (N_12483,N_11034,N_10007);
or U12484 (N_12484,N_9937,N_11144);
nand U12485 (N_12485,N_10883,N_9411);
or U12486 (N_12486,N_9307,N_9162);
nor U12487 (N_12487,N_10840,N_11421);
or U12488 (N_12488,N_9612,N_10835);
nor U12489 (N_12489,N_11064,N_10240);
and U12490 (N_12490,N_10251,N_10652);
or U12491 (N_12491,N_9793,N_9340);
and U12492 (N_12492,N_11607,N_11810);
xor U12493 (N_12493,N_9083,N_10624);
and U12494 (N_12494,N_10989,N_10476);
and U12495 (N_12495,N_10105,N_11622);
or U12496 (N_12496,N_9316,N_9134);
nor U12497 (N_12497,N_11506,N_9389);
nand U12498 (N_12498,N_11059,N_11367);
or U12499 (N_12499,N_11424,N_11413);
or U12500 (N_12500,N_11277,N_9775);
nor U12501 (N_12501,N_11565,N_11558);
or U12502 (N_12502,N_10310,N_10215);
and U12503 (N_12503,N_9762,N_11756);
nor U12504 (N_12504,N_10903,N_10895);
and U12505 (N_12505,N_9055,N_9714);
or U12506 (N_12506,N_11965,N_10027);
or U12507 (N_12507,N_10567,N_10454);
nand U12508 (N_12508,N_11865,N_9986);
nand U12509 (N_12509,N_11140,N_10053);
or U12510 (N_12510,N_9412,N_10626);
nor U12511 (N_12511,N_10440,N_9382);
nand U12512 (N_12512,N_10926,N_10284);
or U12513 (N_12513,N_10754,N_9160);
and U12514 (N_12514,N_11888,N_9289);
and U12515 (N_12515,N_10072,N_11004);
xnor U12516 (N_12516,N_11328,N_9752);
and U12517 (N_12517,N_10994,N_10405);
nand U12518 (N_12518,N_9392,N_9577);
nand U12519 (N_12519,N_10349,N_11280);
nor U12520 (N_12520,N_9831,N_9308);
nand U12521 (N_12521,N_9914,N_9268);
nand U12522 (N_12522,N_9672,N_9946);
or U12523 (N_12523,N_11753,N_11858);
nor U12524 (N_12524,N_10106,N_9206);
or U12525 (N_12525,N_9715,N_10838);
and U12526 (N_12526,N_11946,N_9486);
and U12527 (N_12527,N_11085,N_10620);
or U12528 (N_12528,N_9192,N_9909);
and U12529 (N_12529,N_11062,N_11171);
or U12530 (N_12530,N_9791,N_9606);
xor U12531 (N_12531,N_11624,N_11783);
nand U12532 (N_12532,N_10818,N_11508);
and U12533 (N_12533,N_9964,N_11448);
nor U12534 (N_12534,N_9779,N_9111);
or U12535 (N_12535,N_10812,N_10180);
nand U12536 (N_12536,N_10168,N_10059);
and U12537 (N_12537,N_10186,N_10370);
xnor U12538 (N_12538,N_10427,N_9652);
nor U12539 (N_12539,N_10424,N_11427);
and U12540 (N_12540,N_10610,N_10112);
or U12541 (N_12541,N_9071,N_9003);
xor U12542 (N_12542,N_11431,N_9537);
and U12543 (N_12543,N_9487,N_10458);
or U12544 (N_12544,N_9706,N_9846);
and U12545 (N_12545,N_9651,N_9832);
nand U12546 (N_12546,N_9265,N_10128);
nor U12547 (N_12547,N_9571,N_9820);
nand U12548 (N_12548,N_10158,N_10352);
and U12549 (N_12549,N_11921,N_9481);
and U12550 (N_12550,N_11285,N_10494);
and U12551 (N_12551,N_10258,N_11048);
nor U12552 (N_12552,N_11669,N_9852);
nor U12553 (N_12553,N_9842,N_11312);
or U12554 (N_12554,N_11437,N_9357);
or U12555 (N_12555,N_9953,N_9050);
or U12556 (N_12556,N_9979,N_10094);
or U12557 (N_12557,N_11916,N_9182);
and U12558 (N_12558,N_10943,N_10004);
nand U12559 (N_12559,N_10161,N_9185);
nor U12560 (N_12560,N_9458,N_9320);
or U12561 (N_12561,N_11839,N_10699);
and U12562 (N_12562,N_10507,N_10324);
or U12563 (N_12563,N_9588,N_11094);
or U12564 (N_12564,N_10023,N_11901);
and U12565 (N_12565,N_10491,N_9351);
nor U12566 (N_12566,N_9993,N_10103);
and U12567 (N_12567,N_9859,N_10082);
or U12568 (N_12568,N_10911,N_11330);
nand U12569 (N_12569,N_11952,N_11138);
nor U12570 (N_12570,N_9478,N_9029);
or U12571 (N_12571,N_9030,N_10335);
nand U12572 (N_12572,N_9167,N_9041);
nor U12573 (N_12573,N_11837,N_9660);
or U12574 (N_12574,N_11379,N_9566);
or U12575 (N_12575,N_11084,N_11845);
or U12576 (N_12576,N_9475,N_10906);
nor U12577 (N_12577,N_11656,N_10807);
and U12578 (N_12578,N_11691,N_10361);
or U12579 (N_12579,N_11385,N_11885);
nand U12580 (N_12580,N_11718,N_10387);
or U12581 (N_12581,N_10898,N_11588);
or U12582 (N_12582,N_10485,N_10343);
xnor U12583 (N_12583,N_10359,N_11822);
nor U12584 (N_12584,N_10568,N_10212);
xor U12585 (N_12585,N_10500,N_9395);
nand U12586 (N_12586,N_9885,N_9226);
nor U12587 (N_12587,N_10077,N_9168);
and U12588 (N_12588,N_11801,N_11615);
nor U12589 (N_12589,N_9498,N_9324);
nand U12590 (N_12590,N_9892,N_9836);
nor U12591 (N_12591,N_9135,N_9704);
and U12592 (N_12592,N_10417,N_11847);
or U12593 (N_12593,N_11661,N_10131);
and U12594 (N_12594,N_10685,N_9976);
and U12595 (N_12595,N_10130,N_10904);
and U12596 (N_12596,N_11802,N_11353);
and U12597 (N_12597,N_9371,N_10630);
nor U12598 (N_12598,N_11345,N_9284);
and U12599 (N_12599,N_11469,N_10680);
or U12600 (N_12600,N_9439,N_10772);
or U12601 (N_12601,N_10283,N_10234);
nor U12602 (N_12602,N_10220,N_9932);
or U12603 (N_12603,N_9420,N_9631);
xor U12604 (N_12604,N_10831,N_10982);
and U12605 (N_12605,N_10374,N_10200);
nor U12606 (N_12606,N_11552,N_10811);
and U12607 (N_12607,N_10649,N_10902);
nor U12608 (N_12608,N_10697,N_9376);
and U12609 (N_12609,N_10993,N_9150);
nor U12610 (N_12610,N_10139,N_10269);
nand U12611 (N_12611,N_10965,N_9018);
nand U12612 (N_12612,N_9061,N_9133);
or U12613 (N_12613,N_9367,N_9818);
nand U12614 (N_12614,N_10331,N_9491);
and U12615 (N_12615,N_10550,N_9620);
xor U12616 (N_12616,N_9377,N_10541);
nor U12617 (N_12617,N_11297,N_10117);
or U12618 (N_12618,N_10057,N_9532);
or U12619 (N_12619,N_10410,N_10646);
nor U12620 (N_12620,N_11428,N_9548);
and U12621 (N_12621,N_9346,N_11208);
or U12622 (N_12622,N_10634,N_10488);
and U12623 (N_12623,N_9051,N_11602);
nand U12624 (N_12624,N_9100,N_11737);
and U12625 (N_12625,N_9669,N_11902);
and U12626 (N_12626,N_9729,N_11497);
or U12627 (N_12627,N_10379,N_10888);
nor U12628 (N_12628,N_10376,N_10189);
and U12629 (N_12629,N_11990,N_10322);
or U12630 (N_12630,N_11623,N_11252);
nor U12631 (N_12631,N_9764,N_11848);
nand U12632 (N_12632,N_9028,N_10218);
and U12633 (N_12633,N_9608,N_10510);
and U12634 (N_12634,N_10214,N_10882);
nor U12635 (N_12635,N_10066,N_11149);
nand U12636 (N_12636,N_11445,N_10092);
nor U12637 (N_12637,N_10086,N_11708);
or U12638 (N_12638,N_11647,N_9113);
or U12639 (N_12639,N_9335,N_9699);
nand U12640 (N_12640,N_9634,N_10546);
nand U12641 (N_12641,N_11396,N_9593);
and U12642 (N_12642,N_11959,N_11198);
nor U12643 (N_12643,N_9687,N_10010);
nand U12644 (N_12644,N_10774,N_11135);
nand U12645 (N_12645,N_9887,N_10893);
nor U12646 (N_12646,N_9124,N_9466);
or U12647 (N_12647,N_9952,N_10942);
nand U12648 (N_12648,N_10918,N_11372);
nor U12649 (N_12649,N_10616,N_9535);
and U12650 (N_12650,N_11056,N_11216);
and U12651 (N_12651,N_9586,N_10768);
and U12652 (N_12652,N_11455,N_9596);
and U12653 (N_12653,N_10632,N_11698);
and U12654 (N_12654,N_10418,N_10262);
or U12655 (N_12655,N_9928,N_11097);
nor U12656 (N_12656,N_11803,N_11892);
xnor U12657 (N_12657,N_10509,N_11092);
and U12658 (N_12658,N_9686,N_9052);
nor U12659 (N_12659,N_10899,N_10633);
or U12660 (N_12660,N_11366,N_11011);
nor U12661 (N_12661,N_10625,N_9583);
nand U12662 (N_12662,N_11710,N_10371);
nor U12663 (N_12663,N_11939,N_10905);
nor U12664 (N_12664,N_11707,N_9505);
or U12665 (N_12665,N_10102,N_10928);
nand U12666 (N_12666,N_11314,N_9383);
or U12667 (N_12667,N_10869,N_10243);
nand U12668 (N_12668,N_10028,N_10466);
nor U12669 (N_12669,N_9880,N_9587);
or U12670 (N_12670,N_9375,N_9516);
and U12671 (N_12671,N_9110,N_9149);
or U12672 (N_12672,N_9048,N_10746);
and U12673 (N_12673,N_9726,N_9163);
nor U12674 (N_12674,N_10332,N_10605);
or U12675 (N_12675,N_11262,N_9821);
and U12676 (N_12676,N_11388,N_11211);
and U12677 (N_12677,N_10621,N_9839);
or U12678 (N_12678,N_9570,N_9585);
or U12679 (N_12679,N_10923,N_11709);
or U12680 (N_12680,N_11080,N_11697);
nor U12681 (N_12681,N_11417,N_11355);
and U12682 (N_12682,N_9722,N_10983);
and U12683 (N_12683,N_9644,N_10022);
and U12684 (N_12684,N_10457,N_11182);
nor U12685 (N_12685,N_10890,N_10841);
xor U12686 (N_12686,N_11917,N_10592);
nor U12687 (N_12687,N_9435,N_9283);
nor U12688 (N_12688,N_9691,N_9700);
or U12689 (N_12689,N_11705,N_10939);
nand U12690 (N_12690,N_11387,N_10976);
nor U12691 (N_12691,N_10365,N_9193);
or U12692 (N_12692,N_9116,N_11580);
or U12693 (N_12693,N_9900,N_11680);
nor U12694 (N_12694,N_10008,N_10338);
nor U12695 (N_12695,N_9142,N_9230);
nor U12696 (N_12696,N_10705,N_11982);
xnor U12697 (N_12697,N_11278,N_10978);
nand U12698 (N_12698,N_11818,N_9948);
nor U12699 (N_12699,N_9858,N_10005);
nand U12700 (N_12700,N_11426,N_11693);
and U12701 (N_12701,N_10429,N_11403);
or U12702 (N_12702,N_9974,N_11266);
nand U12703 (N_12703,N_11932,N_9648);
and U12704 (N_12704,N_11009,N_9637);
and U12705 (N_12705,N_11804,N_10100);
nor U12706 (N_12706,N_9493,N_11743);
nor U12707 (N_12707,N_9973,N_10820);
and U12708 (N_12708,N_10076,N_9751);
nor U12709 (N_12709,N_9370,N_10600);
and U12710 (N_12710,N_11627,N_11825);
nand U12711 (N_12711,N_11653,N_9153);
nor U12712 (N_12712,N_11055,N_11023);
nand U12713 (N_12713,N_9318,N_10119);
and U12714 (N_12714,N_9957,N_11478);
nand U12715 (N_12715,N_10393,N_11450);
and U12716 (N_12716,N_10179,N_9488);
and U12717 (N_12717,N_11081,N_11543);
nand U12718 (N_12718,N_11868,N_11028);
nand U12719 (N_12719,N_11202,N_9541);
nand U12720 (N_12720,N_10829,N_10991);
nand U12721 (N_12721,N_11988,N_10786);
nand U12722 (N_12722,N_9044,N_11012);
and U12723 (N_12723,N_9888,N_10502);
or U12724 (N_12724,N_11184,N_9430);
or U12725 (N_12725,N_11465,N_10329);
nand U12726 (N_12726,N_11324,N_11221);
nor U12727 (N_12727,N_10935,N_11595);
nor U12728 (N_12728,N_9152,N_10052);
or U12729 (N_12729,N_9733,N_11146);
nand U12730 (N_12730,N_10089,N_10998);
nand U12731 (N_12731,N_11728,N_11393);
nor U12732 (N_12732,N_11003,N_10795);
and U12733 (N_12733,N_9074,N_9469);
and U12734 (N_12734,N_10401,N_10659);
and U12735 (N_12735,N_10887,N_9219);
or U12736 (N_12736,N_10444,N_9590);
and U12737 (N_12737,N_11666,N_11389);
or U12738 (N_12738,N_11717,N_11954);
nor U12739 (N_12739,N_11773,N_10162);
or U12740 (N_12740,N_9602,N_10278);
and U12741 (N_12741,N_11454,N_10769);
nand U12742 (N_12742,N_11704,N_10049);
or U12743 (N_12743,N_9437,N_11912);
nand U12744 (N_12744,N_10526,N_10793);
nor U12745 (N_12745,N_9445,N_10530);
nor U12746 (N_12746,N_9350,N_9698);
xnor U12747 (N_12747,N_9984,N_11651);
nand U12748 (N_12748,N_11104,N_11619);
or U12749 (N_12749,N_10981,N_10885);
nor U12750 (N_12750,N_9961,N_9007);
or U12751 (N_12751,N_11338,N_10722);
or U12752 (N_12752,N_9862,N_9520);
nand U12753 (N_12753,N_11352,N_11673);
nand U12754 (N_12754,N_9743,N_11566);
xnor U12755 (N_12755,N_11360,N_10116);
and U12756 (N_12756,N_11606,N_9433);
nor U12757 (N_12757,N_9421,N_11122);
or U12758 (N_12758,N_9721,N_10695);
or U12759 (N_12759,N_10581,N_10582);
nand U12760 (N_12760,N_10480,N_9385);
or U12761 (N_12761,N_9629,N_9279);
nor U12762 (N_12762,N_10003,N_10238);
or U12763 (N_12763,N_11113,N_11382);
nand U12764 (N_12764,N_10160,N_9908);
or U12765 (N_12765,N_11378,N_11224);
nor U12766 (N_12766,N_10570,N_9002);
and U12767 (N_12767,N_10423,N_10419);
nand U12768 (N_12768,N_11864,N_10293);
xnor U12769 (N_12769,N_11924,N_11546);
nand U12770 (N_12770,N_9067,N_11120);
nand U12771 (N_12771,N_9146,N_9966);
or U12772 (N_12772,N_11925,N_9202);
or U12773 (N_12773,N_9526,N_10783);
nor U12774 (N_12774,N_10539,N_10641);
nor U12775 (N_12775,N_9078,N_10114);
or U12776 (N_12776,N_9328,N_9473);
nand U12777 (N_12777,N_9099,N_9759);
or U12778 (N_12778,N_9552,N_11050);
nand U12779 (N_12779,N_9692,N_9132);
or U12780 (N_12780,N_9409,N_10392);
and U12781 (N_12781,N_9361,N_11492);
nor U12782 (N_12782,N_11794,N_9557);
nor U12783 (N_12783,N_11668,N_11263);
xor U12784 (N_12784,N_11160,N_10360);
xnor U12785 (N_12785,N_11716,N_9069);
nand U12786 (N_12786,N_11600,N_10267);
nand U12787 (N_12787,N_10825,N_11218);
nand U12788 (N_12788,N_10314,N_9757);
nor U12789 (N_12789,N_9023,N_9636);
or U12790 (N_12790,N_9465,N_11026);
nand U12791 (N_12791,N_10736,N_11215);
or U12792 (N_12792,N_9252,N_9910);
xnor U12793 (N_12793,N_9085,N_9529);
or U12794 (N_12794,N_10462,N_11745);
nor U12795 (N_12795,N_11438,N_9456);
or U12796 (N_12796,N_11458,N_9501);
nor U12797 (N_12797,N_11567,N_10744);
or U12798 (N_12798,N_10787,N_9426);
nor U12799 (N_12799,N_10780,N_10345);
or U12800 (N_12800,N_9710,N_10308);
and U12801 (N_12801,N_9565,N_9630);
nand U12802 (N_12802,N_10881,N_10737);
nand U12803 (N_12803,N_11255,N_11729);
xor U12804 (N_12804,N_10828,N_11507);
or U12805 (N_12805,N_11196,N_10728);
nor U12806 (N_12806,N_10095,N_10197);
and U12807 (N_12807,N_11170,N_9828);
or U12808 (N_12808,N_11501,N_10517);
nor U12809 (N_12809,N_10266,N_11134);
nor U12810 (N_12810,N_9243,N_9920);
or U12811 (N_12811,N_9676,N_9084);
and U12812 (N_12812,N_9261,N_9155);
or U12813 (N_12813,N_11014,N_9214);
nand U12814 (N_12814,N_9665,N_9049);
nand U12815 (N_12815,N_11045,N_11066);
and U12816 (N_12816,N_10601,N_10588);
and U12817 (N_12817,N_11576,N_9617);
nand U12818 (N_12818,N_11746,N_9525);
and U12819 (N_12819,N_10087,N_10512);
and U12820 (N_12820,N_11305,N_10426);
and U12821 (N_12821,N_11531,N_11880);
nor U12822 (N_12822,N_9555,N_10074);
and U12823 (N_12823,N_10244,N_11984);
or U12824 (N_12824,N_11613,N_11571);
or U12825 (N_12825,N_10934,N_11049);
nand U12826 (N_12826,N_9806,N_9286);
or U12827 (N_12827,N_9638,N_11304);
xnor U12828 (N_12828,N_11997,N_9718);
nor U12829 (N_12829,N_9073,N_9345);
nor U12830 (N_12830,N_11275,N_10213);
nand U12831 (N_12831,N_10463,N_10202);
nand U12832 (N_12832,N_10229,N_10689);
and U12833 (N_12833,N_9463,N_9242);
or U12834 (N_12834,N_10474,N_9233);
nor U12835 (N_12835,N_9601,N_10622);
or U12836 (N_12836,N_11635,N_11809);
nor U12837 (N_12837,N_11446,N_11220);
nor U12838 (N_12838,N_10090,N_9272);
and U12839 (N_12839,N_11713,N_11614);
or U12840 (N_12840,N_9054,N_11024);
or U12841 (N_12841,N_9255,N_10927);
and U12842 (N_12842,N_11523,N_10518);
or U12843 (N_12843,N_10915,N_9917);
nand U12844 (N_12844,N_9915,N_11719);
or U12845 (N_12845,N_9104,N_9967);
or U12846 (N_12846,N_10063,N_9874);
nand U12847 (N_12847,N_9374,N_10000);
nor U12848 (N_12848,N_11612,N_11910);
nand U12849 (N_12849,N_11374,N_11712);
nand U12850 (N_12850,N_9227,N_11351);
nor U12851 (N_12851,N_9912,N_9017);
nand U12852 (N_12852,N_11987,N_10872);
nor U12853 (N_12853,N_11075,N_9447);
nor U12854 (N_12854,N_11951,N_11771);
nand U12855 (N_12855,N_10388,N_10549);
nand U12856 (N_12856,N_10759,N_9780);
nand U12857 (N_12857,N_11829,N_9933);
or U12858 (N_12858,N_11569,N_9442);
or U12859 (N_12859,N_9197,N_10201);
or U12860 (N_12860,N_11131,N_10675);
or U12861 (N_12861,N_10261,N_9807);
or U12862 (N_12862,N_11812,N_11103);
or U12863 (N_12863,N_9690,N_10740);
nor U12864 (N_12864,N_10947,N_10702);
nand U12865 (N_12865,N_9166,N_10650);
nor U12866 (N_12866,N_10029,N_11115);
and U12867 (N_12867,N_11650,N_11700);
nor U12868 (N_12868,N_10483,N_9461);
and U12869 (N_12869,N_9545,N_9671);
or U12870 (N_12870,N_11585,N_9145);
and U12871 (N_12871,N_9560,N_10232);
or U12872 (N_12872,N_9489,N_11166);
nor U12873 (N_12873,N_11030,N_9719);
nand U12874 (N_12874,N_10758,N_10174);
or U12875 (N_12875,N_10900,N_10227);
and U12876 (N_12876,N_9628,N_9674);
nor U12877 (N_12877,N_11109,N_10033);
nor U12878 (N_12878,N_10816,N_9641);
xor U12879 (N_12879,N_11481,N_11395);
or U12880 (N_12880,N_9077,N_10273);
nor U12881 (N_12881,N_9878,N_11638);
nand U12882 (N_12882,N_11974,N_9837);
nand U12883 (N_12883,N_9408,N_9039);
or U12884 (N_12884,N_10070,N_11036);
nand U12885 (N_12885,N_11646,N_11963);
and U12886 (N_12886,N_11204,N_11797);
or U12887 (N_12887,N_9200,N_10224);
nor U12888 (N_12888,N_10207,N_11978);
nand U12889 (N_12889,N_10537,N_9983);
or U12890 (N_12890,N_10553,N_9165);
nand U12891 (N_12891,N_9216,N_9090);
nand U12892 (N_12892,N_11579,N_10430);
nor U12893 (N_12893,N_9911,N_11758);
nor U12894 (N_12894,N_9926,N_11587);
or U12895 (N_12895,N_11405,N_11483);
or U12896 (N_12896,N_11444,N_11341);
and U12897 (N_12897,N_9213,N_10948);
nor U12898 (N_12898,N_11502,N_11547);
or U12899 (N_12899,N_11748,N_9302);
nand U12900 (N_12900,N_10551,N_9455);
nand U12901 (N_12901,N_10021,N_11128);
xnor U12902 (N_12902,N_9112,N_11329);
nor U12903 (N_12903,N_11769,N_10286);
nor U12904 (N_12904,N_9237,N_10864);
and U12905 (N_12905,N_9410,N_9334);
and U12906 (N_12906,N_11112,N_9388);
nand U12907 (N_12907,N_9534,N_10727);
or U12908 (N_12908,N_10751,N_10481);
nand U12909 (N_12909,N_10467,N_10839);
nand U12910 (N_12910,N_9773,N_11678);
nor U12911 (N_12911,N_9860,N_10955);
nand U12912 (N_12912,N_9604,N_10933);
and U12913 (N_12913,N_11744,N_11260);
nand U12914 (N_12914,N_9679,N_10607);
and U12915 (N_12915,N_9336,N_10874);
and U12916 (N_12916,N_10334,N_11768);
xor U12917 (N_12917,N_11111,N_9689);
and U12918 (N_12918,N_10827,N_10673);
and U12919 (N_12919,N_10017,N_9748);
or U12920 (N_12920,N_11933,N_9436);
and U12921 (N_12921,N_9396,N_10134);
nand U12922 (N_12922,N_9955,N_11363);
and U12923 (N_12923,N_11654,N_10664);
or U12924 (N_12924,N_9796,N_10490);
and U12925 (N_12925,N_9288,N_9708);
nor U12926 (N_12926,N_10140,N_10713);
nor U12927 (N_12927,N_11993,N_10554);
nand U12928 (N_12928,N_10901,N_10385);
and U12929 (N_12929,N_11893,N_11384);
nand U12930 (N_12930,N_10858,N_11249);
nand U12931 (N_12931,N_11878,N_10235);
or U12932 (N_12932,N_11896,N_11333);
or U12933 (N_12933,N_11430,N_9238);
nor U12934 (N_12934,N_9217,N_11076);
or U12935 (N_12935,N_9939,N_9038);
and U12936 (N_12936,N_10313,N_11377);
xnor U12937 (N_12937,N_11798,N_11676);
and U12938 (N_12938,N_9281,N_10446);
or U12939 (N_12939,N_9797,N_10850);
xnor U12940 (N_12940,N_11861,N_10637);
or U12941 (N_12941,N_11043,N_10499);
or U12942 (N_12942,N_10614,N_10190);
nand U12943 (N_12943,N_11449,N_9999);
nor U12944 (N_12944,N_9639,N_9581);
nand U12945 (N_12945,N_9598,N_9490);
and U12946 (N_12946,N_11575,N_11392);
nor U12947 (N_12947,N_9795,N_9404);
and U12948 (N_12948,N_9977,N_9633);
nor U12949 (N_12949,N_11958,N_11976);
nand U12950 (N_12950,N_11604,N_10118);
or U12951 (N_12951,N_9658,N_9470);
nand U12952 (N_12952,N_11827,N_9502);
and U12953 (N_12953,N_11882,N_11287);
nand U12954 (N_12954,N_11692,N_10097);
nand U12955 (N_12955,N_11340,N_10975);
nor U12956 (N_12956,N_10604,N_9697);
or U12957 (N_12957,N_10056,N_9760);
nand U12958 (N_12958,N_10666,N_11684);
nor U12959 (N_12959,N_9626,N_10815);
nand U12960 (N_12960,N_11957,N_10757);
or U12961 (N_12961,N_10111,N_10303);
nor U12962 (N_12962,N_10437,N_11037);
nor U12963 (N_12963,N_9131,N_11824);
and U12964 (N_12964,N_11657,N_10836);
nand U12965 (N_12965,N_9766,N_10245);
and U12966 (N_12966,N_10967,N_9512);
nand U12967 (N_12967,N_9425,N_9186);
nor U12968 (N_12968,N_9724,N_11488);
and U12969 (N_12969,N_10805,N_9225);
nor U12970 (N_12970,N_11686,N_10326);
and U12971 (N_12971,N_9696,N_9817);
or U12972 (N_12972,N_11145,N_11894);
and U12973 (N_12973,N_10677,N_9504);
or U12974 (N_12974,N_11306,N_10721);
nand U12975 (N_12975,N_10845,N_9610);
and U12976 (N_12976,N_11346,N_11257);
or U12977 (N_12977,N_9331,N_11476);
and U12978 (N_12978,N_9935,N_11069);
and U12979 (N_12979,N_10079,N_11766);
nand U12980 (N_12980,N_10448,N_11941);
nand U12981 (N_12981,N_11172,N_11649);
nand U12982 (N_12982,N_11577,N_11225);
and U12983 (N_12983,N_9758,N_9855);
nand U12984 (N_12984,N_9140,N_10676);
nor U12985 (N_12985,N_10913,N_11290);
or U12986 (N_12986,N_11598,N_11630);
nand U12987 (N_12987,N_9240,N_11190);
and U12988 (N_12988,N_11420,N_9680);
and U12989 (N_12989,N_11940,N_11741);
or U12990 (N_12990,N_9081,N_11930);
nor U12991 (N_12991,N_10651,N_9179);
xnor U12992 (N_12992,N_10167,N_10497);
nand U12993 (N_12993,N_10799,N_9451);
and U12994 (N_12994,N_9025,N_10973);
nor U12995 (N_12995,N_10834,N_11913);
or U12996 (N_12996,N_11060,N_10724);
or U12997 (N_12997,N_11423,N_10287);
nand U12998 (N_12998,N_11070,N_10734);
nor U12999 (N_12999,N_9277,N_10233);
or U13000 (N_13000,N_10970,N_9865);
nand U13001 (N_13001,N_11947,N_11119);
nand U13002 (N_13002,N_9485,N_11261);
or U13003 (N_13003,N_11327,N_9782);
nor U13004 (N_13004,N_11253,N_11189);
or U13005 (N_13005,N_9424,N_11555);
xnor U13006 (N_13006,N_9769,N_11452);
or U13007 (N_13007,N_10081,N_11980);
nand U13008 (N_13008,N_11041,N_11125);
nor U13009 (N_13009,N_10715,N_11181);
or U13010 (N_13010,N_10400,N_10719);
and U13011 (N_13011,N_11212,N_11156);
nand U13012 (N_13012,N_9459,N_9812);
and U13013 (N_13013,N_11631,N_11227);
nand U13014 (N_13014,N_10961,N_9923);
and U13015 (N_13015,N_10136,N_10806);
nor U13016 (N_13016,N_10312,N_9138);
nand U13017 (N_13017,N_9761,N_11703);
and U13018 (N_13018,N_9884,N_9930);
and U13019 (N_13019,N_9264,N_11909);
nand U13020 (N_13020,N_10842,N_10249);
nor U13021 (N_13021,N_9785,N_10682);
or U13022 (N_13022,N_9882,N_9978);
nand U13023 (N_13023,N_9872,N_10595);
or U13024 (N_13024,N_9448,N_9843);
or U13025 (N_13025,N_10011,N_9918);
or U13026 (N_13026,N_9826,N_10153);
nor U13027 (N_13027,N_9319,N_10577);
nor U13028 (N_13028,N_11130,N_11079);
and U13029 (N_13029,N_9540,N_9944);
and U13030 (N_13030,N_10849,N_11644);
and U13031 (N_13031,N_9899,N_9199);
or U13032 (N_13032,N_10306,N_9118);
nor U13033 (N_13033,N_10525,N_11365);
nand U13034 (N_13034,N_11992,N_11301);
or U13035 (N_13035,N_10876,N_11443);
nor U13036 (N_13036,N_9312,N_10085);
nor U13037 (N_13037,N_11303,N_10185);
or U13038 (N_13038,N_11436,N_10018);
and U13039 (N_13039,N_9850,N_11006);
nor U13040 (N_13040,N_10513,N_11044);
or U13041 (N_13041,N_10319,N_10316);
nor U13042 (N_13042,N_10433,N_11849);
and U13043 (N_13043,N_9354,N_10700);
nor U13044 (N_13044,N_10558,N_11564);
nand U13045 (N_13045,N_11755,N_11872);
or U13046 (N_13046,N_10062,N_11906);
and U13047 (N_13047,N_11991,N_9969);
or U13048 (N_13048,N_9783,N_11474);
and U13049 (N_13049,N_9338,N_10391);
nor U13050 (N_13050,N_11890,N_9258);
or U13051 (N_13051,N_9231,N_9732);
and U13052 (N_13052,N_9457,N_9798);
or U13053 (N_13053,N_11039,N_9207);
xnor U13054 (N_13054,N_11573,N_9008);
xnor U13055 (N_13055,N_9968,N_10256);
or U13056 (N_13056,N_10988,N_11323);
nor U13057 (N_13057,N_10048,N_10584);
nor U13058 (N_13058,N_11230,N_9379);
nor U13059 (N_13059,N_9249,N_10367);
nor U13060 (N_13060,N_9954,N_11534);
or U13061 (N_13061,N_11636,N_11696);
or U13062 (N_13062,N_11553,N_11873);
and U13063 (N_13063,N_10470,N_11239);
and U13064 (N_13064,N_9778,N_11539);
or U13065 (N_13065,N_11702,N_10528);
and U13066 (N_13066,N_9825,N_10127);
or U13067 (N_13067,N_11375,N_9889);
or U13068 (N_13068,N_10006,N_9594);
or U13069 (N_13069,N_11163,N_10654);
nor U13070 (N_13070,N_10672,N_11515);
nand U13071 (N_13071,N_9321,N_11150);
nor U13072 (N_13072,N_10718,N_11967);
nor U13073 (N_13073,N_11077,N_11029);
nor U13074 (N_13074,N_11986,N_10060);
or U13075 (N_13075,N_10784,N_11608);
and U13076 (N_13076,N_9088,N_11001);
or U13077 (N_13077,N_11254,N_10617);
nand U13078 (N_13078,N_9428,N_10962);
nor U13079 (N_13079,N_9879,N_9542);
nor U13080 (N_13080,N_10456,N_10250);
or U13081 (N_13081,N_10789,N_11002);
or U13082 (N_13082,N_11632,N_10193);
nor U13083 (N_13083,N_10237,N_9254);
or U13084 (N_13084,N_9154,N_11578);
and U13085 (N_13085,N_10779,N_10855);
and U13086 (N_13086,N_11817,N_10920);
and U13087 (N_13087,N_9042,N_10298);
or U13088 (N_13088,N_11889,N_11641);
or U13089 (N_13089,N_9296,N_9109);
or U13090 (N_13090,N_10394,N_9108);
xnor U13091 (N_13091,N_11597,N_11779);
and U13092 (N_13092,N_11859,N_11761);
or U13093 (N_13093,N_10561,N_11416);
nand U13094 (N_13094,N_9819,N_10794);
and U13095 (N_13095,N_9829,N_9159);
and U13096 (N_13096,N_9173,N_10045);
or U13097 (N_13097,N_9675,N_11591);
nand U13098 (N_13098,N_11082,N_11556);
nand U13099 (N_13099,N_9989,N_10945);
nand U13100 (N_13100,N_10956,N_11067);
and U13101 (N_13101,N_9212,N_11482);
nand U13102 (N_13102,N_10460,N_10723);
or U13103 (N_13103,N_10046,N_10569);
nor U13104 (N_13104,N_10980,N_10344);
xor U13105 (N_13105,N_10716,N_11593);
xnor U13106 (N_13106,N_11985,N_11210);
nor U13107 (N_13107,N_9399,N_9627);
nand U13108 (N_13108,N_11949,N_11618);
and U13109 (N_13109,N_10776,N_11911);
nand U13110 (N_13110,N_11923,N_9736);
nor U13111 (N_13111,N_11295,N_11732);
and U13112 (N_13112,N_10897,N_9156);
nor U13113 (N_13113,N_9136,N_10347);
nor U13114 (N_13114,N_11434,N_9076);
xnor U13115 (N_13115,N_10492,N_9484);
or U13116 (N_13116,N_11747,N_9992);
or U13117 (N_13117,N_10108,N_10445);
nand U13118 (N_13118,N_9343,N_9373);
or U13119 (N_13119,N_9731,N_10589);
nor U13120 (N_13120,N_9949,N_11466);
xnor U13121 (N_13121,N_10348,N_11457);
nand U13122 (N_13122,N_9508,N_11962);
and U13123 (N_13123,N_10498,N_9624);
and U13124 (N_13124,N_10752,N_11774);
nor U13125 (N_13125,N_10946,N_10636);
and U13126 (N_13126,N_9188,N_10692);
nand U13127 (N_13127,N_10767,N_11948);
and U13128 (N_13128,N_9522,N_9739);
nor U13129 (N_13129,N_9270,N_11540);
nand U13130 (N_13130,N_9929,N_10019);
nor U13131 (N_13131,N_11720,N_9378);
or U13132 (N_13132,N_11008,N_9497);
and U13133 (N_13133,N_10873,N_10346);
or U13134 (N_13134,N_10653,N_9293);
nand U13135 (N_13135,N_11541,N_9358);
or U13136 (N_13136,N_10792,N_10195);
or U13137 (N_13137,N_9251,N_9921);
and U13138 (N_13138,N_10024,N_10323);
nand U13139 (N_13139,N_11964,N_10931);
or U13140 (N_13140,N_11551,N_11274);
nor U13141 (N_13141,N_11599,N_11315);
and U13142 (N_13142,N_11371,N_11013);
and U13143 (N_13143,N_11088,N_10543);
or U13144 (N_13144,N_10148,N_10176);
and U13145 (N_13145,N_11782,N_10110);
and U13146 (N_13146,N_10459,N_10871);
and U13147 (N_13147,N_10782,N_11981);
xnor U13148 (N_13148,N_9897,N_9851);
nor U13149 (N_13149,N_9033,N_10944);
nor U13150 (N_13150,N_9943,N_10765);
or U13151 (N_13151,N_11525,N_9536);
nor U13152 (N_13152,N_10113,N_11786);
or U13153 (N_13153,N_10615,N_11485);
or U13154 (N_13154,N_11222,N_10362);
and U13155 (N_13155,N_9006,N_9822);
and U13156 (N_13156,N_10341,N_9072);
or U13157 (N_13157,N_11369,N_10696);
nor U13158 (N_13158,N_11226,N_11318);
nand U13159 (N_13159,N_9427,N_11999);
or U13160 (N_13160,N_9429,N_11869);
xnor U13161 (N_13161,N_11307,N_9985);
or U13162 (N_13162,N_10555,N_9177);
nand U13163 (N_13163,N_10506,N_10790);
or U13164 (N_13164,N_9621,N_10473);
nor U13165 (N_13165,N_11032,N_10196);
and U13166 (N_13166,N_11244,N_11862);
or U13167 (N_13167,N_11061,N_9924);
or U13168 (N_13168,N_10848,N_9107);
and U13169 (N_13169,N_11057,N_9464);
or U13170 (N_13170,N_11381,N_9745);
nor U13171 (N_13171,N_10302,N_9582);
nand U13172 (N_13172,N_9297,N_11998);
nor U13173 (N_13173,N_9734,N_9250);
and U13174 (N_13174,N_9001,N_10487);
or U13175 (N_13175,N_11137,N_11611);
and U13176 (N_13176,N_9663,N_11183);
nand U13177 (N_13177,N_9867,N_11296);
or U13178 (N_13178,N_10281,N_9705);
nand U13179 (N_13179,N_9303,N_11751);
or U13180 (N_13180,N_11106,N_9827);
and U13181 (N_13181,N_10889,N_11610);
nor U13182 (N_13182,N_9415,N_9128);
nand U13183 (N_13183,N_9533,N_10606);
or U13184 (N_13184,N_11090,N_10354);
and U13185 (N_13185,N_9763,N_11672);
nor U13186 (N_13186,N_9482,N_10358);
and U13187 (N_13187,N_10320,N_10986);
nand U13188 (N_13188,N_10386,N_10822);
and U13189 (N_13189,N_10465,N_10922);
or U13190 (N_13190,N_11559,N_9106);
nand U13191 (N_13191,N_10378,N_9086);
or U13192 (N_13192,N_11238,N_10037);
and U13193 (N_13193,N_10073,N_9543);
and U13194 (N_13194,N_9661,N_10778);
nor U13195 (N_13195,N_11811,N_10276);
nand U13196 (N_13196,N_10241,N_9419);
and U13197 (N_13197,N_11176,N_11236);
and U13198 (N_13198,N_9659,N_11645);
and U13199 (N_13199,N_10534,N_10950);
and U13200 (N_13200,N_11177,N_9417);
nand U13201 (N_13201,N_10522,N_9737);
and U13202 (N_13202,N_11409,N_11596);
nor U13203 (N_13203,N_9950,N_9713);
and U13204 (N_13204,N_10151,N_9119);
or U13205 (N_13205,N_11159,N_10169);
or U13206 (N_13206,N_11308,N_10425);
nor U13207 (N_13207,N_9082,N_11391);
and U13208 (N_13208,N_9317,N_10938);
or U13209 (N_13209,N_9089,N_10203);
nor U13210 (N_13210,N_9789,N_11425);
xor U13211 (N_13211,N_10738,N_11944);
nor U13212 (N_13212,N_10091,N_10691);
and U13213 (N_13213,N_10863,N_10412);
nor U13214 (N_13214,N_11453,N_9332);
nor U13215 (N_13215,N_10451,N_9151);
and U13216 (N_13216,N_11820,N_9962);
nand U13217 (N_13217,N_10536,N_11078);
nand U13218 (N_13218,N_11479,N_11854);
or U13219 (N_13219,N_11251,N_10563);
and U13220 (N_13220,N_10670,N_11537);
nand U13221 (N_13221,N_9741,N_9863);
and U13222 (N_13222,N_9688,N_11956);
or U13223 (N_13223,N_10503,N_9161);
nor U13224 (N_13224,N_11228,N_11256);
nor U13225 (N_13225,N_10032,N_10693);
nor U13226 (N_13226,N_11095,N_11386);
or U13227 (N_13227,N_9275,N_11005);
or U13228 (N_13228,N_11831,N_9712);
nor U13229 (N_13229,N_10263,N_9527);
nand U13230 (N_13230,N_10455,N_9246);
nand U13231 (N_13231,N_11339,N_9364);
nand U13232 (N_13232,N_9440,N_11877);
or U13233 (N_13233,N_10047,N_9804);
and U13234 (N_13234,N_10205,N_9901);
and U13235 (N_13235,N_9325,N_11953);
or U13236 (N_13236,N_11724,N_9830);
nand U13237 (N_13237,N_9034,N_11663);
nand U13238 (N_13238,N_11229,N_9642);
nand U13239 (N_13239,N_10586,N_9247);
xnor U13240 (N_13240,N_11155,N_9864);
nor U13241 (N_13241,N_11178,N_10051);
nand U13242 (N_13242,N_11681,N_10317);
or U13243 (N_13243,N_11971,N_9059);
and U13244 (N_13244,N_9753,N_9368);
nand U13245 (N_13245,N_10297,N_9685);
and U13246 (N_13246,N_9480,N_11522);
and U13247 (N_13247,N_9203,N_10710);
or U13248 (N_13248,N_10992,N_10987);
nand U13249 (N_13249,N_9787,N_10808);
and U13250 (N_13250,N_10275,N_11918);
nor U13251 (N_13251,N_9513,N_11765);
or U13252 (N_13252,N_10643,N_10357);
and U13253 (N_13253,N_11996,N_9040);
nor U13254 (N_13254,N_11380,N_9114);
nor U13255 (N_13255,N_11807,N_9229);
nor U13256 (N_13256,N_11404,N_9720);
nand U13257 (N_13257,N_11781,N_9204);
nand U13258 (N_13258,N_11289,N_10002);
nand U13259 (N_13259,N_10230,N_11258);
or U13260 (N_13260,N_11772,N_11194);
and U13261 (N_13261,N_11322,N_9538);
or U13262 (N_13262,N_10802,N_10814);
and U13263 (N_13263,N_10246,N_9591);
nor U13264 (N_13264,N_11875,N_11089);
nor U13265 (N_13265,N_11433,N_9026);
nand U13266 (N_13266,N_9972,N_9313);
xor U13267 (N_13267,N_11071,N_11821);
nand U13268 (N_13268,N_10590,N_9622);
nand U13269 (N_13269,N_9956,N_11418);
or U13270 (N_13270,N_11291,N_9666);
and U13271 (N_13271,N_9856,N_11625);
nand U13272 (N_13272,N_9333,N_10609);
nor U13273 (N_13273,N_11826,N_11642);
nor U13274 (N_13274,N_9121,N_11520);
nand U13275 (N_13275,N_11493,N_11528);
nor U13276 (N_13276,N_9794,N_11938);
and U13277 (N_13277,N_9434,N_9127);
nand U13278 (N_13278,N_10851,N_9322);
and U13279 (N_13279,N_10963,N_11500);
nor U13280 (N_13280,N_11574,N_11264);
nor U13281 (N_13281,N_9468,N_9824);
or U13282 (N_13282,N_11390,N_11118);
nand U13283 (N_13283,N_11884,N_11529);
nor U13284 (N_13284,N_10566,N_9640);
nand U13285 (N_13285,N_11456,N_9158);
or U13286 (N_13286,N_10748,N_11406);
nor U13287 (N_13287,N_10104,N_11344);
nand U13288 (N_13288,N_10801,N_10844);
nand U13289 (N_13289,N_9903,N_10545);
nand U13290 (N_13290,N_10395,N_10133);
and U13291 (N_13291,N_9190,N_9295);
nor U13292 (N_13292,N_11521,N_11835);
or U13293 (N_13293,N_9519,N_10709);
or U13294 (N_13294,N_10532,N_10187);
or U13295 (N_13295,N_11628,N_11139);
nor U13296 (N_13296,N_9450,N_10511);
and U13297 (N_13297,N_11674,N_9619);
nand U13298 (N_13298,N_10271,N_11414);
nand U13299 (N_13299,N_11020,N_10730);
and U13300 (N_13300,N_9958,N_9895);
nand U13301 (N_13301,N_9960,N_10411);
or U13302 (N_13302,N_10209,N_11659);
or U13303 (N_13303,N_11370,N_10635);
nand U13304 (N_13304,N_11943,N_9228);
nor U13305 (N_13305,N_9164,N_9945);
nand U13306 (N_13306,N_10529,N_9035);
xnor U13307 (N_13307,N_11842,N_10064);
nand U13308 (N_13308,N_11589,N_11442);
or U13309 (N_13309,N_11775,N_9309);
nand U13310 (N_13310,N_10088,N_10867);
nor U13311 (N_13311,N_11342,N_10166);
nor U13312 (N_13312,N_11361,N_10422);
or U13313 (N_13313,N_10038,N_9891);
nand U13314 (N_13314,N_11429,N_9653);
xnor U13315 (N_13315,N_9996,N_10406);
nor U13316 (N_13316,N_10075,N_11620);
nand U13317 (N_13317,N_10030,N_9881);
and U13318 (N_13318,N_10587,N_9844);
nor U13319 (N_13319,N_11265,N_9799);
nor U13320 (N_13320,N_10403,N_11063);
nand U13321 (N_13321,N_11685,N_9386);
and U13322 (N_13322,N_9032,N_9187);
xor U13323 (N_13323,N_9181,N_11694);
or U13324 (N_13324,N_11789,N_10315);
or U13325 (N_13325,N_10741,N_10080);
nand U13326 (N_13326,N_9245,N_11815);
or U13327 (N_13327,N_9329,N_11509);
nand U13328 (N_13328,N_9323,N_9599);
and U13329 (N_13329,N_9327,N_11660);
nand U13330 (N_13330,N_10192,N_9394);
nor U13331 (N_13331,N_10669,N_9805);
or U13332 (N_13332,N_11706,N_10436);
or U13333 (N_13333,N_9925,N_10735);
nand U13334 (N_13334,N_9681,N_9730);
or U13335 (N_13335,N_10797,N_11283);
nor U13336 (N_13336,N_9562,N_9300);
nor U13337 (N_13337,N_10311,N_11844);
and U13338 (N_13338,N_10917,N_9353);
nor U13339 (N_13339,N_9441,N_10199);
or U13340 (N_13340,N_11883,N_10846);
nand U13341 (N_13341,N_10557,N_11544);
nor U13342 (N_13342,N_10449,N_10542);
nor U13343 (N_13343,N_11851,N_10039);
nor U13344 (N_13344,N_9274,N_9091);
or U13345 (N_13345,N_10325,N_9905);
nor U13346 (N_13346,N_9947,N_10291);
nand U13347 (N_13347,N_9580,N_10328);
nor U13348 (N_13348,N_9711,N_10399);
nand U13349 (N_13349,N_11526,N_10290);
or U13350 (N_13350,N_10843,N_9873);
nand U13351 (N_13351,N_10138,N_11209);
or U13352 (N_13352,N_10135,N_10120);
nor U13353 (N_13353,N_10688,N_11634);
nor U13354 (N_13354,N_11025,N_11494);
nand U13355 (N_13355,N_9314,N_11617);
nand U13356 (N_13356,N_11871,N_11054);
nand U13357 (N_13357,N_9673,N_11435);
nand U13358 (N_13358,N_10381,N_9728);
nor U13359 (N_13359,N_9365,N_11180);
and U13360 (N_13360,N_10853,N_11068);
nor U13361 (N_13361,N_10122,N_9942);
and U13362 (N_13362,N_9647,N_10698);
nor U13363 (N_13363,N_9196,N_11268);
nand U13364 (N_13364,N_10720,N_9662);
nor U13365 (N_13365,N_9013,N_9667);
nor U13366 (N_13366,N_10109,N_10552);
nand U13367 (N_13367,N_9716,N_10098);
nor U13368 (N_13368,N_9814,N_10574);
nand U13369 (N_13369,N_9507,N_11926);
or U13370 (N_13370,N_10711,N_11968);
or U13371 (N_13371,N_10547,N_10628);
and U13372 (N_13372,N_10559,N_9198);
and U13373 (N_13373,N_10661,N_11411);
nor U13374 (N_13374,N_11590,N_11292);
or U13375 (N_13375,N_11349,N_9558);
and U13376 (N_13376,N_9390,N_11472);
nand U13377 (N_13377,N_9657,N_11690);
nand U13378 (N_13378,N_10318,N_11234);
and U13379 (N_13379,N_11757,N_10914);
nor U13380 (N_13380,N_9305,N_11053);
nor U13381 (N_13381,N_9747,N_10966);
nor U13382 (N_13382,N_9020,N_11907);
and U13383 (N_13383,N_10879,N_10484);
or U13384 (N_13384,N_11147,N_11532);
nor U13385 (N_13385,N_10222,N_9369);
and U13386 (N_13386,N_10562,N_11519);
xnor U13387 (N_13387,N_11535,N_11723);
or U13388 (N_13388,N_9616,N_11373);
nor U13389 (N_13389,N_9380,N_10226);
nand U13390 (N_13390,N_9511,N_10678);
nand U13391 (N_13391,N_9079,N_10701);
xor U13392 (N_13392,N_11294,N_9304);
nand U13393 (N_13393,N_11007,N_10183);
or U13394 (N_13394,N_9494,N_10355);
nor U13395 (N_13395,N_9551,N_9348);
nor U13396 (N_13396,N_10194,N_9531);
nand U13397 (N_13397,N_11136,N_11701);
nand U13398 (N_13398,N_9356,N_9600);
and U13399 (N_13399,N_10957,N_9422);
or U13400 (N_13400,N_11332,N_11248);
nand U13401 (N_13401,N_10450,N_10575);
and U13402 (N_13402,N_11286,N_10152);
nor U13403 (N_13403,N_9105,N_10219);
nand U13404 (N_13404,N_10612,N_10154);
or U13405 (N_13405,N_10031,N_11816);
and U13406 (N_13406,N_11832,N_10438);
nor U13407 (N_13407,N_9815,N_9257);
and U13408 (N_13408,N_11407,N_9359);
and U13409 (N_13409,N_9623,N_10932);
nor U13410 (N_13410,N_11903,N_11548);
nand U13411 (N_13411,N_11823,N_10729);
nand U13412 (N_13412,N_10404,N_10540);
or U13413 (N_13413,N_11321,N_10611);
or U13414 (N_13414,N_11358,N_11470);
or U13415 (N_13415,N_11126,N_9472);
xnor U13416 (N_13416,N_9201,N_9094);
nor U13417 (N_13417,N_10439,N_10977);
nand U13418 (N_13418,N_11853,N_9027);
or U13419 (N_13419,N_9005,N_9772);
and U13420 (N_13420,N_9546,N_9092);
and U13421 (N_13421,N_10707,N_10184);
nand U13422 (N_13422,N_11655,N_10277);
nor U13423 (N_13423,N_11093,N_10416);
nand U13424 (N_13424,N_9523,N_10990);
and U13425 (N_13425,N_9232,N_11484);
and U13426 (N_13426,N_9416,N_9876);
nor U13427 (N_13427,N_11279,N_10383);
xnor U13428 (N_13428,N_9635,N_9065);
and U13429 (N_13429,N_9057,N_10461);
nor U13430 (N_13430,N_11259,N_10257);
nor U13431 (N_13431,N_10788,N_9655);
or U13432 (N_13432,N_9997,N_10204);
and U13433 (N_13433,N_9853,N_10854);
nor U13434 (N_13434,N_11536,N_11293);
nand U13435 (N_13435,N_11742,N_9717);
or U13436 (N_13436,N_9740,N_10107);
nand U13437 (N_13437,N_10706,N_9553);
nand U13438 (N_13438,N_10940,N_10859);
and U13439 (N_13439,N_10146,N_9808);
or U13440 (N_13440,N_10242,N_11165);
and U13441 (N_13441,N_10907,N_9045);
nor U13442 (N_13442,N_9362,N_11586);
or U13443 (N_13443,N_9175,N_10658);
or U13444 (N_13444,N_10434,N_10985);
nor U13445 (N_13445,N_10132,N_10043);
or U13446 (N_13446,N_11459,N_11233);
or U13447 (N_13447,N_9840,N_11935);
or U13448 (N_13448,N_9285,N_10364);
nand U13449 (N_13449,N_9414,N_9896);
nand U13450 (N_13450,N_11019,N_10228);
and U13451 (N_13451,N_11105,N_10402);
and U13452 (N_13452,N_11018,N_9838);
or U13453 (N_13453,N_11489,N_9058);
and U13454 (N_13454,N_11245,N_11031);
nand U13455 (N_13455,N_10813,N_11401);
nor U13456 (N_13456,N_9019,N_10773);
or U13457 (N_13457,N_9126,N_10280);
and U13458 (N_13458,N_9310,N_11282);
or U13459 (N_13459,N_10868,N_9139);
and U13460 (N_13460,N_11397,N_9991);
nand U13461 (N_13461,N_9746,N_11185);
nor U13462 (N_13462,N_11752,N_11791);
nand U13463 (N_13463,N_10025,N_9530);
or U13464 (N_13464,N_9650,N_10684);
nor U13465 (N_13465,N_11677,N_9987);
nor U13466 (N_13466,N_9360,N_10785);
or U13467 (N_13467,N_10150,N_11945);
or U13468 (N_13468,N_11790,N_10413);
or U13469 (N_13469,N_11473,N_11995);
nand U13470 (N_13470,N_11462,N_9768);
nand U13471 (N_13471,N_9000,N_11788);
and U13472 (N_13472,N_11151,N_10464);
and U13473 (N_13473,N_11320,N_10044);
or U13474 (N_13474,N_10667,N_9191);
nand U13475 (N_13475,N_9342,N_10657);
and U13476 (N_13476,N_10067,N_10571);
nor U13477 (N_13477,N_11298,N_11499);
nand U13478 (N_13478,N_11169,N_10145);
and U13479 (N_13479,N_10282,N_11191);
or U13480 (N_13480,N_11348,N_10093);
or U13481 (N_13481,N_9299,N_10810);
and U13482 (N_13482,N_9096,N_11042);
nor U13483 (N_13483,N_9235,N_10599);
nand U13484 (N_13484,N_10959,N_10254);
and U13485 (N_13485,N_10225,N_10259);
xnor U13486 (N_13486,N_10770,N_9467);
or U13487 (N_13487,N_11288,N_9770);
and U13488 (N_13488,N_9547,N_10629);
nand U13489 (N_13489,N_10505,N_10299);
nand U13490 (N_13490,N_10001,N_9618);
nor U13491 (N_13491,N_9087,N_11785);
and U13492 (N_13492,N_10265,N_10288);
nand U13493 (N_13493,N_11583,N_11866);
nor U13494 (N_13494,N_10084,N_11727);
and U13495 (N_13495,N_10377,N_11051);
or U13496 (N_13496,N_11247,N_11762);
and U13497 (N_13497,N_11664,N_11814);
nor U13498 (N_13498,N_10408,N_11518);
or U13499 (N_13499,N_11415,N_11633);
nor U13500 (N_13500,N_10256,N_9305);
nand U13501 (N_13501,N_9661,N_10325);
nor U13502 (N_13502,N_10557,N_9120);
xor U13503 (N_13503,N_11474,N_9699);
nand U13504 (N_13504,N_10346,N_10272);
nand U13505 (N_13505,N_11161,N_9116);
nand U13506 (N_13506,N_10114,N_9887);
and U13507 (N_13507,N_11234,N_10595);
nand U13508 (N_13508,N_9070,N_11103);
nor U13509 (N_13509,N_10503,N_11004);
nand U13510 (N_13510,N_10415,N_11160);
and U13511 (N_13511,N_11234,N_9643);
nand U13512 (N_13512,N_10316,N_11116);
and U13513 (N_13513,N_10289,N_11502);
nor U13514 (N_13514,N_11885,N_10527);
and U13515 (N_13515,N_10387,N_11491);
nand U13516 (N_13516,N_9402,N_11871);
and U13517 (N_13517,N_9612,N_11140);
or U13518 (N_13518,N_11127,N_9319);
and U13519 (N_13519,N_11984,N_10258);
and U13520 (N_13520,N_10112,N_10323);
nand U13521 (N_13521,N_9888,N_9048);
and U13522 (N_13522,N_9715,N_10901);
and U13523 (N_13523,N_9110,N_10247);
nand U13524 (N_13524,N_10547,N_11783);
and U13525 (N_13525,N_10988,N_11041);
nor U13526 (N_13526,N_11759,N_10290);
and U13527 (N_13527,N_11926,N_9487);
nand U13528 (N_13528,N_10967,N_11787);
or U13529 (N_13529,N_10920,N_11352);
and U13530 (N_13530,N_9870,N_11916);
and U13531 (N_13531,N_11255,N_9919);
and U13532 (N_13532,N_11803,N_11630);
and U13533 (N_13533,N_11880,N_9872);
and U13534 (N_13534,N_9312,N_9536);
nand U13535 (N_13535,N_9403,N_11185);
and U13536 (N_13536,N_10228,N_11758);
nand U13537 (N_13537,N_10491,N_9155);
or U13538 (N_13538,N_11339,N_10834);
and U13539 (N_13539,N_11533,N_9987);
and U13540 (N_13540,N_9828,N_9760);
or U13541 (N_13541,N_11952,N_10722);
nand U13542 (N_13542,N_10387,N_9338);
and U13543 (N_13543,N_10217,N_11527);
xor U13544 (N_13544,N_10260,N_11285);
or U13545 (N_13545,N_9607,N_11958);
or U13546 (N_13546,N_10270,N_11034);
and U13547 (N_13547,N_10678,N_11497);
or U13548 (N_13548,N_9326,N_9798);
nor U13549 (N_13549,N_11617,N_10097);
or U13550 (N_13550,N_11823,N_10221);
or U13551 (N_13551,N_9436,N_11520);
or U13552 (N_13552,N_9726,N_11447);
or U13553 (N_13553,N_11577,N_11241);
and U13554 (N_13554,N_11865,N_9365);
or U13555 (N_13555,N_10717,N_9051);
nand U13556 (N_13556,N_11030,N_9340);
nor U13557 (N_13557,N_10114,N_11630);
nor U13558 (N_13558,N_11382,N_9115);
or U13559 (N_13559,N_10069,N_9106);
nand U13560 (N_13560,N_11066,N_9757);
and U13561 (N_13561,N_10001,N_9901);
nand U13562 (N_13562,N_10658,N_9134);
nand U13563 (N_13563,N_11230,N_11587);
or U13564 (N_13564,N_11294,N_9410);
or U13565 (N_13565,N_11783,N_11790);
or U13566 (N_13566,N_9966,N_11176);
nor U13567 (N_13567,N_9435,N_10235);
nor U13568 (N_13568,N_11126,N_11352);
nand U13569 (N_13569,N_10959,N_10537);
or U13570 (N_13570,N_11969,N_11314);
and U13571 (N_13571,N_11269,N_9791);
or U13572 (N_13572,N_10910,N_10123);
or U13573 (N_13573,N_10140,N_11789);
or U13574 (N_13574,N_11017,N_9686);
or U13575 (N_13575,N_9673,N_9419);
or U13576 (N_13576,N_10058,N_11067);
nor U13577 (N_13577,N_9482,N_9512);
nor U13578 (N_13578,N_11690,N_10246);
nand U13579 (N_13579,N_9946,N_9909);
and U13580 (N_13580,N_9002,N_9827);
nor U13581 (N_13581,N_9458,N_10643);
nor U13582 (N_13582,N_11969,N_11435);
or U13583 (N_13583,N_10552,N_11448);
nand U13584 (N_13584,N_9662,N_10845);
nand U13585 (N_13585,N_11700,N_9697);
nand U13586 (N_13586,N_10714,N_9308);
or U13587 (N_13587,N_10706,N_10798);
nand U13588 (N_13588,N_11335,N_9763);
or U13589 (N_13589,N_9030,N_10075);
or U13590 (N_13590,N_11291,N_9539);
and U13591 (N_13591,N_10139,N_9191);
or U13592 (N_13592,N_10857,N_10779);
xnor U13593 (N_13593,N_9991,N_11186);
and U13594 (N_13594,N_10252,N_10198);
nor U13595 (N_13595,N_9905,N_9677);
and U13596 (N_13596,N_9568,N_10358);
nand U13597 (N_13597,N_11283,N_10359);
nor U13598 (N_13598,N_11129,N_9380);
or U13599 (N_13599,N_11846,N_11366);
and U13600 (N_13600,N_11554,N_10030);
nand U13601 (N_13601,N_11137,N_9602);
nor U13602 (N_13602,N_9504,N_11417);
xnor U13603 (N_13603,N_10257,N_10442);
and U13604 (N_13604,N_11977,N_9046);
nand U13605 (N_13605,N_10980,N_11636);
nand U13606 (N_13606,N_10874,N_10740);
nand U13607 (N_13607,N_10138,N_9285);
nand U13608 (N_13608,N_11895,N_9726);
nand U13609 (N_13609,N_10561,N_9710);
and U13610 (N_13610,N_11866,N_10417);
nand U13611 (N_13611,N_11151,N_11833);
nor U13612 (N_13612,N_11121,N_9708);
or U13613 (N_13613,N_11326,N_10264);
or U13614 (N_13614,N_10501,N_9556);
nor U13615 (N_13615,N_11281,N_11823);
and U13616 (N_13616,N_10974,N_9914);
or U13617 (N_13617,N_10935,N_10031);
nor U13618 (N_13618,N_10466,N_10899);
nand U13619 (N_13619,N_11967,N_9318);
nand U13620 (N_13620,N_11653,N_9550);
or U13621 (N_13621,N_11458,N_11636);
and U13622 (N_13622,N_10249,N_10132);
or U13623 (N_13623,N_10806,N_9423);
or U13624 (N_13624,N_10234,N_10737);
nand U13625 (N_13625,N_10410,N_9374);
and U13626 (N_13626,N_11448,N_10236);
and U13627 (N_13627,N_11316,N_10884);
xnor U13628 (N_13628,N_10079,N_10350);
or U13629 (N_13629,N_11958,N_9806);
and U13630 (N_13630,N_10670,N_11958);
and U13631 (N_13631,N_11523,N_11676);
and U13632 (N_13632,N_9328,N_10071);
or U13633 (N_13633,N_11041,N_10391);
or U13634 (N_13634,N_11834,N_9114);
nor U13635 (N_13635,N_9575,N_9538);
or U13636 (N_13636,N_11549,N_9700);
or U13637 (N_13637,N_10663,N_9063);
nand U13638 (N_13638,N_10758,N_10470);
and U13639 (N_13639,N_9929,N_9416);
nand U13640 (N_13640,N_9291,N_9564);
and U13641 (N_13641,N_11092,N_9332);
nor U13642 (N_13642,N_10545,N_10195);
and U13643 (N_13643,N_10987,N_11209);
nand U13644 (N_13644,N_10855,N_10518);
and U13645 (N_13645,N_10994,N_9870);
and U13646 (N_13646,N_9293,N_11913);
nand U13647 (N_13647,N_9824,N_11251);
nor U13648 (N_13648,N_11387,N_10883);
and U13649 (N_13649,N_9584,N_10203);
or U13650 (N_13650,N_11235,N_9646);
or U13651 (N_13651,N_9950,N_11412);
xor U13652 (N_13652,N_10456,N_9565);
and U13653 (N_13653,N_11456,N_11569);
nor U13654 (N_13654,N_10929,N_9167);
or U13655 (N_13655,N_10641,N_11574);
nand U13656 (N_13656,N_11343,N_11370);
and U13657 (N_13657,N_10776,N_10610);
nor U13658 (N_13658,N_9767,N_10747);
nor U13659 (N_13659,N_11079,N_9460);
nand U13660 (N_13660,N_9247,N_11877);
nand U13661 (N_13661,N_11648,N_9984);
nor U13662 (N_13662,N_9364,N_9200);
and U13663 (N_13663,N_11494,N_10304);
nand U13664 (N_13664,N_9690,N_9273);
nor U13665 (N_13665,N_9043,N_9228);
nand U13666 (N_13666,N_10745,N_10991);
nand U13667 (N_13667,N_9257,N_11002);
and U13668 (N_13668,N_9308,N_11602);
or U13669 (N_13669,N_10088,N_10126);
xnor U13670 (N_13670,N_10154,N_10116);
or U13671 (N_13671,N_11182,N_11105);
or U13672 (N_13672,N_9296,N_10497);
nor U13673 (N_13673,N_11373,N_9933);
or U13674 (N_13674,N_9271,N_11679);
and U13675 (N_13675,N_10592,N_9283);
or U13676 (N_13676,N_9714,N_9707);
and U13677 (N_13677,N_9819,N_11860);
or U13678 (N_13678,N_10927,N_9408);
nor U13679 (N_13679,N_10577,N_10845);
nor U13680 (N_13680,N_9520,N_11168);
and U13681 (N_13681,N_9947,N_9349);
nand U13682 (N_13682,N_11158,N_10748);
nor U13683 (N_13683,N_11952,N_9810);
nor U13684 (N_13684,N_11951,N_10018);
nor U13685 (N_13685,N_10197,N_9233);
nand U13686 (N_13686,N_9237,N_9044);
and U13687 (N_13687,N_11447,N_9264);
or U13688 (N_13688,N_11425,N_10084);
nand U13689 (N_13689,N_11144,N_11028);
nor U13690 (N_13690,N_10477,N_11013);
or U13691 (N_13691,N_11824,N_11940);
or U13692 (N_13692,N_9721,N_9165);
and U13693 (N_13693,N_11345,N_10633);
nor U13694 (N_13694,N_9608,N_10605);
and U13695 (N_13695,N_11369,N_9057);
nor U13696 (N_13696,N_10875,N_10269);
nand U13697 (N_13697,N_11526,N_11802);
xor U13698 (N_13698,N_9023,N_11228);
nor U13699 (N_13699,N_11231,N_10814);
nor U13700 (N_13700,N_9556,N_11083);
nand U13701 (N_13701,N_11400,N_11818);
nor U13702 (N_13702,N_10627,N_9637);
nand U13703 (N_13703,N_9293,N_10057);
nor U13704 (N_13704,N_9267,N_10706);
nor U13705 (N_13705,N_11000,N_9301);
nand U13706 (N_13706,N_10154,N_11009);
nand U13707 (N_13707,N_11950,N_11487);
xor U13708 (N_13708,N_11770,N_10939);
and U13709 (N_13709,N_10448,N_9878);
nor U13710 (N_13710,N_11817,N_11750);
nor U13711 (N_13711,N_10621,N_9139);
or U13712 (N_13712,N_10858,N_9615);
or U13713 (N_13713,N_9357,N_10897);
nor U13714 (N_13714,N_11532,N_11257);
nand U13715 (N_13715,N_11777,N_11857);
and U13716 (N_13716,N_9232,N_10168);
or U13717 (N_13717,N_10976,N_9590);
nand U13718 (N_13718,N_10378,N_11809);
nor U13719 (N_13719,N_10837,N_11685);
nand U13720 (N_13720,N_10424,N_11463);
and U13721 (N_13721,N_9217,N_11210);
or U13722 (N_13722,N_11130,N_11595);
and U13723 (N_13723,N_11917,N_11295);
or U13724 (N_13724,N_10594,N_9383);
or U13725 (N_13725,N_11923,N_11958);
nor U13726 (N_13726,N_9415,N_9066);
or U13727 (N_13727,N_9846,N_10727);
and U13728 (N_13728,N_10843,N_11265);
nand U13729 (N_13729,N_11306,N_9744);
nand U13730 (N_13730,N_11562,N_11771);
nor U13731 (N_13731,N_9457,N_10783);
and U13732 (N_13732,N_9009,N_11236);
and U13733 (N_13733,N_10423,N_10224);
and U13734 (N_13734,N_10137,N_10752);
xor U13735 (N_13735,N_11560,N_11829);
or U13736 (N_13736,N_9097,N_9707);
nor U13737 (N_13737,N_10599,N_9411);
nor U13738 (N_13738,N_11546,N_10157);
or U13739 (N_13739,N_9858,N_11037);
and U13740 (N_13740,N_9860,N_9760);
and U13741 (N_13741,N_9409,N_11386);
and U13742 (N_13742,N_9413,N_11479);
or U13743 (N_13743,N_11721,N_10529);
or U13744 (N_13744,N_10798,N_10756);
nand U13745 (N_13745,N_9525,N_10680);
or U13746 (N_13746,N_10998,N_10748);
and U13747 (N_13747,N_11204,N_10561);
nand U13748 (N_13748,N_11490,N_9564);
nand U13749 (N_13749,N_11881,N_10779);
nand U13750 (N_13750,N_11058,N_9662);
nand U13751 (N_13751,N_11033,N_11155);
nor U13752 (N_13752,N_11538,N_10178);
and U13753 (N_13753,N_9472,N_9813);
or U13754 (N_13754,N_9804,N_10957);
xnor U13755 (N_13755,N_11421,N_9109);
nand U13756 (N_13756,N_9253,N_9724);
nand U13757 (N_13757,N_10028,N_11522);
nand U13758 (N_13758,N_10914,N_9125);
nor U13759 (N_13759,N_9607,N_11608);
nand U13760 (N_13760,N_10161,N_10236);
or U13761 (N_13761,N_10846,N_9364);
nand U13762 (N_13762,N_9326,N_9938);
and U13763 (N_13763,N_10205,N_9198);
nor U13764 (N_13764,N_10959,N_11908);
nor U13765 (N_13765,N_9971,N_9830);
or U13766 (N_13766,N_10387,N_10472);
nor U13767 (N_13767,N_11175,N_11671);
or U13768 (N_13768,N_11410,N_9964);
nand U13769 (N_13769,N_11094,N_9489);
nor U13770 (N_13770,N_9641,N_9271);
and U13771 (N_13771,N_9425,N_9918);
and U13772 (N_13772,N_11821,N_11713);
or U13773 (N_13773,N_9228,N_11728);
nand U13774 (N_13774,N_10659,N_9358);
and U13775 (N_13775,N_10531,N_11925);
and U13776 (N_13776,N_10791,N_10282);
or U13777 (N_13777,N_11418,N_9004);
and U13778 (N_13778,N_9233,N_10572);
and U13779 (N_13779,N_11414,N_10133);
and U13780 (N_13780,N_9041,N_11886);
nand U13781 (N_13781,N_10370,N_9497);
or U13782 (N_13782,N_11957,N_10619);
nand U13783 (N_13783,N_10405,N_9320);
and U13784 (N_13784,N_11601,N_10234);
nand U13785 (N_13785,N_9645,N_11468);
and U13786 (N_13786,N_11302,N_11800);
nor U13787 (N_13787,N_10962,N_9458);
or U13788 (N_13788,N_9675,N_11715);
and U13789 (N_13789,N_11699,N_10691);
and U13790 (N_13790,N_9721,N_9991);
nand U13791 (N_13791,N_11871,N_9151);
nor U13792 (N_13792,N_10386,N_10581);
nor U13793 (N_13793,N_11839,N_11662);
nor U13794 (N_13794,N_10642,N_10390);
nor U13795 (N_13795,N_9052,N_9878);
nor U13796 (N_13796,N_10911,N_10218);
or U13797 (N_13797,N_11849,N_9502);
nand U13798 (N_13798,N_9805,N_10616);
or U13799 (N_13799,N_10220,N_9414);
or U13800 (N_13800,N_11073,N_9269);
or U13801 (N_13801,N_10520,N_11818);
and U13802 (N_13802,N_10588,N_11447);
nor U13803 (N_13803,N_11223,N_10822);
nor U13804 (N_13804,N_11928,N_9857);
or U13805 (N_13805,N_9505,N_9892);
nor U13806 (N_13806,N_10407,N_11893);
nor U13807 (N_13807,N_11639,N_11679);
nor U13808 (N_13808,N_11953,N_11167);
or U13809 (N_13809,N_10469,N_10186);
nand U13810 (N_13810,N_10510,N_10847);
nand U13811 (N_13811,N_9699,N_11738);
nor U13812 (N_13812,N_10470,N_10637);
or U13813 (N_13813,N_9954,N_10776);
and U13814 (N_13814,N_11150,N_9781);
or U13815 (N_13815,N_9336,N_11579);
nand U13816 (N_13816,N_10924,N_9539);
or U13817 (N_13817,N_11767,N_9943);
nand U13818 (N_13818,N_9262,N_11968);
and U13819 (N_13819,N_10778,N_10407);
nor U13820 (N_13820,N_9092,N_9955);
and U13821 (N_13821,N_10216,N_9655);
or U13822 (N_13822,N_9988,N_11706);
nor U13823 (N_13823,N_9117,N_11320);
nor U13824 (N_13824,N_10585,N_11833);
xnor U13825 (N_13825,N_9315,N_10132);
or U13826 (N_13826,N_11842,N_9858);
or U13827 (N_13827,N_10257,N_9769);
or U13828 (N_13828,N_10195,N_9363);
or U13829 (N_13829,N_11894,N_9655);
and U13830 (N_13830,N_10207,N_9504);
and U13831 (N_13831,N_9996,N_11054);
or U13832 (N_13832,N_9172,N_11729);
nor U13833 (N_13833,N_11691,N_10717);
and U13834 (N_13834,N_11416,N_11550);
and U13835 (N_13835,N_9294,N_11164);
and U13836 (N_13836,N_11881,N_9642);
and U13837 (N_13837,N_10799,N_9915);
xor U13838 (N_13838,N_11860,N_10009);
xor U13839 (N_13839,N_10908,N_10717);
nor U13840 (N_13840,N_9634,N_9530);
or U13841 (N_13841,N_11825,N_11397);
nand U13842 (N_13842,N_10400,N_10654);
or U13843 (N_13843,N_10669,N_10985);
and U13844 (N_13844,N_10967,N_9235);
nor U13845 (N_13845,N_9756,N_11740);
nor U13846 (N_13846,N_9619,N_9210);
nor U13847 (N_13847,N_9889,N_11154);
nor U13848 (N_13848,N_9309,N_11977);
and U13849 (N_13849,N_10525,N_9679);
nor U13850 (N_13850,N_9851,N_10198);
and U13851 (N_13851,N_11948,N_11735);
and U13852 (N_13852,N_10685,N_10422);
and U13853 (N_13853,N_11801,N_9130);
or U13854 (N_13854,N_11247,N_9771);
and U13855 (N_13855,N_10171,N_11027);
and U13856 (N_13856,N_10803,N_9673);
nand U13857 (N_13857,N_10664,N_10412);
or U13858 (N_13858,N_10867,N_9496);
and U13859 (N_13859,N_9114,N_9527);
nand U13860 (N_13860,N_10398,N_11790);
or U13861 (N_13861,N_9686,N_9821);
nand U13862 (N_13862,N_10004,N_9714);
or U13863 (N_13863,N_10555,N_10314);
and U13864 (N_13864,N_9691,N_11886);
and U13865 (N_13865,N_9025,N_11259);
and U13866 (N_13866,N_10128,N_9643);
or U13867 (N_13867,N_9875,N_10017);
or U13868 (N_13868,N_10929,N_11604);
nand U13869 (N_13869,N_9158,N_9159);
or U13870 (N_13870,N_10519,N_10057);
xor U13871 (N_13871,N_10005,N_9677);
nor U13872 (N_13872,N_9676,N_11264);
nand U13873 (N_13873,N_9224,N_10103);
nor U13874 (N_13874,N_9194,N_10708);
nor U13875 (N_13875,N_10663,N_10889);
or U13876 (N_13876,N_10306,N_9076);
nand U13877 (N_13877,N_11016,N_10216);
and U13878 (N_13878,N_11519,N_9111);
nand U13879 (N_13879,N_11618,N_11965);
or U13880 (N_13880,N_9921,N_9894);
or U13881 (N_13881,N_9542,N_11960);
nand U13882 (N_13882,N_10621,N_11832);
xnor U13883 (N_13883,N_10371,N_10796);
and U13884 (N_13884,N_11644,N_9538);
nand U13885 (N_13885,N_11162,N_10678);
nor U13886 (N_13886,N_11050,N_9417);
nor U13887 (N_13887,N_9282,N_10867);
and U13888 (N_13888,N_10418,N_9793);
nor U13889 (N_13889,N_11615,N_10259);
nor U13890 (N_13890,N_10811,N_10541);
nand U13891 (N_13891,N_9382,N_9042);
and U13892 (N_13892,N_9144,N_10887);
nand U13893 (N_13893,N_9408,N_11527);
nor U13894 (N_13894,N_9221,N_10200);
nor U13895 (N_13895,N_9952,N_10689);
nand U13896 (N_13896,N_10567,N_10612);
or U13897 (N_13897,N_9627,N_9689);
nand U13898 (N_13898,N_9358,N_11344);
and U13899 (N_13899,N_11656,N_9846);
nand U13900 (N_13900,N_11446,N_9299);
or U13901 (N_13901,N_11387,N_11830);
nor U13902 (N_13902,N_10667,N_10015);
nor U13903 (N_13903,N_11079,N_9858);
nor U13904 (N_13904,N_11825,N_9179);
or U13905 (N_13905,N_11231,N_11095);
or U13906 (N_13906,N_11112,N_9431);
or U13907 (N_13907,N_10273,N_11042);
and U13908 (N_13908,N_10604,N_9263);
nor U13909 (N_13909,N_10490,N_10105);
and U13910 (N_13910,N_11245,N_10399);
or U13911 (N_13911,N_10818,N_9356);
nand U13912 (N_13912,N_10706,N_11170);
nor U13913 (N_13913,N_9608,N_9036);
nand U13914 (N_13914,N_10684,N_10140);
xor U13915 (N_13915,N_10598,N_10109);
and U13916 (N_13916,N_10882,N_9025);
or U13917 (N_13917,N_11211,N_9728);
nor U13918 (N_13918,N_10882,N_10839);
nor U13919 (N_13919,N_10308,N_9162);
and U13920 (N_13920,N_11649,N_9542);
or U13921 (N_13921,N_9161,N_10269);
or U13922 (N_13922,N_11923,N_9850);
nand U13923 (N_13923,N_10290,N_9538);
nand U13924 (N_13924,N_10066,N_11552);
nand U13925 (N_13925,N_10969,N_9570);
or U13926 (N_13926,N_9302,N_10088);
or U13927 (N_13927,N_9518,N_9656);
or U13928 (N_13928,N_10138,N_10483);
and U13929 (N_13929,N_10952,N_10420);
nor U13930 (N_13930,N_9199,N_9758);
nand U13931 (N_13931,N_11986,N_9007);
nor U13932 (N_13932,N_11511,N_9075);
or U13933 (N_13933,N_10929,N_11893);
or U13934 (N_13934,N_9202,N_11629);
nor U13935 (N_13935,N_11532,N_11881);
nand U13936 (N_13936,N_11684,N_10256);
or U13937 (N_13937,N_11613,N_9083);
xnor U13938 (N_13938,N_9678,N_10099);
and U13939 (N_13939,N_9761,N_10157);
and U13940 (N_13940,N_9360,N_11254);
nand U13941 (N_13941,N_9800,N_11523);
and U13942 (N_13942,N_9645,N_10104);
and U13943 (N_13943,N_11755,N_10742);
nand U13944 (N_13944,N_9139,N_11405);
or U13945 (N_13945,N_11396,N_11285);
nor U13946 (N_13946,N_9066,N_11863);
or U13947 (N_13947,N_9615,N_11549);
nand U13948 (N_13948,N_9353,N_9229);
or U13949 (N_13949,N_10235,N_9953);
and U13950 (N_13950,N_9925,N_11316);
or U13951 (N_13951,N_10019,N_11571);
nand U13952 (N_13952,N_9876,N_10748);
nor U13953 (N_13953,N_11960,N_10412);
nand U13954 (N_13954,N_9269,N_11048);
or U13955 (N_13955,N_10819,N_11493);
or U13956 (N_13956,N_11663,N_11630);
nand U13957 (N_13957,N_9271,N_10048);
and U13958 (N_13958,N_11533,N_9507);
nand U13959 (N_13959,N_9774,N_9711);
or U13960 (N_13960,N_9671,N_11053);
nand U13961 (N_13961,N_10512,N_11155);
or U13962 (N_13962,N_9924,N_11979);
nor U13963 (N_13963,N_10644,N_11327);
or U13964 (N_13964,N_9177,N_10186);
and U13965 (N_13965,N_10521,N_11042);
or U13966 (N_13966,N_10412,N_10229);
nor U13967 (N_13967,N_11336,N_11223);
and U13968 (N_13968,N_11052,N_10257);
xor U13969 (N_13969,N_10636,N_10911);
nand U13970 (N_13970,N_11890,N_9410);
and U13971 (N_13971,N_9589,N_10442);
or U13972 (N_13972,N_10209,N_10126);
nor U13973 (N_13973,N_11622,N_10608);
nor U13974 (N_13974,N_9199,N_10255);
nand U13975 (N_13975,N_11330,N_11530);
nand U13976 (N_13976,N_9423,N_9272);
or U13977 (N_13977,N_9395,N_9391);
nor U13978 (N_13978,N_9998,N_10171);
or U13979 (N_13979,N_10736,N_10467);
nand U13980 (N_13980,N_9630,N_10916);
nand U13981 (N_13981,N_9747,N_11561);
or U13982 (N_13982,N_9329,N_11180);
or U13983 (N_13983,N_9862,N_9221);
and U13984 (N_13984,N_10855,N_11835);
nor U13985 (N_13985,N_10313,N_10624);
and U13986 (N_13986,N_11893,N_11037);
nor U13987 (N_13987,N_9289,N_9515);
nor U13988 (N_13988,N_11696,N_10432);
nor U13989 (N_13989,N_11288,N_10871);
nor U13990 (N_13990,N_11066,N_10560);
or U13991 (N_13991,N_9126,N_9526);
or U13992 (N_13992,N_10435,N_10611);
or U13993 (N_13993,N_9123,N_11069);
nand U13994 (N_13994,N_11772,N_11182);
and U13995 (N_13995,N_10785,N_9611);
nand U13996 (N_13996,N_11734,N_9851);
nand U13997 (N_13997,N_11835,N_11552);
and U13998 (N_13998,N_9637,N_11738);
nand U13999 (N_13999,N_9696,N_11039);
nor U14000 (N_14000,N_9184,N_10742);
and U14001 (N_14001,N_11603,N_9885);
and U14002 (N_14002,N_11018,N_9512);
or U14003 (N_14003,N_9224,N_9899);
and U14004 (N_14004,N_10771,N_11494);
nand U14005 (N_14005,N_9002,N_10044);
and U14006 (N_14006,N_9005,N_11001);
nor U14007 (N_14007,N_10345,N_10644);
nand U14008 (N_14008,N_9866,N_9146);
nand U14009 (N_14009,N_9370,N_9080);
or U14010 (N_14010,N_11523,N_10400);
or U14011 (N_14011,N_10336,N_9567);
nor U14012 (N_14012,N_10458,N_9243);
nor U14013 (N_14013,N_11125,N_9433);
or U14014 (N_14014,N_9438,N_10064);
or U14015 (N_14015,N_9674,N_9801);
and U14016 (N_14016,N_9993,N_10363);
nand U14017 (N_14017,N_9011,N_11295);
or U14018 (N_14018,N_9774,N_11853);
or U14019 (N_14019,N_10681,N_11328);
or U14020 (N_14020,N_11146,N_9331);
nand U14021 (N_14021,N_11328,N_10047);
nor U14022 (N_14022,N_11948,N_10674);
xnor U14023 (N_14023,N_9269,N_11303);
nand U14024 (N_14024,N_10177,N_10484);
nor U14025 (N_14025,N_11214,N_9933);
or U14026 (N_14026,N_11108,N_10818);
nor U14027 (N_14027,N_11089,N_9019);
nor U14028 (N_14028,N_10120,N_10233);
and U14029 (N_14029,N_10592,N_9660);
and U14030 (N_14030,N_11549,N_10873);
xnor U14031 (N_14031,N_11568,N_10684);
nor U14032 (N_14032,N_10809,N_11505);
or U14033 (N_14033,N_10189,N_9851);
and U14034 (N_14034,N_9962,N_11753);
nand U14035 (N_14035,N_9932,N_11230);
nor U14036 (N_14036,N_11612,N_9432);
xor U14037 (N_14037,N_10901,N_11590);
or U14038 (N_14038,N_10352,N_9666);
and U14039 (N_14039,N_11957,N_10730);
nand U14040 (N_14040,N_11667,N_10572);
or U14041 (N_14041,N_9912,N_10836);
nand U14042 (N_14042,N_10194,N_11852);
or U14043 (N_14043,N_9063,N_9305);
nor U14044 (N_14044,N_10712,N_11280);
nand U14045 (N_14045,N_11550,N_11025);
nand U14046 (N_14046,N_11587,N_10716);
or U14047 (N_14047,N_10532,N_11932);
nor U14048 (N_14048,N_11719,N_10616);
and U14049 (N_14049,N_9744,N_11135);
nand U14050 (N_14050,N_9387,N_10306);
or U14051 (N_14051,N_11711,N_9414);
or U14052 (N_14052,N_10322,N_10604);
or U14053 (N_14053,N_11856,N_10982);
nand U14054 (N_14054,N_10252,N_10096);
or U14055 (N_14055,N_10383,N_10048);
nor U14056 (N_14056,N_10197,N_10784);
nand U14057 (N_14057,N_9628,N_9909);
nor U14058 (N_14058,N_11809,N_11714);
nor U14059 (N_14059,N_10622,N_10794);
nand U14060 (N_14060,N_11679,N_10040);
xnor U14061 (N_14061,N_10165,N_10604);
and U14062 (N_14062,N_9125,N_10068);
nand U14063 (N_14063,N_9314,N_9624);
or U14064 (N_14064,N_11693,N_9676);
or U14065 (N_14065,N_11967,N_9126);
nor U14066 (N_14066,N_10954,N_9983);
or U14067 (N_14067,N_11366,N_10573);
nand U14068 (N_14068,N_11486,N_11030);
or U14069 (N_14069,N_10372,N_10111);
nor U14070 (N_14070,N_9532,N_10955);
nor U14071 (N_14071,N_11698,N_9479);
nor U14072 (N_14072,N_11510,N_10612);
and U14073 (N_14073,N_10849,N_9245);
nor U14074 (N_14074,N_11626,N_10292);
or U14075 (N_14075,N_11743,N_10557);
nand U14076 (N_14076,N_10435,N_10807);
and U14077 (N_14077,N_9873,N_11141);
nand U14078 (N_14078,N_9589,N_11362);
nand U14079 (N_14079,N_10849,N_11444);
and U14080 (N_14080,N_9782,N_10557);
nand U14081 (N_14081,N_9128,N_10923);
and U14082 (N_14082,N_11194,N_10715);
nor U14083 (N_14083,N_11444,N_9690);
nand U14084 (N_14084,N_9053,N_9382);
or U14085 (N_14085,N_11579,N_10068);
and U14086 (N_14086,N_11970,N_9939);
and U14087 (N_14087,N_10883,N_11914);
and U14088 (N_14088,N_10757,N_9798);
nand U14089 (N_14089,N_11164,N_11965);
or U14090 (N_14090,N_10216,N_10634);
nand U14091 (N_14091,N_10874,N_9158);
nor U14092 (N_14092,N_9149,N_11055);
and U14093 (N_14093,N_9287,N_9245);
nor U14094 (N_14094,N_11502,N_9451);
nor U14095 (N_14095,N_9678,N_11314);
nand U14096 (N_14096,N_10494,N_9570);
or U14097 (N_14097,N_9239,N_10842);
and U14098 (N_14098,N_10382,N_9182);
and U14099 (N_14099,N_10710,N_11604);
or U14100 (N_14100,N_10159,N_11086);
and U14101 (N_14101,N_10479,N_9948);
nor U14102 (N_14102,N_10266,N_10262);
nand U14103 (N_14103,N_9706,N_10263);
nor U14104 (N_14104,N_9477,N_10783);
nor U14105 (N_14105,N_9095,N_10117);
and U14106 (N_14106,N_11341,N_9390);
and U14107 (N_14107,N_9766,N_11036);
nor U14108 (N_14108,N_11403,N_10015);
and U14109 (N_14109,N_11310,N_11347);
nor U14110 (N_14110,N_10260,N_11693);
nor U14111 (N_14111,N_11233,N_9674);
nor U14112 (N_14112,N_11623,N_11034);
and U14113 (N_14113,N_10026,N_9146);
or U14114 (N_14114,N_9726,N_9442);
and U14115 (N_14115,N_11467,N_11950);
nor U14116 (N_14116,N_10401,N_9703);
nand U14117 (N_14117,N_9361,N_10027);
or U14118 (N_14118,N_11817,N_11556);
nand U14119 (N_14119,N_11426,N_9186);
or U14120 (N_14120,N_9574,N_9231);
or U14121 (N_14121,N_11923,N_9551);
or U14122 (N_14122,N_9055,N_11374);
nand U14123 (N_14123,N_10496,N_10507);
or U14124 (N_14124,N_10105,N_10545);
xnor U14125 (N_14125,N_9837,N_10011);
and U14126 (N_14126,N_11597,N_9193);
nor U14127 (N_14127,N_9807,N_11117);
nor U14128 (N_14128,N_11451,N_9956);
or U14129 (N_14129,N_10762,N_11830);
nand U14130 (N_14130,N_10117,N_9950);
nand U14131 (N_14131,N_9409,N_10433);
or U14132 (N_14132,N_9559,N_9565);
nor U14133 (N_14133,N_10800,N_10233);
nand U14134 (N_14134,N_11784,N_9518);
xnor U14135 (N_14135,N_10687,N_9009);
nand U14136 (N_14136,N_9143,N_9918);
or U14137 (N_14137,N_11145,N_11889);
nor U14138 (N_14138,N_11268,N_11147);
nand U14139 (N_14139,N_10145,N_9082);
nand U14140 (N_14140,N_10273,N_9083);
nor U14141 (N_14141,N_11753,N_10274);
nand U14142 (N_14142,N_11383,N_10569);
nor U14143 (N_14143,N_11915,N_10579);
or U14144 (N_14144,N_10846,N_9620);
nor U14145 (N_14145,N_9059,N_11126);
nand U14146 (N_14146,N_11424,N_11511);
or U14147 (N_14147,N_9380,N_9471);
nor U14148 (N_14148,N_10292,N_9385);
xnor U14149 (N_14149,N_11673,N_10522);
and U14150 (N_14150,N_10332,N_10009);
and U14151 (N_14151,N_11027,N_10732);
nor U14152 (N_14152,N_9415,N_10204);
nor U14153 (N_14153,N_10219,N_10399);
nor U14154 (N_14154,N_9818,N_10515);
nor U14155 (N_14155,N_11638,N_10198);
or U14156 (N_14156,N_10468,N_9526);
nor U14157 (N_14157,N_10717,N_10688);
nand U14158 (N_14158,N_11356,N_9450);
nand U14159 (N_14159,N_11180,N_9356);
or U14160 (N_14160,N_10834,N_10150);
or U14161 (N_14161,N_10712,N_10157);
and U14162 (N_14162,N_11239,N_9426);
nor U14163 (N_14163,N_9715,N_10568);
and U14164 (N_14164,N_10189,N_9034);
nor U14165 (N_14165,N_11868,N_10634);
and U14166 (N_14166,N_10434,N_11837);
nor U14167 (N_14167,N_10493,N_11602);
nor U14168 (N_14168,N_9315,N_10698);
nand U14169 (N_14169,N_10123,N_10620);
and U14170 (N_14170,N_10413,N_11868);
nor U14171 (N_14171,N_10180,N_9366);
and U14172 (N_14172,N_11468,N_9717);
nand U14173 (N_14173,N_9452,N_9323);
or U14174 (N_14174,N_9805,N_9211);
or U14175 (N_14175,N_9733,N_11757);
nand U14176 (N_14176,N_10945,N_11191);
nand U14177 (N_14177,N_11269,N_9162);
nor U14178 (N_14178,N_9062,N_10528);
nor U14179 (N_14179,N_10283,N_10199);
and U14180 (N_14180,N_11337,N_11869);
and U14181 (N_14181,N_10689,N_11097);
and U14182 (N_14182,N_10544,N_10228);
or U14183 (N_14183,N_9880,N_9524);
or U14184 (N_14184,N_9155,N_9863);
nor U14185 (N_14185,N_9326,N_9009);
and U14186 (N_14186,N_11122,N_10191);
nand U14187 (N_14187,N_9943,N_9364);
nand U14188 (N_14188,N_9616,N_11369);
or U14189 (N_14189,N_9133,N_11772);
or U14190 (N_14190,N_9445,N_11915);
nor U14191 (N_14191,N_9616,N_9778);
nand U14192 (N_14192,N_9189,N_9691);
and U14193 (N_14193,N_10698,N_9560);
and U14194 (N_14194,N_9569,N_11017);
nor U14195 (N_14195,N_10139,N_11740);
or U14196 (N_14196,N_11251,N_11800);
xnor U14197 (N_14197,N_9124,N_11559);
nor U14198 (N_14198,N_11733,N_9827);
xnor U14199 (N_14199,N_11793,N_10667);
nand U14200 (N_14200,N_10056,N_11107);
or U14201 (N_14201,N_11225,N_9598);
nor U14202 (N_14202,N_10894,N_10058);
nand U14203 (N_14203,N_11657,N_10746);
and U14204 (N_14204,N_10075,N_11183);
or U14205 (N_14205,N_11778,N_9354);
and U14206 (N_14206,N_10076,N_9936);
and U14207 (N_14207,N_11894,N_10378);
nor U14208 (N_14208,N_9326,N_9317);
nor U14209 (N_14209,N_10958,N_11041);
and U14210 (N_14210,N_10606,N_9569);
nand U14211 (N_14211,N_10263,N_9494);
or U14212 (N_14212,N_11104,N_9299);
or U14213 (N_14213,N_9410,N_10133);
nand U14214 (N_14214,N_11688,N_10792);
nor U14215 (N_14215,N_9453,N_9870);
nand U14216 (N_14216,N_10747,N_10666);
nor U14217 (N_14217,N_10566,N_9681);
and U14218 (N_14218,N_9693,N_11134);
nand U14219 (N_14219,N_11744,N_10576);
nand U14220 (N_14220,N_10224,N_9151);
or U14221 (N_14221,N_9766,N_9314);
or U14222 (N_14222,N_9177,N_9042);
nand U14223 (N_14223,N_11940,N_11232);
nor U14224 (N_14224,N_11685,N_11563);
or U14225 (N_14225,N_10136,N_11517);
and U14226 (N_14226,N_9266,N_11054);
or U14227 (N_14227,N_9772,N_9192);
or U14228 (N_14228,N_9400,N_11399);
or U14229 (N_14229,N_9584,N_10045);
nand U14230 (N_14230,N_9524,N_11438);
xnor U14231 (N_14231,N_10335,N_9458);
nor U14232 (N_14232,N_9969,N_11684);
and U14233 (N_14233,N_10958,N_11218);
and U14234 (N_14234,N_10025,N_10823);
nand U14235 (N_14235,N_10648,N_9193);
nand U14236 (N_14236,N_9988,N_11218);
or U14237 (N_14237,N_11293,N_11546);
nand U14238 (N_14238,N_10863,N_11310);
or U14239 (N_14239,N_10672,N_10843);
nor U14240 (N_14240,N_9193,N_10645);
xnor U14241 (N_14241,N_10008,N_9539);
and U14242 (N_14242,N_9129,N_10585);
or U14243 (N_14243,N_9358,N_10620);
nand U14244 (N_14244,N_9186,N_10698);
nand U14245 (N_14245,N_11604,N_9591);
or U14246 (N_14246,N_9586,N_10358);
nand U14247 (N_14247,N_9683,N_9692);
nand U14248 (N_14248,N_10802,N_10832);
or U14249 (N_14249,N_11316,N_11456);
nand U14250 (N_14250,N_10029,N_11719);
and U14251 (N_14251,N_9684,N_11876);
nor U14252 (N_14252,N_9280,N_11672);
and U14253 (N_14253,N_11267,N_11763);
nand U14254 (N_14254,N_9691,N_10272);
and U14255 (N_14255,N_11992,N_11599);
nor U14256 (N_14256,N_11462,N_11890);
nor U14257 (N_14257,N_10624,N_11525);
xnor U14258 (N_14258,N_9316,N_9714);
or U14259 (N_14259,N_9686,N_11129);
or U14260 (N_14260,N_10521,N_9722);
nand U14261 (N_14261,N_9419,N_9006);
or U14262 (N_14262,N_11959,N_9779);
and U14263 (N_14263,N_10975,N_9233);
nor U14264 (N_14264,N_11493,N_11358);
or U14265 (N_14265,N_11487,N_11145);
nand U14266 (N_14266,N_10649,N_9381);
nor U14267 (N_14267,N_10516,N_9427);
and U14268 (N_14268,N_9033,N_11873);
nor U14269 (N_14269,N_11938,N_11952);
or U14270 (N_14270,N_10280,N_10090);
or U14271 (N_14271,N_11656,N_9749);
and U14272 (N_14272,N_10810,N_11632);
and U14273 (N_14273,N_11666,N_11779);
or U14274 (N_14274,N_10493,N_11210);
or U14275 (N_14275,N_11993,N_11161);
or U14276 (N_14276,N_11083,N_9584);
and U14277 (N_14277,N_9984,N_10576);
nand U14278 (N_14278,N_11894,N_9882);
nor U14279 (N_14279,N_11241,N_10135);
and U14280 (N_14280,N_9785,N_10576);
or U14281 (N_14281,N_11301,N_9104);
nor U14282 (N_14282,N_11452,N_9176);
and U14283 (N_14283,N_10516,N_11784);
and U14284 (N_14284,N_9584,N_10388);
or U14285 (N_14285,N_10148,N_10240);
and U14286 (N_14286,N_11318,N_9677);
and U14287 (N_14287,N_9063,N_9167);
or U14288 (N_14288,N_9798,N_10646);
nor U14289 (N_14289,N_11623,N_11341);
or U14290 (N_14290,N_9527,N_11673);
or U14291 (N_14291,N_10219,N_11081);
nor U14292 (N_14292,N_9703,N_10128);
and U14293 (N_14293,N_11621,N_9193);
nand U14294 (N_14294,N_10674,N_9988);
nor U14295 (N_14295,N_10283,N_9842);
and U14296 (N_14296,N_9721,N_11776);
nor U14297 (N_14297,N_9875,N_10697);
nand U14298 (N_14298,N_9378,N_11067);
nand U14299 (N_14299,N_10615,N_11293);
and U14300 (N_14300,N_9635,N_9262);
nand U14301 (N_14301,N_10549,N_10495);
xor U14302 (N_14302,N_11321,N_9915);
nand U14303 (N_14303,N_10082,N_10181);
nand U14304 (N_14304,N_10633,N_9328);
xor U14305 (N_14305,N_9098,N_10745);
and U14306 (N_14306,N_10451,N_10294);
or U14307 (N_14307,N_10294,N_10873);
or U14308 (N_14308,N_11695,N_11082);
or U14309 (N_14309,N_10759,N_10995);
nor U14310 (N_14310,N_10112,N_9152);
nor U14311 (N_14311,N_10055,N_9495);
nand U14312 (N_14312,N_11658,N_9783);
nand U14313 (N_14313,N_9716,N_11871);
nor U14314 (N_14314,N_10392,N_9558);
or U14315 (N_14315,N_9890,N_9620);
and U14316 (N_14316,N_9009,N_9759);
nor U14317 (N_14317,N_11022,N_9972);
or U14318 (N_14318,N_11252,N_11521);
or U14319 (N_14319,N_10734,N_10496);
and U14320 (N_14320,N_11767,N_10797);
and U14321 (N_14321,N_9832,N_10473);
nor U14322 (N_14322,N_9071,N_11290);
or U14323 (N_14323,N_9913,N_11546);
or U14324 (N_14324,N_11013,N_11317);
and U14325 (N_14325,N_9357,N_10752);
or U14326 (N_14326,N_10449,N_9762);
and U14327 (N_14327,N_10473,N_9033);
nor U14328 (N_14328,N_9035,N_10888);
and U14329 (N_14329,N_9561,N_11622);
nand U14330 (N_14330,N_11372,N_9229);
nor U14331 (N_14331,N_9062,N_9492);
nor U14332 (N_14332,N_9784,N_9628);
or U14333 (N_14333,N_11465,N_9719);
nand U14334 (N_14334,N_11792,N_10472);
and U14335 (N_14335,N_9849,N_10231);
or U14336 (N_14336,N_9670,N_11436);
nand U14337 (N_14337,N_11132,N_10005);
and U14338 (N_14338,N_10323,N_9553);
and U14339 (N_14339,N_9145,N_9666);
nor U14340 (N_14340,N_10520,N_10273);
or U14341 (N_14341,N_10664,N_10173);
nand U14342 (N_14342,N_11520,N_9999);
nor U14343 (N_14343,N_9613,N_10803);
or U14344 (N_14344,N_10938,N_11515);
and U14345 (N_14345,N_11907,N_10382);
and U14346 (N_14346,N_10911,N_9044);
xnor U14347 (N_14347,N_9240,N_11568);
or U14348 (N_14348,N_11876,N_9381);
nand U14349 (N_14349,N_11401,N_10939);
nand U14350 (N_14350,N_11494,N_11511);
nor U14351 (N_14351,N_9220,N_9543);
nand U14352 (N_14352,N_11514,N_11117);
or U14353 (N_14353,N_10497,N_9705);
nand U14354 (N_14354,N_9723,N_11836);
nor U14355 (N_14355,N_9346,N_11282);
and U14356 (N_14356,N_9258,N_10041);
or U14357 (N_14357,N_9222,N_11745);
nand U14358 (N_14358,N_9378,N_9065);
nor U14359 (N_14359,N_10693,N_10550);
nor U14360 (N_14360,N_9160,N_9017);
or U14361 (N_14361,N_11983,N_11659);
nand U14362 (N_14362,N_9608,N_9294);
and U14363 (N_14363,N_11868,N_9839);
or U14364 (N_14364,N_11049,N_11770);
or U14365 (N_14365,N_11219,N_11714);
and U14366 (N_14366,N_9163,N_9036);
and U14367 (N_14367,N_10188,N_9799);
nand U14368 (N_14368,N_11074,N_10102);
and U14369 (N_14369,N_9639,N_10119);
nand U14370 (N_14370,N_11812,N_10663);
or U14371 (N_14371,N_10405,N_9770);
nand U14372 (N_14372,N_11214,N_11345);
nand U14373 (N_14373,N_10281,N_10489);
nand U14374 (N_14374,N_9760,N_10960);
nor U14375 (N_14375,N_11089,N_11664);
or U14376 (N_14376,N_9185,N_9251);
nand U14377 (N_14377,N_11851,N_9775);
nor U14378 (N_14378,N_9078,N_10323);
nand U14379 (N_14379,N_11107,N_11706);
nand U14380 (N_14380,N_11858,N_10735);
or U14381 (N_14381,N_11375,N_9211);
nand U14382 (N_14382,N_9266,N_9101);
and U14383 (N_14383,N_11333,N_9493);
and U14384 (N_14384,N_9110,N_9390);
nor U14385 (N_14385,N_11756,N_11869);
and U14386 (N_14386,N_10130,N_10359);
nand U14387 (N_14387,N_11246,N_9136);
nand U14388 (N_14388,N_10712,N_10477);
and U14389 (N_14389,N_9905,N_10123);
nor U14390 (N_14390,N_9739,N_11232);
or U14391 (N_14391,N_9385,N_9043);
or U14392 (N_14392,N_10327,N_11891);
and U14393 (N_14393,N_10433,N_10025);
nand U14394 (N_14394,N_10415,N_11736);
nand U14395 (N_14395,N_9871,N_11896);
nand U14396 (N_14396,N_9319,N_10004);
nand U14397 (N_14397,N_10157,N_9959);
or U14398 (N_14398,N_11001,N_9942);
nor U14399 (N_14399,N_9973,N_9017);
nor U14400 (N_14400,N_9242,N_9250);
or U14401 (N_14401,N_10129,N_9357);
or U14402 (N_14402,N_10372,N_9550);
or U14403 (N_14403,N_10846,N_10792);
nand U14404 (N_14404,N_11203,N_9518);
nand U14405 (N_14405,N_10430,N_9197);
and U14406 (N_14406,N_9493,N_11698);
nand U14407 (N_14407,N_9648,N_9176);
xor U14408 (N_14408,N_11575,N_11517);
nor U14409 (N_14409,N_10124,N_9531);
nor U14410 (N_14410,N_11768,N_11433);
nor U14411 (N_14411,N_10804,N_9256);
nor U14412 (N_14412,N_9745,N_10319);
or U14413 (N_14413,N_9411,N_11608);
nor U14414 (N_14414,N_10216,N_11602);
nand U14415 (N_14415,N_11545,N_11098);
or U14416 (N_14416,N_9975,N_10434);
nand U14417 (N_14417,N_10020,N_10514);
and U14418 (N_14418,N_11127,N_9883);
nand U14419 (N_14419,N_9801,N_10048);
nor U14420 (N_14420,N_11221,N_10808);
and U14421 (N_14421,N_9554,N_11634);
and U14422 (N_14422,N_9993,N_9128);
nand U14423 (N_14423,N_9758,N_10146);
nand U14424 (N_14424,N_11471,N_10981);
and U14425 (N_14425,N_9711,N_10918);
nand U14426 (N_14426,N_10147,N_11600);
and U14427 (N_14427,N_10757,N_10968);
nand U14428 (N_14428,N_10216,N_9149);
and U14429 (N_14429,N_11237,N_11335);
and U14430 (N_14430,N_9075,N_10816);
nand U14431 (N_14431,N_11770,N_11124);
and U14432 (N_14432,N_9060,N_11668);
and U14433 (N_14433,N_9360,N_11148);
nor U14434 (N_14434,N_10906,N_9158);
and U14435 (N_14435,N_10315,N_11712);
nor U14436 (N_14436,N_9173,N_9611);
nor U14437 (N_14437,N_11106,N_10256);
or U14438 (N_14438,N_9667,N_10706);
nand U14439 (N_14439,N_10900,N_11119);
or U14440 (N_14440,N_9056,N_11065);
nor U14441 (N_14441,N_9849,N_10015);
and U14442 (N_14442,N_9039,N_9801);
nor U14443 (N_14443,N_11319,N_10363);
xor U14444 (N_14444,N_10387,N_10722);
and U14445 (N_14445,N_10495,N_10385);
nand U14446 (N_14446,N_11506,N_11198);
nor U14447 (N_14447,N_11631,N_11008);
and U14448 (N_14448,N_10588,N_11509);
nand U14449 (N_14449,N_11159,N_11707);
and U14450 (N_14450,N_9314,N_10693);
nand U14451 (N_14451,N_9263,N_10760);
and U14452 (N_14452,N_11003,N_9582);
nor U14453 (N_14453,N_11966,N_9870);
or U14454 (N_14454,N_11653,N_10181);
or U14455 (N_14455,N_9264,N_10614);
nor U14456 (N_14456,N_10252,N_9743);
nand U14457 (N_14457,N_10411,N_10828);
or U14458 (N_14458,N_10533,N_9979);
nand U14459 (N_14459,N_9679,N_11245);
nor U14460 (N_14460,N_11610,N_9917);
nor U14461 (N_14461,N_11052,N_9199);
and U14462 (N_14462,N_11873,N_11236);
and U14463 (N_14463,N_11359,N_11847);
nor U14464 (N_14464,N_10756,N_9431);
and U14465 (N_14465,N_9203,N_9279);
nor U14466 (N_14466,N_9311,N_10475);
nand U14467 (N_14467,N_11116,N_11608);
nand U14468 (N_14468,N_11257,N_10790);
nor U14469 (N_14469,N_11860,N_9070);
nor U14470 (N_14470,N_10847,N_10630);
nand U14471 (N_14471,N_9459,N_11365);
nand U14472 (N_14472,N_11534,N_10000);
nand U14473 (N_14473,N_9562,N_11402);
nor U14474 (N_14474,N_11142,N_11568);
nor U14475 (N_14475,N_10388,N_9612);
nor U14476 (N_14476,N_10498,N_11370);
nand U14477 (N_14477,N_9513,N_9732);
or U14478 (N_14478,N_10502,N_10121);
or U14479 (N_14479,N_9957,N_10559);
or U14480 (N_14480,N_9066,N_11041);
and U14481 (N_14481,N_10746,N_9997);
nand U14482 (N_14482,N_11609,N_10443);
nor U14483 (N_14483,N_11008,N_9618);
and U14484 (N_14484,N_9150,N_11869);
nor U14485 (N_14485,N_10023,N_9727);
nand U14486 (N_14486,N_9689,N_11084);
or U14487 (N_14487,N_11150,N_10624);
or U14488 (N_14488,N_9495,N_11965);
nand U14489 (N_14489,N_10797,N_9257);
nand U14490 (N_14490,N_9347,N_10208);
or U14491 (N_14491,N_11582,N_9765);
or U14492 (N_14492,N_9085,N_11860);
or U14493 (N_14493,N_9539,N_10121);
nand U14494 (N_14494,N_9419,N_9960);
nand U14495 (N_14495,N_10927,N_11673);
or U14496 (N_14496,N_11020,N_10120);
or U14497 (N_14497,N_11175,N_10642);
and U14498 (N_14498,N_9318,N_11276);
nor U14499 (N_14499,N_11227,N_10981);
xnor U14500 (N_14500,N_10712,N_10231);
nand U14501 (N_14501,N_9784,N_11563);
and U14502 (N_14502,N_9543,N_10000);
nand U14503 (N_14503,N_11962,N_10151);
and U14504 (N_14504,N_9360,N_11812);
nand U14505 (N_14505,N_9551,N_11630);
or U14506 (N_14506,N_9113,N_11552);
nand U14507 (N_14507,N_11823,N_11825);
xor U14508 (N_14508,N_9980,N_10600);
nand U14509 (N_14509,N_10370,N_10925);
nor U14510 (N_14510,N_10263,N_11249);
nor U14511 (N_14511,N_9446,N_10972);
nand U14512 (N_14512,N_9247,N_11996);
and U14513 (N_14513,N_10157,N_10077);
nor U14514 (N_14514,N_11669,N_11778);
nor U14515 (N_14515,N_10719,N_9663);
and U14516 (N_14516,N_9130,N_11769);
xnor U14517 (N_14517,N_10928,N_10778);
and U14518 (N_14518,N_11247,N_11119);
nand U14519 (N_14519,N_9583,N_11126);
nand U14520 (N_14520,N_10452,N_11352);
and U14521 (N_14521,N_9912,N_10815);
nor U14522 (N_14522,N_10005,N_9161);
nand U14523 (N_14523,N_9523,N_10313);
nor U14524 (N_14524,N_9375,N_11659);
nand U14525 (N_14525,N_11250,N_9377);
xnor U14526 (N_14526,N_11853,N_9108);
and U14527 (N_14527,N_10556,N_9124);
nor U14528 (N_14528,N_9701,N_10986);
or U14529 (N_14529,N_9975,N_9115);
nand U14530 (N_14530,N_11314,N_9486);
nor U14531 (N_14531,N_10773,N_11343);
xor U14532 (N_14532,N_9934,N_11185);
and U14533 (N_14533,N_10995,N_11188);
nand U14534 (N_14534,N_9258,N_10978);
or U14535 (N_14535,N_9497,N_9005);
nor U14536 (N_14536,N_10126,N_10861);
or U14537 (N_14537,N_9426,N_9946);
nor U14538 (N_14538,N_9922,N_10540);
and U14539 (N_14539,N_9120,N_10242);
xnor U14540 (N_14540,N_9120,N_9394);
nor U14541 (N_14541,N_9579,N_10379);
and U14542 (N_14542,N_9331,N_9501);
nand U14543 (N_14543,N_9735,N_11084);
nand U14544 (N_14544,N_11406,N_11303);
nor U14545 (N_14545,N_10075,N_11041);
and U14546 (N_14546,N_10865,N_11255);
nor U14547 (N_14547,N_11122,N_11868);
and U14548 (N_14548,N_9470,N_10868);
and U14549 (N_14549,N_9448,N_11924);
nand U14550 (N_14550,N_10739,N_9393);
nor U14551 (N_14551,N_11065,N_11107);
or U14552 (N_14552,N_11465,N_9878);
or U14553 (N_14553,N_11410,N_10640);
nand U14554 (N_14554,N_11082,N_9887);
nor U14555 (N_14555,N_11279,N_11452);
nand U14556 (N_14556,N_10303,N_11787);
nor U14557 (N_14557,N_10621,N_9144);
and U14558 (N_14558,N_10843,N_10499);
or U14559 (N_14559,N_9066,N_11352);
nand U14560 (N_14560,N_9071,N_10461);
or U14561 (N_14561,N_10942,N_10932);
or U14562 (N_14562,N_11517,N_10361);
and U14563 (N_14563,N_11229,N_10068);
nand U14564 (N_14564,N_10538,N_10271);
and U14565 (N_14565,N_11021,N_11514);
or U14566 (N_14566,N_11327,N_11202);
or U14567 (N_14567,N_10999,N_11153);
nor U14568 (N_14568,N_10180,N_11547);
and U14569 (N_14569,N_11808,N_9012);
nand U14570 (N_14570,N_9478,N_10449);
nor U14571 (N_14571,N_10691,N_9754);
nand U14572 (N_14572,N_11954,N_9989);
nand U14573 (N_14573,N_10602,N_11655);
and U14574 (N_14574,N_9883,N_10083);
nor U14575 (N_14575,N_9603,N_9113);
nor U14576 (N_14576,N_11863,N_9225);
and U14577 (N_14577,N_9063,N_11597);
and U14578 (N_14578,N_9558,N_10381);
nand U14579 (N_14579,N_10762,N_9355);
or U14580 (N_14580,N_9538,N_11115);
and U14581 (N_14581,N_9953,N_10036);
nand U14582 (N_14582,N_10955,N_9669);
or U14583 (N_14583,N_9396,N_9371);
and U14584 (N_14584,N_10759,N_11377);
or U14585 (N_14585,N_10997,N_9426);
nand U14586 (N_14586,N_9548,N_10869);
nor U14587 (N_14587,N_11496,N_11197);
nor U14588 (N_14588,N_10179,N_11095);
nor U14589 (N_14589,N_11949,N_10324);
nor U14590 (N_14590,N_11206,N_9569);
and U14591 (N_14591,N_11947,N_10839);
or U14592 (N_14592,N_10909,N_11297);
or U14593 (N_14593,N_11772,N_9544);
or U14594 (N_14594,N_10439,N_9538);
nor U14595 (N_14595,N_11089,N_9788);
nor U14596 (N_14596,N_9783,N_10264);
nand U14597 (N_14597,N_11088,N_10967);
or U14598 (N_14598,N_10125,N_11347);
and U14599 (N_14599,N_9144,N_10517);
nor U14600 (N_14600,N_11722,N_9769);
or U14601 (N_14601,N_10149,N_9426);
nor U14602 (N_14602,N_11815,N_10327);
and U14603 (N_14603,N_9322,N_9398);
nor U14604 (N_14604,N_9224,N_9264);
nand U14605 (N_14605,N_10463,N_11883);
or U14606 (N_14606,N_10951,N_9511);
nor U14607 (N_14607,N_9685,N_11932);
or U14608 (N_14608,N_11837,N_10060);
and U14609 (N_14609,N_10160,N_11596);
nor U14610 (N_14610,N_9733,N_9796);
and U14611 (N_14611,N_10014,N_9568);
and U14612 (N_14612,N_10748,N_10863);
and U14613 (N_14613,N_10713,N_11079);
nor U14614 (N_14614,N_9014,N_10295);
and U14615 (N_14615,N_10337,N_9853);
or U14616 (N_14616,N_10670,N_10436);
or U14617 (N_14617,N_11079,N_9009);
and U14618 (N_14618,N_9950,N_10166);
nor U14619 (N_14619,N_10751,N_11733);
nor U14620 (N_14620,N_9464,N_11953);
or U14621 (N_14621,N_9587,N_10894);
or U14622 (N_14622,N_10588,N_11227);
nand U14623 (N_14623,N_9240,N_10597);
and U14624 (N_14624,N_10196,N_10218);
nand U14625 (N_14625,N_11642,N_10634);
nor U14626 (N_14626,N_11875,N_10468);
nand U14627 (N_14627,N_9653,N_9085);
nand U14628 (N_14628,N_10941,N_9185);
and U14629 (N_14629,N_9565,N_11260);
or U14630 (N_14630,N_11298,N_11003);
nand U14631 (N_14631,N_11506,N_9874);
or U14632 (N_14632,N_10324,N_10783);
nor U14633 (N_14633,N_10380,N_10436);
and U14634 (N_14634,N_11519,N_10476);
nand U14635 (N_14635,N_10255,N_11120);
and U14636 (N_14636,N_9541,N_9702);
or U14637 (N_14637,N_11376,N_9033);
nor U14638 (N_14638,N_9389,N_10109);
or U14639 (N_14639,N_10397,N_11092);
nand U14640 (N_14640,N_10563,N_11694);
nand U14641 (N_14641,N_11593,N_9879);
and U14642 (N_14642,N_10369,N_11013);
or U14643 (N_14643,N_9264,N_10593);
and U14644 (N_14644,N_11208,N_9803);
nor U14645 (N_14645,N_10986,N_9488);
nand U14646 (N_14646,N_11825,N_10502);
or U14647 (N_14647,N_9732,N_11465);
and U14648 (N_14648,N_9466,N_9685);
nand U14649 (N_14649,N_11593,N_10500);
and U14650 (N_14650,N_10453,N_10672);
nor U14651 (N_14651,N_9399,N_10103);
nor U14652 (N_14652,N_10827,N_9077);
or U14653 (N_14653,N_10963,N_9560);
nand U14654 (N_14654,N_10762,N_10879);
or U14655 (N_14655,N_11668,N_10125);
nand U14656 (N_14656,N_11030,N_10845);
nand U14657 (N_14657,N_9065,N_11144);
and U14658 (N_14658,N_10353,N_11274);
or U14659 (N_14659,N_11018,N_11155);
or U14660 (N_14660,N_9778,N_10270);
nand U14661 (N_14661,N_10728,N_10765);
nor U14662 (N_14662,N_11520,N_9618);
nor U14663 (N_14663,N_9922,N_9862);
nor U14664 (N_14664,N_10082,N_10148);
nand U14665 (N_14665,N_11802,N_11393);
or U14666 (N_14666,N_9799,N_10293);
xnor U14667 (N_14667,N_11102,N_11975);
or U14668 (N_14668,N_10646,N_9174);
nor U14669 (N_14669,N_10937,N_10146);
nor U14670 (N_14670,N_9645,N_11065);
nand U14671 (N_14671,N_9042,N_9697);
and U14672 (N_14672,N_11289,N_11531);
nor U14673 (N_14673,N_11408,N_10254);
and U14674 (N_14674,N_11222,N_10922);
or U14675 (N_14675,N_11422,N_10509);
and U14676 (N_14676,N_10270,N_11274);
nand U14677 (N_14677,N_11784,N_10893);
and U14678 (N_14678,N_11212,N_10734);
nand U14679 (N_14679,N_9493,N_11874);
or U14680 (N_14680,N_9398,N_10542);
or U14681 (N_14681,N_9421,N_9745);
nor U14682 (N_14682,N_9927,N_9413);
nor U14683 (N_14683,N_10700,N_9758);
or U14684 (N_14684,N_11759,N_11242);
nor U14685 (N_14685,N_10486,N_11769);
nand U14686 (N_14686,N_9616,N_10440);
nand U14687 (N_14687,N_9880,N_9157);
nand U14688 (N_14688,N_9459,N_9039);
nand U14689 (N_14689,N_10118,N_9941);
xnor U14690 (N_14690,N_10917,N_11850);
nor U14691 (N_14691,N_9473,N_11015);
nand U14692 (N_14692,N_11104,N_11832);
or U14693 (N_14693,N_9970,N_11351);
nand U14694 (N_14694,N_11901,N_11015);
nor U14695 (N_14695,N_11876,N_10268);
nand U14696 (N_14696,N_11414,N_10249);
nand U14697 (N_14697,N_9018,N_9587);
nor U14698 (N_14698,N_11713,N_11880);
and U14699 (N_14699,N_10123,N_10554);
and U14700 (N_14700,N_10917,N_11061);
and U14701 (N_14701,N_10467,N_10249);
and U14702 (N_14702,N_9606,N_11679);
nand U14703 (N_14703,N_9303,N_9767);
nand U14704 (N_14704,N_9676,N_9430);
or U14705 (N_14705,N_9331,N_11002);
nand U14706 (N_14706,N_9289,N_11206);
nand U14707 (N_14707,N_11832,N_10988);
or U14708 (N_14708,N_9900,N_10028);
and U14709 (N_14709,N_9086,N_9576);
and U14710 (N_14710,N_10645,N_11904);
nor U14711 (N_14711,N_11174,N_10401);
nand U14712 (N_14712,N_9100,N_9277);
and U14713 (N_14713,N_10495,N_11031);
nor U14714 (N_14714,N_10522,N_11611);
or U14715 (N_14715,N_11197,N_11165);
and U14716 (N_14716,N_10597,N_9982);
and U14717 (N_14717,N_11494,N_11572);
nor U14718 (N_14718,N_9091,N_10408);
or U14719 (N_14719,N_11251,N_11948);
or U14720 (N_14720,N_11244,N_11065);
nand U14721 (N_14721,N_9001,N_9082);
nand U14722 (N_14722,N_10490,N_9709);
nor U14723 (N_14723,N_9863,N_10186);
and U14724 (N_14724,N_10834,N_10568);
or U14725 (N_14725,N_11820,N_11915);
and U14726 (N_14726,N_10382,N_9532);
nand U14727 (N_14727,N_9039,N_11904);
nor U14728 (N_14728,N_9948,N_11731);
and U14729 (N_14729,N_10128,N_10377);
xnor U14730 (N_14730,N_9714,N_11092);
nand U14731 (N_14731,N_9396,N_9603);
nand U14732 (N_14732,N_9948,N_9827);
nor U14733 (N_14733,N_10586,N_11519);
nor U14734 (N_14734,N_9054,N_9043);
nand U14735 (N_14735,N_10467,N_10654);
nor U14736 (N_14736,N_10524,N_9382);
or U14737 (N_14737,N_10749,N_10696);
and U14738 (N_14738,N_10110,N_9964);
nand U14739 (N_14739,N_9949,N_10612);
nor U14740 (N_14740,N_10040,N_11801);
nand U14741 (N_14741,N_10720,N_10900);
nand U14742 (N_14742,N_9809,N_10713);
nand U14743 (N_14743,N_10739,N_10345);
or U14744 (N_14744,N_10247,N_11946);
and U14745 (N_14745,N_9671,N_10353);
or U14746 (N_14746,N_9022,N_11037);
or U14747 (N_14747,N_9170,N_10825);
nor U14748 (N_14748,N_9881,N_11326);
nand U14749 (N_14749,N_9737,N_10746);
nand U14750 (N_14750,N_10731,N_11063);
xor U14751 (N_14751,N_9382,N_10785);
and U14752 (N_14752,N_11032,N_9276);
or U14753 (N_14753,N_10071,N_11151);
or U14754 (N_14754,N_11211,N_10896);
or U14755 (N_14755,N_11388,N_9023);
nand U14756 (N_14756,N_9027,N_10983);
and U14757 (N_14757,N_9679,N_9351);
and U14758 (N_14758,N_11138,N_9481);
or U14759 (N_14759,N_10301,N_10328);
or U14760 (N_14760,N_10051,N_11851);
nor U14761 (N_14761,N_11169,N_10315);
nor U14762 (N_14762,N_10958,N_9708);
or U14763 (N_14763,N_9968,N_10512);
xor U14764 (N_14764,N_11833,N_9755);
nand U14765 (N_14765,N_11570,N_9524);
and U14766 (N_14766,N_10100,N_9706);
or U14767 (N_14767,N_9977,N_9089);
xor U14768 (N_14768,N_10774,N_9111);
nor U14769 (N_14769,N_10767,N_9931);
and U14770 (N_14770,N_9316,N_9445);
nand U14771 (N_14771,N_10799,N_11750);
and U14772 (N_14772,N_11136,N_9560);
or U14773 (N_14773,N_10085,N_11874);
and U14774 (N_14774,N_9243,N_10020);
or U14775 (N_14775,N_10945,N_10865);
xnor U14776 (N_14776,N_11497,N_11942);
nand U14777 (N_14777,N_9309,N_10718);
nor U14778 (N_14778,N_11519,N_10393);
nand U14779 (N_14779,N_9086,N_9195);
nand U14780 (N_14780,N_9992,N_11173);
nor U14781 (N_14781,N_11100,N_9664);
nand U14782 (N_14782,N_9641,N_9666);
or U14783 (N_14783,N_9861,N_10774);
nor U14784 (N_14784,N_11569,N_10413);
nor U14785 (N_14785,N_9543,N_10093);
or U14786 (N_14786,N_9745,N_9833);
and U14787 (N_14787,N_9441,N_9604);
and U14788 (N_14788,N_10628,N_9175);
nand U14789 (N_14789,N_11620,N_11197);
or U14790 (N_14790,N_10228,N_10382);
nor U14791 (N_14791,N_11926,N_10016);
nand U14792 (N_14792,N_10423,N_11822);
and U14793 (N_14793,N_9521,N_11865);
and U14794 (N_14794,N_10840,N_10557);
nand U14795 (N_14795,N_9423,N_10466);
and U14796 (N_14796,N_9430,N_11479);
nor U14797 (N_14797,N_11963,N_11793);
nand U14798 (N_14798,N_9782,N_9943);
and U14799 (N_14799,N_11477,N_9692);
nor U14800 (N_14800,N_11481,N_9688);
or U14801 (N_14801,N_10692,N_10151);
or U14802 (N_14802,N_10258,N_9209);
xnor U14803 (N_14803,N_10877,N_9750);
nor U14804 (N_14804,N_11770,N_11726);
and U14805 (N_14805,N_10117,N_11627);
and U14806 (N_14806,N_9757,N_11163);
nor U14807 (N_14807,N_9783,N_11959);
nor U14808 (N_14808,N_11513,N_10735);
nand U14809 (N_14809,N_9260,N_11429);
and U14810 (N_14810,N_10249,N_10635);
xnor U14811 (N_14811,N_9509,N_10051);
nand U14812 (N_14812,N_9310,N_11894);
nor U14813 (N_14813,N_11137,N_10654);
xor U14814 (N_14814,N_10785,N_10650);
or U14815 (N_14815,N_11048,N_11629);
nand U14816 (N_14816,N_10396,N_9096);
nor U14817 (N_14817,N_9934,N_9048);
and U14818 (N_14818,N_10091,N_11776);
and U14819 (N_14819,N_11638,N_10530);
nor U14820 (N_14820,N_9219,N_11883);
nand U14821 (N_14821,N_10100,N_11194);
nor U14822 (N_14822,N_10803,N_9810);
nand U14823 (N_14823,N_9375,N_10500);
nor U14824 (N_14824,N_9276,N_9263);
nand U14825 (N_14825,N_10897,N_10789);
or U14826 (N_14826,N_11181,N_10611);
xnor U14827 (N_14827,N_11342,N_10651);
and U14828 (N_14828,N_10871,N_10451);
nand U14829 (N_14829,N_11907,N_11338);
nor U14830 (N_14830,N_9417,N_9548);
and U14831 (N_14831,N_9811,N_10245);
nor U14832 (N_14832,N_11133,N_11602);
and U14833 (N_14833,N_11240,N_9325);
nor U14834 (N_14834,N_10021,N_11416);
or U14835 (N_14835,N_11211,N_9563);
and U14836 (N_14836,N_11340,N_10724);
xor U14837 (N_14837,N_11416,N_9436);
and U14838 (N_14838,N_10635,N_10983);
or U14839 (N_14839,N_9156,N_10569);
and U14840 (N_14840,N_9855,N_11083);
nor U14841 (N_14841,N_10681,N_11643);
or U14842 (N_14842,N_9351,N_10563);
nand U14843 (N_14843,N_10720,N_11125);
nand U14844 (N_14844,N_9883,N_11356);
and U14845 (N_14845,N_9479,N_9878);
nand U14846 (N_14846,N_11611,N_9881);
and U14847 (N_14847,N_9295,N_11339);
xnor U14848 (N_14848,N_10719,N_10094);
and U14849 (N_14849,N_11099,N_10432);
nor U14850 (N_14850,N_9732,N_11252);
and U14851 (N_14851,N_9392,N_11950);
nand U14852 (N_14852,N_10360,N_9702);
or U14853 (N_14853,N_9224,N_11633);
nand U14854 (N_14854,N_11801,N_10355);
nor U14855 (N_14855,N_9458,N_11333);
nor U14856 (N_14856,N_11984,N_9826);
nor U14857 (N_14857,N_10802,N_11765);
or U14858 (N_14858,N_11849,N_10512);
and U14859 (N_14859,N_9484,N_10818);
nand U14860 (N_14860,N_10682,N_10155);
and U14861 (N_14861,N_11598,N_9295);
or U14862 (N_14862,N_10106,N_10674);
or U14863 (N_14863,N_9443,N_10492);
nor U14864 (N_14864,N_9645,N_10822);
and U14865 (N_14865,N_9117,N_10996);
nand U14866 (N_14866,N_9985,N_9814);
nor U14867 (N_14867,N_9458,N_9400);
and U14868 (N_14868,N_10839,N_9650);
and U14869 (N_14869,N_11566,N_10121);
nor U14870 (N_14870,N_9461,N_10902);
nor U14871 (N_14871,N_11400,N_10233);
and U14872 (N_14872,N_9567,N_10425);
nand U14873 (N_14873,N_10131,N_9576);
nor U14874 (N_14874,N_9535,N_10820);
nand U14875 (N_14875,N_10583,N_11695);
and U14876 (N_14876,N_10234,N_10575);
or U14877 (N_14877,N_10746,N_9999);
nor U14878 (N_14878,N_11518,N_9319);
nor U14879 (N_14879,N_10211,N_9027);
or U14880 (N_14880,N_10735,N_10845);
nand U14881 (N_14881,N_10022,N_10893);
or U14882 (N_14882,N_9891,N_11903);
or U14883 (N_14883,N_10662,N_10125);
and U14884 (N_14884,N_11242,N_11705);
nand U14885 (N_14885,N_9577,N_11679);
or U14886 (N_14886,N_10589,N_9777);
nand U14887 (N_14887,N_10732,N_10091);
nor U14888 (N_14888,N_11249,N_10075);
nand U14889 (N_14889,N_11876,N_9865);
nor U14890 (N_14890,N_9680,N_9921);
and U14891 (N_14891,N_9819,N_10540);
nand U14892 (N_14892,N_9379,N_9366);
nor U14893 (N_14893,N_10775,N_11029);
nor U14894 (N_14894,N_11432,N_9877);
or U14895 (N_14895,N_11386,N_9930);
and U14896 (N_14896,N_10111,N_10439);
or U14897 (N_14897,N_10860,N_10821);
nand U14898 (N_14898,N_11084,N_11232);
nor U14899 (N_14899,N_9418,N_10409);
or U14900 (N_14900,N_11639,N_11199);
nand U14901 (N_14901,N_11779,N_10800);
or U14902 (N_14902,N_9477,N_11178);
nand U14903 (N_14903,N_11277,N_11170);
and U14904 (N_14904,N_9630,N_11229);
and U14905 (N_14905,N_9397,N_9539);
nand U14906 (N_14906,N_11647,N_9699);
or U14907 (N_14907,N_10096,N_11948);
nor U14908 (N_14908,N_10813,N_10109);
nor U14909 (N_14909,N_10314,N_10863);
nor U14910 (N_14910,N_11016,N_11558);
and U14911 (N_14911,N_10293,N_9281);
or U14912 (N_14912,N_11097,N_9080);
nand U14913 (N_14913,N_10914,N_10652);
nand U14914 (N_14914,N_10491,N_11845);
and U14915 (N_14915,N_10264,N_9886);
nand U14916 (N_14916,N_10672,N_10510);
nand U14917 (N_14917,N_9848,N_10018);
nor U14918 (N_14918,N_9209,N_9566);
nand U14919 (N_14919,N_11992,N_11715);
and U14920 (N_14920,N_9447,N_10988);
and U14921 (N_14921,N_9674,N_9442);
nand U14922 (N_14922,N_11623,N_10816);
nand U14923 (N_14923,N_11032,N_9931);
nor U14924 (N_14924,N_11502,N_9432);
nor U14925 (N_14925,N_10099,N_9054);
and U14926 (N_14926,N_11584,N_9263);
or U14927 (N_14927,N_10362,N_11347);
nand U14928 (N_14928,N_11457,N_11677);
nor U14929 (N_14929,N_11156,N_11654);
or U14930 (N_14930,N_9858,N_9673);
and U14931 (N_14931,N_11126,N_10717);
or U14932 (N_14932,N_9532,N_11466);
nand U14933 (N_14933,N_9949,N_9917);
and U14934 (N_14934,N_10392,N_11015);
or U14935 (N_14935,N_11595,N_11912);
and U14936 (N_14936,N_9520,N_10580);
and U14937 (N_14937,N_9746,N_9640);
or U14938 (N_14938,N_10685,N_10070);
nor U14939 (N_14939,N_10054,N_9450);
or U14940 (N_14940,N_11977,N_11483);
nor U14941 (N_14941,N_10383,N_10875);
nor U14942 (N_14942,N_9524,N_10899);
nand U14943 (N_14943,N_10903,N_11376);
and U14944 (N_14944,N_10584,N_10073);
nor U14945 (N_14945,N_9659,N_10237);
nor U14946 (N_14946,N_11040,N_10833);
and U14947 (N_14947,N_11417,N_9088);
and U14948 (N_14948,N_11862,N_10270);
xnor U14949 (N_14949,N_11943,N_10226);
and U14950 (N_14950,N_10045,N_10866);
and U14951 (N_14951,N_9719,N_11882);
or U14952 (N_14952,N_11772,N_9076);
nand U14953 (N_14953,N_10044,N_10097);
and U14954 (N_14954,N_9579,N_9777);
and U14955 (N_14955,N_9876,N_9266);
nand U14956 (N_14956,N_11788,N_10566);
or U14957 (N_14957,N_9022,N_11632);
nand U14958 (N_14958,N_9815,N_11321);
nor U14959 (N_14959,N_10381,N_9035);
nand U14960 (N_14960,N_10724,N_9565);
nand U14961 (N_14961,N_10435,N_10593);
or U14962 (N_14962,N_9891,N_10187);
and U14963 (N_14963,N_11549,N_11652);
nand U14964 (N_14964,N_9852,N_11452);
nand U14965 (N_14965,N_9769,N_11519);
and U14966 (N_14966,N_9876,N_10201);
nand U14967 (N_14967,N_10718,N_10462);
and U14968 (N_14968,N_11186,N_9497);
nand U14969 (N_14969,N_9349,N_10433);
nand U14970 (N_14970,N_10135,N_11537);
and U14971 (N_14971,N_11482,N_9077);
and U14972 (N_14972,N_9610,N_9142);
and U14973 (N_14973,N_10925,N_10590);
nand U14974 (N_14974,N_11349,N_9989);
nand U14975 (N_14975,N_10751,N_11667);
or U14976 (N_14976,N_10527,N_9088);
and U14977 (N_14977,N_11630,N_10200);
nand U14978 (N_14978,N_9417,N_9682);
nor U14979 (N_14979,N_9255,N_10451);
or U14980 (N_14980,N_10148,N_9839);
nor U14981 (N_14981,N_11218,N_9823);
nor U14982 (N_14982,N_11396,N_11534);
nor U14983 (N_14983,N_10014,N_11348);
or U14984 (N_14984,N_9322,N_9741);
nand U14985 (N_14985,N_11386,N_10822);
and U14986 (N_14986,N_10233,N_9733);
nor U14987 (N_14987,N_10421,N_11378);
nand U14988 (N_14988,N_9924,N_9393);
or U14989 (N_14989,N_9697,N_11397);
and U14990 (N_14990,N_10673,N_10914);
nand U14991 (N_14991,N_10294,N_11123);
or U14992 (N_14992,N_10560,N_11242);
and U14993 (N_14993,N_9356,N_11165);
nor U14994 (N_14994,N_9213,N_10362);
or U14995 (N_14995,N_10793,N_11889);
or U14996 (N_14996,N_11305,N_10318);
nor U14997 (N_14997,N_10440,N_11235);
or U14998 (N_14998,N_10987,N_9385);
nor U14999 (N_14999,N_10314,N_10201);
and UO_0 (O_0,N_12836,N_12136);
nor UO_1 (O_1,N_14964,N_13870);
nor UO_2 (O_2,N_12875,N_12396);
and UO_3 (O_3,N_12929,N_14644);
and UO_4 (O_4,N_13972,N_12627);
nor UO_5 (O_5,N_13196,N_14294);
nand UO_6 (O_6,N_12079,N_14550);
or UO_7 (O_7,N_14234,N_13046);
nor UO_8 (O_8,N_13065,N_12403);
nor UO_9 (O_9,N_12541,N_12475);
nor UO_10 (O_10,N_14021,N_12550);
nor UO_11 (O_11,N_14230,N_14766);
nor UO_12 (O_12,N_12869,N_12733);
and UO_13 (O_13,N_13515,N_14499);
nand UO_14 (O_14,N_14582,N_14354);
or UO_15 (O_15,N_12834,N_14761);
or UO_16 (O_16,N_13357,N_12582);
or UO_17 (O_17,N_13689,N_14738);
or UO_18 (O_18,N_14064,N_12747);
and UO_19 (O_19,N_14993,N_12116);
nand UO_20 (O_20,N_12957,N_13560);
nor UO_21 (O_21,N_12431,N_13545);
nor UO_22 (O_22,N_12255,N_13098);
xor UO_23 (O_23,N_12793,N_13340);
nor UO_24 (O_24,N_14327,N_14741);
or UO_25 (O_25,N_14673,N_13599);
and UO_26 (O_26,N_14503,N_12878);
nor UO_27 (O_27,N_12858,N_14840);
nand UO_28 (O_28,N_13147,N_13947);
or UO_29 (O_29,N_13057,N_13408);
nand UO_30 (O_30,N_13320,N_14219);
nor UO_31 (O_31,N_13937,N_14472);
nor UO_32 (O_32,N_12166,N_13486);
and UO_33 (O_33,N_12633,N_13701);
nand UO_34 (O_34,N_12820,N_13558);
or UO_35 (O_35,N_13038,N_12822);
nor UO_36 (O_36,N_13698,N_12441);
or UO_37 (O_37,N_12080,N_14085);
and UO_38 (O_38,N_12837,N_13479);
nor UO_39 (O_39,N_12902,N_12742);
nor UO_40 (O_40,N_14433,N_13799);
and UO_41 (O_41,N_12446,N_13395);
nand UO_42 (O_42,N_13430,N_14537);
nor UO_43 (O_43,N_14058,N_14783);
nor UO_44 (O_44,N_14057,N_14083);
or UO_45 (O_45,N_14259,N_14142);
or UO_46 (O_46,N_12385,N_14310);
nand UO_47 (O_47,N_13148,N_13686);
nand UO_48 (O_48,N_14596,N_13235);
and UO_49 (O_49,N_12104,N_13043);
and UO_50 (O_50,N_12915,N_14179);
or UO_51 (O_51,N_14031,N_13469);
or UO_52 (O_52,N_14937,N_14255);
nor UO_53 (O_53,N_12603,N_14697);
and UO_54 (O_54,N_12358,N_12783);
and UO_55 (O_55,N_12273,N_12043);
nand UO_56 (O_56,N_12295,N_14606);
and UO_57 (O_57,N_14584,N_13151);
and UO_58 (O_58,N_12500,N_14041);
and UO_59 (O_59,N_13164,N_12367);
xor UO_60 (O_60,N_13574,N_13814);
nand UO_61 (O_61,N_13021,N_14396);
nor UO_62 (O_62,N_14850,N_14658);
nand UO_63 (O_63,N_12901,N_13627);
and UO_64 (O_64,N_12111,N_14857);
nand UO_65 (O_65,N_13391,N_12590);
nor UO_66 (O_66,N_13883,N_13623);
nor UO_67 (O_67,N_14579,N_12652);
or UO_68 (O_68,N_13210,N_12845);
or UO_69 (O_69,N_14136,N_14954);
and UO_70 (O_70,N_14634,N_13743);
or UO_71 (O_71,N_14067,N_14316);
nor UO_72 (O_72,N_13637,N_14710);
nand UO_73 (O_73,N_13154,N_12331);
and UO_74 (O_74,N_12968,N_12135);
or UO_75 (O_75,N_12730,N_12756);
nor UO_76 (O_76,N_14305,N_14613);
or UO_77 (O_77,N_13314,N_12674);
and UO_78 (O_78,N_13795,N_12320);
nor UO_79 (O_79,N_12490,N_14553);
and UO_80 (O_80,N_14301,N_13872);
and UO_81 (O_81,N_14029,N_13393);
nand UO_82 (O_82,N_13311,N_13174);
or UO_83 (O_83,N_13012,N_14888);
nand UO_84 (O_84,N_13004,N_12433);
nor UO_85 (O_85,N_14967,N_13081);
nor UO_86 (O_86,N_12705,N_14286);
xor UO_87 (O_87,N_14638,N_12530);
or UO_88 (O_88,N_12734,N_14557);
or UO_89 (O_89,N_13646,N_13326);
nand UO_90 (O_90,N_14307,N_14914);
or UO_91 (O_91,N_14285,N_14877);
and UO_92 (O_92,N_13626,N_13252);
nor UO_93 (O_93,N_12567,N_13504);
nand UO_94 (O_94,N_13944,N_14966);
or UO_95 (O_95,N_14635,N_14719);
nor UO_96 (O_96,N_12791,N_13280);
nand UO_97 (O_97,N_12059,N_14180);
nand UO_98 (O_98,N_12168,N_13173);
or UO_99 (O_99,N_12860,N_12555);
nand UO_100 (O_100,N_14818,N_13633);
xor UO_101 (O_101,N_12425,N_14916);
nand UO_102 (O_102,N_14284,N_13533);
or UO_103 (O_103,N_14560,N_12174);
nand UO_104 (O_104,N_12948,N_13699);
nand UO_105 (O_105,N_12937,N_12106);
nor UO_106 (O_106,N_13918,N_14545);
and UO_107 (O_107,N_14485,N_13309);
nor UO_108 (O_108,N_13386,N_14032);
and UO_109 (O_109,N_14432,N_13593);
or UO_110 (O_110,N_12527,N_12127);
and UO_111 (O_111,N_14716,N_12888);
and UO_112 (O_112,N_14100,N_13956);
nor UO_113 (O_113,N_14073,N_14607);
or UO_114 (O_114,N_13133,N_12017);
nor UO_115 (O_115,N_12788,N_12177);
nor UO_116 (O_116,N_12884,N_14043);
nand UO_117 (O_117,N_13206,N_13374);
nand UO_118 (O_118,N_12741,N_14858);
or UO_119 (O_119,N_12246,N_13092);
nand UO_120 (O_120,N_13788,N_14325);
and UO_121 (O_121,N_14124,N_14308);
nor UO_122 (O_122,N_13645,N_14754);
and UO_123 (O_123,N_14657,N_12140);
and UO_124 (O_124,N_14614,N_14098);
and UO_125 (O_125,N_13505,N_14177);
nand UO_126 (O_126,N_13201,N_13267);
nand UO_127 (O_127,N_12903,N_14455);
or UO_128 (O_128,N_12006,N_12839);
and UO_129 (O_129,N_14563,N_13261);
or UO_130 (O_130,N_12090,N_14737);
or UO_131 (O_131,N_13105,N_12890);
or UO_132 (O_132,N_12546,N_12608);
nand UO_133 (O_133,N_13705,N_14496);
and UO_134 (O_134,N_14681,N_14702);
and UO_135 (O_135,N_12397,N_14734);
nor UO_136 (O_136,N_14399,N_13327);
nand UO_137 (O_137,N_12443,N_12923);
nand UO_138 (O_138,N_13367,N_12525);
nand UO_139 (O_139,N_14045,N_13602);
nor UO_140 (O_140,N_12574,N_13632);
nand UO_141 (O_141,N_14805,N_14933);
and UO_142 (O_142,N_12028,N_13496);
nor UO_143 (O_143,N_12581,N_12970);
nor UO_144 (O_144,N_14290,N_13217);
nand UO_145 (O_145,N_12014,N_12969);
nor UO_146 (O_146,N_14689,N_14152);
and UO_147 (O_147,N_12719,N_14210);
or UO_148 (O_148,N_12812,N_13498);
nor UO_149 (O_149,N_13338,N_14254);
nand UO_150 (O_150,N_14072,N_14438);
nand UO_151 (O_151,N_12231,N_12900);
or UO_152 (O_152,N_12941,N_13375);
or UO_153 (O_153,N_13616,N_13955);
nor UO_154 (O_154,N_14413,N_14151);
nor UO_155 (O_155,N_14982,N_12328);
and UO_156 (O_156,N_12815,N_14165);
nor UO_157 (O_157,N_14450,N_12348);
or UO_158 (O_158,N_14642,N_14027);
nor UO_159 (O_159,N_13824,N_14975);
and UO_160 (O_160,N_13125,N_14283);
and UO_161 (O_161,N_14037,N_13119);
nor UO_162 (O_162,N_13005,N_14922);
nor UO_163 (O_163,N_12847,N_13380);
nor UO_164 (O_164,N_14726,N_12195);
nor UO_165 (O_165,N_14971,N_14852);
or UO_166 (O_166,N_14267,N_14470);
nor UO_167 (O_167,N_13313,N_12067);
nand UO_168 (O_168,N_12473,N_12298);
nor UO_169 (O_169,N_14686,N_12657);
and UO_170 (O_170,N_13047,N_12818);
nor UO_171 (O_171,N_13040,N_13575);
nor UO_172 (O_172,N_13432,N_14848);
and UO_173 (O_173,N_14279,N_13774);
and UO_174 (O_174,N_12047,N_13964);
and UO_175 (O_175,N_13262,N_12735);
and UO_176 (O_176,N_14289,N_14728);
xnor UO_177 (O_177,N_12726,N_12096);
nand UO_178 (O_178,N_13145,N_14081);
nand UO_179 (O_179,N_12487,N_14640);
and UO_180 (O_180,N_13833,N_13707);
and UO_181 (O_181,N_12885,N_12798);
nor UO_182 (O_182,N_14256,N_12459);
nor UO_183 (O_183,N_14419,N_14976);
or UO_184 (O_184,N_14712,N_14587);
nor UO_185 (O_185,N_12631,N_13511);
nor UO_186 (O_186,N_14422,N_12270);
nor UO_187 (O_187,N_14175,N_12628);
or UO_188 (O_188,N_12737,N_14725);
xnor UO_189 (O_189,N_13735,N_13979);
or UO_190 (O_190,N_13869,N_13329);
nor UO_191 (O_191,N_12542,N_12517);
nand UO_192 (O_192,N_12873,N_14655);
nand UO_193 (O_193,N_14739,N_13926);
or UO_194 (O_194,N_12887,N_12029);
nor UO_195 (O_195,N_14304,N_12290);
nor UO_196 (O_196,N_13132,N_13683);
or UO_197 (O_197,N_13700,N_12368);
nand UO_198 (O_198,N_14816,N_12215);
nand UO_199 (O_199,N_12663,N_13237);
nand UO_200 (O_200,N_13389,N_13304);
or UO_201 (O_201,N_12825,N_14841);
and UO_202 (O_202,N_13346,N_12986);
and UO_203 (O_203,N_13225,N_12691);
nor UO_204 (O_204,N_14363,N_14102);
nor UO_205 (O_205,N_12149,N_13130);
nand UO_206 (O_206,N_14787,N_14352);
and UO_207 (O_207,N_12131,N_14174);
and UO_208 (O_208,N_14919,N_12019);
or UO_209 (O_209,N_13172,N_12641);
and UO_210 (O_210,N_13243,N_13382);
and UO_211 (O_211,N_13620,N_13288);
or UO_212 (O_212,N_14262,N_14694);
and UO_213 (O_213,N_12399,N_13428);
or UO_214 (O_214,N_13333,N_13856);
or UO_215 (O_215,N_14763,N_14544);
and UO_216 (O_216,N_14534,N_14660);
or UO_217 (O_217,N_13268,N_14382);
nand UO_218 (O_218,N_13975,N_13527);
and UO_219 (O_219,N_14000,N_13846);
and UO_220 (O_220,N_14384,N_14389);
nor UO_221 (O_221,N_12237,N_14520);
and UO_222 (O_222,N_12982,N_12926);
nor UO_223 (O_223,N_13512,N_12304);
or UO_224 (O_224,N_12416,N_14931);
and UO_225 (O_225,N_13205,N_12949);
nand UO_226 (O_226,N_12418,N_14208);
or UO_227 (O_227,N_13485,N_12714);
nor UO_228 (O_228,N_14135,N_12088);
or UO_229 (O_229,N_14198,N_14344);
and UO_230 (O_230,N_14099,N_14762);
nand UO_231 (O_231,N_13231,N_14918);
and UO_232 (O_232,N_14893,N_14809);
and UO_233 (O_233,N_12240,N_13638);
nor UO_234 (O_234,N_14406,N_12553);
nand UO_235 (O_235,N_12132,N_13952);
or UO_236 (O_236,N_14025,N_13019);
nor UO_237 (O_237,N_12423,N_12649);
and UO_238 (O_238,N_14828,N_13783);
nand UO_239 (O_239,N_12789,N_14778);
or UO_240 (O_240,N_14276,N_13358);
and UO_241 (O_241,N_14690,N_14409);
nand UO_242 (O_242,N_13807,N_14672);
nor UO_243 (O_243,N_14353,N_14249);
or UO_244 (O_244,N_14968,N_14610);
or UO_245 (O_245,N_12024,N_12376);
nor UO_246 (O_246,N_14329,N_12849);
and UO_247 (O_247,N_14890,N_14070);
and UO_248 (O_248,N_13448,N_13353);
or UO_249 (O_249,N_13661,N_14404);
and UO_250 (O_250,N_13658,N_12424);
xor UO_251 (O_251,N_12402,N_12523);
and UO_252 (O_252,N_12703,N_12575);
nor UO_253 (O_253,N_12062,N_14700);
nor UO_254 (O_254,N_12752,N_12061);
nor UO_255 (O_255,N_13143,N_14357);
or UO_256 (O_256,N_12597,N_14956);
and UO_257 (O_257,N_12053,N_13998);
xor UO_258 (O_258,N_14882,N_14132);
or UO_259 (O_259,N_12563,N_12154);
and UO_260 (O_260,N_12465,N_12564);
and UO_261 (O_261,N_13166,N_14653);
and UO_262 (O_262,N_14282,N_13837);
or UO_263 (O_263,N_14911,N_13880);
or UO_264 (O_264,N_14771,N_12738);
and UO_265 (O_265,N_14999,N_12119);
or UO_266 (O_266,N_12928,N_14471);
or UO_267 (O_267,N_14648,N_13829);
nor UO_268 (O_268,N_14552,N_14748);
or UO_269 (O_269,N_12232,N_12813);
and UO_270 (O_270,N_13903,N_14693);
nor UO_271 (O_271,N_13923,N_13414);
and UO_272 (O_272,N_14402,N_14424);
nor UO_273 (O_273,N_14541,N_12374);
or UO_274 (O_274,N_14351,N_14312);
nand UO_275 (O_275,N_13887,N_13761);
nor UO_276 (O_276,N_13269,N_14337);
nand UO_277 (O_277,N_14793,N_14113);
or UO_278 (O_278,N_14239,N_12327);
and UO_279 (O_279,N_12591,N_13376);
or UO_280 (O_280,N_14313,N_12005);
nor UO_281 (O_281,N_12770,N_13223);
nor UO_282 (O_282,N_13874,N_14757);
or UO_283 (O_283,N_14426,N_14167);
or UO_284 (O_284,N_13844,N_14695);
nand UO_285 (O_285,N_12921,N_13577);
and UO_286 (O_286,N_14183,N_12409);
or UO_287 (O_287,N_14874,N_12211);
nor UO_288 (O_288,N_13266,N_13753);
or UO_289 (O_289,N_14133,N_12623);
and UO_290 (O_290,N_14631,N_13347);
or UO_291 (O_291,N_13877,N_14838);
nor UO_292 (O_292,N_13471,N_14707);
and UO_293 (O_293,N_12700,N_14985);
and UO_294 (O_294,N_13191,N_13949);
and UO_295 (O_295,N_12513,N_13286);
nor UO_296 (O_296,N_13895,N_13715);
nand UO_297 (O_297,N_12435,N_12023);
nand UO_298 (O_298,N_13051,N_13158);
xnor UO_299 (O_299,N_13866,N_12158);
nor UO_300 (O_300,N_12412,N_14457);
and UO_301 (O_301,N_13335,N_12334);
nor UO_302 (O_302,N_14833,N_12238);
or UO_303 (O_303,N_13033,N_14140);
and UO_304 (O_304,N_12044,N_13981);
or UO_305 (O_305,N_13028,N_12613);
nand UO_306 (O_306,N_12463,N_14190);
or UO_307 (O_307,N_12662,N_13483);
or UO_308 (O_308,N_14427,N_12365);
nor UO_309 (O_309,N_12528,N_13230);
or UO_310 (O_310,N_14575,N_12538);
nor UO_311 (O_311,N_13199,N_13216);
nor UO_312 (O_312,N_12081,N_13908);
nor UO_313 (O_313,N_14188,N_12020);
and UO_314 (O_314,N_13458,N_12919);
and UO_315 (O_315,N_13214,N_13094);
nor UO_316 (O_316,N_14498,N_12583);
or UO_317 (O_317,N_13589,N_12366);
nor UO_318 (O_318,N_14277,N_13138);
and UO_319 (O_319,N_12739,N_13780);
nor UO_320 (O_320,N_14274,N_13111);
nand UO_321 (O_321,N_14191,N_14950);
nand UO_322 (O_322,N_14374,N_12655);
or UO_323 (O_323,N_13211,N_13927);
nand UO_324 (O_324,N_14220,N_14578);
and UO_325 (O_325,N_14163,N_14388);
xor UO_326 (O_326,N_14530,N_12980);
or UO_327 (O_327,N_13372,N_13531);
and UO_328 (O_328,N_14297,N_13178);
and UO_329 (O_329,N_12850,N_14901);
and UO_330 (O_330,N_12973,N_13818);
and UO_331 (O_331,N_14633,N_13023);
nor UO_332 (O_332,N_14595,N_13849);
xnor UO_333 (O_333,N_12797,N_14233);
nand UO_334 (O_334,N_12569,N_14094);
nor UO_335 (O_335,N_12417,N_14097);
nor UO_336 (O_336,N_12579,N_13924);
or UO_337 (O_337,N_13289,N_13350);
and UO_338 (O_338,N_12436,N_14115);
or UO_339 (O_339,N_12727,N_14405);
nand UO_340 (O_340,N_12592,N_12796);
xor UO_341 (O_341,N_14831,N_12274);
nand UO_342 (O_342,N_12689,N_14643);
or UO_343 (O_343,N_12160,N_13366);
and UO_344 (O_344,N_14080,N_12557);
or UO_345 (O_345,N_13757,N_14125);
or UO_346 (O_346,N_13000,N_12344);
and UO_347 (O_347,N_12282,N_13624);
nand UO_348 (O_348,N_14126,N_12066);
nand UO_349 (O_349,N_14941,N_14367);
or UO_350 (O_350,N_13508,N_12675);
nor UO_351 (O_351,N_13711,N_12315);
nor UO_352 (O_352,N_12978,N_12883);
or UO_353 (O_353,N_12207,N_13187);
nand UO_354 (O_354,N_12805,N_14536);
or UO_355 (O_355,N_12469,N_12307);
nand UO_356 (O_356,N_14765,N_13596);
nand UO_357 (O_357,N_13087,N_13169);
or UO_358 (O_358,N_12682,N_14205);
nor UO_359 (O_359,N_13122,N_13284);
and UO_360 (O_360,N_13819,N_14444);
and UO_361 (O_361,N_14265,N_12408);
nor UO_362 (O_362,N_13739,N_13054);
and UO_363 (O_363,N_13969,N_13960);
nor UO_364 (O_364,N_12755,N_12971);
and UO_365 (O_365,N_14299,N_14987);
or UO_366 (O_366,N_12352,N_14245);
and UO_367 (O_367,N_14446,N_13195);
nor UO_368 (O_368,N_13867,N_12084);
nor UO_369 (O_369,N_13826,N_14755);
nor UO_370 (O_370,N_13062,N_13406);
or UO_371 (O_371,N_14360,N_13635);
and UO_372 (O_372,N_12256,N_14480);
and UO_373 (O_373,N_12802,N_14416);
and UO_374 (O_374,N_13665,N_12519);
nor UO_375 (O_375,N_13968,N_12203);
nor UO_376 (O_376,N_14410,N_14323);
xnor UO_377 (O_377,N_13907,N_13929);
and UO_378 (O_378,N_13659,N_14318);
xnor UO_379 (O_379,N_14768,N_13948);
or UO_380 (O_380,N_12959,N_14244);
nor UO_381 (O_381,N_13896,N_12323);
nand UO_382 (O_382,N_13352,N_13666);
nor UO_383 (O_383,N_14714,N_13011);
and UO_384 (O_384,N_12013,N_12117);
nor UO_385 (O_385,N_14088,N_13032);
and UO_386 (O_386,N_14970,N_13830);
or UO_387 (O_387,N_13800,N_12434);
nor UO_388 (O_388,N_13290,N_12831);
or UO_389 (O_389,N_12483,N_13928);
and UO_390 (O_390,N_14129,N_12065);
and UO_391 (O_391,N_13524,N_13369);
nor UO_392 (O_392,N_12379,N_14696);
or UO_393 (O_393,N_12317,N_14128);
nor UO_394 (O_394,N_13002,N_14494);
or UO_395 (O_395,N_13114,N_12015);
and UO_396 (O_396,N_14887,N_12985);
nand UO_397 (O_397,N_13559,N_13962);
or UO_398 (O_398,N_13283,N_14039);
and UO_399 (O_399,N_14692,N_14292);
nand UO_400 (O_400,N_13464,N_12782);
or UO_401 (O_401,N_13112,N_14232);
nor UO_402 (O_402,N_13653,N_14053);
and UO_403 (O_403,N_13355,N_14623);
and UO_404 (O_404,N_14618,N_13936);
or UO_405 (O_405,N_12731,N_13052);
nand UO_406 (O_406,N_13823,N_14456);
nand UO_407 (O_407,N_13398,N_12272);
and UO_408 (O_408,N_12279,N_14273);
and UO_409 (O_409,N_12181,N_14028);
nor UO_410 (O_410,N_12234,N_12069);
and UO_411 (O_411,N_14980,N_12872);
nand UO_412 (O_412,N_12100,N_12035);
or UO_413 (O_413,N_13091,N_14153);
and UO_414 (O_414,N_12002,N_12909);
or UO_415 (O_415,N_14065,N_12593);
or UO_416 (O_416,N_12164,N_12746);
or UO_417 (O_417,N_13601,N_13249);
and UO_418 (O_418,N_12637,N_13457);
or UO_419 (O_419,N_13538,N_13449);
and UO_420 (O_420,N_12251,N_14863);
and UO_421 (O_421,N_14724,N_14150);
and UO_422 (O_422,N_12640,N_14935);
nor UO_423 (O_423,N_13368,N_13299);
nor UO_424 (O_424,N_12498,N_13827);
nor UO_425 (O_425,N_13769,N_14050);
and UO_426 (O_426,N_12497,N_13770);
and UO_427 (O_427,N_14845,N_14439);
nor UO_428 (O_428,N_12007,N_12499);
nor UO_429 (O_429,N_13762,N_12151);
nand UO_430 (O_430,N_12075,N_13958);
nand UO_431 (O_431,N_12091,N_13241);
nor UO_432 (O_432,N_14797,N_12855);
nor UO_433 (O_433,N_12192,N_13344);
and UO_434 (O_434,N_12810,N_12912);
or UO_435 (O_435,N_14779,N_14012);
nor UO_436 (O_436,N_14952,N_14669);
or UO_437 (O_437,N_14780,N_14280);
or UO_438 (O_438,N_14972,N_12233);
nor UO_439 (O_439,N_13781,N_13418);
and UO_440 (O_440,N_14068,N_14341);
nor UO_441 (O_441,N_12283,N_12225);
and UO_442 (O_442,N_12994,N_13050);
and UO_443 (O_443,N_12389,N_14711);
nor UO_444 (O_444,N_14158,N_13131);
and UO_445 (O_445,N_14293,N_12202);
nor UO_446 (O_446,N_12764,N_12997);
xnor UO_447 (O_447,N_13808,N_13640);
nor UO_448 (O_448,N_12388,N_14300);
nand UO_449 (O_449,N_12670,N_12205);
or UO_450 (O_450,N_12276,N_12321);
or UO_451 (O_451,N_14359,N_14176);
and UO_452 (O_452,N_12524,N_13815);
and UO_453 (O_453,N_14875,N_12312);
or UO_454 (O_454,N_12182,N_13541);
and UO_455 (O_455,N_14609,N_13069);
and UO_456 (O_456,N_12543,N_13010);
nand UO_457 (O_457,N_12570,N_13411);
or UO_458 (O_458,N_12128,N_12607);
nand UO_459 (O_459,N_12963,N_12578);
nor UO_460 (O_460,N_14769,N_14910);
and UO_461 (O_461,N_13614,N_14311);
or UO_462 (O_462,N_14788,N_13322);
or UO_463 (O_463,N_14646,N_14706);
nor UO_464 (O_464,N_14790,N_14899);
or UO_465 (O_465,N_14731,N_14047);
nand UO_466 (O_466,N_13410,N_14435);
or UO_467 (O_467,N_14322,N_12484);
nor UO_468 (O_468,N_13873,N_14548);
nand UO_469 (O_469,N_13443,N_12584);
nand UO_470 (O_470,N_12865,N_13097);
nor UO_471 (O_471,N_12573,N_13994);
or UO_472 (O_472,N_12058,N_12843);
and UO_473 (O_473,N_12595,N_12363);
nand UO_474 (O_474,N_13441,N_14851);
nand UO_475 (O_475,N_14730,N_14004);
and UO_476 (O_476,N_13782,N_12511);
nor UO_477 (O_477,N_12426,N_12462);
or UO_478 (O_478,N_13759,N_14026);
or UO_479 (O_479,N_12341,N_14758);
or UO_480 (O_480,N_13549,N_13392);
or UO_481 (O_481,N_12615,N_13473);
nand UO_482 (O_482,N_14022,N_12085);
nor UO_483 (O_483,N_14760,N_13006);
or UO_484 (O_484,N_14934,N_14248);
nor UO_485 (O_485,N_12620,N_13951);
and UO_486 (O_486,N_12410,N_13692);
and UO_487 (O_487,N_14824,N_14889);
or UO_488 (O_488,N_13622,N_14001);
and UO_489 (O_489,N_14222,N_14194);
nor UO_490 (O_490,N_13048,N_14112);
and UO_491 (O_491,N_14509,N_13484);
nor UO_492 (O_492,N_12210,N_14871);
nand UO_493 (O_493,N_13186,N_13228);
or UO_494 (O_494,N_13536,N_14465);
nand UO_495 (O_495,N_14171,N_13470);
nor UO_496 (O_496,N_14143,N_14017);
nor UO_497 (O_497,N_14429,N_12961);
xor UO_498 (O_498,N_12302,N_13920);
or UO_499 (O_499,N_12522,N_13842);
nand UO_500 (O_500,N_14597,N_14782);
nand UO_501 (O_501,N_14802,N_12713);
nor UO_502 (O_502,N_13922,N_13631);
and UO_503 (O_503,N_14879,N_12046);
nor UO_504 (O_504,N_12297,N_12057);
nand UO_505 (O_505,N_13584,N_12618);
or UO_506 (O_506,N_14084,N_12337);
nand UO_507 (O_507,N_12976,N_13984);
nand UO_508 (O_508,N_12999,N_13976);
or UO_509 (O_509,N_14843,N_12535);
nor UO_510 (O_510,N_13478,N_13185);
nand UO_511 (O_511,N_12897,N_14856);
nor UO_512 (O_512,N_14598,N_13985);
and UO_513 (O_513,N_12082,N_14974);
nor UO_514 (O_514,N_14504,N_13255);
nor UO_515 (O_515,N_12137,N_14870);
nand UO_516 (O_516,N_14988,N_13259);
or UO_517 (O_517,N_12089,N_14679);
or UO_518 (O_518,N_12588,N_13194);
nand UO_519 (O_519,N_13360,N_13477);
nand UO_520 (O_520,N_14555,N_14767);
nor UO_521 (O_521,N_14071,N_14990);
nand UO_522 (O_522,N_14258,N_13089);
or UO_523 (O_523,N_13696,N_12656);
and UO_524 (O_524,N_14253,N_13784);
xor UO_525 (O_525,N_12074,N_13404);
nand UO_526 (O_526,N_12134,N_12179);
nand UO_527 (O_527,N_12281,N_13466);
or UO_528 (O_528,N_12454,N_14269);
or UO_529 (O_529,N_13727,N_13897);
nor UO_530 (O_530,N_13650,N_14287);
nand UO_531 (O_531,N_12621,N_12152);
nor UO_532 (O_532,N_12718,N_12247);
nand UO_533 (O_533,N_13563,N_14491);
and UO_534 (O_534,N_13945,N_13450);
or UO_535 (O_535,N_12988,N_12153);
nor UO_536 (O_536,N_12816,N_13697);
nor UO_537 (O_537,N_13383,N_12646);
and UO_538 (O_538,N_12068,N_14298);
nand UO_539 (O_539,N_13888,N_12003);
nand UO_540 (O_540,N_13071,N_12930);
nor UO_541 (O_541,N_13644,N_13433);
nand UO_542 (O_542,N_14948,N_12293);
nand UO_543 (O_543,N_12060,N_14807);
xnor UO_544 (O_544,N_13176,N_12138);
or UO_545 (O_545,N_14009,N_13664);
nand UO_546 (O_546,N_13649,N_13370);
nand UO_547 (O_547,N_12708,N_13642);
nor UO_548 (O_548,N_14773,N_14583);
and UO_549 (O_549,N_14146,N_13475);
and UO_550 (O_550,N_13207,N_12639);
and UO_551 (O_551,N_12846,N_13103);
nor UO_552 (O_552,N_13305,N_12678);
nand UO_553 (O_553,N_12226,N_13371);
and UO_554 (O_554,N_13323,N_12905);
or UO_555 (O_555,N_13253,N_13966);
and UO_556 (O_556,N_12697,N_14223);
nand UO_557 (O_557,N_14377,N_13177);
nor UO_558 (O_558,N_12228,N_13902);
or UO_559 (O_559,N_12840,N_14199);
nor UO_560 (O_560,N_13617,N_14362);
nand UO_561 (O_561,N_12979,N_12223);
nand UO_562 (O_562,N_12776,N_12311);
or UO_563 (O_563,N_14998,N_12357);
or UO_564 (O_564,N_14086,N_14184);
and UO_565 (O_565,N_12904,N_14202);
nand UO_566 (O_566,N_12178,N_14319);
nor UO_567 (O_567,N_14625,N_14204);
and UO_568 (O_568,N_12668,N_14139);
nor UO_569 (O_569,N_13362,N_13108);
nor UO_570 (O_570,N_14173,N_12432);
nor UO_571 (O_571,N_12732,N_13020);
xnor UO_572 (O_572,N_12684,N_12894);
nor UO_573 (O_573,N_12105,N_12685);
nand UO_574 (O_574,N_13342,N_12457);
nand UO_575 (O_575,N_14896,N_13317);
nand UO_576 (O_576,N_12638,N_13193);
or UO_577 (O_577,N_13116,N_14735);
or UO_578 (O_578,N_13212,N_14869);
and UO_579 (O_579,N_14109,N_12173);
or UO_580 (O_580,N_12495,N_14428);
and UO_581 (O_581,N_14529,N_13572);
nor UO_582 (O_582,N_12141,N_13239);
nor UO_583 (O_583,N_14532,N_13643);
nor UO_584 (O_584,N_12616,N_12956);
nand UO_585 (O_585,N_13655,N_12853);
nor UO_586 (O_586,N_13641,N_13754);
and UO_587 (O_587,N_13274,N_13017);
and UO_588 (O_588,N_13986,N_13034);
nor UO_589 (O_589,N_14556,N_12186);
nor UO_590 (O_590,N_14395,N_13328);
nor UO_591 (O_591,N_14543,N_13060);
nor UO_592 (O_592,N_13789,N_12572);
or UO_593 (O_593,N_14386,N_12466);
nand UO_594 (O_594,N_14926,N_12109);
and UO_595 (O_595,N_13009,N_12717);
nor UO_596 (O_596,N_14263,N_14822);
or UO_597 (O_597,N_13894,N_12350);
nor UO_598 (O_598,N_14819,N_14002);
or UO_599 (O_599,N_12220,N_13625);
or UO_600 (O_600,N_12129,N_13805);
nor UO_601 (O_601,N_14006,N_13090);
or UO_602 (O_602,N_12896,N_14718);
nor UO_603 (O_603,N_14630,N_13691);
nor UO_604 (O_604,N_14915,N_12165);
nor UO_605 (O_605,N_14034,N_12353);
nor UO_606 (O_606,N_12660,N_14929);
and UO_607 (O_607,N_14015,N_14364);
nor UO_608 (O_608,N_14701,N_13270);
nand UO_609 (O_609,N_14250,N_13082);
or UO_610 (O_610,N_13459,N_14581);
or UO_611 (O_611,N_12870,N_14798);
xnor UO_612 (O_612,N_13240,N_12139);
and UO_613 (O_613,N_13227,N_14592);
nor UO_614 (O_614,N_14913,N_12325);
or UO_615 (O_615,N_13709,N_13356);
nor UO_616 (O_616,N_12993,N_14355);
or UO_617 (O_617,N_13295,N_14243);
nand UO_618 (O_618,N_14574,N_12481);
or UO_619 (O_619,N_13750,N_12841);
nand UO_620 (O_620,N_13198,N_13794);
nor UO_621 (O_621,N_13919,N_14953);
nor UO_622 (O_622,N_12683,N_13868);
nor UO_623 (O_623,N_14649,N_13124);
or UO_624 (O_624,N_12038,N_13771);
nand UO_625 (O_625,N_13308,N_12042);
and UO_626 (O_626,N_13592,N_14775);
xnor UO_627 (O_627,N_12811,N_12720);
and UO_628 (O_628,N_14288,N_12171);
nand UO_629 (O_629,N_13016,N_13480);
nand UO_630 (O_630,N_14678,N_14441);
and UO_631 (O_631,N_12102,N_14401);
nor UO_632 (O_632,N_14569,N_12867);
nor UO_633 (O_633,N_12659,N_12666);
nor UO_634 (O_634,N_14492,N_14240);
or UO_635 (O_635,N_13115,N_14121);
and UO_636 (O_636,N_13570,N_13123);
or UO_637 (O_637,N_13053,N_12219);
or UO_638 (O_638,N_13067,N_13397);
and UO_639 (O_639,N_12144,N_13760);
nand UO_640 (O_640,N_14434,N_13461);
or UO_641 (O_641,N_12933,N_12771);
or UO_642 (O_642,N_13787,N_14523);
nand UO_643 (O_643,N_14593,N_12438);
nor UO_644 (O_644,N_13117,N_12785);
and UO_645 (O_645,N_13882,N_14049);
nand UO_646 (O_646,N_12194,N_12198);
nand UO_647 (O_647,N_14385,N_14616);
nor UO_648 (O_648,N_14366,N_13736);
nand UO_649 (O_649,N_12781,N_12030);
nand UO_650 (O_650,N_12474,N_12958);
and UO_651 (O_651,N_12953,N_14155);
or UO_652 (O_652,N_14209,N_14839);
nand UO_653 (O_653,N_12650,N_14235);
and UO_654 (O_654,N_13694,N_12318);
nor UO_655 (O_655,N_13066,N_14949);
nand UO_656 (O_656,N_14275,N_14347);
or UO_657 (O_657,N_13312,N_13492);
nor UO_658 (O_658,N_14117,N_12492);
or UO_659 (O_659,N_14580,N_12695);
and UO_660 (O_660,N_12995,N_13835);
or UO_661 (O_661,N_12387,N_13516);
and UO_662 (O_662,N_13146,N_14508);
or UO_663 (O_663,N_14781,N_14983);
or UO_664 (O_664,N_14376,N_13424);
nor UO_665 (O_665,N_14772,N_12838);
and UO_666 (O_666,N_12534,N_13113);
and UO_667 (O_667,N_14200,N_13991);
nand UO_668 (O_668,N_12120,N_13710);
or UO_669 (O_669,N_13950,N_14008);
and UO_670 (O_670,N_13501,N_13597);
and UO_671 (O_671,N_14484,N_13165);
and UO_672 (O_672,N_14189,N_14270);
nand UO_673 (O_673,N_13544,N_12163);
or UO_674 (O_674,N_14181,N_13493);
or UO_675 (O_675,N_14897,N_13238);
and UO_676 (O_676,N_12259,N_14342);
or UO_677 (O_677,N_13126,N_14114);
nor UO_678 (O_678,N_14221,N_12532);
nand UO_679 (O_679,N_12086,N_12442);
nand UO_680 (O_680,N_14519,N_12309);
nand UO_681 (O_681,N_12842,N_13722);
nand UO_682 (O_682,N_13245,N_13845);
and UO_683 (O_683,N_13224,N_12193);
nor UO_684 (O_684,N_14063,N_13965);
nor UO_685 (O_685,N_13881,N_13530);
nand UO_686 (O_686,N_14059,N_13300);
and UO_687 (O_687,N_12300,N_14829);
or UO_688 (O_688,N_14837,N_13183);
nand UO_689 (O_689,N_13550,N_14554);
nand UO_690 (O_690,N_13068,N_12817);
or UO_691 (O_691,N_13413,N_14803);
nor UO_692 (O_692,N_12794,N_14522);
nand UO_693 (O_693,N_14753,N_12429);
xnor UO_694 (O_694,N_14666,N_14608);
nor UO_695 (O_695,N_14601,N_12461);
nand UO_696 (O_696,N_13264,N_12748);
nor UO_697 (O_697,N_14637,N_13579);
and UO_698 (O_698,N_14390,N_14817);
nand UO_699 (O_699,N_13135,N_13244);
nor UO_700 (O_700,N_13909,N_13831);
nor UO_701 (O_701,N_14886,N_13378);
and UO_702 (O_702,N_13452,N_12694);
and UO_703 (O_703,N_13911,N_14420);
nor UO_704 (O_704,N_12394,N_14977);
nor UO_705 (O_705,N_12863,N_14381);
nand UO_706 (O_706,N_12634,N_14564);
and UO_707 (O_707,N_12258,N_12644);
nor UO_708 (O_708,N_14729,N_13776);
nor UO_709 (O_709,N_13741,N_14568);
nand UO_710 (O_710,N_13379,N_12072);
and UO_711 (O_711,N_13063,N_12033);
and UO_712 (O_712,N_12489,N_12911);
xnor UO_713 (O_713,N_12955,N_14717);
or UO_714 (O_714,N_13445,N_12510);
or UO_715 (O_715,N_13042,N_14500);
nor UO_716 (O_716,N_12221,N_14826);
nand UO_717 (O_717,N_14880,N_13134);
and UO_718 (O_718,N_14789,N_14495);
or UO_719 (O_719,N_13749,N_14501);
and UO_720 (O_720,N_13820,N_13772);
nand UO_721 (O_721,N_13656,N_13906);
and UO_722 (O_722,N_13403,N_14713);
nand UO_723 (O_723,N_13939,N_14627);
nand UO_724 (O_724,N_14013,N_13296);
nor UO_725 (O_725,N_13488,N_12183);
nor UO_726 (O_726,N_14349,N_12886);
nor UO_727 (O_727,N_14825,N_13619);
nor UO_728 (O_728,N_13732,N_13891);
nor UO_729 (O_729,N_12095,N_14612);
nor UO_730 (O_730,N_14884,N_12243);
and UO_731 (O_731,N_14218,N_13978);
xor UO_732 (O_732,N_14488,N_14699);
nor UO_733 (O_733,N_14827,N_13963);
and UO_734 (O_734,N_14978,N_13910);
nand UO_735 (O_735,N_13786,N_14516);
nand UO_736 (O_736,N_13843,N_12347);
or UO_737 (O_737,N_14836,N_12548);
nand UO_738 (O_738,N_13423,N_14195);
and UO_739 (O_739,N_12448,N_13556);
nor UO_740 (O_740,N_13070,N_12048);
or UO_741 (O_741,N_14481,N_14431);
nor UO_742 (O_742,N_12913,N_14108);
or UO_743 (O_743,N_12265,N_14561);
nor UO_744 (O_744,N_12686,N_13610);
and UO_745 (O_745,N_12502,N_12452);
nand UO_746 (O_746,N_14995,N_13365);
or UO_747 (O_747,N_13429,N_12340);
nor UO_748 (O_748,N_12121,N_13802);
or UO_749 (O_749,N_13218,N_14938);
nor UO_750 (O_750,N_12824,N_13077);
or UO_751 (O_751,N_14774,N_13307);
nor UO_752 (O_752,N_14003,N_12829);
nand UO_753 (O_753,N_13569,N_14475);
nand UO_754 (O_754,N_14296,N_12455);
and UO_755 (O_755,N_14445,N_14946);
nor UO_756 (O_756,N_12339,N_13106);
nor UO_757 (O_757,N_14844,N_12250);
nor UO_758 (O_758,N_13157,N_12935);
nor UO_759 (O_759,N_12244,N_14535);
nand UO_760 (O_760,N_14577,N_14559);
and UO_761 (O_761,N_13221,N_14489);
nor UO_762 (O_762,N_14105,N_14197);
nand UO_763 (O_763,N_12951,N_12882);
and UO_764 (O_764,N_13039,N_12333);
or UO_765 (O_765,N_12063,N_12806);
nand UO_766 (O_766,N_13405,N_12504);
and UO_767 (O_767,N_13578,N_13763);
or UO_768 (O_768,N_12440,N_13525);
and UO_769 (O_769,N_12010,N_14463);
nor UO_770 (O_770,N_14345,N_13297);
or UO_771 (O_771,N_13061,N_13861);
nand UO_772 (O_772,N_13684,N_14973);
and UO_773 (O_773,N_14663,N_14647);
and UO_774 (O_774,N_14749,N_14961);
nand UO_775 (O_775,N_12382,N_12464);
nor UO_776 (O_776,N_13534,N_13339);
and UO_777 (O_777,N_13745,N_14425);
nor UO_778 (O_778,N_13425,N_13607);
and UO_779 (O_779,N_13110,N_12145);
nand UO_780 (O_780,N_14078,N_13022);
or UO_781 (O_781,N_12778,N_12977);
or UO_782 (O_782,N_13639,N_13292);
or UO_783 (O_783,N_12594,N_13959);
and UO_784 (O_784,N_13407,N_12724);
xnor UO_785 (O_785,N_13319,N_13674);
or UO_786 (O_786,N_12908,N_13044);
xnor UO_787 (O_787,N_13100,N_13129);
nand UO_788 (O_788,N_12150,N_14268);
or UO_789 (O_789,N_13209,N_13208);
nand UO_790 (O_790,N_12406,N_13865);
or UO_791 (O_791,N_14392,N_12395);
and UO_792 (O_792,N_14830,N_14620);
or UO_793 (O_793,N_14014,N_14866);
and UO_794 (O_794,N_13351,N_12450);
nor UO_795 (O_795,N_14947,N_12142);
nor UO_796 (O_796,N_14722,N_12614);
or UO_797 (O_797,N_13420,N_13942);
or UO_798 (O_798,N_12159,N_13162);
and UO_799 (O_799,N_14928,N_14905);
xnor UO_800 (O_800,N_14603,N_13744);
or UO_801 (O_801,N_14046,N_12856);
or UO_802 (O_802,N_12449,N_12336);
nor UO_803 (O_803,N_13168,N_14303);
or UO_804 (O_804,N_12110,N_13598);
nand UO_805 (O_805,N_14252,N_14131);
nor UO_806 (O_806,N_13109,N_14261);
or UO_807 (O_807,N_14358,N_13803);
or UO_808 (O_808,N_13029,N_14149);
or UO_809 (O_809,N_13878,N_12172);
or UO_810 (O_810,N_13680,N_13465);
and UO_811 (O_811,N_14038,N_14709);
nand UO_812 (O_812,N_13437,N_12108);
and UO_813 (O_813,N_14164,N_14521);
nor UO_814 (O_814,N_14170,N_12236);
nor UO_815 (O_815,N_13704,N_12795);
nand UO_816 (O_816,N_13427,N_12671);
nand UO_817 (O_817,N_13507,N_14502);
nand UO_818 (O_818,N_12216,N_13594);
nor UO_819 (O_819,N_12826,N_14517);
nor UO_820 (O_820,N_14111,N_12253);
nand UO_821 (O_821,N_12830,N_13730);
nor UO_822 (O_822,N_13716,N_13236);
nor UO_823 (O_823,N_12415,N_12126);
or UO_824 (O_824,N_13777,N_13003);
or UO_825 (O_825,N_13555,N_14799);
or UO_826 (O_826,N_14743,N_14506);
nand UO_827 (O_827,N_13987,N_12322);
nand UO_828 (O_828,N_13520,N_13670);
or UO_829 (O_829,N_14943,N_12218);
or UO_830 (O_830,N_13828,N_12775);
or UO_831 (O_831,N_12891,N_13864);
or UO_832 (O_832,N_13875,N_14468);
and UO_833 (O_833,N_12585,N_13318);
nor UO_834 (O_834,N_12460,N_12673);
or UO_835 (O_835,N_13163,N_14370);
nand UO_836 (O_836,N_12516,N_12699);
or UO_837 (O_837,N_13073,N_12343);
or UO_838 (O_838,N_14476,N_13293);
nor UO_839 (O_839,N_13669,N_14531);
or UO_840 (O_840,N_14936,N_12445);
nand UO_841 (O_841,N_12767,N_14225);
nor UO_842 (O_842,N_14116,N_12169);
nand UO_843 (O_843,N_12576,N_13728);
nand UO_844 (O_844,N_14137,N_14562);
nand UO_845 (O_845,N_13673,N_12468);
xor UO_846 (O_846,N_12199,N_13086);
or UO_847 (O_847,N_12710,N_14216);
and UO_848 (O_848,N_13007,N_14505);
nand UO_849 (O_849,N_13434,N_13088);
or UO_850 (O_850,N_13159,N_12078);
or UO_851 (O_851,N_13860,N_13899);
nor UO_852 (O_852,N_13499,N_13233);
nor UO_853 (O_853,N_13419,N_12346);
or UO_854 (O_854,N_14295,N_13136);
nor UO_855 (O_855,N_14795,N_12917);
nand UO_856 (O_856,N_13588,N_12390);
xor UO_857 (O_857,N_12654,N_12861);
xor UO_858 (O_858,N_12052,N_14670);
and UO_859 (O_859,N_12001,N_13615);
and UO_860 (O_860,N_14343,N_13825);
or UO_861 (O_861,N_13415,N_13542);
nand UO_862 (O_862,N_12972,N_13812);
or UO_863 (O_863,N_12547,N_12965);
nand UO_864 (O_864,N_13834,N_12906);
or UO_865 (O_865,N_14820,N_14076);
nor UO_866 (O_866,N_12774,N_14461);
nor UO_867 (O_867,N_13015,N_13539);
or UO_868 (O_868,N_14493,N_14867);
nand UO_869 (O_869,N_14525,N_13582);
or UO_870 (O_870,N_13446,N_12687);
nand UO_871 (O_871,N_13997,N_12611);
and UO_872 (O_872,N_13988,N_12568);
and UO_873 (O_873,N_12437,N_14215);
nand UO_874 (O_874,N_13621,N_13447);
and UO_875 (O_875,N_13765,N_12653);
nand UO_876 (O_876,N_12864,N_12520);
nand UO_877 (O_877,N_12766,N_14639);
nor UO_878 (O_878,N_13336,N_14346);
nor UO_879 (O_879,N_14551,N_13756);
and UO_880 (O_880,N_14721,N_14033);
and UO_881 (O_881,N_14147,N_13586);
nand UO_882 (O_882,N_14056,N_12565);
nor UO_883 (O_883,N_14664,N_12299);
nand UO_884 (O_884,N_13190,N_14237);
and UO_885 (O_885,N_14035,N_12990);
nor UO_886 (O_886,N_12496,N_14339);
and UO_887 (O_887,N_12763,N_12112);
or UO_888 (O_888,N_12130,N_13310);
and UO_889 (O_889,N_14148,N_12123);
nor UO_890 (O_890,N_13848,N_12101);
or UO_891 (O_891,N_13729,N_14744);
and UO_892 (O_892,N_13247,N_14172);
nor UO_893 (O_893,N_12740,N_12037);
nor UO_894 (O_894,N_12189,N_13348);
or UO_895 (O_895,N_14407,N_13141);
nand UO_896 (O_896,N_14868,N_13734);
and UO_897 (O_897,N_14549,N_13455);
nand UO_898 (O_898,N_14214,N_13862);
and UO_899 (O_899,N_12196,N_12488);
and UO_900 (O_900,N_12624,N_12939);
nand UO_901 (O_901,N_12918,N_12361);
nor UO_902 (O_902,N_14813,N_13453);
nand UO_903 (O_903,N_13595,N_13535);
or UO_904 (O_904,N_12777,N_14540);
nor UO_905 (O_905,N_13271,N_13941);
and UO_906 (O_906,N_13137,N_14120);
nand UO_907 (O_907,N_14186,N_13442);
and UO_908 (O_908,N_12143,N_14641);
nand UO_909 (O_909,N_12049,N_14842);
nand UO_910 (O_910,N_12125,N_14732);
and UO_911 (O_911,N_13609,N_12260);
nand UO_912 (O_912,N_12827,N_12676);
or UO_913 (O_913,N_12204,N_13388);
nor UO_914 (O_914,N_14212,N_13546);
and UO_915 (O_915,N_13265,N_13045);
and UO_916 (O_916,N_12094,N_12866);
nand UO_917 (O_917,N_14951,N_13973);
or UO_918 (O_918,N_12893,N_12898);
nand UO_919 (O_919,N_12025,N_12041);
and UO_920 (O_920,N_12422,N_12277);
nor UO_921 (O_921,N_12521,N_13491);
nand UO_922 (O_922,N_13526,N_12600);
and UO_923 (O_923,N_13127,N_12083);
nor UO_924 (O_924,N_14331,N_12879);
nor UO_925 (O_925,N_13494,N_14372);
and UO_926 (O_926,N_12780,N_14145);
nand UO_927 (O_927,N_14792,N_12630);
nand UO_928 (O_928,N_13345,N_14118);
or UO_929 (O_929,N_13917,N_14090);
nand UO_930 (O_930,N_14864,N_14996);
nor UO_931 (O_931,N_12375,N_12874);
and UO_932 (O_932,N_14161,N_12814);
nor UO_933 (O_933,N_12706,N_14103);
or UO_934 (O_934,N_14368,N_12208);
nor UO_935 (O_935,N_14745,N_13273);
nor UO_936 (O_936,N_13489,N_13275);
nand UO_937 (O_937,N_14611,N_13721);
and UO_938 (O_938,N_14051,N_13170);
or UO_939 (O_939,N_14213,N_12161);
nand UO_940 (O_940,N_14906,N_12790);
nor UO_941 (O_941,N_13013,N_14326);
and UO_942 (O_942,N_12617,N_12544);
nand UO_943 (O_943,N_12914,N_13041);
nor UO_944 (O_944,N_14241,N_12239);
nor UO_945 (O_945,N_12113,N_14442);
nor UO_946 (O_946,N_12643,N_12819);
nand UO_947 (O_947,N_14885,N_12938);
and UO_948 (O_948,N_12754,N_12355);
or UO_949 (O_949,N_14742,N_14281);
nand UO_950 (O_950,N_12451,N_13840);
nand UO_951 (O_951,N_12787,N_14691);
and UO_952 (O_952,N_12197,N_13142);
nand UO_953 (O_953,N_13591,N_14572);
nand UO_954 (O_954,N_12213,N_12945);
and UO_955 (O_955,N_12723,N_14242);
nand UO_956 (O_956,N_12987,N_13059);
nand UO_957 (O_957,N_13886,N_14853);
or UO_958 (O_958,N_12967,N_14558);
or UO_959 (O_959,N_14872,N_13075);
or UO_960 (O_960,N_14821,N_12146);
nand UO_961 (O_961,N_14048,N_13713);
nand UO_962 (O_962,N_12479,N_13813);
nor UO_963 (O_963,N_14378,N_13657);
nor UO_964 (O_964,N_13587,N_12952);
or UO_965 (O_965,N_12765,N_14624);
or UO_966 (O_966,N_14477,N_12356);
nand UO_967 (O_967,N_12736,N_13202);
nand UO_968 (O_968,N_14656,N_12093);
and UO_969 (O_969,N_14777,N_14011);
nand UO_970 (O_970,N_13719,N_12745);
nor UO_971 (O_971,N_13731,N_13387);
nor UO_972 (O_972,N_14066,N_12974);
nand UO_973 (O_973,N_12503,N_14527);
nor UO_974 (O_974,N_12916,N_12288);
nand UO_975 (O_975,N_14981,N_13885);
nand UO_976 (O_976,N_12688,N_13892);
nor UO_977 (O_977,N_12533,N_14203);
nand UO_978 (O_978,N_12807,N_14547);
nand UO_979 (O_979,N_13733,N_14862);
nand UO_980 (O_980,N_13140,N_13748);
or UO_981 (O_981,N_13260,N_14615);
and UO_982 (O_982,N_13337,N_14079);
nor UO_983 (O_983,N_13568,N_13226);
and UO_984 (O_984,N_14104,N_12241);
nor UO_985 (O_985,N_13085,N_13529);
nor UO_986 (O_986,N_14567,N_13648);
nor UO_987 (O_987,N_14883,N_13540);
or UO_988 (O_988,N_12491,N_13334);
nor UO_989 (O_989,N_14160,N_12447);
nor UO_990 (O_990,N_14082,N_12757);
and UO_991 (O_991,N_14462,N_14217);
nor UO_992 (O_992,N_12964,N_12895);
nor UO_993 (O_993,N_13703,N_13482);
and UO_994 (O_994,N_13647,N_12439);
nand UO_995 (O_995,N_13024,N_13532);
and UO_996 (O_996,N_12536,N_12349);
nor UO_997 (O_997,N_12261,N_12133);
and UO_998 (O_998,N_14005,N_14794);
nor UO_999 (O_999,N_14421,N_13500);
nand UO_1000 (O_1000,N_14588,N_14459);
xor UO_1001 (O_1001,N_14945,N_13930);
or UO_1002 (O_1002,N_14272,N_14984);
nand UO_1003 (O_1003,N_13832,N_13604);
nor UO_1004 (O_1004,N_13916,N_12301);
nor UO_1005 (O_1005,N_12217,N_12823);
and UO_1006 (O_1006,N_14211,N_13321);
or UO_1007 (O_1007,N_12661,N_14892);
and UO_1008 (O_1008,N_12430,N_14846);
nor UO_1009 (O_1009,N_13331,N_14626);
or UO_1010 (O_1010,N_12266,N_12097);
or UO_1011 (O_1011,N_14600,N_13618);
nor UO_1012 (O_1012,N_12269,N_14182);
and UO_1013 (O_1013,N_14667,N_13682);
or UO_1014 (O_1014,N_14291,N_12821);
nor UO_1015 (O_1015,N_12022,N_12876);
nand UO_1016 (O_1016,N_13758,N_13943);
nor UO_1017 (O_1017,N_12257,N_13583);
nand UO_1018 (O_1018,N_14069,N_13742);
nor UO_1019 (O_1019,N_14565,N_13636);
nor UO_1020 (O_1020,N_13612,N_14430);
nor UO_1021 (O_1021,N_14962,N_14226);
xnor UO_1022 (O_1022,N_13853,N_14727);
nor UO_1023 (O_1023,N_14418,N_13444);
nor UO_1024 (O_1024,N_12018,N_14698);
or UO_1025 (O_1025,N_14904,N_13562);
nand UO_1026 (O_1026,N_14330,N_14628);
or UO_1027 (O_1027,N_12268,N_14024);
nand UO_1028 (O_1028,N_14849,N_12229);
nand UO_1029 (O_1029,N_12744,N_14650);
nor UO_1030 (O_1030,N_12004,N_13821);
nand UO_1031 (O_1031,N_13893,N_13553);
nor UO_1032 (O_1032,N_13416,N_14570);
and UO_1033 (O_1033,N_13058,N_14091);
nor UO_1034 (O_1034,N_12098,N_12751);
or UO_1035 (O_1035,N_13566,N_14224);
or UO_1036 (O_1036,N_13785,N_12835);
or UO_1037 (O_1037,N_12857,N_13101);
nand UO_1038 (O_1038,N_13855,N_14238);
and UO_1039 (O_1039,N_12954,N_14814);
nand UO_1040 (O_1040,N_12305,N_13651);
or UO_1041 (O_1041,N_14458,N_13315);
or UO_1042 (O_1042,N_12147,N_14524);
or UO_1043 (O_1043,N_12925,N_12984);
and UO_1044 (O_1044,N_12626,N_13871);
or UO_1045 (O_1045,N_13890,N_12677);
and UO_1046 (O_1046,N_12619,N_13608);
and UO_1047 (O_1047,N_13031,N_14632);
or UO_1048 (O_1048,N_14207,N_13188);
xnor UO_1049 (O_1049,N_13431,N_14723);
and UO_1050 (O_1050,N_14398,N_12507);
nor UO_1051 (O_1051,N_12118,N_13502);
nand UO_1052 (O_1052,N_12848,N_14127);
and UO_1053 (O_1053,N_12571,N_14806);
and UO_1054 (O_1054,N_13778,N_12039);
nand UO_1055 (O_1055,N_14900,N_14661);
xnor UO_1056 (O_1056,N_12804,N_14784);
and UO_1057 (O_1057,N_14590,N_12506);
and UO_1058 (O_1058,N_12854,N_12749);
nor UO_1059 (O_1059,N_12707,N_13961);
and UO_1060 (O_1060,N_14835,N_13688);
or UO_1061 (O_1061,N_12214,N_14873);
or UO_1062 (O_1062,N_13667,N_13863);
nand UO_1063 (O_1063,N_13600,N_13977);
nor UO_1064 (O_1064,N_12589,N_12587);
or UO_1065 (O_1065,N_13629,N_13055);
nor UO_1066 (O_1066,N_13456,N_13213);
and UO_1067 (O_1067,N_13150,N_13551);
xnor UO_1068 (O_1068,N_12962,N_14271);
nor UO_1069 (O_1069,N_12808,N_14940);
or UO_1070 (O_1070,N_13301,N_14383);
nand UO_1071 (O_1071,N_14397,N_12625);
or UO_1072 (O_1072,N_13580,N_13573);
or UO_1073 (O_1073,N_14651,N_13102);
nor UO_1074 (O_1074,N_12552,N_12009);
or UO_1075 (O_1075,N_14328,N_14538);
or UO_1076 (O_1076,N_12045,N_12758);
or UO_1077 (O_1077,N_13276,N_12801);
nor UO_1078 (O_1078,N_12947,N_13695);
nor UO_1079 (O_1079,N_13078,N_12235);
and UO_1080 (O_1080,N_13263,N_12514);
nand UO_1081 (O_1081,N_14539,N_14454);
and UO_1082 (O_1082,N_13161,N_12635);
nand UO_1083 (O_1083,N_12201,N_12427);
and UO_1084 (O_1084,N_14585,N_13454);
nand UO_1085 (O_1085,N_12762,N_13401);
and UO_1086 (O_1086,N_12728,N_14365);
nor UO_1087 (O_1087,N_12586,N_14703);
nand UO_1088 (O_1088,N_12667,N_12910);
or UO_1089 (O_1089,N_12632,N_12271);
nand UO_1090 (O_1090,N_13564,N_12378);
or UO_1091 (O_1091,N_13278,N_12486);
and UO_1092 (O_1092,N_12622,N_14054);
or UO_1093 (O_1093,N_12768,N_12050);
or UO_1094 (O_1094,N_13200,N_12651);
and UO_1095 (O_1095,N_13706,N_12285);
nor UO_1096 (O_1096,N_13611,N_14469);
nand UO_1097 (O_1097,N_13723,N_14036);
nor UO_1098 (O_1098,N_12393,N_12362);
xnor UO_1099 (O_1099,N_13281,N_14589);
or UO_1100 (O_1100,N_14684,N_14400);
or UO_1101 (O_1101,N_12026,N_13938);
nor UO_1102 (O_1102,N_12114,N_14859);
nor UO_1103 (O_1103,N_14379,N_12176);
or UO_1104 (O_1104,N_14654,N_12016);
nand UO_1105 (O_1105,N_14201,N_13676);
nor UO_1106 (O_1106,N_14992,N_13472);
nand UO_1107 (O_1107,N_13585,N_13438);
nand UO_1108 (O_1108,N_12453,N_14055);
or UO_1109 (O_1109,N_12881,N_12725);
nor UO_1110 (O_1110,N_12577,N_12722);
nand UO_1111 (O_1111,N_12055,N_12155);
nor UO_1112 (O_1112,N_13687,N_13083);
and UO_1113 (O_1113,N_13001,N_14228);
or UO_1114 (O_1114,N_14629,N_14979);
nand UO_1115 (O_1115,N_14605,N_12012);
nand UO_1116 (O_1116,N_14619,N_14119);
nand UO_1117 (O_1117,N_13139,N_12335);
or UO_1118 (O_1118,N_13279,N_14020);
and UO_1119 (O_1119,N_14676,N_14497);
and UO_1120 (O_1120,N_13495,N_12832);
nand UO_1121 (O_1121,N_12868,N_12373);
and UO_1122 (O_1122,N_12753,N_13693);
and UO_1123 (O_1123,N_14955,N_14602);
nor UO_1124 (O_1124,N_12596,N_14808);
nor UO_1125 (O_1125,N_14408,N_13993);
and UO_1126 (O_1126,N_12636,N_14662);
and UO_1127 (O_1127,N_13439,N_12693);
nand UO_1128 (O_1128,N_14156,N_13652);
or UO_1129 (O_1129,N_13084,N_12245);
and UO_1130 (O_1130,N_12760,N_14007);
and UO_1131 (O_1131,N_14865,N_13232);
nand UO_1132 (O_1132,N_12073,N_14878);
nor UO_1133 (O_1133,N_12407,N_12540);
nor UO_1134 (O_1134,N_13672,N_13836);
and UO_1135 (O_1135,N_13940,N_13931);
nand UO_1136 (O_1136,N_14440,N_13324);
nand UO_1137 (O_1137,N_14854,N_13654);
and UO_1138 (O_1138,N_12554,N_13847);
nor UO_1139 (O_1139,N_13361,N_13487);
and UO_1140 (O_1140,N_13412,N_14942);
or UO_1141 (O_1141,N_12476,N_12669);
or UO_1142 (O_1142,N_13118,N_12681);
and UO_1143 (O_1143,N_14192,N_14834);
nand UO_1144 (O_1144,N_12404,N_14921);
and UO_1145 (O_1145,N_14747,N_13915);
and UO_1146 (O_1146,N_13933,N_12478);
nand UO_1147 (O_1147,N_12701,N_13773);
nand UO_1148 (O_1148,N_12924,N_12946);
or UO_1149 (O_1149,N_12076,N_12609);
or UO_1150 (O_1150,N_13390,N_14674);
and UO_1151 (O_1151,N_14997,N_14944);
nor UO_1152 (O_1152,N_13714,N_13992);
nand UO_1153 (O_1153,N_14815,N_13189);
and UO_1154 (O_1154,N_13913,N_14016);
or UO_1155 (O_1155,N_12369,N_13999);
nand UO_1156 (O_1156,N_14482,N_12314);
nor UO_1157 (O_1157,N_13282,N_13752);
nor UO_1158 (O_1158,N_12377,N_14042);
or UO_1159 (O_1159,N_13468,N_13675);
nor UO_1160 (O_1160,N_12800,N_13571);
and UO_1161 (O_1161,N_13792,N_14687);
xnor UO_1162 (O_1162,N_14720,N_13074);
nand UO_1163 (O_1163,N_12099,N_14044);
or UO_1164 (O_1164,N_14075,N_13422);
nand UO_1165 (O_1165,N_12485,N_13026);
and UO_1166 (O_1166,N_14264,N_13630);
or UO_1167 (O_1167,N_12287,N_13996);
nand UO_1168 (O_1168,N_13876,N_13076);
or UO_1169 (O_1169,N_14236,N_13179);
nor UO_1170 (O_1170,N_12224,N_14144);
and UO_1171 (O_1171,N_13399,N_12467);
or UO_1172 (O_1172,N_13234,N_14881);
and UO_1173 (O_1173,N_13810,N_14487);
nand UO_1174 (O_1174,N_14740,N_13726);
nor UO_1175 (O_1175,N_12877,N_14668);
or UO_1176 (O_1176,N_12992,N_12381);
nor UO_1177 (O_1177,N_13049,N_14861);
nand UO_1178 (O_1178,N_12604,N_12580);
nor UO_1179 (O_1179,N_12329,N_14415);
and UO_1180 (O_1180,N_14157,N_13537);
nand UO_1181 (O_1181,N_13552,N_12784);
nor UO_1182 (O_1182,N_14621,N_13481);
or UO_1183 (O_1183,N_14925,N_12103);
or UO_1184 (O_1184,N_14989,N_14986);
or UO_1185 (O_1185,N_14770,N_12531);
nand UO_1186 (O_1186,N_14168,N_12034);
nand UO_1187 (O_1187,N_12537,N_13590);
and UO_1188 (O_1188,N_14518,N_13798);
or UO_1189 (O_1189,N_14336,N_14087);
or UO_1190 (O_1190,N_13246,N_12401);
or UO_1191 (O_1191,N_13152,N_13613);
or UO_1192 (O_1192,N_13144,N_13149);
or UO_1193 (O_1193,N_13606,N_13095);
and UO_1194 (O_1194,N_12989,N_13775);
or UO_1195 (O_1195,N_14736,N_13181);
nor UO_1196 (O_1196,N_13547,N_13287);
and UO_1197 (O_1197,N_13628,N_14909);
nor UO_1198 (O_1198,N_12380,N_13242);
xor UO_1199 (O_1199,N_14246,N_12124);
nand UO_1200 (O_1200,N_14466,N_12679);
and UO_1201 (O_1201,N_12338,N_12036);
nor UO_1202 (O_1202,N_13793,N_12880);
nor UO_1203 (O_1203,N_13251,N_14394);
or UO_1204 (O_1204,N_14023,N_14490);
or UO_1205 (O_1205,N_13018,N_13277);
or UO_1206 (O_1206,N_14573,N_14451);
and UO_1207 (O_1207,N_12187,N_13192);
and UO_1208 (O_1208,N_14939,N_12480);
nor UO_1209 (O_1209,N_14486,N_13385);
and UO_1210 (O_1210,N_13156,N_13354);
and UO_1211 (O_1211,N_14894,N_12779);
and UO_1212 (O_1212,N_13222,N_13436);
nand UO_1213 (O_1213,N_12284,N_14957);
xnor UO_1214 (O_1214,N_13463,N_13008);
or UO_1215 (O_1215,N_12364,N_12562);
nor UO_1216 (O_1216,N_13025,N_13080);
or UO_1217 (O_1217,N_14473,N_13476);
nand UO_1218 (O_1218,N_14912,N_14478);
nand UO_1219 (O_1219,N_12716,N_13203);
nor UO_1220 (O_1220,N_13107,N_12077);
nand UO_1221 (O_1221,N_12698,N_14018);
and UO_1222 (O_1222,N_13851,N_13497);
nor UO_1223 (O_1223,N_12709,N_12115);
xnor UO_1224 (O_1224,N_14832,N_13490);
or UO_1225 (O_1225,N_14645,N_13791);
or UO_1226 (O_1226,N_13298,N_13768);
nor UO_1227 (O_1227,N_12743,N_12310);
nor UO_1228 (O_1228,N_14594,N_14095);
and UO_1229 (O_1229,N_14335,N_14811);
nand UO_1230 (O_1230,N_13898,N_12263);
or UO_1231 (O_1231,N_14196,N_12056);
or UO_1232 (O_1232,N_13989,N_14074);
nor UO_1233 (O_1233,N_12792,N_12966);
nand UO_1234 (O_1234,N_12011,N_13426);
nor UO_1235 (O_1235,N_12773,N_12702);
nand UO_1236 (O_1236,N_13712,N_13879);
nand UO_1237 (O_1237,N_14791,N_14257);
and UO_1238 (O_1238,N_13737,N_13718);
nand UO_1239 (O_1239,N_12539,N_14959);
and UO_1240 (O_1240,N_14965,N_12712);
and UO_1241 (O_1241,N_12852,N_13677);
xnor UO_1242 (O_1242,N_14350,N_14361);
nand UO_1243 (O_1243,N_14908,N_13171);
xor UO_1244 (O_1244,N_14903,N_12162);
nand UO_1245 (O_1245,N_13204,N_13220);
nor UO_1246 (O_1246,N_14138,N_14715);
or UO_1247 (O_1247,N_14159,N_14752);
nor UO_1248 (O_1248,N_13528,N_14040);
or UO_1249 (O_1249,N_13932,N_14591);
and UO_1250 (O_1250,N_14334,N_12167);
nor UO_1251 (O_1251,N_13364,N_14107);
nand UO_1252 (O_1252,N_14708,N_13751);
and UO_1253 (O_1253,N_12759,N_13971);
or UO_1254 (O_1254,N_12871,N_14542);
and UO_1255 (O_1255,N_13035,N_12645);
or UO_1256 (O_1256,N_13806,N_12936);
nand UO_1257 (O_1257,N_13660,N_12008);
xnor UO_1258 (O_1258,N_12209,N_13603);
nor UO_1259 (O_1259,N_12360,N_12658);
and UO_1260 (O_1260,N_12704,N_14533);
and UO_1261 (O_1261,N_13841,N_13513);
nor UO_1262 (O_1262,N_12294,N_14019);
and UO_1263 (O_1263,N_13254,N_13359);
nor UO_1264 (O_1264,N_12286,N_12844);
or UO_1265 (O_1265,N_14526,N_13079);
nor UO_1266 (O_1266,N_13671,N_14528);
xnor UO_1267 (O_1267,N_12932,N_13934);
nand UO_1268 (O_1268,N_14786,N_13121);
nor UO_1269 (O_1269,N_12262,N_14162);
nand UO_1270 (O_1270,N_14683,N_13850);
and UO_1271 (O_1271,N_14860,N_14096);
xnor UO_1272 (O_1272,N_12518,N_14320);
or UO_1273 (O_1273,N_14178,N_14010);
and UO_1274 (O_1274,N_12983,N_13316);
nand UO_1275 (O_1275,N_13858,N_12680);
nand UO_1276 (O_1276,N_12070,N_12560);
and UO_1277 (O_1277,N_14375,N_13967);
nand UO_1278 (O_1278,N_13889,N_12400);
nor UO_1279 (O_1279,N_13248,N_14206);
nand UO_1280 (O_1280,N_14187,N_13519);
nand UO_1281 (O_1281,N_14566,N_12428);
nand UO_1282 (O_1282,N_14920,N_13363);
and UO_1283 (O_1283,N_14447,N_12107);
or UO_1284 (O_1284,N_14796,N_12559);
or UO_1285 (O_1285,N_14750,N_14134);
xnor UO_1286 (O_1286,N_13377,N_14823);
nor UO_1287 (O_1287,N_13990,N_12021);
and UO_1288 (O_1288,N_13839,N_12027);
or UO_1289 (O_1289,N_12991,N_12031);
nor UO_1290 (O_1290,N_13514,N_13717);
nor UO_1291 (O_1291,N_14479,N_13014);
or UO_1292 (O_1292,N_12950,N_14801);
nor UO_1293 (O_1293,N_12405,N_12648);
nand UO_1294 (O_1294,N_12566,N_13804);
nand UO_1295 (O_1295,N_13027,N_12512);
nor UO_1296 (O_1296,N_12319,N_12599);
nand UO_1297 (O_1297,N_12692,N_14266);
nor UO_1298 (O_1298,N_14902,N_13905);
nand UO_1299 (O_1299,N_14154,N_14412);
or UO_1300 (O_1300,N_12482,N_12000);
and UO_1301 (O_1301,N_14776,N_13523);
or UO_1302 (O_1302,N_14960,N_14994);
and UO_1303 (O_1303,N_13435,N_12175);
or UO_1304 (O_1304,N_13554,N_12384);
xnor UO_1305 (O_1305,N_14764,N_14847);
nor UO_1306 (O_1306,N_14576,N_13854);
nand UO_1307 (O_1307,N_13954,N_12242);
or UO_1308 (O_1308,N_12545,N_13790);
and UO_1309 (O_1309,N_12303,N_13921);
or UO_1310 (O_1310,N_12157,N_14812);
nor UO_1311 (O_1311,N_14448,N_12330);
and UO_1312 (O_1312,N_14927,N_13258);
and UO_1313 (O_1313,N_12392,N_13175);
or UO_1314 (O_1314,N_13702,N_14704);
and UO_1315 (O_1315,N_13720,N_13072);
and UO_1316 (O_1316,N_14932,N_13197);
and UO_1317 (O_1317,N_14130,N_14309);
nand UO_1318 (O_1318,N_12769,N_14437);
nand UO_1319 (O_1319,N_14474,N_14452);
and UO_1320 (O_1320,N_13451,N_13506);
xnor UO_1321 (O_1321,N_12927,N_14306);
or UO_1322 (O_1322,N_12526,N_12509);
or UO_1323 (O_1323,N_12715,N_12212);
or UO_1324 (O_1324,N_13884,N_12421);
nor UO_1325 (O_1325,N_13462,N_13809);
nand UO_1326 (O_1326,N_13801,N_14991);
or UO_1327 (O_1327,N_14251,N_13509);
and UO_1328 (O_1328,N_12254,N_13576);
nor UO_1329 (O_1329,N_12598,N_14751);
nand UO_1330 (O_1330,N_13634,N_13565);
or UO_1331 (O_1331,N_14891,N_13384);
or UO_1332 (O_1332,N_12606,N_12332);
nand UO_1333 (O_1333,N_12558,N_12372);
or UO_1334 (O_1334,N_13543,N_14077);
nand UO_1335 (O_1335,N_13341,N_12200);
or UO_1336 (O_1336,N_13343,N_12943);
nand UO_1337 (O_1337,N_12230,N_13901);
nand UO_1338 (O_1338,N_12180,N_12612);
and UO_1339 (O_1339,N_12345,N_12252);
or UO_1340 (O_1340,N_12602,N_14380);
and UO_1341 (O_1341,N_13250,N_13725);
and UO_1342 (O_1342,N_12296,N_13567);
nand UO_1343 (O_1343,N_13229,N_13400);
nand UO_1344 (O_1344,N_12170,N_12359);
xnor UO_1345 (O_1345,N_13332,N_13970);
and UO_1346 (O_1346,N_14617,N_13767);
nor UO_1347 (O_1347,N_12472,N_13474);
nor UO_1348 (O_1348,N_14371,N_12354);
nand UO_1349 (O_1349,N_14089,N_12665);
or UO_1350 (O_1350,N_13064,N_13325);
nor UO_1351 (O_1351,N_13816,N_13946);
nand UO_1352 (O_1352,N_13120,N_14052);
or UO_1353 (O_1353,N_14746,N_14930);
and UO_1354 (O_1354,N_14110,N_12508);
nor UO_1355 (O_1355,N_12267,N_14453);
nor UO_1356 (O_1356,N_14665,N_13548);
nand UO_1357 (O_1357,N_12551,N_12629);
and UO_1358 (O_1358,N_12556,N_12386);
nor UO_1359 (O_1359,N_12931,N_14512);
or UO_1360 (O_1360,N_12892,N_12185);
nor UO_1361 (O_1361,N_14671,N_12064);
or UO_1362 (O_1362,N_12414,N_14785);
and UO_1363 (O_1363,N_12316,N_14680);
and UO_1364 (O_1364,N_12122,N_13167);
nor UO_1365 (O_1365,N_13518,N_14369);
nand UO_1366 (O_1366,N_13605,N_13099);
nand UO_1367 (O_1367,N_14193,N_13982);
nor UO_1368 (O_1368,N_13935,N_13467);
and UO_1369 (O_1369,N_14756,N_14387);
or UO_1370 (O_1370,N_14464,N_14682);
nand UO_1371 (O_1371,N_12920,N_14515);
or UO_1372 (O_1372,N_13440,N_12248);
and UO_1373 (O_1373,N_14436,N_12529);
or UO_1374 (O_1374,N_12561,N_14800);
and UO_1375 (O_1375,N_12605,N_14229);
nand UO_1376 (O_1376,N_13373,N_12998);
nor UO_1377 (O_1377,N_12996,N_12505);
or UO_1378 (O_1378,N_14122,N_13128);
and UO_1379 (O_1379,N_12799,N_14675);
nor UO_1380 (O_1380,N_12370,N_14101);
and UO_1381 (O_1381,N_14332,N_12206);
nand UO_1382 (O_1382,N_13797,N_13285);
and UO_1383 (O_1383,N_14278,N_12383);
or UO_1384 (O_1384,N_14924,N_14231);
or UO_1385 (O_1385,N_14317,N_14393);
and UO_1386 (O_1386,N_14062,N_13396);
nor UO_1387 (O_1387,N_13668,N_13957);
or UO_1388 (O_1388,N_12313,N_14414);
nand UO_1389 (O_1389,N_13974,N_14141);
and UO_1390 (O_1390,N_13182,N_14356);
or UO_1391 (O_1391,N_12371,N_12444);
or UO_1392 (O_1392,N_12907,N_12342);
nand UO_1393 (O_1393,N_14514,N_13779);
and UO_1394 (O_1394,N_13303,N_12859);
nor UO_1395 (O_1395,N_14907,N_12729);
and UO_1396 (O_1396,N_13859,N_12851);
nor UO_1397 (O_1397,N_14348,N_13037);
or UO_1398 (O_1398,N_12889,N_13857);
or UO_1399 (O_1399,N_13724,N_13912);
nand UO_1400 (O_1400,N_12227,N_12601);
nor UO_1401 (O_1401,N_13104,N_12470);
and UO_1402 (O_1402,N_13257,N_13421);
or UO_1403 (O_1403,N_12803,N_12672);
nand UO_1404 (O_1404,N_14604,N_13402);
or UO_1405 (O_1405,N_13900,N_12275);
xor UO_1406 (O_1406,N_12188,N_13764);
or UO_1407 (O_1407,N_14895,N_12249);
or UO_1408 (O_1408,N_12190,N_13409);
and UO_1409 (O_1409,N_12280,N_14622);
or UO_1410 (O_1410,N_14963,N_14169);
nor UO_1411 (O_1411,N_13153,N_12398);
nor UO_1412 (O_1412,N_13983,N_12862);
or UO_1413 (O_1413,N_12391,N_12156);
nand UO_1414 (O_1414,N_12981,N_13294);
and UO_1415 (O_1415,N_12549,N_14636);
nand UO_1416 (O_1416,N_14123,N_12690);
nor UO_1417 (O_1417,N_12711,N_13747);
nand UO_1418 (O_1418,N_14333,N_14324);
and UO_1419 (O_1419,N_14417,N_13678);
nor UO_1420 (O_1420,N_14391,N_12750);
or UO_1421 (O_1421,N_14060,N_14314);
nand UO_1422 (O_1422,N_13679,N_13460);
nor UO_1423 (O_1423,N_14106,N_12610);
or UO_1424 (O_1424,N_12413,N_12515);
nor UO_1425 (O_1425,N_12833,N_12289);
and UO_1426 (O_1426,N_12420,N_13766);
and UO_1427 (O_1427,N_13036,N_13030);
or UO_1428 (O_1428,N_13510,N_14092);
and UO_1429 (O_1429,N_13746,N_14510);
and UO_1430 (O_1430,N_13096,N_13522);
xor UO_1431 (O_1431,N_14659,N_12291);
nand UO_1432 (O_1432,N_14483,N_12899);
and UO_1433 (O_1433,N_14688,N_12493);
nor UO_1434 (O_1434,N_14969,N_12411);
nand UO_1435 (O_1435,N_14855,N_13056);
and UO_1436 (O_1436,N_13291,N_12040);
or UO_1437 (O_1437,N_13521,N_13093);
nor UO_1438 (O_1438,N_14511,N_12222);
nand UO_1439 (O_1439,N_13796,N_12191);
or UO_1440 (O_1440,N_14373,N_12501);
or UO_1441 (O_1441,N_12264,N_14876);
or UO_1442 (O_1442,N_12647,N_14185);
or UO_1443 (O_1443,N_14705,N_14260);
nand UO_1444 (O_1444,N_13852,N_14093);
and UO_1445 (O_1445,N_14652,N_13256);
nor UO_1446 (O_1446,N_13306,N_13272);
or UO_1447 (O_1447,N_14030,N_14449);
nand UO_1448 (O_1448,N_14677,N_14403);
nor UO_1449 (O_1449,N_13581,N_14227);
nand UO_1450 (O_1450,N_12306,N_14443);
xor UO_1451 (O_1451,N_12664,N_14423);
nand UO_1452 (O_1452,N_12054,N_14546);
or UO_1453 (O_1453,N_12071,N_13184);
and UO_1454 (O_1454,N_12934,N_13690);
and UO_1455 (O_1455,N_12975,N_14898);
and UO_1456 (O_1456,N_13330,N_13681);
and UO_1457 (O_1457,N_12786,N_13215);
nor UO_1458 (O_1458,N_12471,N_13663);
nor UO_1459 (O_1459,N_13180,N_13822);
and UO_1460 (O_1460,N_12184,N_12942);
nor UO_1461 (O_1461,N_13980,N_12087);
nand UO_1462 (O_1462,N_14411,N_12092);
or UO_1463 (O_1463,N_13904,N_13349);
and UO_1464 (O_1464,N_14338,N_14467);
xnor UO_1465 (O_1465,N_12278,N_13561);
and UO_1466 (O_1466,N_14923,N_13219);
and UO_1467 (O_1467,N_14685,N_13517);
nor UO_1468 (O_1468,N_14460,N_12696);
and UO_1469 (O_1469,N_14958,N_14061);
or UO_1470 (O_1470,N_14302,N_12494);
nor UO_1471 (O_1471,N_13925,N_14804);
nand UO_1472 (O_1472,N_12458,N_13755);
or UO_1473 (O_1473,N_12419,N_12960);
nor UO_1474 (O_1474,N_14513,N_14321);
nand UO_1475 (O_1475,N_14340,N_14247);
xor UO_1476 (O_1476,N_14917,N_12922);
nand UO_1477 (O_1477,N_13160,N_12772);
or UO_1478 (O_1478,N_13662,N_12051);
and UO_1479 (O_1479,N_12308,N_13417);
nor UO_1480 (O_1480,N_13685,N_12761);
nand UO_1481 (O_1481,N_13155,N_13740);
or UO_1482 (O_1482,N_12828,N_12032);
and UO_1483 (O_1483,N_13811,N_14586);
nor UO_1484 (O_1484,N_12642,N_12148);
or UO_1485 (O_1485,N_12809,N_13302);
or UO_1486 (O_1486,N_12292,N_14315);
nand UO_1487 (O_1487,N_13995,N_12326);
nor UO_1488 (O_1488,N_13557,N_12477);
nor UO_1489 (O_1489,N_13817,N_12721);
nand UO_1490 (O_1490,N_12351,N_12324);
nor UO_1491 (O_1491,N_13953,N_13394);
nand UO_1492 (O_1492,N_14810,N_13838);
nor UO_1493 (O_1493,N_13708,N_12456);
nor UO_1494 (O_1494,N_14759,N_14166);
nor UO_1495 (O_1495,N_14733,N_13381);
nand UO_1496 (O_1496,N_14507,N_14571);
nor UO_1497 (O_1497,N_14599,N_13503);
nand UO_1498 (O_1498,N_12940,N_12944);
and UO_1499 (O_1499,N_13914,N_13738);
or UO_1500 (O_1500,N_14288,N_12634);
and UO_1501 (O_1501,N_14821,N_13707);
nand UO_1502 (O_1502,N_13309,N_14495);
or UO_1503 (O_1503,N_14465,N_13011);
nor UO_1504 (O_1504,N_14002,N_12202);
nor UO_1505 (O_1505,N_13593,N_12912);
or UO_1506 (O_1506,N_13869,N_14950);
nor UO_1507 (O_1507,N_13371,N_14093);
nor UO_1508 (O_1508,N_13053,N_13722);
nor UO_1509 (O_1509,N_12709,N_14618);
or UO_1510 (O_1510,N_14990,N_14067);
nor UO_1511 (O_1511,N_12069,N_14257);
nand UO_1512 (O_1512,N_13002,N_12421);
or UO_1513 (O_1513,N_13240,N_13716);
or UO_1514 (O_1514,N_13789,N_12273);
nand UO_1515 (O_1515,N_12795,N_13685);
nor UO_1516 (O_1516,N_14703,N_14527);
nand UO_1517 (O_1517,N_14906,N_14513);
or UO_1518 (O_1518,N_13770,N_12066);
or UO_1519 (O_1519,N_14700,N_13495);
nand UO_1520 (O_1520,N_12604,N_13872);
and UO_1521 (O_1521,N_14439,N_14274);
or UO_1522 (O_1522,N_13402,N_14599);
or UO_1523 (O_1523,N_12912,N_14131);
and UO_1524 (O_1524,N_12461,N_12508);
nand UO_1525 (O_1525,N_13774,N_12206);
or UO_1526 (O_1526,N_14986,N_14381);
nor UO_1527 (O_1527,N_12709,N_12456);
nor UO_1528 (O_1528,N_13997,N_14809);
nor UO_1529 (O_1529,N_13690,N_13201);
and UO_1530 (O_1530,N_12357,N_13951);
nand UO_1531 (O_1531,N_13425,N_14585);
nor UO_1532 (O_1532,N_14578,N_13084);
nand UO_1533 (O_1533,N_12696,N_13062);
nand UO_1534 (O_1534,N_12954,N_12480);
or UO_1535 (O_1535,N_14677,N_14569);
nand UO_1536 (O_1536,N_13462,N_14443);
nand UO_1537 (O_1537,N_12019,N_12772);
and UO_1538 (O_1538,N_14993,N_12595);
and UO_1539 (O_1539,N_14082,N_14718);
or UO_1540 (O_1540,N_12267,N_12637);
nor UO_1541 (O_1541,N_13513,N_13749);
and UO_1542 (O_1542,N_12918,N_14317);
and UO_1543 (O_1543,N_13960,N_13153);
or UO_1544 (O_1544,N_14204,N_14684);
or UO_1545 (O_1545,N_14645,N_14948);
nand UO_1546 (O_1546,N_14817,N_13009);
and UO_1547 (O_1547,N_12760,N_13611);
or UO_1548 (O_1548,N_12808,N_13272);
and UO_1549 (O_1549,N_13314,N_14454);
or UO_1550 (O_1550,N_14375,N_14564);
nor UO_1551 (O_1551,N_13357,N_13167);
nor UO_1552 (O_1552,N_13909,N_14963);
nand UO_1553 (O_1553,N_13367,N_13749);
nor UO_1554 (O_1554,N_12616,N_14093);
and UO_1555 (O_1555,N_13469,N_13974);
or UO_1556 (O_1556,N_13714,N_14191);
or UO_1557 (O_1557,N_12547,N_14924);
nand UO_1558 (O_1558,N_13441,N_13575);
or UO_1559 (O_1559,N_12100,N_12671);
and UO_1560 (O_1560,N_13084,N_13452);
and UO_1561 (O_1561,N_14192,N_14579);
and UO_1562 (O_1562,N_13357,N_13409);
or UO_1563 (O_1563,N_14760,N_12817);
and UO_1564 (O_1564,N_14047,N_14715);
nand UO_1565 (O_1565,N_13097,N_14687);
nand UO_1566 (O_1566,N_12367,N_12511);
or UO_1567 (O_1567,N_13301,N_12602);
nand UO_1568 (O_1568,N_14715,N_13700);
nor UO_1569 (O_1569,N_12387,N_12721);
and UO_1570 (O_1570,N_13303,N_12326);
nor UO_1571 (O_1571,N_14262,N_12979);
and UO_1572 (O_1572,N_12632,N_14385);
nand UO_1573 (O_1573,N_14830,N_13171);
nor UO_1574 (O_1574,N_14900,N_13329);
nand UO_1575 (O_1575,N_13066,N_14336);
nor UO_1576 (O_1576,N_14347,N_13711);
or UO_1577 (O_1577,N_14023,N_13655);
or UO_1578 (O_1578,N_14768,N_14771);
or UO_1579 (O_1579,N_12624,N_12946);
and UO_1580 (O_1580,N_12778,N_12377);
nor UO_1581 (O_1581,N_14372,N_12775);
nor UO_1582 (O_1582,N_13558,N_12141);
nor UO_1583 (O_1583,N_14874,N_14782);
nand UO_1584 (O_1584,N_14034,N_13833);
and UO_1585 (O_1585,N_14462,N_13475);
and UO_1586 (O_1586,N_12780,N_13216);
nor UO_1587 (O_1587,N_12446,N_14155);
nor UO_1588 (O_1588,N_12771,N_14635);
and UO_1589 (O_1589,N_12179,N_14387);
nor UO_1590 (O_1590,N_14423,N_13826);
nand UO_1591 (O_1591,N_14148,N_14859);
nand UO_1592 (O_1592,N_14715,N_12309);
nor UO_1593 (O_1593,N_12378,N_12820);
nor UO_1594 (O_1594,N_13799,N_13215);
and UO_1595 (O_1595,N_12855,N_13752);
or UO_1596 (O_1596,N_12785,N_12861);
or UO_1597 (O_1597,N_13782,N_12264);
nand UO_1598 (O_1598,N_13469,N_13292);
nor UO_1599 (O_1599,N_14132,N_14893);
nand UO_1600 (O_1600,N_13480,N_14686);
and UO_1601 (O_1601,N_14432,N_13692);
and UO_1602 (O_1602,N_12416,N_13912);
xnor UO_1603 (O_1603,N_12969,N_13823);
or UO_1604 (O_1604,N_12516,N_13062);
and UO_1605 (O_1605,N_12008,N_14492);
or UO_1606 (O_1606,N_12376,N_14678);
nor UO_1607 (O_1607,N_14097,N_13910);
nand UO_1608 (O_1608,N_14188,N_12910);
nand UO_1609 (O_1609,N_12244,N_12319);
nor UO_1610 (O_1610,N_12550,N_14029);
nor UO_1611 (O_1611,N_14724,N_14371);
and UO_1612 (O_1612,N_14583,N_13334);
nand UO_1613 (O_1613,N_13110,N_13115);
xor UO_1614 (O_1614,N_14615,N_12617);
and UO_1615 (O_1615,N_12452,N_12389);
or UO_1616 (O_1616,N_14891,N_12679);
and UO_1617 (O_1617,N_13297,N_13885);
or UO_1618 (O_1618,N_13219,N_12403);
and UO_1619 (O_1619,N_14181,N_13047);
nor UO_1620 (O_1620,N_13144,N_14875);
or UO_1621 (O_1621,N_13217,N_14534);
and UO_1622 (O_1622,N_13382,N_12879);
nand UO_1623 (O_1623,N_13505,N_12731);
nand UO_1624 (O_1624,N_12968,N_12466);
or UO_1625 (O_1625,N_14581,N_14569);
nor UO_1626 (O_1626,N_13013,N_14037);
nand UO_1627 (O_1627,N_12345,N_14231);
nor UO_1628 (O_1628,N_12214,N_13579);
and UO_1629 (O_1629,N_13395,N_13061);
and UO_1630 (O_1630,N_12220,N_14008);
nand UO_1631 (O_1631,N_14191,N_13640);
and UO_1632 (O_1632,N_13405,N_12064);
and UO_1633 (O_1633,N_12972,N_14019);
xor UO_1634 (O_1634,N_14274,N_13686);
nor UO_1635 (O_1635,N_14660,N_13522);
nor UO_1636 (O_1636,N_12296,N_12334);
nand UO_1637 (O_1637,N_14233,N_13229);
nand UO_1638 (O_1638,N_13035,N_13275);
or UO_1639 (O_1639,N_12774,N_12150);
and UO_1640 (O_1640,N_13032,N_12532);
or UO_1641 (O_1641,N_14602,N_12652);
or UO_1642 (O_1642,N_14047,N_13410);
nand UO_1643 (O_1643,N_12884,N_12194);
or UO_1644 (O_1644,N_12867,N_14128);
nor UO_1645 (O_1645,N_14534,N_12406);
and UO_1646 (O_1646,N_12373,N_13081);
or UO_1647 (O_1647,N_13982,N_13037);
nor UO_1648 (O_1648,N_13612,N_13760);
nand UO_1649 (O_1649,N_12773,N_13261);
and UO_1650 (O_1650,N_13772,N_12271);
and UO_1651 (O_1651,N_13458,N_12903);
nand UO_1652 (O_1652,N_12240,N_13747);
and UO_1653 (O_1653,N_14715,N_12074);
and UO_1654 (O_1654,N_12997,N_12234);
nor UO_1655 (O_1655,N_12087,N_13025);
or UO_1656 (O_1656,N_14658,N_12306);
and UO_1657 (O_1657,N_13273,N_13014);
and UO_1658 (O_1658,N_12948,N_14739);
or UO_1659 (O_1659,N_14830,N_13182);
and UO_1660 (O_1660,N_13355,N_13697);
and UO_1661 (O_1661,N_12119,N_12850);
nor UO_1662 (O_1662,N_14980,N_12509);
nor UO_1663 (O_1663,N_14094,N_13242);
or UO_1664 (O_1664,N_13574,N_14159);
or UO_1665 (O_1665,N_12573,N_14590);
or UO_1666 (O_1666,N_12169,N_14399);
or UO_1667 (O_1667,N_12769,N_12047);
nand UO_1668 (O_1668,N_12008,N_13920);
or UO_1669 (O_1669,N_14911,N_14164);
and UO_1670 (O_1670,N_12527,N_14959);
or UO_1671 (O_1671,N_14653,N_13127);
nand UO_1672 (O_1672,N_13519,N_14502);
and UO_1673 (O_1673,N_13017,N_12600);
nand UO_1674 (O_1674,N_14563,N_12607);
and UO_1675 (O_1675,N_13628,N_14065);
or UO_1676 (O_1676,N_14457,N_13424);
or UO_1677 (O_1677,N_12761,N_13540);
nor UO_1678 (O_1678,N_13802,N_12556);
or UO_1679 (O_1679,N_13183,N_12613);
nand UO_1680 (O_1680,N_14517,N_13203);
and UO_1681 (O_1681,N_14840,N_13951);
or UO_1682 (O_1682,N_13136,N_12349);
or UO_1683 (O_1683,N_13982,N_13175);
xor UO_1684 (O_1684,N_12552,N_13020);
and UO_1685 (O_1685,N_13706,N_14382);
xor UO_1686 (O_1686,N_12264,N_12112);
nand UO_1687 (O_1687,N_12245,N_13102);
nor UO_1688 (O_1688,N_14398,N_12381);
nand UO_1689 (O_1689,N_13878,N_13696);
or UO_1690 (O_1690,N_13488,N_12070);
or UO_1691 (O_1691,N_14174,N_12714);
and UO_1692 (O_1692,N_13454,N_13360);
nor UO_1693 (O_1693,N_14361,N_14782);
nand UO_1694 (O_1694,N_12575,N_13898);
nand UO_1695 (O_1695,N_14129,N_12409);
xnor UO_1696 (O_1696,N_13436,N_14404);
nand UO_1697 (O_1697,N_14924,N_13373);
nor UO_1698 (O_1698,N_13256,N_12396);
nand UO_1699 (O_1699,N_13334,N_12317);
nand UO_1700 (O_1700,N_12876,N_13040);
nor UO_1701 (O_1701,N_12275,N_12762);
nand UO_1702 (O_1702,N_14263,N_13661);
and UO_1703 (O_1703,N_13820,N_14259);
nand UO_1704 (O_1704,N_14198,N_12912);
nand UO_1705 (O_1705,N_13986,N_14563);
or UO_1706 (O_1706,N_14585,N_12749);
or UO_1707 (O_1707,N_13902,N_14399);
nor UO_1708 (O_1708,N_13969,N_12909);
nand UO_1709 (O_1709,N_12979,N_12740);
and UO_1710 (O_1710,N_14389,N_14775);
nand UO_1711 (O_1711,N_13387,N_14886);
xor UO_1712 (O_1712,N_12670,N_12497);
and UO_1713 (O_1713,N_12570,N_14727);
and UO_1714 (O_1714,N_13578,N_14872);
or UO_1715 (O_1715,N_13946,N_14194);
or UO_1716 (O_1716,N_12243,N_13468);
or UO_1717 (O_1717,N_12920,N_13368);
nand UO_1718 (O_1718,N_13585,N_13028);
and UO_1719 (O_1719,N_14229,N_13363);
nor UO_1720 (O_1720,N_14003,N_14156);
nand UO_1721 (O_1721,N_13261,N_14167);
nor UO_1722 (O_1722,N_12529,N_13777);
or UO_1723 (O_1723,N_12844,N_13221);
nor UO_1724 (O_1724,N_13509,N_12576);
nand UO_1725 (O_1725,N_12844,N_14307);
or UO_1726 (O_1726,N_13995,N_13683);
or UO_1727 (O_1727,N_12790,N_13447);
nor UO_1728 (O_1728,N_13265,N_12917);
or UO_1729 (O_1729,N_12837,N_13342);
nor UO_1730 (O_1730,N_12461,N_13560);
xor UO_1731 (O_1731,N_13673,N_14807);
nor UO_1732 (O_1732,N_14274,N_13442);
or UO_1733 (O_1733,N_14413,N_12444);
or UO_1734 (O_1734,N_12054,N_14339);
nor UO_1735 (O_1735,N_14858,N_12256);
nor UO_1736 (O_1736,N_12781,N_13446);
nand UO_1737 (O_1737,N_14424,N_14917);
or UO_1738 (O_1738,N_14229,N_12827);
nor UO_1739 (O_1739,N_14103,N_13212);
nor UO_1740 (O_1740,N_13202,N_14047);
nor UO_1741 (O_1741,N_13217,N_12205);
or UO_1742 (O_1742,N_14541,N_13157);
and UO_1743 (O_1743,N_14255,N_13225);
or UO_1744 (O_1744,N_14753,N_12165);
and UO_1745 (O_1745,N_13894,N_12097);
nand UO_1746 (O_1746,N_14312,N_14146);
nand UO_1747 (O_1747,N_14663,N_13512);
nor UO_1748 (O_1748,N_14821,N_12698);
or UO_1749 (O_1749,N_12101,N_12207);
or UO_1750 (O_1750,N_14015,N_14592);
and UO_1751 (O_1751,N_14590,N_12137);
nand UO_1752 (O_1752,N_12427,N_12452);
nor UO_1753 (O_1753,N_14780,N_12245);
nand UO_1754 (O_1754,N_13194,N_13941);
or UO_1755 (O_1755,N_14942,N_12351);
and UO_1756 (O_1756,N_14658,N_13624);
and UO_1757 (O_1757,N_13619,N_14462);
or UO_1758 (O_1758,N_13701,N_14716);
xnor UO_1759 (O_1759,N_13573,N_12168);
nor UO_1760 (O_1760,N_13733,N_14778);
or UO_1761 (O_1761,N_13481,N_13277);
and UO_1762 (O_1762,N_12474,N_12584);
nand UO_1763 (O_1763,N_13620,N_14580);
and UO_1764 (O_1764,N_14563,N_14532);
nor UO_1765 (O_1765,N_13469,N_13837);
or UO_1766 (O_1766,N_12049,N_14951);
and UO_1767 (O_1767,N_14972,N_12950);
nand UO_1768 (O_1768,N_12705,N_12183);
nor UO_1769 (O_1769,N_14186,N_13949);
and UO_1770 (O_1770,N_13940,N_13692);
or UO_1771 (O_1771,N_13078,N_12307);
or UO_1772 (O_1772,N_13153,N_14084);
and UO_1773 (O_1773,N_13667,N_12338);
and UO_1774 (O_1774,N_12255,N_14144);
or UO_1775 (O_1775,N_13817,N_14648);
xor UO_1776 (O_1776,N_13701,N_14573);
and UO_1777 (O_1777,N_12547,N_13970);
nand UO_1778 (O_1778,N_12164,N_14810);
nor UO_1779 (O_1779,N_12384,N_13074);
or UO_1780 (O_1780,N_12285,N_13927);
nand UO_1781 (O_1781,N_13935,N_12081);
or UO_1782 (O_1782,N_14818,N_12250);
nor UO_1783 (O_1783,N_14021,N_12729);
or UO_1784 (O_1784,N_13324,N_14038);
and UO_1785 (O_1785,N_14434,N_13165);
xnor UO_1786 (O_1786,N_12379,N_12195);
nand UO_1787 (O_1787,N_12809,N_13988);
nand UO_1788 (O_1788,N_14525,N_12724);
or UO_1789 (O_1789,N_13514,N_14986);
nand UO_1790 (O_1790,N_12467,N_13736);
nand UO_1791 (O_1791,N_12234,N_13469);
nand UO_1792 (O_1792,N_13059,N_14816);
nand UO_1793 (O_1793,N_14008,N_13109);
nor UO_1794 (O_1794,N_12912,N_13608);
nand UO_1795 (O_1795,N_14576,N_12314);
or UO_1796 (O_1796,N_13665,N_14556);
nor UO_1797 (O_1797,N_13855,N_14940);
nand UO_1798 (O_1798,N_12872,N_13839);
or UO_1799 (O_1799,N_12015,N_14775);
nand UO_1800 (O_1800,N_12819,N_12359);
or UO_1801 (O_1801,N_14837,N_14916);
nand UO_1802 (O_1802,N_12194,N_12390);
nand UO_1803 (O_1803,N_12805,N_14476);
nor UO_1804 (O_1804,N_14343,N_12863);
nor UO_1805 (O_1805,N_13465,N_14313);
or UO_1806 (O_1806,N_13439,N_13145);
or UO_1807 (O_1807,N_13935,N_13619);
and UO_1808 (O_1808,N_12148,N_14500);
nand UO_1809 (O_1809,N_12974,N_12012);
or UO_1810 (O_1810,N_13077,N_12360);
or UO_1811 (O_1811,N_12890,N_12303);
nand UO_1812 (O_1812,N_12765,N_14724);
nand UO_1813 (O_1813,N_14111,N_12368);
nor UO_1814 (O_1814,N_14286,N_14895);
nand UO_1815 (O_1815,N_14529,N_13191);
nor UO_1816 (O_1816,N_14188,N_14495);
nor UO_1817 (O_1817,N_13679,N_14785);
and UO_1818 (O_1818,N_14140,N_12862);
nand UO_1819 (O_1819,N_12432,N_14707);
nor UO_1820 (O_1820,N_13332,N_12173);
nor UO_1821 (O_1821,N_14829,N_13294);
and UO_1822 (O_1822,N_12229,N_13892);
or UO_1823 (O_1823,N_14489,N_12022);
nand UO_1824 (O_1824,N_13905,N_14618);
nor UO_1825 (O_1825,N_13351,N_12153);
or UO_1826 (O_1826,N_12503,N_14519);
and UO_1827 (O_1827,N_12340,N_13992);
nor UO_1828 (O_1828,N_12615,N_13923);
nand UO_1829 (O_1829,N_13201,N_12736);
and UO_1830 (O_1830,N_12354,N_12545);
or UO_1831 (O_1831,N_13402,N_13572);
and UO_1832 (O_1832,N_12613,N_14495);
nor UO_1833 (O_1833,N_13023,N_13001);
nor UO_1834 (O_1834,N_12876,N_14216);
nor UO_1835 (O_1835,N_12679,N_13005);
or UO_1836 (O_1836,N_13634,N_13971);
xor UO_1837 (O_1837,N_13729,N_12014);
nor UO_1838 (O_1838,N_13251,N_14741);
nor UO_1839 (O_1839,N_14982,N_13481);
and UO_1840 (O_1840,N_13026,N_12992);
xor UO_1841 (O_1841,N_12852,N_13994);
or UO_1842 (O_1842,N_13669,N_13202);
or UO_1843 (O_1843,N_13715,N_14066);
nor UO_1844 (O_1844,N_12639,N_13358);
or UO_1845 (O_1845,N_13286,N_13184);
nor UO_1846 (O_1846,N_12607,N_13852);
xor UO_1847 (O_1847,N_13475,N_12799);
nand UO_1848 (O_1848,N_14699,N_13381);
nand UO_1849 (O_1849,N_13095,N_13156);
nand UO_1850 (O_1850,N_12014,N_14874);
nor UO_1851 (O_1851,N_14084,N_14559);
nand UO_1852 (O_1852,N_14267,N_13448);
nand UO_1853 (O_1853,N_14286,N_12714);
or UO_1854 (O_1854,N_13155,N_14269);
nor UO_1855 (O_1855,N_14750,N_14483);
nor UO_1856 (O_1856,N_13236,N_12974);
nand UO_1857 (O_1857,N_14691,N_12250);
or UO_1858 (O_1858,N_14303,N_14232);
and UO_1859 (O_1859,N_14284,N_12642);
or UO_1860 (O_1860,N_12446,N_13979);
and UO_1861 (O_1861,N_14887,N_13297);
or UO_1862 (O_1862,N_13996,N_14945);
or UO_1863 (O_1863,N_13871,N_12279);
nor UO_1864 (O_1864,N_12833,N_12122);
and UO_1865 (O_1865,N_13442,N_12209);
nand UO_1866 (O_1866,N_12132,N_12026);
or UO_1867 (O_1867,N_13712,N_14625);
nor UO_1868 (O_1868,N_12515,N_12036);
or UO_1869 (O_1869,N_12598,N_12864);
or UO_1870 (O_1870,N_14087,N_13789);
xor UO_1871 (O_1871,N_13071,N_12995);
or UO_1872 (O_1872,N_12877,N_14273);
nor UO_1873 (O_1873,N_14371,N_13359);
nand UO_1874 (O_1874,N_12837,N_12216);
or UO_1875 (O_1875,N_14041,N_12103);
nand UO_1876 (O_1876,N_13783,N_13522);
nand UO_1877 (O_1877,N_12210,N_14675);
nor UO_1878 (O_1878,N_12561,N_14963);
and UO_1879 (O_1879,N_14991,N_12233);
and UO_1880 (O_1880,N_13286,N_13487);
xor UO_1881 (O_1881,N_13968,N_14356);
or UO_1882 (O_1882,N_12183,N_14409);
and UO_1883 (O_1883,N_13611,N_13145);
nor UO_1884 (O_1884,N_12427,N_13256);
nor UO_1885 (O_1885,N_13419,N_13969);
or UO_1886 (O_1886,N_12318,N_14108);
and UO_1887 (O_1887,N_13786,N_14020);
nor UO_1888 (O_1888,N_14673,N_12668);
or UO_1889 (O_1889,N_14200,N_13988);
or UO_1890 (O_1890,N_14328,N_12440);
nand UO_1891 (O_1891,N_12916,N_13039);
nand UO_1892 (O_1892,N_12549,N_14872);
nor UO_1893 (O_1893,N_13042,N_13038);
or UO_1894 (O_1894,N_14386,N_14469);
nand UO_1895 (O_1895,N_13244,N_14261);
or UO_1896 (O_1896,N_14440,N_13942);
nor UO_1897 (O_1897,N_14590,N_14363);
nand UO_1898 (O_1898,N_14117,N_14544);
and UO_1899 (O_1899,N_13231,N_14358);
nor UO_1900 (O_1900,N_12602,N_13551);
nand UO_1901 (O_1901,N_14393,N_14817);
or UO_1902 (O_1902,N_14562,N_13076);
nand UO_1903 (O_1903,N_13584,N_12720);
nand UO_1904 (O_1904,N_13330,N_13883);
or UO_1905 (O_1905,N_13275,N_12821);
or UO_1906 (O_1906,N_14886,N_12990);
nor UO_1907 (O_1907,N_13502,N_12898);
or UO_1908 (O_1908,N_13790,N_12080);
nand UO_1909 (O_1909,N_14014,N_12255);
or UO_1910 (O_1910,N_13105,N_12607);
or UO_1911 (O_1911,N_12304,N_12142);
and UO_1912 (O_1912,N_12317,N_12748);
nor UO_1913 (O_1913,N_13900,N_13429);
xor UO_1914 (O_1914,N_12932,N_13251);
nand UO_1915 (O_1915,N_13433,N_13440);
nor UO_1916 (O_1916,N_13747,N_13411);
and UO_1917 (O_1917,N_12377,N_14908);
or UO_1918 (O_1918,N_12698,N_13221);
or UO_1919 (O_1919,N_13899,N_14454);
or UO_1920 (O_1920,N_13455,N_14755);
nor UO_1921 (O_1921,N_14677,N_12631);
and UO_1922 (O_1922,N_13532,N_14400);
nand UO_1923 (O_1923,N_12084,N_13944);
or UO_1924 (O_1924,N_12769,N_12451);
or UO_1925 (O_1925,N_12503,N_13416);
and UO_1926 (O_1926,N_14709,N_13268);
or UO_1927 (O_1927,N_14582,N_12559);
and UO_1928 (O_1928,N_13712,N_14587);
nand UO_1929 (O_1929,N_14574,N_12322);
or UO_1930 (O_1930,N_14861,N_14635);
nand UO_1931 (O_1931,N_14840,N_13968);
nor UO_1932 (O_1932,N_13665,N_13915);
nor UO_1933 (O_1933,N_14631,N_14109);
xor UO_1934 (O_1934,N_13647,N_13925);
nand UO_1935 (O_1935,N_12524,N_13491);
nor UO_1936 (O_1936,N_12992,N_13606);
nor UO_1937 (O_1937,N_13452,N_13228);
nor UO_1938 (O_1938,N_12417,N_14528);
nor UO_1939 (O_1939,N_14765,N_12690);
nor UO_1940 (O_1940,N_13050,N_14671);
or UO_1941 (O_1941,N_13555,N_14561);
nor UO_1942 (O_1942,N_14091,N_12505);
nand UO_1943 (O_1943,N_14110,N_14962);
xnor UO_1944 (O_1944,N_13647,N_12544);
or UO_1945 (O_1945,N_14637,N_14800);
and UO_1946 (O_1946,N_12355,N_13679);
nor UO_1947 (O_1947,N_14774,N_12930);
nand UO_1948 (O_1948,N_14415,N_14120);
nor UO_1949 (O_1949,N_12029,N_13981);
and UO_1950 (O_1950,N_12619,N_14142);
nand UO_1951 (O_1951,N_12091,N_13633);
nand UO_1952 (O_1952,N_14774,N_14390);
nand UO_1953 (O_1953,N_14154,N_13655);
nand UO_1954 (O_1954,N_13851,N_13118);
nand UO_1955 (O_1955,N_13648,N_12678);
nand UO_1956 (O_1956,N_14751,N_14413);
nor UO_1957 (O_1957,N_13699,N_14933);
and UO_1958 (O_1958,N_14146,N_14608);
nand UO_1959 (O_1959,N_13512,N_12759);
nand UO_1960 (O_1960,N_13778,N_14357);
and UO_1961 (O_1961,N_14551,N_12658);
nand UO_1962 (O_1962,N_12798,N_14884);
nand UO_1963 (O_1963,N_13945,N_14115);
or UO_1964 (O_1964,N_12566,N_14411);
nand UO_1965 (O_1965,N_14912,N_14122);
or UO_1966 (O_1966,N_13559,N_13988);
nor UO_1967 (O_1967,N_14647,N_12759);
nor UO_1968 (O_1968,N_13559,N_14792);
nor UO_1969 (O_1969,N_13700,N_12277);
nand UO_1970 (O_1970,N_12124,N_13071);
nor UO_1971 (O_1971,N_14377,N_14946);
nor UO_1972 (O_1972,N_14320,N_14127);
and UO_1973 (O_1973,N_12958,N_12560);
xnor UO_1974 (O_1974,N_13123,N_12724);
nand UO_1975 (O_1975,N_14070,N_12074);
nand UO_1976 (O_1976,N_14648,N_14616);
nor UO_1977 (O_1977,N_14962,N_12149);
or UO_1978 (O_1978,N_14454,N_13309);
nor UO_1979 (O_1979,N_14201,N_14523);
or UO_1980 (O_1980,N_14340,N_14689);
nor UO_1981 (O_1981,N_12914,N_13573);
and UO_1982 (O_1982,N_14257,N_14594);
or UO_1983 (O_1983,N_13317,N_12444);
nor UO_1984 (O_1984,N_13013,N_13829);
and UO_1985 (O_1985,N_14880,N_13724);
xor UO_1986 (O_1986,N_14732,N_12584);
nand UO_1987 (O_1987,N_13338,N_13790);
or UO_1988 (O_1988,N_14170,N_13444);
or UO_1989 (O_1989,N_12834,N_12389);
nor UO_1990 (O_1990,N_13988,N_13162);
nor UO_1991 (O_1991,N_14571,N_14564);
nand UO_1992 (O_1992,N_12823,N_13422);
and UO_1993 (O_1993,N_13864,N_13343);
and UO_1994 (O_1994,N_14278,N_12634);
or UO_1995 (O_1995,N_14851,N_13719);
and UO_1996 (O_1996,N_12589,N_14752);
nand UO_1997 (O_1997,N_12717,N_13503);
nor UO_1998 (O_1998,N_14991,N_12858);
or UO_1999 (O_1999,N_14416,N_14519);
endmodule