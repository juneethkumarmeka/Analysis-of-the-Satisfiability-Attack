module basic_1000_10000_1500_100_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_236,In_821);
xnor U1 (N_1,In_329,In_13);
and U2 (N_2,In_356,In_415);
nand U3 (N_3,In_85,In_538);
or U4 (N_4,In_286,In_611);
nor U5 (N_5,In_498,In_327);
nor U6 (N_6,In_715,In_685);
and U7 (N_7,In_517,In_207);
and U8 (N_8,In_271,In_185);
and U9 (N_9,In_805,In_164);
and U10 (N_10,In_942,In_229);
and U11 (N_11,In_870,In_167);
and U12 (N_12,In_874,In_144);
nand U13 (N_13,In_350,In_456);
xor U14 (N_14,In_422,In_769);
and U15 (N_15,In_375,In_804);
nor U16 (N_16,In_206,In_364);
nor U17 (N_17,In_400,In_59);
or U18 (N_18,In_783,In_664);
nor U19 (N_19,In_270,In_312);
nand U20 (N_20,In_103,In_79);
or U21 (N_21,In_503,In_153);
nor U22 (N_22,In_829,In_626);
xnor U23 (N_23,In_396,In_40);
xnor U24 (N_24,In_293,In_116);
or U25 (N_25,In_418,In_20);
and U26 (N_26,In_162,In_780);
nor U27 (N_27,In_64,In_537);
or U28 (N_28,In_986,In_864);
nand U29 (N_29,In_359,In_738);
nand U30 (N_30,In_845,In_266);
nand U31 (N_31,In_392,In_512);
nor U32 (N_32,In_652,In_377);
xor U33 (N_33,In_226,In_402);
nand U34 (N_34,In_490,In_281);
nand U35 (N_35,In_478,In_467);
xor U36 (N_36,In_315,In_260);
xor U37 (N_37,In_218,In_848);
xnor U38 (N_38,In_925,In_311);
and U39 (N_39,In_758,In_27);
and U40 (N_40,In_307,In_360);
nor U41 (N_41,In_952,In_799);
xor U42 (N_42,In_58,In_775);
and U43 (N_43,In_972,In_343);
and U44 (N_44,In_161,In_555);
nand U45 (N_45,In_105,In_599);
nand U46 (N_46,In_106,In_460);
xor U47 (N_47,In_317,In_10);
nor U48 (N_48,In_981,In_3);
xor U49 (N_49,In_133,In_568);
or U50 (N_50,In_160,In_628);
xnor U51 (N_51,In_548,In_589);
or U52 (N_52,In_171,In_722);
and U53 (N_53,In_872,In_806);
xnor U54 (N_54,In_527,In_752);
and U55 (N_55,In_917,In_618);
xnor U56 (N_56,In_62,In_647);
xnor U57 (N_57,In_807,In_929);
nor U58 (N_58,In_259,In_693);
and U59 (N_59,In_533,In_150);
or U60 (N_60,In_609,In_563);
and U61 (N_61,In_119,In_697);
nand U62 (N_62,In_766,In_48);
xor U63 (N_63,In_253,In_221);
and U64 (N_64,In_849,In_531);
xnor U65 (N_65,In_959,In_802);
or U66 (N_66,In_211,In_678);
xnor U67 (N_67,In_889,In_84);
xnor U68 (N_68,In_567,In_607);
xnor U69 (N_69,In_523,In_267);
xor U70 (N_70,In_876,In_55);
nor U71 (N_71,In_910,In_616);
or U72 (N_72,In_19,In_112);
and U73 (N_73,In_737,In_690);
xor U74 (N_74,In_262,In_99);
nand U75 (N_75,In_574,In_322);
and U76 (N_76,In_152,In_433);
nor U77 (N_77,In_502,In_970);
nand U78 (N_78,In_443,In_447);
and U79 (N_79,In_827,In_214);
nand U80 (N_80,In_473,In_645);
nor U81 (N_81,In_554,In_485);
or U82 (N_82,In_923,In_822);
and U83 (N_83,In_406,In_543);
or U84 (N_84,In_50,In_801);
and U85 (N_85,In_767,In_118);
xnor U86 (N_86,In_840,In_908);
nand U87 (N_87,In_898,In_384);
or U88 (N_88,In_299,In_386);
nand U89 (N_89,In_366,In_71);
nand U90 (N_90,In_276,In_409);
or U91 (N_91,In_593,In_838);
xnor U92 (N_92,In_324,In_508);
nor U93 (N_93,In_689,In_184);
nand U94 (N_94,In_9,In_622);
nor U95 (N_95,In_136,In_17);
or U96 (N_96,In_306,In_950);
and U97 (N_97,In_8,In_565);
and U98 (N_98,In_818,In_886);
nand U99 (N_99,In_35,In_643);
nand U100 (N_100,In_420,In_181);
or U101 (N_101,In_137,In_368);
nor U102 (N_102,N_92,N_13);
and U103 (N_103,In_638,In_608);
nand U104 (N_104,In_397,In_149);
nor U105 (N_105,In_586,In_798);
nand U106 (N_106,In_916,In_345);
nor U107 (N_107,In_896,In_82);
xnor U108 (N_108,In_782,In_138);
nor U109 (N_109,In_158,N_86);
or U110 (N_110,In_835,In_23);
and U111 (N_111,In_398,In_772);
nor U112 (N_112,In_269,In_587);
nand U113 (N_113,In_698,In_56);
and U114 (N_114,N_62,In_865);
and U115 (N_115,In_123,In_468);
xnor U116 (N_116,In_768,In_279);
and U117 (N_117,In_474,N_36);
nor U118 (N_118,In_948,N_46);
and U119 (N_119,In_483,In_985);
and U120 (N_120,In_884,In_475);
xor U121 (N_121,In_790,In_755);
nand U122 (N_122,In_900,In_337);
xnor U123 (N_123,In_14,In_53);
xnor U124 (N_124,In_330,In_815);
nand U125 (N_125,In_931,In_197);
nand U126 (N_126,In_18,In_499);
and U127 (N_127,In_63,In_993);
nand U128 (N_128,In_189,In_951);
nand U129 (N_129,N_72,In_895);
xnor U130 (N_130,In_182,In_724);
and U131 (N_131,In_296,In_282);
xnor U132 (N_132,In_705,In_551);
and U133 (N_133,In_450,In_342);
nor U134 (N_134,In_151,In_630);
and U135 (N_135,In_225,In_275);
xor U136 (N_136,In_476,In_719);
nand U137 (N_137,In_393,In_428);
nor U138 (N_138,In_170,In_379);
nand U139 (N_139,In_712,In_223);
nor U140 (N_140,In_67,In_547);
xnor U141 (N_141,In_290,In_122);
or U142 (N_142,In_853,In_542);
nand U143 (N_143,In_388,In_370);
and U144 (N_144,In_836,In_613);
nor U145 (N_145,In_961,In_410);
nor U146 (N_146,In_76,In_159);
nand U147 (N_147,In_156,In_661);
nor U148 (N_148,In_172,In_187);
xnor U149 (N_149,In_990,In_803);
nor U150 (N_150,In_129,In_493);
or U151 (N_151,N_84,In_124);
xor U152 (N_152,In_100,In_629);
nor U153 (N_153,N_77,In_938);
xor U154 (N_154,In_102,N_50);
nand U155 (N_155,In_749,In_614);
or U156 (N_156,In_301,In_4);
or U157 (N_157,In_524,In_36);
or U158 (N_158,In_696,In_978);
xor U159 (N_159,In_559,In_659);
xnor U160 (N_160,In_148,In_877);
xnor U161 (N_161,In_11,In_581);
and U162 (N_162,In_539,N_39);
and U163 (N_163,In_54,In_871);
nor U164 (N_164,In_25,In_703);
xor U165 (N_165,In_510,N_11);
nand U166 (N_166,In_486,In_556);
xnor U167 (N_167,N_45,In_319);
or U168 (N_168,In_175,In_147);
nand U169 (N_169,In_640,In_96);
or U170 (N_170,In_432,In_511);
nor U171 (N_171,In_302,In_209);
and U172 (N_172,In_280,In_395);
nor U173 (N_173,N_75,In_882);
nand U174 (N_174,In_174,In_245);
nor U175 (N_175,N_26,In_419);
and U176 (N_176,In_577,In_146);
nor U177 (N_177,In_177,In_520);
and U178 (N_178,In_930,In_892);
nand U179 (N_179,In_940,In_387);
nand U180 (N_180,In_438,In_120);
and U181 (N_181,In_466,In_842);
xnor U182 (N_182,N_16,In_489);
and U183 (N_183,In_331,In_869);
nand U184 (N_184,In_190,In_653);
or U185 (N_185,In_166,In_810);
nor U186 (N_186,In_74,In_371);
nand U187 (N_187,N_93,N_17);
and U188 (N_188,In_561,In_335);
and U189 (N_189,In_268,In_505);
and U190 (N_190,In_374,In_451);
nor U191 (N_191,N_14,N_9);
or U192 (N_192,In_132,In_204);
or U193 (N_193,In_352,In_816);
xnor U194 (N_194,In_414,In_636);
or U195 (N_195,In_716,In_394);
xor U196 (N_196,In_742,In_721);
nor U197 (N_197,In_602,In_179);
and U198 (N_198,In_771,In_662);
and U199 (N_199,In_580,In_788);
nand U200 (N_200,In_213,In_744);
xnor U201 (N_201,N_168,In_700);
xor U202 (N_202,N_181,In_30);
xnor U203 (N_203,In_686,N_174);
xor U204 (N_204,N_189,In_339);
nand U205 (N_205,N_167,In_348);
xnor U206 (N_206,N_135,N_192);
nand U207 (N_207,In_710,In_544);
and U208 (N_208,N_111,N_106);
xnor U209 (N_209,In_726,In_252);
and U210 (N_210,In_462,In_287);
and U211 (N_211,In_528,N_137);
nor U212 (N_212,In_656,In_671);
nor U213 (N_213,In_93,In_596);
or U214 (N_214,In_308,In_362);
nor U215 (N_215,In_911,In_817);
nand U216 (N_216,In_968,N_198);
or U217 (N_217,N_34,In_789);
nor U218 (N_218,In_960,In_458);
and U219 (N_219,N_128,In_429);
nor U220 (N_220,N_43,In_606);
nand U221 (N_221,In_761,In_902);
or U222 (N_222,N_37,In_828);
and U223 (N_223,In_261,In_695);
nor U224 (N_224,In_453,In_918);
xnor U225 (N_225,N_78,In_479);
nand U226 (N_226,In_868,In_417);
and U227 (N_227,In_127,In_663);
nor U228 (N_228,In_249,In_504);
nand U229 (N_229,N_79,N_186);
xnor U230 (N_230,In_756,In_101);
nor U231 (N_231,In_991,N_47);
or U232 (N_232,In_617,In_78);
and U233 (N_233,N_175,In_883);
and U234 (N_234,N_147,In_651);
or U235 (N_235,In_341,In_141);
and U236 (N_236,In_196,N_6);
or U237 (N_237,In_436,In_532);
xnor U238 (N_238,In_347,In_944);
nor U239 (N_239,In_47,In_774);
and U240 (N_240,In_186,In_957);
nor U241 (N_241,In_830,In_391);
and U242 (N_242,In_655,N_146);
nor U243 (N_243,In_70,In_846);
or U244 (N_244,In_294,In_192);
or U245 (N_245,In_292,In_578);
nand U246 (N_246,In_757,In_157);
or U247 (N_247,In_413,In_979);
nor U248 (N_248,N_41,N_171);
nor U249 (N_249,In_22,In_107);
or U250 (N_250,In_740,In_612);
and U251 (N_251,In_21,In_935);
and U252 (N_252,In_878,N_159);
nand U253 (N_253,In_759,In_24);
nand U254 (N_254,N_20,In_632);
xor U255 (N_255,In_831,In_346);
xnor U256 (N_256,In_235,In_255);
nand U257 (N_257,N_114,N_53);
xor U258 (N_258,In_987,In_472);
nor U259 (N_259,N_191,In_316);
nand U260 (N_260,In_811,In_604);
and U261 (N_261,In_90,In_201);
and U262 (N_262,In_125,In_954);
or U263 (N_263,In_355,N_5);
nor U264 (N_264,In_674,In_692);
nand U265 (N_265,In_369,In_191);
or U266 (N_266,In_927,In_378);
xor U267 (N_267,N_38,In_873);
and U268 (N_268,In_477,In_974);
and U269 (N_269,In_668,In_284);
or U270 (N_270,In_176,N_81);
and U271 (N_271,In_649,In_385);
xor U272 (N_272,In_560,In_318);
xnor U273 (N_273,In_143,In_16);
nor U274 (N_274,In_754,In_155);
xnor U275 (N_275,In_603,In_449);
or U276 (N_276,N_153,In_509);
nor U277 (N_277,In_309,In_257);
or U278 (N_278,N_185,In_901);
nand U279 (N_279,In_38,In_733);
and U280 (N_280,In_401,In_855);
or U281 (N_281,In_860,In_130);
or U282 (N_282,In_247,N_113);
nand U283 (N_283,In_183,In_224);
nor U284 (N_284,In_964,In_424);
and U285 (N_285,In_820,In_718);
and U286 (N_286,In_195,N_118);
xnor U287 (N_287,In_46,In_169);
or U288 (N_288,N_49,In_494);
nand U289 (N_289,N_109,In_514);
and U290 (N_290,In_792,In_441);
nor U291 (N_291,N_193,In_328);
xor U292 (N_292,In_234,N_58);
and U293 (N_293,In_670,In_562);
nand U294 (N_294,N_42,In_875);
and U295 (N_295,In_34,In_357);
nor U296 (N_296,In_248,In_305);
xor U297 (N_297,In_228,N_184);
and U298 (N_298,In_363,In_905);
and U299 (N_299,In_937,In_826);
nand U300 (N_300,N_95,In_939);
or U301 (N_301,In_26,In_781);
nor U302 (N_302,In_646,In_484);
nand U303 (N_303,In_77,In_427);
nor U304 (N_304,N_233,In_814);
nand U305 (N_305,In_241,In_277);
nor U306 (N_306,In_861,In_32);
and U307 (N_307,N_110,In_773);
nor U308 (N_308,In_44,In_51);
nand U309 (N_309,In_576,N_12);
nor U310 (N_310,In_880,In_361);
xnor U311 (N_311,In_941,In_654);
xnor U312 (N_312,In_857,In_976);
nor U313 (N_313,N_33,In_500);
or U314 (N_314,In_212,In_240);
or U315 (N_315,In_126,In_1);
or U316 (N_316,In_140,In_966);
or U317 (N_317,In_208,In_445);
or U318 (N_318,In_549,In_854);
and U319 (N_319,In_859,N_166);
xor U320 (N_320,In_442,N_277);
and U321 (N_321,N_25,N_120);
or U322 (N_322,In_83,In_725);
nor U323 (N_323,N_226,In_566);
xor U324 (N_324,In_809,In_862);
or U325 (N_325,In_334,N_297);
nor U326 (N_326,N_276,In_732);
xnor U327 (N_327,In_367,In_230);
and U328 (N_328,N_152,In_682);
nand U329 (N_329,N_270,In_627);
or U330 (N_330,In_243,N_157);
and U331 (N_331,In_457,N_23);
xnor U332 (N_332,N_48,In_743);
and U333 (N_333,N_31,In_634);
xnor U334 (N_334,In_897,In_791);
nor U335 (N_335,In_463,In_597);
or U336 (N_336,In_582,N_99);
nand U337 (N_337,In_75,In_326);
and U338 (N_338,In_45,N_150);
nand U339 (N_339,In_992,In_39);
xor U340 (N_340,In_701,N_125);
nor U341 (N_341,In_676,In_426);
xor U342 (N_342,N_288,In_12);
and U343 (N_343,N_71,In_748);
nand U344 (N_344,N_66,N_57);
or U345 (N_345,In_142,N_249);
nor U346 (N_346,In_833,N_214);
or U347 (N_347,In_323,In_601);
xor U348 (N_348,In_336,N_104);
and U349 (N_349,N_201,In_982);
and U350 (N_350,In_303,In_736);
nor U351 (N_351,In_265,N_236);
or U352 (N_352,In_88,N_63);
nor U353 (N_353,In_879,In_104);
and U354 (N_354,N_68,N_40);
or U355 (N_355,In_111,In_52);
nand U356 (N_356,N_67,N_80);
or U357 (N_357,In_746,In_666);
and U358 (N_358,In_794,In_920);
xor U359 (N_359,In_907,In_321);
nor U360 (N_360,In_975,N_211);
xnor U361 (N_361,N_140,In_254);
nor U362 (N_362,N_69,N_7);
nor U363 (N_363,In_852,In_863);
xor U364 (N_364,In_60,In_965);
xor U365 (N_365,N_292,N_161);
nor U366 (N_366,N_238,In_633);
nand U367 (N_367,In_837,In_541);
nand U368 (N_368,N_30,In_605);
nand U369 (N_369,In_765,In_258);
xnor U370 (N_370,N_232,N_101);
nand U371 (N_371,In_376,N_209);
and U372 (N_372,In_238,In_890);
nand U373 (N_373,In_439,N_172);
or U374 (N_374,In_304,In_620);
xnor U375 (N_375,N_246,In_999);
xor U376 (N_376,In_635,In_344);
nor U377 (N_377,In_711,In_550);
nand U378 (N_378,In_980,In_988);
nor U379 (N_379,In_314,In_325);
and U380 (N_380,N_182,N_266);
nand U381 (N_381,In_29,In_958);
nor U382 (N_382,In_465,In_117);
nand U383 (N_383,In_847,In_914);
and U384 (N_384,In_501,In_516);
nor U385 (N_385,In_683,In_909);
xor U386 (N_386,In_219,In_913);
nor U387 (N_387,N_218,N_289);
and U388 (N_388,In_272,In_495);
xnor U389 (N_389,N_247,In_953);
xnor U390 (N_390,N_261,In_313);
xor U391 (N_391,In_232,In_65);
nor U392 (N_392,N_235,In_730);
nor U393 (N_393,In_89,In_471);
xor U394 (N_394,In_924,In_320);
nor U395 (N_395,N_196,In_881);
and U396 (N_396,In_785,N_83);
nand U397 (N_397,N_87,N_284);
nor U398 (N_398,In_291,N_165);
xor U399 (N_399,N_177,In_506);
xnor U400 (N_400,N_307,In_57);
xnor U401 (N_401,In_131,In_519);
nor U402 (N_402,In_932,In_242);
nor U403 (N_403,In_273,In_669);
xor U404 (N_404,N_205,N_132);
nand U405 (N_405,In_354,N_204);
or U406 (N_406,N_367,N_18);
and U407 (N_407,In_893,In_694);
and U408 (N_408,In_778,In_592);
and U409 (N_409,In_677,In_899);
or U410 (N_410,In_750,In_996);
xor U411 (N_411,In_572,N_350);
xor U412 (N_412,In_198,In_298);
nor U413 (N_413,In_380,N_241);
xnor U414 (N_414,In_997,In_588);
and U415 (N_415,N_117,N_283);
nand U416 (N_416,In_154,N_351);
nand U417 (N_417,N_100,N_316);
xnor U418 (N_418,N_24,In_403);
and U419 (N_419,N_74,N_298);
nor U420 (N_420,N_317,N_88);
xnor U421 (N_421,N_134,In_239);
and U422 (N_422,N_206,N_338);
nor U423 (N_423,In_358,In_787);
nor U424 (N_424,N_334,N_59);
xor U425 (N_425,In_558,N_286);
nand U426 (N_426,In_973,In_188);
or U427 (N_427,In_844,In_885);
or U428 (N_428,N_390,In_658);
and U429 (N_429,In_797,N_269);
xor U430 (N_430,N_333,N_279);
xnor U431 (N_431,In_95,N_61);
or U432 (N_432,In_283,In_145);
nand U433 (N_433,N_239,N_155);
or U434 (N_434,N_178,In_679);
nor U435 (N_435,N_136,In_675);
xor U436 (N_436,N_399,In_583);
nand U437 (N_437,N_341,In_297);
nor U438 (N_438,N_313,N_151);
or U439 (N_439,N_223,In_28);
and U440 (N_440,In_856,N_240);
nand U441 (N_441,N_127,N_309);
or U442 (N_442,In_430,N_319);
nand U443 (N_443,In_776,N_396);
nand U444 (N_444,In_673,N_143);
nor U445 (N_445,In_753,In_793);
and U446 (N_446,N_144,In_621);
and U447 (N_447,In_637,N_392);
xor U448 (N_448,In_699,In_382);
xnor U449 (N_449,In_530,In_557);
xor U450 (N_450,N_354,In_405);
xor U451 (N_451,N_295,N_44);
nand U452 (N_452,In_42,In_200);
xnor U453 (N_453,In_452,N_229);
nand U454 (N_454,In_513,N_332);
or U455 (N_455,In_850,N_360);
xnor U456 (N_456,In_194,N_262);
nor U457 (N_457,In_912,In_251);
or U458 (N_458,In_745,N_123);
and U459 (N_459,In_569,In_529);
xor U460 (N_460,In_631,In_165);
nor U461 (N_461,In_824,N_369);
nand U462 (N_462,N_325,In_421);
xor U463 (N_463,N_320,In_446);
nand U464 (N_464,In_222,N_56);
nand U465 (N_465,In_278,N_265);
xnor U466 (N_466,N_52,N_170);
nor U467 (N_467,In_764,N_112);
nor U468 (N_468,N_387,N_373);
xor U469 (N_469,In_440,N_398);
nand U470 (N_470,N_271,N_115);
or U471 (N_471,In_922,N_345);
or U472 (N_472,N_180,N_329);
xor U473 (N_473,In_665,N_199);
or U474 (N_474,In_416,N_89);
and U475 (N_475,In_15,N_324);
or U476 (N_476,N_234,N_363);
or U477 (N_477,N_382,In_739);
and U478 (N_478,In_625,N_336);
or U479 (N_479,In_33,In_41);
and U480 (N_480,N_176,N_15);
nand U481 (N_481,N_179,In_199);
and U482 (N_482,N_94,N_195);
nor U483 (N_483,N_308,N_393);
nand U484 (N_484,In_720,In_546);
nor U485 (N_485,N_0,In_573);
xor U486 (N_486,N_251,N_85);
or U487 (N_487,N_359,In_867);
xnor U488 (N_488,In_115,N_255);
nor U489 (N_489,In_926,In_969);
xor U490 (N_490,N_312,In_87);
nand U491 (N_491,N_344,N_156);
or U492 (N_492,N_340,N_342);
nand U493 (N_493,N_158,N_349);
or U494 (N_494,N_194,N_323);
nand U495 (N_495,In_786,In_365);
xnor U496 (N_496,N_372,N_303);
xor U497 (N_497,In_437,In_956);
or U498 (N_498,In_984,In_947);
xor U499 (N_499,N_35,N_357);
xor U500 (N_500,N_365,In_688);
or U501 (N_501,N_202,In_600);
xor U502 (N_502,N_141,N_448);
nor U503 (N_503,N_389,N_221);
nor U504 (N_504,In_372,In_709);
and U505 (N_505,In_591,N_210);
nand U506 (N_506,N_272,In_98);
xor U507 (N_507,In_714,N_267);
and U508 (N_508,In_747,In_215);
xnor U509 (N_509,In_338,N_483);
nand U510 (N_510,In_73,N_21);
xor U511 (N_511,N_302,N_374);
or U512 (N_512,In_946,In_610);
nand U513 (N_513,In_300,N_429);
or U514 (N_514,In_295,N_318);
nor U515 (N_515,N_133,N_426);
and U516 (N_516,In_431,N_339);
or U517 (N_517,N_274,N_479);
and U518 (N_518,N_413,In_49);
nand U519 (N_519,In_921,N_290);
xor U520 (N_520,N_215,In_459);
or U521 (N_521,In_515,N_328);
nor U522 (N_522,In_285,N_105);
nor U523 (N_523,N_60,In_680);
and U524 (N_524,In_760,N_462);
xnor U525 (N_525,N_273,In_858);
nor U526 (N_526,N_465,In_72);
xor U527 (N_527,N_242,N_348);
and U528 (N_528,In_841,N_404);
xor U529 (N_529,In_480,In_728);
or U530 (N_530,In_507,In_707);
nor U531 (N_531,N_446,In_274);
xnor U532 (N_532,In_288,In_983);
nand U533 (N_533,N_162,N_436);
nand U534 (N_534,N_482,N_478);
nor U535 (N_535,In_735,N_256);
nor U536 (N_536,N_213,In_998);
nand U537 (N_537,In_383,In_43);
nand U538 (N_538,N_441,In_891);
xnor U539 (N_539,In_575,N_403);
or U540 (N_540,N_439,In_231);
nand U541 (N_541,In_644,N_268);
and U542 (N_542,N_327,N_119);
nor U543 (N_543,N_200,N_492);
nand U544 (N_544,N_103,In_193);
nor U545 (N_545,N_169,N_461);
nand U546 (N_546,N_391,In_619);
nand U547 (N_547,In_340,In_37);
nand U548 (N_548,N_469,In_639);
or U549 (N_549,N_2,In_763);
or U550 (N_550,N_455,N_411);
and U551 (N_551,N_484,N_454);
and U552 (N_552,N_460,In_933);
xnor U553 (N_553,In_971,N_243);
nor U554 (N_554,N_386,N_430);
and U555 (N_555,In_995,In_110);
or U556 (N_556,N_414,In_681);
nor U557 (N_557,In_487,N_107);
or U558 (N_558,In_784,N_22);
nand U559 (N_559,In_220,In_80);
or U560 (N_560,N_96,N_432);
nand U561 (N_561,In_904,In_425);
nor U562 (N_562,N_420,N_129);
xor U563 (N_563,In_482,N_90);
xnor U564 (N_564,N_122,In_570);
or U565 (N_565,In_173,In_843);
xor U566 (N_566,In_641,N_331);
nor U567 (N_567,N_287,N_263);
nor U568 (N_568,In_713,N_124);
nor U569 (N_569,N_379,In_660);
nor U570 (N_570,N_400,N_438);
nor U571 (N_571,N_138,In_351);
xor U572 (N_572,N_378,In_642);
nand U573 (N_573,N_10,In_203);
xnor U574 (N_574,In_919,In_246);
xnor U575 (N_575,In_564,In_594);
nand U576 (N_576,In_977,N_346);
xnor U577 (N_577,N_91,In_615);
nand U578 (N_578,In_66,N_294);
nor U579 (N_579,N_160,N_375);
nand U580 (N_580,N_65,N_183);
xor U581 (N_581,In_461,N_330);
xnor U582 (N_582,N_417,In_134);
nor U583 (N_583,In_411,In_444);
nand U584 (N_584,In_455,N_1);
or U585 (N_585,N_364,In_202);
nand U586 (N_586,In_454,N_437);
or U587 (N_587,N_275,In_894);
or U588 (N_588,In_256,N_447);
nand U589 (N_589,In_751,N_402);
nor U590 (N_590,N_370,N_139);
and U591 (N_591,N_498,In_887);
and U592 (N_592,In_552,N_416);
nor U593 (N_593,N_384,N_190);
nand U594 (N_594,N_8,In_404);
nand U595 (N_595,N_347,In_381);
nand U596 (N_596,In_813,N_377);
nor U597 (N_597,N_335,In_332);
xnor U598 (N_598,N_231,N_296);
xnor U599 (N_599,N_278,N_409);
xnor U600 (N_600,N_493,N_575);
nand U601 (N_601,In_915,N_587);
nand U602 (N_602,In_623,In_244);
nor U603 (N_603,N_578,In_657);
nand U604 (N_604,N_457,N_544);
nand U605 (N_605,N_584,N_579);
xnor U606 (N_606,In_31,In_349);
or U607 (N_607,In_139,N_442);
nand U608 (N_608,N_187,N_518);
nor U609 (N_609,In_967,N_428);
nor U610 (N_610,N_521,N_486);
nand U611 (N_611,In_109,N_451);
nor U612 (N_612,N_27,In_163);
or U613 (N_613,N_252,N_154);
nand U614 (N_614,In_464,N_553);
nand U615 (N_615,In_373,N_300);
and U616 (N_616,In_69,N_467);
and U617 (N_617,In_553,In_708);
or U618 (N_618,N_488,In_571);
nor U619 (N_619,In_989,In_525);
xor U620 (N_620,In_779,N_590);
and U621 (N_621,In_702,In_492);
nand U622 (N_622,N_496,N_550);
nor U623 (N_623,In_86,N_130);
nand U624 (N_624,N_97,In_706);
xor U625 (N_625,N_499,N_554);
nor U626 (N_626,In_590,N_538);
and U627 (N_627,N_456,N_376);
xnor U628 (N_628,N_519,In_536);
xor U629 (N_629,N_371,In_389);
or U630 (N_630,N_539,N_507);
or U631 (N_631,In_2,N_32);
or U632 (N_632,N_452,N_285);
or U633 (N_633,N_401,N_491);
or U634 (N_634,N_573,In_834);
nor U635 (N_635,In_777,In_81);
nor U636 (N_636,N_314,N_116);
xnor U637 (N_637,N_572,N_163);
nor U638 (N_638,N_212,In_94);
nor U639 (N_639,N_3,N_470);
nand U640 (N_640,N_562,N_450);
nor U641 (N_641,N_54,In_399);
xnor U642 (N_642,N_512,In_97);
and U643 (N_643,In_928,In_650);
or U644 (N_644,N_583,N_108);
and U645 (N_645,In_825,N_245);
nand U646 (N_646,In_121,In_545);
nand U647 (N_647,N_299,N_406);
nand U648 (N_648,In_691,N_528);
nor U649 (N_649,N_547,In_135);
nand U650 (N_650,In_61,N_495);
and U651 (N_651,N_595,In_819);
nand U652 (N_652,In_7,In_949);
xnor U653 (N_653,N_381,In_481);
and U654 (N_654,N_321,N_412);
nand U655 (N_655,In_113,N_506);
or U656 (N_656,In_734,N_366);
nor U657 (N_657,In_210,In_648);
or U658 (N_658,In_68,N_407);
nor U659 (N_659,N_585,In_390);
or U660 (N_660,N_570,In_526);
and U661 (N_661,In_448,In_92);
nor U662 (N_662,N_475,N_237);
and U663 (N_663,N_565,In_180);
xor U664 (N_664,N_281,N_217);
or U665 (N_665,N_468,In_672);
nor U666 (N_666,N_310,N_551);
or U667 (N_667,In_227,In_497);
nand U668 (N_668,N_569,N_592);
and U669 (N_669,N_421,N_533);
and U670 (N_670,N_197,N_435);
and U671 (N_671,N_541,N_586);
or U672 (N_672,N_301,N_520);
xor U673 (N_673,In_488,N_394);
nand U674 (N_674,In_795,In_667);
and U675 (N_675,N_427,In_5);
nand U676 (N_676,N_545,N_561);
or U677 (N_677,N_445,In_906);
and U678 (N_678,N_126,N_556);
nand U679 (N_679,N_424,N_216);
nand U680 (N_680,In_108,N_443);
or U681 (N_681,N_304,N_524);
nand U682 (N_682,N_244,In_114);
nand U683 (N_683,N_593,N_222);
xor U684 (N_684,N_380,In_470);
and U685 (N_685,In_540,N_361);
or U686 (N_686,N_322,N_315);
nand U687 (N_687,N_28,N_4);
and U688 (N_688,N_574,In_823);
or U689 (N_689,N_531,N_464);
xor U690 (N_690,N_415,N_326);
xnor U691 (N_691,In_808,In_333);
and U692 (N_692,N_343,N_358);
or U693 (N_693,N_282,N_431);
and U694 (N_694,N_537,N_29);
xnor U695 (N_695,N_337,N_503);
xor U696 (N_696,In_584,In_800);
nor U697 (N_697,N_425,N_385);
nand U698 (N_698,N_422,N_581);
nor U699 (N_699,In_469,In_168);
nand U700 (N_700,N_480,N_440);
or U701 (N_701,In_741,N_667);
nor U702 (N_702,N_397,N_557);
xor U703 (N_703,N_641,In_518);
nor U704 (N_704,N_674,N_250);
and U705 (N_705,In_178,N_500);
nor U706 (N_706,N_352,N_149);
xor U707 (N_707,N_527,N_559);
xor U708 (N_708,N_73,In_289);
nor U709 (N_709,N_611,N_614);
and U710 (N_710,In_412,In_729);
nand U711 (N_711,In_263,N_259);
nor U712 (N_712,N_487,N_98);
xor U713 (N_713,N_355,In_535);
and U714 (N_714,N_501,N_410);
and U715 (N_715,N_449,N_145);
xor U716 (N_716,N_254,In_936);
nor U717 (N_717,In_687,N_549);
nand U718 (N_718,N_697,N_616);
nor U719 (N_719,N_603,N_591);
and U720 (N_720,N_645,N_504);
or U721 (N_721,In_237,N_532);
and U722 (N_722,N_517,N_636);
and U723 (N_723,N_693,N_459);
nor U724 (N_724,In_310,N_694);
nor U725 (N_725,N_672,In_496);
nand U726 (N_726,N_513,N_660);
nand U727 (N_727,N_598,N_423);
or U728 (N_728,In_962,N_264);
and U729 (N_729,N_612,In_522);
nor U730 (N_730,N_654,N_188);
or U731 (N_731,N_485,In_91);
or U732 (N_732,N_220,N_664);
nand U733 (N_733,N_418,N_311);
nand U734 (N_734,N_563,N_653);
xnor U735 (N_735,In_812,N_610);
xor U736 (N_736,N_643,N_669);
nand U737 (N_737,N_602,N_514);
xnor U738 (N_738,N_502,N_628);
and U739 (N_739,N_682,N_82);
nand U740 (N_740,N_681,N_474);
xor U741 (N_741,N_698,N_463);
and U742 (N_742,N_625,N_473);
nand U743 (N_743,N_687,N_511);
xnor U744 (N_744,In_6,N_227);
nor U745 (N_745,N_651,N_476);
xnor U746 (N_746,N_609,N_691);
and U747 (N_747,N_228,N_607);
or U748 (N_748,N_618,N_526);
nand U749 (N_749,In_963,N_55);
xor U750 (N_750,N_203,N_555);
or U751 (N_751,N_640,In_423);
or U752 (N_752,N_515,N_588);
xnor U753 (N_753,N_634,N_601);
nor U754 (N_754,N_639,N_629);
nor U755 (N_755,N_657,N_293);
and U756 (N_756,N_64,In_435);
nand U757 (N_757,N_617,In_762);
nand U758 (N_758,N_580,N_655);
xor U759 (N_759,N_564,N_540);
xnor U760 (N_760,N_577,N_408);
nand U761 (N_761,N_692,N_675);
nand U762 (N_762,In_994,In_624);
nand U763 (N_763,N_121,N_665);
and U764 (N_764,N_248,N_142);
nor U765 (N_765,N_471,N_353);
nand U766 (N_766,N_395,N_635);
and U767 (N_767,N_552,N_542);
xor U768 (N_768,N_566,N_477);
nand U769 (N_769,N_207,N_419);
xnor U770 (N_770,N_490,In_521);
or U771 (N_771,N_505,N_508);
or U772 (N_772,N_668,N_102);
or U773 (N_773,In_866,In_727);
nor U774 (N_774,N_649,In_250);
xor U775 (N_775,N_224,N_679);
xor U776 (N_776,N_663,N_652);
and U777 (N_777,N_620,N_622);
or U778 (N_778,In_851,N_633);
or U779 (N_779,N_646,N_567);
xnor U780 (N_780,N_383,N_472);
and U781 (N_781,N_280,N_536);
or U782 (N_782,In_534,In_704);
or U783 (N_783,N_525,N_489);
nand U784 (N_784,N_666,N_671);
nand U785 (N_785,N_230,N_173);
and U786 (N_786,In_945,N_529);
and U787 (N_787,In_233,In_491);
or U788 (N_788,N_619,N_560);
nand U789 (N_789,In_128,N_305);
or U790 (N_790,In_585,In_903);
nor U791 (N_791,N_650,In_353);
nor U792 (N_792,N_637,N_219);
nor U793 (N_793,N_688,N_70);
nor U794 (N_794,N_684,N_659);
xnor U795 (N_795,N_568,N_535);
nand U796 (N_796,N_453,N_51);
nor U797 (N_797,N_683,N_680);
nand U798 (N_798,N_670,N_600);
or U799 (N_799,N_606,N_631);
and U800 (N_800,N_673,N_716);
nand U801 (N_801,N_76,N_208);
or U802 (N_802,N_605,In_731);
or U803 (N_803,N_621,N_701);
xor U804 (N_804,N_608,In_595);
and U805 (N_805,N_509,N_795);
xnor U806 (N_806,N_703,N_728);
and U807 (N_807,N_783,N_799);
and U808 (N_808,N_759,N_780);
nor U809 (N_809,N_790,N_738);
and U810 (N_810,N_772,In_407);
nor U811 (N_811,N_597,N_604);
nand U812 (N_812,N_709,In_955);
xnor U813 (N_813,N_741,N_702);
nor U814 (N_814,N_690,In_796);
and U815 (N_815,N_720,N_696);
xor U816 (N_816,N_746,N_757);
nor U817 (N_817,N_534,N_707);
xnor U818 (N_818,N_466,N_797);
and U819 (N_819,N_761,N_750);
or U820 (N_820,In_217,N_724);
xor U821 (N_821,N_723,N_792);
xnor U822 (N_822,N_433,N_530);
nor U823 (N_823,N_762,In_684);
nand U824 (N_824,N_596,N_497);
or U825 (N_825,N_781,N_516);
xor U826 (N_826,N_768,N_736);
nand U827 (N_827,N_253,N_726);
or U828 (N_828,N_787,N_747);
and U829 (N_829,N_644,N_705);
nor U830 (N_830,N_779,N_405);
nand U831 (N_831,N_624,N_777);
nor U832 (N_832,N_725,N_767);
nor U833 (N_833,In_888,N_599);
nor U834 (N_834,N_793,N_689);
xnor U835 (N_835,N_789,N_754);
or U836 (N_836,N_714,N_753);
xor U837 (N_837,In_598,N_548);
nor U838 (N_838,N_615,N_522);
xnor U839 (N_839,N_745,N_388);
nand U840 (N_840,N_735,N_582);
and U841 (N_841,N_648,N_678);
nor U842 (N_842,In_717,N_571);
nor U843 (N_843,N_258,In_934);
nand U844 (N_844,N_730,N_785);
nand U845 (N_845,In_408,N_19);
nor U846 (N_846,N_306,N_719);
nand U847 (N_847,N_594,N_737);
or U848 (N_848,In_205,N_729);
xor U849 (N_849,N_710,N_782);
nand U850 (N_850,N_773,N_642);
and U851 (N_851,In_434,In_723);
nor U852 (N_852,N_613,N_647);
xor U853 (N_853,N_775,N_362);
xnor U854 (N_854,N_676,In_264);
nand U855 (N_855,N_764,In_0);
or U856 (N_856,In_943,N_706);
nor U857 (N_857,N_704,N_630);
nor U858 (N_858,N_623,N_434);
xnor U859 (N_859,N_291,N_774);
xor U860 (N_860,N_791,N_756);
or U861 (N_861,N_257,N_148);
nand U862 (N_862,N_677,N_765);
nor U863 (N_863,N_458,N_794);
and U864 (N_864,N_732,N_748);
nor U865 (N_865,N_708,In_832);
nor U866 (N_866,N_721,N_722);
nand U867 (N_867,N_751,N_632);
nand U868 (N_868,N_718,N_356);
nor U869 (N_869,N_700,In_770);
nor U870 (N_870,N_744,N_711);
or U871 (N_871,N_739,N_784);
xor U872 (N_872,N_638,N_656);
nand U873 (N_873,N_523,N_546);
xnor U874 (N_874,N_731,N_444);
or U875 (N_875,N_717,N_769);
xnor U876 (N_876,N_368,N_760);
xnor U877 (N_877,N_743,N_798);
or U878 (N_878,N_778,N_712);
xor U879 (N_879,N_543,N_558);
nand U880 (N_880,N_627,N_734);
or U881 (N_881,N_589,N_661);
or U882 (N_882,N_225,N_788);
xnor U883 (N_883,N_758,N_662);
nand U884 (N_884,In_579,N_576);
nand U885 (N_885,N_796,N_763);
and U886 (N_886,N_742,N_695);
nor U887 (N_887,N_733,N_770);
and U888 (N_888,N_740,N_766);
xnor U889 (N_889,N_776,N_686);
or U890 (N_890,N_699,N_131);
nand U891 (N_891,N_749,N_510);
nor U892 (N_892,N_771,N_494);
or U893 (N_893,N_626,In_839);
or U894 (N_894,In_216,N_164);
and U895 (N_895,N_658,N_727);
xor U896 (N_896,N_685,N_713);
nor U897 (N_897,N_481,N_786);
nand U898 (N_898,N_755,N_752);
xor U899 (N_899,N_260,N_715);
nor U900 (N_900,N_809,N_804);
or U901 (N_901,N_841,N_877);
xor U902 (N_902,N_824,N_836);
nor U903 (N_903,N_899,N_888);
xor U904 (N_904,N_813,N_886);
nor U905 (N_905,N_801,N_851);
xor U906 (N_906,N_843,N_846);
xnor U907 (N_907,N_893,N_839);
nand U908 (N_908,N_811,N_815);
or U909 (N_909,N_870,N_818);
and U910 (N_910,N_891,N_897);
xnor U911 (N_911,N_837,N_829);
nand U912 (N_912,N_802,N_834);
and U913 (N_913,N_867,N_814);
xnor U914 (N_914,N_825,N_828);
and U915 (N_915,N_817,N_847);
nor U916 (N_916,N_878,N_889);
and U917 (N_917,N_859,N_807);
nand U918 (N_918,N_882,N_842);
nor U919 (N_919,N_805,N_863);
nor U920 (N_920,N_850,N_885);
nor U921 (N_921,N_861,N_864);
nand U922 (N_922,N_819,N_879);
xnor U923 (N_923,N_865,N_810);
or U924 (N_924,N_890,N_803);
nand U925 (N_925,N_873,N_855);
or U926 (N_926,N_898,N_830);
and U927 (N_927,N_883,N_816);
nand U928 (N_928,N_826,N_880);
and U929 (N_929,N_822,N_869);
nand U930 (N_930,N_832,N_812);
and U931 (N_931,N_894,N_868);
xor U932 (N_932,N_876,N_854);
xor U933 (N_933,N_866,N_833);
nand U934 (N_934,N_844,N_871);
or U935 (N_935,N_896,N_872);
nor U936 (N_936,N_875,N_820);
or U937 (N_937,N_853,N_856);
and U938 (N_938,N_831,N_849);
nand U939 (N_939,N_845,N_821);
and U940 (N_940,N_848,N_887);
and U941 (N_941,N_835,N_800);
nand U942 (N_942,N_808,N_881);
and U943 (N_943,N_852,N_838);
and U944 (N_944,N_858,N_823);
nand U945 (N_945,N_827,N_895);
nand U946 (N_946,N_860,N_884);
and U947 (N_947,N_892,N_874);
and U948 (N_948,N_840,N_806);
and U949 (N_949,N_857,N_862);
nor U950 (N_950,N_853,N_805);
nor U951 (N_951,N_836,N_865);
xnor U952 (N_952,N_811,N_885);
xor U953 (N_953,N_875,N_822);
nand U954 (N_954,N_884,N_886);
nor U955 (N_955,N_854,N_821);
or U956 (N_956,N_833,N_868);
xnor U957 (N_957,N_815,N_896);
nand U958 (N_958,N_848,N_821);
or U959 (N_959,N_806,N_883);
xor U960 (N_960,N_812,N_891);
and U961 (N_961,N_868,N_800);
nand U962 (N_962,N_898,N_877);
nand U963 (N_963,N_874,N_887);
and U964 (N_964,N_889,N_812);
xnor U965 (N_965,N_843,N_899);
nor U966 (N_966,N_859,N_873);
xor U967 (N_967,N_889,N_881);
xnor U968 (N_968,N_886,N_848);
and U969 (N_969,N_880,N_837);
xnor U970 (N_970,N_819,N_826);
or U971 (N_971,N_818,N_803);
nand U972 (N_972,N_885,N_894);
nand U973 (N_973,N_850,N_826);
nor U974 (N_974,N_828,N_814);
and U975 (N_975,N_827,N_884);
nor U976 (N_976,N_845,N_843);
xnor U977 (N_977,N_891,N_871);
nand U978 (N_978,N_800,N_841);
or U979 (N_979,N_806,N_821);
nor U980 (N_980,N_849,N_899);
nand U981 (N_981,N_863,N_846);
nor U982 (N_982,N_840,N_803);
or U983 (N_983,N_887,N_833);
nand U984 (N_984,N_896,N_878);
xnor U985 (N_985,N_815,N_820);
nor U986 (N_986,N_860,N_804);
and U987 (N_987,N_815,N_817);
nand U988 (N_988,N_877,N_859);
xnor U989 (N_989,N_872,N_856);
and U990 (N_990,N_884,N_848);
or U991 (N_991,N_840,N_874);
and U992 (N_992,N_823,N_874);
nor U993 (N_993,N_865,N_870);
and U994 (N_994,N_842,N_873);
or U995 (N_995,N_822,N_893);
or U996 (N_996,N_898,N_883);
or U997 (N_997,N_881,N_800);
or U998 (N_998,N_862,N_832);
nand U999 (N_999,N_812,N_814);
and U1000 (N_1000,N_983,N_907);
or U1001 (N_1001,N_992,N_958);
nor U1002 (N_1002,N_903,N_905);
nor U1003 (N_1003,N_960,N_924);
nand U1004 (N_1004,N_955,N_953);
nand U1005 (N_1005,N_912,N_936);
xnor U1006 (N_1006,N_949,N_984);
nor U1007 (N_1007,N_978,N_969);
nand U1008 (N_1008,N_980,N_997);
nor U1009 (N_1009,N_922,N_971);
nand U1010 (N_1010,N_935,N_947);
nor U1011 (N_1011,N_916,N_996);
nor U1012 (N_1012,N_986,N_909);
xnor U1013 (N_1013,N_999,N_933);
and U1014 (N_1014,N_956,N_906);
nand U1015 (N_1015,N_928,N_917);
or U1016 (N_1016,N_993,N_923);
xnor U1017 (N_1017,N_946,N_930);
xor U1018 (N_1018,N_942,N_902);
or U1019 (N_1019,N_913,N_944);
and U1020 (N_1020,N_951,N_979);
nand U1021 (N_1021,N_914,N_904);
and U1022 (N_1022,N_990,N_976);
nor U1023 (N_1023,N_966,N_900);
or U1024 (N_1024,N_987,N_967);
or U1025 (N_1025,N_926,N_988);
xor U1026 (N_1026,N_931,N_981);
nand U1027 (N_1027,N_945,N_994);
nor U1028 (N_1028,N_985,N_968);
and U1029 (N_1029,N_974,N_952);
nor U1030 (N_1030,N_973,N_937);
and U1031 (N_1031,N_925,N_910);
or U1032 (N_1032,N_957,N_901);
nand U1033 (N_1033,N_939,N_915);
or U1034 (N_1034,N_977,N_998);
nor U1035 (N_1035,N_921,N_950);
xnor U1036 (N_1036,N_920,N_963);
xor U1037 (N_1037,N_964,N_932);
or U1038 (N_1038,N_911,N_982);
or U1039 (N_1039,N_908,N_961);
nand U1040 (N_1040,N_927,N_918);
xnor U1041 (N_1041,N_959,N_941);
xor U1042 (N_1042,N_943,N_989);
or U1043 (N_1043,N_938,N_975);
xnor U1044 (N_1044,N_954,N_972);
xor U1045 (N_1045,N_995,N_929);
xor U1046 (N_1046,N_934,N_965);
or U1047 (N_1047,N_970,N_940);
nor U1048 (N_1048,N_948,N_919);
and U1049 (N_1049,N_991,N_962);
nand U1050 (N_1050,N_992,N_988);
xor U1051 (N_1051,N_950,N_962);
or U1052 (N_1052,N_989,N_909);
nor U1053 (N_1053,N_932,N_913);
nor U1054 (N_1054,N_988,N_904);
xnor U1055 (N_1055,N_943,N_930);
nor U1056 (N_1056,N_987,N_937);
nand U1057 (N_1057,N_942,N_956);
nand U1058 (N_1058,N_917,N_941);
and U1059 (N_1059,N_942,N_951);
and U1060 (N_1060,N_962,N_916);
nand U1061 (N_1061,N_981,N_945);
xnor U1062 (N_1062,N_945,N_936);
xor U1063 (N_1063,N_991,N_922);
nor U1064 (N_1064,N_974,N_915);
xnor U1065 (N_1065,N_927,N_942);
and U1066 (N_1066,N_951,N_937);
xor U1067 (N_1067,N_934,N_967);
nand U1068 (N_1068,N_948,N_968);
nand U1069 (N_1069,N_968,N_952);
and U1070 (N_1070,N_927,N_980);
or U1071 (N_1071,N_999,N_952);
or U1072 (N_1072,N_946,N_974);
nor U1073 (N_1073,N_975,N_980);
or U1074 (N_1074,N_919,N_917);
and U1075 (N_1075,N_976,N_986);
or U1076 (N_1076,N_929,N_976);
or U1077 (N_1077,N_942,N_926);
or U1078 (N_1078,N_921,N_973);
xnor U1079 (N_1079,N_998,N_917);
and U1080 (N_1080,N_959,N_977);
xor U1081 (N_1081,N_957,N_978);
or U1082 (N_1082,N_953,N_972);
or U1083 (N_1083,N_965,N_926);
and U1084 (N_1084,N_964,N_986);
nand U1085 (N_1085,N_902,N_948);
and U1086 (N_1086,N_997,N_992);
nand U1087 (N_1087,N_924,N_962);
nand U1088 (N_1088,N_950,N_989);
xnor U1089 (N_1089,N_955,N_942);
and U1090 (N_1090,N_918,N_925);
nor U1091 (N_1091,N_999,N_980);
and U1092 (N_1092,N_901,N_991);
and U1093 (N_1093,N_986,N_958);
and U1094 (N_1094,N_937,N_945);
nor U1095 (N_1095,N_945,N_955);
nand U1096 (N_1096,N_938,N_967);
or U1097 (N_1097,N_959,N_991);
nand U1098 (N_1098,N_971,N_947);
or U1099 (N_1099,N_941,N_991);
and U1100 (N_1100,N_1060,N_1068);
xor U1101 (N_1101,N_1045,N_1094);
and U1102 (N_1102,N_1095,N_1000);
or U1103 (N_1103,N_1013,N_1080);
nor U1104 (N_1104,N_1021,N_1078);
nor U1105 (N_1105,N_1066,N_1026);
or U1106 (N_1106,N_1003,N_1099);
nand U1107 (N_1107,N_1065,N_1008);
and U1108 (N_1108,N_1028,N_1057);
and U1109 (N_1109,N_1022,N_1074);
or U1110 (N_1110,N_1047,N_1070);
and U1111 (N_1111,N_1044,N_1035);
or U1112 (N_1112,N_1048,N_1061);
or U1113 (N_1113,N_1043,N_1017);
and U1114 (N_1114,N_1001,N_1031);
nand U1115 (N_1115,N_1064,N_1071);
and U1116 (N_1116,N_1073,N_1011);
and U1117 (N_1117,N_1058,N_1072);
or U1118 (N_1118,N_1020,N_1086);
nand U1119 (N_1119,N_1093,N_1069);
nor U1120 (N_1120,N_1004,N_1040);
nor U1121 (N_1121,N_1038,N_1027);
or U1122 (N_1122,N_1087,N_1075);
nor U1123 (N_1123,N_1052,N_1090);
nor U1124 (N_1124,N_1067,N_1056);
xor U1125 (N_1125,N_1092,N_1012);
nor U1126 (N_1126,N_1054,N_1025);
and U1127 (N_1127,N_1029,N_1024);
or U1128 (N_1128,N_1051,N_1023);
or U1129 (N_1129,N_1033,N_1042);
and U1130 (N_1130,N_1007,N_1085);
or U1131 (N_1131,N_1050,N_1082);
nor U1132 (N_1132,N_1005,N_1032);
nand U1133 (N_1133,N_1006,N_1059);
nand U1134 (N_1134,N_1097,N_1019);
or U1135 (N_1135,N_1076,N_1039);
or U1136 (N_1136,N_1015,N_1062);
or U1137 (N_1137,N_1010,N_1049);
xnor U1138 (N_1138,N_1081,N_1037);
and U1139 (N_1139,N_1016,N_1083);
and U1140 (N_1140,N_1053,N_1055);
or U1141 (N_1141,N_1084,N_1036);
or U1142 (N_1142,N_1091,N_1014);
xor U1143 (N_1143,N_1098,N_1079);
nand U1144 (N_1144,N_1034,N_1089);
xor U1145 (N_1145,N_1096,N_1046);
nand U1146 (N_1146,N_1002,N_1030);
nand U1147 (N_1147,N_1077,N_1018);
and U1148 (N_1148,N_1041,N_1063);
nand U1149 (N_1149,N_1009,N_1088);
or U1150 (N_1150,N_1090,N_1018);
and U1151 (N_1151,N_1035,N_1081);
nor U1152 (N_1152,N_1095,N_1087);
or U1153 (N_1153,N_1011,N_1094);
nor U1154 (N_1154,N_1064,N_1081);
xor U1155 (N_1155,N_1044,N_1008);
nand U1156 (N_1156,N_1077,N_1020);
nor U1157 (N_1157,N_1065,N_1079);
nand U1158 (N_1158,N_1095,N_1060);
nor U1159 (N_1159,N_1094,N_1027);
xor U1160 (N_1160,N_1051,N_1033);
nor U1161 (N_1161,N_1008,N_1085);
nand U1162 (N_1162,N_1093,N_1086);
nand U1163 (N_1163,N_1006,N_1091);
nand U1164 (N_1164,N_1081,N_1059);
or U1165 (N_1165,N_1072,N_1049);
xor U1166 (N_1166,N_1050,N_1065);
and U1167 (N_1167,N_1049,N_1095);
or U1168 (N_1168,N_1085,N_1035);
xnor U1169 (N_1169,N_1035,N_1042);
and U1170 (N_1170,N_1049,N_1016);
nor U1171 (N_1171,N_1051,N_1090);
xnor U1172 (N_1172,N_1043,N_1088);
xor U1173 (N_1173,N_1069,N_1075);
xor U1174 (N_1174,N_1058,N_1022);
nand U1175 (N_1175,N_1026,N_1027);
or U1176 (N_1176,N_1028,N_1066);
nor U1177 (N_1177,N_1083,N_1074);
and U1178 (N_1178,N_1096,N_1024);
or U1179 (N_1179,N_1072,N_1004);
and U1180 (N_1180,N_1035,N_1097);
nand U1181 (N_1181,N_1090,N_1068);
nand U1182 (N_1182,N_1079,N_1052);
nor U1183 (N_1183,N_1089,N_1025);
and U1184 (N_1184,N_1085,N_1090);
and U1185 (N_1185,N_1071,N_1061);
and U1186 (N_1186,N_1067,N_1006);
nand U1187 (N_1187,N_1082,N_1044);
and U1188 (N_1188,N_1031,N_1024);
or U1189 (N_1189,N_1084,N_1044);
xor U1190 (N_1190,N_1071,N_1010);
nand U1191 (N_1191,N_1031,N_1035);
or U1192 (N_1192,N_1028,N_1072);
nor U1193 (N_1193,N_1014,N_1028);
nand U1194 (N_1194,N_1068,N_1064);
xor U1195 (N_1195,N_1041,N_1029);
and U1196 (N_1196,N_1089,N_1062);
xnor U1197 (N_1197,N_1028,N_1015);
nand U1198 (N_1198,N_1058,N_1012);
xor U1199 (N_1199,N_1059,N_1035);
xor U1200 (N_1200,N_1178,N_1153);
nand U1201 (N_1201,N_1129,N_1179);
and U1202 (N_1202,N_1181,N_1110);
and U1203 (N_1203,N_1194,N_1190);
nand U1204 (N_1204,N_1133,N_1112);
nor U1205 (N_1205,N_1191,N_1162);
nor U1206 (N_1206,N_1103,N_1121);
xor U1207 (N_1207,N_1119,N_1108);
nand U1208 (N_1208,N_1107,N_1171);
xnor U1209 (N_1209,N_1196,N_1188);
nand U1210 (N_1210,N_1138,N_1137);
nor U1211 (N_1211,N_1167,N_1117);
or U1212 (N_1212,N_1114,N_1172);
nor U1213 (N_1213,N_1157,N_1173);
nand U1214 (N_1214,N_1141,N_1126);
nor U1215 (N_1215,N_1120,N_1101);
nand U1216 (N_1216,N_1128,N_1116);
nand U1217 (N_1217,N_1113,N_1140);
xor U1218 (N_1218,N_1160,N_1192);
nor U1219 (N_1219,N_1104,N_1195);
and U1220 (N_1220,N_1131,N_1100);
nand U1221 (N_1221,N_1127,N_1151);
nor U1222 (N_1222,N_1132,N_1136);
or U1223 (N_1223,N_1145,N_1161);
nor U1224 (N_1224,N_1142,N_1135);
nor U1225 (N_1225,N_1111,N_1124);
and U1226 (N_1226,N_1187,N_1182);
xnor U1227 (N_1227,N_1122,N_1154);
nand U1228 (N_1228,N_1193,N_1146);
or U1229 (N_1229,N_1165,N_1176);
xor U1230 (N_1230,N_1105,N_1170);
nor U1231 (N_1231,N_1148,N_1174);
or U1232 (N_1232,N_1183,N_1115);
or U1233 (N_1233,N_1155,N_1144);
nor U1234 (N_1234,N_1185,N_1177);
xnor U1235 (N_1235,N_1123,N_1106);
nor U1236 (N_1236,N_1147,N_1125);
or U1237 (N_1237,N_1149,N_1197);
xor U1238 (N_1238,N_1198,N_1109);
and U1239 (N_1239,N_1186,N_1102);
and U1240 (N_1240,N_1134,N_1199);
xor U1241 (N_1241,N_1164,N_1130);
nor U1242 (N_1242,N_1166,N_1169);
and U1243 (N_1243,N_1175,N_1168);
or U1244 (N_1244,N_1150,N_1184);
xnor U1245 (N_1245,N_1180,N_1163);
or U1246 (N_1246,N_1159,N_1189);
xor U1247 (N_1247,N_1156,N_1152);
nor U1248 (N_1248,N_1143,N_1158);
nand U1249 (N_1249,N_1118,N_1139);
nor U1250 (N_1250,N_1165,N_1161);
nor U1251 (N_1251,N_1180,N_1192);
nand U1252 (N_1252,N_1165,N_1151);
nand U1253 (N_1253,N_1133,N_1140);
xor U1254 (N_1254,N_1111,N_1129);
xor U1255 (N_1255,N_1164,N_1126);
or U1256 (N_1256,N_1189,N_1147);
xnor U1257 (N_1257,N_1198,N_1148);
xor U1258 (N_1258,N_1117,N_1190);
or U1259 (N_1259,N_1140,N_1152);
or U1260 (N_1260,N_1152,N_1177);
nand U1261 (N_1261,N_1170,N_1142);
nand U1262 (N_1262,N_1169,N_1107);
nor U1263 (N_1263,N_1127,N_1113);
and U1264 (N_1264,N_1126,N_1158);
nand U1265 (N_1265,N_1113,N_1198);
xnor U1266 (N_1266,N_1155,N_1187);
nand U1267 (N_1267,N_1139,N_1184);
and U1268 (N_1268,N_1142,N_1136);
and U1269 (N_1269,N_1179,N_1130);
xor U1270 (N_1270,N_1121,N_1194);
and U1271 (N_1271,N_1144,N_1132);
xor U1272 (N_1272,N_1196,N_1159);
nor U1273 (N_1273,N_1180,N_1140);
nand U1274 (N_1274,N_1198,N_1190);
and U1275 (N_1275,N_1171,N_1130);
nand U1276 (N_1276,N_1104,N_1156);
and U1277 (N_1277,N_1113,N_1183);
xor U1278 (N_1278,N_1124,N_1107);
or U1279 (N_1279,N_1145,N_1134);
or U1280 (N_1280,N_1139,N_1199);
nand U1281 (N_1281,N_1186,N_1101);
xor U1282 (N_1282,N_1190,N_1122);
nand U1283 (N_1283,N_1170,N_1151);
nor U1284 (N_1284,N_1116,N_1191);
nand U1285 (N_1285,N_1185,N_1158);
xnor U1286 (N_1286,N_1107,N_1100);
or U1287 (N_1287,N_1117,N_1191);
and U1288 (N_1288,N_1182,N_1184);
nand U1289 (N_1289,N_1102,N_1177);
xor U1290 (N_1290,N_1172,N_1107);
xor U1291 (N_1291,N_1107,N_1144);
and U1292 (N_1292,N_1127,N_1179);
or U1293 (N_1293,N_1153,N_1129);
and U1294 (N_1294,N_1131,N_1103);
xor U1295 (N_1295,N_1108,N_1139);
and U1296 (N_1296,N_1143,N_1107);
nor U1297 (N_1297,N_1154,N_1128);
or U1298 (N_1298,N_1153,N_1111);
or U1299 (N_1299,N_1135,N_1166);
xnor U1300 (N_1300,N_1295,N_1298);
and U1301 (N_1301,N_1260,N_1216);
nor U1302 (N_1302,N_1207,N_1246);
nor U1303 (N_1303,N_1258,N_1244);
nor U1304 (N_1304,N_1236,N_1203);
nand U1305 (N_1305,N_1233,N_1250);
or U1306 (N_1306,N_1297,N_1217);
nand U1307 (N_1307,N_1200,N_1286);
xor U1308 (N_1308,N_1221,N_1256);
xnor U1309 (N_1309,N_1213,N_1225);
xnor U1310 (N_1310,N_1230,N_1211);
nand U1311 (N_1311,N_1210,N_1204);
xnor U1312 (N_1312,N_1280,N_1271);
nor U1313 (N_1313,N_1231,N_1290);
or U1314 (N_1314,N_1284,N_1257);
and U1315 (N_1315,N_1288,N_1292);
nand U1316 (N_1316,N_1259,N_1261);
nor U1317 (N_1317,N_1267,N_1220);
xor U1318 (N_1318,N_1278,N_1239);
and U1319 (N_1319,N_1249,N_1223);
or U1320 (N_1320,N_1289,N_1287);
and U1321 (N_1321,N_1265,N_1266);
nor U1322 (N_1322,N_1206,N_1219);
and U1323 (N_1323,N_1205,N_1283);
or U1324 (N_1324,N_1224,N_1228);
and U1325 (N_1325,N_1272,N_1227);
and U1326 (N_1326,N_1247,N_1296);
and U1327 (N_1327,N_1299,N_1214);
nand U1328 (N_1328,N_1282,N_1281);
xor U1329 (N_1329,N_1234,N_1215);
or U1330 (N_1330,N_1201,N_1273);
or U1331 (N_1331,N_1263,N_1240);
xnor U1332 (N_1332,N_1232,N_1218);
and U1333 (N_1333,N_1253,N_1208);
xor U1334 (N_1334,N_1274,N_1277);
or U1335 (N_1335,N_1243,N_1255);
nand U1336 (N_1336,N_1241,N_1270);
and U1337 (N_1337,N_1242,N_1276);
nor U1338 (N_1338,N_1212,N_1251);
nor U1339 (N_1339,N_1229,N_1245);
or U1340 (N_1340,N_1291,N_1202);
nor U1341 (N_1341,N_1238,N_1294);
and U1342 (N_1342,N_1269,N_1209);
and U1343 (N_1343,N_1248,N_1252);
xor U1344 (N_1344,N_1237,N_1235);
xor U1345 (N_1345,N_1275,N_1262);
nand U1346 (N_1346,N_1293,N_1279);
and U1347 (N_1347,N_1264,N_1268);
nand U1348 (N_1348,N_1226,N_1285);
xor U1349 (N_1349,N_1254,N_1222);
nand U1350 (N_1350,N_1285,N_1217);
or U1351 (N_1351,N_1230,N_1281);
and U1352 (N_1352,N_1205,N_1248);
nand U1353 (N_1353,N_1225,N_1279);
nand U1354 (N_1354,N_1277,N_1221);
and U1355 (N_1355,N_1211,N_1266);
nand U1356 (N_1356,N_1293,N_1251);
xnor U1357 (N_1357,N_1236,N_1294);
xor U1358 (N_1358,N_1286,N_1209);
xnor U1359 (N_1359,N_1227,N_1250);
xor U1360 (N_1360,N_1250,N_1256);
nor U1361 (N_1361,N_1255,N_1249);
nand U1362 (N_1362,N_1252,N_1295);
and U1363 (N_1363,N_1263,N_1243);
or U1364 (N_1364,N_1292,N_1228);
nor U1365 (N_1365,N_1210,N_1237);
or U1366 (N_1366,N_1243,N_1264);
xor U1367 (N_1367,N_1229,N_1298);
xor U1368 (N_1368,N_1288,N_1213);
and U1369 (N_1369,N_1200,N_1250);
nor U1370 (N_1370,N_1234,N_1276);
and U1371 (N_1371,N_1222,N_1224);
nand U1372 (N_1372,N_1240,N_1250);
and U1373 (N_1373,N_1205,N_1218);
or U1374 (N_1374,N_1220,N_1244);
nor U1375 (N_1375,N_1217,N_1291);
xnor U1376 (N_1376,N_1210,N_1270);
nor U1377 (N_1377,N_1296,N_1230);
xor U1378 (N_1378,N_1234,N_1273);
or U1379 (N_1379,N_1206,N_1226);
nand U1380 (N_1380,N_1209,N_1276);
nor U1381 (N_1381,N_1256,N_1280);
nand U1382 (N_1382,N_1224,N_1233);
xnor U1383 (N_1383,N_1210,N_1213);
nand U1384 (N_1384,N_1208,N_1295);
nand U1385 (N_1385,N_1225,N_1235);
or U1386 (N_1386,N_1293,N_1289);
or U1387 (N_1387,N_1232,N_1248);
xnor U1388 (N_1388,N_1255,N_1234);
and U1389 (N_1389,N_1202,N_1229);
nor U1390 (N_1390,N_1260,N_1206);
or U1391 (N_1391,N_1207,N_1266);
nor U1392 (N_1392,N_1207,N_1256);
xor U1393 (N_1393,N_1213,N_1247);
or U1394 (N_1394,N_1286,N_1277);
nor U1395 (N_1395,N_1262,N_1249);
nand U1396 (N_1396,N_1239,N_1292);
or U1397 (N_1397,N_1210,N_1223);
nand U1398 (N_1398,N_1281,N_1278);
nor U1399 (N_1399,N_1205,N_1268);
and U1400 (N_1400,N_1386,N_1310);
nor U1401 (N_1401,N_1338,N_1396);
xor U1402 (N_1402,N_1346,N_1336);
nand U1403 (N_1403,N_1351,N_1332);
xor U1404 (N_1404,N_1365,N_1307);
xnor U1405 (N_1405,N_1334,N_1363);
and U1406 (N_1406,N_1316,N_1357);
or U1407 (N_1407,N_1350,N_1313);
nand U1408 (N_1408,N_1319,N_1368);
nor U1409 (N_1409,N_1388,N_1366);
nand U1410 (N_1410,N_1306,N_1371);
nand U1411 (N_1411,N_1303,N_1374);
or U1412 (N_1412,N_1300,N_1343);
or U1413 (N_1413,N_1328,N_1387);
or U1414 (N_1414,N_1331,N_1393);
xnor U1415 (N_1415,N_1376,N_1337);
and U1416 (N_1416,N_1390,N_1324);
and U1417 (N_1417,N_1384,N_1380);
and U1418 (N_1418,N_1301,N_1308);
and U1419 (N_1419,N_1381,N_1317);
nor U1420 (N_1420,N_1330,N_1392);
nand U1421 (N_1421,N_1359,N_1318);
nor U1422 (N_1422,N_1391,N_1394);
xnor U1423 (N_1423,N_1344,N_1397);
and U1424 (N_1424,N_1341,N_1339);
or U1425 (N_1425,N_1398,N_1321);
or U1426 (N_1426,N_1342,N_1352);
or U1427 (N_1427,N_1362,N_1304);
nor U1428 (N_1428,N_1358,N_1340);
nand U1429 (N_1429,N_1314,N_1311);
or U1430 (N_1430,N_1375,N_1320);
and U1431 (N_1431,N_1309,N_1305);
or U1432 (N_1432,N_1372,N_1353);
nor U1433 (N_1433,N_1399,N_1335);
nor U1434 (N_1434,N_1329,N_1345);
nand U1435 (N_1435,N_1348,N_1354);
xnor U1436 (N_1436,N_1373,N_1385);
nand U1437 (N_1437,N_1349,N_1325);
nand U1438 (N_1438,N_1322,N_1347);
or U1439 (N_1439,N_1356,N_1379);
nand U1440 (N_1440,N_1364,N_1315);
and U1441 (N_1441,N_1312,N_1361);
or U1442 (N_1442,N_1395,N_1377);
or U1443 (N_1443,N_1382,N_1355);
xnor U1444 (N_1444,N_1369,N_1302);
nor U1445 (N_1445,N_1378,N_1360);
and U1446 (N_1446,N_1333,N_1370);
and U1447 (N_1447,N_1326,N_1327);
xor U1448 (N_1448,N_1389,N_1323);
nand U1449 (N_1449,N_1367,N_1383);
xnor U1450 (N_1450,N_1338,N_1313);
xnor U1451 (N_1451,N_1314,N_1306);
nand U1452 (N_1452,N_1357,N_1328);
nand U1453 (N_1453,N_1340,N_1390);
or U1454 (N_1454,N_1331,N_1373);
and U1455 (N_1455,N_1385,N_1312);
nand U1456 (N_1456,N_1329,N_1308);
and U1457 (N_1457,N_1362,N_1307);
nor U1458 (N_1458,N_1309,N_1310);
or U1459 (N_1459,N_1311,N_1342);
nor U1460 (N_1460,N_1381,N_1323);
nor U1461 (N_1461,N_1362,N_1397);
or U1462 (N_1462,N_1303,N_1357);
nor U1463 (N_1463,N_1323,N_1376);
nand U1464 (N_1464,N_1341,N_1349);
nand U1465 (N_1465,N_1326,N_1398);
nor U1466 (N_1466,N_1325,N_1326);
nor U1467 (N_1467,N_1363,N_1314);
and U1468 (N_1468,N_1374,N_1313);
xnor U1469 (N_1469,N_1352,N_1319);
nand U1470 (N_1470,N_1379,N_1349);
and U1471 (N_1471,N_1396,N_1361);
and U1472 (N_1472,N_1399,N_1315);
nor U1473 (N_1473,N_1354,N_1369);
xor U1474 (N_1474,N_1344,N_1301);
xor U1475 (N_1475,N_1365,N_1379);
or U1476 (N_1476,N_1337,N_1384);
nor U1477 (N_1477,N_1393,N_1390);
xnor U1478 (N_1478,N_1325,N_1389);
nor U1479 (N_1479,N_1312,N_1398);
nand U1480 (N_1480,N_1320,N_1354);
and U1481 (N_1481,N_1356,N_1355);
and U1482 (N_1482,N_1354,N_1318);
nand U1483 (N_1483,N_1357,N_1321);
nand U1484 (N_1484,N_1329,N_1307);
nand U1485 (N_1485,N_1305,N_1375);
or U1486 (N_1486,N_1361,N_1300);
nand U1487 (N_1487,N_1392,N_1344);
xor U1488 (N_1488,N_1381,N_1346);
and U1489 (N_1489,N_1302,N_1326);
nor U1490 (N_1490,N_1370,N_1346);
nor U1491 (N_1491,N_1304,N_1375);
or U1492 (N_1492,N_1363,N_1318);
or U1493 (N_1493,N_1323,N_1303);
nand U1494 (N_1494,N_1354,N_1386);
xnor U1495 (N_1495,N_1333,N_1377);
or U1496 (N_1496,N_1309,N_1382);
xor U1497 (N_1497,N_1320,N_1338);
nand U1498 (N_1498,N_1333,N_1303);
and U1499 (N_1499,N_1339,N_1314);
and U1500 (N_1500,N_1482,N_1421);
nor U1501 (N_1501,N_1403,N_1490);
xnor U1502 (N_1502,N_1466,N_1461);
and U1503 (N_1503,N_1440,N_1494);
and U1504 (N_1504,N_1439,N_1429);
nand U1505 (N_1505,N_1408,N_1432);
and U1506 (N_1506,N_1474,N_1471);
xnor U1507 (N_1507,N_1450,N_1484);
nand U1508 (N_1508,N_1468,N_1460);
and U1509 (N_1509,N_1485,N_1472);
xnor U1510 (N_1510,N_1449,N_1411);
xor U1511 (N_1511,N_1420,N_1441);
xnor U1512 (N_1512,N_1454,N_1480);
nand U1513 (N_1513,N_1469,N_1402);
nand U1514 (N_1514,N_1462,N_1426);
and U1515 (N_1515,N_1434,N_1478);
nor U1516 (N_1516,N_1491,N_1400);
or U1517 (N_1517,N_1487,N_1419);
xor U1518 (N_1518,N_1412,N_1442);
nand U1519 (N_1519,N_1464,N_1495);
or U1520 (N_1520,N_1430,N_1413);
and U1521 (N_1521,N_1455,N_1467);
nand U1522 (N_1522,N_1404,N_1473);
nand U1523 (N_1523,N_1477,N_1458);
or U1524 (N_1524,N_1418,N_1447);
or U1525 (N_1525,N_1407,N_1481);
and U1526 (N_1526,N_1486,N_1415);
nor U1527 (N_1527,N_1446,N_1499);
or U1528 (N_1528,N_1451,N_1463);
nand U1529 (N_1529,N_1417,N_1433);
nand U1530 (N_1530,N_1456,N_1410);
nor U1531 (N_1531,N_1444,N_1488);
or U1532 (N_1532,N_1475,N_1483);
and U1533 (N_1533,N_1459,N_1496);
xor U1534 (N_1534,N_1414,N_1435);
and U1535 (N_1535,N_1465,N_1428);
nor U1536 (N_1536,N_1416,N_1425);
xor U1537 (N_1537,N_1453,N_1427);
xor U1538 (N_1538,N_1422,N_1479);
nand U1539 (N_1539,N_1424,N_1438);
or U1540 (N_1540,N_1452,N_1470);
xnor U1541 (N_1541,N_1409,N_1445);
nand U1542 (N_1542,N_1492,N_1498);
and U1543 (N_1543,N_1406,N_1448);
xnor U1544 (N_1544,N_1457,N_1497);
and U1545 (N_1545,N_1423,N_1443);
nor U1546 (N_1546,N_1401,N_1476);
xor U1547 (N_1547,N_1431,N_1436);
or U1548 (N_1548,N_1405,N_1489);
and U1549 (N_1549,N_1437,N_1493);
or U1550 (N_1550,N_1469,N_1463);
nor U1551 (N_1551,N_1463,N_1409);
xnor U1552 (N_1552,N_1476,N_1414);
and U1553 (N_1553,N_1424,N_1447);
and U1554 (N_1554,N_1451,N_1494);
nand U1555 (N_1555,N_1477,N_1426);
xor U1556 (N_1556,N_1421,N_1450);
nand U1557 (N_1557,N_1455,N_1472);
nor U1558 (N_1558,N_1404,N_1445);
nor U1559 (N_1559,N_1462,N_1464);
or U1560 (N_1560,N_1443,N_1433);
nor U1561 (N_1561,N_1453,N_1488);
and U1562 (N_1562,N_1499,N_1452);
or U1563 (N_1563,N_1488,N_1415);
nor U1564 (N_1564,N_1460,N_1435);
and U1565 (N_1565,N_1408,N_1454);
and U1566 (N_1566,N_1464,N_1461);
nor U1567 (N_1567,N_1482,N_1445);
and U1568 (N_1568,N_1470,N_1403);
or U1569 (N_1569,N_1466,N_1408);
xnor U1570 (N_1570,N_1456,N_1427);
or U1571 (N_1571,N_1404,N_1455);
and U1572 (N_1572,N_1449,N_1454);
xnor U1573 (N_1573,N_1407,N_1488);
and U1574 (N_1574,N_1498,N_1414);
xnor U1575 (N_1575,N_1450,N_1423);
nand U1576 (N_1576,N_1464,N_1426);
nand U1577 (N_1577,N_1412,N_1406);
xnor U1578 (N_1578,N_1455,N_1438);
or U1579 (N_1579,N_1425,N_1402);
xor U1580 (N_1580,N_1408,N_1440);
nand U1581 (N_1581,N_1490,N_1498);
nand U1582 (N_1582,N_1413,N_1458);
nor U1583 (N_1583,N_1478,N_1487);
and U1584 (N_1584,N_1411,N_1491);
and U1585 (N_1585,N_1477,N_1405);
or U1586 (N_1586,N_1445,N_1441);
nor U1587 (N_1587,N_1405,N_1482);
nand U1588 (N_1588,N_1443,N_1450);
and U1589 (N_1589,N_1455,N_1421);
nand U1590 (N_1590,N_1477,N_1401);
nand U1591 (N_1591,N_1446,N_1437);
or U1592 (N_1592,N_1499,N_1498);
xnor U1593 (N_1593,N_1436,N_1471);
nand U1594 (N_1594,N_1480,N_1489);
nor U1595 (N_1595,N_1481,N_1406);
nand U1596 (N_1596,N_1420,N_1483);
and U1597 (N_1597,N_1472,N_1412);
xor U1598 (N_1598,N_1410,N_1422);
or U1599 (N_1599,N_1489,N_1472);
xnor U1600 (N_1600,N_1517,N_1588);
xnor U1601 (N_1601,N_1572,N_1528);
or U1602 (N_1602,N_1554,N_1555);
xor U1603 (N_1603,N_1573,N_1585);
nor U1604 (N_1604,N_1567,N_1538);
nand U1605 (N_1605,N_1575,N_1563);
and U1606 (N_1606,N_1594,N_1531);
or U1607 (N_1607,N_1597,N_1542);
and U1608 (N_1608,N_1532,N_1503);
xor U1609 (N_1609,N_1521,N_1514);
xor U1610 (N_1610,N_1509,N_1508);
nand U1611 (N_1611,N_1586,N_1539);
nor U1612 (N_1612,N_1535,N_1504);
and U1613 (N_1613,N_1560,N_1571);
or U1614 (N_1614,N_1502,N_1598);
and U1615 (N_1615,N_1537,N_1582);
nand U1616 (N_1616,N_1518,N_1536);
or U1617 (N_1617,N_1548,N_1595);
and U1618 (N_1618,N_1546,N_1553);
nand U1619 (N_1619,N_1559,N_1564);
xor U1620 (N_1620,N_1556,N_1534);
nor U1621 (N_1621,N_1526,N_1576);
or U1622 (N_1622,N_1519,N_1550);
xor U1623 (N_1623,N_1561,N_1589);
xnor U1624 (N_1624,N_1558,N_1583);
nand U1625 (N_1625,N_1525,N_1501);
nand U1626 (N_1626,N_1510,N_1520);
nor U1627 (N_1627,N_1557,N_1513);
nor U1628 (N_1628,N_1581,N_1590);
nand U1629 (N_1629,N_1569,N_1545);
nor U1630 (N_1630,N_1579,N_1527);
nand U1631 (N_1631,N_1544,N_1593);
xnor U1632 (N_1632,N_1577,N_1511);
xnor U1633 (N_1633,N_1530,N_1515);
or U1634 (N_1634,N_1533,N_1591);
nor U1635 (N_1635,N_1574,N_1578);
xor U1636 (N_1636,N_1524,N_1505);
or U1637 (N_1637,N_1547,N_1543);
nor U1638 (N_1638,N_1549,N_1523);
nor U1639 (N_1639,N_1587,N_1592);
xor U1640 (N_1640,N_1580,N_1516);
or U1641 (N_1641,N_1552,N_1522);
xor U1642 (N_1642,N_1596,N_1566);
or U1643 (N_1643,N_1599,N_1570);
or U1644 (N_1644,N_1565,N_1540);
nor U1645 (N_1645,N_1584,N_1562);
xnor U1646 (N_1646,N_1507,N_1500);
or U1647 (N_1647,N_1512,N_1551);
and U1648 (N_1648,N_1541,N_1568);
and U1649 (N_1649,N_1529,N_1506);
nor U1650 (N_1650,N_1553,N_1547);
nand U1651 (N_1651,N_1500,N_1508);
nor U1652 (N_1652,N_1525,N_1596);
and U1653 (N_1653,N_1525,N_1533);
nor U1654 (N_1654,N_1503,N_1595);
and U1655 (N_1655,N_1513,N_1545);
nand U1656 (N_1656,N_1597,N_1529);
or U1657 (N_1657,N_1503,N_1593);
or U1658 (N_1658,N_1567,N_1505);
or U1659 (N_1659,N_1581,N_1599);
or U1660 (N_1660,N_1544,N_1598);
nand U1661 (N_1661,N_1583,N_1546);
nand U1662 (N_1662,N_1555,N_1514);
xor U1663 (N_1663,N_1520,N_1559);
and U1664 (N_1664,N_1582,N_1532);
and U1665 (N_1665,N_1539,N_1564);
xnor U1666 (N_1666,N_1584,N_1515);
nand U1667 (N_1667,N_1564,N_1520);
xor U1668 (N_1668,N_1559,N_1589);
and U1669 (N_1669,N_1555,N_1552);
nand U1670 (N_1670,N_1557,N_1554);
xnor U1671 (N_1671,N_1536,N_1514);
nor U1672 (N_1672,N_1517,N_1536);
nor U1673 (N_1673,N_1557,N_1543);
and U1674 (N_1674,N_1510,N_1551);
nand U1675 (N_1675,N_1550,N_1523);
nor U1676 (N_1676,N_1536,N_1504);
xnor U1677 (N_1677,N_1564,N_1555);
xnor U1678 (N_1678,N_1557,N_1529);
or U1679 (N_1679,N_1505,N_1528);
and U1680 (N_1680,N_1544,N_1513);
nor U1681 (N_1681,N_1561,N_1516);
xnor U1682 (N_1682,N_1511,N_1548);
nand U1683 (N_1683,N_1556,N_1532);
nor U1684 (N_1684,N_1587,N_1552);
and U1685 (N_1685,N_1549,N_1511);
nor U1686 (N_1686,N_1543,N_1556);
or U1687 (N_1687,N_1596,N_1578);
or U1688 (N_1688,N_1559,N_1540);
and U1689 (N_1689,N_1580,N_1534);
or U1690 (N_1690,N_1577,N_1512);
nor U1691 (N_1691,N_1575,N_1592);
and U1692 (N_1692,N_1567,N_1569);
or U1693 (N_1693,N_1502,N_1590);
nor U1694 (N_1694,N_1529,N_1553);
or U1695 (N_1695,N_1552,N_1584);
and U1696 (N_1696,N_1581,N_1524);
xor U1697 (N_1697,N_1549,N_1518);
nor U1698 (N_1698,N_1514,N_1515);
xnor U1699 (N_1699,N_1586,N_1530);
and U1700 (N_1700,N_1665,N_1669);
or U1701 (N_1701,N_1659,N_1617);
or U1702 (N_1702,N_1662,N_1676);
and U1703 (N_1703,N_1697,N_1605);
nand U1704 (N_1704,N_1642,N_1638);
xor U1705 (N_1705,N_1683,N_1633);
nor U1706 (N_1706,N_1609,N_1623);
and U1707 (N_1707,N_1691,N_1645);
xor U1708 (N_1708,N_1626,N_1644);
and U1709 (N_1709,N_1603,N_1621);
and U1710 (N_1710,N_1639,N_1654);
nor U1711 (N_1711,N_1622,N_1646);
nor U1712 (N_1712,N_1661,N_1643);
nand U1713 (N_1713,N_1684,N_1655);
xor U1714 (N_1714,N_1616,N_1651);
xor U1715 (N_1715,N_1673,N_1658);
nand U1716 (N_1716,N_1677,N_1660);
nor U1717 (N_1717,N_1624,N_1694);
xor U1718 (N_1718,N_1688,N_1640);
or U1719 (N_1719,N_1664,N_1618);
or U1720 (N_1720,N_1612,N_1674);
nand U1721 (N_1721,N_1620,N_1671);
nor U1722 (N_1722,N_1601,N_1656);
and U1723 (N_1723,N_1629,N_1670);
and U1724 (N_1724,N_1647,N_1649);
or U1725 (N_1725,N_1687,N_1695);
or U1726 (N_1726,N_1680,N_1614);
xnor U1727 (N_1727,N_1698,N_1692);
and U1728 (N_1728,N_1630,N_1636);
nand U1729 (N_1729,N_1667,N_1600);
xnor U1730 (N_1730,N_1602,N_1619);
or U1731 (N_1731,N_1610,N_1634);
nor U1732 (N_1732,N_1625,N_1689);
xnor U1733 (N_1733,N_1657,N_1604);
or U1734 (N_1734,N_1699,N_1666);
nand U1735 (N_1735,N_1693,N_1615);
xor U1736 (N_1736,N_1650,N_1696);
nor U1737 (N_1737,N_1608,N_1682);
and U1738 (N_1738,N_1653,N_1678);
nand U1739 (N_1739,N_1631,N_1635);
or U1740 (N_1740,N_1611,N_1663);
and U1741 (N_1741,N_1681,N_1607);
nand U1742 (N_1742,N_1672,N_1613);
or U1743 (N_1743,N_1652,N_1675);
and U1744 (N_1744,N_1632,N_1637);
xor U1745 (N_1745,N_1690,N_1606);
or U1746 (N_1746,N_1648,N_1679);
xnor U1747 (N_1747,N_1628,N_1668);
and U1748 (N_1748,N_1641,N_1627);
xnor U1749 (N_1749,N_1685,N_1686);
nor U1750 (N_1750,N_1619,N_1664);
nand U1751 (N_1751,N_1662,N_1621);
nand U1752 (N_1752,N_1608,N_1652);
nand U1753 (N_1753,N_1620,N_1659);
and U1754 (N_1754,N_1614,N_1687);
nor U1755 (N_1755,N_1607,N_1619);
or U1756 (N_1756,N_1699,N_1611);
xnor U1757 (N_1757,N_1634,N_1651);
nand U1758 (N_1758,N_1688,N_1695);
nand U1759 (N_1759,N_1677,N_1617);
xnor U1760 (N_1760,N_1684,N_1646);
and U1761 (N_1761,N_1689,N_1690);
nor U1762 (N_1762,N_1694,N_1683);
and U1763 (N_1763,N_1632,N_1613);
xor U1764 (N_1764,N_1695,N_1622);
and U1765 (N_1765,N_1630,N_1660);
xor U1766 (N_1766,N_1699,N_1634);
nand U1767 (N_1767,N_1680,N_1686);
nor U1768 (N_1768,N_1635,N_1602);
nor U1769 (N_1769,N_1608,N_1638);
or U1770 (N_1770,N_1639,N_1679);
xor U1771 (N_1771,N_1652,N_1685);
nand U1772 (N_1772,N_1666,N_1618);
or U1773 (N_1773,N_1651,N_1686);
xnor U1774 (N_1774,N_1658,N_1682);
nor U1775 (N_1775,N_1663,N_1614);
nor U1776 (N_1776,N_1651,N_1683);
xnor U1777 (N_1777,N_1659,N_1693);
or U1778 (N_1778,N_1645,N_1697);
nand U1779 (N_1779,N_1654,N_1613);
or U1780 (N_1780,N_1636,N_1643);
nand U1781 (N_1781,N_1648,N_1610);
nand U1782 (N_1782,N_1621,N_1620);
or U1783 (N_1783,N_1669,N_1698);
or U1784 (N_1784,N_1683,N_1614);
nor U1785 (N_1785,N_1636,N_1625);
xor U1786 (N_1786,N_1671,N_1696);
or U1787 (N_1787,N_1646,N_1669);
nor U1788 (N_1788,N_1655,N_1640);
xor U1789 (N_1789,N_1603,N_1673);
and U1790 (N_1790,N_1663,N_1664);
and U1791 (N_1791,N_1674,N_1666);
and U1792 (N_1792,N_1694,N_1600);
or U1793 (N_1793,N_1639,N_1673);
xor U1794 (N_1794,N_1613,N_1642);
or U1795 (N_1795,N_1652,N_1632);
nand U1796 (N_1796,N_1606,N_1688);
nand U1797 (N_1797,N_1601,N_1693);
nand U1798 (N_1798,N_1671,N_1635);
nor U1799 (N_1799,N_1684,N_1617);
xor U1800 (N_1800,N_1748,N_1715);
xor U1801 (N_1801,N_1722,N_1728);
or U1802 (N_1802,N_1778,N_1753);
xor U1803 (N_1803,N_1763,N_1777);
nand U1804 (N_1804,N_1794,N_1786);
nand U1805 (N_1805,N_1745,N_1711);
and U1806 (N_1806,N_1717,N_1706);
and U1807 (N_1807,N_1771,N_1754);
or U1808 (N_1808,N_1795,N_1770);
xor U1809 (N_1809,N_1732,N_1756);
nor U1810 (N_1810,N_1784,N_1734);
or U1811 (N_1811,N_1727,N_1791);
nand U1812 (N_1812,N_1767,N_1792);
or U1813 (N_1813,N_1743,N_1721);
or U1814 (N_1814,N_1713,N_1768);
nor U1815 (N_1815,N_1700,N_1789);
nand U1816 (N_1816,N_1729,N_1796);
nor U1817 (N_1817,N_1774,N_1779);
or U1818 (N_1818,N_1709,N_1781);
xnor U1819 (N_1819,N_1737,N_1747);
nor U1820 (N_1820,N_1765,N_1735);
xor U1821 (N_1821,N_1787,N_1723);
or U1822 (N_1822,N_1764,N_1757);
and U1823 (N_1823,N_1704,N_1798);
nand U1824 (N_1824,N_1755,N_1769);
nand U1825 (N_1825,N_1710,N_1733);
or U1826 (N_1826,N_1760,N_1707);
xor U1827 (N_1827,N_1758,N_1714);
nor U1828 (N_1828,N_1730,N_1797);
and U1829 (N_1829,N_1742,N_1744);
xor U1830 (N_1830,N_1785,N_1708);
or U1831 (N_1831,N_1750,N_1776);
nor U1832 (N_1832,N_1740,N_1759);
xnor U1833 (N_1833,N_1718,N_1703);
nand U1834 (N_1834,N_1724,N_1783);
nor U1835 (N_1835,N_1788,N_1799);
xor U1836 (N_1836,N_1775,N_1782);
nor U1837 (N_1837,N_1766,N_1719);
and U1838 (N_1838,N_1793,N_1772);
or U1839 (N_1839,N_1741,N_1739);
and U1840 (N_1840,N_1780,N_1716);
or U1841 (N_1841,N_1761,N_1705);
nand U1842 (N_1842,N_1720,N_1731);
xor U1843 (N_1843,N_1762,N_1738);
xor U1844 (N_1844,N_1749,N_1712);
and U1845 (N_1845,N_1701,N_1746);
nor U1846 (N_1846,N_1702,N_1726);
xnor U1847 (N_1847,N_1790,N_1725);
nor U1848 (N_1848,N_1773,N_1751);
xnor U1849 (N_1849,N_1752,N_1736);
nor U1850 (N_1850,N_1704,N_1707);
and U1851 (N_1851,N_1787,N_1763);
xnor U1852 (N_1852,N_1793,N_1777);
and U1853 (N_1853,N_1740,N_1739);
nand U1854 (N_1854,N_1757,N_1720);
or U1855 (N_1855,N_1772,N_1779);
nand U1856 (N_1856,N_1784,N_1703);
nor U1857 (N_1857,N_1760,N_1753);
and U1858 (N_1858,N_1757,N_1745);
and U1859 (N_1859,N_1722,N_1727);
and U1860 (N_1860,N_1791,N_1710);
or U1861 (N_1861,N_1751,N_1715);
and U1862 (N_1862,N_1748,N_1702);
nor U1863 (N_1863,N_1723,N_1737);
and U1864 (N_1864,N_1700,N_1717);
and U1865 (N_1865,N_1725,N_1759);
nor U1866 (N_1866,N_1717,N_1715);
nor U1867 (N_1867,N_1700,N_1763);
and U1868 (N_1868,N_1740,N_1786);
nor U1869 (N_1869,N_1700,N_1798);
and U1870 (N_1870,N_1727,N_1758);
nand U1871 (N_1871,N_1701,N_1725);
or U1872 (N_1872,N_1754,N_1749);
xor U1873 (N_1873,N_1731,N_1757);
xnor U1874 (N_1874,N_1776,N_1758);
nand U1875 (N_1875,N_1730,N_1746);
xor U1876 (N_1876,N_1743,N_1783);
nand U1877 (N_1877,N_1762,N_1707);
nand U1878 (N_1878,N_1751,N_1752);
or U1879 (N_1879,N_1705,N_1731);
xnor U1880 (N_1880,N_1733,N_1716);
nand U1881 (N_1881,N_1758,N_1747);
nor U1882 (N_1882,N_1703,N_1721);
nor U1883 (N_1883,N_1752,N_1763);
nor U1884 (N_1884,N_1714,N_1761);
nor U1885 (N_1885,N_1743,N_1750);
or U1886 (N_1886,N_1794,N_1747);
xor U1887 (N_1887,N_1760,N_1752);
xnor U1888 (N_1888,N_1720,N_1735);
nor U1889 (N_1889,N_1733,N_1760);
xor U1890 (N_1890,N_1783,N_1785);
and U1891 (N_1891,N_1762,N_1761);
and U1892 (N_1892,N_1741,N_1738);
nand U1893 (N_1893,N_1708,N_1741);
nand U1894 (N_1894,N_1734,N_1776);
nor U1895 (N_1895,N_1753,N_1702);
nor U1896 (N_1896,N_1753,N_1711);
xnor U1897 (N_1897,N_1726,N_1740);
xnor U1898 (N_1898,N_1727,N_1751);
nand U1899 (N_1899,N_1700,N_1765);
and U1900 (N_1900,N_1882,N_1861);
nand U1901 (N_1901,N_1862,N_1875);
or U1902 (N_1902,N_1838,N_1823);
and U1903 (N_1903,N_1824,N_1820);
nand U1904 (N_1904,N_1804,N_1858);
nor U1905 (N_1905,N_1822,N_1819);
or U1906 (N_1906,N_1869,N_1899);
xnor U1907 (N_1907,N_1857,N_1868);
nand U1908 (N_1908,N_1839,N_1860);
xnor U1909 (N_1909,N_1801,N_1855);
nor U1910 (N_1910,N_1817,N_1851);
or U1911 (N_1911,N_1888,N_1828);
and U1912 (N_1912,N_1848,N_1846);
and U1913 (N_1913,N_1845,N_1864);
nor U1914 (N_1914,N_1863,N_1884);
xor U1915 (N_1915,N_1898,N_1895);
or U1916 (N_1916,N_1853,N_1890);
xor U1917 (N_1917,N_1897,N_1811);
nand U1918 (N_1918,N_1825,N_1810);
xnor U1919 (N_1919,N_1836,N_1800);
xor U1920 (N_1920,N_1808,N_1889);
or U1921 (N_1921,N_1877,N_1805);
or U1922 (N_1922,N_1809,N_1852);
nor U1923 (N_1923,N_1840,N_1854);
xor U1924 (N_1924,N_1886,N_1872);
nor U1925 (N_1925,N_1849,N_1813);
nor U1926 (N_1926,N_1885,N_1803);
or U1927 (N_1927,N_1831,N_1871);
nand U1928 (N_1928,N_1834,N_1850);
xor U1929 (N_1929,N_1835,N_1806);
nand U1930 (N_1930,N_1880,N_1896);
nor U1931 (N_1931,N_1878,N_1879);
nor U1932 (N_1932,N_1826,N_1802);
nand U1933 (N_1933,N_1867,N_1837);
or U1934 (N_1934,N_1842,N_1829);
xor U1935 (N_1935,N_1816,N_1859);
xnor U1936 (N_1936,N_1873,N_1812);
and U1937 (N_1937,N_1815,N_1892);
or U1938 (N_1938,N_1827,N_1844);
and U1939 (N_1939,N_1870,N_1893);
nand U1940 (N_1940,N_1881,N_1818);
xor U1941 (N_1941,N_1866,N_1814);
or U1942 (N_1942,N_1894,N_1883);
or U1943 (N_1943,N_1887,N_1876);
and U1944 (N_1944,N_1833,N_1874);
or U1945 (N_1945,N_1832,N_1847);
nor U1946 (N_1946,N_1821,N_1807);
or U1947 (N_1947,N_1830,N_1865);
xor U1948 (N_1948,N_1856,N_1843);
nor U1949 (N_1949,N_1891,N_1841);
and U1950 (N_1950,N_1896,N_1828);
xor U1951 (N_1951,N_1899,N_1888);
or U1952 (N_1952,N_1803,N_1842);
nand U1953 (N_1953,N_1857,N_1858);
or U1954 (N_1954,N_1835,N_1842);
xor U1955 (N_1955,N_1885,N_1877);
xor U1956 (N_1956,N_1895,N_1867);
nand U1957 (N_1957,N_1854,N_1838);
nor U1958 (N_1958,N_1808,N_1843);
nand U1959 (N_1959,N_1855,N_1876);
nor U1960 (N_1960,N_1845,N_1809);
nor U1961 (N_1961,N_1867,N_1839);
xnor U1962 (N_1962,N_1838,N_1856);
or U1963 (N_1963,N_1848,N_1821);
nand U1964 (N_1964,N_1820,N_1880);
and U1965 (N_1965,N_1825,N_1875);
and U1966 (N_1966,N_1847,N_1867);
or U1967 (N_1967,N_1877,N_1870);
and U1968 (N_1968,N_1868,N_1802);
nor U1969 (N_1969,N_1814,N_1842);
nand U1970 (N_1970,N_1846,N_1875);
or U1971 (N_1971,N_1887,N_1872);
nand U1972 (N_1972,N_1856,N_1887);
or U1973 (N_1973,N_1813,N_1808);
xor U1974 (N_1974,N_1811,N_1812);
nor U1975 (N_1975,N_1897,N_1844);
xor U1976 (N_1976,N_1818,N_1805);
or U1977 (N_1977,N_1844,N_1890);
and U1978 (N_1978,N_1883,N_1882);
and U1979 (N_1979,N_1815,N_1857);
xor U1980 (N_1980,N_1884,N_1854);
or U1981 (N_1981,N_1862,N_1853);
or U1982 (N_1982,N_1851,N_1877);
and U1983 (N_1983,N_1853,N_1814);
xor U1984 (N_1984,N_1896,N_1852);
or U1985 (N_1985,N_1875,N_1828);
or U1986 (N_1986,N_1822,N_1839);
nand U1987 (N_1987,N_1875,N_1826);
or U1988 (N_1988,N_1809,N_1812);
or U1989 (N_1989,N_1832,N_1826);
xor U1990 (N_1990,N_1834,N_1808);
or U1991 (N_1991,N_1852,N_1834);
nor U1992 (N_1992,N_1825,N_1899);
or U1993 (N_1993,N_1800,N_1813);
nor U1994 (N_1994,N_1842,N_1850);
xnor U1995 (N_1995,N_1824,N_1815);
nor U1996 (N_1996,N_1844,N_1878);
nor U1997 (N_1997,N_1854,N_1830);
nor U1998 (N_1998,N_1895,N_1809);
or U1999 (N_1999,N_1860,N_1882);
xnor U2000 (N_2000,N_1938,N_1949);
nor U2001 (N_2001,N_1964,N_1986);
or U2002 (N_2002,N_1961,N_1925);
nor U2003 (N_2003,N_1943,N_1910);
and U2004 (N_2004,N_1977,N_1981);
nor U2005 (N_2005,N_1931,N_1967);
or U2006 (N_2006,N_1979,N_1958);
or U2007 (N_2007,N_1971,N_1996);
and U2008 (N_2008,N_1987,N_1901);
and U2009 (N_2009,N_1907,N_1904);
or U2010 (N_2010,N_1930,N_1980);
nand U2011 (N_2011,N_1911,N_1973);
or U2012 (N_2012,N_1959,N_1997);
and U2013 (N_2013,N_1976,N_1950);
nand U2014 (N_2014,N_1975,N_1966);
nor U2015 (N_2015,N_1955,N_1913);
nand U2016 (N_2016,N_1903,N_1927);
nand U2017 (N_2017,N_1909,N_1928);
xor U2018 (N_2018,N_1933,N_1972);
xnor U2019 (N_2019,N_1999,N_1984);
and U2020 (N_2020,N_1923,N_1952);
xnor U2021 (N_2021,N_1990,N_1926);
xnor U2022 (N_2022,N_1932,N_1939);
nand U2023 (N_2023,N_1991,N_1920);
and U2024 (N_2024,N_1902,N_1936);
and U2025 (N_2025,N_1929,N_1970);
and U2026 (N_2026,N_1962,N_1945);
and U2027 (N_2027,N_1934,N_1942);
nor U2028 (N_2028,N_1935,N_1941);
and U2029 (N_2029,N_1994,N_1916);
nor U2030 (N_2030,N_1906,N_1978);
nand U2031 (N_2031,N_1944,N_1917);
and U2032 (N_2032,N_1946,N_1993);
nor U2033 (N_2033,N_1956,N_1969);
and U2034 (N_2034,N_1951,N_1982);
and U2035 (N_2035,N_1914,N_1948);
or U2036 (N_2036,N_1988,N_1924);
or U2037 (N_2037,N_1992,N_1998);
nor U2038 (N_2038,N_1937,N_1900);
and U2039 (N_2039,N_1947,N_1908);
xor U2040 (N_2040,N_1915,N_1919);
or U2041 (N_2041,N_1983,N_1953);
nor U2042 (N_2042,N_1954,N_1968);
nand U2043 (N_2043,N_1965,N_1940);
or U2044 (N_2044,N_1912,N_1918);
nor U2045 (N_2045,N_1921,N_1905);
and U2046 (N_2046,N_1957,N_1960);
nand U2047 (N_2047,N_1995,N_1963);
or U2048 (N_2048,N_1989,N_1922);
nand U2049 (N_2049,N_1985,N_1974);
xnor U2050 (N_2050,N_1954,N_1955);
xor U2051 (N_2051,N_1989,N_1987);
nand U2052 (N_2052,N_1978,N_1993);
nor U2053 (N_2053,N_1985,N_1969);
or U2054 (N_2054,N_1953,N_1954);
xnor U2055 (N_2055,N_1903,N_1991);
and U2056 (N_2056,N_1922,N_1948);
xnor U2057 (N_2057,N_1998,N_1991);
or U2058 (N_2058,N_1924,N_1987);
xor U2059 (N_2059,N_1921,N_1988);
nor U2060 (N_2060,N_1964,N_1989);
nor U2061 (N_2061,N_1985,N_1904);
and U2062 (N_2062,N_1952,N_1929);
xnor U2063 (N_2063,N_1935,N_1903);
nand U2064 (N_2064,N_1929,N_1994);
nor U2065 (N_2065,N_1990,N_1903);
nor U2066 (N_2066,N_1935,N_1917);
xor U2067 (N_2067,N_1972,N_1939);
nand U2068 (N_2068,N_1999,N_1958);
and U2069 (N_2069,N_1914,N_1980);
or U2070 (N_2070,N_1931,N_1957);
and U2071 (N_2071,N_1977,N_1929);
nand U2072 (N_2072,N_1988,N_1980);
nand U2073 (N_2073,N_1965,N_1946);
xnor U2074 (N_2074,N_1913,N_1968);
xnor U2075 (N_2075,N_1912,N_1985);
nor U2076 (N_2076,N_1990,N_1975);
or U2077 (N_2077,N_1934,N_1945);
nand U2078 (N_2078,N_1970,N_1990);
nand U2079 (N_2079,N_1954,N_1988);
xnor U2080 (N_2080,N_1999,N_1923);
nand U2081 (N_2081,N_1960,N_1908);
xnor U2082 (N_2082,N_1989,N_1961);
or U2083 (N_2083,N_1954,N_1978);
xor U2084 (N_2084,N_1969,N_1918);
nand U2085 (N_2085,N_1973,N_1905);
nor U2086 (N_2086,N_1902,N_1997);
xor U2087 (N_2087,N_1965,N_1950);
nor U2088 (N_2088,N_1933,N_1950);
and U2089 (N_2089,N_1988,N_1968);
xor U2090 (N_2090,N_1935,N_1956);
xnor U2091 (N_2091,N_1991,N_1965);
nor U2092 (N_2092,N_1981,N_1947);
xnor U2093 (N_2093,N_1976,N_1974);
nand U2094 (N_2094,N_1913,N_1961);
and U2095 (N_2095,N_1934,N_1925);
and U2096 (N_2096,N_1973,N_1961);
nor U2097 (N_2097,N_1908,N_1980);
and U2098 (N_2098,N_1982,N_1954);
nand U2099 (N_2099,N_1944,N_1953);
nor U2100 (N_2100,N_2058,N_2076);
or U2101 (N_2101,N_2068,N_2046);
or U2102 (N_2102,N_2002,N_2008);
nand U2103 (N_2103,N_2088,N_2092);
nor U2104 (N_2104,N_2000,N_2014);
xor U2105 (N_2105,N_2079,N_2077);
nand U2106 (N_2106,N_2063,N_2034);
nor U2107 (N_2107,N_2031,N_2074);
xnor U2108 (N_2108,N_2015,N_2086);
xor U2109 (N_2109,N_2065,N_2051);
or U2110 (N_2110,N_2085,N_2026);
xor U2111 (N_2111,N_2061,N_2030);
xnor U2112 (N_2112,N_2055,N_2094);
or U2113 (N_2113,N_2072,N_2042);
nand U2114 (N_2114,N_2048,N_2007);
nor U2115 (N_2115,N_2067,N_2043);
nor U2116 (N_2116,N_2040,N_2084);
nand U2117 (N_2117,N_2097,N_2064);
nor U2118 (N_2118,N_2047,N_2090);
nor U2119 (N_2119,N_2075,N_2069);
nor U2120 (N_2120,N_2022,N_2087);
xor U2121 (N_2121,N_2095,N_2033);
or U2122 (N_2122,N_2004,N_2078);
and U2123 (N_2123,N_2039,N_2093);
xor U2124 (N_2124,N_2081,N_2021);
or U2125 (N_2125,N_2049,N_2013);
or U2126 (N_2126,N_2035,N_2003);
or U2127 (N_2127,N_2037,N_2032);
nor U2128 (N_2128,N_2073,N_2062);
or U2129 (N_2129,N_2044,N_2091);
nand U2130 (N_2130,N_2029,N_2019);
nand U2131 (N_2131,N_2050,N_2010);
xor U2132 (N_2132,N_2012,N_2009);
nand U2133 (N_2133,N_2099,N_2083);
and U2134 (N_2134,N_2070,N_2001);
xor U2135 (N_2135,N_2027,N_2082);
nand U2136 (N_2136,N_2016,N_2071);
xnor U2137 (N_2137,N_2036,N_2098);
xor U2138 (N_2138,N_2011,N_2024);
and U2139 (N_2139,N_2025,N_2038);
and U2140 (N_2140,N_2018,N_2089);
or U2141 (N_2141,N_2096,N_2060);
or U2142 (N_2142,N_2052,N_2066);
and U2143 (N_2143,N_2041,N_2020);
nand U2144 (N_2144,N_2005,N_2017);
nand U2145 (N_2145,N_2059,N_2080);
xnor U2146 (N_2146,N_2045,N_2056);
or U2147 (N_2147,N_2054,N_2023);
nor U2148 (N_2148,N_2057,N_2006);
and U2149 (N_2149,N_2053,N_2028);
and U2150 (N_2150,N_2053,N_2049);
and U2151 (N_2151,N_2096,N_2080);
nor U2152 (N_2152,N_2083,N_2063);
nand U2153 (N_2153,N_2077,N_2050);
nor U2154 (N_2154,N_2079,N_2074);
nand U2155 (N_2155,N_2092,N_2078);
and U2156 (N_2156,N_2097,N_2062);
nand U2157 (N_2157,N_2070,N_2022);
and U2158 (N_2158,N_2040,N_2019);
nand U2159 (N_2159,N_2049,N_2006);
nor U2160 (N_2160,N_2044,N_2045);
nor U2161 (N_2161,N_2025,N_2019);
xor U2162 (N_2162,N_2090,N_2053);
and U2163 (N_2163,N_2022,N_2057);
nand U2164 (N_2164,N_2086,N_2065);
nand U2165 (N_2165,N_2036,N_2034);
or U2166 (N_2166,N_2062,N_2012);
nand U2167 (N_2167,N_2007,N_2078);
nand U2168 (N_2168,N_2095,N_2016);
xnor U2169 (N_2169,N_2015,N_2002);
or U2170 (N_2170,N_2058,N_2072);
or U2171 (N_2171,N_2048,N_2024);
xnor U2172 (N_2172,N_2014,N_2022);
and U2173 (N_2173,N_2093,N_2060);
and U2174 (N_2174,N_2030,N_2056);
or U2175 (N_2175,N_2073,N_2059);
nor U2176 (N_2176,N_2048,N_2021);
nor U2177 (N_2177,N_2097,N_2080);
nand U2178 (N_2178,N_2025,N_2043);
and U2179 (N_2179,N_2055,N_2013);
nand U2180 (N_2180,N_2046,N_2069);
xor U2181 (N_2181,N_2053,N_2041);
xor U2182 (N_2182,N_2081,N_2099);
and U2183 (N_2183,N_2074,N_2056);
nor U2184 (N_2184,N_2053,N_2075);
xor U2185 (N_2185,N_2084,N_2092);
nor U2186 (N_2186,N_2011,N_2029);
xnor U2187 (N_2187,N_2040,N_2035);
or U2188 (N_2188,N_2005,N_2085);
xnor U2189 (N_2189,N_2002,N_2048);
and U2190 (N_2190,N_2084,N_2067);
xor U2191 (N_2191,N_2040,N_2029);
xor U2192 (N_2192,N_2035,N_2096);
xor U2193 (N_2193,N_2004,N_2088);
nand U2194 (N_2194,N_2049,N_2034);
nor U2195 (N_2195,N_2015,N_2052);
or U2196 (N_2196,N_2026,N_2001);
nand U2197 (N_2197,N_2090,N_2096);
nor U2198 (N_2198,N_2096,N_2038);
and U2199 (N_2199,N_2025,N_2048);
xnor U2200 (N_2200,N_2151,N_2193);
nand U2201 (N_2201,N_2172,N_2167);
xnor U2202 (N_2202,N_2181,N_2187);
xor U2203 (N_2203,N_2109,N_2182);
xnor U2204 (N_2204,N_2122,N_2143);
nand U2205 (N_2205,N_2178,N_2190);
nor U2206 (N_2206,N_2173,N_2161);
or U2207 (N_2207,N_2148,N_2123);
nand U2208 (N_2208,N_2136,N_2170);
nand U2209 (N_2209,N_2121,N_2105);
or U2210 (N_2210,N_2176,N_2150);
nor U2211 (N_2211,N_2189,N_2169);
nand U2212 (N_2212,N_2112,N_2164);
xor U2213 (N_2213,N_2179,N_2101);
xor U2214 (N_2214,N_2126,N_2145);
nor U2215 (N_2215,N_2129,N_2132);
and U2216 (N_2216,N_2199,N_2130);
xnor U2217 (N_2217,N_2156,N_2183);
and U2218 (N_2218,N_2124,N_2120);
nand U2219 (N_2219,N_2157,N_2144);
and U2220 (N_2220,N_2117,N_2175);
or U2221 (N_2221,N_2133,N_2106);
or U2222 (N_2222,N_2163,N_2196);
and U2223 (N_2223,N_2100,N_2166);
or U2224 (N_2224,N_2110,N_2138);
nor U2225 (N_2225,N_2174,N_2191);
and U2226 (N_2226,N_2168,N_2195);
nand U2227 (N_2227,N_2188,N_2140);
nand U2228 (N_2228,N_2131,N_2116);
nand U2229 (N_2229,N_2160,N_2111);
or U2230 (N_2230,N_2184,N_2108);
or U2231 (N_2231,N_2162,N_2142);
nor U2232 (N_2232,N_2113,N_2127);
or U2233 (N_2233,N_2139,N_2134);
or U2234 (N_2234,N_2192,N_2165);
xnor U2235 (N_2235,N_2158,N_2186);
nand U2236 (N_2236,N_2180,N_2118);
and U2237 (N_2237,N_2104,N_2159);
nand U2238 (N_2238,N_2177,N_2115);
or U2239 (N_2239,N_2198,N_2135);
xor U2240 (N_2240,N_2128,N_2153);
xnor U2241 (N_2241,N_2137,N_2102);
nor U2242 (N_2242,N_2154,N_2103);
xor U2243 (N_2243,N_2194,N_2149);
xnor U2244 (N_2244,N_2146,N_2171);
nand U2245 (N_2245,N_2185,N_2152);
xor U2246 (N_2246,N_2125,N_2155);
and U2247 (N_2247,N_2119,N_2141);
nand U2248 (N_2248,N_2147,N_2107);
or U2249 (N_2249,N_2197,N_2114);
nand U2250 (N_2250,N_2102,N_2115);
nor U2251 (N_2251,N_2140,N_2161);
or U2252 (N_2252,N_2135,N_2123);
and U2253 (N_2253,N_2179,N_2119);
nor U2254 (N_2254,N_2158,N_2115);
and U2255 (N_2255,N_2126,N_2147);
nand U2256 (N_2256,N_2130,N_2107);
and U2257 (N_2257,N_2118,N_2125);
nand U2258 (N_2258,N_2129,N_2166);
or U2259 (N_2259,N_2137,N_2186);
nor U2260 (N_2260,N_2101,N_2132);
and U2261 (N_2261,N_2196,N_2198);
xnor U2262 (N_2262,N_2143,N_2195);
or U2263 (N_2263,N_2127,N_2129);
nand U2264 (N_2264,N_2141,N_2112);
or U2265 (N_2265,N_2134,N_2159);
nor U2266 (N_2266,N_2172,N_2163);
or U2267 (N_2267,N_2188,N_2128);
or U2268 (N_2268,N_2150,N_2126);
xnor U2269 (N_2269,N_2161,N_2188);
xor U2270 (N_2270,N_2178,N_2116);
nand U2271 (N_2271,N_2168,N_2143);
nor U2272 (N_2272,N_2188,N_2172);
and U2273 (N_2273,N_2142,N_2182);
nand U2274 (N_2274,N_2145,N_2184);
nor U2275 (N_2275,N_2193,N_2120);
or U2276 (N_2276,N_2162,N_2143);
or U2277 (N_2277,N_2191,N_2136);
or U2278 (N_2278,N_2181,N_2152);
or U2279 (N_2279,N_2194,N_2190);
nor U2280 (N_2280,N_2187,N_2124);
and U2281 (N_2281,N_2118,N_2193);
or U2282 (N_2282,N_2132,N_2155);
or U2283 (N_2283,N_2185,N_2155);
and U2284 (N_2284,N_2194,N_2137);
xnor U2285 (N_2285,N_2181,N_2132);
nand U2286 (N_2286,N_2174,N_2149);
nand U2287 (N_2287,N_2174,N_2115);
nor U2288 (N_2288,N_2150,N_2189);
or U2289 (N_2289,N_2179,N_2121);
or U2290 (N_2290,N_2143,N_2152);
or U2291 (N_2291,N_2169,N_2190);
or U2292 (N_2292,N_2189,N_2151);
nand U2293 (N_2293,N_2156,N_2103);
and U2294 (N_2294,N_2147,N_2184);
and U2295 (N_2295,N_2120,N_2190);
xnor U2296 (N_2296,N_2101,N_2162);
xnor U2297 (N_2297,N_2121,N_2196);
nand U2298 (N_2298,N_2161,N_2184);
or U2299 (N_2299,N_2100,N_2130);
nor U2300 (N_2300,N_2264,N_2260);
xor U2301 (N_2301,N_2276,N_2233);
and U2302 (N_2302,N_2299,N_2250);
and U2303 (N_2303,N_2211,N_2222);
xnor U2304 (N_2304,N_2247,N_2218);
and U2305 (N_2305,N_2283,N_2279);
nand U2306 (N_2306,N_2241,N_2293);
nor U2307 (N_2307,N_2217,N_2243);
nor U2308 (N_2308,N_2280,N_2263);
nor U2309 (N_2309,N_2288,N_2226);
or U2310 (N_2310,N_2254,N_2207);
or U2311 (N_2311,N_2261,N_2285);
or U2312 (N_2312,N_2215,N_2290);
or U2313 (N_2313,N_2259,N_2213);
and U2314 (N_2314,N_2229,N_2271);
xor U2315 (N_2315,N_2219,N_2227);
and U2316 (N_2316,N_2231,N_2204);
and U2317 (N_2317,N_2224,N_2291);
and U2318 (N_2318,N_2235,N_2223);
and U2319 (N_2319,N_2277,N_2282);
xnor U2320 (N_2320,N_2286,N_2203);
and U2321 (N_2321,N_2267,N_2240);
and U2322 (N_2322,N_2232,N_2274);
nor U2323 (N_2323,N_2273,N_2257);
nand U2324 (N_2324,N_2214,N_2230);
nor U2325 (N_2325,N_2201,N_2256);
nor U2326 (N_2326,N_2200,N_2294);
nor U2327 (N_2327,N_2298,N_2252);
or U2328 (N_2328,N_2202,N_2237);
nand U2329 (N_2329,N_2284,N_2212);
nand U2330 (N_2330,N_2205,N_2249);
nand U2331 (N_2331,N_2281,N_2295);
or U2332 (N_2332,N_2278,N_2251);
and U2333 (N_2333,N_2221,N_2228);
and U2334 (N_2334,N_2236,N_2253);
nand U2335 (N_2335,N_2225,N_2289);
nand U2336 (N_2336,N_2268,N_2220);
nor U2337 (N_2337,N_2244,N_2269);
or U2338 (N_2338,N_2296,N_2209);
and U2339 (N_2339,N_2265,N_2292);
and U2340 (N_2340,N_2297,N_2248);
xnor U2341 (N_2341,N_2255,N_2238);
nor U2342 (N_2342,N_2287,N_2262);
and U2343 (N_2343,N_2206,N_2266);
nor U2344 (N_2344,N_2216,N_2245);
xnor U2345 (N_2345,N_2210,N_2272);
nand U2346 (N_2346,N_2242,N_2258);
nand U2347 (N_2347,N_2234,N_2239);
and U2348 (N_2348,N_2246,N_2270);
xnor U2349 (N_2349,N_2275,N_2208);
nor U2350 (N_2350,N_2251,N_2222);
nand U2351 (N_2351,N_2297,N_2296);
or U2352 (N_2352,N_2247,N_2221);
nor U2353 (N_2353,N_2233,N_2210);
or U2354 (N_2354,N_2238,N_2231);
nand U2355 (N_2355,N_2250,N_2298);
nand U2356 (N_2356,N_2272,N_2205);
or U2357 (N_2357,N_2254,N_2267);
nand U2358 (N_2358,N_2215,N_2237);
xor U2359 (N_2359,N_2299,N_2242);
or U2360 (N_2360,N_2276,N_2268);
and U2361 (N_2361,N_2259,N_2206);
and U2362 (N_2362,N_2235,N_2224);
nor U2363 (N_2363,N_2205,N_2217);
nor U2364 (N_2364,N_2226,N_2238);
nand U2365 (N_2365,N_2211,N_2203);
and U2366 (N_2366,N_2219,N_2286);
nor U2367 (N_2367,N_2287,N_2249);
nor U2368 (N_2368,N_2201,N_2253);
xnor U2369 (N_2369,N_2211,N_2291);
xnor U2370 (N_2370,N_2209,N_2215);
nand U2371 (N_2371,N_2225,N_2295);
or U2372 (N_2372,N_2283,N_2271);
nor U2373 (N_2373,N_2201,N_2224);
nor U2374 (N_2374,N_2267,N_2234);
or U2375 (N_2375,N_2280,N_2292);
and U2376 (N_2376,N_2269,N_2208);
and U2377 (N_2377,N_2244,N_2234);
nand U2378 (N_2378,N_2229,N_2270);
and U2379 (N_2379,N_2259,N_2204);
and U2380 (N_2380,N_2246,N_2283);
nand U2381 (N_2381,N_2290,N_2277);
xor U2382 (N_2382,N_2273,N_2205);
and U2383 (N_2383,N_2205,N_2246);
nor U2384 (N_2384,N_2241,N_2216);
xnor U2385 (N_2385,N_2291,N_2241);
xnor U2386 (N_2386,N_2275,N_2268);
and U2387 (N_2387,N_2234,N_2299);
and U2388 (N_2388,N_2242,N_2235);
or U2389 (N_2389,N_2252,N_2289);
xor U2390 (N_2390,N_2297,N_2242);
or U2391 (N_2391,N_2256,N_2203);
xor U2392 (N_2392,N_2227,N_2203);
or U2393 (N_2393,N_2223,N_2273);
or U2394 (N_2394,N_2245,N_2274);
xor U2395 (N_2395,N_2294,N_2268);
nand U2396 (N_2396,N_2234,N_2264);
and U2397 (N_2397,N_2284,N_2261);
nand U2398 (N_2398,N_2280,N_2288);
nand U2399 (N_2399,N_2235,N_2204);
or U2400 (N_2400,N_2313,N_2315);
nand U2401 (N_2401,N_2346,N_2379);
nand U2402 (N_2402,N_2368,N_2345);
xor U2403 (N_2403,N_2356,N_2318);
nand U2404 (N_2404,N_2386,N_2344);
nor U2405 (N_2405,N_2321,N_2335);
nor U2406 (N_2406,N_2337,N_2389);
nor U2407 (N_2407,N_2308,N_2365);
xor U2408 (N_2408,N_2314,N_2397);
nand U2409 (N_2409,N_2363,N_2347);
and U2410 (N_2410,N_2310,N_2342);
nand U2411 (N_2411,N_2305,N_2327);
nand U2412 (N_2412,N_2361,N_2384);
nor U2413 (N_2413,N_2392,N_2309);
or U2414 (N_2414,N_2317,N_2353);
nor U2415 (N_2415,N_2364,N_2352);
or U2416 (N_2416,N_2398,N_2326);
nand U2417 (N_2417,N_2330,N_2380);
nor U2418 (N_2418,N_2374,N_2362);
xnor U2419 (N_2419,N_2329,N_2372);
xnor U2420 (N_2420,N_2311,N_2385);
and U2421 (N_2421,N_2307,N_2328);
or U2422 (N_2422,N_2358,N_2304);
nand U2423 (N_2423,N_2332,N_2338);
or U2424 (N_2424,N_2333,N_2323);
nor U2425 (N_2425,N_2302,N_2360);
or U2426 (N_2426,N_2391,N_2322);
or U2427 (N_2427,N_2339,N_2301);
and U2428 (N_2428,N_2319,N_2331);
and U2429 (N_2429,N_2343,N_2367);
xor U2430 (N_2430,N_2348,N_2394);
or U2431 (N_2431,N_2354,N_2383);
and U2432 (N_2432,N_2350,N_2371);
nor U2433 (N_2433,N_2366,N_2312);
and U2434 (N_2434,N_2351,N_2390);
xor U2435 (N_2435,N_2316,N_2306);
xor U2436 (N_2436,N_2396,N_2375);
nor U2437 (N_2437,N_2370,N_2359);
and U2438 (N_2438,N_2393,N_2377);
or U2439 (N_2439,N_2325,N_2376);
nand U2440 (N_2440,N_2300,N_2349);
xor U2441 (N_2441,N_2382,N_2336);
or U2442 (N_2442,N_2320,N_2355);
xor U2443 (N_2443,N_2378,N_2357);
xor U2444 (N_2444,N_2324,N_2395);
and U2445 (N_2445,N_2399,N_2373);
xor U2446 (N_2446,N_2387,N_2334);
or U2447 (N_2447,N_2388,N_2341);
xor U2448 (N_2448,N_2369,N_2303);
and U2449 (N_2449,N_2381,N_2340);
and U2450 (N_2450,N_2367,N_2352);
nor U2451 (N_2451,N_2345,N_2365);
and U2452 (N_2452,N_2323,N_2327);
nor U2453 (N_2453,N_2390,N_2388);
or U2454 (N_2454,N_2382,N_2361);
or U2455 (N_2455,N_2397,N_2396);
nor U2456 (N_2456,N_2337,N_2351);
or U2457 (N_2457,N_2363,N_2309);
and U2458 (N_2458,N_2367,N_2378);
nor U2459 (N_2459,N_2308,N_2306);
or U2460 (N_2460,N_2326,N_2343);
nor U2461 (N_2461,N_2377,N_2358);
or U2462 (N_2462,N_2366,N_2387);
or U2463 (N_2463,N_2365,N_2355);
xor U2464 (N_2464,N_2326,N_2381);
nand U2465 (N_2465,N_2391,N_2386);
and U2466 (N_2466,N_2337,N_2304);
xor U2467 (N_2467,N_2381,N_2364);
nor U2468 (N_2468,N_2374,N_2303);
nand U2469 (N_2469,N_2396,N_2303);
xnor U2470 (N_2470,N_2346,N_2373);
and U2471 (N_2471,N_2372,N_2383);
nand U2472 (N_2472,N_2313,N_2393);
nor U2473 (N_2473,N_2354,N_2323);
nand U2474 (N_2474,N_2377,N_2334);
and U2475 (N_2475,N_2344,N_2356);
xnor U2476 (N_2476,N_2315,N_2302);
and U2477 (N_2477,N_2355,N_2366);
nor U2478 (N_2478,N_2376,N_2378);
or U2479 (N_2479,N_2368,N_2367);
xnor U2480 (N_2480,N_2398,N_2382);
nor U2481 (N_2481,N_2345,N_2361);
or U2482 (N_2482,N_2378,N_2366);
nand U2483 (N_2483,N_2359,N_2330);
xor U2484 (N_2484,N_2311,N_2365);
nor U2485 (N_2485,N_2367,N_2335);
nand U2486 (N_2486,N_2359,N_2347);
or U2487 (N_2487,N_2394,N_2364);
xnor U2488 (N_2488,N_2340,N_2376);
or U2489 (N_2489,N_2327,N_2370);
xnor U2490 (N_2490,N_2345,N_2320);
xnor U2491 (N_2491,N_2359,N_2381);
and U2492 (N_2492,N_2357,N_2304);
nand U2493 (N_2493,N_2365,N_2351);
nor U2494 (N_2494,N_2315,N_2324);
and U2495 (N_2495,N_2348,N_2300);
nand U2496 (N_2496,N_2318,N_2309);
nor U2497 (N_2497,N_2348,N_2310);
xor U2498 (N_2498,N_2388,N_2366);
xor U2499 (N_2499,N_2386,N_2371);
or U2500 (N_2500,N_2489,N_2474);
nand U2501 (N_2501,N_2496,N_2476);
nor U2502 (N_2502,N_2462,N_2475);
nor U2503 (N_2503,N_2408,N_2486);
nand U2504 (N_2504,N_2451,N_2491);
nand U2505 (N_2505,N_2416,N_2469);
xnor U2506 (N_2506,N_2472,N_2498);
xor U2507 (N_2507,N_2425,N_2490);
and U2508 (N_2508,N_2485,N_2477);
nor U2509 (N_2509,N_2484,N_2463);
and U2510 (N_2510,N_2403,N_2483);
or U2511 (N_2511,N_2481,N_2423);
nand U2512 (N_2512,N_2420,N_2443);
nand U2513 (N_2513,N_2402,N_2410);
xnor U2514 (N_2514,N_2428,N_2455);
xnor U2515 (N_2515,N_2406,N_2440);
or U2516 (N_2516,N_2456,N_2465);
or U2517 (N_2517,N_2473,N_2479);
or U2518 (N_2518,N_2409,N_2436);
or U2519 (N_2519,N_2494,N_2499);
nand U2520 (N_2520,N_2422,N_2431);
nand U2521 (N_2521,N_2411,N_2487);
xor U2522 (N_2522,N_2464,N_2450);
and U2523 (N_2523,N_2407,N_2445);
xor U2524 (N_2524,N_2497,N_2400);
nor U2525 (N_2525,N_2466,N_2429);
nor U2526 (N_2526,N_2424,N_2433);
xor U2527 (N_2527,N_2453,N_2404);
and U2528 (N_2528,N_2467,N_2492);
or U2529 (N_2529,N_2418,N_2495);
nor U2530 (N_2530,N_2401,N_2435);
and U2531 (N_2531,N_2441,N_2430);
xnor U2532 (N_2532,N_2405,N_2426);
or U2533 (N_2533,N_2412,N_2461);
nand U2534 (N_2534,N_2470,N_2421);
and U2535 (N_2535,N_2471,N_2413);
nand U2536 (N_2536,N_2468,N_2458);
or U2537 (N_2537,N_2419,N_2448);
nand U2538 (N_2538,N_2442,N_2460);
xnor U2539 (N_2539,N_2493,N_2459);
xnor U2540 (N_2540,N_2482,N_2452);
and U2541 (N_2541,N_2454,N_2444);
or U2542 (N_2542,N_2480,N_2478);
and U2543 (N_2543,N_2432,N_2439);
and U2544 (N_2544,N_2417,N_2414);
nand U2545 (N_2545,N_2457,N_2449);
nor U2546 (N_2546,N_2447,N_2434);
nor U2547 (N_2547,N_2427,N_2488);
and U2548 (N_2548,N_2446,N_2437);
or U2549 (N_2549,N_2438,N_2415);
and U2550 (N_2550,N_2413,N_2420);
xnor U2551 (N_2551,N_2494,N_2464);
nand U2552 (N_2552,N_2400,N_2449);
nand U2553 (N_2553,N_2403,N_2463);
nor U2554 (N_2554,N_2490,N_2476);
nand U2555 (N_2555,N_2416,N_2455);
or U2556 (N_2556,N_2450,N_2428);
nor U2557 (N_2557,N_2425,N_2499);
or U2558 (N_2558,N_2493,N_2435);
xor U2559 (N_2559,N_2487,N_2496);
nor U2560 (N_2560,N_2461,N_2410);
nand U2561 (N_2561,N_2433,N_2473);
nor U2562 (N_2562,N_2467,N_2406);
or U2563 (N_2563,N_2403,N_2417);
nor U2564 (N_2564,N_2472,N_2410);
xor U2565 (N_2565,N_2481,N_2483);
nand U2566 (N_2566,N_2442,N_2441);
nand U2567 (N_2567,N_2497,N_2408);
xnor U2568 (N_2568,N_2466,N_2483);
nand U2569 (N_2569,N_2494,N_2470);
nand U2570 (N_2570,N_2480,N_2435);
and U2571 (N_2571,N_2460,N_2450);
or U2572 (N_2572,N_2471,N_2420);
nand U2573 (N_2573,N_2457,N_2458);
or U2574 (N_2574,N_2472,N_2466);
nand U2575 (N_2575,N_2493,N_2431);
nand U2576 (N_2576,N_2442,N_2469);
xor U2577 (N_2577,N_2479,N_2477);
or U2578 (N_2578,N_2490,N_2435);
xnor U2579 (N_2579,N_2485,N_2463);
or U2580 (N_2580,N_2412,N_2411);
nand U2581 (N_2581,N_2451,N_2407);
nand U2582 (N_2582,N_2417,N_2419);
nand U2583 (N_2583,N_2411,N_2493);
xor U2584 (N_2584,N_2453,N_2493);
nand U2585 (N_2585,N_2472,N_2461);
and U2586 (N_2586,N_2422,N_2480);
nor U2587 (N_2587,N_2411,N_2497);
nand U2588 (N_2588,N_2458,N_2428);
or U2589 (N_2589,N_2426,N_2442);
xnor U2590 (N_2590,N_2478,N_2420);
or U2591 (N_2591,N_2492,N_2429);
nor U2592 (N_2592,N_2458,N_2459);
or U2593 (N_2593,N_2427,N_2411);
or U2594 (N_2594,N_2434,N_2471);
xor U2595 (N_2595,N_2498,N_2403);
or U2596 (N_2596,N_2416,N_2479);
nor U2597 (N_2597,N_2420,N_2451);
xor U2598 (N_2598,N_2454,N_2469);
nand U2599 (N_2599,N_2404,N_2497);
and U2600 (N_2600,N_2568,N_2572);
nor U2601 (N_2601,N_2569,N_2592);
nand U2602 (N_2602,N_2594,N_2528);
or U2603 (N_2603,N_2520,N_2586);
nand U2604 (N_2604,N_2553,N_2554);
or U2605 (N_2605,N_2575,N_2567);
or U2606 (N_2606,N_2580,N_2534);
nand U2607 (N_2607,N_2555,N_2591);
nand U2608 (N_2608,N_2563,N_2544);
nor U2609 (N_2609,N_2570,N_2518);
and U2610 (N_2610,N_2542,N_2502);
nor U2611 (N_2611,N_2516,N_2582);
xor U2612 (N_2612,N_2585,N_2579);
or U2613 (N_2613,N_2538,N_2515);
and U2614 (N_2614,N_2505,N_2501);
nor U2615 (N_2615,N_2548,N_2531);
nor U2616 (N_2616,N_2540,N_2512);
or U2617 (N_2617,N_2551,N_2508);
or U2618 (N_2618,N_2509,N_2577);
nor U2619 (N_2619,N_2561,N_2549);
nand U2620 (N_2620,N_2559,N_2574);
and U2621 (N_2621,N_2526,N_2584);
nand U2622 (N_2622,N_2557,N_2535);
and U2623 (N_2623,N_2500,N_2504);
nor U2624 (N_2624,N_2599,N_2545);
xnor U2625 (N_2625,N_2558,N_2524);
nor U2626 (N_2626,N_2598,N_2552);
nand U2627 (N_2627,N_2506,N_2587);
nor U2628 (N_2628,N_2543,N_2550);
nand U2629 (N_2629,N_2547,N_2573);
or U2630 (N_2630,N_2503,N_2522);
and U2631 (N_2631,N_2593,N_2578);
or U2632 (N_2632,N_2536,N_2541);
xnor U2633 (N_2633,N_2589,N_2537);
or U2634 (N_2634,N_2533,N_2560);
xor U2635 (N_2635,N_2562,N_2511);
xor U2636 (N_2636,N_2596,N_2525);
or U2637 (N_2637,N_2595,N_2565);
xnor U2638 (N_2638,N_2510,N_2517);
nor U2639 (N_2639,N_2566,N_2521);
and U2640 (N_2640,N_2581,N_2527);
or U2641 (N_2641,N_2539,N_2529);
xor U2642 (N_2642,N_2546,N_2530);
xnor U2643 (N_2643,N_2576,N_2507);
nand U2644 (N_2644,N_2523,N_2590);
and U2645 (N_2645,N_2564,N_2571);
xnor U2646 (N_2646,N_2532,N_2514);
nand U2647 (N_2647,N_2597,N_2513);
nand U2648 (N_2648,N_2556,N_2519);
nor U2649 (N_2649,N_2588,N_2583);
and U2650 (N_2650,N_2557,N_2514);
nand U2651 (N_2651,N_2551,N_2596);
and U2652 (N_2652,N_2545,N_2524);
xor U2653 (N_2653,N_2577,N_2545);
nand U2654 (N_2654,N_2539,N_2511);
nand U2655 (N_2655,N_2528,N_2553);
and U2656 (N_2656,N_2550,N_2568);
nand U2657 (N_2657,N_2552,N_2577);
and U2658 (N_2658,N_2595,N_2548);
and U2659 (N_2659,N_2575,N_2580);
or U2660 (N_2660,N_2572,N_2564);
and U2661 (N_2661,N_2511,N_2593);
or U2662 (N_2662,N_2546,N_2512);
nand U2663 (N_2663,N_2511,N_2525);
and U2664 (N_2664,N_2520,N_2522);
or U2665 (N_2665,N_2598,N_2507);
and U2666 (N_2666,N_2508,N_2565);
and U2667 (N_2667,N_2568,N_2577);
or U2668 (N_2668,N_2595,N_2578);
xnor U2669 (N_2669,N_2569,N_2580);
nor U2670 (N_2670,N_2599,N_2559);
nor U2671 (N_2671,N_2541,N_2564);
and U2672 (N_2672,N_2503,N_2543);
xnor U2673 (N_2673,N_2503,N_2512);
nand U2674 (N_2674,N_2551,N_2588);
xor U2675 (N_2675,N_2542,N_2561);
or U2676 (N_2676,N_2547,N_2524);
or U2677 (N_2677,N_2510,N_2579);
nand U2678 (N_2678,N_2512,N_2572);
nand U2679 (N_2679,N_2514,N_2525);
nor U2680 (N_2680,N_2520,N_2571);
nand U2681 (N_2681,N_2582,N_2548);
nor U2682 (N_2682,N_2530,N_2543);
nor U2683 (N_2683,N_2558,N_2551);
xnor U2684 (N_2684,N_2552,N_2511);
and U2685 (N_2685,N_2522,N_2563);
xor U2686 (N_2686,N_2577,N_2587);
nor U2687 (N_2687,N_2552,N_2531);
or U2688 (N_2688,N_2514,N_2524);
nand U2689 (N_2689,N_2599,N_2504);
nor U2690 (N_2690,N_2535,N_2545);
xor U2691 (N_2691,N_2530,N_2519);
nand U2692 (N_2692,N_2559,N_2580);
and U2693 (N_2693,N_2558,N_2552);
nand U2694 (N_2694,N_2511,N_2561);
and U2695 (N_2695,N_2588,N_2506);
nor U2696 (N_2696,N_2507,N_2500);
xnor U2697 (N_2697,N_2538,N_2580);
nand U2698 (N_2698,N_2539,N_2544);
xor U2699 (N_2699,N_2577,N_2512);
or U2700 (N_2700,N_2625,N_2656);
or U2701 (N_2701,N_2604,N_2694);
and U2702 (N_2702,N_2675,N_2678);
and U2703 (N_2703,N_2697,N_2676);
nand U2704 (N_2704,N_2651,N_2617);
xnor U2705 (N_2705,N_2623,N_2627);
or U2706 (N_2706,N_2612,N_2693);
xor U2707 (N_2707,N_2618,N_2661);
nor U2708 (N_2708,N_2631,N_2696);
and U2709 (N_2709,N_2664,N_2674);
nand U2710 (N_2710,N_2621,N_2673);
xnor U2711 (N_2711,N_2633,N_2607);
and U2712 (N_2712,N_2622,N_2648);
nand U2713 (N_2713,N_2605,N_2616);
nand U2714 (N_2714,N_2657,N_2613);
nand U2715 (N_2715,N_2681,N_2644);
nand U2716 (N_2716,N_2615,N_2635);
and U2717 (N_2717,N_2611,N_2677);
or U2718 (N_2718,N_2649,N_2610);
nor U2719 (N_2719,N_2655,N_2663);
or U2720 (N_2720,N_2640,N_2667);
nand U2721 (N_2721,N_2628,N_2669);
nand U2722 (N_2722,N_2683,N_2636);
or U2723 (N_2723,N_2698,N_2629);
and U2724 (N_2724,N_2659,N_2603);
or U2725 (N_2725,N_2614,N_2642);
and U2726 (N_2726,N_2684,N_2679);
or U2727 (N_2727,N_2699,N_2637);
and U2728 (N_2728,N_2602,N_2634);
nand U2729 (N_2729,N_2639,N_2650);
and U2730 (N_2730,N_2660,N_2666);
and U2731 (N_2731,N_2658,N_2695);
nor U2732 (N_2732,N_2665,N_2626);
and U2733 (N_2733,N_2671,N_2662);
and U2734 (N_2734,N_2672,N_2686);
or U2735 (N_2735,N_2630,N_2653);
or U2736 (N_2736,N_2647,N_2620);
nor U2737 (N_2737,N_2643,N_2609);
nand U2738 (N_2738,N_2687,N_2654);
and U2739 (N_2739,N_2688,N_2606);
or U2740 (N_2740,N_2619,N_2624);
xnor U2741 (N_2741,N_2680,N_2601);
or U2742 (N_2742,N_2646,N_2641);
and U2743 (N_2743,N_2689,N_2632);
xor U2744 (N_2744,N_2690,N_2682);
nor U2745 (N_2745,N_2600,N_2645);
or U2746 (N_2746,N_2670,N_2685);
nand U2747 (N_2747,N_2638,N_2608);
xnor U2748 (N_2748,N_2652,N_2668);
and U2749 (N_2749,N_2692,N_2691);
nor U2750 (N_2750,N_2679,N_2699);
and U2751 (N_2751,N_2605,N_2606);
nor U2752 (N_2752,N_2664,N_2655);
nor U2753 (N_2753,N_2646,N_2623);
nor U2754 (N_2754,N_2672,N_2627);
and U2755 (N_2755,N_2645,N_2630);
nor U2756 (N_2756,N_2685,N_2634);
xor U2757 (N_2757,N_2637,N_2685);
nand U2758 (N_2758,N_2670,N_2636);
xnor U2759 (N_2759,N_2636,N_2682);
nand U2760 (N_2760,N_2627,N_2628);
nor U2761 (N_2761,N_2610,N_2607);
and U2762 (N_2762,N_2660,N_2645);
nand U2763 (N_2763,N_2684,N_2636);
nand U2764 (N_2764,N_2610,N_2655);
xnor U2765 (N_2765,N_2695,N_2604);
nor U2766 (N_2766,N_2659,N_2636);
xor U2767 (N_2767,N_2653,N_2692);
xnor U2768 (N_2768,N_2627,N_2694);
nor U2769 (N_2769,N_2609,N_2695);
or U2770 (N_2770,N_2677,N_2645);
xor U2771 (N_2771,N_2690,N_2697);
nand U2772 (N_2772,N_2666,N_2693);
nand U2773 (N_2773,N_2651,N_2653);
xor U2774 (N_2774,N_2632,N_2665);
and U2775 (N_2775,N_2625,N_2693);
or U2776 (N_2776,N_2616,N_2601);
or U2777 (N_2777,N_2656,N_2692);
and U2778 (N_2778,N_2696,N_2626);
or U2779 (N_2779,N_2620,N_2675);
or U2780 (N_2780,N_2671,N_2630);
xor U2781 (N_2781,N_2658,N_2631);
xnor U2782 (N_2782,N_2642,N_2652);
and U2783 (N_2783,N_2612,N_2651);
or U2784 (N_2784,N_2637,N_2630);
nand U2785 (N_2785,N_2618,N_2602);
and U2786 (N_2786,N_2680,N_2642);
nand U2787 (N_2787,N_2622,N_2657);
nand U2788 (N_2788,N_2644,N_2676);
nand U2789 (N_2789,N_2682,N_2627);
or U2790 (N_2790,N_2656,N_2642);
and U2791 (N_2791,N_2682,N_2613);
nand U2792 (N_2792,N_2686,N_2602);
xor U2793 (N_2793,N_2683,N_2670);
and U2794 (N_2794,N_2625,N_2678);
nor U2795 (N_2795,N_2607,N_2669);
nor U2796 (N_2796,N_2652,N_2694);
xnor U2797 (N_2797,N_2637,N_2664);
nor U2798 (N_2798,N_2674,N_2673);
and U2799 (N_2799,N_2652,N_2686);
and U2800 (N_2800,N_2780,N_2746);
xor U2801 (N_2801,N_2768,N_2748);
xnor U2802 (N_2802,N_2759,N_2792);
or U2803 (N_2803,N_2794,N_2715);
nand U2804 (N_2804,N_2770,N_2772);
and U2805 (N_2805,N_2717,N_2743);
nand U2806 (N_2806,N_2752,N_2790);
nor U2807 (N_2807,N_2731,N_2703);
and U2808 (N_2808,N_2791,N_2756);
xnor U2809 (N_2809,N_2749,N_2753);
or U2810 (N_2810,N_2718,N_2741);
nor U2811 (N_2811,N_2775,N_2757);
or U2812 (N_2812,N_2719,N_2742);
xnor U2813 (N_2813,N_2789,N_2706);
nor U2814 (N_2814,N_2773,N_2744);
nor U2815 (N_2815,N_2722,N_2798);
or U2816 (N_2816,N_2782,N_2734);
nand U2817 (N_2817,N_2755,N_2745);
and U2818 (N_2818,N_2716,N_2728);
xnor U2819 (N_2819,N_2760,N_2705);
or U2820 (N_2820,N_2785,N_2727);
and U2821 (N_2821,N_2712,N_2771);
nand U2822 (N_2822,N_2729,N_2737);
nor U2823 (N_2823,N_2767,N_2764);
or U2824 (N_2824,N_2709,N_2776);
nand U2825 (N_2825,N_2786,N_2788);
nor U2826 (N_2826,N_2799,N_2751);
nor U2827 (N_2827,N_2740,N_2702);
xnor U2828 (N_2828,N_2779,N_2713);
xor U2829 (N_2829,N_2750,N_2781);
xor U2830 (N_2830,N_2714,N_2730);
nand U2831 (N_2831,N_2784,N_2738);
or U2832 (N_2832,N_2778,N_2723);
and U2833 (N_2833,N_2747,N_2766);
nor U2834 (N_2834,N_2787,N_2701);
and U2835 (N_2835,N_2704,N_2707);
nand U2836 (N_2836,N_2769,N_2700);
nand U2837 (N_2837,N_2795,N_2720);
nand U2838 (N_2838,N_2758,N_2754);
or U2839 (N_2839,N_2777,N_2724);
nor U2840 (N_2840,N_2761,N_2774);
or U2841 (N_2841,N_2783,N_2726);
or U2842 (N_2842,N_2796,N_2735);
or U2843 (N_2843,N_2711,N_2763);
and U2844 (N_2844,N_2765,N_2721);
and U2845 (N_2845,N_2732,N_2797);
nand U2846 (N_2846,N_2736,N_2733);
and U2847 (N_2847,N_2793,N_2708);
xor U2848 (N_2848,N_2739,N_2710);
xor U2849 (N_2849,N_2725,N_2762);
or U2850 (N_2850,N_2778,N_2725);
and U2851 (N_2851,N_2708,N_2755);
nand U2852 (N_2852,N_2787,N_2798);
nor U2853 (N_2853,N_2755,N_2747);
nand U2854 (N_2854,N_2763,N_2770);
xor U2855 (N_2855,N_2770,N_2738);
and U2856 (N_2856,N_2739,N_2795);
xnor U2857 (N_2857,N_2746,N_2745);
nor U2858 (N_2858,N_2706,N_2741);
xnor U2859 (N_2859,N_2731,N_2798);
xnor U2860 (N_2860,N_2702,N_2797);
xor U2861 (N_2861,N_2744,N_2783);
and U2862 (N_2862,N_2709,N_2758);
xnor U2863 (N_2863,N_2729,N_2786);
xnor U2864 (N_2864,N_2787,N_2727);
and U2865 (N_2865,N_2725,N_2759);
xnor U2866 (N_2866,N_2732,N_2710);
nor U2867 (N_2867,N_2754,N_2750);
or U2868 (N_2868,N_2720,N_2776);
or U2869 (N_2869,N_2762,N_2774);
nor U2870 (N_2870,N_2798,N_2758);
and U2871 (N_2871,N_2719,N_2705);
and U2872 (N_2872,N_2706,N_2769);
nor U2873 (N_2873,N_2735,N_2758);
and U2874 (N_2874,N_2767,N_2760);
and U2875 (N_2875,N_2764,N_2752);
nor U2876 (N_2876,N_2742,N_2739);
nor U2877 (N_2877,N_2721,N_2764);
and U2878 (N_2878,N_2765,N_2743);
xor U2879 (N_2879,N_2778,N_2787);
nor U2880 (N_2880,N_2779,N_2705);
nand U2881 (N_2881,N_2728,N_2710);
and U2882 (N_2882,N_2716,N_2734);
nand U2883 (N_2883,N_2730,N_2725);
nor U2884 (N_2884,N_2756,N_2743);
or U2885 (N_2885,N_2756,N_2757);
nor U2886 (N_2886,N_2705,N_2724);
nand U2887 (N_2887,N_2708,N_2726);
and U2888 (N_2888,N_2768,N_2716);
nor U2889 (N_2889,N_2774,N_2760);
nand U2890 (N_2890,N_2783,N_2738);
nor U2891 (N_2891,N_2746,N_2717);
xor U2892 (N_2892,N_2747,N_2733);
nand U2893 (N_2893,N_2791,N_2718);
xor U2894 (N_2894,N_2724,N_2713);
or U2895 (N_2895,N_2713,N_2711);
and U2896 (N_2896,N_2703,N_2727);
nand U2897 (N_2897,N_2778,N_2724);
xnor U2898 (N_2898,N_2793,N_2763);
nand U2899 (N_2899,N_2736,N_2723);
xnor U2900 (N_2900,N_2858,N_2828);
and U2901 (N_2901,N_2817,N_2804);
nor U2902 (N_2902,N_2882,N_2899);
xnor U2903 (N_2903,N_2810,N_2811);
nand U2904 (N_2904,N_2879,N_2873);
nand U2905 (N_2905,N_2809,N_2830);
or U2906 (N_2906,N_2876,N_2853);
and U2907 (N_2907,N_2813,N_2863);
nand U2908 (N_2908,N_2869,N_2886);
and U2909 (N_2909,N_2815,N_2812);
or U2910 (N_2910,N_2861,N_2803);
xor U2911 (N_2911,N_2832,N_2884);
nand U2912 (N_2912,N_2857,N_2829);
and U2913 (N_2913,N_2872,N_2868);
xor U2914 (N_2914,N_2881,N_2859);
nand U2915 (N_2915,N_2888,N_2844);
and U2916 (N_2916,N_2845,N_2854);
xor U2917 (N_2917,N_2852,N_2898);
nor U2918 (N_2918,N_2864,N_2891);
or U2919 (N_2919,N_2826,N_2802);
or U2920 (N_2920,N_2820,N_2897);
xnor U2921 (N_2921,N_2831,N_2850);
nor U2922 (N_2922,N_2877,N_2893);
nand U2923 (N_2923,N_2800,N_2822);
or U2924 (N_2924,N_2819,N_2806);
nor U2925 (N_2925,N_2875,N_2894);
or U2926 (N_2926,N_2838,N_2827);
nand U2927 (N_2927,N_2878,N_2833);
or U2928 (N_2928,N_2895,N_2842);
nand U2929 (N_2929,N_2835,N_2890);
or U2930 (N_2930,N_2801,N_2846);
and U2931 (N_2931,N_2818,N_2865);
nor U2932 (N_2932,N_2885,N_2814);
nor U2933 (N_2933,N_2837,N_2834);
and U2934 (N_2934,N_2847,N_2862);
nor U2935 (N_2935,N_2892,N_2889);
or U2936 (N_2936,N_2807,N_2839);
or U2937 (N_2937,N_2887,N_2824);
or U2938 (N_2938,N_2866,N_2871);
nor U2939 (N_2939,N_2851,N_2823);
or U2940 (N_2940,N_2855,N_2836);
and U2941 (N_2941,N_2821,N_2870);
xnor U2942 (N_2942,N_2805,N_2860);
nand U2943 (N_2943,N_2896,N_2840);
nand U2944 (N_2944,N_2841,N_2848);
or U2945 (N_2945,N_2808,N_2883);
xnor U2946 (N_2946,N_2816,N_2867);
or U2947 (N_2947,N_2843,N_2856);
xnor U2948 (N_2948,N_2849,N_2880);
nor U2949 (N_2949,N_2874,N_2825);
nand U2950 (N_2950,N_2816,N_2801);
nand U2951 (N_2951,N_2806,N_2853);
and U2952 (N_2952,N_2885,N_2822);
or U2953 (N_2953,N_2868,N_2807);
nor U2954 (N_2954,N_2834,N_2821);
xor U2955 (N_2955,N_2822,N_2871);
and U2956 (N_2956,N_2824,N_2859);
and U2957 (N_2957,N_2894,N_2800);
and U2958 (N_2958,N_2829,N_2818);
nand U2959 (N_2959,N_2847,N_2813);
and U2960 (N_2960,N_2870,N_2819);
or U2961 (N_2961,N_2848,N_2861);
xor U2962 (N_2962,N_2839,N_2826);
nor U2963 (N_2963,N_2842,N_2835);
or U2964 (N_2964,N_2860,N_2870);
xnor U2965 (N_2965,N_2898,N_2809);
nor U2966 (N_2966,N_2831,N_2846);
nand U2967 (N_2967,N_2830,N_2886);
or U2968 (N_2968,N_2835,N_2868);
and U2969 (N_2969,N_2857,N_2850);
xor U2970 (N_2970,N_2833,N_2859);
and U2971 (N_2971,N_2859,N_2826);
nand U2972 (N_2972,N_2869,N_2885);
and U2973 (N_2973,N_2825,N_2885);
and U2974 (N_2974,N_2822,N_2880);
and U2975 (N_2975,N_2800,N_2805);
nand U2976 (N_2976,N_2801,N_2894);
nand U2977 (N_2977,N_2895,N_2835);
nor U2978 (N_2978,N_2831,N_2897);
or U2979 (N_2979,N_2811,N_2843);
nor U2980 (N_2980,N_2856,N_2837);
and U2981 (N_2981,N_2821,N_2847);
nand U2982 (N_2982,N_2811,N_2877);
nor U2983 (N_2983,N_2885,N_2856);
nor U2984 (N_2984,N_2805,N_2893);
or U2985 (N_2985,N_2827,N_2834);
or U2986 (N_2986,N_2869,N_2847);
and U2987 (N_2987,N_2803,N_2878);
and U2988 (N_2988,N_2815,N_2869);
or U2989 (N_2989,N_2820,N_2862);
xnor U2990 (N_2990,N_2890,N_2810);
xnor U2991 (N_2991,N_2842,N_2859);
nand U2992 (N_2992,N_2815,N_2838);
xnor U2993 (N_2993,N_2835,N_2833);
xor U2994 (N_2994,N_2838,N_2817);
and U2995 (N_2995,N_2884,N_2800);
nand U2996 (N_2996,N_2885,N_2886);
xnor U2997 (N_2997,N_2835,N_2859);
and U2998 (N_2998,N_2821,N_2874);
and U2999 (N_2999,N_2825,N_2848);
xor U3000 (N_3000,N_2911,N_2950);
or U3001 (N_3001,N_2971,N_2906);
and U3002 (N_3002,N_2914,N_2976);
xnor U3003 (N_3003,N_2931,N_2942);
or U3004 (N_3004,N_2980,N_2915);
xor U3005 (N_3005,N_2917,N_2945);
xor U3006 (N_3006,N_2969,N_2987);
nor U3007 (N_3007,N_2975,N_2966);
and U3008 (N_3008,N_2955,N_2959);
nand U3009 (N_3009,N_2968,N_2948);
nor U3010 (N_3010,N_2903,N_2933);
or U3011 (N_3011,N_2956,N_2900);
or U3012 (N_3012,N_2994,N_2918);
nor U3013 (N_3013,N_2916,N_2992);
nor U3014 (N_3014,N_2929,N_2977);
nor U3015 (N_3015,N_2961,N_2951);
nand U3016 (N_3016,N_2995,N_2937);
xor U3017 (N_3017,N_2946,N_2943);
or U3018 (N_3018,N_2963,N_2960);
nand U3019 (N_3019,N_2909,N_2949);
and U3020 (N_3020,N_2979,N_2940);
nor U3021 (N_3021,N_2954,N_2953);
and U3022 (N_3022,N_2985,N_2988);
or U3023 (N_3023,N_2962,N_2934);
or U3024 (N_3024,N_2908,N_2913);
and U3025 (N_3025,N_2907,N_2905);
nand U3026 (N_3026,N_2996,N_2998);
or U3027 (N_3027,N_2997,N_2935);
nand U3028 (N_3028,N_2967,N_2970);
nand U3029 (N_3029,N_2930,N_2964);
and U3030 (N_3030,N_2981,N_2904);
nand U3031 (N_3031,N_2919,N_2901);
nand U3032 (N_3032,N_2989,N_2982);
nand U3033 (N_3033,N_2983,N_2986);
xnor U3034 (N_3034,N_2938,N_2974);
or U3035 (N_3035,N_2921,N_2958);
nor U3036 (N_3036,N_2912,N_2952);
nor U3037 (N_3037,N_2925,N_2972);
nor U3038 (N_3038,N_2923,N_2941);
xnor U3039 (N_3039,N_2973,N_2932);
nand U3040 (N_3040,N_2990,N_2902);
xnor U3041 (N_3041,N_2920,N_2984);
xor U3042 (N_3042,N_2924,N_2926);
nand U3043 (N_3043,N_2910,N_2965);
and U3044 (N_3044,N_2999,N_2939);
and U3045 (N_3045,N_2928,N_2922);
or U3046 (N_3046,N_2978,N_2944);
or U3047 (N_3047,N_2957,N_2947);
nor U3048 (N_3048,N_2991,N_2993);
nand U3049 (N_3049,N_2936,N_2927);
nand U3050 (N_3050,N_2972,N_2977);
nand U3051 (N_3051,N_2911,N_2920);
and U3052 (N_3052,N_2979,N_2973);
nand U3053 (N_3053,N_2968,N_2935);
nor U3054 (N_3054,N_2916,N_2902);
nor U3055 (N_3055,N_2923,N_2956);
nor U3056 (N_3056,N_2915,N_2954);
nor U3057 (N_3057,N_2932,N_2960);
nand U3058 (N_3058,N_2915,N_2957);
nand U3059 (N_3059,N_2908,N_2946);
and U3060 (N_3060,N_2987,N_2952);
xor U3061 (N_3061,N_2924,N_2987);
and U3062 (N_3062,N_2909,N_2934);
nor U3063 (N_3063,N_2934,N_2956);
nor U3064 (N_3064,N_2940,N_2959);
and U3065 (N_3065,N_2987,N_2933);
nor U3066 (N_3066,N_2977,N_2962);
xor U3067 (N_3067,N_2962,N_2933);
xnor U3068 (N_3068,N_2902,N_2933);
and U3069 (N_3069,N_2925,N_2932);
and U3070 (N_3070,N_2933,N_2980);
nor U3071 (N_3071,N_2971,N_2933);
nor U3072 (N_3072,N_2978,N_2902);
nand U3073 (N_3073,N_2908,N_2999);
or U3074 (N_3074,N_2950,N_2945);
or U3075 (N_3075,N_2953,N_2946);
xor U3076 (N_3076,N_2908,N_2934);
nand U3077 (N_3077,N_2925,N_2917);
nor U3078 (N_3078,N_2927,N_2995);
and U3079 (N_3079,N_2952,N_2955);
or U3080 (N_3080,N_2930,N_2973);
and U3081 (N_3081,N_2906,N_2986);
nor U3082 (N_3082,N_2917,N_2918);
nor U3083 (N_3083,N_2907,N_2998);
nand U3084 (N_3084,N_2939,N_2913);
nor U3085 (N_3085,N_2956,N_2955);
nor U3086 (N_3086,N_2952,N_2905);
or U3087 (N_3087,N_2944,N_2986);
or U3088 (N_3088,N_2909,N_2937);
xnor U3089 (N_3089,N_2921,N_2915);
or U3090 (N_3090,N_2918,N_2929);
or U3091 (N_3091,N_2917,N_2904);
nand U3092 (N_3092,N_2950,N_2968);
and U3093 (N_3093,N_2954,N_2988);
nor U3094 (N_3094,N_2911,N_2931);
or U3095 (N_3095,N_2904,N_2978);
and U3096 (N_3096,N_2976,N_2919);
nor U3097 (N_3097,N_2934,N_2915);
and U3098 (N_3098,N_2949,N_2998);
or U3099 (N_3099,N_2902,N_2982);
xnor U3100 (N_3100,N_3085,N_3006);
xor U3101 (N_3101,N_3048,N_3038);
xor U3102 (N_3102,N_3062,N_3044);
and U3103 (N_3103,N_3002,N_3087);
nor U3104 (N_3104,N_3036,N_3058);
and U3105 (N_3105,N_3080,N_3015);
or U3106 (N_3106,N_3041,N_3081);
nor U3107 (N_3107,N_3095,N_3074);
nor U3108 (N_3108,N_3027,N_3089);
xnor U3109 (N_3109,N_3012,N_3020);
nor U3110 (N_3110,N_3028,N_3025);
and U3111 (N_3111,N_3014,N_3098);
or U3112 (N_3112,N_3059,N_3088);
xnor U3113 (N_3113,N_3021,N_3051);
xor U3114 (N_3114,N_3086,N_3071);
and U3115 (N_3115,N_3037,N_3091);
xnor U3116 (N_3116,N_3068,N_3061);
nand U3117 (N_3117,N_3073,N_3032);
and U3118 (N_3118,N_3056,N_3023);
xor U3119 (N_3119,N_3093,N_3026);
xor U3120 (N_3120,N_3016,N_3053);
xor U3121 (N_3121,N_3035,N_3039);
nand U3122 (N_3122,N_3001,N_3034);
nand U3123 (N_3123,N_3007,N_3043);
nand U3124 (N_3124,N_3049,N_3009);
xor U3125 (N_3125,N_3090,N_3013);
xor U3126 (N_3126,N_3094,N_3065);
and U3127 (N_3127,N_3045,N_3047);
nand U3128 (N_3128,N_3054,N_3077);
or U3129 (N_3129,N_3079,N_3030);
nand U3130 (N_3130,N_3092,N_3097);
and U3131 (N_3131,N_3033,N_3050);
or U3132 (N_3132,N_3042,N_3017);
xnor U3133 (N_3133,N_3010,N_3083);
xor U3134 (N_3134,N_3072,N_3067);
and U3135 (N_3135,N_3075,N_3022);
xor U3136 (N_3136,N_3076,N_3063);
and U3137 (N_3137,N_3040,N_3070);
xor U3138 (N_3138,N_3031,N_3099);
and U3139 (N_3139,N_3008,N_3069);
and U3140 (N_3140,N_3003,N_3078);
nor U3141 (N_3141,N_3024,N_3046);
or U3142 (N_3142,N_3055,N_3004);
nand U3143 (N_3143,N_3000,N_3018);
nand U3144 (N_3144,N_3060,N_3052);
and U3145 (N_3145,N_3084,N_3011);
and U3146 (N_3146,N_3082,N_3005);
nand U3147 (N_3147,N_3029,N_3096);
nand U3148 (N_3148,N_3064,N_3057);
nor U3149 (N_3149,N_3066,N_3019);
nand U3150 (N_3150,N_3081,N_3005);
nand U3151 (N_3151,N_3053,N_3086);
or U3152 (N_3152,N_3038,N_3074);
xnor U3153 (N_3153,N_3036,N_3056);
or U3154 (N_3154,N_3053,N_3064);
nand U3155 (N_3155,N_3010,N_3063);
xor U3156 (N_3156,N_3066,N_3018);
nand U3157 (N_3157,N_3091,N_3016);
xor U3158 (N_3158,N_3032,N_3055);
or U3159 (N_3159,N_3014,N_3086);
or U3160 (N_3160,N_3093,N_3034);
nand U3161 (N_3161,N_3033,N_3017);
and U3162 (N_3162,N_3059,N_3081);
or U3163 (N_3163,N_3057,N_3027);
xnor U3164 (N_3164,N_3094,N_3017);
nor U3165 (N_3165,N_3002,N_3023);
or U3166 (N_3166,N_3031,N_3092);
or U3167 (N_3167,N_3076,N_3014);
or U3168 (N_3168,N_3033,N_3066);
and U3169 (N_3169,N_3048,N_3060);
and U3170 (N_3170,N_3011,N_3030);
nand U3171 (N_3171,N_3013,N_3093);
nand U3172 (N_3172,N_3020,N_3053);
xor U3173 (N_3173,N_3093,N_3009);
nor U3174 (N_3174,N_3071,N_3088);
nor U3175 (N_3175,N_3027,N_3003);
xnor U3176 (N_3176,N_3039,N_3070);
and U3177 (N_3177,N_3083,N_3033);
or U3178 (N_3178,N_3096,N_3036);
or U3179 (N_3179,N_3035,N_3013);
or U3180 (N_3180,N_3086,N_3018);
and U3181 (N_3181,N_3023,N_3057);
xor U3182 (N_3182,N_3045,N_3087);
nor U3183 (N_3183,N_3004,N_3021);
xor U3184 (N_3184,N_3024,N_3050);
xor U3185 (N_3185,N_3046,N_3044);
and U3186 (N_3186,N_3090,N_3050);
nand U3187 (N_3187,N_3032,N_3018);
or U3188 (N_3188,N_3090,N_3033);
or U3189 (N_3189,N_3099,N_3053);
xnor U3190 (N_3190,N_3081,N_3033);
nand U3191 (N_3191,N_3045,N_3020);
or U3192 (N_3192,N_3003,N_3028);
xnor U3193 (N_3193,N_3051,N_3034);
nand U3194 (N_3194,N_3045,N_3070);
xor U3195 (N_3195,N_3062,N_3050);
nand U3196 (N_3196,N_3085,N_3000);
nor U3197 (N_3197,N_3025,N_3063);
and U3198 (N_3198,N_3035,N_3050);
nor U3199 (N_3199,N_3057,N_3032);
xor U3200 (N_3200,N_3192,N_3131);
or U3201 (N_3201,N_3154,N_3105);
and U3202 (N_3202,N_3178,N_3185);
and U3203 (N_3203,N_3125,N_3115);
and U3204 (N_3204,N_3111,N_3110);
nand U3205 (N_3205,N_3177,N_3103);
nor U3206 (N_3206,N_3187,N_3104);
and U3207 (N_3207,N_3174,N_3123);
xor U3208 (N_3208,N_3138,N_3194);
and U3209 (N_3209,N_3183,N_3188);
nor U3210 (N_3210,N_3151,N_3164);
and U3211 (N_3211,N_3150,N_3118);
xor U3212 (N_3212,N_3160,N_3112);
nand U3213 (N_3213,N_3173,N_3158);
or U3214 (N_3214,N_3133,N_3152);
and U3215 (N_3215,N_3153,N_3163);
or U3216 (N_3216,N_3147,N_3184);
and U3217 (N_3217,N_3132,N_3137);
and U3218 (N_3218,N_3175,N_3180);
nor U3219 (N_3219,N_3100,N_3195);
nand U3220 (N_3220,N_3146,N_3142);
or U3221 (N_3221,N_3108,N_3120);
nor U3222 (N_3222,N_3161,N_3168);
nor U3223 (N_3223,N_3196,N_3186);
nor U3224 (N_3224,N_3141,N_3181);
nand U3225 (N_3225,N_3106,N_3189);
xor U3226 (N_3226,N_3198,N_3128);
and U3227 (N_3227,N_3162,N_3170);
nor U3228 (N_3228,N_3172,N_3157);
nand U3229 (N_3229,N_3199,N_3193);
or U3230 (N_3230,N_3136,N_3109);
xnor U3231 (N_3231,N_3121,N_3159);
nand U3232 (N_3232,N_3130,N_3140);
xor U3233 (N_3233,N_3191,N_3139);
nor U3234 (N_3234,N_3190,N_3127);
nand U3235 (N_3235,N_3126,N_3129);
xor U3236 (N_3236,N_3165,N_3124);
and U3237 (N_3237,N_3135,N_3114);
nand U3238 (N_3238,N_3119,N_3143);
and U3239 (N_3239,N_3101,N_3117);
or U3240 (N_3240,N_3156,N_3113);
or U3241 (N_3241,N_3166,N_3144);
nor U3242 (N_3242,N_3197,N_3149);
xor U3243 (N_3243,N_3171,N_3167);
or U3244 (N_3244,N_3102,N_3107);
nor U3245 (N_3245,N_3148,N_3179);
or U3246 (N_3246,N_3182,N_3145);
nand U3247 (N_3247,N_3155,N_3134);
nand U3248 (N_3248,N_3116,N_3169);
nand U3249 (N_3249,N_3176,N_3122);
nand U3250 (N_3250,N_3127,N_3132);
xor U3251 (N_3251,N_3103,N_3104);
and U3252 (N_3252,N_3180,N_3135);
nor U3253 (N_3253,N_3158,N_3155);
and U3254 (N_3254,N_3158,N_3146);
nor U3255 (N_3255,N_3167,N_3122);
or U3256 (N_3256,N_3120,N_3190);
or U3257 (N_3257,N_3149,N_3151);
nor U3258 (N_3258,N_3176,N_3110);
and U3259 (N_3259,N_3142,N_3173);
and U3260 (N_3260,N_3102,N_3159);
or U3261 (N_3261,N_3100,N_3112);
nand U3262 (N_3262,N_3147,N_3109);
and U3263 (N_3263,N_3142,N_3144);
and U3264 (N_3264,N_3172,N_3155);
nand U3265 (N_3265,N_3148,N_3110);
xnor U3266 (N_3266,N_3103,N_3135);
nor U3267 (N_3267,N_3166,N_3106);
and U3268 (N_3268,N_3110,N_3122);
nand U3269 (N_3269,N_3130,N_3177);
xnor U3270 (N_3270,N_3152,N_3129);
nor U3271 (N_3271,N_3103,N_3140);
xnor U3272 (N_3272,N_3124,N_3129);
and U3273 (N_3273,N_3149,N_3193);
and U3274 (N_3274,N_3120,N_3151);
and U3275 (N_3275,N_3128,N_3145);
xor U3276 (N_3276,N_3106,N_3172);
nand U3277 (N_3277,N_3177,N_3105);
or U3278 (N_3278,N_3117,N_3135);
nor U3279 (N_3279,N_3110,N_3142);
or U3280 (N_3280,N_3100,N_3163);
xor U3281 (N_3281,N_3104,N_3195);
nor U3282 (N_3282,N_3113,N_3158);
nand U3283 (N_3283,N_3154,N_3130);
and U3284 (N_3284,N_3138,N_3139);
nor U3285 (N_3285,N_3105,N_3122);
and U3286 (N_3286,N_3166,N_3172);
and U3287 (N_3287,N_3176,N_3113);
xor U3288 (N_3288,N_3138,N_3148);
xnor U3289 (N_3289,N_3113,N_3167);
nor U3290 (N_3290,N_3132,N_3154);
and U3291 (N_3291,N_3111,N_3140);
and U3292 (N_3292,N_3153,N_3116);
nand U3293 (N_3293,N_3101,N_3164);
nor U3294 (N_3294,N_3157,N_3106);
nand U3295 (N_3295,N_3182,N_3115);
nand U3296 (N_3296,N_3138,N_3130);
and U3297 (N_3297,N_3100,N_3156);
or U3298 (N_3298,N_3163,N_3184);
nand U3299 (N_3299,N_3159,N_3128);
xnor U3300 (N_3300,N_3253,N_3245);
and U3301 (N_3301,N_3215,N_3238);
xnor U3302 (N_3302,N_3243,N_3225);
and U3303 (N_3303,N_3205,N_3230);
nand U3304 (N_3304,N_3224,N_3278);
xor U3305 (N_3305,N_3261,N_3202);
nand U3306 (N_3306,N_3209,N_3216);
nor U3307 (N_3307,N_3212,N_3268);
nand U3308 (N_3308,N_3242,N_3281);
nor U3309 (N_3309,N_3201,N_3291);
nor U3310 (N_3310,N_3249,N_3221);
and U3311 (N_3311,N_3297,N_3274);
nor U3312 (N_3312,N_3271,N_3246);
and U3313 (N_3313,N_3257,N_3284);
and U3314 (N_3314,N_3295,N_3267);
nand U3315 (N_3315,N_3208,N_3247);
nand U3316 (N_3316,N_3256,N_3254);
or U3317 (N_3317,N_3235,N_3207);
and U3318 (N_3318,N_3232,N_3236);
nor U3319 (N_3319,N_3227,N_3229);
nand U3320 (N_3320,N_3283,N_3270);
or U3321 (N_3321,N_3282,N_3237);
xor U3322 (N_3322,N_3258,N_3259);
nand U3323 (N_3323,N_3203,N_3260);
nand U3324 (N_3324,N_3285,N_3288);
or U3325 (N_3325,N_3277,N_3231);
nor U3326 (N_3326,N_3290,N_3248);
or U3327 (N_3327,N_3293,N_3223);
nor U3328 (N_3328,N_3286,N_3273);
nand U3329 (N_3329,N_3250,N_3269);
nand U3330 (N_3330,N_3265,N_3228);
nor U3331 (N_3331,N_3206,N_3280);
nor U3332 (N_3332,N_3294,N_3255);
or U3333 (N_3333,N_3275,N_3211);
xnor U3334 (N_3334,N_3276,N_3226);
or U3335 (N_3335,N_3262,N_3204);
or U3336 (N_3336,N_3210,N_3214);
xnor U3337 (N_3337,N_3289,N_3200);
nor U3338 (N_3338,N_3252,N_3264);
and U3339 (N_3339,N_3240,N_3222);
xnor U3340 (N_3340,N_3244,N_3217);
nor U3341 (N_3341,N_3233,N_3251);
or U3342 (N_3342,N_3220,N_3241);
or U3343 (N_3343,N_3292,N_3213);
xnor U3344 (N_3344,N_3279,N_3234);
nand U3345 (N_3345,N_3272,N_3298);
nor U3346 (N_3346,N_3263,N_3218);
nand U3347 (N_3347,N_3219,N_3239);
nand U3348 (N_3348,N_3299,N_3287);
xnor U3349 (N_3349,N_3296,N_3266);
xor U3350 (N_3350,N_3225,N_3230);
and U3351 (N_3351,N_3259,N_3275);
xor U3352 (N_3352,N_3261,N_3230);
nand U3353 (N_3353,N_3207,N_3277);
xor U3354 (N_3354,N_3273,N_3223);
nand U3355 (N_3355,N_3269,N_3227);
and U3356 (N_3356,N_3224,N_3257);
nor U3357 (N_3357,N_3261,N_3242);
and U3358 (N_3358,N_3247,N_3241);
xor U3359 (N_3359,N_3213,N_3254);
xor U3360 (N_3360,N_3229,N_3266);
nand U3361 (N_3361,N_3287,N_3258);
nor U3362 (N_3362,N_3274,N_3241);
and U3363 (N_3363,N_3287,N_3214);
nor U3364 (N_3364,N_3225,N_3283);
xor U3365 (N_3365,N_3267,N_3255);
or U3366 (N_3366,N_3236,N_3226);
nor U3367 (N_3367,N_3234,N_3252);
xor U3368 (N_3368,N_3243,N_3222);
or U3369 (N_3369,N_3255,N_3242);
nor U3370 (N_3370,N_3238,N_3204);
and U3371 (N_3371,N_3255,N_3264);
xor U3372 (N_3372,N_3230,N_3258);
and U3373 (N_3373,N_3269,N_3298);
or U3374 (N_3374,N_3209,N_3258);
nor U3375 (N_3375,N_3263,N_3228);
nand U3376 (N_3376,N_3220,N_3249);
or U3377 (N_3377,N_3269,N_3208);
and U3378 (N_3378,N_3248,N_3247);
xnor U3379 (N_3379,N_3220,N_3224);
nand U3380 (N_3380,N_3284,N_3269);
and U3381 (N_3381,N_3252,N_3296);
and U3382 (N_3382,N_3234,N_3206);
or U3383 (N_3383,N_3212,N_3295);
and U3384 (N_3384,N_3294,N_3276);
nor U3385 (N_3385,N_3275,N_3221);
nand U3386 (N_3386,N_3221,N_3293);
or U3387 (N_3387,N_3299,N_3258);
and U3388 (N_3388,N_3229,N_3282);
and U3389 (N_3389,N_3273,N_3207);
or U3390 (N_3390,N_3248,N_3259);
nand U3391 (N_3391,N_3267,N_3247);
nand U3392 (N_3392,N_3267,N_3260);
or U3393 (N_3393,N_3297,N_3206);
nor U3394 (N_3394,N_3214,N_3288);
nand U3395 (N_3395,N_3204,N_3276);
nand U3396 (N_3396,N_3277,N_3206);
xnor U3397 (N_3397,N_3234,N_3220);
xnor U3398 (N_3398,N_3269,N_3205);
or U3399 (N_3399,N_3281,N_3210);
or U3400 (N_3400,N_3340,N_3360);
nand U3401 (N_3401,N_3312,N_3338);
nand U3402 (N_3402,N_3379,N_3365);
nor U3403 (N_3403,N_3374,N_3352);
and U3404 (N_3404,N_3333,N_3362);
nand U3405 (N_3405,N_3334,N_3372);
and U3406 (N_3406,N_3316,N_3383);
or U3407 (N_3407,N_3310,N_3339);
nand U3408 (N_3408,N_3341,N_3397);
nand U3409 (N_3409,N_3353,N_3395);
nand U3410 (N_3410,N_3344,N_3371);
nor U3411 (N_3411,N_3399,N_3394);
nor U3412 (N_3412,N_3331,N_3375);
xnor U3413 (N_3413,N_3386,N_3382);
or U3414 (N_3414,N_3350,N_3357);
or U3415 (N_3415,N_3358,N_3311);
and U3416 (N_3416,N_3346,N_3359);
xor U3417 (N_3417,N_3324,N_3369);
xnor U3418 (N_3418,N_3345,N_3396);
nand U3419 (N_3419,N_3349,N_3364);
xnor U3420 (N_3420,N_3335,N_3351);
and U3421 (N_3421,N_3332,N_3309);
nor U3422 (N_3422,N_3322,N_3388);
xnor U3423 (N_3423,N_3308,N_3329);
or U3424 (N_3424,N_3323,N_3366);
or U3425 (N_3425,N_3342,N_3327);
nand U3426 (N_3426,N_3302,N_3398);
and U3427 (N_3427,N_3385,N_3361);
xor U3428 (N_3428,N_3393,N_3336);
and U3429 (N_3429,N_3389,N_3320);
xnor U3430 (N_3430,N_3300,N_3392);
and U3431 (N_3431,N_3367,N_3315);
and U3432 (N_3432,N_3378,N_3380);
nor U3433 (N_3433,N_3368,N_3347);
nand U3434 (N_3434,N_3370,N_3355);
nor U3435 (N_3435,N_3391,N_3314);
or U3436 (N_3436,N_3301,N_3307);
xnor U3437 (N_3437,N_3373,N_3337);
xnor U3438 (N_3438,N_3363,N_3330);
nand U3439 (N_3439,N_3313,N_3356);
and U3440 (N_3440,N_3328,N_3303);
xor U3441 (N_3441,N_3376,N_3390);
xor U3442 (N_3442,N_3306,N_3377);
nand U3443 (N_3443,N_3325,N_3305);
or U3444 (N_3444,N_3321,N_3381);
and U3445 (N_3445,N_3343,N_3348);
and U3446 (N_3446,N_3387,N_3317);
nor U3447 (N_3447,N_3384,N_3319);
nor U3448 (N_3448,N_3354,N_3318);
nor U3449 (N_3449,N_3304,N_3326);
nand U3450 (N_3450,N_3319,N_3302);
nor U3451 (N_3451,N_3324,N_3315);
nor U3452 (N_3452,N_3363,N_3328);
and U3453 (N_3453,N_3356,N_3365);
or U3454 (N_3454,N_3310,N_3324);
and U3455 (N_3455,N_3300,N_3351);
and U3456 (N_3456,N_3339,N_3321);
nand U3457 (N_3457,N_3337,N_3388);
and U3458 (N_3458,N_3321,N_3379);
and U3459 (N_3459,N_3364,N_3376);
nor U3460 (N_3460,N_3342,N_3375);
or U3461 (N_3461,N_3380,N_3306);
and U3462 (N_3462,N_3392,N_3343);
nor U3463 (N_3463,N_3326,N_3392);
nand U3464 (N_3464,N_3387,N_3305);
and U3465 (N_3465,N_3381,N_3309);
and U3466 (N_3466,N_3309,N_3340);
xnor U3467 (N_3467,N_3372,N_3313);
nor U3468 (N_3468,N_3346,N_3380);
and U3469 (N_3469,N_3357,N_3342);
or U3470 (N_3470,N_3384,N_3336);
and U3471 (N_3471,N_3329,N_3370);
nor U3472 (N_3472,N_3303,N_3381);
xor U3473 (N_3473,N_3347,N_3342);
nor U3474 (N_3474,N_3319,N_3355);
or U3475 (N_3475,N_3369,N_3377);
and U3476 (N_3476,N_3364,N_3318);
or U3477 (N_3477,N_3357,N_3338);
nor U3478 (N_3478,N_3375,N_3350);
or U3479 (N_3479,N_3323,N_3331);
or U3480 (N_3480,N_3392,N_3314);
and U3481 (N_3481,N_3306,N_3333);
or U3482 (N_3482,N_3392,N_3336);
nand U3483 (N_3483,N_3308,N_3376);
and U3484 (N_3484,N_3351,N_3394);
or U3485 (N_3485,N_3327,N_3348);
or U3486 (N_3486,N_3376,N_3341);
or U3487 (N_3487,N_3368,N_3361);
nor U3488 (N_3488,N_3375,N_3328);
nand U3489 (N_3489,N_3364,N_3353);
and U3490 (N_3490,N_3364,N_3350);
xnor U3491 (N_3491,N_3385,N_3331);
xor U3492 (N_3492,N_3328,N_3321);
nor U3493 (N_3493,N_3311,N_3325);
xor U3494 (N_3494,N_3391,N_3319);
nor U3495 (N_3495,N_3330,N_3332);
xnor U3496 (N_3496,N_3358,N_3321);
and U3497 (N_3497,N_3302,N_3358);
nand U3498 (N_3498,N_3356,N_3388);
xnor U3499 (N_3499,N_3357,N_3309);
nor U3500 (N_3500,N_3471,N_3478);
and U3501 (N_3501,N_3442,N_3408);
xor U3502 (N_3502,N_3410,N_3402);
nand U3503 (N_3503,N_3400,N_3464);
and U3504 (N_3504,N_3436,N_3462);
nand U3505 (N_3505,N_3456,N_3492);
nor U3506 (N_3506,N_3495,N_3484);
nor U3507 (N_3507,N_3485,N_3433);
nand U3508 (N_3508,N_3474,N_3458);
and U3509 (N_3509,N_3438,N_3445);
xnor U3510 (N_3510,N_3424,N_3435);
and U3511 (N_3511,N_3472,N_3488);
nor U3512 (N_3512,N_3443,N_3430);
nand U3513 (N_3513,N_3461,N_3457);
xnor U3514 (N_3514,N_3429,N_3440);
or U3515 (N_3515,N_3480,N_3441);
and U3516 (N_3516,N_3418,N_3446);
nand U3517 (N_3517,N_3467,N_3466);
nor U3518 (N_3518,N_3494,N_3487);
or U3519 (N_3519,N_3482,N_3475);
nand U3520 (N_3520,N_3401,N_3451);
or U3521 (N_3521,N_3431,N_3499);
nand U3522 (N_3522,N_3416,N_3444);
nand U3523 (N_3523,N_3496,N_3497);
nor U3524 (N_3524,N_3407,N_3498);
nand U3525 (N_3525,N_3450,N_3449);
or U3526 (N_3526,N_3465,N_3422);
and U3527 (N_3527,N_3426,N_3493);
nor U3528 (N_3528,N_3406,N_3491);
xnor U3529 (N_3529,N_3414,N_3486);
nand U3530 (N_3530,N_3481,N_3409);
or U3531 (N_3531,N_3477,N_3448);
and U3532 (N_3532,N_3427,N_3454);
nand U3533 (N_3533,N_3420,N_3455);
nor U3534 (N_3534,N_3453,N_3476);
and U3535 (N_3535,N_3421,N_3404);
xor U3536 (N_3536,N_3437,N_3468);
or U3537 (N_3537,N_3425,N_3469);
nand U3538 (N_3538,N_3403,N_3473);
nand U3539 (N_3539,N_3479,N_3460);
nor U3540 (N_3540,N_3452,N_3447);
or U3541 (N_3541,N_3490,N_3423);
nor U3542 (N_3542,N_3417,N_3483);
or U3543 (N_3543,N_3405,N_3434);
nand U3544 (N_3544,N_3470,N_3411);
xor U3545 (N_3545,N_3439,N_3415);
and U3546 (N_3546,N_3428,N_3432);
nor U3547 (N_3547,N_3459,N_3463);
nor U3548 (N_3548,N_3413,N_3412);
nand U3549 (N_3549,N_3419,N_3489);
xnor U3550 (N_3550,N_3429,N_3486);
or U3551 (N_3551,N_3422,N_3400);
xnor U3552 (N_3552,N_3474,N_3468);
xnor U3553 (N_3553,N_3403,N_3439);
xor U3554 (N_3554,N_3419,N_3461);
or U3555 (N_3555,N_3486,N_3436);
and U3556 (N_3556,N_3407,N_3431);
and U3557 (N_3557,N_3477,N_3466);
xor U3558 (N_3558,N_3480,N_3460);
nand U3559 (N_3559,N_3411,N_3472);
xor U3560 (N_3560,N_3474,N_3489);
nand U3561 (N_3561,N_3430,N_3405);
and U3562 (N_3562,N_3428,N_3429);
xor U3563 (N_3563,N_3490,N_3404);
xnor U3564 (N_3564,N_3432,N_3421);
xnor U3565 (N_3565,N_3456,N_3444);
and U3566 (N_3566,N_3448,N_3443);
or U3567 (N_3567,N_3421,N_3442);
or U3568 (N_3568,N_3437,N_3462);
xnor U3569 (N_3569,N_3423,N_3426);
xnor U3570 (N_3570,N_3467,N_3410);
or U3571 (N_3571,N_3467,N_3465);
nor U3572 (N_3572,N_3425,N_3437);
and U3573 (N_3573,N_3449,N_3485);
nand U3574 (N_3574,N_3413,N_3499);
and U3575 (N_3575,N_3449,N_3461);
nand U3576 (N_3576,N_3442,N_3440);
and U3577 (N_3577,N_3473,N_3416);
nand U3578 (N_3578,N_3449,N_3454);
xnor U3579 (N_3579,N_3401,N_3468);
and U3580 (N_3580,N_3451,N_3434);
nor U3581 (N_3581,N_3465,N_3468);
or U3582 (N_3582,N_3480,N_3479);
and U3583 (N_3583,N_3486,N_3476);
and U3584 (N_3584,N_3426,N_3481);
nor U3585 (N_3585,N_3438,N_3456);
or U3586 (N_3586,N_3489,N_3442);
and U3587 (N_3587,N_3498,N_3493);
xnor U3588 (N_3588,N_3498,N_3460);
or U3589 (N_3589,N_3428,N_3437);
xor U3590 (N_3590,N_3471,N_3434);
nor U3591 (N_3591,N_3493,N_3419);
xnor U3592 (N_3592,N_3428,N_3445);
or U3593 (N_3593,N_3404,N_3488);
nor U3594 (N_3594,N_3459,N_3471);
and U3595 (N_3595,N_3432,N_3420);
and U3596 (N_3596,N_3434,N_3403);
xnor U3597 (N_3597,N_3462,N_3482);
or U3598 (N_3598,N_3438,N_3479);
nor U3599 (N_3599,N_3404,N_3482);
nand U3600 (N_3600,N_3583,N_3515);
nor U3601 (N_3601,N_3523,N_3526);
nor U3602 (N_3602,N_3538,N_3550);
nand U3603 (N_3603,N_3534,N_3537);
or U3604 (N_3604,N_3572,N_3511);
nor U3605 (N_3605,N_3553,N_3564);
and U3606 (N_3606,N_3546,N_3578);
xnor U3607 (N_3607,N_3576,N_3591);
xor U3608 (N_3608,N_3547,N_3584);
or U3609 (N_3609,N_3504,N_3574);
nor U3610 (N_3610,N_3517,N_3575);
nand U3611 (N_3611,N_3516,N_3530);
or U3612 (N_3612,N_3585,N_3542);
xnor U3613 (N_3613,N_3503,N_3598);
or U3614 (N_3614,N_3580,N_3502);
and U3615 (N_3615,N_3589,N_3563);
nor U3616 (N_3616,N_3567,N_3577);
nand U3617 (N_3617,N_3558,N_3548);
nor U3618 (N_3618,N_3596,N_3554);
or U3619 (N_3619,N_3532,N_3560);
or U3620 (N_3620,N_3568,N_3509);
nand U3621 (N_3621,N_3529,N_3559);
xnor U3622 (N_3622,N_3527,N_3522);
or U3623 (N_3623,N_3571,N_3587);
and U3624 (N_3624,N_3549,N_3531);
and U3625 (N_3625,N_3544,N_3590);
or U3626 (N_3626,N_3566,N_3552);
and U3627 (N_3627,N_3524,N_3599);
xor U3628 (N_3628,N_3555,N_3581);
nand U3629 (N_3629,N_3521,N_3597);
xnor U3630 (N_3630,N_3582,N_3557);
and U3631 (N_3631,N_3540,N_3592);
and U3632 (N_3632,N_3506,N_3565);
nand U3633 (N_3633,N_3586,N_3543);
xor U3634 (N_3634,N_3519,N_3501);
and U3635 (N_3635,N_3541,N_3545);
nand U3636 (N_3636,N_3595,N_3508);
nor U3637 (N_3637,N_3507,N_3533);
nor U3638 (N_3638,N_3536,N_3520);
or U3639 (N_3639,N_3562,N_3539);
nand U3640 (N_3640,N_3561,N_3535);
xnor U3641 (N_3641,N_3588,N_3513);
xnor U3642 (N_3642,N_3593,N_3570);
nor U3643 (N_3643,N_3500,N_3556);
or U3644 (N_3644,N_3594,N_3579);
nor U3645 (N_3645,N_3528,N_3505);
or U3646 (N_3646,N_3551,N_3514);
or U3647 (N_3647,N_3569,N_3525);
nand U3648 (N_3648,N_3518,N_3573);
nand U3649 (N_3649,N_3512,N_3510);
or U3650 (N_3650,N_3544,N_3531);
nand U3651 (N_3651,N_3516,N_3513);
or U3652 (N_3652,N_3550,N_3586);
nand U3653 (N_3653,N_3592,N_3508);
nor U3654 (N_3654,N_3583,N_3597);
and U3655 (N_3655,N_3574,N_3592);
and U3656 (N_3656,N_3574,N_3581);
and U3657 (N_3657,N_3554,N_3565);
xor U3658 (N_3658,N_3579,N_3572);
nor U3659 (N_3659,N_3562,N_3559);
nand U3660 (N_3660,N_3563,N_3534);
nor U3661 (N_3661,N_3584,N_3537);
and U3662 (N_3662,N_3576,N_3558);
or U3663 (N_3663,N_3505,N_3593);
xnor U3664 (N_3664,N_3502,N_3550);
nor U3665 (N_3665,N_3506,N_3545);
nand U3666 (N_3666,N_3575,N_3539);
or U3667 (N_3667,N_3562,N_3528);
and U3668 (N_3668,N_3566,N_3567);
nor U3669 (N_3669,N_3577,N_3557);
or U3670 (N_3670,N_3509,N_3563);
xor U3671 (N_3671,N_3576,N_3518);
nand U3672 (N_3672,N_3504,N_3593);
xnor U3673 (N_3673,N_3576,N_3594);
nor U3674 (N_3674,N_3557,N_3524);
and U3675 (N_3675,N_3514,N_3576);
and U3676 (N_3676,N_3543,N_3530);
nor U3677 (N_3677,N_3557,N_3586);
nor U3678 (N_3678,N_3528,N_3523);
and U3679 (N_3679,N_3504,N_3577);
xnor U3680 (N_3680,N_3541,N_3536);
nor U3681 (N_3681,N_3562,N_3556);
or U3682 (N_3682,N_3513,N_3573);
or U3683 (N_3683,N_3544,N_3512);
nor U3684 (N_3684,N_3506,N_3533);
nor U3685 (N_3685,N_3505,N_3571);
nor U3686 (N_3686,N_3535,N_3562);
or U3687 (N_3687,N_3505,N_3501);
nor U3688 (N_3688,N_3510,N_3592);
xnor U3689 (N_3689,N_3552,N_3506);
nand U3690 (N_3690,N_3529,N_3511);
xor U3691 (N_3691,N_3533,N_3544);
or U3692 (N_3692,N_3596,N_3593);
and U3693 (N_3693,N_3580,N_3528);
or U3694 (N_3694,N_3574,N_3540);
xnor U3695 (N_3695,N_3538,N_3517);
xor U3696 (N_3696,N_3541,N_3568);
or U3697 (N_3697,N_3586,N_3598);
xnor U3698 (N_3698,N_3587,N_3540);
nor U3699 (N_3699,N_3559,N_3545);
nor U3700 (N_3700,N_3626,N_3681);
or U3701 (N_3701,N_3669,N_3678);
nor U3702 (N_3702,N_3676,N_3611);
and U3703 (N_3703,N_3692,N_3685);
nor U3704 (N_3704,N_3697,N_3684);
nor U3705 (N_3705,N_3629,N_3666);
and U3706 (N_3706,N_3677,N_3696);
or U3707 (N_3707,N_3699,N_3693);
nand U3708 (N_3708,N_3672,N_3671);
nor U3709 (N_3709,N_3660,N_3646);
nand U3710 (N_3710,N_3689,N_3682);
nor U3711 (N_3711,N_3627,N_3680);
xnor U3712 (N_3712,N_3606,N_3670);
and U3713 (N_3713,N_3619,N_3600);
or U3714 (N_3714,N_3601,N_3673);
and U3715 (N_3715,N_3620,N_3634);
or U3716 (N_3716,N_3690,N_3665);
xnor U3717 (N_3717,N_3625,N_3624);
nand U3718 (N_3718,N_3605,N_3657);
or U3719 (N_3719,N_3663,N_3694);
nor U3720 (N_3720,N_3635,N_3630);
and U3721 (N_3721,N_3641,N_3609);
and U3722 (N_3722,N_3652,N_3686);
xnor U3723 (N_3723,N_3623,N_3645);
nand U3724 (N_3724,N_3698,N_3612);
or U3725 (N_3725,N_3644,N_3662);
xnor U3726 (N_3726,N_3658,N_3667);
nand U3727 (N_3727,N_3616,N_3618);
nor U3728 (N_3728,N_3633,N_3631);
or U3729 (N_3729,N_3642,N_3691);
and U3730 (N_3730,N_3607,N_3659);
or U3731 (N_3731,N_3639,N_3650);
or U3732 (N_3732,N_3622,N_3608);
or U3733 (N_3733,N_3674,N_3655);
xor U3734 (N_3734,N_3661,N_3604);
nand U3735 (N_3735,N_3648,N_3664);
nor U3736 (N_3736,N_3688,N_3603);
and U3737 (N_3737,N_3628,N_3617);
or U3738 (N_3738,N_3654,N_3679);
or U3739 (N_3739,N_3695,N_3614);
xnor U3740 (N_3740,N_3653,N_3637);
nor U3741 (N_3741,N_3675,N_3621);
nand U3742 (N_3742,N_3683,N_3643);
or U3743 (N_3743,N_3647,N_3602);
or U3744 (N_3744,N_3610,N_3687);
nor U3745 (N_3745,N_3613,N_3651);
nor U3746 (N_3746,N_3640,N_3656);
xnor U3747 (N_3747,N_3636,N_3668);
or U3748 (N_3748,N_3649,N_3638);
nand U3749 (N_3749,N_3615,N_3632);
or U3750 (N_3750,N_3644,N_3699);
or U3751 (N_3751,N_3670,N_3643);
and U3752 (N_3752,N_3692,N_3622);
and U3753 (N_3753,N_3632,N_3654);
nand U3754 (N_3754,N_3610,N_3601);
and U3755 (N_3755,N_3655,N_3697);
or U3756 (N_3756,N_3617,N_3613);
or U3757 (N_3757,N_3676,N_3660);
xor U3758 (N_3758,N_3646,N_3620);
xnor U3759 (N_3759,N_3612,N_3673);
and U3760 (N_3760,N_3639,N_3672);
and U3761 (N_3761,N_3662,N_3657);
nand U3762 (N_3762,N_3613,N_3600);
nor U3763 (N_3763,N_3641,N_3676);
nor U3764 (N_3764,N_3600,N_3699);
and U3765 (N_3765,N_3642,N_3612);
xnor U3766 (N_3766,N_3612,N_3611);
nand U3767 (N_3767,N_3646,N_3681);
and U3768 (N_3768,N_3656,N_3692);
xor U3769 (N_3769,N_3644,N_3668);
or U3770 (N_3770,N_3698,N_3669);
or U3771 (N_3771,N_3662,N_3618);
or U3772 (N_3772,N_3683,N_3657);
xor U3773 (N_3773,N_3616,N_3653);
or U3774 (N_3774,N_3689,N_3695);
xnor U3775 (N_3775,N_3644,N_3663);
xnor U3776 (N_3776,N_3695,N_3694);
nand U3777 (N_3777,N_3691,N_3648);
nor U3778 (N_3778,N_3635,N_3698);
nor U3779 (N_3779,N_3633,N_3668);
xor U3780 (N_3780,N_3606,N_3650);
nand U3781 (N_3781,N_3656,N_3665);
or U3782 (N_3782,N_3619,N_3601);
nand U3783 (N_3783,N_3661,N_3659);
nor U3784 (N_3784,N_3694,N_3628);
nand U3785 (N_3785,N_3658,N_3601);
xor U3786 (N_3786,N_3685,N_3668);
nand U3787 (N_3787,N_3627,N_3622);
and U3788 (N_3788,N_3623,N_3676);
nor U3789 (N_3789,N_3601,N_3607);
or U3790 (N_3790,N_3626,N_3678);
nand U3791 (N_3791,N_3616,N_3692);
nand U3792 (N_3792,N_3639,N_3633);
and U3793 (N_3793,N_3682,N_3638);
xnor U3794 (N_3794,N_3637,N_3649);
and U3795 (N_3795,N_3639,N_3651);
nand U3796 (N_3796,N_3675,N_3651);
or U3797 (N_3797,N_3618,N_3619);
xor U3798 (N_3798,N_3604,N_3636);
nor U3799 (N_3799,N_3639,N_3616);
nand U3800 (N_3800,N_3792,N_3722);
nor U3801 (N_3801,N_3707,N_3791);
xnor U3802 (N_3802,N_3750,N_3795);
and U3803 (N_3803,N_3769,N_3766);
nand U3804 (N_3804,N_3744,N_3763);
nand U3805 (N_3805,N_3786,N_3742);
and U3806 (N_3806,N_3737,N_3727);
and U3807 (N_3807,N_3701,N_3772);
nor U3808 (N_3808,N_3709,N_3756);
and U3809 (N_3809,N_3732,N_3782);
and U3810 (N_3810,N_3771,N_3787);
and U3811 (N_3811,N_3710,N_3778);
nor U3812 (N_3812,N_3779,N_3748);
nor U3813 (N_3813,N_3754,N_3726);
and U3814 (N_3814,N_3774,N_3735);
xor U3815 (N_3815,N_3780,N_3704);
nand U3816 (N_3816,N_3755,N_3764);
nand U3817 (N_3817,N_3738,N_3720);
or U3818 (N_3818,N_3719,N_3775);
and U3819 (N_3819,N_3739,N_3776);
nand U3820 (N_3820,N_3729,N_3794);
or U3821 (N_3821,N_3751,N_3700);
nor U3822 (N_3822,N_3702,N_3741);
xnor U3823 (N_3823,N_3784,N_3789);
nand U3824 (N_3824,N_3743,N_3797);
and U3825 (N_3825,N_3762,N_3734);
or U3826 (N_3826,N_3768,N_3712);
nand U3827 (N_3827,N_3714,N_3749);
or U3828 (N_3828,N_3798,N_3716);
nor U3829 (N_3829,N_3736,N_3746);
nand U3830 (N_3830,N_3713,N_3731);
nand U3831 (N_3831,N_3783,N_3745);
and U3832 (N_3832,N_3703,N_3781);
or U3833 (N_3833,N_3705,N_3721);
nor U3834 (N_3834,N_3770,N_3752);
nor U3835 (N_3835,N_3796,N_3747);
xnor U3836 (N_3836,N_3767,N_3759);
and U3837 (N_3837,N_3730,N_3717);
nor U3838 (N_3838,N_3788,N_3785);
and U3839 (N_3839,N_3740,N_3708);
nand U3840 (N_3840,N_3799,N_3777);
or U3841 (N_3841,N_3733,N_3724);
or U3842 (N_3842,N_3773,N_3718);
and U3843 (N_3843,N_3715,N_3790);
and U3844 (N_3844,N_3711,N_3760);
and U3845 (N_3845,N_3758,N_3793);
xnor U3846 (N_3846,N_3725,N_3753);
nor U3847 (N_3847,N_3761,N_3765);
and U3848 (N_3848,N_3706,N_3757);
and U3849 (N_3849,N_3728,N_3723);
and U3850 (N_3850,N_3724,N_3744);
nor U3851 (N_3851,N_3708,N_3792);
nand U3852 (N_3852,N_3719,N_3704);
or U3853 (N_3853,N_3759,N_3793);
nor U3854 (N_3854,N_3731,N_3759);
xnor U3855 (N_3855,N_3752,N_3722);
xnor U3856 (N_3856,N_3780,N_3725);
nor U3857 (N_3857,N_3700,N_3763);
nor U3858 (N_3858,N_3739,N_3762);
and U3859 (N_3859,N_3774,N_3707);
nor U3860 (N_3860,N_3786,N_3727);
or U3861 (N_3861,N_3736,N_3790);
or U3862 (N_3862,N_3795,N_3758);
xor U3863 (N_3863,N_3724,N_3759);
or U3864 (N_3864,N_3780,N_3709);
xor U3865 (N_3865,N_3783,N_3715);
and U3866 (N_3866,N_3798,N_3735);
nor U3867 (N_3867,N_3733,N_3715);
xnor U3868 (N_3868,N_3798,N_3763);
nor U3869 (N_3869,N_3775,N_3730);
or U3870 (N_3870,N_3722,N_3708);
and U3871 (N_3871,N_3731,N_3732);
or U3872 (N_3872,N_3764,N_3714);
xnor U3873 (N_3873,N_3772,N_3707);
nand U3874 (N_3874,N_3715,N_3754);
and U3875 (N_3875,N_3743,N_3744);
xnor U3876 (N_3876,N_3793,N_3752);
nand U3877 (N_3877,N_3790,N_3737);
nand U3878 (N_3878,N_3786,N_3710);
nand U3879 (N_3879,N_3713,N_3771);
and U3880 (N_3880,N_3731,N_3799);
or U3881 (N_3881,N_3731,N_3778);
and U3882 (N_3882,N_3717,N_3710);
nand U3883 (N_3883,N_3740,N_3753);
nand U3884 (N_3884,N_3773,N_3702);
and U3885 (N_3885,N_3722,N_3774);
and U3886 (N_3886,N_3792,N_3783);
nor U3887 (N_3887,N_3790,N_3781);
nand U3888 (N_3888,N_3719,N_3776);
xor U3889 (N_3889,N_3738,N_3764);
or U3890 (N_3890,N_3787,N_3741);
nand U3891 (N_3891,N_3738,N_3778);
xor U3892 (N_3892,N_3712,N_3779);
xor U3893 (N_3893,N_3711,N_3745);
and U3894 (N_3894,N_3718,N_3792);
or U3895 (N_3895,N_3725,N_3737);
nand U3896 (N_3896,N_3771,N_3795);
xor U3897 (N_3897,N_3778,N_3746);
and U3898 (N_3898,N_3794,N_3720);
xor U3899 (N_3899,N_3780,N_3754);
or U3900 (N_3900,N_3868,N_3890);
nand U3901 (N_3901,N_3881,N_3845);
nor U3902 (N_3902,N_3863,N_3824);
and U3903 (N_3903,N_3838,N_3805);
nand U3904 (N_3904,N_3807,N_3814);
or U3905 (N_3905,N_3813,N_3857);
nand U3906 (N_3906,N_3836,N_3806);
xor U3907 (N_3907,N_3865,N_3802);
or U3908 (N_3908,N_3848,N_3833);
xor U3909 (N_3909,N_3843,N_3842);
nor U3910 (N_3910,N_3839,N_3866);
nor U3911 (N_3911,N_3841,N_3849);
and U3912 (N_3912,N_3827,N_3856);
and U3913 (N_3913,N_3860,N_3879);
nor U3914 (N_3914,N_3819,N_3877);
or U3915 (N_3915,N_3809,N_3855);
xnor U3916 (N_3916,N_3891,N_3864);
and U3917 (N_3917,N_3889,N_3851);
nand U3918 (N_3918,N_3886,N_3822);
xnor U3919 (N_3919,N_3835,N_3818);
nand U3920 (N_3920,N_3896,N_3898);
nand U3921 (N_3921,N_3895,N_3852);
and U3922 (N_3922,N_3808,N_3844);
nand U3923 (N_3923,N_3894,N_3837);
and U3924 (N_3924,N_3801,N_3825);
nor U3925 (N_3925,N_3840,N_3867);
nor U3926 (N_3926,N_3892,N_3899);
or U3927 (N_3927,N_3884,N_3880);
nor U3928 (N_3928,N_3893,N_3815);
xor U3929 (N_3929,N_3832,N_3823);
or U3930 (N_3930,N_3873,N_3834);
xnor U3931 (N_3931,N_3828,N_3826);
or U3932 (N_3932,N_3811,N_3817);
or U3933 (N_3933,N_3821,N_3876);
or U3934 (N_3934,N_3810,N_3859);
and U3935 (N_3935,N_3897,N_3846);
nand U3936 (N_3936,N_3847,N_3820);
and U3937 (N_3937,N_3885,N_3871);
or U3938 (N_3938,N_3858,N_3869);
and U3939 (N_3939,N_3862,N_3831);
or U3940 (N_3940,N_3816,N_3870);
nand U3941 (N_3941,N_3878,N_3803);
or U3942 (N_3942,N_3829,N_3887);
or U3943 (N_3943,N_3854,N_3888);
and U3944 (N_3944,N_3853,N_3872);
xor U3945 (N_3945,N_3804,N_3875);
nor U3946 (N_3946,N_3883,N_3861);
and U3947 (N_3947,N_3850,N_3830);
and U3948 (N_3948,N_3874,N_3882);
and U3949 (N_3949,N_3800,N_3812);
nand U3950 (N_3950,N_3862,N_3838);
and U3951 (N_3951,N_3891,N_3834);
nor U3952 (N_3952,N_3876,N_3813);
and U3953 (N_3953,N_3829,N_3861);
and U3954 (N_3954,N_3837,N_3864);
nor U3955 (N_3955,N_3897,N_3894);
and U3956 (N_3956,N_3843,N_3810);
and U3957 (N_3957,N_3801,N_3813);
nor U3958 (N_3958,N_3823,N_3827);
nand U3959 (N_3959,N_3833,N_3856);
nor U3960 (N_3960,N_3829,N_3879);
and U3961 (N_3961,N_3834,N_3829);
and U3962 (N_3962,N_3808,N_3851);
and U3963 (N_3963,N_3839,N_3890);
nand U3964 (N_3964,N_3810,N_3886);
nor U3965 (N_3965,N_3864,N_3819);
nor U3966 (N_3966,N_3869,N_3845);
xnor U3967 (N_3967,N_3876,N_3883);
nor U3968 (N_3968,N_3806,N_3898);
xor U3969 (N_3969,N_3892,N_3862);
and U3970 (N_3970,N_3816,N_3892);
xor U3971 (N_3971,N_3848,N_3864);
or U3972 (N_3972,N_3821,N_3816);
and U3973 (N_3973,N_3882,N_3807);
nand U3974 (N_3974,N_3895,N_3892);
xnor U3975 (N_3975,N_3868,N_3851);
nand U3976 (N_3976,N_3800,N_3848);
nor U3977 (N_3977,N_3832,N_3877);
or U3978 (N_3978,N_3806,N_3894);
nor U3979 (N_3979,N_3805,N_3849);
or U3980 (N_3980,N_3805,N_3888);
nor U3981 (N_3981,N_3808,N_3856);
nor U3982 (N_3982,N_3860,N_3861);
and U3983 (N_3983,N_3880,N_3892);
or U3984 (N_3984,N_3840,N_3875);
and U3985 (N_3985,N_3881,N_3817);
nand U3986 (N_3986,N_3831,N_3881);
or U3987 (N_3987,N_3810,N_3840);
nand U3988 (N_3988,N_3898,N_3819);
or U3989 (N_3989,N_3843,N_3846);
nor U3990 (N_3990,N_3808,N_3894);
or U3991 (N_3991,N_3894,N_3863);
or U3992 (N_3992,N_3899,N_3806);
nand U3993 (N_3993,N_3830,N_3812);
and U3994 (N_3994,N_3836,N_3849);
nor U3995 (N_3995,N_3834,N_3882);
nand U3996 (N_3996,N_3834,N_3899);
nor U3997 (N_3997,N_3821,N_3861);
and U3998 (N_3998,N_3806,N_3868);
or U3999 (N_3999,N_3827,N_3836);
nor U4000 (N_4000,N_3963,N_3986);
or U4001 (N_4001,N_3935,N_3911);
xor U4002 (N_4002,N_3999,N_3989);
nand U4003 (N_4003,N_3974,N_3907);
xnor U4004 (N_4004,N_3943,N_3958);
nor U4005 (N_4005,N_3921,N_3924);
nand U4006 (N_4006,N_3933,N_3998);
xnor U4007 (N_4007,N_3917,N_3923);
xor U4008 (N_4008,N_3932,N_3970);
nor U4009 (N_4009,N_3922,N_3903);
or U4010 (N_4010,N_3987,N_3950);
or U4011 (N_4011,N_3995,N_3957);
nand U4012 (N_4012,N_3983,N_3914);
and U4013 (N_4013,N_3956,N_3955);
nor U4014 (N_4014,N_3901,N_3945);
or U4015 (N_4015,N_3908,N_3996);
xor U4016 (N_4016,N_3949,N_3962);
xnor U4017 (N_4017,N_3969,N_3942);
xnor U4018 (N_4018,N_3941,N_3971);
nand U4019 (N_4019,N_3973,N_3991);
or U4020 (N_4020,N_3906,N_3994);
and U4021 (N_4021,N_3925,N_3967);
xor U4022 (N_4022,N_3910,N_3912);
nand U4023 (N_4023,N_3927,N_3988);
nand U4024 (N_4024,N_3959,N_3938);
nor U4025 (N_4025,N_3940,N_3937);
nand U4026 (N_4026,N_3965,N_3936);
xnor U4027 (N_4027,N_3905,N_3972);
nor U4028 (N_4028,N_3930,N_3966);
or U4029 (N_4029,N_3968,N_3928);
or U4030 (N_4030,N_3980,N_3953);
nand U4031 (N_4031,N_3997,N_3992);
or U4032 (N_4032,N_3990,N_3944);
nand U4033 (N_4033,N_3929,N_3920);
or U4034 (N_4034,N_3954,N_3961);
and U4035 (N_4035,N_3916,N_3919);
xor U4036 (N_4036,N_3948,N_3946);
nand U4037 (N_4037,N_3964,N_3926);
nand U4038 (N_4038,N_3952,N_3984);
xnor U4039 (N_4039,N_3981,N_3978);
or U4040 (N_4040,N_3918,N_3909);
nand U4041 (N_4041,N_3947,N_3985);
and U4042 (N_4042,N_3982,N_3951);
nand U4043 (N_4043,N_3939,N_3913);
or U4044 (N_4044,N_3993,N_3934);
nand U4045 (N_4045,N_3900,N_3960);
nand U4046 (N_4046,N_3979,N_3977);
nor U4047 (N_4047,N_3976,N_3915);
nand U4048 (N_4048,N_3975,N_3902);
nor U4049 (N_4049,N_3904,N_3931);
and U4050 (N_4050,N_3983,N_3930);
xnor U4051 (N_4051,N_3908,N_3935);
and U4052 (N_4052,N_3954,N_3921);
nor U4053 (N_4053,N_3977,N_3909);
xor U4054 (N_4054,N_3937,N_3967);
nand U4055 (N_4055,N_3997,N_3933);
xnor U4056 (N_4056,N_3990,N_3974);
nor U4057 (N_4057,N_3954,N_3948);
or U4058 (N_4058,N_3968,N_3902);
or U4059 (N_4059,N_3954,N_3934);
nor U4060 (N_4060,N_3914,N_3958);
nand U4061 (N_4061,N_3905,N_3998);
nor U4062 (N_4062,N_3919,N_3945);
nor U4063 (N_4063,N_3960,N_3964);
xnor U4064 (N_4064,N_3931,N_3994);
and U4065 (N_4065,N_3985,N_3936);
xnor U4066 (N_4066,N_3940,N_3999);
or U4067 (N_4067,N_3918,N_3931);
or U4068 (N_4068,N_3953,N_3988);
xor U4069 (N_4069,N_3986,N_3990);
or U4070 (N_4070,N_3914,N_3987);
nand U4071 (N_4071,N_3969,N_3936);
and U4072 (N_4072,N_3983,N_3985);
nor U4073 (N_4073,N_3935,N_3925);
and U4074 (N_4074,N_3920,N_3997);
xor U4075 (N_4075,N_3987,N_3915);
xnor U4076 (N_4076,N_3900,N_3909);
nor U4077 (N_4077,N_3921,N_3935);
nor U4078 (N_4078,N_3908,N_3959);
nor U4079 (N_4079,N_3941,N_3962);
nand U4080 (N_4080,N_3936,N_3962);
and U4081 (N_4081,N_3944,N_3995);
nand U4082 (N_4082,N_3909,N_3942);
xor U4083 (N_4083,N_3953,N_3970);
xor U4084 (N_4084,N_3983,N_3918);
and U4085 (N_4085,N_3907,N_3931);
or U4086 (N_4086,N_3942,N_3991);
xor U4087 (N_4087,N_3970,N_3914);
nor U4088 (N_4088,N_3921,N_3962);
or U4089 (N_4089,N_3920,N_3966);
xnor U4090 (N_4090,N_3995,N_3966);
xnor U4091 (N_4091,N_3913,N_3917);
xor U4092 (N_4092,N_3955,N_3922);
nand U4093 (N_4093,N_3997,N_3969);
nor U4094 (N_4094,N_3994,N_3955);
xor U4095 (N_4095,N_3906,N_3956);
or U4096 (N_4096,N_3993,N_3927);
or U4097 (N_4097,N_3912,N_3962);
xnor U4098 (N_4098,N_3987,N_3911);
and U4099 (N_4099,N_3997,N_3994);
or U4100 (N_4100,N_4037,N_4010);
or U4101 (N_4101,N_4040,N_4005);
or U4102 (N_4102,N_4086,N_4053);
nand U4103 (N_4103,N_4016,N_4057);
or U4104 (N_4104,N_4050,N_4009);
or U4105 (N_4105,N_4007,N_4004);
xnor U4106 (N_4106,N_4030,N_4041);
nor U4107 (N_4107,N_4008,N_4018);
xor U4108 (N_4108,N_4022,N_4043);
and U4109 (N_4109,N_4074,N_4025);
or U4110 (N_4110,N_4046,N_4036);
and U4111 (N_4111,N_4024,N_4061);
nor U4112 (N_4112,N_4000,N_4003);
nor U4113 (N_4113,N_4035,N_4071);
xnor U4114 (N_4114,N_4048,N_4082);
and U4115 (N_4115,N_4002,N_4027);
nor U4116 (N_4116,N_4012,N_4015);
and U4117 (N_4117,N_4031,N_4094);
and U4118 (N_4118,N_4073,N_4059);
nand U4119 (N_4119,N_4032,N_4044);
or U4120 (N_4120,N_4079,N_4011);
xor U4121 (N_4121,N_4078,N_4014);
and U4122 (N_4122,N_4090,N_4070);
or U4123 (N_4123,N_4063,N_4098);
and U4124 (N_4124,N_4077,N_4069);
nor U4125 (N_4125,N_4034,N_4042);
xor U4126 (N_4126,N_4029,N_4020);
or U4127 (N_4127,N_4092,N_4064);
or U4128 (N_4128,N_4023,N_4072);
or U4129 (N_4129,N_4038,N_4095);
nor U4130 (N_4130,N_4013,N_4099);
nor U4131 (N_4131,N_4055,N_4084);
and U4132 (N_4132,N_4066,N_4028);
and U4133 (N_4133,N_4096,N_4075);
nand U4134 (N_4134,N_4093,N_4087);
xor U4135 (N_4135,N_4017,N_4056);
nor U4136 (N_4136,N_4047,N_4076);
or U4137 (N_4137,N_4058,N_4068);
and U4138 (N_4138,N_4067,N_4054);
and U4139 (N_4139,N_4019,N_4045);
or U4140 (N_4140,N_4097,N_4083);
nor U4141 (N_4141,N_4051,N_4033);
or U4142 (N_4142,N_4049,N_4091);
xor U4143 (N_4143,N_4085,N_4001);
and U4144 (N_4144,N_4081,N_4065);
nand U4145 (N_4145,N_4062,N_4006);
or U4146 (N_4146,N_4039,N_4060);
nor U4147 (N_4147,N_4089,N_4026);
or U4148 (N_4148,N_4088,N_4052);
or U4149 (N_4149,N_4080,N_4021);
or U4150 (N_4150,N_4004,N_4082);
xnor U4151 (N_4151,N_4016,N_4075);
nand U4152 (N_4152,N_4035,N_4068);
xnor U4153 (N_4153,N_4084,N_4013);
nor U4154 (N_4154,N_4057,N_4052);
xor U4155 (N_4155,N_4080,N_4042);
or U4156 (N_4156,N_4038,N_4042);
or U4157 (N_4157,N_4097,N_4069);
and U4158 (N_4158,N_4037,N_4050);
xnor U4159 (N_4159,N_4014,N_4064);
and U4160 (N_4160,N_4072,N_4008);
and U4161 (N_4161,N_4054,N_4077);
and U4162 (N_4162,N_4029,N_4024);
nor U4163 (N_4163,N_4076,N_4082);
and U4164 (N_4164,N_4073,N_4090);
nor U4165 (N_4165,N_4010,N_4027);
nand U4166 (N_4166,N_4016,N_4047);
nor U4167 (N_4167,N_4068,N_4072);
and U4168 (N_4168,N_4014,N_4088);
or U4169 (N_4169,N_4016,N_4097);
or U4170 (N_4170,N_4031,N_4066);
and U4171 (N_4171,N_4034,N_4097);
xnor U4172 (N_4172,N_4085,N_4062);
nor U4173 (N_4173,N_4053,N_4031);
or U4174 (N_4174,N_4039,N_4002);
xnor U4175 (N_4175,N_4057,N_4027);
nand U4176 (N_4176,N_4018,N_4086);
nand U4177 (N_4177,N_4089,N_4075);
and U4178 (N_4178,N_4052,N_4067);
xnor U4179 (N_4179,N_4081,N_4098);
nand U4180 (N_4180,N_4087,N_4057);
xnor U4181 (N_4181,N_4056,N_4060);
xor U4182 (N_4182,N_4060,N_4035);
nor U4183 (N_4183,N_4070,N_4053);
nor U4184 (N_4184,N_4089,N_4055);
nand U4185 (N_4185,N_4090,N_4057);
and U4186 (N_4186,N_4001,N_4019);
xor U4187 (N_4187,N_4093,N_4066);
nor U4188 (N_4188,N_4045,N_4088);
nor U4189 (N_4189,N_4032,N_4029);
and U4190 (N_4190,N_4025,N_4098);
nor U4191 (N_4191,N_4048,N_4005);
or U4192 (N_4192,N_4039,N_4071);
xor U4193 (N_4193,N_4025,N_4011);
xor U4194 (N_4194,N_4089,N_4095);
xor U4195 (N_4195,N_4004,N_4069);
or U4196 (N_4196,N_4008,N_4007);
xor U4197 (N_4197,N_4029,N_4074);
nand U4198 (N_4198,N_4004,N_4038);
and U4199 (N_4199,N_4098,N_4097);
nand U4200 (N_4200,N_4130,N_4177);
or U4201 (N_4201,N_4142,N_4192);
and U4202 (N_4202,N_4126,N_4162);
nand U4203 (N_4203,N_4128,N_4140);
or U4204 (N_4204,N_4199,N_4188);
nand U4205 (N_4205,N_4152,N_4138);
and U4206 (N_4206,N_4191,N_4182);
nor U4207 (N_4207,N_4195,N_4119);
nor U4208 (N_4208,N_4186,N_4171);
nand U4209 (N_4209,N_4127,N_4106);
nor U4210 (N_4210,N_4159,N_4144);
nand U4211 (N_4211,N_4150,N_4133);
or U4212 (N_4212,N_4143,N_4170);
or U4213 (N_4213,N_4103,N_4167);
and U4214 (N_4214,N_4173,N_4181);
xnor U4215 (N_4215,N_4109,N_4184);
and U4216 (N_4216,N_4116,N_4120);
and U4217 (N_4217,N_4125,N_4166);
and U4218 (N_4218,N_4132,N_4165);
xor U4219 (N_4219,N_4175,N_4131);
or U4220 (N_4220,N_4174,N_4198);
and U4221 (N_4221,N_4164,N_4112);
nand U4222 (N_4222,N_4169,N_4108);
xnor U4223 (N_4223,N_4100,N_4118);
xor U4224 (N_4224,N_4123,N_4161);
nor U4225 (N_4225,N_4141,N_4190);
or U4226 (N_4226,N_4113,N_4104);
nand U4227 (N_4227,N_4136,N_4135);
nor U4228 (N_4228,N_4151,N_4115);
xor U4229 (N_4229,N_4160,N_4155);
or U4230 (N_4230,N_4197,N_4137);
nand U4231 (N_4231,N_4156,N_4179);
nor U4232 (N_4232,N_4111,N_4180);
and U4233 (N_4233,N_4110,N_4193);
and U4234 (N_4234,N_4158,N_4153);
nor U4235 (N_4235,N_4107,N_4185);
or U4236 (N_4236,N_4154,N_4168);
xor U4237 (N_4237,N_4178,N_4148);
and U4238 (N_4238,N_4157,N_4176);
and U4239 (N_4239,N_4139,N_4117);
nor U4240 (N_4240,N_4145,N_4194);
xnor U4241 (N_4241,N_4121,N_4163);
xnor U4242 (N_4242,N_4149,N_4196);
or U4243 (N_4243,N_4134,N_4122);
xor U4244 (N_4244,N_4101,N_4129);
xor U4245 (N_4245,N_4146,N_4124);
nand U4246 (N_4246,N_4189,N_4147);
or U4247 (N_4247,N_4187,N_4105);
or U4248 (N_4248,N_4114,N_4102);
or U4249 (N_4249,N_4183,N_4172);
nand U4250 (N_4250,N_4187,N_4191);
nor U4251 (N_4251,N_4162,N_4189);
xnor U4252 (N_4252,N_4143,N_4122);
and U4253 (N_4253,N_4134,N_4136);
nand U4254 (N_4254,N_4118,N_4171);
nor U4255 (N_4255,N_4171,N_4182);
xnor U4256 (N_4256,N_4151,N_4105);
nor U4257 (N_4257,N_4149,N_4110);
nand U4258 (N_4258,N_4128,N_4175);
and U4259 (N_4259,N_4151,N_4163);
nor U4260 (N_4260,N_4114,N_4186);
nor U4261 (N_4261,N_4185,N_4180);
xor U4262 (N_4262,N_4140,N_4187);
nor U4263 (N_4263,N_4170,N_4180);
xnor U4264 (N_4264,N_4166,N_4164);
and U4265 (N_4265,N_4124,N_4162);
nor U4266 (N_4266,N_4190,N_4134);
and U4267 (N_4267,N_4159,N_4103);
and U4268 (N_4268,N_4169,N_4145);
nor U4269 (N_4269,N_4117,N_4112);
xnor U4270 (N_4270,N_4144,N_4168);
and U4271 (N_4271,N_4106,N_4157);
nand U4272 (N_4272,N_4121,N_4141);
and U4273 (N_4273,N_4118,N_4179);
xor U4274 (N_4274,N_4130,N_4112);
xnor U4275 (N_4275,N_4182,N_4115);
or U4276 (N_4276,N_4118,N_4144);
and U4277 (N_4277,N_4138,N_4133);
and U4278 (N_4278,N_4110,N_4172);
or U4279 (N_4279,N_4117,N_4191);
xor U4280 (N_4280,N_4112,N_4121);
or U4281 (N_4281,N_4119,N_4183);
xnor U4282 (N_4282,N_4116,N_4105);
nor U4283 (N_4283,N_4127,N_4199);
nor U4284 (N_4284,N_4113,N_4161);
nand U4285 (N_4285,N_4134,N_4141);
nor U4286 (N_4286,N_4177,N_4163);
nor U4287 (N_4287,N_4125,N_4168);
nand U4288 (N_4288,N_4180,N_4154);
nor U4289 (N_4289,N_4101,N_4167);
and U4290 (N_4290,N_4143,N_4165);
nand U4291 (N_4291,N_4114,N_4108);
nor U4292 (N_4292,N_4173,N_4126);
and U4293 (N_4293,N_4159,N_4194);
nor U4294 (N_4294,N_4193,N_4139);
xor U4295 (N_4295,N_4198,N_4185);
xor U4296 (N_4296,N_4115,N_4167);
nor U4297 (N_4297,N_4181,N_4150);
xnor U4298 (N_4298,N_4168,N_4170);
nand U4299 (N_4299,N_4195,N_4116);
and U4300 (N_4300,N_4215,N_4259);
xor U4301 (N_4301,N_4288,N_4230);
or U4302 (N_4302,N_4278,N_4260);
or U4303 (N_4303,N_4249,N_4258);
nand U4304 (N_4304,N_4236,N_4297);
nand U4305 (N_4305,N_4248,N_4290);
nor U4306 (N_4306,N_4298,N_4267);
nand U4307 (N_4307,N_4294,N_4211);
xnor U4308 (N_4308,N_4292,N_4268);
and U4309 (N_4309,N_4242,N_4206);
or U4310 (N_4310,N_4254,N_4296);
or U4311 (N_4311,N_4270,N_4272);
nor U4312 (N_4312,N_4266,N_4223);
nand U4313 (N_4313,N_4205,N_4280);
and U4314 (N_4314,N_4276,N_4226);
or U4315 (N_4315,N_4253,N_4228);
xor U4316 (N_4316,N_4208,N_4295);
nand U4317 (N_4317,N_4289,N_4257);
and U4318 (N_4318,N_4227,N_4293);
xor U4319 (N_4319,N_4202,N_4201);
and U4320 (N_4320,N_4274,N_4240);
or U4321 (N_4321,N_4221,N_4222);
nor U4322 (N_4322,N_4216,N_4243);
xor U4323 (N_4323,N_4250,N_4233);
xnor U4324 (N_4324,N_4209,N_4286);
nand U4325 (N_4325,N_4231,N_4265);
nor U4326 (N_4326,N_4203,N_4252);
or U4327 (N_4327,N_4282,N_4234);
xnor U4328 (N_4328,N_4291,N_4251);
and U4329 (N_4329,N_4281,N_4247);
nand U4330 (N_4330,N_4264,N_4207);
xnor U4331 (N_4331,N_4220,N_4244);
nor U4332 (N_4332,N_4273,N_4269);
nand U4333 (N_4333,N_4214,N_4279);
xnor U4334 (N_4334,N_4241,N_4218);
nand U4335 (N_4335,N_4262,N_4237);
xnor U4336 (N_4336,N_4275,N_4246);
xnor U4337 (N_4337,N_4287,N_4225);
nor U4338 (N_4338,N_4229,N_4239);
xor U4339 (N_4339,N_4285,N_4217);
xor U4340 (N_4340,N_4219,N_4213);
or U4341 (N_4341,N_4284,N_4255);
xnor U4342 (N_4342,N_4238,N_4224);
and U4343 (N_4343,N_4277,N_4210);
nor U4344 (N_4344,N_4235,N_4256);
or U4345 (N_4345,N_4263,N_4204);
nand U4346 (N_4346,N_4232,N_4212);
xor U4347 (N_4347,N_4271,N_4261);
and U4348 (N_4348,N_4299,N_4283);
nor U4349 (N_4349,N_4200,N_4245);
nor U4350 (N_4350,N_4283,N_4274);
or U4351 (N_4351,N_4218,N_4233);
and U4352 (N_4352,N_4259,N_4234);
and U4353 (N_4353,N_4207,N_4244);
nand U4354 (N_4354,N_4219,N_4237);
or U4355 (N_4355,N_4260,N_4259);
nand U4356 (N_4356,N_4289,N_4225);
nor U4357 (N_4357,N_4268,N_4233);
or U4358 (N_4358,N_4299,N_4251);
nor U4359 (N_4359,N_4259,N_4236);
nand U4360 (N_4360,N_4223,N_4262);
or U4361 (N_4361,N_4235,N_4250);
nand U4362 (N_4362,N_4232,N_4241);
nor U4363 (N_4363,N_4228,N_4235);
and U4364 (N_4364,N_4289,N_4226);
nand U4365 (N_4365,N_4210,N_4265);
or U4366 (N_4366,N_4282,N_4204);
or U4367 (N_4367,N_4284,N_4258);
or U4368 (N_4368,N_4295,N_4235);
and U4369 (N_4369,N_4285,N_4226);
or U4370 (N_4370,N_4244,N_4227);
xnor U4371 (N_4371,N_4264,N_4217);
or U4372 (N_4372,N_4240,N_4217);
and U4373 (N_4373,N_4281,N_4284);
or U4374 (N_4374,N_4238,N_4287);
nand U4375 (N_4375,N_4222,N_4217);
nor U4376 (N_4376,N_4201,N_4249);
nor U4377 (N_4377,N_4268,N_4281);
nand U4378 (N_4378,N_4279,N_4286);
xor U4379 (N_4379,N_4211,N_4263);
xor U4380 (N_4380,N_4272,N_4275);
and U4381 (N_4381,N_4221,N_4211);
nor U4382 (N_4382,N_4238,N_4291);
or U4383 (N_4383,N_4225,N_4224);
or U4384 (N_4384,N_4281,N_4252);
and U4385 (N_4385,N_4231,N_4232);
and U4386 (N_4386,N_4294,N_4298);
or U4387 (N_4387,N_4222,N_4254);
nand U4388 (N_4388,N_4290,N_4278);
xor U4389 (N_4389,N_4259,N_4277);
and U4390 (N_4390,N_4218,N_4246);
xnor U4391 (N_4391,N_4249,N_4266);
xnor U4392 (N_4392,N_4265,N_4298);
nand U4393 (N_4393,N_4223,N_4269);
or U4394 (N_4394,N_4257,N_4298);
nand U4395 (N_4395,N_4246,N_4245);
nand U4396 (N_4396,N_4283,N_4225);
nand U4397 (N_4397,N_4275,N_4274);
or U4398 (N_4398,N_4209,N_4262);
xnor U4399 (N_4399,N_4258,N_4264);
and U4400 (N_4400,N_4342,N_4307);
xor U4401 (N_4401,N_4371,N_4399);
nor U4402 (N_4402,N_4340,N_4329);
or U4403 (N_4403,N_4373,N_4352);
xor U4404 (N_4404,N_4345,N_4368);
or U4405 (N_4405,N_4360,N_4387);
xnor U4406 (N_4406,N_4395,N_4322);
xnor U4407 (N_4407,N_4300,N_4388);
nand U4408 (N_4408,N_4335,N_4364);
nand U4409 (N_4409,N_4353,N_4386);
xnor U4410 (N_4410,N_4319,N_4372);
and U4411 (N_4411,N_4347,N_4376);
or U4412 (N_4412,N_4325,N_4312);
xnor U4413 (N_4413,N_4354,N_4332);
xnor U4414 (N_4414,N_4357,N_4370);
or U4415 (N_4415,N_4350,N_4391);
xor U4416 (N_4416,N_4301,N_4378);
and U4417 (N_4417,N_4381,N_4383);
or U4418 (N_4418,N_4308,N_4306);
nand U4419 (N_4419,N_4356,N_4330);
and U4420 (N_4420,N_4361,N_4334);
nand U4421 (N_4421,N_4321,N_4327);
or U4422 (N_4422,N_4393,N_4346);
xnor U4423 (N_4423,N_4315,N_4389);
nand U4424 (N_4424,N_4310,N_4358);
or U4425 (N_4425,N_4366,N_4365);
or U4426 (N_4426,N_4323,N_4328);
or U4427 (N_4427,N_4359,N_4318);
nand U4428 (N_4428,N_4343,N_4336);
nor U4429 (N_4429,N_4397,N_4331);
or U4430 (N_4430,N_4324,N_4320);
xor U4431 (N_4431,N_4398,N_4379);
nand U4432 (N_4432,N_4384,N_4374);
nor U4433 (N_4433,N_4304,N_4305);
nand U4434 (N_4434,N_4349,N_4369);
xor U4435 (N_4435,N_4348,N_4333);
or U4436 (N_4436,N_4392,N_4311);
or U4437 (N_4437,N_4351,N_4394);
nand U4438 (N_4438,N_4385,N_4338);
nor U4439 (N_4439,N_4344,N_4337);
nand U4440 (N_4440,N_4363,N_4390);
and U4441 (N_4441,N_4326,N_4355);
nor U4442 (N_4442,N_4317,N_4375);
and U4443 (N_4443,N_4377,N_4396);
nor U4444 (N_4444,N_4314,N_4339);
and U4445 (N_4445,N_4341,N_4309);
or U4446 (N_4446,N_4316,N_4362);
and U4447 (N_4447,N_4302,N_4380);
nor U4448 (N_4448,N_4303,N_4382);
and U4449 (N_4449,N_4313,N_4367);
xor U4450 (N_4450,N_4350,N_4305);
or U4451 (N_4451,N_4303,N_4388);
nand U4452 (N_4452,N_4342,N_4383);
nor U4453 (N_4453,N_4313,N_4331);
xor U4454 (N_4454,N_4334,N_4388);
and U4455 (N_4455,N_4395,N_4325);
nand U4456 (N_4456,N_4357,N_4399);
nand U4457 (N_4457,N_4326,N_4311);
or U4458 (N_4458,N_4390,N_4377);
nor U4459 (N_4459,N_4312,N_4346);
and U4460 (N_4460,N_4325,N_4338);
nor U4461 (N_4461,N_4378,N_4341);
nand U4462 (N_4462,N_4333,N_4398);
or U4463 (N_4463,N_4312,N_4379);
or U4464 (N_4464,N_4318,N_4368);
nor U4465 (N_4465,N_4345,N_4374);
nand U4466 (N_4466,N_4314,N_4391);
or U4467 (N_4467,N_4383,N_4370);
nand U4468 (N_4468,N_4306,N_4376);
and U4469 (N_4469,N_4365,N_4349);
xnor U4470 (N_4470,N_4303,N_4326);
nor U4471 (N_4471,N_4322,N_4329);
nor U4472 (N_4472,N_4333,N_4357);
and U4473 (N_4473,N_4321,N_4346);
and U4474 (N_4474,N_4356,N_4361);
nor U4475 (N_4475,N_4332,N_4326);
or U4476 (N_4476,N_4335,N_4315);
xnor U4477 (N_4477,N_4310,N_4325);
or U4478 (N_4478,N_4383,N_4333);
nor U4479 (N_4479,N_4360,N_4346);
nor U4480 (N_4480,N_4333,N_4312);
nand U4481 (N_4481,N_4395,N_4332);
nand U4482 (N_4482,N_4321,N_4340);
xor U4483 (N_4483,N_4351,N_4329);
nand U4484 (N_4484,N_4319,N_4317);
nor U4485 (N_4485,N_4377,N_4333);
or U4486 (N_4486,N_4311,N_4302);
or U4487 (N_4487,N_4391,N_4334);
nand U4488 (N_4488,N_4390,N_4366);
or U4489 (N_4489,N_4318,N_4302);
and U4490 (N_4490,N_4306,N_4357);
or U4491 (N_4491,N_4306,N_4301);
nor U4492 (N_4492,N_4346,N_4304);
nand U4493 (N_4493,N_4329,N_4374);
xor U4494 (N_4494,N_4371,N_4340);
and U4495 (N_4495,N_4379,N_4397);
nand U4496 (N_4496,N_4399,N_4365);
nand U4497 (N_4497,N_4305,N_4393);
xnor U4498 (N_4498,N_4332,N_4316);
and U4499 (N_4499,N_4341,N_4307);
nor U4500 (N_4500,N_4428,N_4492);
nand U4501 (N_4501,N_4448,N_4493);
nor U4502 (N_4502,N_4478,N_4435);
nor U4503 (N_4503,N_4452,N_4429);
and U4504 (N_4504,N_4461,N_4446);
xnor U4505 (N_4505,N_4410,N_4472);
xor U4506 (N_4506,N_4409,N_4479);
nor U4507 (N_4507,N_4496,N_4473);
nor U4508 (N_4508,N_4484,N_4455);
nand U4509 (N_4509,N_4457,N_4412);
and U4510 (N_4510,N_4453,N_4405);
xor U4511 (N_4511,N_4474,N_4463);
xnor U4512 (N_4512,N_4411,N_4456);
nand U4513 (N_4513,N_4494,N_4481);
nor U4514 (N_4514,N_4407,N_4499);
nand U4515 (N_4515,N_4486,N_4424);
nand U4516 (N_4516,N_4400,N_4430);
nor U4517 (N_4517,N_4498,N_4449);
and U4518 (N_4518,N_4417,N_4459);
and U4519 (N_4519,N_4489,N_4445);
xor U4520 (N_4520,N_4427,N_4482);
nor U4521 (N_4521,N_4423,N_4433);
or U4522 (N_4522,N_4415,N_4416);
and U4523 (N_4523,N_4434,N_4404);
and U4524 (N_4524,N_4476,N_4485);
and U4525 (N_4525,N_4418,N_4437);
xor U4526 (N_4526,N_4419,N_4439);
and U4527 (N_4527,N_4471,N_4401);
and U4528 (N_4528,N_4444,N_4441);
nor U4529 (N_4529,N_4464,N_4477);
and U4530 (N_4530,N_4413,N_4432);
and U4531 (N_4531,N_4497,N_4425);
and U4532 (N_4532,N_4470,N_4402);
or U4533 (N_4533,N_4462,N_4440);
or U4534 (N_4534,N_4431,N_4460);
and U4535 (N_4535,N_4403,N_4480);
xor U4536 (N_4536,N_4450,N_4422);
and U4537 (N_4537,N_4458,N_4469);
xor U4538 (N_4538,N_4443,N_4436);
nand U4539 (N_4539,N_4447,N_4414);
or U4540 (N_4540,N_4475,N_4483);
or U4541 (N_4541,N_4468,N_4490);
xor U4542 (N_4542,N_4454,N_4466);
nor U4543 (N_4543,N_4491,N_4421);
nor U4544 (N_4544,N_4426,N_4451);
or U4545 (N_4545,N_4420,N_4408);
nor U4546 (N_4546,N_4487,N_4438);
and U4547 (N_4547,N_4495,N_4467);
nand U4548 (N_4548,N_4488,N_4406);
nand U4549 (N_4549,N_4465,N_4442);
and U4550 (N_4550,N_4494,N_4486);
and U4551 (N_4551,N_4463,N_4415);
or U4552 (N_4552,N_4467,N_4479);
or U4553 (N_4553,N_4426,N_4458);
and U4554 (N_4554,N_4442,N_4486);
xor U4555 (N_4555,N_4454,N_4487);
and U4556 (N_4556,N_4454,N_4497);
or U4557 (N_4557,N_4441,N_4438);
and U4558 (N_4558,N_4490,N_4402);
nand U4559 (N_4559,N_4436,N_4474);
and U4560 (N_4560,N_4474,N_4429);
nor U4561 (N_4561,N_4490,N_4441);
and U4562 (N_4562,N_4491,N_4438);
xnor U4563 (N_4563,N_4444,N_4446);
and U4564 (N_4564,N_4454,N_4485);
or U4565 (N_4565,N_4449,N_4488);
nand U4566 (N_4566,N_4400,N_4418);
or U4567 (N_4567,N_4405,N_4492);
xor U4568 (N_4568,N_4434,N_4492);
nor U4569 (N_4569,N_4499,N_4476);
nor U4570 (N_4570,N_4412,N_4447);
or U4571 (N_4571,N_4447,N_4434);
nand U4572 (N_4572,N_4474,N_4499);
or U4573 (N_4573,N_4459,N_4456);
xnor U4574 (N_4574,N_4471,N_4494);
and U4575 (N_4575,N_4447,N_4437);
nand U4576 (N_4576,N_4490,N_4464);
xnor U4577 (N_4577,N_4446,N_4420);
nand U4578 (N_4578,N_4487,N_4451);
and U4579 (N_4579,N_4434,N_4414);
and U4580 (N_4580,N_4425,N_4435);
nor U4581 (N_4581,N_4456,N_4439);
and U4582 (N_4582,N_4477,N_4440);
or U4583 (N_4583,N_4470,N_4492);
and U4584 (N_4584,N_4421,N_4482);
nand U4585 (N_4585,N_4499,N_4411);
nor U4586 (N_4586,N_4412,N_4462);
xnor U4587 (N_4587,N_4481,N_4404);
nand U4588 (N_4588,N_4401,N_4488);
xor U4589 (N_4589,N_4434,N_4473);
and U4590 (N_4590,N_4485,N_4437);
nor U4591 (N_4591,N_4471,N_4438);
and U4592 (N_4592,N_4457,N_4431);
xnor U4593 (N_4593,N_4401,N_4464);
xnor U4594 (N_4594,N_4480,N_4448);
or U4595 (N_4595,N_4448,N_4429);
or U4596 (N_4596,N_4444,N_4417);
nor U4597 (N_4597,N_4497,N_4469);
or U4598 (N_4598,N_4406,N_4445);
and U4599 (N_4599,N_4420,N_4449);
nor U4600 (N_4600,N_4566,N_4564);
nand U4601 (N_4601,N_4568,N_4562);
nand U4602 (N_4602,N_4529,N_4575);
or U4603 (N_4603,N_4527,N_4550);
xnor U4604 (N_4604,N_4547,N_4573);
nor U4605 (N_4605,N_4531,N_4509);
or U4606 (N_4606,N_4572,N_4544);
xor U4607 (N_4607,N_4511,N_4570);
nor U4608 (N_4608,N_4596,N_4519);
or U4609 (N_4609,N_4538,N_4551);
or U4610 (N_4610,N_4589,N_4567);
or U4611 (N_4611,N_4552,N_4591);
nor U4612 (N_4612,N_4534,N_4579);
and U4613 (N_4613,N_4555,N_4599);
nor U4614 (N_4614,N_4588,N_4530);
or U4615 (N_4615,N_4597,N_4593);
or U4616 (N_4616,N_4574,N_4561);
xor U4617 (N_4617,N_4520,N_4554);
and U4618 (N_4618,N_4517,N_4576);
nor U4619 (N_4619,N_4585,N_4523);
and U4620 (N_4620,N_4540,N_4556);
xor U4621 (N_4621,N_4553,N_4542);
nand U4622 (N_4622,N_4533,N_4512);
nand U4623 (N_4623,N_4528,N_4515);
xor U4624 (N_4624,N_4595,N_4543);
nand U4625 (N_4625,N_4569,N_4581);
xnor U4626 (N_4626,N_4526,N_4563);
xor U4627 (N_4627,N_4598,N_4522);
xor U4628 (N_4628,N_4587,N_4514);
nand U4629 (N_4629,N_4541,N_4504);
nor U4630 (N_4630,N_4505,N_4594);
nand U4631 (N_4631,N_4560,N_4586);
nor U4632 (N_4632,N_4508,N_4592);
nor U4633 (N_4633,N_4500,N_4532);
and U4634 (N_4634,N_4536,N_4545);
or U4635 (N_4635,N_4513,N_4583);
and U4636 (N_4636,N_4571,N_4578);
xnor U4637 (N_4637,N_4503,N_4525);
nand U4638 (N_4638,N_4584,N_4501);
or U4639 (N_4639,N_4502,N_4559);
and U4640 (N_4640,N_4516,N_4548);
and U4641 (N_4641,N_4535,N_4565);
nor U4642 (N_4642,N_4549,N_4580);
and U4643 (N_4643,N_4507,N_4539);
and U4644 (N_4644,N_4518,N_4546);
and U4645 (N_4645,N_4521,N_4590);
or U4646 (N_4646,N_4506,N_4582);
nor U4647 (N_4647,N_4537,N_4524);
and U4648 (N_4648,N_4577,N_4510);
or U4649 (N_4649,N_4558,N_4557);
or U4650 (N_4650,N_4595,N_4536);
and U4651 (N_4651,N_4594,N_4575);
nand U4652 (N_4652,N_4566,N_4540);
and U4653 (N_4653,N_4508,N_4519);
nand U4654 (N_4654,N_4568,N_4563);
or U4655 (N_4655,N_4537,N_4593);
and U4656 (N_4656,N_4585,N_4540);
nor U4657 (N_4657,N_4565,N_4504);
nor U4658 (N_4658,N_4518,N_4569);
nor U4659 (N_4659,N_4577,N_4507);
nand U4660 (N_4660,N_4537,N_4529);
xnor U4661 (N_4661,N_4535,N_4591);
xor U4662 (N_4662,N_4562,N_4516);
nand U4663 (N_4663,N_4530,N_4566);
or U4664 (N_4664,N_4581,N_4547);
xnor U4665 (N_4665,N_4548,N_4518);
or U4666 (N_4666,N_4516,N_4531);
nand U4667 (N_4667,N_4504,N_4523);
and U4668 (N_4668,N_4568,N_4500);
nor U4669 (N_4669,N_4598,N_4571);
and U4670 (N_4670,N_4583,N_4535);
and U4671 (N_4671,N_4543,N_4537);
and U4672 (N_4672,N_4599,N_4518);
or U4673 (N_4673,N_4530,N_4547);
or U4674 (N_4674,N_4552,N_4574);
xor U4675 (N_4675,N_4560,N_4575);
or U4676 (N_4676,N_4516,N_4583);
xnor U4677 (N_4677,N_4538,N_4571);
nor U4678 (N_4678,N_4535,N_4556);
and U4679 (N_4679,N_4511,N_4514);
xnor U4680 (N_4680,N_4550,N_4562);
or U4681 (N_4681,N_4592,N_4582);
nand U4682 (N_4682,N_4566,N_4523);
xor U4683 (N_4683,N_4561,N_4552);
and U4684 (N_4684,N_4505,N_4537);
xor U4685 (N_4685,N_4532,N_4514);
nand U4686 (N_4686,N_4505,N_4572);
nand U4687 (N_4687,N_4525,N_4572);
xnor U4688 (N_4688,N_4547,N_4593);
nand U4689 (N_4689,N_4536,N_4534);
xor U4690 (N_4690,N_4566,N_4500);
and U4691 (N_4691,N_4546,N_4589);
and U4692 (N_4692,N_4587,N_4532);
nand U4693 (N_4693,N_4520,N_4560);
nand U4694 (N_4694,N_4508,N_4588);
nor U4695 (N_4695,N_4556,N_4588);
nor U4696 (N_4696,N_4516,N_4580);
nand U4697 (N_4697,N_4564,N_4582);
nor U4698 (N_4698,N_4571,N_4528);
nor U4699 (N_4699,N_4565,N_4557);
or U4700 (N_4700,N_4669,N_4618);
nor U4701 (N_4701,N_4625,N_4640);
nand U4702 (N_4702,N_4678,N_4606);
nor U4703 (N_4703,N_4603,N_4639);
nor U4704 (N_4704,N_4673,N_4628);
nor U4705 (N_4705,N_4649,N_4605);
xnor U4706 (N_4706,N_4680,N_4665);
nand U4707 (N_4707,N_4683,N_4686);
nand U4708 (N_4708,N_4613,N_4672);
and U4709 (N_4709,N_4635,N_4646);
and U4710 (N_4710,N_4634,N_4632);
nand U4711 (N_4711,N_4664,N_4647);
nand U4712 (N_4712,N_4677,N_4623);
nor U4713 (N_4713,N_4629,N_4653);
and U4714 (N_4714,N_4654,N_4601);
nand U4715 (N_4715,N_4687,N_4690);
nor U4716 (N_4716,N_4688,N_4676);
nand U4717 (N_4717,N_4663,N_4656);
nand U4718 (N_4718,N_4695,N_4626);
nand U4719 (N_4719,N_4636,N_4631);
nor U4720 (N_4720,N_4696,N_4622);
or U4721 (N_4721,N_4602,N_4621);
xor U4722 (N_4722,N_4681,N_4694);
and U4723 (N_4723,N_4652,N_4645);
and U4724 (N_4724,N_4668,N_4644);
or U4725 (N_4725,N_4643,N_4682);
nand U4726 (N_4726,N_4659,N_4692);
or U4727 (N_4727,N_4671,N_4662);
and U4728 (N_4728,N_4675,N_4648);
nor U4729 (N_4729,N_4638,N_4661);
nand U4730 (N_4730,N_4679,N_4615);
or U4731 (N_4731,N_4611,N_4617);
nor U4732 (N_4732,N_4699,N_4641);
and U4733 (N_4733,N_4689,N_4612);
xor U4734 (N_4734,N_4666,N_4658);
nand U4735 (N_4735,N_4651,N_4684);
xor U4736 (N_4736,N_4697,N_4650);
or U4737 (N_4737,N_4616,N_4674);
and U4738 (N_4738,N_4620,N_4619);
nand U4739 (N_4739,N_4633,N_4630);
and U4740 (N_4740,N_4667,N_4607);
nor U4741 (N_4741,N_4604,N_4624);
xnor U4742 (N_4742,N_4660,N_4608);
nor U4743 (N_4743,N_4610,N_4600);
or U4744 (N_4744,N_4670,N_4698);
or U4745 (N_4745,N_4637,N_4655);
xor U4746 (N_4746,N_4642,N_4657);
nor U4747 (N_4747,N_4693,N_4614);
nand U4748 (N_4748,N_4691,N_4609);
xor U4749 (N_4749,N_4685,N_4627);
nand U4750 (N_4750,N_4603,N_4622);
nor U4751 (N_4751,N_4658,N_4627);
nand U4752 (N_4752,N_4669,N_4691);
xor U4753 (N_4753,N_4680,N_4675);
xnor U4754 (N_4754,N_4611,N_4622);
and U4755 (N_4755,N_4611,N_4602);
nand U4756 (N_4756,N_4683,N_4671);
or U4757 (N_4757,N_4671,N_4652);
nand U4758 (N_4758,N_4680,N_4669);
and U4759 (N_4759,N_4697,N_4633);
nand U4760 (N_4760,N_4623,N_4669);
nand U4761 (N_4761,N_4610,N_4612);
nand U4762 (N_4762,N_4686,N_4673);
and U4763 (N_4763,N_4650,N_4678);
and U4764 (N_4764,N_4665,N_4608);
nor U4765 (N_4765,N_4667,N_4674);
or U4766 (N_4766,N_4636,N_4606);
nand U4767 (N_4767,N_4644,N_4624);
and U4768 (N_4768,N_4627,N_4628);
and U4769 (N_4769,N_4696,N_4610);
or U4770 (N_4770,N_4648,N_4622);
nor U4771 (N_4771,N_4697,N_4689);
xor U4772 (N_4772,N_4639,N_4686);
xor U4773 (N_4773,N_4665,N_4666);
or U4774 (N_4774,N_4646,N_4601);
xor U4775 (N_4775,N_4618,N_4607);
nand U4776 (N_4776,N_4668,N_4634);
or U4777 (N_4777,N_4611,N_4680);
nand U4778 (N_4778,N_4606,N_4635);
nand U4779 (N_4779,N_4610,N_4693);
and U4780 (N_4780,N_4629,N_4652);
nand U4781 (N_4781,N_4692,N_4651);
nand U4782 (N_4782,N_4668,N_4654);
nor U4783 (N_4783,N_4645,N_4659);
and U4784 (N_4784,N_4633,N_4610);
nand U4785 (N_4785,N_4633,N_4695);
nor U4786 (N_4786,N_4696,N_4679);
or U4787 (N_4787,N_4690,N_4623);
and U4788 (N_4788,N_4627,N_4612);
nand U4789 (N_4789,N_4632,N_4670);
xnor U4790 (N_4790,N_4669,N_4672);
nor U4791 (N_4791,N_4604,N_4667);
or U4792 (N_4792,N_4675,N_4685);
or U4793 (N_4793,N_4601,N_4645);
nand U4794 (N_4794,N_4687,N_4683);
nor U4795 (N_4795,N_4611,N_4643);
or U4796 (N_4796,N_4655,N_4620);
xor U4797 (N_4797,N_4612,N_4624);
nand U4798 (N_4798,N_4690,N_4645);
or U4799 (N_4799,N_4624,N_4636);
and U4800 (N_4800,N_4777,N_4746);
or U4801 (N_4801,N_4710,N_4780);
nor U4802 (N_4802,N_4721,N_4718);
and U4803 (N_4803,N_4792,N_4707);
nor U4804 (N_4804,N_4788,N_4761);
and U4805 (N_4805,N_4752,N_4742);
nand U4806 (N_4806,N_4776,N_4741);
or U4807 (N_4807,N_4702,N_4728);
and U4808 (N_4808,N_4796,N_4708);
nor U4809 (N_4809,N_4799,N_4745);
nand U4810 (N_4810,N_4743,N_4713);
nand U4811 (N_4811,N_4724,N_4767);
nor U4812 (N_4812,N_4715,N_4773);
xnor U4813 (N_4813,N_4755,N_4781);
and U4814 (N_4814,N_4719,N_4731);
nand U4815 (N_4815,N_4739,N_4768);
nand U4816 (N_4816,N_4734,N_4735);
nor U4817 (N_4817,N_4736,N_4775);
and U4818 (N_4818,N_4720,N_4716);
nor U4819 (N_4819,N_4774,N_4771);
and U4820 (N_4820,N_4758,N_4732);
and U4821 (N_4821,N_4733,N_4712);
xor U4822 (N_4822,N_4766,N_4763);
nor U4823 (N_4823,N_4759,N_4700);
xor U4824 (N_4824,N_4725,N_4782);
nor U4825 (N_4825,N_4765,N_4709);
or U4826 (N_4826,N_4794,N_4714);
and U4827 (N_4827,N_4747,N_4740);
or U4828 (N_4828,N_4701,N_4705);
nand U4829 (N_4829,N_4723,N_4798);
nor U4830 (N_4830,N_4770,N_4711);
xnor U4831 (N_4831,N_4790,N_4787);
nor U4832 (N_4832,N_4791,N_4729);
nand U4833 (N_4833,N_4779,N_4757);
or U4834 (N_4834,N_4762,N_4737);
nand U4835 (N_4835,N_4778,N_4751);
and U4836 (N_4836,N_4756,N_4764);
nor U4837 (N_4837,N_4738,N_4750);
or U4838 (N_4838,N_4703,N_4786);
or U4839 (N_4839,N_4795,N_4706);
nor U4840 (N_4840,N_4772,N_4797);
nor U4841 (N_4841,N_4753,N_4704);
nand U4842 (N_4842,N_4793,N_4784);
nor U4843 (N_4843,N_4730,N_4769);
nand U4844 (N_4844,N_4748,N_4783);
nand U4845 (N_4845,N_4754,N_4717);
nand U4846 (N_4846,N_4760,N_4744);
nand U4847 (N_4847,N_4789,N_4722);
or U4848 (N_4848,N_4749,N_4727);
xnor U4849 (N_4849,N_4785,N_4726);
xnor U4850 (N_4850,N_4762,N_4798);
xor U4851 (N_4851,N_4708,N_4720);
or U4852 (N_4852,N_4729,N_4774);
and U4853 (N_4853,N_4703,N_4702);
or U4854 (N_4854,N_4786,N_4705);
nor U4855 (N_4855,N_4709,N_4730);
and U4856 (N_4856,N_4770,N_4704);
nor U4857 (N_4857,N_4703,N_4745);
nor U4858 (N_4858,N_4722,N_4760);
nor U4859 (N_4859,N_4792,N_4710);
or U4860 (N_4860,N_4746,N_4767);
or U4861 (N_4861,N_4789,N_4716);
xnor U4862 (N_4862,N_4748,N_4773);
nand U4863 (N_4863,N_4796,N_4718);
xnor U4864 (N_4864,N_4729,N_4780);
xnor U4865 (N_4865,N_4727,N_4734);
nor U4866 (N_4866,N_4707,N_4791);
and U4867 (N_4867,N_4778,N_4734);
and U4868 (N_4868,N_4722,N_4798);
nor U4869 (N_4869,N_4792,N_4704);
nand U4870 (N_4870,N_4768,N_4721);
and U4871 (N_4871,N_4706,N_4740);
nor U4872 (N_4872,N_4770,N_4755);
xnor U4873 (N_4873,N_4787,N_4757);
nand U4874 (N_4874,N_4753,N_4756);
nand U4875 (N_4875,N_4794,N_4735);
and U4876 (N_4876,N_4755,N_4771);
or U4877 (N_4877,N_4733,N_4761);
and U4878 (N_4878,N_4712,N_4718);
nor U4879 (N_4879,N_4707,N_4738);
xnor U4880 (N_4880,N_4748,N_4720);
nor U4881 (N_4881,N_4775,N_4754);
and U4882 (N_4882,N_4709,N_4774);
and U4883 (N_4883,N_4707,N_4778);
xor U4884 (N_4884,N_4785,N_4792);
xnor U4885 (N_4885,N_4795,N_4769);
nand U4886 (N_4886,N_4790,N_4732);
xnor U4887 (N_4887,N_4702,N_4757);
and U4888 (N_4888,N_4721,N_4723);
and U4889 (N_4889,N_4742,N_4714);
nand U4890 (N_4890,N_4711,N_4752);
nor U4891 (N_4891,N_4776,N_4761);
nor U4892 (N_4892,N_4710,N_4786);
or U4893 (N_4893,N_4703,N_4706);
nand U4894 (N_4894,N_4786,N_4757);
and U4895 (N_4895,N_4762,N_4760);
xor U4896 (N_4896,N_4734,N_4707);
xnor U4897 (N_4897,N_4758,N_4781);
and U4898 (N_4898,N_4760,N_4765);
or U4899 (N_4899,N_4795,N_4782);
and U4900 (N_4900,N_4838,N_4844);
nand U4901 (N_4901,N_4864,N_4882);
nor U4902 (N_4902,N_4813,N_4860);
nand U4903 (N_4903,N_4862,N_4800);
or U4904 (N_4904,N_4847,N_4898);
nor U4905 (N_4905,N_4894,N_4897);
nand U4906 (N_4906,N_4845,N_4835);
nand U4907 (N_4907,N_4837,N_4805);
or U4908 (N_4908,N_4809,N_4856);
nor U4909 (N_4909,N_4804,N_4827);
and U4910 (N_4910,N_4821,N_4831);
nand U4911 (N_4911,N_4895,N_4857);
nand U4912 (N_4912,N_4874,N_4842);
xor U4913 (N_4913,N_4872,N_4888);
nor U4914 (N_4914,N_4843,N_4848);
xor U4915 (N_4915,N_4893,N_4803);
nand U4916 (N_4916,N_4855,N_4852);
nor U4917 (N_4917,N_4812,N_4858);
or U4918 (N_4918,N_4802,N_4829);
or U4919 (N_4919,N_4836,N_4885);
and U4920 (N_4920,N_4859,N_4818);
or U4921 (N_4921,N_4815,N_4899);
nand U4922 (N_4922,N_4816,N_4849);
and U4923 (N_4923,N_4820,N_4896);
xor U4924 (N_4924,N_4854,N_4887);
xnor U4925 (N_4925,N_4871,N_4890);
nor U4926 (N_4926,N_4825,N_4850);
xor U4927 (N_4927,N_4884,N_4830);
nand U4928 (N_4928,N_4808,N_4870);
nor U4929 (N_4929,N_4891,N_4878);
xnor U4930 (N_4930,N_4863,N_4834);
xnor U4931 (N_4931,N_4806,N_4873);
and U4932 (N_4932,N_4881,N_4832);
xnor U4933 (N_4933,N_4875,N_4892);
and U4934 (N_4934,N_4846,N_4853);
xnor U4935 (N_4935,N_4861,N_4833);
xnor U4936 (N_4936,N_4851,N_4819);
xor U4937 (N_4937,N_4839,N_4801);
xnor U4938 (N_4938,N_4868,N_4889);
or U4939 (N_4939,N_4886,N_4869);
and U4940 (N_4940,N_4807,N_4883);
xnor U4941 (N_4941,N_4817,N_4877);
and U4942 (N_4942,N_4840,N_4814);
and U4943 (N_4943,N_4810,N_4876);
or U4944 (N_4944,N_4828,N_4879);
nor U4945 (N_4945,N_4822,N_4867);
nor U4946 (N_4946,N_4823,N_4865);
or U4947 (N_4947,N_4811,N_4824);
xnor U4948 (N_4948,N_4866,N_4880);
and U4949 (N_4949,N_4841,N_4826);
xor U4950 (N_4950,N_4878,N_4863);
nor U4951 (N_4951,N_4807,N_4839);
nor U4952 (N_4952,N_4867,N_4811);
xnor U4953 (N_4953,N_4882,N_4857);
and U4954 (N_4954,N_4824,N_4849);
or U4955 (N_4955,N_4895,N_4843);
xor U4956 (N_4956,N_4887,N_4835);
nand U4957 (N_4957,N_4877,N_4830);
xnor U4958 (N_4958,N_4807,N_4891);
xor U4959 (N_4959,N_4805,N_4858);
xor U4960 (N_4960,N_4886,N_4851);
or U4961 (N_4961,N_4880,N_4807);
and U4962 (N_4962,N_4817,N_4808);
xor U4963 (N_4963,N_4877,N_4893);
xnor U4964 (N_4964,N_4844,N_4858);
nand U4965 (N_4965,N_4851,N_4840);
xor U4966 (N_4966,N_4826,N_4878);
nand U4967 (N_4967,N_4807,N_4836);
xor U4968 (N_4968,N_4843,N_4855);
nor U4969 (N_4969,N_4820,N_4848);
nand U4970 (N_4970,N_4892,N_4823);
and U4971 (N_4971,N_4827,N_4872);
nand U4972 (N_4972,N_4842,N_4836);
or U4973 (N_4973,N_4814,N_4826);
nor U4974 (N_4974,N_4840,N_4807);
nor U4975 (N_4975,N_4889,N_4894);
xnor U4976 (N_4976,N_4856,N_4814);
and U4977 (N_4977,N_4831,N_4818);
nor U4978 (N_4978,N_4832,N_4894);
and U4979 (N_4979,N_4879,N_4869);
nor U4980 (N_4980,N_4875,N_4898);
nand U4981 (N_4981,N_4859,N_4806);
or U4982 (N_4982,N_4809,N_4804);
xnor U4983 (N_4983,N_4823,N_4880);
nand U4984 (N_4984,N_4827,N_4801);
or U4985 (N_4985,N_4861,N_4841);
xor U4986 (N_4986,N_4816,N_4856);
and U4987 (N_4987,N_4881,N_4857);
xor U4988 (N_4988,N_4818,N_4852);
nor U4989 (N_4989,N_4882,N_4813);
and U4990 (N_4990,N_4825,N_4893);
xor U4991 (N_4991,N_4818,N_4864);
xnor U4992 (N_4992,N_4849,N_4894);
xnor U4993 (N_4993,N_4892,N_4869);
xor U4994 (N_4994,N_4867,N_4865);
or U4995 (N_4995,N_4801,N_4855);
xnor U4996 (N_4996,N_4847,N_4879);
and U4997 (N_4997,N_4847,N_4885);
xor U4998 (N_4998,N_4809,N_4859);
xor U4999 (N_4999,N_4878,N_4836);
xor U5000 (N_5000,N_4991,N_4903);
or U5001 (N_5001,N_4922,N_4921);
xnor U5002 (N_5002,N_4917,N_4976);
nand U5003 (N_5003,N_4910,N_4999);
xnor U5004 (N_5004,N_4931,N_4914);
nor U5005 (N_5005,N_4953,N_4995);
and U5006 (N_5006,N_4924,N_4935);
xnor U5007 (N_5007,N_4959,N_4938);
and U5008 (N_5008,N_4909,N_4988);
nor U5009 (N_5009,N_4945,N_4973);
and U5010 (N_5010,N_4925,N_4955);
and U5011 (N_5011,N_4962,N_4975);
and U5012 (N_5012,N_4947,N_4929);
or U5013 (N_5013,N_4989,N_4930);
xnor U5014 (N_5014,N_4919,N_4985);
or U5015 (N_5015,N_4993,N_4958);
nor U5016 (N_5016,N_4978,N_4932);
xnor U5017 (N_5017,N_4904,N_4972);
or U5018 (N_5018,N_4934,N_4926);
and U5019 (N_5019,N_4918,N_4977);
nand U5020 (N_5020,N_4979,N_4967);
xnor U5021 (N_5021,N_4900,N_4960);
xnor U5022 (N_5022,N_4939,N_4969);
nand U5023 (N_5023,N_4949,N_4964);
or U5024 (N_5024,N_4948,N_4987);
and U5025 (N_5025,N_4946,N_4956);
or U5026 (N_5026,N_4986,N_4998);
nor U5027 (N_5027,N_4923,N_4937);
xnor U5028 (N_5028,N_4920,N_4957);
or U5029 (N_5029,N_4982,N_4952);
or U5030 (N_5030,N_4950,N_4970);
or U5031 (N_5031,N_4983,N_4974);
nand U5032 (N_5032,N_4981,N_4965);
nor U5033 (N_5033,N_4944,N_4936);
xor U5034 (N_5034,N_4966,N_4912);
xor U5035 (N_5035,N_4905,N_4941);
nand U5036 (N_5036,N_4927,N_4901);
nand U5037 (N_5037,N_4968,N_4928);
nand U5038 (N_5038,N_4990,N_4961);
nor U5039 (N_5039,N_4907,N_4954);
nand U5040 (N_5040,N_4913,N_4984);
and U5041 (N_5041,N_4943,N_4933);
nand U5042 (N_5042,N_4942,N_4906);
nor U5043 (N_5043,N_4911,N_4994);
or U5044 (N_5044,N_4915,N_4997);
nor U5045 (N_5045,N_4992,N_4963);
or U5046 (N_5046,N_4980,N_4902);
nor U5047 (N_5047,N_4996,N_4971);
and U5048 (N_5048,N_4951,N_4908);
xor U5049 (N_5049,N_4916,N_4940);
or U5050 (N_5050,N_4961,N_4993);
nand U5051 (N_5051,N_4983,N_4904);
nand U5052 (N_5052,N_4978,N_4977);
nor U5053 (N_5053,N_4929,N_4969);
xnor U5054 (N_5054,N_4958,N_4900);
or U5055 (N_5055,N_4945,N_4905);
and U5056 (N_5056,N_4917,N_4994);
xor U5057 (N_5057,N_4961,N_4934);
nor U5058 (N_5058,N_4955,N_4902);
and U5059 (N_5059,N_4983,N_4959);
nor U5060 (N_5060,N_4996,N_4915);
and U5061 (N_5061,N_4995,N_4976);
nand U5062 (N_5062,N_4940,N_4914);
nor U5063 (N_5063,N_4980,N_4932);
or U5064 (N_5064,N_4982,N_4979);
and U5065 (N_5065,N_4913,N_4935);
and U5066 (N_5066,N_4909,N_4998);
and U5067 (N_5067,N_4956,N_4967);
nor U5068 (N_5068,N_4939,N_4940);
and U5069 (N_5069,N_4940,N_4951);
nand U5070 (N_5070,N_4973,N_4923);
or U5071 (N_5071,N_4999,N_4946);
and U5072 (N_5072,N_4916,N_4963);
nor U5073 (N_5073,N_4977,N_4994);
and U5074 (N_5074,N_4982,N_4976);
nor U5075 (N_5075,N_4913,N_4972);
and U5076 (N_5076,N_4921,N_4983);
nand U5077 (N_5077,N_4977,N_4983);
or U5078 (N_5078,N_4974,N_4969);
xnor U5079 (N_5079,N_4952,N_4979);
nand U5080 (N_5080,N_4998,N_4938);
nand U5081 (N_5081,N_4918,N_4941);
and U5082 (N_5082,N_4932,N_4925);
nand U5083 (N_5083,N_4936,N_4965);
and U5084 (N_5084,N_4950,N_4961);
nor U5085 (N_5085,N_4995,N_4947);
nor U5086 (N_5086,N_4900,N_4945);
nor U5087 (N_5087,N_4992,N_4916);
xnor U5088 (N_5088,N_4966,N_4926);
or U5089 (N_5089,N_4977,N_4906);
nand U5090 (N_5090,N_4958,N_4985);
xor U5091 (N_5091,N_4981,N_4954);
or U5092 (N_5092,N_4905,N_4926);
and U5093 (N_5093,N_4927,N_4975);
xnor U5094 (N_5094,N_4906,N_4929);
nor U5095 (N_5095,N_4931,N_4966);
or U5096 (N_5096,N_4910,N_4998);
or U5097 (N_5097,N_4937,N_4936);
or U5098 (N_5098,N_4968,N_4972);
xor U5099 (N_5099,N_4928,N_4983);
nor U5100 (N_5100,N_5089,N_5016);
xor U5101 (N_5101,N_5045,N_5011);
xor U5102 (N_5102,N_5041,N_5090);
xor U5103 (N_5103,N_5092,N_5023);
and U5104 (N_5104,N_5043,N_5013);
and U5105 (N_5105,N_5010,N_5046);
and U5106 (N_5106,N_5018,N_5082);
xnor U5107 (N_5107,N_5039,N_5002);
xnor U5108 (N_5108,N_5070,N_5052);
nand U5109 (N_5109,N_5063,N_5027);
or U5110 (N_5110,N_5049,N_5038);
nand U5111 (N_5111,N_5095,N_5005);
or U5112 (N_5112,N_5044,N_5079);
xnor U5113 (N_5113,N_5054,N_5067);
or U5114 (N_5114,N_5040,N_5029);
or U5115 (N_5115,N_5077,N_5057);
nor U5116 (N_5116,N_5053,N_5000);
and U5117 (N_5117,N_5083,N_5026);
and U5118 (N_5118,N_5091,N_5012);
or U5119 (N_5119,N_5071,N_5007);
nand U5120 (N_5120,N_5025,N_5003);
or U5121 (N_5121,N_5030,N_5042);
and U5122 (N_5122,N_5058,N_5080);
xnor U5123 (N_5123,N_5055,N_5084);
xnor U5124 (N_5124,N_5078,N_5035);
and U5125 (N_5125,N_5009,N_5097);
or U5126 (N_5126,N_5015,N_5096);
nand U5127 (N_5127,N_5085,N_5069);
or U5128 (N_5128,N_5059,N_5098);
or U5129 (N_5129,N_5047,N_5064);
nor U5130 (N_5130,N_5062,N_5036);
and U5131 (N_5131,N_5094,N_5008);
nor U5132 (N_5132,N_5004,N_5006);
or U5133 (N_5133,N_5031,N_5019);
nor U5134 (N_5134,N_5024,N_5068);
nand U5135 (N_5135,N_5086,N_5066);
xnor U5136 (N_5136,N_5072,N_5074);
xor U5137 (N_5137,N_5014,N_5028);
nor U5138 (N_5138,N_5032,N_5088);
xor U5139 (N_5139,N_5022,N_5034);
nand U5140 (N_5140,N_5065,N_5017);
or U5141 (N_5141,N_5073,N_5037);
or U5142 (N_5142,N_5076,N_5087);
nand U5143 (N_5143,N_5056,N_5001);
or U5144 (N_5144,N_5075,N_5099);
and U5145 (N_5145,N_5050,N_5033);
nor U5146 (N_5146,N_5020,N_5093);
and U5147 (N_5147,N_5021,N_5051);
and U5148 (N_5148,N_5048,N_5061);
or U5149 (N_5149,N_5060,N_5081);
nor U5150 (N_5150,N_5022,N_5027);
xor U5151 (N_5151,N_5025,N_5013);
and U5152 (N_5152,N_5091,N_5037);
and U5153 (N_5153,N_5096,N_5011);
nand U5154 (N_5154,N_5088,N_5028);
nor U5155 (N_5155,N_5035,N_5057);
or U5156 (N_5156,N_5007,N_5064);
or U5157 (N_5157,N_5043,N_5029);
xnor U5158 (N_5158,N_5089,N_5044);
nand U5159 (N_5159,N_5057,N_5069);
xor U5160 (N_5160,N_5058,N_5060);
nor U5161 (N_5161,N_5038,N_5029);
nand U5162 (N_5162,N_5022,N_5082);
or U5163 (N_5163,N_5067,N_5071);
nor U5164 (N_5164,N_5023,N_5078);
and U5165 (N_5165,N_5072,N_5096);
xor U5166 (N_5166,N_5086,N_5070);
or U5167 (N_5167,N_5031,N_5038);
nand U5168 (N_5168,N_5092,N_5060);
nand U5169 (N_5169,N_5036,N_5032);
nand U5170 (N_5170,N_5080,N_5003);
or U5171 (N_5171,N_5035,N_5008);
nor U5172 (N_5172,N_5078,N_5004);
xor U5173 (N_5173,N_5062,N_5086);
nand U5174 (N_5174,N_5099,N_5038);
nand U5175 (N_5175,N_5081,N_5000);
nand U5176 (N_5176,N_5027,N_5039);
xor U5177 (N_5177,N_5067,N_5081);
nor U5178 (N_5178,N_5010,N_5005);
xor U5179 (N_5179,N_5044,N_5005);
xor U5180 (N_5180,N_5093,N_5084);
and U5181 (N_5181,N_5091,N_5013);
or U5182 (N_5182,N_5026,N_5003);
and U5183 (N_5183,N_5019,N_5066);
xor U5184 (N_5184,N_5015,N_5017);
xor U5185 (N_5185,N_5022,N_5010);
nand U5186 (N_5186,N_5014,N_5006);
nor U5187 (N_5187,N_5058,N_5027);
and U5188 (N_5188,N_5016,N_5012);
or U5189 (N_5189,N_5068,N_5016);
and U5190 (N_5190,N_5044,N_5028);
xnor U5191 (N_5191,N_5000,N_5044);
xnor U5192 (N_5192,N_5030,N_5040);
nor U5193 (N_5193,N_5085,N_5086);
nand U5194 (N_5194,N_5066,N_5085);
xnor U5195 (N_5195,N_5053,N_5019);
or U5196 (N_5196,N_5003,N_5081);
nor U5197 (N_5197,N_5056,N_5089);
and U5198 (N_5198,N_5087,N_5007);
and U5199 (N_5199,N_5049,N_5085);
nand U5200 (N_5200,N_5171,N_5184);
nor U5201 (N_5201,N_5190,N_5110);
xnor U5202 (N_5202,N_5128,N_5175);
xnor U5203 (N_5203,N_5138,N_5122);
and U5204 (N_5204,N_5147,N_5141);
nor U5205 (N_5205,N_5105,N_5186);
xnor U5206 (N_5206,N_5130,N_5113);
xor U5207 (N_5207,N_5137,N_5121);
nand U5208 (N_5208,N_5132,N_5109);
xor U5209 (N_5209,N_5158,N_5145);
nand U5210 (N_5210,N_5111,N_5194);
and U5211 (N_5211,N_5102,N_5149);
and U5212 (N_5212,N_5173,N_5142);
xnor U5213 (N_5213,N_5148,N_5101);
or U5214 (N_5214,N_5153,N_5131);
nor U5215 (N_5215,N_5179,N_5104);
xor U5216 (N_5216,N_5151,N_5165);
nor U5217 (N_5217,N_5189,N_5191);
and U5218 (N_5218,N_5188,N_5117);
nor U5219 (N_5219,N_5119,N_5103);
nor U5220 (N_5220,N_5169,N_5164);
nor U5221 (N_5221,N_5181,N_5162);
or U5222 (N_5222,N_5167,N_5154);
nand U5223 (N_5223,N_5125,N_5168);
nand U5224 (N_5224,N_5197,N_5159);
nand U5225 (N_5225,N_5107,N_5116);
and U5226 (N_5226,N_5127,N_5118);
nand U5227 (N_5227,N_5106,N_5174);
and U5228 (N_5228,N_5198,N_5183);
and U5229 (N_5229,N_5156,N_5126);
nor U5230 (N_5230,N_5180,N_5114);
or U5231 (N_5231,N_5170,N_5143);
xnor U5232 (N_5232,N_5140,N_5166);
xnor U5233 (N_5233,N_5195,N_5112);
xor U5234 (N_5234,N_5152,N_5182);
nor U5235 (N_5235,N_5100,N_5124);
xor U5236 (N_5236,N_5146,N_5108);
nor U5237 (N_5237,N_5185,N_5120);
xnor U5238 (N_5238,N_5139,N_5172);
nand U5239 (N_5239,N_5196,N_5115);
xnor U5240 (N_5240,N_5161,N_5187);
nand U5241 (N_5241,N_5144,N_5133);
nor U5242 (N_5242,N_5193,N_5176);
and U5243 (N_5243,N_5178,N_5129);
xor U5244 (N_5244,N_5135,N_5136);
and U5245 (N_5245,N_5150,N_5192);
or U5246 (N_5246,N_5157,N_5160);
xor U5247 (N_5247,N_5123,N_5177);
nor U5248 (N_5248,N_5134,N_5163);
xnor U5249 (N_5249,N_5155,N_5199);
and U5250 (N_5250,N_5199,N_5167);
nand U5251 (N_5251,N_5174,N_5142);
and U5252 (N_5252,N_5198,N_5185);
or U5253 (N_5253,N_5154,N_5144);
nand U5254 (N_5254,N_5161,N_5169);
nand U5255 (N_5255,N_5199,N_5129);
or U5256 (N_5256,N_5155,N_5116);
xor U5257 (N_5257,N_5182,N_5116);
nand U5258 (N_5258,N_5111,N_5101);
xnor U5259 (N_5259,N_5144,N_5155);
nor U5260 (N_5260,N_5159,N_5150);
xor U5261 (N_5261,N_5106,N_5171);
and U5262 (N_5262,N_5137,N_5166);
nor U5263 (N_5263,N_5142,N_5170);
xnor U5264 (N_5264,N_5103,N_5136);
or U5265 (N_5265,N_5126,N_5135);
and U5266 (N_5266,N_5192,N_5121);
or U5267 (N_5267,N_5109,N_5168);
and U5268 (N_5268,N_5108,N_5110);
xnor U5269 (N_5269,N_5157,N_5167);
and U5270 (N_5270,N_5189,N_5103);
xor U5271 (N_5271,N_5123,N_5159);
xnor U5272 (N_5272,N_5122,N_5141);
nor U5273 (N_5273,N_5193,N_5124);
and U5274 (N_5274,N_5123,N_5164);
xnor U5275 (N_5275,N_5104,N_5188);
nor U5276 (N_5276,N_5111,N_5193);
and U5277 (N_5277,N_5176,N_5197);
nand U5278 (N_5278,N_5168,N_5188);
or U5279 (N_5279,N_5111,N_5155);
xnor U5280 (N_5280,N_5106,N_5127);
nor U5281 (N_5281,N_5124,N_5143);
and U5282 (N_5282,N_5181,N_5120);
or U5283 (N_5283,N_5105,N_5104);
nor U5284 (N_5284,N_5126,N_5191);
xor U5285 (N_5285,N_5155,N_5196);
xnor U5286 (N_5286,N_5158,N_5146);
nand U5287 (N_5287,N_5191,N_5146);
or U5288 (N_5288,N_5132,N_5110);
nand U5289 (N_5289,N_5140,N_5199);
nor U5290 (N_5290,N_5171,N_5140);
nand U5291 (N_5291,N_5161,N_5149);
nor U5292 (N_5292,N_5198,N_5108);
and U5293 (N_5293,N_5193,N_5165);
nor U5294 (N_5294,N_5135,N_5113);
nor U5295 (N_5295,N_5163,N_5131);
nor U5296 (N_5296,N_5133,N_5184);
or U5297 (N_5297,N_5117,N_5198);
nand U5298 (N_5298,N_5117,N_5164);
nor U5299 (N_5299,N_5173,N_5187);
xnor U5300 (N_5300,N_5266,N_5254);
or U5301 (N_5301,N_5232,N_5235);
or U5302 (N_5302,N_5230,N_5258);
xnor U5303 (N_5303,N_5221,N_5244);
and U5304 (N_5304,N_5212,N_5259);
and U5305 (N_5305,N_5285,N_5278);
or U5306 (N_5306,N_5224,N_5236);
nor U5307 (N_5307,N_5251,N_5246);
xnor U5308 (N_5308,N_5216,N_5283);
and U5309 (N_5309,N_5286,N_5296);
or U5310 (N_5310,N_5229,N_5217);
nor U5311 (N_5311,N_5215,N_5268);
xnor U5312 (N_5312,N_5276,N_5279);
nor U5313 (N_5313,N_5289,N_5218);
or U5314 (N_5314,N_5274,N_5281);
and U5315 (N_5315,N_5239,N_5257);
nor U5316 (N_5316,N_5242,N_5248);
or U5317 (N_5317,N_5204,N_5243);
nor U5318 (N_5318,N_5203,N_5249);
and U5319 (N_5319,N_5294,N_5264);
xor U5320 (N_5320,N_5270,N_5211);
and U5321 (N_5321,N_5299,N_5247);
or U5322 (N_5322,N_5226,N_5252);
nor U5323 (N_5323,N_5225,N_5222);
nand U5324 (N_5324,N_5260,N_5238);
nand U5325 (N_5325,N_5265,N_5262);
nand U5326 (N_5326,N_5223,N_5263);
and U5327 (N_5327,N_5273,N_5233);
and U5328 (N_5328,N_5220,N_5288);
nand U5329 (N_5329,N_5213,N_5206);
nor U5330 (N_5330,N_5253,N_5231);
or U5331 (N_5331,N_5201,N_5284);
xor U5332 (N_5332,N_5237,N_5292);
xor U5333 (N_5333,N_5291,N_5280);
and U5334 (N_5334,N_5256,N_5269);
xnor U5335 (N_5335,N_5295,N_5272);
and U5336 (N_5336,N_5234,N_5297);
or U5337 (N_5337,N_5227,N_5255);
nand U5338 (N_5338,N_5210,N_5200);
and U5339 (N_5339,N_5298,N_5241);
and U5340 (N_5340,N_5209,N_5207);
and U5341 (N_5341,N_5267,N_5214);
or U5342 (N_5342,N_5290,N_5282);
nand U5343 (N_5343,N_5293,N_5287);
or U5344 (N_5344,N_5275,N_5228);
xor U5345 (N_5345,N_5261,N_5277);
and U5346 (N_5346,N_5240,N_5219);
and U5347 (N_5347,N_5205,N_5250);
xor U5348 (N_5348,N_5271,N_5208);
or U5349 (N_5349,N_5202,N_5245);
nor U5350 (N_5350,N_5290,N_5285);
and U5351 (N_5351,N_5249,N_5235);
nor U5352 (N_5352,N_5228,N_5257);
and U5353 (N_5353,N_5214,N_5293);
xor U5354 (N_5354,N_5206,N_5239);
or U5355 (N_5355,N_5295,N_5286);
nor U5356 (N_5356,N_5200,N_5274);
nor U5357 (N_5357,N_5217,N_5291);
and U5358 (N_5358,N_5216,N_5295);
nor U5359 (N_5359,N_5239,N_5207);
nand U5360 (N_5360,N_5210,N_5203);
and U5361 (N_5361,N_5215,N_5238);
xnor U5362 (N_5362,N_5235,N_5283);
xor U5363 (N_5363,N_5256,N_5280);
nor U5364 (N_5364,N_5280,N_5216);
nor U5365 (N_5365,N_5271,N_5299);
nor U5366 (N_5366,N_5272,N_5218);
nand U5367 (N_5367,N_5239,N_5246);
nand U5368 (N_5368,N_5283,N_5212);
or U5369 (N_5369,N_5215,N_5205);
nand U5370 (N_5370,N_5279,N_5212);
nand U5371 (N_5371,N_5217,N_5214);
nor U5372 (N_5372,N_5227,N_5269);
and U5373 (N_5373,N_5265,N_5217);
or U5374 (N_5374,N_5246,N_5238);
nor U5375 (N_5375,N_5224,N_5294);
and U5376 (N_5376,N_5236,N_5291);
xor U5377 (N_5377,N_5227,N_5206);
or U5378 (N_5378,N_5214,N_5254);
nor U5379 (N_5379,N_5227,N_5273);
nand U5380 (N_5380,N_5270,N_5219);
nand U5381 (N_5381,N_5218,N_5204);
or U5382 (N_5382,N_5263,N_5228);
nor U5383 (N_5383,N_5224,N_5275);
nand U5384 (N_5384,N_5207,N_5241);
and U5385 (N_5385,N_5260,N_5242);
xor U5386 (N_5386,N_5210,N_5287);
and U5387 (N_5387,N_5293,N_5242);
nand U5388 (N_5388,N_5259,N_5222);
nand U5389 (N_5389,N_5258,N_5214);
nand U5390 (N_5390,N_5248,N_5258);
or U5391 (N_5391,N_5266,N_5298);
or U5392 (N_5392,N_5259,N_5203);
nand U5393 (N_5393,N_5249,N_5287);
or U5394 (N_5394,N_5269,N_5223);
nor U5395 (N_5395,N_5224,N_5254);
xor U5396 (N_5396,N_5253,N_5270);
nor U5397 (N_5397,N_5261,N_5299);
and U5398 (N_5398,N_5200,N_5230);
xnor U5399 (N_5399,N_5290,N_5241);
or U5400 (N_5400,N_5355,N_5395);
nor U5401 (N_5401,N_5347,N_5342);
and U5402 (N_5402,N_5374,N_5300);
nand U5403 (N_5403,N_5333,N_5392);
nor U5404 (N_5404,N_5306,N_5324);
and U5405 (N_5405,N_5383,N_5360);
or U5406 (N_5406,N_5315,N_5305);
nor U5407 (N_5407,N_5370,N_5369);
and U5408 (N_5408,N_5385,N_5398);
or U5409 (N_5409,N_5366,N_5314);
nand U5410 (N_5410,N_5323,N_5325);
xnor U5411 (N_5411,N_5361,N_5345);
nor U5412 (N_5412,N_5349,N_5350);
xor U5413 (N_5413,N_5382,N_5362);
nor U5414 (N_5414,N_5312,N_5304);
and U5415 (N_5415,N_5391,N_5353);
nor U5416 (N_5416,N_5338,N_5346);
nor U5417 (N_5417,N_5388,N_5301);
and U5418 (N_5418,N_5379,N_5341);
and U5419 (N_5419,N_5384,N_5386);
or U5420 (N_5420,N_5356,N_5329);
xor U5421 (N_5421,N_5327,N_5380);
nand U5422 (N_5422,N_5319,N_5352);
xnor U5423 (N_5423,N_5310,N_5351);
or U5424 (N_5424,N_5340,N_5344);
nand U5425 (N_5425,N_5317,N_5320);
xnor U5426 (N_5426,N_5322,N_5328);
and U5427 (N_5427,N_5394,N_5358);
nor U5428 (N_5428,N_5390,N_5376);
and U5429 (N_5429,N_5337,N_5316);
nor U5430 (N_5430,N_5359,N_5372);
nand U5431 (N_5431,N_5393,N_5368);
or U5432 (N_5432,N_5321,N_5309);
or U5433 (N_5433,N_5326,N_5330);
xnor U5434 (N_5434,N_5377,N_5364);
and U5435 (N_5435,N_5303,N_5302);
nand U5436 (N_5436,N_5335,N_5343);
xnor U5437 (N_5437,N_5331,N_5357);
nand U5438 (N_5438,N_5365,N_5373);
and U5439 (N_5439,N_5397,N_5332);
nand U5440 (N_5440,N_5371,N_5399);
nand U5441 (N_5441,N_5367,N_5311);
nand U5442 (N_5442,N_5375,N_5336);
nand U5443 (N_5443,N_5396,N_5313);
nand U5444 (N_5444,N_5307,N_5389);
nand U5445 (N_5445,N_5308,N_5387);
nor U5446 (N_5446,N_5339,N_5381);
or U5447 (N_5447,N_5354,N_5318);
and U5448 (N_5448,N_5363,N_5378);
nor U5449 (N_5449,N_5334,N_5348);
xnor U5450 (N_5450,N_5341,N_5375);
and U5451 (N_5451,N_5332,N_5330);
nand U5452 (N_5452,N_5314,N_5352);
nor U5453 (N_5453,N_5324,N_5357);
nor U5454 (N_5454,N_5321,N_5364);
nor U5455 (N_5455,N_5393,N_5373);
nand U5456 (N_5456,N_5394,N_5351);
or U5457 (N_5457,N_5315,N_5350);
xnor U5458 (N_5458,N_5377,N_5384);
nor U5459 (N_5459,N_5363,N_5379);
xor U5460 (N_5460,N_5301,N_5392);
nand U5461 (N_5461,N_5312,N_5394);
nand U5462 (N_5462,N_5325,N_5388);
xnor U5463 (N_5463,N_5389,N_5344);
or U5464 (N_5464,N_5387,N_5357);
nor U5465 (N_5465,N_5319,N_5311);
and U5466 (N_5466,N_5346,N_5320);
or U5467 (N_5467,N_5362,N_5307);
xor U5468 (N_5468,N_5307,N_5382);
and U5469 (N_5469,N_5397,N_5326);
and U5470 (N_5470,N_5350,N_5320);
nand U5471 (N_5471,N_5358,N_5363);
nand U5472 (N_5472,N_5354,N_5361);
nand U5473 (N_5473,N_5387,N_5390);
or U5474 (N_5474,N_5318,N_5370);
nor U5475 (N_5475,N_5363,N_5331);
and U5476 (N_5476,N_5344,N_5357);
nand U5477 (N_5477,N_5317,N_5365);
and U5478 (N_5478,N_5329,N_5304);
nand U5479 (N_5479,N_5308,N_5348);
nor U5480 (N_5480,N_5360,N_5357);
xor U5481 (N_5481,N_5368,N_5374);
nor U5482 (N_5482,N_5357,N_5389);
or U5483 (N_5483,N_5347,N_5379);
xor U5484 (N_5484,N_5317,N_5393);
nand U5485 (N_5485,N_5386,N_5358);
and U5486 (N_5486,N_5326,N_5375);
nor U5487 (N_5487,N_5340,N_5398);
xor U5488 (N_5488,N_5372,N_5369);
xor U5489 (N_5489,N_5304,N_5381);
nand U5490 (N_5490,N_5363,N_5341);
xnor U5491 (N_5491,N_5393,N_5376);
or U5492 (N_5492,N_5364,N_5333);
and U5493 (N_5493,N_5381,N_5370);
or U5494 (N_5494,N_5344,N_5341);
nand U5495 (N_5495,N_5357,N_5309);
nand U5496 (N_5496,N_5309,N_5326);
nand U5497 (N_5497,N_5396,N_5347);
nand U5498 (N_5498,N_5397,N_5301);
and U5499 (N_5499,N_5372,N_5322);
and U5500 (N_5500,N_5415,N_5449);
xnor U5501 (N_5501,N_5416,N_5440);
nand U5502 (N_5502,N_5492,N_5453);
and U5503 (N_5503,N_5470,N_5475);
or U5504 (N_5504,N_5457,N_5438);
nor U5505 (N_5505,N_5464,N_5456);
nor U5506 (N_5506,N_5497,N_5458);
nand U5507 (N_5507,N_5404,N_5444);
and U5508 (N_5508,N_5473,N_5491);
and U5509 (N_5509,N_5454,N_5448);
and U5510 (N_5510,N_5402,N_5485);
or U5511 (N_5511,N_5467,N_5437);
nor U5512 (N_5512,N_5496,N_5451);
nand U5513 (N_5513,N_5407,N_5487);
nor U5514 (N_5514,N_5498,N_5461);
and U5515 (N_5515,N_5429,N_5433);
nor U5516 (N_5516,N_5495,N_5455);
and U5517 (N_5517,N_5428,N_5476);
and U5518 (N_5518,N_5410,N_5431);
or U5519 (N_5519,N_5468,N_5452);
nand U5520 (N_5520,N_5427,N_5447);
nand U5521 (N_5521,N_5441,N_5401);
nand U5522 (N_5522,N_5414,N_5430);
nand U5523 (N_5523,N_5479,N_5423);
xor U5524 (N_5524,N_5499,N_5432);
nor U5525 (N_5525,N_5465,N_5488);
nor U5526 (N_5526,N_5445,N_5460);
xor U5527 (N_5527,N_5493,N_5434);
nor U5528 (N_5528,N_5443,N_5463);
or U5529 (N_5529,N_5450,N_5481);
xor U5530 (N_5530,N_5419,N_5486);
xor U5531 (N_5531,N_5409,N_5474);
nor U5532 (N_5532,N_5436,N_5459);
and U5533 (N_5533,N_5466,N_5490);
and U5534 (N_5534,N_5421,N_5417);
xor U5535 (N_5535,N_5469,N_5425);
or U5536 (N_5536,N_5439,N_5462);
or U5537 (N_5537,N_5413,N_5424);
xnor U5538 (N_5538,N_5406,N_5483);
and U5539 (N_5539,N_5484,N_5420);
nand U5540 (N_5540,N_5442,N_5403);
or U5541 (N_5541,N_5411,N_5477);
nor U5542 (N_5542,N_5435,N_5471);
and U5543 (N_5543,N_5482,N_5494);
nand U5544 (N_5544,N_5489,N_5400);
xor U5545 (N_5545,N_5418,N_5478);
nand U5546 (N_5546,N_5412,N_5422);
xnor U5547 (N_5547,N_5405,N_5408);
nand U5548 (N_5548,N_5472,N_5426);
nor U5549 (N_5549,N_5480,N_5446);
xor U5550 (N_5550,N_5409,N_5406);
xnor U5551 (N_5551,N_5405,N_5412);
nor U5552 (N_5552,N_5480,N_5408);
and U5553 (N_5553,N_5408,N_5427);
xor U5554 (N_5554,N_5499,N_5427);
nor U5555 (N_5555,N_5465,N_5454);
or U5556 (N_5556,N_5479,N_5487);
xor U5557 (N_5557,N_5445,N_5414);
nand U5558 (N_5558,N_5419,N_5404);
xnor U5559 (N_5559,N_5481,N_5420);
nand U5560 (N_5560,N_5449,N_5472);
or U5561 (N_5561,N_5497,N_5409);
or U5562 (N_5562,N_5433,N_5420);
nand U5563 (N_5563,N_5494,N_5479);
nor U5564 (N_5564,N_5427,N_5483);
or U5565 (N_5565,N_5423,N_5480);
xnor U5566 (N_5566,N_5430,N_5418);
and U5567 (N_5567,N_5490,N_5419);
or U5568 (N_5568,N_5471,N_5473);
nand U5569 (N_5569,N_5483,N_5481);
and U5570 (N_5570,N_5460,N_5482);
xor U5571 (N_5571,N_5401,N_5431);
or U5572 (N_5572,N_5410,N_5414);
nor U5573 (N_5573,N_5445,N_5452);
nand U5574 (N_5574,N_5415,N_5472);
nor U5575 (N_5575,N_5475,N_5441);
nor U5576 (N_5576,N_5402,N_5405);
nand U5577 (N_5577,N_5429,N_5443);
nand U5578 (N_5578,N_5484,N_5490);
and U5579 (N_5579,N_5416,N_5436);
xnor U5580 (N_5580,N_5498,N_5468);
nor U5581 (N_5581,N_5438,N_5477);
and U5582 (N_5582,N_5440,N_5432);
or U5583 (N_5583,N_5401,N_5495);
nand U5584 (N_5584,N_5462,N_5419);
or U5585 (N_5585,N_5493,N_5482);
or U5586 (N_5586,N_5428,N_5456);
nor U5587 (N_5587,N_5494,N_5415);
and U5588 (N_5588,N_5433,N_5470);
nand U5589 (N_5589,N_5430,N_5435);
nor U5590 (N_5590,N_5495,N_5445);
and U5591 (N_5591,N_5469,N_5468);
and U5592 (N_5592,N_5472,N_5402);
nand U5593 (N_5593,N_5423,N_5403);
xnor U5594 (N_5594,N_5496,N_5475);
xnor U5595 (N_5595,N_5471,N_5424);
or U5596 (N_5596,N_5484,N_5494);
xor U5597 (N_5597,N_5406,N_5476);
xnor U5598 (N_5598,N_5432,N_5481);
and U5599 (N_5599,N_5495,N_5457);
xor U5600 (N_5600,N_5528,N_5553);
nand U5601 (N_5601,N_5506,N_5526);
nor U5602 (N_5602,N_5519,N_5598);
nand U5603 (N_5603,N_5576,N_5539);
and U5604 (N_5604,N_5515,N_5579);
nand U5605 (N_5605,N_5572,N_5500);
nor U5606 (N_5606,N_5554,N_5585);
or U5607 (N_5607,N_5547,N_5516);
xor U5608 (N_5608,N_5563,N_5592);
or U5609 (N_5609,N_5545,N_5591);
and U5610 (N_5610,N_5502,N_5533);
xnor U5611 (N_5611,N_5548,N_5508);
nor U5612 (N_5612,N_5571,N_5577);
and U5613 (N_5613,N_5543,N_5514);
and U5614 (N_5614,N_5521,N_5595);
nand U5615 (N_5615,N_5504,N_5555);
nand U5616 (N_5616,N_5527,N_5549);
nand U5617 (N_5617,N_5501,N_5520);
xor U5618 (N_5618,N_5535,N_5558);
xor U5619 (N_5619,N_5540,N_5581);
xor U5620 (N_5620,N_5580,N_5525);
nor U5621 (N_5621,N_5560,N_5534);
or U5622 (N_5622,N_5578,N_5518);
nor U5623 (N_5623,N_5510,N_5513);
nor U5624 (N_5624,N_5582,N_5556);
xor U5625 (N_5625,N_5562,N_5568);
or U5626 (N_5626,N_5524,N_5590);
nand U5627 (N_5627,N_5541,N_5569);
nor U5628 (N_5628,N_5511,N_5536);
xor U5629 (N_5629,N_5588,N_5542);
nor U5630 (N_5630,N_5546,N_5584);
or U5631 (N_5631,N_5559,N_5538);
nand U5632 (N_5632,N_5551,N_5523);
xnor U5633 (N_5633,N_5550,N_5594);
xnor U5634 (N_5634,N_5509,N_5599);
and U5635 (N_5635,N_5532,N_5531);
or U5636 (N_5636,N_5574,N_5561);
nand U5637 (N_5637,N_5583,N_5589);
or U5638 (N_5638,N_5557,N_5596);
and U5639 (N_5639,N_5529,N_5587);
and U5640 (N_5640,N_5570,N_5522);
and U5641 (N_5641,N_5505,N_5597);
and U5642 (N_5642,N_5573,N_5512);
or U5643 (N_5643,N_5530,N_5517);
xor U5644 (N_5644,N_5503,N_5593);
or U5645 (N_5645,N_5567,N_5564);
nor U5646 (N_5646,N_5575,N_5507);
or U5647 (N_5647,N_5552,N_5565);
and U5648 (N_5648,N_5586,N_5566);
nor U5649 (N_5649,N_5544,N_5537);
and U5650 (N_5650,N_5589,N_5511);
nor U5651 (N_5651,N_5529,N_5514);
xnor U5652 (N_5652,N_5516,N_5511);
nor U5653 (N_5653,N_5538,N_5592);
nand U5654 (N_5654,N_5580,N_5565);
and U5655 (N_5655,N_5548,N_5578);
nor U5656 (N_5656,N_5503,N_5571);
xnor U5657 (N_5657,N_5540,N_5563);
nand U5658 (N_5658,N_5528,N_5541);
xnor U5659 (N_5659,N_5549,N_5529);
xor U5660 (N_5660,N_5555,N_5543);
xnor U5661 (N_5661,N_5544,N_5583);
or U5662 (N_5662,N_5504,N_5545);
nand U5663 (N_5663,N_5501,N_5548);
or U5664 (N_5664,N_5502,N_5543);
or U5665 (N_5665,N_5516,N_5523);
and U5666 (N_5666,N_5567,N_5576);
and U5667 (N_5667,N_5520,N_5516);
nand U5668 (N_5668,N_5575,N_5562);
nor U5669 (N_5669,N_5516,N_5510);
and U5670 (N_5670,N_5515,N_5537);
nand U5671 (N_5671,N_5506,N_5585);
and U5672 (N_5672,N_5501,N_5510);
xnor U5673 (N_5673,N_5592,N_5599);
xor U5674 (N_5674,N_5524,N_5592);
nand U5675 (N_5675,N_5513,N_5595);
nor U5676 (N_5676,N_5509,N_5594);
nor U5677 (N_5677,N_5559,N_5512);
nor U5678 (N_5678,N_5510,N_5571);
nand U5679 (N_5679,N_5590,N_5596);
nor U5680 (N_5680,N_5535,N_5541);
nand U5681 (N_5681,N_5518,N_5572);
or U5682 (N_5682,N_5505,N_5555);
and U5683 (N_5683,N_5532,N_5542);
nand U5684 (N_5684,N_5552,N_5593);
or U5685 (N_5685,N_5527,N_5581);
xnor U5686 (N_5686,N_5564,N_5581);
or U5687 (N_5687,N_5599,N_5530);
nor U5688 (N_5688,N_5508,N_5562);
xnor U5689 (N_5689,N_5530,N_5597);
nor U5690 (N_5690,N_5597,N_5585);
xnor U5691 (N_5691,N_5563,N_5506);
nand U5692 (N_5692,N_5531,N_5577);
xor U5693 (N_5693,N_5587,N_5531);
xnor U5694 (N_5694,N_5553,N_5509);
xnor U5695 (N_5695,N_5546,N_5542);
nor U5696 (N_5696,N_5556,N_5522);
xor U5697 (N_5697,N_5536,N_5505);
xnor U5698 (N_5698,N_5576,N_5521);
or U5699 (N_5699,N_5531,N_5525);
nand U5700 (N_5700,N_5631,N_5654);
and U5701 (N_5701,N_5648,N_5665);
and U5702 (N_5702,N_5640,N_5687);
nor U5703 (N_5703,N_5608,N_5616);
or U5704 (N_5704,N_5697,N_5638);
or U5705 (N_5705,N_5604,N_5698);
nand U5706 (N_5706,N_5689,N_5642);
nand U5707 (N_5707,N_5683,N_5680);
or U5708 (N_5708,N_5669,N_5603);
xnor U5709 (N_5709,N_5660,N_5601);
xnor U5710 (N_5710,N_5613,N_5637);
xor U5711 (N_5711,N_5627,N_5668);
xnor U5712 (N_5712,N_5691,N_5670);
nand U5713 (N_5713,N_5686,N_5624);
nand U5714 (N_5714,N_5647,N_5611);
or U5715 (N_5715,N_5646,N_5652);
nor U5716 (N_5716,N_5690,N_5623);
and U5717 (N_5717,N_5664,N_5674);
and U5718 (N_5718,N_5612,N_5633);
nand U5719 (N_5719,N_5658,N_5681);
nand U5720 (N_5720,N_5606,N_5653);
or U5721 (N_5721,N_5610,N_5671);
nand U5722 (N_5722,N_5656,N_5626);
xnor U5723 (N_5723,N_5661,N_5639);
xor U5724 (N_5724,N_5684,N_5672);
nor U5725 (N_5725,N_5659,N_5645);
and U5726 (N_5726,N_5618,N_5625);
xor U5727 (N_5727,N_5657,N_5676);
nor U5728 (N_5728,N_5615,N_5644);
or U5729 (N_5729,N_5692,N_5609);
xnor U5730 (N_5730,N_5650,N_5602);
or U5731 (N_5731,N_5628,N_5649);
or U5732 (N_5732,N_5677,N_5643);
nand U5733 (N_5733,N_5600,N_5634);
xor U5734 (N_5734,N_5630,N_5675);
or U5735 (N_5735,N_5666,N_5685);
nor U5736 (N_5736,N_5622,N_5632);
nor U5737 (N_5737,N_5635,N_5629);
nor U5738 (N_5738,N_5655,N_5651);
and U5739 (N_5739,N_5682,N_5673);
and U5740 (N_5740,N_5621,N_5678);
nand U5741 (N_5741,N_5641,N_5694);
xnor U5742 (N_5742,N_5620,N_5679);
and U5743 (N_5743,N_5662,N_5607);
or U5744 (N_5744,N_5667,N_5663);
or U5745 (N_5745,N_5617,N_5614);
nor U5746 (N_5746,N_5695,N_5699);
nor U5747 (N_5747,N_5619,N_5693);
or U5748 (N_5748,N_5688,N_5605);
nand U5749 (N_5749,N_5696,N_5636);
nor U5750 (N_5750,N_5690,N_5694);
nor U5751 (N_5751,N_5658,N_5618);
xnor U5752 (N_5752,N_5672,N_5608);
nand U5753 (N_5753,N_5606,N_5603);
and U5754 (N_5754,N_5602,N_5672);
xor U5755 (N_5755,N_5640,N_5685);
nand U5756 (N_5756,N_5614,N_5622);
nand U5757 (N_5757,N_5621,N_5647);
and U5758 (N_5758,N_5665,N_5673);
and U5759 (N_5759,N_5636,N_5690);
and U5760 (N_5760,N_5673,N_5679);
nand U5761 (N_5761,N_5653,N_5645);
nor U5762 (N_5762,N_5640,N_5613);
or U5763 (N_5763,N_5610,N_5638);
nand U5764 (N_5764,N_5645,N_5691);
nor U5765 (N_5765,N_5649,N_5616);
xnor U5766 (N_5766,N_5698,N_5681);
nand U5767 (N_5767,N_5682,N_5680);
or U5768 (N_5768,N_5697,N_5657);
xnor U5769 (N_5769,N_5605,N_5616);
nor U5770 (N_5770,N_5636,N_5609);
or U5771 (N_5771,N_5614,N_5661);
and U5772 (N_5772,N_5619,N_5661);
and U5773 (N_5773,N_5697,N_5679);
and U5774 (N_5774,N_5657,N_5693);
xor U5775 (N_5775,N_5616,N_5662);
or U5776 (N_5776,N_5654,N_5658);
or U5777 (N_5777,N_5665,N_5696);
xnor U5778 (N_5778,N_5635,N_5666);
nor U5779 (N_5779,N_5640,N_5641);
nor U5780 (N_5780,N_5611,N_5615);
nand U5781 (N_5781,N_5649,N_5627);
nor U5782 (N_5782,N_5695,N_5654);
nor U5783 (N_5783,N_5603,N_5605);
nand U5784 (N_5784,N_5679,N_5642);
or U5785 (N_5785,N_5675,N_5685);
and U5786 (N_5786,N_5662,N_5668);
nand U5787 (N_5787,N_5633,N_5656);
xnor U5788 (N_5788,N_5614,N_5697);
nor U5789 (N_5789,N_5646,N_5686);
and U5790 (N_5790,N_5680,N_5618);
nand U5791 (N_5791,N_5689,N_5698);
nor U5792 (N_5792,N_5684,N_5651);
nand U5793 (N_5793,N_5687,N_5604);
xor U5794 (N_5794,N_5686,N_5652);
nand U5795 (N_5795,N_5640,N_5614);
and U5796 (N_5796,N_5611,N_5624);
and U5797 (N_5797,N_5689,N_5658);
nor U5798 (N_5798,N_5618,N_5631);
or U5799 (N_5799,N_5656,N_5655);
nor U5800 (N_5800,N_5712,N_5744);
nor U5801 (N_5801,N_5741,N_5732);
and U5802 (N_5802,N_5725,N_5792);
nand U5803 (N_5803,N_5774,N_5770);
nand U5804 (N_5804,N_5747,N_5786);
nand U5805 (N_5805,N_5748,N_5745);
nand U5806 (N_5806,N_5709,N_5779);
nor U5807 (N_5807,N_5739,N_5737);
or U5808 (N_5808,N_5705,N_5798);
nor U5809 (N_5809,N_5775,N_5730);
and U5810 (N_5810,N_5754,N_5704);
nor U5811 (N_5811,N_5794,N_5715);
and U5812 (N_5812,N_5752,N_5778);
xnor U5813 (N_5813,N_5766,N_5700);
nor U5814 (N_5814,N_5764,N_5729);
nor U5815 (N_5815,N_5762,N_5784);
xor U5816 (N_5816,N_5783,N_5789);
and U5817 (N_5817,N_5785,N_5795);
nand U5818 (N_5818,N_5793,N_5791);
xnor U5819 (N_5819,N_5788,N_5753);
or U5820 (N_5820,N_5735,N_5726);
and U5821 (N_5821,N_5782,N_5714);
nand U5822 (N_5822,N_5799,N_5767);
nand U5823 (N_5823,N_5727,N_5746);
and U5824 (N_5824,N_5731,N_5743);
xor U5825 (N_5825,N_5713,N_5742);
or U5826 (N_5826,N_5710,N_5734);
or U5827 (N_5827,N_5755,N_5711);
nor U5828 (N_5828,N_5757,N_5776);
nor U5829 (N_5829,N_5708,N_5736);
xor U5830 (N_5830,N_5772,N_5733);
or U5831 (N_5831,N_5750,N_5756);
xnor U5832 (N_5832,N_5781,N_5777);
nor U5833 (N_5833,N_5706,N_5724);
nor U5834 (N_5834,N_5761,N_5768);
or U5835 (N_5835,N_5787,N_5719);
xnor U5836 (N_5836,N_5716,N_5749);
and U5837 (N_5837,N_5723,N_5717);
and U5838 (N_5838,N_5797,N_5703);
and U5839 (N_5839,N_5701,N_5773);
nand U5840 (N_5840,N_5769,N_5751);
xor U5841 (N_5841,N_5738,N_5728);
and U5842 (N_5842,N_5718,N_5722);
or U5843 (N_5843,N_5707,N_5771);
or U5844 (N_5844,N_5780,N_5720);
nand U5845 (N_5845,N_5760,N_5790);
nand U5846 (N_5846,N_5796,N_5759);
xor U5847 (N_5847,N_5740,N_5765);
nand U5848 (N_5848,N_5763,N_5758);
and U5849 (N_5849,N_5721,N_5702);
and U5850 (N_5850,N_5782,N_5717);
or U5851 (N_5851,N_5715,N_5728);
and U5852 (N_5852,N_5737,N_5748);
or U5853 (N_5853,N_5747,N_5776);
nand U5854 (N_5854,N_5743,N_5768);
and U5855 (N_5855,N_5762,N_5782);
and U5856 (N_5856,N_5786,N_5726);
xnor U5857 (N_5857,N_5752,N_5798);
nand U5858 (N_5858,N_5745,N_5718);
and U5859 (N_5859,N_5799,N_5748);
nor U5860 (N_5860,N_5753,N_5706);
or U5861 (N_5861,N_5739,N_5781);
and U5862 (N_5862,N_5722,N_5713);
nand U5863 (N_5863,N_5799,N_5792);
or U5864 (N_5864,N_5726,N_5729);
nand U5865 (N_5865,N_5788,N_5718);
xnor U5866 (N_5866,N_5754,N_5736);
nor U5867 (N_5867,N_5767,N_5717);
nor U5868 (N_5868,N_5777,N_5720);
nand U5869 (N_5869,N_5778,N_5731);
nor U5870 (N_5870,N_5794,N_5798);
nor U5871 (N_5871,N_5713,N_5778);
and U5872 (N_5872,N_5753,N_5776);
and U5873 (N_5873,N_5742,N_5779);
nand U5874 (N_5874,N_5700,N_5707);
and U5875 (N_5875,N_5777,N_5791);
and U5876 (N_5876,N_5728,N_5791);
nor U5877 (N_5877,N_5726,N_5711);
nor U5878 (N_5878,N_5738,N_5735);
nor U5879 (N_5879,N_5701,N_5724);
or U5880 (N_5880,N_5783,N_5712);
nor U5881 (N_5881,N_5766,N_5736);
nor U5882 (N_5882,N_5759,N_5719);
nor U5883 (N_5883,N_5736,N_5730);
xnor U5884 (N_5884,N_5761,N_5755);
nand U5885 (N_5885,N_5779,N_5757);
nor U5886 (N_5886,N_5733,N_5758);
nand U5887 (N_5887,N_5709,N_5772);
or U5888 (N_5888,N_5757,N_5777);
nand U5889 (N_5889,N_5769,N_5712);
or U5890 (N_5890,N_5710,N_5769);
or U5891 (N_5891,N_5767,N_5798);
or U5892 (N_5892,N_5787,N_5721);
and U5893 (N_5893,N_5717,N_5752);
xnor U5894 (N_5894,N_5715,N_5724);
xor U5895 (N_5895,N_5772,N_5735);
nand U5896 (N_5896,N_5783,N_5715);
xor U5897 (N_5897,N_5794,N_5734);
xnor U5898 (N_5898,N_5761,N_5758);
xnor U5899 (N_5899,N_5791,N_5731);
and U5900 (N_5900,N_5897,N_5803);
or U5901 (N_5901,N_5896,N_5879);
nor U5902 (N_5902,N_5863,N_5886);
nand U5903 (N_5903,N_5836,N_5817);
and U5904 (N_5904,N_5864,N_5839);
and U5905 (N_5905,N_5831,N_5837);
and U5906 (N_5906,N_5812,N_5804);
or U5907 (N_5907,N_5846,N_5834);
and U5908 (N_5908,N_5881,N_5856);
xnor U5909 (N_5909,N_5830,N_5867);
and U5910 (N_5910,N_5811,N_5891);
nor U5911 (N_5911,N_5809,N_5857);
xor U5912 (N_5912,N_5825,N_5816);
nand U5913 (N_5913,N_5885,N_5823);
nand U5914 (N_5914,N_5875,N_5848);
xnor U5915 (N_5915,N_5873,N_5806);
and U5916 (N_5916,N_5843,N_5888);
or U5917 (N_5917,N_5835,N_5824);
nor U5918 (N_5918,N_5854,N_5847);
nor U5919 (N_5919,N_5820,N_5884);
nand U5920 (N_5920,N_5850,N_5871);
or U5921 (N_5921,N_5899,N_5865);
and U5922 (N_5922,N_5898,N_5853);
nor U5923 (N_5923,N_5890,N_5892);
xnor U5924 (N_5924,N_5874,N_5828);
and U5925 (N_5925,N_5819,N_5876);
or U5926 (N_5926,N_5813,N_5869);
nor U5927 (N_5927,N_5844,N_5895);
and U5928 (N_5928,N_5807,N_5838);
or U5929 (N_5929,N_5849,N_5887);
nand U5930 (N_5930,N_5829,N_5827);
nand U5931 (N_5931,N_5851,N_5859);
or U5932 (N_5932,N_5818,N_5832);
xnor U5933 (N_5933,N_5852,N_5808);
nand U5934 (N_5934,N_5815,N_5814);
xnor U5935 (N_5935,N_5810,N_5860);
nor U5936 (N_5936,N_5858,N_5841);
or U5937 (N_5937,N_5870,N_5868);
and U5938 (N_5938,N_5826,N_5889);
nand U5939 (N_5939,N_5883,N_5877);
and U5940 (N_5940,N_5880,N_5822);
and U5941 (N_5941,N_5893,N_5862);
nand U5942 (N_5942,N_5845,N_5855);
nand U5943 (N_5943,N_5878,N_5894);
nor U5944 (N_5944,N_5833,N_5801);
xor U5945 (N_5945,N_5872,N_5866);
nor U5946 (N_5946,N_5840,N_5800);
xnor U5947 (N_5947,N_5802,N_5842);
and U5948 (N_5948,N_5861,N_5882);
xnor U5949 (N_5949,N_5821,N_5805);
nand U5950 (N_5950,N_5873,N_5813);
nand U5951 (N_5951,N_5859,N_5871);
xor U5952 (N_5952,N_5840,N_5851);
nor U5953 (N_5953,N_5846,N_5848);
and U5954 (N_5954,N_5845,N_5840);
or U5955 (N_5955,N_5800,N_5848);
xnor U5956 (N_5956,N_5818,N_5876);
or U5957 (N_5957,N_5844,N_5815);
and U5958 (N_5958,N_5815,N_5810);
xnor U5959 (N_5959,N_5876,N_5827);
and U5960 (N_5960,N_5895,N_5856);
and U5961 (N_5961,N_5891,N_5831);
xor U5962 (N_5962,N_5883,N_5860);
or U5963 (N_5963,N_5866,N_5899);
or U5964 (N_5964,N_5863,N_5813);
or U5965 (N_5965,N_5850,N_5840);
and U5966 (N_5966,N_5864,N_5811);
or U5967 (N_5967,N_5839,N_5852);
xnor U5968 (N_5968,N_5840,N_5807);
nand U5969 (N_5969,N_5824,N_5896);
nor U5970 (N_5970,N_5842,N_5883);
and U5971 (N_5971,N_5815,N_5822);
or U5972 (N_5972,N_5890,N_5849);
xnor U5973 (N_5973,N_5805,N_5808);
or U5974 (N_5974,N_5870,N_5822);
nor U5975 (N_5975,N_5873,N_5893);
and U5976 (N_5976,N_5820,N_5861);
nand U5977 (N_5977,N_5809,N_5820);
and U5978 (N_5978,N_5822,N_5869);
xor U5979 (N_5979,N_5827,N_5808);
nor U5980 (N_5980,N_5861,N_5866);
and U5981 (N_5981,N_5801,N_5803);
nand U5982 (N_5982,N_5842,N_5854);
nor U5983 (N_5983,N_5815,N_5881);
nor U5984 (N_5984,N_5830,N_5827);
or U5985 (N_5985,N_5876,N_5885);
or U5986 (N_5986,N_5849,N_5865);
xor U5987 (N_5987,N_5817,N_5800);
and U5988 (N_5988,N_5824,N_5814);
nor U5989 (N_5989,N_5830,N_5865);
nand U5990 (N_5990,N_5827,N_5814);
nor U5991 (N_5991,N_5898,N_5863);
and U5992 (N_5992,N_5811,N_5889);
nor U5993 (N_5993,N_5889,N_5806);
and U5994 (N_5994,N_5877,N_5894);
xor U5995 (N_5995,N_5865,N_5898);
and U5996 (N_5996,N_5832,N_5800);
nor U5997 (N_5997,N_5836,N_5871);
nor U5998 (N_5998,N_5893,N_5817);
nor U5999 (N_5999,N_5876,N_5810);
and U6000 (N_6000,N_5948,N_5980);
nor U6001 (N_6001,N_5909,N_5957);
or U6002 (N_6002,N_5992,N_5907);
nand U6003 (N_6003,N_5950,N_5986);
and U6004 (N_6004,N_5922,N_5943);
nor U6005 (N_6005,N_5997,N_5955);
or U6006 (N_6006,N_5915,N_5998);
nand U6007 (N_6007,N_5938,N_5919);
xnor U6008 (N_6008,N_5987,N_5990);
nor U6009 (N_6009,N_5913,N_5927);
and U6010 (N_6010,N_5973,N_5903);
nor U6011 (N_6011,N_5952,N_5969);
nor U6012 (N_6012,N_5901,N_5984);
and U6013 (N_6013,N_5941,N_5974);
xor U6014 (N_6014,N_5908,N_5911);
and U6015 (N_6015,N_5976,N_5921);
and U6016 (N_6016,N_5964,N_5942);
xnor U6017 (N_6017,N_5925,N_5929);
and U6018 (N_6018,N_5972,N_5991);
nor U6019 (N_6019,N_5981,N_5928);
nand U6020 (N_6020,N_5989,N_5902);
nand U6021 (N_6021,N_5954,N_5958);
or U6022 (N_6022,N_5996,N_5906);
xnor U6023 (N_6023,N_5959,N_5914);
and U6024 (N_6024,N_5988,N_5904);
and U6025 (N_6025,N_5978,N_5905);
or U6026 (N_6026,N_5961,N_5960);
xnor U6027 (N_6027,N_5912,N_5993);
or U6028 (N_6028,N_5926,N_5946);
or U6029 (N_6029,N_5994,N_5931);
nand U6030 (N_6030,N_5971,N_5949);
nor U6031 (N_6031,N_5933,N_5916);
xnor U6032 (N_6032,N_5965,N_5900);
and U6033 (N_6033,N_5975,N_5985);
nor U6034 (N_6034,N_5999,N_5935);
nand U6035 (N_6035,N_5918,N_5970);
or U6036 (N_6036,N_5977,N_5940);
xor U6037 (N_6037,N_5956,N_5983);
or U6038 (N_6038,N_5924,N_5951);
nor U6039 (N_6039,N_5944,N_5953);
and U6040 (N_6040,N_5982,N_5966);
or U6041 (N_6041,N_5962,N_5968);
nor U6042 (N_6042,N_5923,N_5945);
xor U6043 (N_6043,N_5995,N_5934);
xor U6044 (N_6044,N_5939,N_5932);
nor U6045 (N_6045,N_5937,N_5979);
nor U6046 (N_6046,N_5963,N_5910);
nor U6047 (N_6047,N_5967,N_5936);
nand U6048 (N_6048,N_5920,N_5930);
or U6049 (N_6049,N_5947,N_5917);
nand U6050 (N_6050,N_5947,N_5926);
and U6051 (N_6051,N_5977,N_5988);
nor U6052 (N_6052,N_5972,N_5994);
nand U6053 (N_6053,N_5911,N_5998);
nor U6054 (N_6054,N_5961,N_5949);
and U6055 (N_6055,N_5910,N_5961);
and U6056 (N_6056,N_5952,N_5992);
or U6057 (N_6057,N_5916,N_5999);
nor U6058 (N_6058,N_5940,N_5915);
and U6059 (N_6059,N_5927,N_5906);
nor U6060 (N_6060,N_5929,N_5917);
and U6061 (N_6061,N_5953,N_5950);
nand U6062 (N_6062,N_5931,N_5962);
nand U6063 (N_6063,N_5957,N_5903);
nor U6064 (N_6064,N_5933,N_5982);
and U6065 (N_6065,N_5993,N_5931);
nand U6066 (N_6066,N_5913,N_5991);
nor U6067 (N_6067,N_5997,N_5941);
nor U6068 (N_6068,N_5957,N_5964);
and U6069 (N_6069,N_5937,N_5901);
nand U6070 (N_6070,N_5908,N_5935);
xor U6071 (N_6071,N_5988,N_5993);
or U6072 (N_6072,N_5964,N_5943);
and U6073 (N_6073,N_5958,N_5942);
xnor U6074 (N_6074,N_5945,N_5965);
xnor U6075 (N_6075,N_5914,N_5937);
nand U6076 (N_6076,N_5950,N_5971);
or U6077 (N_6077,N_5940,N_5900);
or U6078 (N_6078,N_5905,N_5912);
nand U6079 (N_6079,N_5989,N_5900);
and U6080 (N_6080,N_5956,N_5981);
or U6081 (N_6081,N_5934,N_5987);
or U6082 (N_6082,N_5974,N_5963);
nand U6083 (N_6083,N_5933,N_5955);
nand U6084 (N_6084,N_5973,N_5982);
and U6085 (N_6085,N_5951,N_5944);
nor U6086 (N_6086,N_5945,N_5934);
nor U6087 (N_6087,N_5964,N_5911);
nand U6088 (N_6088,N_5958,N_5972);
and U6089 (N_6089,N_5958,N_5981);
xor U6090 (N_6090,N_5939,N_5929);
or U6091 (N_6091,N_5922,N_5961);
or U6092 (N_6092,N_5994,N_5966);
and U6093 (N_6093,N_5952,N_5994);
xor U6094 (N_6094,N_5984,N_5934);
nand U6095 (N_6095,N_5995,N_5991);
and U6096 (N_6096,N_5988,N_5995);
xnor U6097 (N_6097,N_5926,N_5973);
xor U6098 (N_6098,N_5986,N_5933);
nor U6099 (N_6099,N_5970,N_5946);
and U6100 (N_6100,N_6025,N_6023);
and U6101 (N_6101,N_6045,N_6068);
nand U6102 (N_6102,N_6087,N_6033);
and U6103 (N_6103,N_6075,N_6035);
xnor U6104 (N_6104,N_6088,N_6002);
and U6105 (N_6105,N_6037,N_6026);
nand U6106 (N_6106,N_6083,N_6006);
or U6107 (N_6107,N_6056,N_6046);
or U6108 (N_6108,N_6061,N_6057);
nor U6109 (N_6109,N_6093,N_6040);
nand U6110 (N_6110,N_6010,N_6030);
xnor U6111 (N_6111,N_6073,N_6001);
or U6112 (N_6112,N_6039,N_6066);
nand U6113 (N_6113,N_6021,N_6022);
nor U6114 (N_6114,N_6012,N_6028);
nor U6115 (N_6115,N_6067,N_6071);
or U6116 (N_6116,N_6034,N_6044);
nand U6117 (N_6117,N_6011,N_6013);
and U6118 (N_6118,N_6097,N_6062);
xnor U6119 (N_6119,N_6047,N_6084);
nand U6120 (N_6120,N_6051,N_6099);
nor U6121 (N_6121,N_6081,N_6052);
and U6122 (N_6122,N_6032,N_6090);
or U6123 (N_6123,N_6082,N_6096);
or U6124 (N_6124,N_6048,N_6038);
or U6125 (N_6125,N_6000,N_6054);
or U6126 (N_6126,N_6092,N_6017);
nand U6127 (N_6127,N_6004,N_6041);
and U6128 (N_6128,N_6086,N_6072);
xor U6129 (N_6129,N_6003,N_6085);
nand U6130 (N_6130,N_6009,N_6027);
and U6131 (N_6131,N_6089,N_6055);
or U6132 (N_6132,N_6078,N_6080);
and U6133 (N_6133,N_6063,N_6005);
or U6134 (N_6134,N_6094,N_6074);
xnor U6135 (N_6135,N_6024,N_6036);
and U6136 (N_6136,N_6015,N_6016);
or U6137 (N_6137,N_6014,N_6019);
nor U6138 (N_6138,N_6079,N_6065);
xor U6139 (N_6139,N_6008,N_6007);
nor U6140 (N_6140,N_6020,N_6031);
nor U6141 (N_6141,N_6049,N_6043);
or U6142 (N_6142,N_6050,N_6069);
and U6143 (N_6143,N_6058,N_6042);
and U6144 (N_6144,N_6060,N_6095);
nor U6145 (N_6145,N_6077,N_6029);
and U6146 (N_6146,N_6059,N_6098);
xnor U6147 (N_6147,N_6064,N_6076);
nor U6148 (N_6148,N_6018,N_6053);
xor U6149 (N_6149,N_6091,N_6070);
nand U6150 (N_6150,N_6057,N_6059);
or U6151 (N_6151,N_6093,N_6085);
or U6152 (N_6152,N_6030,N_6035);
nor U6153 (N_6153,N_6024,N_6096);
and U6154 (N_6154,N_6025,N_6044);
xnor U6155 (N_6155,N_6028,N_6083);
xnor U6156 (N_6156,N_6060,N_6075);
and U6157 (N_6157,N_6078,N_6002);
nand U6158 (N_6158,N_6070,N_6012);
nor U6159 (N_6159,N_6095,N_6059);
nand U6160 (N_6160,N_6008,N_6096);
nand U6161 (N_6161,N_6097,N_6041);
and U6162 (N_6162,N_6049,N_6096);
nor U6163 (N_6163,N_6048,N_6040);
nor U6164 (N_6164,N_6026,N_6085);
nand U6165 (N_6165,N_6049,N_6010);
nand U6166 (N_6166,N_6050,N_6004);
or U6167 (N_6167,N_6046,N_6006);
and U6168 (N_6168,N_6031,N_6003);
and U6169 (N_6169,N_6045,N_6042);
or U6170 (N_6170,N_6048,N_6012);
nor U6171 (N_6171,N_6077,N_6078);
or U6172 (N_6172,N_6004,N_6094);
xor U6173 (N_6173,N_6010,N_6009);
and U6174 (N_6174,N_6053,N_6044);
or U6175 (N_6175,N_6089,N_6073);
nand U6176 (N_6176,N_6035,N_6029);
nand U6177 (N_6177,N_6000,N_6060);
xnor U6178 (N_6178,N_6080,N_6075);
or U6179 (N_6179,N_6018,N_6072);
nor U6180 (N_6180,N_6071,N_6041);
nor U6181 (N_6181,N_6013,N_6025);
nand U6182 (N_6182,N_6099,N_6030);
or U6183 (N_6183,N_6079,N_6055);
and U6184 (N_6184,N_6020,N_6084);
xor U6185 (N_6185,N_6082,N_6088);
and U6186 (N_6186,N_6003,N_6084);
and U6187 (N_6187,N_6002,N_6095);
nor U6188 (N_6188,N_6028,N_6058);
nor U6189 (N_6189,N_6053,N_6054);
nand U6190 (N_6190,N_6010,N_6076);
nor U6191 (N_6191,N_6083,N_6040);
or U6192 (N_6192,N_6063,N_6045);
and U6193 (N_6193,N_6030,N_6050);
and U6194 (N_6194,N_6085,N_6047);
nor U6195 (N_6195,N_6076,N_6035);
xor U6196 (N_6196,N_6032,N_6064);
or U6197 (N_6197,N_6027,N_6023);
or U6198 (N_6198,N_6059,N_6077);
nand U6199 (N_6199,N_6059,N_6019);
nor U6200 (N_6200,N_6123,N_6184);
nor U6201 (N_6201,N_6113,N_6129);
or U6202 (N_6202,N_6159,N_6155);
nor U6203 (N_6203,N_6180,N_6105);
xnor U6204 (N_6204,N_6109,N_6102);
nor U6205 (N_6205,N_6196,N_6191);
or U6206 (N_6206,N_6164,N_6125);
nor U6207 (N_6207,N_6170,N_6117);
or U6208 (N_6208,N_6190,N_6158);
or U6209 (N_6209,N_6130,N_6131);
and U6210 (N_6210,N_6118,N_6141);
nand U6211 (N_6211,N_6168,N_6136);
nor U6212 (N_6212,N_6193,N_6165);
and U6213 (N_6213,N_6150,N_6144);
nand U6214 (N_6214,N_6197,N_6153);
and U6215 (N_6215,N_6101,N_6177);
xnor U6216 (N_6216,N_6186,N_6124);
or U6217 (N_6217,N_6112,N_6192);
or U6218 (N_6218,N_6171,N_6115);
xor U6219 (N_6219,N_6167,N_6198);
or U6220 (N_6220,N_6119,N_6116);
xor U6221 (N_6221,N_6189,N_6140);
nor U6222 (N_6222,N_6135,N_6145);
and U6223 (N_6223,N_6100,N_6178);
or U6224 (N_6224,N_6195,N_6156);
nand U6225 (N_6225,N_6181,N_6187);
xnor U6226 (N_6226,N_6146,N_6160);
nand U6227 (N_6227,N_6128,N_6107);
and U6228 (N_6228,N_6134,N_6110);
or U6229 (N_6229,N_6133,N_6137);
nor U6230 (N_6230,N_6122,N_6157);
nand U6231 (N_6231,N_6174,N_6185);
and U6232 (N_6232,N_6149,N_6114);
and U6233 (N_6233,N_6199,N_6152);
xor U6234 (N_6234,N_6147,N_6188);
nor U6235 (N_6235,N_6106,N_6183);
and U6236 (N_6236,N_6176,N_6161);
or U6237 (N_6237,N_6148,N_6162);
xor U6238 (N_6238,N_6154,N_6120);
or U6239 (N_6239,N_6126,N_6169);
or U6240 (N_6240,N_6179,N_6104);
nor U6241 (N_6241,N_6151,N_6163);
and U6242 (N_6242,N_6194,N_6103);
or U6243 (N_6243,N_6142,N_6132);
and U6244 (N_6244,N_6127,N_6111);
xor U6245 (N_6245,N_6121,N_6166);
or U6246 (N_6246,N_6173,N_6139);
xor U6247 (N_6247,N_6172,N_6175);
nand U6248 (N_6248,N_6108,N_6143);
or U6249 (N_6249,N_6182,N_6138);
nor U6250 (N_6250,N_6119,N_6160);
xor U6251 (N_6251,N_6115,N_6163);
nand U6252 (N_6252,N_6147,N_6101);
xor U6253 (N_6253,N_6124,N_6110);
nand U6254 (N_6254,N_6133,N_6110);
and U6255 (N_6255,N_6147,N_6117);
nand U6256 (N_6256,N_6103,N_6151);
or U6257 (N_6257,N_6166,N_6179);
or U6258 (N_6258,N_6134,N_6135);
nor U6259 (N_6259,N_6124,N_6128);
nand U6260 (N_6260,N_6161,N_6127);
nand U6261 (N_6261,N_6159,N_6183);
xor U6262 (N_6262,N_6173,N_6170);
or U6263 (N_6263,N_6175,N_6154);
nor U6264 (N_6264,N_6159,N_6126);
or U6265 (N_6265,N_6122,N_6181);
xnor U6266 (N_6266,N_6180,N_6190);
nor U6267 (N_6267,N_6197,N_6104);
or U6268 (N_6268,N_6122,N_6192);
xor U6269 (N_6269,N_6168,N_6167);
xor U6270 (N_6270,N_6192,N_6127);
and U6271 (N_6271,N_6113,N_6192);
or U6272 (N_6272,N_6112,N_6133);
or U6273 (N_6273,N_6124,N_6139);
nor U6274 (N_6274,N_6186,N_6107);
and U6275 (N_6275,N_6156,N_6145);
or U6276 (N_6276,N_6102,N_6113);
or U6277 (N_6277,N_6178,N_6167);
and U6278 (N_6278,N_6162,N_6151);
and U6279 (N_6279,N_6135,N_6108);
or U6280 (N_6280,N_6110,N_6197);
or U6281 (N_6281,N_6143,N_6131);
xor U6282 (N_6282,N_6185,N_6179);
or U6283 (N_6283,N_6129,N_6187);
xor U6284 (N_6284,N_6103,N_6154);
or U6285 (N_6285,N_6182,N_6166);
nor U6286 (N_6286,N_6189,N_6145);
or U6287 (N_6287,N_6123,N_6178);
and U6288 (N_6288,N_6168,N_6145);
and U6289 (N_6289,N_6170,N_6168);
nand U6290 (N_6290,N_6143,N_6138);
nand U6291 (N_6291,N_6121,N_6192);
and U6292 (N_6292,N_6162,N_6184);
nand U6293 (N_6293,N_6177,N_6107);
and U6294 (N_6294,N_6111,N_6104);
nor U6295 (N_6295,N_6174,N_6150);
nand U6296 (N_6296,N_6106,N_6148);
nor U6297 (N_6297,N_6106,N_6147);
nor U6298 (N_6298,N_6161,N_6141);
nand U6299 (N_6299,N_6198,N_6166);
nor U6300 (N_6300,N_6201,N_6237);
nand U6301 (N_6301,N_6291,N_6258);
nand U6302 (N_6302,N_6289,N_6299);
nor U6303 (N_6303,N_6228,N_6294);
and U6304 (N_6304,N_6271,N_6281);
and U6305 (N_6305,N_6220,N_6240);
or U6306 (N_6306,N_6266,N_6268);
xor U6307 (N_6307,N_6288,N_6279);
or U6308 (N_6308,N_6254,N_6245);
nand U6309 (N_6309,N_6232,N_6260);
nand U6310 (N_6310,N_6248,N_6287);
or U6311 (N_6311,N_6269,N_6225);
xor U6312 (N_6312,N_6263,N_6223);
nor U6313 (N_6313,N_6253,N_6226);
nand U6314 (N_6314,N_6211,N_6216);
or U6315 (N_6315,N_6249,N_6219);
and U6316 (N_6316,N_6286,N_6290);
nor U6317 (N_6317,N_6292,N_6238);
nand U6318 (N_6318,N_6234,N_6277);
nor U6319 (N_6319,N_6282,N_6231);
nand U6320 (N_6320,N_6212,N_6285);
or U6321 (N_6321,N_6250,N_6205);
or U6322 (N_6322,N_6235,N_6257);
nor U6323 (N_6323,N_6242,N_6200);
or U6324 (N_6324,N_6243,N_6295);
and U6325 (N_6325,N_6241,N_6297);
nand U6326 (N_6326,N_6221,N_6207);
nor U6327 (N_6327,N_6217,N_6274);
nand U6328 (N_6328,N_6236,N_6255);
or U6329 (N_6329,N_6209,N_6204);
or U6330 (N_6330,N_6239,N_6296);
or U6331 (N_6331,N_6213,N_6229);
and U6332 (N_6332,N_6284,N_6283);
nand U6333 (N_6333,N_6218,N_6298);
xnor U6334 (N_6334,N_6233,N_6247);
xnor U6335 (N_6335,N_6224,N_6210);
and U6336 (N_6336,N_6214,N_6270);
and U6337 (N_6337,N_6261,N_6273);
and U6338 (N_6338,N_6252,N_6251);
nor U6339 (N_6339,N_6276,N_6246);
nand U6340 (N_6340,N_6227,N_6244);
and U6341 (N_6341,N_6208,N_6202);
nand U6342 (N_6342,N_6280,N_6230);
nand U6343 (N_6343,N_6262,N_6267);
nand U6344 (N_6344,N_6264,N_6256);
and U6345 (N_6345,N_6275,N_6203);
nand U6346 (N_6346,N_6222,N_6293);
xnor U6347 (N_6347,N_6278,N_6206);
nor U6348 (N_6348,N_6265,N_6272);
xor U6349 (N_6349,N_6259,N_6215);
or U6350 (N_6350,N_6289,N_6248);
nand U6351 (N_6351,N_6233,N_6238);
nor U6352 (N_6352,N_6257,N_6206);
or U6353 (N_6353,N_6201,N_6234);
nor U6354 (N_6354,N_6259,N_6275);
xnor U6355 (N_6355,N_6223,N_6293);
and U6356 (N_6356,N_6213,N_6233);
nor U6357 (N_6357,N_6246,N_6230);
and U6358 (N_6358,N_6290,N_6201);
or U6359 (N_6359,N_6255,N_6216);
or U6360 (N_6360,N_6201,N_6240);
xnor U6361 (N_6361,N_6250,N_6246);
nor U6362 (N_6362,N_6253,N_6283);
nand U6363 (N_6363,N_6252,N_6230);
nand U6364 (N_6364,N_6218,N_6201);
nand U6365 (N_6365,N_6218,N_6213);
nand U6366 (N_6366,N_6288,N_6217);
and U6367 (N_6367,N_6251,N_6233);
and U6368 (N_6368,N_6290,N_6236);
or U6369 (N_6369,N_6201,N_6254);
xnor U6370 (N_6370,N_6292,N_6245);
xnor U6371 (N_6371,N_6230,N_6279);
and U6372 (N_6372,N_6297,N_6249);
and U6373 (N_6373,N_6258,N_6226);
xnor U6374 (N_6374,N_6238,N_6295);
xnor U6375 (N_6375,N_6223,N_6262);
xor U6376 (N_6376,N_6230,N_6261);
xor U6377 (N_6377,N_6291,N_6251);
or U6378 (N_6378,N_6210,N_6250);
and U6379 (N_6379,N_6299,N_6297);
nor U6380 (N_6380,N_6227,N_6222);
xnor U6381 (N_6381,N_6209,N_6215);
nand U6382 (N_6382,N_6223,N_6279);
nand U6383 (N_6383,N_6256,N_6289);
and U6384 (N_6384,N_6261,N_6275);
nor U6385 (N_6385,N_6263,N_6249);
xor U6386 (N_6386,N_6204,N_6230);
or U6387 (N_6387,N_6240,N_6275);
and U6388 (N_6388,N_6288,N_6284);
and U6389 (N_6389,N_6240,N_6211);
nand U6390 (N_6390,N_6284,N_6257);
or U6391 (N_6391,N_6285,N_6244);
nand U6392 (N_6392,N_6205,N_6266);
nand U6393 (N_6393,N_6245,N_6269);
nor U6394 (N_6394,N_6271,N_6273);
nor U6395 (N_6395,N_6217,N_6276);
and U6396 (N_6396,N_6292,N_6266);
nor U6397 (N_6397,N_6219,N_6205);
or U6398 (N_6398,N_6223,N_6282);
and U6399 (N_6399,N_6293,N_6211);
nand U6400 (N_6400,N_6358,N_6329);
xnor U6401 (N_6401,N_6323,N_6379);
nor U6402 (N_6402,N_6387,N_6354);
nand U6403 (N_6403,N_6384,N_6328);
nor U6404 (N_6404,N_6381,N_6349);
nor U6405 (N_6405,N_6334,N_6399);
nor U6406 (N_6406,N_6389,N_6336);
xnor U6407 (N_6407,N_6306,N_6342);
xor U6408 (N_6408,N_6300,N_6353);
nor U6409 (N_6409,N_6348,N_6346);
and U6410 (N_6410,N_6317,N_6377);
and U6411 (N_6411,N_6373,N_6383);
nand U6412 (N_6412,N_6350,N_6397);
and U6413 (N_6413,N_6396,N_6340);
nand U6414 (N_6414,N_6335,N_6364);
or U6415 (N_6415,N_6366,N_6380);
nor U6416 (N_6416,N_6337,N_6347);
and U6417 (N_6417,N_6371,N_6357);
nand U6418 (N_6418,N_6339,N_6311);
or U6419 (N_6419,N_6363,N_6314);
xnor U6420 (N_6420,N_6356,N_6395);
nor U6421 (N_6421,N_6370,N_6375);
nor U6422 (N_6422,N_6326,N_6390);
or U6423 (N_6423,N_6312,N_6322);
or U6424 (N_6424,N_6302,N_6344);
nand U6425 (N_6425,N_6345,N_6325);
nor U6426 (N_6426,N_6318,N_6320);
or U6427 (N_6427,N_6301,N_6360);
nand U6428 (N_6428,N_6332,N_6308);
nand U6429 (N_6429,N_6310,N_6313);
or U6430 (N_6430,N_6385,N_6388);
and U6431 (N_6431,N_6341,N_6382);
or U6432 (N_6432,N_6359,N_6330);
nor U6433 (N_6433,N_6386,N_6338);
nand U6434 (N_6434,N_6352,N_6331);
nor U6435 (N_6435,N_6394,N_6304);
nand U6436 (N_6436,N_6368,N_6361);
nor U6437 (N_6437,N_6324,N_6315);
xor U6438 (N_6438,N_6343,N_6305);
or U6439 (N_6439,N_6392,N_6319);
nand U6440 (N_6440,N_6391,N_6355);
nand U6441 (N_6441,N_6378,N_6362);
or U6442 (N_6442,N_6367,N_6333);
or U6443 (N_6443,N_6374,N_6303);
or U6444 (N_6444,N_6316,N_6398);
xnor U6445 (N_6445,N_6376,N_6393);
nor U6446 (N_6446,N_6365,N_6372);
or U6447 (N_6447,N_6369,N_6309);
nand U6448 (N_6448,N_6327,N_6351);
and U6449 (N_6449,N_6307,N_6321);
xnor U6450 (N_6450,N_6391,N_6320);
nor U6451 (N_6451,N_6366,N_6338);
or U6452 (N_6452,N_6371,N_6340);
nand U6453 (N_6453,N_6304,N_6357);
and U6454 (N_6454,N_6374,N_6359);
nor U6455 (N_6455,N_6394,N_6372);
nand U6456 (N_6456,N_6387,N_6358);
nand U6457 (N_6457,N_6357,N_6359);
or U6458 (N_6458,N_6303,N_6367);
nand U6459 (N_6459,N_6387,N_6395);
nand U6460 (N_6460,N_6313,N_6311);
xor U6461 (N_6461,N_6337,N_6328);
xor U6462 (N_6462,N_6304,N_6342);
xnor U6463 (N_6463,N_6363,N_6396);
nor U6464 (N_6464,N_6378,N_6347);
nand U6465 (N_6465,N_6367,N_6356);
nand U6466 (N_6466,N_6352,N_6316);
nand U6467 (N_6467,N_6330,N_6303);
and U6468 (N_6468,N_6303,N_6333);
or U6469 (N_6469,N_6320,N_6379);
nand U6470 (N_6470,N_6344,N_6351);
nand U6471 (N_6471,N_6396,N_6386);
or U6472 (N_6472,N_6335,N_6388);
and U6473 (N_6473,N_6333,N_6308);
nand U6474 (N_6474,N_6312,N_6349);
xnor U6475 (N_6475,N_6391,N_6399);
nand U6476 (N_6476,N_6391,N_6309);
nand U6477 (N_6477,N_6356,N_6344);
nand U6478 (N_6478,N_6303,N_6380);
and U6479 (N_6479,N_6333,N_6393);
nor U6480 (N_6480,N_6355,N_6319);
nor U6481 (N_6481,N_6352,N_6357);
or U6482 (N_6482,N_6356,N_6382);
nand U6483 (N_6483,N_6392,N_6312);
or U6484 (N_6484,N_6381,N_6352);
nor U6485 (N_6485,N_6319,N_6339);
xor U6486 (N_6486,N_6318,N_6319);
xor U6487 (N_6487,N_6345,N_6362);
nand U6488 (N_6488,N_6348,N_6350);
nor U6489 (N_6489,N_6393,N_6386);
nand U6490 (N_6490,N_6347,N_6306);
nand U6491 (N_6491,N_6392,N_6388);
nor U6492 (N_6492,N_6337,N_6315);
nor U6493 (N_6493,N_6326,N_6301);
xnor U6494 (N_6494,N_6396,N_6393);
nand U6495 (N_6495,N_6331,N_6365);
nor U6496 (N_6496,N_6388,N_6386);
or U6497 (N_6497,N_6397,N_6321);
nor U6498 (N_6498,N_6388,N_6318);
xnor U6499 (N_6499,N_6311,N_6390);
xnor U6500 (N_6500,N_6442,N_6491);
and U6501 (N_6501,N_6476,N_6448);
nand U6502 (N_6502,N_6474,N_6452);
nand U6503 (N_6503,N_6435,N_6450);
nand U6504 (N_6504,N_6464,N_6441);
nor U6505 (N_6505,N_6408,N_6420);
nor U6506 (N_6506,N_6413,N_6456);
or U6507 (N_6507,N_6454,N_6445);
or U6508 (N_6508,N_6449,N_6496);
or U6509 (N_6509,N_6440,N_6467);
nor U6510 (N_6510,N_6418,N_6402);
nand U6511 (N_6511,N_6473,N_6498);
nor U6512 (N_6512,N_6443,N_6490);
nand U6513 (N_6513,N_6499,N_6436);
or U6514 (N_6514,N_6416,N_6478);
and U6515 (N_6515,N_6429,N_6461);
nor U6516 (N_6516,N_6471,N_6486);
and U6517 (N_6517,N_6428,N_6489);
nor U6518 (N_6518,N_6400,N_6434);
and U6519 (N_6519,N_6472,N_6403);
nand U6520 (N_6520,N_6495,N_6477);
or U6521 (N_6521,N_6444,N_6488);
nor U6522 (N_6522,N_6446,N_6417);
or U6523 (N_6523,N_6401,N_6451);
xnor U6524 (N_6524,N_6479,N_6447);
and U6525 (N_6525,N_6484,N_6458);
nor U6526 (N_6526,N_6465,N_6427);
or U6527 (N_6527,N_6480,N_6430);
xor U6528 (N_6528,N_6469,N_6439);
nor U6529 (N_6529,N_6409,N_6415);
or U6530 (N_6530,N_6492,N_6466);
or U6531 (N_6531,N_6482,N_6483);
and U6532 (N_6532,N_6437,N_6406);
and U6533 (N_6533,N_6468,N_6412);
nor U6534 (N_6534,N_6470,N_6410);
xor U6535 (N_6535,N_6485,N_6493);
xnor U6536 (N_6536,N_6481,N_6419);
xnor U6537 (N_6537,N_6455,N_6487);
and U6538 (N_6538,N_6414,N_6423);
xor U6539 (N_6539,N_6475,N_6425);
xnor U6540 (N_6540,N_6433,N_6431);
xor U6541 (N_6541,N_6404,N_6453);
nand U6542 (N_6542,N_6459,N_6411);
and U6543 (N_6543,N_6497,N_6405);
or U6544 (N_6544,N_6422,N_6460);
or U6545 (N_6545,N_6494,N_6407);
nand U6546 (N_6546,N_6424,N_6421);
nand U6547 (N_6547,N_6463,N_6432);
and U6548 (N_6548,N_6462,N_6457);
xor U6549 (N_6549,N_6438,N_6426);
and U6550 (N_6550,N_6401,N_6474);
and U6551 (N_6551,N_6471,N_6420);
xnor U6552 (N_6552,N_6475,N_6406);
nand U6553 (N_6553,N_6403,N_6407);
xor U6554 (N_6554,N_6469,N_6440);
or U6555 (N_6555,N_6407,N_6482);
nor U6556 (N_6556,N_6479,N_6456);
xor U6557 (N_6557,N_6435,N_6425);
and U6558 (N_6558,N_6411,N_6485);
nor U6559 (N_6559,N_6414,N_6479);
nor U6560 (N_6560,N_6405,N_6458);
nor U6561 (N_6561,N_6406,N_6455);
nor U6562 (N_6562,N_6437,N_6461);
and U6563 (N_6563,N_6433,N_6496);
nor U6564 (N_6564,N_6467,N_6430);
nand U6565 (N_6565,N_6476,N_6411);
or U6566 (N_6566,N_6448,N_6443);
nand U6567 (N_6567,N_6459,N_6499);
xnor U6568 (N_6568,N_6449,N_6406);
xor U6569 (N_6569,N_6472,N_6490);
or U6570 (N_6570,N_6407,N_6405);
and U6571 (N_6571,N_6432,N_6470);
nand U6572 (N_6572,N_6419,N_6485);
or U6573 (N_6573,N_6463,N_6409);
xor U6574 (N_6574,N_6472,N_6450);
nor U6575 (N_6575,N_6486,N_6464);
xnor U6576 (N_6576,N_6490,N_6407);
xnor U6577 (N_6577,N_6438,N_6497);
and U6578 (N_6578,N_6466,N_6445);
xnor U6579 (N_6579,N_6433,N_6463);
or U6580 (N_6580,N_6416,N_6417);
nor U6581 (N_6581,N_6494,N_6410);
xnor U6582 (N_6582,N_6408,N_6448);
xor U6583 (N_6583,N_6446,N_6443);
and U6584 (N_6584,N_6421,N_6469);
xor U6585 (N_6585,N_6436,N_6406);
and U6586 (N_6586,N_6402,N_6455);
xnor U6587 (N_6587,N_6453,N_6487);
xnor U6588 (N_6588,N_6472,N_6457);
xor U6589 (N_6589,N_6430,N_6428);
xnor U6590 (N_6590,N_6449,N_6412);
or U6591 (N_6591,N_6480,N_6483);
xnor U6592 (N_6592,N_6457,N_6434);
nor U6593 (N_6593,N_6404,N_6426);
nand U6594 (N_6594,N_6440,N_6456);
nand U6595 (N_6595,N_6498,N_6410);
or U6596 (N_6596,N_6441,N_6483);
or U6597 (N_6597,N_6463,N_6415);
nor U6598 (N_6598,N_6482,N_6432);
or U6599 (N_6599,N_6460,N_6423);
nor U6600 (N_6600,N_6540,N_6589);
and U6601 (N_6601,N_6507,N_6537);
xor U6602 (N_6602,N_6522,N_6547);
nor U6603 (N_6603,N_6519,N_6565);
or U6604 (N_6604,N_6551,N_6593);
and U6605 (N_6605,N_6553,N_6567);
nand U6606 (N_6606,N_6550,N_6587);
nor U6607 (N_6607,N_6581,N_6594);
and U6608 (N_6608,N_6542,N_6583);
nor U6609 (N_6609,N_6541,N_6520);
nand U6610 (N_6610,N_6576,N_6585);
xnor U6611 (N_6611,N_6568,N_6518);
nor U6612 (N_6612,N_6577,N_6500);
or U6613 (N_6613,N_6513,N_6526);
or U6614 (N_6614,N_6562,N_6552);
or U6615 (N_6615,N_6566,N_6554);
and U6616 (N_6616,N_6502,N_6536);
and U6617 (N_6617,N_6514,N_6530);
nand U6618 (N_6618,N_6549,N_6521);
and U6619 (N_6619,N_6591,N_6511);
nor U6620 (N_6620,N_6509,N_6557);
nand U6621 (N_6621,N_6597,N_6525);
nor U6622 (N_6622,N_6501,N_6574);
xnor U6623 (N_6623,N_6586,N_6548);
or U6624 (N_6624,N_6524,N_6598);
nand U6625 (N_6625,N_6506,N_6532);
xor U6626 (N_6626,N_6582,N_6575);
or U6627 (N_6627,N_6544,N_6516);
nor U6628 (N_6628,N_6578,N_6558);
or U6629 (N_6629,N_6564,N_6563);
nand U6630 (N_6630,N_6560,N_6539);
and U6631 (N_6631,N_6571,N_6538);
xor U6632 (N_6632,N_6555,N_6510);
nor U6633 (N_6633,N_6545,N_6599);
and U6634 (N_6634,N_6527,N_6517);
and U6635 (N_6635,N_6570,N_6561);
nand U6636 (N_6636,N_6531,N_6508);
or U6637 (N_6637,N_6503,N_6595);
nor U6638 (N_6638,N_6512,N_6579);
nand U6639 (N_6639,N_6572,N_6573);
or U6640 (N_6640,N_6580,N_6590);
nand U6641 (N_6641,N_6535,N_6592);
nor U6642 (N_6642,N_6534,N_6543);
xor U6643 (N_6643,N_6515,N_6546);
nor U6644 (N_6644,N_6504,N_6528);
xor U6645 (N_6645,N_6596,N_6588);
and U6646 (N_6646,N_6505,N_6556);
and U6647 (N_6647,N_6584,N_6569);
xor U6648 (N_6648,N_6533,N_6559);
nor U6649 (N_6649,N_6523,N_6529);
or U6650 (N_6650,N_6594,N_6585);
or U6651 (N_6651,N_6521,N_6566);
or U6652 (N_6652,N_6522,N_6578);
xnor U6653 (N_6653,N_6579,N_6582);
nand U6654 (N_6654,N_6535,N_6585);
nor U6655 (N_6655,N_6565,N_6550);
xor U6656 (N_6656,N_6557,N_6523);
or U6657 (N_6657,N_6582,N_6545);
and U6658 (N_6658,N_6576,N_6524);
nand U6659 (N_6659,N_6578,N_6565);
nor U6660 (N_6660,N_6597,N_6524);
and U6661 (N_6661,N_6571,N_6533);
xor U6662 (N_6662,N_6566,N_6542);
nand U6663 (N_6663,N_6505,N_6529);
and U6664 (N_6664,N_6517,N_6593);
xor U6665 (N_6665,N_6526,N_6581);
or U6666 (N_6666,N_6581,N_6537);
nor U6667 (N_6667,N_6553,N_6540);
nand U6668 (N_6668,N_6515,N_6584);
or U6669 (N_6669,N_6522,N_6586);
and U6670 (N_6670,N_6586,N_6510);
nor U6671 (N_6671,N_6580,N_6504);
nor U6672 (N_6672,N_6549,N_6522);
xnor U6673 (N_6673,N_6557,N_6524);
or U6674 (N_6674,N_6590,N_6586);
xor U6675 (N_6675,N_6542,N_6512);
and U6676 (N_6676,N_6520,N_6537);
nand U6677 (N_6677,N_6552,N_6517);
and U6678 (N_6678,N_6529,N_6597);
nand U6679 (N_6679,N_6518,N_6508);
nor U6680 (N_6680,N_6545,N_6548);
and U6681 (N_6681,N_6539,N_6567);
or U6682 (N_6682,N_6582,N_6590);
xnor U6683 (N_6683,N_6562,N_6571);
xor U6684 (N_6684,N_6519,N_6514);
or U6685 (N_6685,N_6595,N_6576);
nand U6686 (N_6686,N_6549,N_6540);
or U6687 (N_6687,N_6590,N_6542);
nand U6688 (N_6688,N_6500,N_6593);
nor U6689 (N_6689,N_6562,N_6547);
and U6690 (N_6690,N_6566,N_6578);
or U6691 (N_6691,N_6591,N_6599);
nand U6692 (N_6692,N_6535,N_6587);
and U6693 (N_6693,N_6566,N_6582);
and U6694 (N_6694,N_6596,N_6518);
nor U6695 (N_6695,N_6527,N_6529);
or U6696 (N_6696,N_6552,N_6523);
nand U6697 (N_6697,N_6537,N_6567);
and U6698 (N_6698,N_6582,N_6593);
and U6699 (N_6699,N_6549,N_6568);
nor U6700 (N_6700,N_6612,N_6639);
nor U6701 (N_6701,N_6690,N_6637);
xnor U6702 (N_6702,N_6630,N_6613);
or U6703 (N_6703,N_6627,N_6663);
nor U6704 (N_6704,N_6691,N_6606);
nor U6705 (N_6705,N_6664,N_6638);
nand U6706 (N_6706,N_6635,N_6694);
nor U6707 (N_6707,N_6695,N_6628);
and U6708 (N_6708,N_6699,N_6611);
and U6709 (N_6709,N_6661,N_6678);
or U6710 (N_6710,N_6692,N_6682);
or U6711 (N_6711,N_6684,N_6659);
nand U6712 (N_6712,N_6672,N_6668);
nand U6713 (N_6713,N_6604,N_6620);
nand U6714 (N_6714,N_6636,N_6629);
or U6715 (N_6715,N_6660,N_6669);
xor U6716 (N_6716,N_6646,N_6618);
or U6717 (N_6717,N_6651,N_6674);
or U6718 (N_6718,N_6656,N_6679);
or U6719 (N_6719,N_6688,N_6696);
or U6720 (N_6720,N_6697,N_6677);
and U6721 (N_6721,N_6641,N_6640);
nor U6722 (N_6722,N_6634,N_6645);
nor U6723 (N_6723,N_6654,N_6653);
nand U6724 (N_6724,N_6626,N_6621);
nor U6725 (N_6725,N_6658,N_6631);
nor U6726 (N_6726,N_6676,N_6642);
and U6727 (N_6727,N_6673,N_6644);
and U6728 (N_6728,N_6608,N_6652);
or U6729 (N_6729,N_6648,N_6609);
or U6730 (N_6730,N_6622,N_6685);
and U6731 (N_6731,N_6600,N_6615);
nor U6732 (N_6732,N_6662,N_6625);
xnor U6733 (N_6733,N_6698,N_6671);
or U6734 (N_6734,N_6667,N_6693);
nor U6735 (N_6735,N_6624,N_6632);
xor U6736 (N_6736,N_6601,N_6650);
and U6737 (N_6737,N_6603,N_6617);
nand U6738 (N_6738,N_6683,N_6689);
and U6739 (N_6739,N_6619,N_6665);
xnor U6740 (N_6740,N_6647,N_6607);
and U6741 (N_6741,N_6623,N_6649);
or U6742 (N_6742,N_6657,N_6616);
nand U6743 (N_6743,N_6666,N_6675);
nor U6744 (N_6744,N_6670,N_6643);
or U6745 (N_6745,N_6681,N_6686);
nand U6746 (N_6746,N_6680,N_6655);
nor U6747 (N_6747,N_6602,N_6687);
or U6748 (N_6748,N_6633,N_6614);
or U6749 (N_6749,N_6605,N_6610);
nand U6750 (N_6750,N_6627,N_6616);
nand U6751 (N_6751,N_6683,N_6684);
nor U6752 (N_6752,N_6688,N_6652);
xor U6753 (N_6753,N_6645,N_6678);
nor U6754 (N_6754,N_6695,N_6613);
and U6755 (N_6755,N_6626,N_6672);
xnor U6756 (N_6756,N_6656,N_6662);
and U6757 (N_6757,N_6620,N_6655);
nor U6758 (N_6758,N_6634,N_6684);
nand U6759 (N_6759,N_6619,N_6664);
nand U6760 (N_6760,N_6629,N_6606);
or U6761 (N_6761,N_6647,N_6669);
xnor U6762 (N_6762,N_6645,N_6616);
or U6763 (N_6763,N_6692,N_6601);
or U6764 (N_6764,N_6650,N_6665);
nand U6765 (N_6765,N_6638,N_6690);
or U6766 (N_6766,N_6684,N_6674);
nor U6767 (N_6767,N_6661,N_6696);
nor U6768 (N_6768,N_6600,N_6665);
or U6769 (N_6769,N_6664,N_6694);
xnor U6770 (N_6770,N_6668,N_6657);
or U6771 (N_6771,N_6606,N_6619);
nor U6772 (N_6772,N_6672,N_6685);
nand U6773 (N_6773,N_6653,N_6605);
nand U6774 (N_6774,N_6668,N_6684);
nand U6775 (N_6775,N_6612,N_6684);
nor U6776 (N_6776,N_6674,N_6694);
and U6777 (N_6777,N_6683,N_6628);
nand U6778 (N_6778,N_6664,N_6674);
and U6779 (N_6779,N_6652,N_6648);
nor U6780 (N_6780,N_6642,N_6674);
and U6781 (N_6781,N_6625,N_6615);
and U6782 (N_6782,N_6665,N_6655);
xor U6783 (N_6783,N_6600,N_6675);
nand U6784 (N_6784,N_6697,N_6672);
nor U6785 (N_6785,N_6656,N_6602);
xor U6786 (N_6786,N_6692,N_6688);
xor U6787 (N_6787,N_6606,N_6601);
and U6788 (N_6788,N_6698,N_6629);
nor U6789 (N_6789,N_6630,N_6647);
or U6790 (N_6790,N_6654,N_6696);
nand U6791 (N_6791,N_6654,N_6626);
xor U6792 (N_6792,N_6609,N_6656);
or U6793 (N_6793,N_6655,N_6642);
nand U6794 (N_6794,N_6641,N_6645);
and U6795 (N_6795,N_6658,N_6688);
nor U6796 (N_6796,N_6699,N_6686);
or U6797 (N_6797,N_6685,N_6631);
nor U6798 (N_6798,N_6695,N_6654);
nor U6799 (N_6799,N_6698,N_6645);
and U6800 (N_6800,N_6760,N_6798);
and U6801 (N_6801,N_6796,N_6721);
or U6802 (N_6802,N_6730,N_6712);
nor U6803 (N_6803,N_6701,N_6757);
xor U6804 (N_6804,N_6715,N_6735);
nor U6805 (N_6805,N_6767,N_6719);
and U6806 (N_6806,N_6705,N_6766);
or U6807 (N_6807,N_6770,N_6764);
and U6808 (N_6808,N_6758,N_6744);
nor U6809 (N_6809,N_6709,N_6729);
nand U6810 (N_6810,N_6741,N_6753);
and U6811 (N_6811,N_6771,N_6714);
nand U6812 (N_6812,N_6734,N_6786);
nand U6813 (N_6813,N_6713,N_6752);
nand U6814 (N_6814,N_6780,N_6772);
or U6815 (N_6815,N_6726,N_6728);
nand U6816 (N_6816,N_6756,N_6716);
or U6817 (N_6817,N_6790,N_6788);
and U6818 (N_6818,N_6710,N_6779);
nor U6819 (N_6819,N_6759,N_6738);
or U6820 (N_6820,N_6711,N_6727);
and U6821 (N_6821,N_6795,N_6700);
and U6822 (N_6822,N_6725,N_6782);
nand U6823 (N_6823,N_6704,N_6792);
or U6824 (N_6824,N_6754,N_6748);
xnor U6825 (N_6825,N_6784,N_6775);
xor U6826 (N_6826,N_6736,N_6783);
nor U6827 (N_6827,N_6791,N_6706);
nand U6828 (N_6828,N_6797,N_6743);
xnor U6829 (N_6829,N_6702,N_6750);
xnor U6830 (N_6830,N_6787,N_6740);
or U6831 (N_6831,N_6794,N_6793);
or U6832 (N_6832,N_6703,N_6742);
xor U6833 (N_6833,N_6731,N_6733);
nor U6834 (N_6834,N_6781,N_6747);
nand U6835 (N_6835,N_6799,N_6739);
or U6836 (N_6836,N_6763,N_6707);
nand U6837 (N_6837,N_6724,N_6762);
nand U6838 (N_6838,N_6737,N_6778);
nand U6839 (N_6839,N_6718,N_6745);
nor U6840 (N_6840,N_6720,N_6776);
xor U6841 (N_6841,N_6765,N_6769);
or U6842 (N_6842,N_6749,N_6761);
or U6843 (N_6843,N_6773,N_6717);
and U6844 (N_6844,N_6768,N_6789);
or U6845 (N_6845,N_6708,N_6777);
xor U6846 (N_6846,N_6722,N_6751);
or U6847 (N_6847,N_6755,N_6774);
xor U6848 (N_6848,N_6746,N_6785);
xnor U6849 (N_6849,N_6723,N_6732);
nand U6850 (N_6850,N_6770,N_6727);
nor U6851 (N_6851,N_6762,N_6768);
or U6852 (N_6852,N_6739,N_6769);
xor U6853 (N_6853,N_6708,N_6706);
or U6854 (N_6854,N_6735,N_6747);
xor U6855 (N_6855,N_6764,N_6735);
and U6856 (N_6856,N_6751,N_6725);
nand U6857 (N_6857,N_6770,N_6765);
nor U6858 (N_6858,N_6746,N_6740);
xnor U6859 (N_6859,N_6777,N_6748);
and U6860 (N_6860,N_6733,N_6762);
or U6861 (N_6861,N_6743,N_6786);
nand U6862 (N_6862,N_6770,N_6753);
xor U6863 (N_6863,N_6749,N_6725);
or U6864 (N_6864,N_6762,N_6726);
xor U6865 (N_6865,N_6740,N_6765);
and U6866 (N_6866,N_6783,N_6787);
nor U6867 (N_6867,N_6716,N_6779);
and U6868 (N_6868,N_6733,N_6787);
xnor U6869 (N_6869,N_6725,N_6733);
xnor U6870 (N_6870,N_6759,N_6789);
nand U6871 (N_6871,N_6798,N_6736);
and U6872 (N_6872,N_6767,N_6748);
or U6873 (N_6873,N_6788,N_6784);
or U6874 (N_6874,N_6784,N_6703);
xor U6875 (N_6875,N_6746,N_6725);
nand U6876 (N_6876,N_6704,N_6720);
xor U6877 (N_6877,N_6741,N_6781);
xnor U6878 (N_6878,N_6757,N_6718);
and U6879 (N_6879,N_6792,N_6768);
xnor U6880 (N_6880,N_6771,N_6772);
nor U6881 (N_6881,N_6730,N_6786);
nand U6882 (N_6882,N_6743,N_6767);
xnor U6883 (N_6883,N_6721,N_6744);
nor U6884 (N_6884,N_6701,N_6748);
xor U6885 (N_6885,N_6703,N_6700);
nand U6886 (N_6886,N_6794,N_6733);
xor U6887 (N_6887,N_6756,N_6713);
nor U6888 (N_6888,N_6722,N_6717);
nand U6889 (N_6889,N_6748,N_6757);
and U6890 (N_6890,N_6772,N_6760);
or U6891 (N_6891,N_6791,N_6780);
nand U6892 (N_6892,N_6761,N_6722);
nand U6893 (N_6893,N_6737,N_6731);
nand U6894 (N_6894,N_6777,N_6715);
nand U6895 (N_6895,N_6703,N_6734);
nor U6896 (N_6896,N_6788,N_6773);
nand U6897 (N_6897,N_6729,N_6799);
or U6898 (N_6898,N_6742,N_6769);
nand U6899 (N_6899,N_6796,N_6723);
or U6900 (N_6900,N_6820,N_6870);
or U6901 (N_6901,N_6818,N_6803);
nand U6902 (N_6902,N_6852,N_6865);
nor U6903 (N_6903,N_6888,N_6806);
and U6904 (N_6904,N_6807,N_6810);
xor U6905 (N_6905,N_6883,N_6882);
or U6906 (N_6906,N_6873,N_6838);
and U6907 (N_6907,N_6813,N_6866);
and U6908 (N_6908,N_6841,N_6881);
or U6909 (N_6909,N_6860,N_6899);
and U6910 (N_6910,N_6804,N_6875);
nor U6911 (N_6911,N_6862,N_6809);
or U6912 (N_6912,N_6815,N_6876);
xnor U6913 (N_6913,N_6871,N_6892);
nand U6914 (N_6914,N_6829,N_6808);
and U6915 (N_6915,N_6879,N_6885);
xor U6916 (N_6916,N_6833,N_6834);
nor U6917 (N_6917,N_6880,N_6802);
or U6918 (N_6918,N_6811,N_6821);
xor U6919 (N_6919,N_6824,N_6817);
xnor U6920 (N_6920,N_6835,N_6800);
nor U6921 (N_6921,N_6840,N_6851);
and U6922 (N_6922,N_6891,N_6812);
nor U6923 (N_6923,N_6854,N_6877);
or U6924 (N_6924,N_6826,N_6867);
and U6925 (N_6925,N_6816,N_6842);
nand U6926 (N_6926,N_6889,N_6861);
xnor U6927 (N_6927,N_6832,N_6853);
nor U6928 (N_6928,N_6836,N_6805);
xor U6929 (N_6929,N_6859,N_6801);
and U6930 (N_6930,N_6845,N_6896);
xor U6931 (N_6931,N_6869,N_6872);
nor U6932 (N_6932,N_6890,N_6831);
nand U6933 (N_6933,N_6828,N_6837);
nor U6934 (N_6934,N_6874,N_6897);
nand U6935 (N_6935,N_6893,N_6864);
xnor U6936 (N_6936,N_6878,N_6827);
or U6937 (N_6937,N_6819,N_6868);
xor U6938 (N_6938,N_6886,N_6823);
nor U6939 (N_6939,N_6822,N_6858);
and U6940 (N_6940,N_6825,N_6814);
xnor U6941 (N_6941,N_6898,N_6847);
nand U6942 (N_6942,N_6856,N_6857);
xnor U6943 (N_6943,N_6844,N_6846);
and U6944 (N_6944,N_6830,N_6848);
and U6945 (N_6945,N_6850,N_6884);
or U6946 (N_6946,N_6894,N_6849);
nand U6947 (N_6947,N_6839,N_6887);
or U6948 (N_6948,N_6843,N_6863);
xor U6949 (N_6949,N_6855,N_6895);
or U6950 (N_6950,N_6827,N_6829);
nor U6951 (N_6951,N_6828,N_6819);
and U6952 (N_6952,N_6869,N_6842);
or U6953 (N_6953,N_6861,N_6896);
xnor U6954 (N_6954,N_6890,N_6840);
xor U6955 (N_6955,N_6852,N_6838);
nand U6956 (N_6956,N_6898,N_6864);
xnor U6957 (N_6957,N_6829,N_6893);
xor U6958 (N_6958,N_6868,N_6871);
nand U6959 (N_6959,N_6878,N_6847);
nand U6960 (N_6960,N_6803,N_6800);
nand U6961 (N_6961,N_6836,N_6871);
or U6962 (N_6962,N_6804,N_6871);
or U6963 (N_6963,N_6869,N_6853);
nand U6964 (N_6964,N_6890,N_6872);
nand U6965 (N_6965,N_6854,N_6869);
nand U6966 (N_6966,N_6898,N_6848);
xnor U6967 (N_6967,N_6849,N_6883);
nor U6968 (N_6968,N_6884,N_6879);
and U6969 (N_6969,N_6857,N_6876);
and U6970 (N_6970,N_6893,N_6884);
xnor U6971 (N_6971,N_6855,N_6820);
nand U6972 (N_6972,N_6841,N_6889);
xor U6973 (N_6973,N_6831,N_6843);
xnor U6974 (N_6974,N_6853,N_6858);
or U6975 (N_6975,N_6821,N_6896);
nand U6976 (N_6976,N_6837,N_6827);
or U6977 (N_6977,N_6851,N_6832);
or U6978 (N_6978,N_6899,N_6823);
nand U6979 (N_6979,N_6835,N_6871);
or U6980 (N_6980,N_6854,N_6875);
or U6981 (N_6981,N_6877,N_6875);
and U6982 (N_6982,N_6896,N_6893);
xor U6983 (N_6983,N_6885,N_6839);
nand U6984 (N_6984,N_6803,N_6865);
nor U6985 (N_6985,N_6854,N_6828);
xnor U6986 (N_6986,N_6891,N_6848);
nand U6987 (N_6987,N_6894,N_6824);
or U6988 (N_6988,N_6824,N_6895);
or U6989 (N_6989,N_6830,N_6845);
xor U6990 (N_6990,N_6896,N_6807);
xnor U6991 (N_6991,N_6898,N_6837);
xnor U6992 (N_6992,N_6879,N_6875);
or U6993 (N_6993,N_6891,N_6863);
nand U6994 (N_6994,N_6828,N_6821);
or U6995 (N_6995,N_6854,N_6865);
and U6996 (N_6996,N_6857,N_6877);
and U6997 (N_6997,N_6825,N_6869);
nor U6998 (N_6998,N_6849,N_6870);
nand U6999 (N_6999,N_6853,N_6828);
or U7000 (N_7000,N_6952,N_6970);
nor U7001 (N_7001,N_6995,N_6911);
nand U7002 (N_7002,N_6950,N_6975);
or U7003 (N_7003,N_6993,N_6974);
nor U7004 (N_7004,N_6927,N_6964);
and U7005 (N_7005,N_6939,N_6999);
nand U7006 (N_7006,N_6988,N_6987);
nor U7007 (N_7007,N_6981,N_6976);
nor U7008 (N_7008,N_6957,N_6926);
xnor U7009 (N_7009,N_6990,N_6904);
xor U7010 (N_7010,N_6979,N_6953);
nand U7011 (N_7011,N_6902,N_6934);
and U7012 (N_7012,N_6905,N_6985);
nand U7013 (N_7013,N_6960,N_6932);
or U7014 (N_7014,N_6903,N_6963);
nand U7015 (N_7015,N_6968,N_6977);
nand U7016 (N_7016,N_6966,N_6978);
nand U7017 (N_7017,N_6922,N_6928);
and U7018 (N_7018,N_6980,N_6943);
xnor U7019 (N_7019,N_6984,N_6931);
and U7020 (N_7020,N_6951,N_6910);
or U7021 (N_7021,N_6941,N_6938);
xnor U7022 (N_7022,N_6992,N_6923);
nor U7023 (N_7023,N_6986,N_6913);
xor U7024 (N_7024,N_6973,N_6959);
and U7025 (N_7025,N_6914,N_6940);
nand U7026 (N_7026,N_6949,N_6989);
nand U7027 (N_7027,N_6906,N_6965);
xor U7028 (N_7028,N_6920,N_6945);
xor U7029 (N_7029,N_6936,N_6962);
xor U7030 (N_7030,N_6907,N_6954);
nor U7031 (N_7031,N_6994,N_6935);
xor U7032 (N_7032,N_6915,N_6917);
nand U7033 (N_7033,N_6909,N_6946);
nand U7034 (N_7034,N_6944,N_6958);
and U7035 (N_7035,N_6983,N_6947);
xor U7036 (N_7036,N_6912,N_6982);
xor U7037 (N_7037,N_6972,N_6933);
or U7038 (N_7038,N_6924,N_6948);
and U7039 (N_7039,N_6955,N_6996);
xor U7040 (N_7040,N_6997,N_6908);
or U7041 (N_7041,N_6967,N_6921);
nand U7042 (N_7042,N_6991,N_6971);
or U7043 (N_7043,N_6901,N_6929);
nor U7044 (N_7044,N_6998,N_6918);
xnor U7045 (N_7045,N_6969,N_6961);
and U7046 (N_7046,N_6916,N_6937);
or U7047 (N_7047,N_6900,N_6956);
nand U7048 (N_7048,N_6930,N_6942);
nand U7049 (N_7049,N_6925,N_6919);
nor U7050 (N_7050,N_6959,N_6996);
xnor U7051 (N_7051,N_6945,N_6951);
xor U7052 (N_7052,N_6924,N_6902);
nand U7053 (N_7053,N_6933,N_6908);
nor U7054 (N_7054,N_6994,N_6997);
xnor U7055 (N_7055,N_6983,N_6981);
xor U7056 (N_7056,N_6908,N_6979);
and U7057 (N_7057,N_6942,N_6953);
nand U7058 (N_7058,N_6962,N_6929);
xor U7059 (N_7059,N_6982,N_6911);
xor U7060 (N_7060,N_6910,N_6999);
xnor U7061 (N_7061,N_6907,N_6926);
nand U7062 (N_7062,N_6990,N_6958);
or U7063 (N_7063,N_6922,N_6918);
nor U7064 (N_7064,N_6944,N_6970);
and U7065 (N_7065,N_6956,N_6975);
or U7066 (N_7066,N_6995,N_6946);
and U7067 (N_7067,N_6946,N_6947);
or U7068 (N_7068,N_6909,N_6947);
and U7069 (N_7069,N_6974,N_6927);
and U7070 (N_7070,N_6903,N_6912);
nor U7071 (N_7071,N_6993,N_6988);
and U7072 (N_7072,N_6972,N_6997);
or U7073 (N_7073,N_6951,N_6920);
nand U7074 (N_7074,N_6916,N_6934);
xnor U7075 (N_7075,N_6978,N_6925);
nand U7076 (N_7076,N_6946,N_6928);
or U7077 (N_7077,N_6961,N_6985);
nor U7078 (N_7078,N_6948,N_6976);
or U7079 (N_7079,N_6981,N_6953);
and U7080 (N_7080,N_6939,N_6969);
nand U7081 (N_7081,N_6904,N_6929);
and U7082 (N_7082,N_6903,N_6980);
nand U7083 (N_7083,N_6953,N_6972);
xnor U7084 (N_7084,N_6949,N_6960);
nor U7085 (N_7085,N_6931,N_6953);
nand U7086 (N_7086,N_6906,N_6911);
nor U7087 (N_7087,N_6965,N_6901);
or U7088 (N_7088,N_6956,N_6931);
or U7089 (N_7089,N_6993,N_6947);
xor U7090 (N_7090,N_6979,N_6976);
nand U7091 (N_7091,N_6916,N_6965);
xor U7092 (N_7092,N_6908,N_6929);
nand U7093 (N_7093,N_6916,N_6924);
xnor U7094 (N_7094,N_6975,N_6966);
or U7095 (N_7095,N_6973,N_6936);
or U7096 (N_7096,N_6933,N_6905);
nor U7097 (N_7097,N_6929,N_6967);
nand U7098 (N_7098,N_6927,N_6962);
and U7099 (N_7099,N_6969,N_6974);
or U7100 (N_7100,N_7084,N_7030);
or U7101 (N_7101,N_7071,N_7007);
and U7102 (N_7102,N_7091,N_7047);
xor U7103 (N_7103,N_7093,N_7050);
and U7104 (N_7104,N_7080,N_7060);
or U7105 (N_7105,N_7053,N_7096);
and U7106 (N_7106,N_7057,N_7098);
and U7107 (N_7107,N_7072,N_7032);
nand U7108 (N_7108,N_7068,N_7021);
or U7109 (N_7109,N_7027,N_7038);
xor U7110 (N_7110,N_7042,N_7069);
xor U7111 (N_7111,N_7065,N_7076);
or U7112 (N_7112,N_7097,N_7035);
nor U7113 (N_7113,N_7034,N_7070);
nand U7114 (N_7114,N_7003,N_7043);
nand U7115 (N_7115,N_7005,N_7024);
nand U7116 (N_7116,N_7085,N_7073);
or U7117 (N_7117,N_7082,N_7028);
and U7118 (N_7118,N_7090,N_7013);
and U7119 (N_7119,N_7011,N_7025);
nand U7120 (N_7120,N_7063,N_7015);
nand U7121 (N_7121,N_7040,N_7048);
and U7122 (N_7122,N_7055,N_7052);
xnor U7123 (N_7123,N_7058,N_7078);
or U7124 (N_7124,N_7014,N_7019);
and U7125 (N_7125,N_7089,N_7004);
nor U7126 (N_7126,N_7087,N_7092);
and U7127 (N_7127,N_7099,N_7031);
nand U7128 (N_7128,N_7039,N_7006);
nor U7129 (N_7129,N_7017,N_7051);
xnor U7130 (N_7130,N_7033,N_7020);
or U7131 (N_7131,N_7062,N_7079);
and U7132 (N_7132,N_7054,N_7023);
and U7133 (N_7133,N_7049,N_7064);
nand U7134 (N_7134,N_7041,N_7008);
xnor U7135 (N_7135,N_7010,N_7037);
nor U7136 (N_7136,N_7029,N_7095);
and U7137 (N_7137,N_7012,N_7061);
or U7138 (N_7138,N_7001,N_7086);
nand U7139 (N_7139,N_7067,N_7045);
nor U7140 (N_7140,N_7018,N_7075);
nor U7141 (N_7141,N_7066,N_7081);
or U7142 (N_7142,N_7044,N_7074);
nand U7143 (N_7143,N_7022,N_7059);
or U7144 (N_7144,N_7083,N_7077);
or U7145 (N_7145,N_7016,N_7056);
or U7146 (N_7146,N_7094,N_7036);
nor U7147 (N_7147,N_7000,N_7009);
and U7148 (N_7148,N_7026,N_7046);
nor U7149 (N_7149,N_7002,N_7088);
nand U7150 (N_7150,N_7040,N_7076);
nand U7151 (N_7151,N_7033,N_7023);
or U7152 (N_7152,N_7006,N_7026);
or U7153 (N_7153,N_7053,N_7006);
xor U7154 (N_7154,N_7045,N_7018);
and U7155 (N_7155,N_7082,N_7087);
nand U7156 (N_7156,N_7080,N_7040);
nand U7157 (N_7157,N_7068,N_7017);
and U7158 (N_7158,N_7071,N_7072);
nor U7159 (N_7159,N_7039,N_7083);
nand U7160 (N_7160,N_7074,N_7069);
nand U7161 (N_7161,N_7082,N_7065);
or U7162 (N_7162,N_7029,N_7000);
nor U7163 (N_7163,N_7023,N_7019);
xor U7164 (N_7164,N_7080,N_7095);
nand U7165 (N_7165,N_7016,N_7007);
nor U7166 (N_7166,N_7074,N_7008);
xnor U7167 (N_7167,N_7027,N_7088);
xor U7168 (N_7168,N_7063,N_7085);
nand U7169 (N_7169,N_7026,N_7019);
and U7170 (N_7170,N_7006,N_7024);
xor U7171 (N_7171,N_7038,N_7099);
and U7172 (N_7172,N_7046,N_7018);
nand U7173 (N_7173,N_7086,N_7049);
nand U7174 (N_7174,N_7020,N_7017);
nand U7175 (N_7175,N_7034,N_7073);
nand U7176 (N_7176,N_7069,N_7061);
xnor U7177 (N_7177,N_7022,N_7080);
and U7178 (N_7178,N_7067,N_7035);
or U7179 (N_7179,N_7074,N_7027);
xor U7180 (N_7180,N_7061,N_7083);
or U7181 (N_7181,N_7065,N_7057);
or U7182 (N_7182,N_7074,N_7038);
nor U7183 (N_7183,N_7004,N_7043);
nand U7184 (N_7184,N_7042,N_7082);
nand U7185 (N_7185,N_7095,N_7014);
or U7186 (N_7186,N_7069,N_7081);
nor U7187 (N_7187,N_7082,N_7024);
or U7188 (N_7188,N_7014,N_7068);
nand U7189 (N_7189,N_7080,N_7058);
nor U7190 (N_7190,N_7009,N_7031);
xnor U7191 (N_7191,N_7007,N_7027);
nand U7192 (N_7192,N_7079,N_7012);
and U7193 (N_7193,N_7010,N_7021);
nand U7194 (N_7194,N_7011,N_7015);
nor U7195 (N_7195,N_7090,N_7065);
and U7196 (N_7196,N_7088,N_7075);
and U7197 (N_7197,N_7079,N_7081);
nor U7198 (N_7198,N_7070,N_7077);
or U7199 (N_7199,N_7068,N_7072);
nor U7200 (N_7200,N_7192,N_7133);
nand U7201 (N_7201,N_7138,N_7112);
nand U7202 (N_7202,N_7139,N_7125);
nand U7203 (N_7203,N_7129,N_7175);
nor U7204 (N_7204,N_7187,N_7123);
xnor U7205 (N_7205,N_7135,N_7114);
nand U7206 (N_7206,N_7174,N_7109);
or U7207 (N_7207,N_7136,N_7182);
or U7208 (N_7208,N_7170,N_7195);
nand U7209 (N_7209,N_7106,N_7161);
xor U7210 (N_7210,N_7128,N_7189);
nand U7211 (N_7211,N_7190,N_7113);
nand U7212 (N_7212,N_7107,N_7122);
and U7213 (N_7213,N_7132,N_7126);
nand U7214 (N_7214,N_7159,N_7111);
nor U7215 (N_7215,N_7180,N_7169);
xor U7216 (N_7216,N_7194,N_7179);
nor U7217 (N_7217,N_7117,N_7102);
or U7218 (N_7218,N_7124,N_7100);
or U7219 (N_7219,N_7103,N_7141);
nor U7220 (N_7220,N_7149,N_7166);
nand U7221 (N_7221,N_7156,N_7154);
nand U7222 (N_7222,N_7137,N_7186);
xnor U7223 (N_7223,N_7171,N_7193);
nand U7224 (N_7224,N_7148,N_7188);
nor U7225 (N_7225,N_7116,N_7104);
and U7226 (N_7226,N_7120,N_7172);
and U7227 (N_7227,N_7198,N_7108);
nor U7228 (N_7228,N_7151,N_7176);
or U7229 (N_7229,N_7167,N_7155);
or U7230 (N_7230,N_7150,N_7119);
or U7231 (N_7231,N_7121,N_7157);
nor U7232 (N_7232,N_7164,N_7131);
nand U7233 (N_7233,N_7191,N_7134);
nor U7234 (N_7234,N_7196,N_7105);
and U7235 (N_7235,N_7145,N_7110);
xnor U7236 (N_7236,N_7178,N_7115);
or U7237 (N_7237,N_7165,N_7163);
nand U7238 (N_7238,N_7168,N_7143);
nor U7239 (N_7239,N_7184,N_7177);
xnor U7240 (N_7240,N_7147,N_7185);
xor U7241 (N_7241,N_7144,N_7130);
nor U7242 (N_7242,N_7127,N_7153);
nor U7243 (N_7243,N_7173,N_7183);
nor U7244 (N_7244,N_7140,N_7162);
nor U7245 (N_7245,N_7181,N_7199);
or U7246 (N_7246,N_7146,N_7160);
nand U7247 (N_7247,N_7101,N_7118);
and U7248 (N_7248,N_7152,N_7142);
xnor U7249 (N_7249,N_7197,N_7158);
or U7250 (N_7250,N_7112,N_7157);
or U7251 (N_7251,N_7177,N_7162);
nor U7252 (N_7252,N_7113,N_7108);
and U7253 (N_7253,N_7102,N_7127);
and U7254 (N_7254,N_7144,N_7102);
nand U7255 (N_7255,N_7182,N_7106);
xnor U7256 (N_7256,N_7116,N_7141);
xor U7257 (N_7257,N_7107,N_7136);
or U7258 (N_7258,N_7165,N_7161);
nand U7259 (N_7259,N_7171,N_7139);
xor U7260 (N_7260,N_7134,N_7198);
nor U7261 (N_7261,N_7112,N_7120);
nand U7262 (N_7262,N_7108,N_7127);
nand U7263 (N_7263,N_7127,N_7140);
or U7264 (N_7264,N_7130,N_7185);
xnor U7265 (N_7265,N_7185,N_7112);
nor U7266 (N_7266,N_7180,N_7165);
and U7267 (N_7267,N_7128,N_7165);
and U7268 (N_7268,N_7142,N_7189);
or U7269 (N_7269,N_7185,N_7174);
nor U7270 (N_7270,N_7198,N_7100);
nand U7271 (N_7271,N_7148,N_7165);
and U7272 (N_7272,N_7116,N_7156);
xnor U7273 (N_7273,N_7164,N_7191);
and U7274 (N_7274,N_7114,N_7111);
xnor U7275 (N_7275,N_7113,N_7156);
or U7276 (N_7276,N_7126,N_7112);
and U7277 (N_7277,N_7100,N_7161);
xor U7278 (N_7278,N_7167,N_7178);
or U7279 (N_7279,N_7182,N_7129);
xnor U7280 (N_7280,N_7124,N_7187);
nand U7281 (N_7281,N_7181,N_7187);
xor U7282 (N_7282,N_7173,N_7119);
nand U7283 (N_7283,N_7197,N_7130);
or U7284 (N_7284,N_7134,N_7151);
xnor U7285 (N_7285,N_7197,N_7178);
and U7286 (N_7286,N_7141,N_7113);
nor U7287 (N_7287,N_7140,N_7150);
nand U7288 (N_7288,N_7177,N_7146);
or U7289 (N_7289,N_7183,N_7112);
nor U7290 (N_7290,N_7103,N_7194);
and U7291 (N_7291,N_7163,N_7114);
and U7292 (N_7292,N_7165,N_7107);
or U7293 (N_7293,N_7149,N_7121);
nand U7294 (N_7294,N_7190,N_7171);
nand U7295 (N_7295,N_7147,N_7197);
nand U7296 (N_7296,N_7156,N_7149);
nand U7297 (N_7297,N_7147,N_7130);
or U7298 (N_7298,N_7125,N_7180);
xnor U7299 (N_7299,N_7177,N_7148);
xor U7300 (N_7300,N_7254,N_7208);
nand U7301 (N_7301,N_7211,N_7264);
or U7302 (N_7302,N_7242,N_7227);
nor U7303 (N_7303,N_7219,N_7236);
nor U7304 (N_7304,N_7213,N_7279);
xor U7305 (N_7305,N_7255,N_7241);
xor U7306 (N_7306,N_7200,N_7265);
nor U7307 (N_7307,N_7243,N_7276);
and U7308 (N_7308,N_7287,N_7280);
nor U7309 (N_7309,N_7269,N_7271);
nand U7310 (N_7310,N_7274,N_7253);
and U7311 (N_7311,N_7204,N_7205);
and U7312 (N_7312,N_7220,N_7250);
xnor U7313 (N_7313,N_7215,N_7296);
nand U7314 (N_7314,N_7247,N_7252);
or U7315 (N_7315,N_7240,N_7246);
nand U7316 (N_7316,N_7239,N_7284);
nand U7317 (N_7317,N_7294,N_7212);
nand U7318 (N_7318,N_7231,N_7299);
and U7319 (N_7319,N_7245,N_7267);
nand U7320 (N_7320,N_7295,N_7282);
nand U7321 (N_7321,N_7218,N_7275);
xnor U7322 (N_7322,N_7262,N_7257);
xor U7323 (N_7323,N_7206,N_7283);
and U7324 (N_7324,N_7266,N_7225);
and U7325 (N_7325,N_7288,N_7228);
or U7326 (N_7326,N_7260,N_7207);
or U7327 (N_7327,N_7285,N_7290);
and U7328 (N_7328,N_7298,N_7289);
and U7329 (N_7329,N_7256,N_7235);
or U7330 (N_7330,N_7217,N_7221);
xnor U7331 (N_7331,N_7201,N_7281);
nor U7332 (N_7332,N_7297,N_7238);
nor U7333 (N_7333,N_7293,N_7292);
nand U7334 (N_7334,N_7223,N_7291);
nor U7335 (N_7335,N_7229,N_7248);
nor U7336 (N_7336,N_7210,N_7232);
and U7337 (N_7337,N_7258,N_7286);
xor U7338 (N_7338,N_7234,N_7203);
or U7339 (N_7339,N_7273,N_7216);
nand U7340 (N_7340,N_7272,N_7222);
nand U7341 (N_7341,N_7209,N_7251);
nor U7342 (N_7342,N_7230,N_7226);
and U7343 (N_7343,N_7224,N_7263);
nand U7344 (N_7344,N_7270,N_7202);
nor U7345 (N_7345,N_7244,N_7277);
nand U7346 (N_7346,N_7278,N_7237);
or U7347 (N_7347,N_7259,N_7214);
nand U7348 (N_7348,N_7268,N_7249);
and U7349 (N_7349,N_7233,N_7261);
nand U7350 (N_7350,N_7272,N_7207);
and U7351 (N_7351,N_7274,N_7288);
nand U7352 (N_7352,N_7273,N_7293);
and U7353 (N_7353,N_7262,N_7280);
and U7354 (N_7354,N_7228,N_7289);
or U7355 (N_7355,N_7217,N_7213);
nand U7356 (N_7356,N_7243,N_7206);
or U7357 (N_7357,N_7290,N_7281);
or U7358 (N_7358,N_7256,N_7278);
nor U7359 (N_7359,N_7297,N_7208);
and U7360 (N_7360,N_7245,N_7230);
and U7361 (N_7361,N_7246,N_7297);
nand U7362 (N_7362,N_7262,N_7216);
xor U7363 (N_7363,N_7283,N_7209);
xnor U7364 (N_7364,N_7232,N_7264);
xnor U7365 (N_7365,N_7200,N_7292);
nand U7366 (N_7366,N_7239,N_7243);
nor U7367 (N_7367,N_7229,N_7250);
and U7368 (N_7368,N_7275,N_7276);
nor U7369 (N_7369,N_7258,N_7296);
and U7370 (N_7370,N_7255,N_7261);
nor U7371 (N_7371,N_7224,N_7249);
xor U7372 (N_7372,N_7202,N_7259);
nor U7373 (N_7373,N_7283,N_7256);
nand U7374 (N_7374,N_7208,N_7290);
nand U7375 (N_7375,N_7218,N_7214);
nand U7376 (N_7376,N_7236,N_7271);
xor U7377 (N_7377,N_7282,N_7298);
and U7378 (N_7378,N_7267,N_7203);
xnor U7379 (N_7379,N_7282,N_7284);
nand U7380 (N_7380,N_7268,N_7215);
and U7381 (N_7381,N_7261,N_7224);
nand U7382 (N_7382,N_7203,N_7241);
nor U7383 (N_7383,N_7245,N_7247);
nand U7384 (N_7384,N_7251,N_7244);
or U7385 (N_7385,N_7264,N_7209);
nand U7386 (N_7386,N_7295,N_7287);
or U7387 (N_7387,N_7277,N_7272);
xor U7388 (N_7388,N_7265,N_7205);
or U7389 (N_7389,N_7230,N_7288);
xor U7390 (N_7390,N_7202,N_7214);
xor U7391 (N_7391,N_7223,N_7240);
xor U7392 (N_7392,N_7262,N_7223);
nand U7393 (N_7393,N_7213,N_7262);
nand U7394 (N_7394,N_7200,N_7272);
and U7395 (N_7395,N_7208,N_7294);
or U7396 (N_7396,N_7269,N_7239);
and U7397 (N_7397,N_7207,N_7294);
xnor U7398 (N_7398,N_7288,N_7246);
nand U7399 (N_7399,N_7272,N_7227);
or U7400 (N_7400,N_7301,N_7350);
and U7401 (N_7401,N_7323,N_7374);
nor U7402 (N_7402,N_7351,N_7355);
xor U7403 (N_7403,N_7376,N_7315);
nor U7404 (N_7404,N_7302,N_7331);
nand U7405 (N_7405,N_7396,N_7391);
or U7406 (N_7406,N_7372,N_7380);
nand U7407 (N_7407,N_7347,N_7383);
xor U7408 (N_7408,N_7348,N_7335);
nor U7409 (N_7409,N_7381,N_7363);
nand U7410 (N_7410,N_7308,N_7319);
nor U7411 (N_7411,N_7398,N_7339);
xor U7412 (N_7412,N_7313,N_7316);
and U7413 (N_7413,N_7321,N_7300);
nand U7414 (N_7414,N_7314,N_7371);
or U7415 (N_7415,N_7375,N_7390);
and U7416 (N_7416,N_7329,N_7382);
and U7417 (N_7417,N_7387,N_7340);
or U7418 (N_7418,N_7362,N_7352);
and U7419 (N_7419,N_7395,N_7385);
or U7420 (N_7420,N_7369,N_7333);
or U7421 (N_7421,N_7310,N_7377);
and U7422 (N_7422,N_7334,N_7378);
nand U7423 (N_7423,N_7303,N_7397);
nor U7424 (N_7424,N_7327,N_7336);
or U7425 (N_7425,N_7305,N_7312);
and U7426 (N_7426,N_7367,N_7309);
and U7427 (N_7427,N_7370,N_7328);
or U7428 (N_7428,N_7317,N_7365);
or U7429 (N_7429,N_7359,N_7353);
or U7430 (N_7430,N_7325,N_7364);
or U7431 (N_7431,N_7337,N_7366);
nand U7432 (N_7432,N_7357,N_7356);
xnor U7433 (N_7433,N_7345,N_7384);
and U7434 (N_7434,N_7368,N_7326);
or U7435 (N_7435,N_7322,N_7306);
nor U7436 (N_7436,N_7392,N_7346);
xnor U7437 (N_7437,N_7307,N_7389);
xnor U7438 (N_7438,N_7304,N_7320);
nand U7439 (N_7439,N_7318,N_7349);
nand U7440 (N_7440,N_7386,N_7341);
and U7441 (N_7441,N_7342,N_7311);
and U7442 (N_7442,N_7393,N_7330);
and U7443 (N_7443,N_7373,N_7361);
or U7444 (N_7444,N_7379,N_7388);
nor U7445 (N_7445,N_7394,N_7338);
and U7446 (N_7446,N_7332,N_7343);
nor U7447 (N_7447,N_7344,N_7399);
xnor U7448 (N_7448,N_7358,N_7324);
nand U7449 (N_7449,N_7360,N_7354);
nand U7450 (N_7450,N_7358,N_7302);
or U7451 (N_7451,N_7309,N_7316);
nor U7452 (N_7452,N_7334,N_7392);
and U7453 (N_7453,N_7364,N_7367);
and U7454 (N_7454,N_7389,N_7339);
and U7455 (N_7455,N_7323,N_7383);
xor U7456 (N_7456,N_7376,N_7367);
nand U7457 (N_7457,N_7304,N_7363);
xor U7458 (N_7458,N_7315,N_7354);
nor U7459 (N_7459,N_7375,N_7305);
and U7460 (N_7460,N_7374,N_7385);
xnor U7461 (N_7461,N_7305,N_7324);
and U7462 (N_7462,N_7380,N_7389);
and U7463 (N_7463,N_7363,N_7331);
nand U7464 (N_7464,N_7397,N_7328);
nor U7465 (N_7465,N_7339,N_7347);
nor U7466 (N_7466,N_7385,N_7373);
xnor U7467 (N_7467,N_7373,N_7375);
nand U7468 (N_7468,N_7348,N_7317);
nand U7469 (N_7469,N_7328,N_7357);
nor U7470 (N_7470,N_7346,N_7364);
nor U7471 (N_7471,N_7311,N_7312);
nand U7472 (N_7472,N_7356,N_7378);
or U7473 (N_7473,N_7347,N_7378);
and U7474 (N_7474,N_7319,N_7392);
nand U7475 (N_7475,N_7300,N_7355);
nor U7476 (N_7476,N_7382,N_7359);
nor U7477 (N_7477,N_7307,N_7316);
or U7478 (N_7478,N_7356,N_7306);
nand U7479 (N_7479,N_7314,N_7367);
nand U7480 (N_7480,N_7323,N_7355);
or U7481 (N_7481,N_7371,N_7366);
xnor U7482 (N_7482,N_7304,N_7377);
nor U7483 (N_7483,N_7348,N_7371);
and U7484 (N_7484,N_7320,N_7365);
nor U7485 (N_7485,N_7312,N_7308);
nor U7486 (N_7486,N_7364,N_7311);
and U7487 (N_7487,N_7361,N_7335);
or U7488 (N_7488,N_7393,N_7363);
nand U7489 (N_7489,N_7312,N_7302);
xnor U7490 (N_7490,N_7363,N_7379);
xnor U7491 (N_7491,N_7365,N_7381);
nand U7492 (N_7492,N_7386,N_7343);
or U7493 (N_7493,N_7303,N_7323);
nor U7494 (N_7494,N_7376,N_7381);
nor U7495 (N_7495,N_7333,N_7392);
nand U7496 (N_7496,N_7354,N_7308);
and U7497 (N_7497,N_7317,N_7344);
and U7498 (N_7498,N_7311,N_7386);
and U7499 (N_7499,N_7391,N_7367);
and U7500 (N_7500,N_7491,N_7439);
xor U7501 (N_7501,N_7458,N_7450);
nor U7502 (N_7502,N_7484,N_7457);
nor U7503 (N_7503,N_7452,N_7485);
or U7504 (N_7504,N_7433,N_7462);
xor U7505 (N_7505,N_7414,N_7468);
xor U7506 (N_7506,N_7422,N_7463);
and U7507 (N_7507,N_7478,N_7460);
and U7508 (N_7508,N_7406,N_7493);
xor U7509 (N_7509,N_7486,N_7425);
and U7510 (N_7510,N_7446,N_7426);
and U7511 (N_7511,N_7476,N_7455);
or U7512 (N_7512,N_7488,N_7445);
nor U7513 (N_7513,N_7404,N_7411);
xor U7514 (N_7514,N_7444,N_7400);
nand U7515 (N_7515,N_7499,N_7447);
and U7516 (N_7516,N_7456,N_7441);
nor U7517 (N_7517,N_7496,N_7436);
or U7518 (N_7518,N_7492,N_7442);
and U7519 (N_7519,N_7453,N_7495);
or U7520 (N_7520,N_7483,N_7479);
xor U7521 (N_7521,N_7418,N_7465);
or U7522 (N_7522,N_7497,N_7469);
or U7523 (N_7523,N_7417,N_7423);
xor U7524 (N_7524,N_7430,N_7474);
xnor U7525 (N_7525,N_7494,N_7473);
nand U7526 (N_7526,N_7427,N_7403);
xor U7527 (N_7527,N_7466,N_7470);
or U7528 (N_7528,N_7489,N_7448);
or U7529 (N_7529,N_7419,N_7407);
nand U7530 (N_7530,N_7472,N_7482);
nor U7531 (N_7531,N_7421,N_7424);
nand U7532 (N_7532,N_7416,N_7487);
and U7533 (N_7533,N_7402,N_7428);
xor U7534 (N_7534,N_7408,N_7432);
nor U7535 (N_7535,N_7449,N_7401);
or U7536 (N_7536,N_7498,N_7459);
and U7537 (N_7537,N_7475,N_7415);
nor U7538 (N_7538,N_7440,N_7454);
and U7539 (N_7539,N_7477,N_7420);
or U7540 (N_7540,N_7435,N_7451);
nor U7541 (N_7541,N_7437,N_7410);
nor U7542 (N_7542,N_7405,N_7431);
nor U7543 (N_7543,N_7434,N_7467);
or U7544 (N_7544,N_7490,N_7429);
xor U7545 (N_7545,N_7413,N_7409);
nand U7546 (N_7546,N_7461,N_7471);
and U7547 (N_7547,N_7438,N_7480);
and U7548 (N_7548,N_7443,N_7481);
and U7549 (N_7549,N_7464,N_7412);
and U7550 (N_7550,N_7469,N_7419);
nand U7551 (N_7551,N_7464,N_7468);
nor U7552 (N_7552,N_7442,N_7432);
or U7553 (N_7553,N_7405,N_7456);
nor U7554 (N_7554,N_7464,N_7489);
nand U7555 (N_7555,N_7403,N_7471);
nor U7556 (N_7556,N_7435,N_7429);
xor U7557 (N_7557,N_7478,N_7466);
or U7558 (N_7558,N_7438,N_7402);
or U7559 (N_7559,N_7438,N_7442);
xor U7560 (N_7560,N_7491,N_7447);
and U7561 (N_7561,N_7434,N_7437);
nor U7562 (N_7562,N_7431,N_7448);
nand U7563 (N_7563,N_7498,N_7469);
xor U7564 (N_7564,N_7441,N_7478);
and U7565 (N_7565,N_7451,N_7412);
xnor U7566 (N_7566,N_7467,N_7411);
and U7567 (N_7567,N_7457,N_7424);
nand U7568 (N_7568,N_7416,N_7439);
nor U7569 (N_7569,N_7497,N_7473);
or U7570 (N_7570,N_7482,N_7421);
nand U7571 (N_7571,N_7474,N_7428);
nand U7572 (N_7572,N_7456,N_7447);
nor U7573 (N_7573,N_7402,N_7467);
nor U7574 (N_7574,N_7418,N_7429);
or U7575 (N_7575,N_7460,N_7405);
nand U7576 (N_7576,N_7463,N_7490);
and U7577 (N_7577,N_7467,N_7407);
nor U7578 (N_7578,N_7446,N_7443);
nor U7579 (N_7579,N_7464,N_7430);
or U7580 (N_7580,N_7494,N_7402);
nor U7581 (N_7581,N_7406,N_7460);
nor U7582 (N_7582,N_7401,N_7422);
xor U7583 (N_7583,N_7487,N_7403);
and U7584 (N_7584,N_7467,N_7460);
or U7585 (N_7585,N_7423,N_7414);
nand U7586 (N_7586,N_7425,N_7437);
xnor U7587 (N_7587,N_7462,N_7471);
nand U7588 (N_7588,N_7471,N_7478);
nand U7589 (N_7589,N_7401,N_7493);
or U7590 (N_7590,N_7432,N_7409);
nand U7591 (N_7591,N_7424,N_7407);
and U7592 (N_7592,N_7441,N_7403);
or U7593 (N_7593,N_7473,N_7443);
or U7594 (N_7594,N_7478,N_7444);
nor U7595 (N_7595,N_7475,N_7433);
or U7596 (N_7596,N_7448,N_7473);
nand U7597 (N_7597,N_7498,N_7453);
nor U7598 (N_7598,N_7456,N_7462);
and U7599 (N_7599,N_7414,N_7460);
and U7600 (N_7600,N_7533,N_7582);
or U7601 (N_7601,N_7585,N_7511);
nor U7602 (N_7602,N_7581,N_7532);
or U7603 (N_7603,N_7561,N_7593);
nor U7604 (N_7604,N_7525,N_7571);
or U7605 (N_7605,N_7507,N_7558);
and U7606 (N_7606,N_7543,N_7526);
nor U7607 (N_7607,N_7512,N_7565);
nand U7608 (N_7608,N_7550,N_7544);
or U7609 (N_7609,N_7503,N_7519);
nand U7610 (N_7610,N_7523,N_7570);
and U7611 (N_7611,N_7516,N_7520);
nor U7612 (N_7612,N_7549,N_7597);
nor U7613 (N_7613,N_7573,N_7552);
nor U7614 (N_7614,N_7510,N_7566);
nand U7615 (N_7615,N_7595,N_7502);
or U7616 (N_7616,N_7531,N_7513);
or U7617 (N_7617,N_7500,N_7509);
nand U7618 (N_7618,N_7546,N_7563);
and U7619 (N_7619,N_7564,N_7567);
nand U7620 (N_7620,N_7517,N_7578);
nand U7621 (N_7621,N_7522,N_7540);
nand U7622 (N_7622,N_7579,N_7588);
and U7623 (N_7623,N_7591,N_7534);
and U7624 (N_7624,N_7535,N_7548);
nor U7625 (N_7625,N_7530,N_7528);
xnor U7626 (N_7626,N_7592,N_7587);
nand U7627 (N_7627,N_7584,N_7537);
and U7628 (N_7628,N_7576,N_7508);
and U7629 (N_7629,N_7547,N_7521);
and U7630 (N_7630,N_7554,N_7504);
xor U7631 (N_7631,N_7557,N_7583);
and U7632 (N_7632,N_7524,N_7560);
nand U7633 (N_7633,N_7577,N_7539);
nor U7634 (N_7634,N_7586,N_7596);
and U7635 (N_7635,N_7551,N_7514);
xnor U7636 (N_7636,N_7594,N_7559);
or U7637 (N_7637,N_7574,N_7553);
nand U7638 (N_7638,N_7501,N_7556);
nor U7639 (N_7639,N_7555,N_7542);
or U7640 (N_7640,N_7505,N_7589);
and U7641 (N_7641,N_7562,N_7572);
and U7642 (N_7642,N_7598,N_7527);
or U7643 (N_7643,N_7529,N_7506);
nand U7644 (N_7644,N_7541,N_7599);
and U7645 (N_7645,N_7569,N_7568);
xor U7646 (N_7646,N_7580,N_7536);
nand U7647 (N_7647,N_7538,N_7575);
xnor U7648 (N_7648,N_7545,N_7590);
nand U7649 (N_7649,N_7518,N_7515);
nor U7650 (N_7650,N_7535,N_7571);
or U7651 (N_7651,N_7508,N_7510);
and U7652 (N_7652,N_7592,N_7541);
or U7653 (N_7653,N_7537,N_7501);
and U7654 (N_7654,N_7506,N_7569);
or U7655 (N_7655,N_7581,N_7554);
xor U7656 (N_7656,N_7591,N_7510);
xnor U7657 (N_7657,N_7586,N_7549);
or U7658 (N_7658,N_7545,N_7522);
nand U7659 (N_7659,N_7509,N_7555);
nand U7660 (N_7660,N_7506,N_7540);
nor U7661 (N_7661,N_7553,N_7547);
nand U7662 (N_7662,N_7561,N_7546);
xor U7663 (N_7663,N_7501,N_7578);
nor U7664 (N_7664,N_7539,N_7541);
and U7665 (N_7665,N_7504,N_7564);
or U7666 (N_7666,N_7557,N_7513);
nand U7667 (N_7667,N_7544,N_7594);
nand U7668 (N_7668,N_7516,N_7564);
nor U7669 (N_7669,N_7574,N_7589);
or U7670 (N_7670,N_7534,N_7545);
xor U7671 (N_7671,N_7525,N_7514);
nor U7672 (N_7672,N_7585,N_7509);
or U7673 (N_7673,N_7591,N_7519);
or U7674 (N_7674,N_7595,N_7598);
nand U7675 (N_7675,N_7589,N_7545);
xor U7676 (N_7676,N_7596,N_7567);
nand U7677 (N_7677,N_7505,N_7515);
and U7678 (N_7678,N_7585,N_7515);
or U7679 (N_7679,N_7593,N_7567);
and U7680 (N_7680,N_7557,N_7582);
xnor U7681 (N_7681,N_7586,N_7540);
and U7682 (N_7682,N_7562,N_7502);
xnor U7683 (N_7683,N_7526,N_7569);
xor U7684 (N_7684,N_7589,N_7538);
or U7685 (N_7685,N_7545,N_7549);
xor U7686 (N_7686,N_7553,N_7543);
or U7687 (N_7687,N_7526,N_7550);
nand U7688 (N_7688,N_7569,N_7515);
nand U7689 (N_7689,N_7541,N_7508);
or U7690 (N_7690,N_7534,N_7502);
nor U7691 (N_7691,N_7514,N_7561);
nand U7692 (N_7692,N_7590,N_7573);
xnor U7693 (N_7693,N_7595,N_7566);
nor U7694 (N_7694,N_7519,N_7572);
or U7695 (N_7695,N_7557,N_7569);
and U7696 (N_7696,N_7547,N_7574);
and U7697 (N_7697,N_7591,N_7529);
xor U7698 (N_7698,N_7572,N_7507);
nand U7699 (N_7699,N_7529,N_7526);
xnor U7700 (N_7700,N_7687,N_7601);
and U7701 (N_7701,N_7673,N_7678);
and U7702 (N_7702,N_7690,N_7681);
nor U7703 (N_7703,N_7609,N_7607);
xnor U7704 (N_7704,N_7668,N_7671);
nand U7705 (N_7705,N_7651,N_7691);
nand U7706 (N_7706,N_7646,N_7656);
nand U7707 (N_7707,N_7647,N_7659);
nor U7708 (N_7708,N_7652,N_7698);
and U7709 (N_7709,N_7641,N_7686);
xnor U7710 (N_7710,N_7664,N_7680);
nand U7711 (N_7711,N_7618,N_7674);
nor U7712 (N_7712,N_7670,N_7682);
nand U7713 (N_7713,N_7643,N_7653);
and U7714 (N_7714,N_7612,N_7662);
nand U7715 (N_7715,N_7634,N_7620);
nor U7716 (N_7716,N_7637,N_7611);
or U7717 (N_7717,N_7688,N_7639);
xor U7718 (N_7718,N_7636,N_7632);
xor U7719 (N_7719,N_7603,N_7615);
nand U7720 (N_7720,N_7638,N_7606);
or U7721 (N_7721,N_7622,N_7642);
nor U7722 (N_7722,N_7667,N_7616);
xnor U7723 (N_7723,N_7677,N_7627);
nand U7724 (N_7724,N_7679,N_7663);
nor U7725 (N_7725,N_7640,N_7655);
nand U7726 (N_7726,N_7649,N_7631);
nand U7727 (N_7727,N_7657,N_7619);
or U7728 (N_7728,N_7604,N_7605);
or U7729 (N_7729,N_7683,N_7602);
and U7730 (N_7730,N_7661,N_7676);
and U7731 (N_7731,N_7623,N_7675);
or U7732 (N_7732,N_7669,N_7648);
xor U7733 (N_7733,N_7692,N_7621);
and U7734 (N_7734,N_7624,N_7697);
xor U7735 (N_7735,N_7617,N_7654);
or U7736 (N_7736,N_7625,N_7608);
and U7737 (N_7737,N_7645,N_7630);
or U7738 (N_7738,N_7665,N_7626);
nor U7739 (N_7739,N_7658,N_7614);
nor U7740 (N_7740,N_7635,N_7600);
or U7741 (N_7741,N_7629,N_7628);
and U7742 (N_7742,N_7685,N_7666);
nor U7743 (N_7743,N_7644,N_7696);
nor U7744 (N_7744,N_7610,N_7660);
nand U7745 (N_7745,N_7694,N_7672);
or U7746 (N_7746,N_7650,N_7689);
nand U7747 (N_7747,N_7613,N_7695);
or U7748 (N_7748,N_7633,N_7684);
or U7749 (N_7749,N_7699,N_7693);
nor U7750 (N_7750,N_7643,N_7686);
nand U7751 (N_7751,N_7647,N_7673);
xnor U7752 (N_7752,N_7636,N_7644);
and U7753 (N_7753,N_7693,N_7652);
nand U7754 (N_7754,N_7672,N_7651);
and U7755 (N_7755,N_7652,N_7675);
nor U7756 (N_7756,N_7604,N_7695);
xnor U7757 (N_7757,N_7622,N_7658);
or U7758 (N_7758,N_7629,N_7665);
nor U7759 (N_7759,N_7641,N_7673);
xor U7760 (N_7760,N_7600,N_7671);
nor U7761 (N_7761,N_7638,N_7601);
or U7762 (N_7762,N_7662,N_7629);
and U7763 (N_7763,N_7645,N_7615);
or U7764 (N_7764,N_7696,N_7664);
nor U7765 (N_7765,N_7672,N_7646);
nand U7766 (N_7766,N_7657,N_7620);
nor U7767 (N_7767,N_7626,N_7604);
xnor U7768 (N_7768,N_7631,N_7670);
and U7769 (N_7769,N_7681,N_7696);
or U7770 (N_7770,N_7648,N_7627);
nand U7771 (N_7771,N_7616,N_7652);
xor U7772 (N_7772,N_7624,N_7636);
and U7773 (N_7773,N_7629,N_7694);
and U7774 (N_7774,N_7636,N_7615);
nand U7775 (N_7775,N_7667,N_7614);
and U7776 (N_7776,N_7616,N_7647);
or U7777 (N_7777,N_7622,N_7675);
nand U7778 (N_7778,N_7642,N_7614);
and U7779 (N_7779,N_7670,N_7664);
nand U7780 (N_7780,N_7606,N_7619);
nand U7781 (N_7781,N_7660,N_7637);
and U7782 (N_7782,N_7614,N_7676);
or U7783 (N_7783,N_7686,N_7674);
xnor U7784 (N_7784,N_7624,N_7665);
and U7785 (N_7785,N_7632,N_7627);
or U7786 (N_7786,N_7626,N_7660);
nor U7787 (N_7787,N_7626,N_7631);
or U7788 (N_7788,N_7610,N_7665);
nand U7789 (N_7789,N_7684,N_7646);
or U7790 (N_7790,N_7603,N_7688);
xor U7791 (N_7791,N_7688,N_7658);
xnor U7792 (N_7792,N_7604,N_7694);
nand U7793 (N_7793,N_7637,N_7644);
nor U7794 (N_7794,N_7645,N_7609);
xor U7795 (N_7795,N_7600,N_7664);
or U7796 (N_7796,N_7686,N_7687);
nor U7797 (N_7797,N_7610,N_7638);
nor U7798 (N_7798,N_7634,N_7610);
nand U7799 (N_7799,N_7657,N_7647);
nor U7800 (N_7800,N_7737,N_7786);
nand U7801 (N_7801,N_7727,N_7718);
nor U7802 (N_7802,N_7798,N_7736);
and U7803 (N_7803,N_7754,N_7759);
xnor U7804 (N_7804,N_7717,N_7799);
or U7805 (N_7805,N_7733,N_7794);
xnor U7806 (N_7806,N_7795,N_7729);
nand U7807 (N_7807,N_7761,N_7793);
or U7808 (N_7808,N_7721,N_7735);
or U7809 (N_7809,N_7738,N_7712);
xor U7810 (N_7810,N_7762,N_7748);
or U7811 (N_7811,N_7775,N_7760);
nor U7812 (N_7812,N_7705,N_7790);
nand U7813 (N_7813,N_7700,N_7785);
and U7814 (N_7814,N_7773,N_7777);
xnor U7815 (N_7815,N_7708,N_7728);
and U7816 (N_7816,N_7703,N_7742);
and U7817 (N_7817,N_7766,N_7743);
or U7818 (N_7818,N_7778,N_7715);
nand U7819 (N_7819,N_7725,N_7780);
nor U7820 (N_7820,N_7765,N_7769);
or U7821 (N_7821,N_7797,N_7749);
nand U7822 (N_7822,N_7767,N_7764);
and U7823 (N_7823,N_7789,N_7731);
and U7824 (N_7824,N_7787,N_7763);
and U7825 (N_7825,N_7746,N_7758);
xor U7826 (N_7826,N_7755,N_7788);
and U7827 (N_7827,N_7770,N_7740);
nand U7828 (N_7828,N_7796,N_7732);
or U7829 (N_7829,N_7713,N_7719);
nor U7830 (N_7830,N_7706,N_7783);
nand U7831 (N_7831,N_7702,N_7753);
and U7832 (N_7832,N_7784,N_7776);
xnor U7833 (N_7833,N_7709,N_7774);
nor U7834 (N_7834,N_7714,N_7739);
nor U7835 (N_7835,N_7722,N_7704);
and U7836 (N_7836,N_7716,N_7747);
xor U7837 (N_7837,N_7791,N_7781);
and U7838 (N_7838,N_7710,N_7792);
and U7839 (N_7839,N_7744,N_7745);
nand U7840 (N_7840,N_7720,N_7711);
or U7841 (N_7841,N_7734,N_7779);
xor U7842 (N_7842,N_7768,N_7723);
or U7843 (N_7843,N_7771,N_7752);
nand U7844 (N_7844,N_7772,N_7724);
and U7845 (N_7845,N_7707,N_7757);
nand U7846 (N_7846,N_7756,N_7751);
or U7847 (N_7847,N_7726,N_7782);
nor U7848 (N_7848,N_7750,N_7730);
xor U7849 (N_7849,N_7741,N_7701);
and U7850 (N_7850,N_7718,N_7748);
xor U7851 (N_7851,N_7722,N_7700);
nand U7852 (N_7852,N_7768,N_7788);
nor U7853 (N_7853,N_7783,N_7772);
and U7854 (N_7854,N_7781,N_7774);
nand U7855 (N_7855,N_7730,N_7736);
and U7856 (N_7856,N_7793,N_7797);
and U7857 (N_7857,N_7730,N_7788);
xnor U7858 (N_7858,N_7753,N_7740);
and U7859 (N_7859,N_7731,N_7759);
nor U7860 (N_7860,N_7777,N_7794);
nor U7861 (N_7861,N_7705,N_7769);
and U7862 (N_7862,N_7772,N_7720);
nand U7863 (N_7863,N_7733,N_7700);
nor U7864 (N_7864,N_7761,N_7730);
nor U7865 (N_7865,N_7722,N_7760);
or U7866 (N_7866,N_7776,N_7714);
nor U7867 (N_7867,N_7732,N_7740);
nand U7868 (N_7868,N_7766,N_7752);
nand U7869 (N_7869,N_7796,N_7792);
nor U7870 (N_7870,N_7779,N_7797);
nand U7871 (N_7871,N_7749,N_7730);
and U7872 (N_7872,N_7797,N_7765);
xor U7873 (N_7873,N_7704,N_7757);
nor U7874 (N_7874,N_7754,N_7797);
xnor U7875 (N_7875,N_7745,N_7720);
and U7876 (N_7876,N_7733,N_7766);
nor U7877 (N_7877,N_7780,N_7773);
or U7878 (N_7878,N_7753,N_7723);
nor U7879 (N_7879,N_7772,N_7719);
nor U7880 (N_7880,N_7712,N_7762);
nor U7881 (N_7881,N_7781,N_7727);
or U7882 (N_7882,N_7750,N_7712);
nor U7883 (N_7883,N_7796,N_7790);
nor U7884 (N_7884,N_7797,N_7729);
nor U7885 (N_7885,N_7772,N_7705);
xnor U7886 (N_7886,N_7766,N_7793);
or U7887 (N_7887,N_7768,N_7783);
xnor U7888 (N_7888,N_7760,N_7761);
nand U7889 (N_7889,N_7754,N_7783);
or U7890 (N_7890,N_7769,N_7748);
or U7891 (N_7891,N_7717,N_7731);
nand U7892 (N_7892,N_7772,N_7730);
or U7893 (N_7893,N_7793,N_7784);
nor U7894 (N_7894,N_7747,N_7705);
nor U7895 (N_7895,N_7785,N_7798);
nor U7896 (N_7896,N_7720,N_7727);
and U7897 (N_7897,N_7791,N_7785);
xor U7898 (N_7898,N_7761,N_7701);
or U7899 (N_7899,N_7751,N_7777);
and U7900 (N_7900,N_7864,N_7889);
nand U7901 (N_7901,N_7828,N_7833);
nand U7902 (N_7902,N_7810,N_7884);
nor U7903 (N_7903,N_7862,N_7869);
xnor U7904 (N_7904,N_7826,N_7841);
and U7905 (N_7905,N_7888,N_7866);
nor U7906 (N_7906,N_7835,N_7806);
and U7907 (N_7907,N_7830,N_7894);
nor U7908 (N_7908,N_7844,N_7876);
or U7909 (N_7909,N_7870,N_7867);
xor U7910 (N_7910,N_7813,N_7858);
xnor U7911 (N_7911,N_7851,N_7850);
xnor U7912 (N_7912,N_7831,N_7892);
and U7913 (N_7913,N_7857,N_7834);
nand U7914 (N_7914,N_7803,N_7837);
or U7915 (N_7915,N_7800,N_7887);
nor U7916 (N_7916,N_7821,N_7861);
nand U7917 (N_7917,N_7839,N_7883);
nor U7918 (N_7918,N_7874,N_7815);
nand U7919 (N_7919,N_7875,N_7873);
nand U7920 (N_7920,N_7898,N_7896);
or U7921 (N_7921,N_7849,N_7880);
or U7922 (N_7922,N_7863,N_7824);
and U7923 (N_7923,N_7853,N_7865);
and U7924 (N_7924,N_7878,N_7817);
nand U7925 (N_7925,N_7871,N_7872);
nor U7926 (N_7926,N_7802,N_7882);
and U7927 (N_7927,N_7805,N_7809);
or U7928 (N_7928,N_7801,N_7842);
xnor U7929 (N_7929,N_7845,N_7856);
or U7930 (N_7930,N_7804,N_7860);
and U7931 (N_7931,N_7825,N_7893);
nand U7932 (N_7932,N_7895,N_7832);
nand U7933 (N_7933,N_7897,N_7885);
nor U7934 (N_7934,N_7812,N_7846);
or U7935 (N_7935,N_7822,N_7848);
nand U7936 (N_7936,N_7840,N_7899);
and U7937 (N_7937,N_7881,N_7854);
nand U7938 (N_7938,N_7819,N_7836);
nor U7939 (N_7939,N_7843,N_7808);
and U7940 (N_7940,N_7811,N_7829);
nand U7941 (N_7941,N_7891,N_7852);
or U7942 (N_7942,N_7877,N_7886);
nor U7943 (N_7943,N_7859,N_7816);
nor U7944 (N_7944,N_7890,N_7847);
and U7945 (N_7945,N_7818,N_7814);
and U7946 (N_7946,N_7820,N_7879);
and U7947 (N_7947,N_7823,N_7807);
nand U7948 (N_7948,N_7868,N_7855);
xnor U7949 (N_7949,N_7827,N_7838);
and U7950 (N_7950,N_7866,N_7805);
or U7951 (N_7951,N_7854,N_7806);
or U7952 (N_7952,N_7868,N_7866);
xor U7953 (N_7953,N_7899,N_7835);
xnor U7954 (N_7954,N_7887,N_7842);
xnor U7955 (N_7955,N_7810,N_7868);
or U7956 (N_7956,N_7847,N_7894);
nand U7957 (N_7957,N_7852,N_7860);
or U7958 (N_7958,N_7842,N_7877);
and U7959 (N_7959,N_7873,N_7883);
and U7960 (N_7960,N_7876,N_7858);
xnor U7961 (N_7961,N_7843,N_7883);
xnor U7962 (N_7962,N_7801,N_7885);
or U7963 (N_7963,N_7865,N_7841);
and U7964 (N_7964,N_7808,N_7852);
and U7965 (N_7965,N_7813,N_7849);
xnor U7966 (N_7966,N_7808,N_7856);
nor U7967 (N_7967,N_7860,N_7849);
nor U7968 (N_7968,N_7870,N_7871);
nand U7969 (N_7969,N_7871,N_7844);
nor U7970 (N_7970,N_7857,N_7888);
and U7971 (N_7971,N_7811,N_7860);
nand U7972 (N_7972,N_7871,N_7847);
nor U7973 (N_7973,N_7861,N_7828);
or U7974 (N_7974,N_7844,N_7843);
xor U7975 (N_7975,N_7857,N_7867);
xnor U7976 (N_7976,N_7866,N_7875);
nand U7977 (N_7977,N_7832,N_7867);
xor U7978 (N_7978,N_7882,N_7815);
xnor U7979 (N_7979,N_7825,N_7854);
and U7980 (N_7980,N_7828,N_7864);
or U7981 (N_7981,N_7804,N_7814);
and U7982 (N_7982,N_7802,N_7826);
and U7983 (N_7983,N_7857,N_7861);
or U7984 (N_7984,N_7870,N_7842);
or U7985 (N_7985,N_7826,N_7878);
xor U7986 (N_7986,N_7897,N_7837);
xnor U7987 (N_7987,N_7879,N_7859);
xor U7988 (N_7988,N_7866,N_7865);
nand U7989 (N_7989,N_7863,N_7831);
xor U7990 (N_7990,N_7859,N_7845);
nor U7991 (N_7991,N_7867,N_7843);
nor U7992 (N_7992,N_7830,N_7860);
nor U7993 (N_7993,N_7831,N_7814);
or U7994 (N_7994,N_7842,N_7807);
or U7995 (N_7995,N_7846,N_7821);
xnor U7996 (N_7996,N_7895,N_7824);
nand U7997 (N_7997,N_7871,N_7873);
xnor U7998 (N_7998,N_7852,N_7828);
and U7999 (N_7999,N_7886,N_7821);
xor U8000 (N_8000,N_7952,N_7968);
nor U8001 (N_8001,N_7941,N_7918);
nand U8002 (N_8002,N_7922,N_7917);
nor U8003 (N_8003,N_7940,N_7919);
xnor U8004 (N_8004,N_7951,N_7955);
nor U8005 (N_8005,N_7975,N_7921);
xnor U8006 (N_8006,N_7993,N_7936);
xnor U8007 (N_8007,N_7932,N_7973);
nand U8008 (N_8008,N_7907,N_7915);
nor U8009 (N_8009,N_7946,N_7999);
nand U8010 (N_8010,N_7930,N_7981);
or U8011 (N_8011,N_7995,N_7929);
and U8012 (N_8012,N_7954,N_7984);
and U8013 (N_8013,N_7970,N_7923);
xnor U8014 (N_8014,N_7909,N_7961);
and U8015 (N_8015,N_7964,N_7926);
nand U8016 (N_8016,N_7953,N_7938);
or U8017 (N_8017,N_7945,N_7966);
nor U8018 (N_8018,N_7979,N_7957);
nor U8019 (N_8019,N_7972,N_7959);
nor U8020 (N_8020,N_7904,N_7914);
nor U8021 (N_8021,N_7965,N_7960);
and U8022 (N_8022,N_7991,N_7990);
nand U8023 (N_8023,N_7937,N_7971);
nor U8024 (N_8024,N_7974,N_7916);
nor U8025 (N_8025,N_7982,N_7977);
and U8026 (N_8026,N_7901,N_7978);
or U8027 (N_8027,N_7996,N_7943);
or U8028 (N_8028,N_7949,N_7950);
xor U8029 (N_8029,N_7902,N_7933);
or U8030 (N_8030,N_7927,N_7958);
and U8031 (N_8031,N_7903,N_7994);
nor U8032 (N_8032,N_7913,N_7985);
and U8033 (N_8033,N_7942,N_7910);
nor U8034 (N_8034,N_7905,N_7956);
xor U8035 (N_8035,N_7948,N_7988);
xnor U8036 (N_8036,N_7983,N_7925);
nor U8037 (N_8037,N_7906,N_7911);
or U8038 (N_8038,N_7992,N_7986);
nor U8039 (N_8039,N_7997,N_7998);
nor U8040 (N_8040,N_7931,N_7920);
xor U8041 (N_8041,N_7967,N_7939);
nand U8042 (N_8042,N_7980,N_7924);
or U8043 (N_8043,N_7944,N_7908);
nor U8044 (N_8044,N_7900,N_7969);
xnor U8045 (N_8045,N_7962,N_7976);
or U8046 (N_8046,N_7935,N_7934);
or U8047 (N_8047,N_7947,N_7912);
and U8048 (N_8048,N_7928,N_7989);
and U8049 (N_8049,N_7987,N_7963);
nor U8050 (N_8050,N_7966,N_7929);
nand U8051 (N_8051,N_7946,N_7974);
and U8052 (N_8052,N_7912,N_7916);
xor U8053 (N_8053,N_7922,N_7973);
xnor U8054 (N_8054,N_7911,N_7982);
nor U8055 (N_8055,N_7916,N_7946);
nand U8056 (N_8056,N_7909,N_7916);
nand U8057 (N_8057,N_7950,N_7957);
and U8058 (N_8058,N_7991,N_7903);
and U8059 (N_8059,N_7934,N_7985);
nand U8060 (N_8060,N_7952,N_7935);
xnor U8061 (N_8061,N_7992,N_7989);
or U8062 (N_8062,N_7934,N_7923);
and U8063 (N_8063,N_7905,N_7918);
xor U8064 (N_8064,N_7957,N_7926);
xnor U8065 (N_8065,N_7966,N_7959);
and U8066 (N_8066,N_7900,N_7917);
nand U8067 (N_8067,N_7982,N_7983);
or U8068 (N_8068,N_7976,N_7975);
nor U8069 (N_8069,N_7934,N_7942);
or U8070 (N_8070,N_7997,N_7958);
nand U8071 (N_8071,N_7952,N_7957);
and U8072 (N_8072,N_7997,N_7966);
nand U8073 (N_8073,N_7979,N_7932);
nor U8074 (N_8074,N_7941,N_7933);
nand U8075 (N_8075,N_7941,N_7970);
nor U8076 (N_8076,N_7913,N_7992);
nor U8077 (N_8077,N_7930,N_7931);
and U8078 (N_8078,N_7950,N_7970);
or U8079 (N_8079,N_7997,N_7946);
nor U8080 (N_8080,N_7922,N_7956);
xor U8081 (N_8081,N_7946,N_7931);
and U8082 (N_8082,N_7912,N_7962);
xnor U8083 (N_8083,N_7974,N_7950);
or U8084 (N_8084,N_7951,N_7908);
or U8085 (N_8085,N_7946,N_7993);
nor U8086 (N_8086,N_7935,N_7982);
nor U8087 (N_8087,N_7948,N_7998);
nand U8088 (N_8088,N_7962,N_7918);
or U8089 (N_8089,N_7941,N_7973);
or U8090 (N_8090,N_7935,N_7990);
or U8091 (N_8091,N_7969,N_7919);
nand U8092 (N_8092,N_7959,N_7957);
xor U8093 (N_8093,N_7975,N_7971);
and U8094 (N_8094,N_7993,N_7920);
nand U8095 (N_8095,N_7924,N_7926);
xnor U8096 (N_8096,N_7991,N_7914);
and U8097 (N_8097,N_7959,N_7964);
nor U8098 (N_8098,N_7929,N_7992);
nor U8099 (N_8099,N_7990,N_7995);
and U8100 (N_8100,N_8095,N_8044);
nor U8101 (N_8101,N_8078,N_8002);
or U8102 (N_8102,N_8080,N_8068);
and U8103 (N_8103,N_8086,N_8008);
nand U8104 (N_8104,N_8003,N_8041);
nor U8105 (N_8105,N_8094,N_8035);
nor U8106 (N_8106,N_8097,N_8067);
nand U8107 (N_8107,N_8069,N_8022);
and U8108 (N_8108,N_8064,N_8016);
nor U8109 (N_8109,N_8063,N_8027);
xnor U8110 (N_8110,N_8015,N_8024);
and U8111 (N_8111,N_8023,N_8053);
nor U8112 (N_8112,N_8004,N_8032);
and U8113 (N_8113,N_8087,N_8089);
and U8114 (N_8114,N_8037,N_8059);
xor U8115 (N_8115,N_8062,N_8017);
xor U8116 (N_8116,N_8021,N_8051);
or U8117 (N_8117,N_8034,N_8077);
nor U8118 (N_8118,N_8036,N_8043);
nand U8119 (N_8119,N_8075,N_8061);
or U8120 (N_8120,N_8005,N_8093);
xnor U8121 (N_8121,N_8085,N_8091);
nor U8122 (N_8122,N_8014,N_8030);
xor U8123 (N_8123,N_8048,N_8049);
nor U8124 (N_8124,N_8056,N_8052);
and U8125 (N_8125,N_8009,N_8012);
xor U8126 (N_8126,N_8007,N_8001);
xor U8127 (N_8127,N_8065,N_8082);
or U8128 (N_8128,N_8029,N_8047);
nand U8129 (N_8129,N_8031,N_8019);
nor U8130 (N_8130,N_8045,N_8033);
or U8131 (N_8131,N_8028,N_8073);
and U8132 (N_8132,N_8079,N_8020);
xnor U8133 (N_8133,N_8088,N_8096);
xor U8134 (N_8134,N_8070,N_8025);
or U8135 (N_8135,N_8084,N_8092);
xnor U8136 (N_8136,N_8010,N_8060);
nor U8137 (N_8137,N_8011,N_8076);
and U8138 (N_8138,N_8098,N_8000);
nor U8139 (N_8139,N_8006,N_8057);
nand U8140 (N_8140,N_8026,N_8083);
nand U8141 (N_8141,N_8039,N_8071);
xnor U8142 (N_8142,N_8081,N_8040);
nand U8143 (N_8143,N_8072,N_8018);
or U8144 (N_8144,N_8046,N_8074);
xor U8145 (N_8145,N_8050,N_8099);
or U8146 (N_8146,N_8013,N_8058);
and U8147 (N_8147,N_8066,N_8090);
nand U8148 (N_8148,N_8055,N_8054);
or U8149 (N_8149,N_8042,N_8038);
or U8150 (N_8150,N_8000,N_8083);
and U8151 (N_8151,N_8023,N_8015);
and U8152 (N_8152,N_8036,N_8042);
and U8153 (N_8153,N_8081,N_8031);
nor U8154 (N_8154,N_8032,N_8005);
or U8155 (N_8155,N_8016,N_8072);
or U8156 (N_8156,N_8031,N_8013);
xor U8157 (N_8157,N_8044,N_8060);
and U8158 (N_8158,N_8025,N_8048);
nand U8159 (N_8159,N_8003,N_8030);
nor U8160 (N_8160,N_8082,N_8005);
or U8161 (N_8161,N_8091,N_8075);
and U8162 (N_8162,N_8040,N_8072);
xnor U8163 (N_8163,N_8057,N_8003);
or U8164 (N_8164,N_8064,N_8069);
nor U8165 (N_8165,N_8034,N_8047);
nor U8166 (N_8166,N_8083,N_8071);
nand U8167 (N_8167,N_8050,N_8079);
or U8168 (N_8168,N_8010,N_8041);
and U8169 (N_8169,N_8016,N_8074);
nor U8170 (N_8170,N_8012,N_8056);
or U8171 (N_8171,N_8072,N_8083);
and U8172 (N_8172,N_8051,N_8007);
and U8173 (N_8173,N_8065,N_8000);
nand U8174 (N_8174,N_8040,N_8083);
nand U8175 (N_8175,N_8047,N_8033);
nand U8176 (N_8176,N_8050,N_8015);
or U8177 (N_8177,N_8022,N_8075);
nand U8178 (N_8178,N_8031,N_8009);
xnor U8179 (N_8179,N_8062,N_8008);
or U8180 (N_8180,N_8093,N_8014);
or U8181 (N_8181,N_8073,N_8067);
nor U8182 (N_8182,N_8020,N_8058);
xor U8183 (N_8183,N_8078,N_8042);
and U8184 (N_8184,N_8016,N_8040);
or U8185 (N_8185,N_8041,N_8075);
and U8186 (N_8186,N_8025,N_8023);
and U8187 (N_8187,N_8057,N_8021);
xor U8188 (N_8188,N_8035,N_8053);
and U8189 (N_8189,N_8003,N_8031);
or U8190 (N_8190,N_8085,N_8076);
and U8191 (N_8191,N_8063,N_8038);
nand U8192 (N_8192,N_8095,N_8052);
nor U8193 (N_8193,N_8059,N_8051);
nand U8194 (N_8194,N_8000,N_8006);
xor U8195 (N_8195,N_8054,N_8084);
nand U8196 (N_8196,N_8064,N_8020);
and U8197 (N_8197,N_8010,N_8093);
and U8198 (N_8198,N_8088,N_8070);
nor U8199 (N_8199,N_8000,N_8074);
xnor U8200 (N_8200,N_8156,N_8172);
and U8201 (N_8201,N_8146,N_8121);
or U8202 (N_8202,N_8168,N_8179);
or U8203 (N_8203,N_8135,N_8176);
nand U8204 (N_8204,N_8151,N_8161);
xnor U8205 (N_8205,N_8171,N_8196);
and U8206 (N_8206,N_8189,N_8180);
nand U8207 (N_8207,N_8192,N_8134);
nand U8208 (N_8208,N_8108,N_8109);
or U8209 (N_8209,N_8154,N_8152);
xor U8210 (N_8210,N_8184,N_8194);
nand U8211 (N_8211,N_8131,N_8102);
and U8212 (N_8212,N_8186,N_8193);
nor U8213 (N_8213,N_8169,N_8130);
nor U8214 (N_8214,N_8181,N_8188);
xnor U8215 (N_8215,N_8199,N_8110);
or U8216 (N_8216,N_8111,N_8187);
nor U8217 (N_8217,N_8117,N_8128);
xor U8218 (N_8218,N_8133,N_8162);
nand U8219 (N_8219,N_8198,N_8174);
or U8220 (N_8220,N_8126,N_8153);
nor U8221 (N_8221,N_8182,N_8101);
and U8222 (N_8222,N_8167,N_8159);
xnor U8223 (N_8223,N_8140,N_8175);
xor U8224 (N_8224,N_8118,N_8112);
nor U8225 (N_8225,N_8104,N_8183);
nand U8226 (N_8226,N_8141,N_8165);
nor U8227 (N_8227,N_8157,N_8164);
and U8228 (N_8228,N_8163,N_8139);
nand U8229 (N_8229,N_8143,N_8103);
xor U8230 (N_8230,N_8177,N_8113);
nand U8231 (N_8231,N_8116,N_8166);
nor U8232 (N_8232,N_8124,N_8107);
and U8233 (N_8233,N_8123,N_8195);
xnor U8234 (N_8234,N_8160,N_8190);
nor U8235 (N_8235,N_8149,N_8142);
nand U8236 (N_8236,N_8106,N_8125);
nor U8237 (N_8237,N_8145,N_8105);
nand U8238 (N_8238,N_8136,N_8197);
and U8239 (N_8239,N_8129,N_8120);
nand U8240 (N_8240,N_8127,N_8178);
nand U8241 (N_8241,N_8137,N_8100);
nand U8242 (N_8242,N_8185,N_8147);
xor U8243 (N_8243,N_8170,N_8122);
or U8244 (N_8244,N_8158,N_8191);
and U8245 (N_8245,N_8173,N_8148);
xnor U8246 (N_8246,N_8155,N_8119);
nand U8247 (N_8247,N_8150,N_8132);
or U8248 (N_8248,N_8138,N_8144);
nand U8249 (N_8249,N_8115,N_8114);
or U8250 (N_8250,N_8114,N_8154);
nand U8251 (N_8251,N_8132,N_8105);
and U8252 (N_8252,N_8155,N_8152);
nor U8253 (N_8253,N_8168,N_8152);
and U8254 (N_8254,N_8118,N_8190);
xor U8255 (N_8255,N_8156,N_8153);
nand U8256 (N_8256,N_8174,N_8191);
nor U8257 (N_8257,N_8121,N_8116);
nand U8258 (N_8258,N_8195,N_8171);
nand U8259 (N_8259,N_8114,N_8145);
nand U8260 (N_8260,N_8153,N_8189);
and U8261 (N_8261,N_8162,N_8187);
nand U8262 (N_8262,N_8171,N_8138);
nor U8263 (N_8263,N_8191,N_8175);
or U8264 (N_8264,N_8133,N_8119);
xor U8265 (N_8265,N_8150,N_8102);
or U8266 (N_8266,N_8190,N_8104);
and U8267 (N_8267,N_8193,N_8184);
nor U8268 (N_8268,N_8133,N_8172);
and U8269 (N_8269,N_8184,N_8158);
nor U8270 (N_8270,N_8186,N_8110);
or U8271 (N_8271,N_8179,N_8153);
nor U8272 (N_8272,N_8125,N_8169);
nor U8273 (N_8273,N_8116,N_8185);
and U8274 (N_8274,N_8167,N_8158);
or U8275 (N_8275,N_8184,N_8157);
or U8276 (N_8276,N_8109,N_8193);
nand U8277 (N_8277,N_8110,N_8166);
xnor U8278 (N_8278,N_8101,N_8129);
xnor U8279 (N_8279,N_8139,N_8171);
and U8280 (N_8280,N_8182,N_8150);
or U8281 (N_8281,N_8168,N_8135);
nor U8282 (N_8282,N_8125,N_8130);
or U8283 (N_8283,N_8172,N_8157);
nand U8284 (N_8284,N_8183,N_8133);
nor U8285 (N_8285,N_8148,N_8159);
nand U8286 (N_8286,N_8172,N_8192);
nand U8287 (N_8287,N_8192,N_8100);
and U8288 (N_8288,N_8114,N_8186);
and U8289 (N_8289,N_8105,N_8174);
nor U8290 (N_8290,N_8104,N_8133);
and U8291 (N_8291,N_8199,N_8160);
nand U8292 (N_8292,N_8116,N_8180);
and U8293 (N_8293,N_8133,N_8171);
nor U8294 (N_8294,N_8101,N_8159);
xnor U8295 (N_8295,N_8111,N_8110);
xnor U8296 (N_8296,N_8105,N_8108);
and U8297 (N_8297,N_8130,N_8192);
xor U8298 (N_8298,N_8141,N_8175);
nand U8299 (N_8299,N_8119,N_8165);
or U8300 (N_8300,N_8237,N_8233);
or U8301 (N_8301,N_8217,N_8297);
nand U8302 (N_8302,N_8220,N_8223);
nand U8303 (N_8303,N_8242,N_8203);
or U8304 (N_8304,N_8290,N_8244);
nand U8305 (N_8305,N_8208,N_8224);
or U8306 (N_8306,N_8238,N_8270);
xnor U8307 (N_8307,N_8235,N_8205);
and U8308 (N_8308,N_8286,N_8200);
and U8309 (N_8309,N_8225,N_8213);
or U8310 (N_8310,N_8264,N_8262);
xnor U8311 (N_8311,N_8261,N_8280);
and U8312 (N_8312,N_8253,N_8201);
nor U8313 (N_8313,N_8230,N_8231);
or U8314 (N_8314,N_8239,N_8245);
xor U8315 (N_8315,N_8275,N_8243);
or U8316 (N_8316,N_8295,N_8278);
and U8317 (N_8317,N_8226,N_8218);
nand U8318 (N_8318,N_8271,N_8246);
nor U8319 (N_8319,N_8296,N_8299);
xor U8320 (N_8320,N_8294,N_8206);
and U8321 (N_8321,N_8209,N_8283);
and U8322 (N_8322,N_8202,N_8268);
and U8323 (N_8323,N_8236,N_8255);
or U8324 (N_8324,N_8256,N_8211);
and U8325 (N_8325,N_8274,N_8219);
xor U8326 (N_8326,N_8227,N_8287);
or U8327 (N_8327,N_8252,N_8291);
nand U8328 (N_8328,N_8298,N_8241);
nand U8329 (N_8329,N_8207,N_8234);
nand U8330 (N_8330,N_8288,N_8282);
or U8331 (N_8331,N_8221,N_8279);
nand U8332 (N_8332,N_8272,N_8266);
or U8333 (N_8333,N_8240,N_8258);
and U8334 (N_8334,N_8222,N_8285);
or U8335 (N_8335,N_8284,N_8263);
and U8336 (N_8336,N_8277,N_8232);
or U8337 (N_8337,N_8292,N_8216);
xnor U8338 (N_8338,N_8254,N_8289);
or U8339 (N_8339,N_8257,N_8260);
nor U8340 (N_8340,N_8250,N_8249);
nand U8341 (N_8341,N_8247,N_8281);
and U8342 (N_8342,N_8293,N_8214);
or U8343 (N_8343,N_8228,N_8229);
nand U8344 (N_8344,N_8210,N_8265);
or U8345 (N_8345,N_8204,N_8267);
xnor U8346 (N_8346,N_8215,N_8276);
xnor U8347 (N_8347,N_8269,N_8251);
xnor U8348 (N_8348,N_8259,N_8248);
or U8349 (N_8349,N_8212,N_8273);
nand U8350 (N_8350,N_8291,N_8247);
xnor U8351 (N_8351,N_8286,N_8245);
xnor U8352 (N_8352,N_8284,N_8212);
nand U8353 (N_8353,N_8262,N_8285);
and U8354 (N_8354,N_8220,N_8263);
xnor U8355 (N_8355,N_8201,N_8205);
and U8356 (N_8356,N_8212,N_8202);
nor U8357 (N_8357,N_8221,N_8285);
or U8358 (N_8358,N_8276,N_8212);
nor U8359 (N_8359,N_8282,N_8204);
xnor U8360 (N_8360,N_8292,N_8242);
and U8361 (N_8361,N_8249,N_8281);
nand U8362 (N_8362,N_8233,N_8223);
and U8363 (N_8363,N_8211,N_8209);
nor U8364 (N_8364,N_8266,N_8281);
nand U8365 (N_8365,N_8289,N_8241);
xor U8366 (N_8366,N_8284,N_8216);
nor U8367 (N_8367,N_8276,N_8244);
nand U8368 (N_8368,N_8205,N_8258);
nor U8369 (N_8369,N_8235,N_8239);
nor U8370 (N_8370,N_8265,N_8233);
nor U8371 (N_8371,N_8292,N_8255);
and U8372 (N_8372,N_8215,N_8246);
and U8373 (N_8373,N_8288,N_8233);
nand U8374 (N_8374,N_8278,N_8227);
nand U8375 (N_8375,N_8277,N_8250);
nand U8376 (N_8376,N_8216,N_8219);
nand U8377 (N_8377,N_8286,N_8223);
nand U8378 (N_8378,N_8217,N_8201);
nor U8379 (N_8379,N_8200,N_8278);
and U8380 (N_8380,N_8200,N_8237);
or U8381 (N_8381,N_8236,N_8211);
nand U8382 (N_8382,N_8289,N_8265);
nand U8383 (N_8383,N_8285,N_8213);
nand U8384 (N_8384,N_8248,N_8299);
xnor U8385 (N_8385,N_8238,N_8231);
xor U8386 (N_8386,N_8201,N_8285);
nand U8387 (N_8387,N_8280,N_8247);
nand U8388 (N_8388,N_8207,N_8236);
nand U8389 (N_8389,N_8234,N_8264);
xor U8390 (N_8390,N_8267,N_8257);
nor U8391 (N_8391,N_8217,N_8232);
and U8392 (N_8392,N_8271,N_8267);
xnor U8393 (N_8393,N_8232,N_8238);
nand U8394 (N_8394,N_8212,N_8245);
xor U8395 (N_8395,N_8264,N_8240);
nor U8396 (N_8396,N_8247,N_8226);
nor U8397 (N_8397,N_8205,N_8239);
or U8398 (N_8398,N_8215,N_8288);
and U8399 (N_8399,N_8231,N_8285);
nand U8400 (N_8400,N_8382,N_8303);
or U8401 (N_8401,N_8386,N_8347);
or U8402 (N_8402,N_8327,N_8341);
or U8403 (N_8403,N_8322,N_8392);
nor U8404 (N_8404,N_8393,N_8329);
nand U8405 (N_8405,N_8311,N_8333);
and U8406 (N_8406,N_8371,N_8312);
nand U8407 (N_8407,N_8361,N_8375);
nor U8408 (N_8408,N_8318,N_8346);
xnor U8409 (N_8409,N_8326,N_8328);
or U8410 (N_8410,N_8359,N_8300);
xnor U8411 (N_8411,N_8350,N_8352);
nor U8412 (N_8412,N_8301,N_8332);
and U8413 (N_8413,N_8377,N_8306);
nand U8414 (N_8414,N_8321,N_8372);
or U8415 (N_8415,N_8395,N_8317);
xor U8416 (N_8416,N_8309,N_8367);
xnor U8417 (N_8417,N_8307,N_8384);
xor U8418 (N_8418,N_8310,N_8340);
xor U8419 (N_8419,N_8353,N_8302);
nand U8420 (N_8420,N_8345,N_8348);
nor U8421 (N_8421,N_8381,N_8315);
nand U8422 (N_8422,N_8373,N_8383);
or U8423 (N_8423,N_8308,N_8385);
nand U8424 (N_8424,N_8396,N_8399);
and U8425 (N_8425,N_8380,N_8370);
or U8426 (N_8426,N_8360,N_8314);
nor U8427 (N_8427,N_8368,N_8320);
nor U8428 (N_8428,N_8313,N_8351);
and U8429 (N_8429,N_8358,N_8379);
and U8430 (N_8430,N_8388,N_8394);
nand U8431 (N_8431,N_8305,N_8319);
nand U8432 (N_8432,N_8391,N_8374);
xnor U8433 (N_8433,N_8363,N_8356);
xnor U8434 (N_8434,N_8366,N_8316);
nand U8435 (N_8435,N_8397,N_8338);
xnor U8436 (N_8436,N_8325,N_8398);
or U8437 (N_8437,N_8365,N_8344);
and U8438 (N_8438,N_8335,N_8343);
nand U8439 (N_8439,N_8337,N_8357);
or U8440 (N_8440,N_8349,N_8369);
nand U8441 (N_8441,N_8336,N_8362);
xnor U8442 (N_8442,N_8304,N_8339);
and U8443 (N_8443,N_8342,N_8323);
xor U8444 (N_8444,N_8330,N_8355);
and U8445 (N_8445,N_8354,N_8378);
nand U8446 (N_8446,N_8364,N_8376);
and U8447 (N_8447,N_8331,N_8387);
xnor U8448 (N_8448,N_8334,N_8324);
nand U8449 (N_8449,N_8390,N_8389);
and U8450 (N_8450,N_8374,N_8367);
nor U8451 (N_8451,N_8324,N_8381);
or U8452 (N_8452,N_8390,N_8322);
or U8453 (N_8453,N_8354,N_8382);
or U8454 (N_8454,N_8380,N_8333);
or U8455 (N_8455,N_8374,N_8380);
nor U8456 (N_8456,N_8321,N_8354);
xnor U8457 (N_8457,N_8398,N_8384);
and U8458 (N_8458,N_8394,N_8389);
nor U8459 (N_8459,N_8338,N_8391);
or U8460 (N_8460,N_8315,N_8393);
nor U8461 (N_8461,N_8374,N_8356);
xnor U8462 (N_8462,N_8355,N_8366);
and U8463 (N_8463,N_8310,N_8388);
xnor U8464 (N_8464,N_8317,N_8349);
and U8465 (N_8465,N_8325,N_8349);
nor U8466 (N_8466,N_8396,N_8384);
and U8467 (N_8467,N_8349,N_8366);
nor U8468 (N_8468,N_8311,N_8345);
nor U8469 (N_8469,N_8344,N_8351);
or U8470 (N_8470,N_8340,N_8391);
nor U8471 (N_8471,N_8306,N_8327);
nor U8472 (N_8472,N_8384,N_8319);
nand U8473 (N_8473,N_8368,N_8339);
nor U8474 (N_8474,N_8365,N_8317);
and U8475 (N_8475,N_8360,N_8367);
nor U8476 (N_8476,N_8331,N_8351);
or U8477 (N_8477,N_8330,N_8352);
and U8478 (N_8478,N_8390,N_8336);
nor U8479 (N_8479,N_8343,N_8370);
and U8480 (N_8480,N_8338,N_8310);
and U8481 (N_8481,N_8329,N_8352);
nand U8482 (N_8482,N_8390,N_8381);
nor U8483 (N_8483,N_8305,N_8355);
or U8484 (N_8484,N_8368,N_8315);
nor U8485 (N_8485,N_8320,N_8398);
xnor U8486 (N_8486,N_8351,N_8372);
nand U8487 (N_8487,N_8307,N_8378);
xor U8488 (N_8488,N_8366,N_8362);
nand U8489 (N_8489,N_8385,N_8353);
xnor U8490 (N_8490,N_8359,N_8306);
nand U8491 (N_8491,N_8394,N_8355);
nor U8492 (N_8492,N_8399,N_8310);
nand U8493 (N_8493,N_8355,N_8391);
nor U8494 (N_8494,N_8300,N_8304);
or U8495 (N_8495,N_8366,N_8385);
nand U8496 (N_8496,N_8302,N_8307);
nand U8497 (N_8497,N_8363,N_8328);
or U8498 (N_8498,N_8335,N_8331);
xor U8499 (N_8499,N_8308,N_8357);
nor U8500 (N_8500,N_8490,N_8416);
nor U8501 (N_8501,N_8432,N_8443);
xnor U8502 (N_8502,N_8447,N_8483);
or U8503 (N_8503,N_8491,N_8473);
xnor U8504 (N_8504,N_8472,N_8444);
nor U8505 (N_8505,N_8462,N_8409);
and U8506 (N_8506,N_8486,N_8478);
and U8507 (N_8507,N_8487,N_8411);
nand U8508 (N_8508,N_8435,N_8434);
nand U8509 (N_8509,N_8440,N_8496);
nand U8510 (N_8510,N_8467,N_8420);
nand U8511 (N_8511,N_8461,N_8446);
or U8512 (N_8512,N_8419,N_8463);
nand U8513 (N_8513,N_8406,N_8415);
or U8514 (N_8514,N_8404,N_8497);
xor U8515 (N_8515,N_8466,N_8481);
nor U8516 (N_8516,N_8430,N_8427);
xor U8517 (N_8517,N_8412,N_8422);
or U8518 (N_8518,N_8499,N_8421);
or U8519 (N_8519,N_8408,N_8417);
nand U8520 (N_8520,N_8464,N_8450);
or U8521 (N_8521,N_8477,N_8445);
and U8522 (N_8522,N_8448,N_8468);
and U8523 (N_8523,N_8433,N_8480);
nor U8524 (N_8524,N_8413,N_8405);
nor U8525 (N_8525,N_8470,N_8469);
nor U8526 (N_8526,N_8451,N_8459);
or U8527 (N_8527,N_8476,N_8424);
and U8528 (N_8528,N_8400,N_8475);
nor U8529 (N_8529,N_8493,N_8489);
nor U8530 (N_8530,N_8453,N_8403);
xor U8531 (N_8531,N_8438,N_8402);
and U8532 (N_8532,N_8455,N_8439);
nand U8533 (N_8533,N_8401,N_8441);
or U8534 (N_8534,N_8485,N_8425);
and U8535 (N_8535,N_8431,N_8407);
and U8536 (N_8536,N_8423,N_8498);
nor U8537 (N_8537,N_8479,N_8471);
nand U8538 (N_8538,N_8437,N_8488);
xor U8539 (N_8539,N_8457,N_8442);
and U8540 (N_8540,N_8494,N_8449);
and U8541 (N_8541,N_8458,N_8482);
nand U8542 (N_8542,N_8484,N_8495);
or U8543 (N_8543,N_8429,N_8492);
and U8544 (N_8544,N_8452,N_8428);
and U8545 (N_8545,N_8460,N_8410);
xor U8546 (N_8546,N_8418,N_8465);
xor U8547 (N_8547,N_8456,N_8436);
nor U8548 (N_8548,N_8474,N_8454);
nand U8549 (N_8549,N_8414,N_8426);
or U8550 (N_8550,N_8482,N_8463);
or U8551 (N_8551,N_8449,N_8458);
nor U8552 (N_8552,N_8440,N_8404);
and U8553 (N_8553,N_8494,N_8439);
or U8554 (N_8554,N_8412,N_8458);
and U8555 (N_8555,N_8473,N_8449);
or U8556 (N_8556,N_8427,N_8401);
xor U8557 (N_8557,N_8476,N_8417);
nand U8558 (N_8558,N_8405,N_8469);
or U8559 (N_8559,N_8478,N_8455);
and U8560 (N_8560,N_8468,N_8490);
xor U8561 (N_8561,N_8454,N_8436);
and U8562 (N_8562,N_8495,N_8475);
or U8563 (N_8563,N_8493,N_8481);
xor U8564 (N_8564,N_8477,N_8466);
xnor U8565 (N_8565,N_8411,N_8465);
nand U8566 (N_8566,N_8461,N_8448);
xor U8567 (N_8567,N_8420,N_8425);
and U8568 (N_8568,N_8402,N_8479);
nor U8569 (N_8569,N_8458,N_8453);
xnor U8570 (N_8570,N_8453,N_8464);
nor U8571 (N_8571,N_8447,N_8445);
xor U8572 (N_8572,N_8466,N_8419);
and U8573 (N_8573,N_8495,N_8479);
nor U8574 (N_8574,N_8471,N_8421);
or U8575 (N_8575,N_8489,N_8488);
or U8576 (N_8576,N_8496,N_8428);
nor U8577 (N_8577,N_8445,N_8452);
or U8578 (N_8578,N_8476,N_8498);
xnor U8579 (N_8579,N_8439,N_8452);
xnor U8580 (N_8580,N_8444,N_8471);
and U8581 (N_8581,N_8404,N_8491);
nor U8582 (N_8582,N_8414,N_8466);
or U8583 (N_8583,N_8457,N_8421);
or U8584 (N_8584,N_8451,N_8410);
xnor U8585 (N_8585,N_8446,N_8451);
or U8586 (N_8586,N_8426,N_8434);
or U8587 (N_8587,N_8498,N_8458);
and U8588 (N_8588,N_8407,N_8451);
and U8589 (N_8589,N_8411,N_8484);
or U8590 (N_8590,N_8457,N_8461);
nor U8591 (N_8591,N_8441,N_8410);
xnor U8592 (N_8592,N_8417,N_8433);
or U8593 (N_8593,N_8477,N_8417);
and U8594 (N_8594,N_8470,N_8448);
nand U8595 (N_8595,N_8476,N_8453);
xnor U8596 (N_8596,N_8470,N_8435);
and U8597 (N_8597,N_8401,N_8421);
nand U8598 (N_8598,N_8412,N_8429);
and U8599 (N_8599,N_8475,N_8438);
nor U8600 (N_8600,N_8502,N_8586);
nand U8601 (N_8601,N_8564,N_8595);
nor U8602 (N_8602,N_8545,N_8528);
and U8603 (N_8603,N_8517,N_8525);
and U8604 (N_8604,N_8506,N_8533);
nor U8605 (N_8605,N_8509,N_8562);
xor U8606 (N_8606,N_8513,N_8596);
or U8607 (N_8607,N_8561,N_8578);
xnor U8608 (N_8608,N_8585,N_8527);
nand U8609 (N_8609,N_8551,N_8598);
and U8610 (N_8610,N_8531,N_8558);
nor U8611 (N_8611,N_8589,N_8504);
xnor U8612 (N_8612,N_8535,N_8550);
and U8613 (N_8613,N_8519,N_8510);
and U8614 (N_8614,N_8554,N_8581);
nor U8615 (N_8615,N_8524,N_8518);
or U8616 (N_8616,N_8583,N_8505);
nor U8617 (N_8617,N_8571,N_8594);
xnor U8618 (N_8618,N_8568,N_8591);
or U8619 (N_8619,N_8534,N_8542);
nand U8620 (N_8620,N_8567,N_8529);
nand U8621 (N_8621,N_8597,N_8569);
or U8622 (N_8622,N_8566,N_8556);
xor U8623 (N_8623,N_8526,N_8584);
or U8624 (N_8624,N_8557,N_8570);
or U8625 (N_8625,N_8532,N_8559);
xnor U8626 (N_8626,N_8563,N_8541);
nor U8627 (N_8627,N_8579,N_8514);
and U8628 (N_8628,N_8565,N_8580);
xor U8629 (N_8629,N_8590,N_8592);
and U8630 (N_8630,N_8512,N_8549);
nor U8631 (N_8631,N_8588,N_8523);
xor U8632 (N_8632,N_8544,N_8515);
or U8633 (N_8633,N_8501,N_8560);
or U8634 (N_8634,N_8511,N_8508);
xor U8635 (N_8635,N_8548,N_8547);
or U8636 (N_8636,N_8516,N_8507);
or U8637 (N_8637,N_8500,N_8573);
or U8638 (N_8638,N_8582,N_8593);
or U8639 (N_8639,N_8599,N_8546);
or U8640 (N_8640,N_8538,N_8540);
and U8641 (N_8641,N_8577,N_8503);
nor U8642 (N_8642,N_8553,N_8520);
xnor U8643 (N_8643,N_8575,N_8539);
or U8644 (N_8644,N_8522,N_8574);
xor U8645 (N_8645,N_8530,N_8572);
or U8646 (N_8646,N_8555,N_8521);
xnor U8647 (N_8647,N_8576,N_8552);
and U8648 (N_8648,N_8543,N_8587);
xor U8649 (N_8649,N_8536,N_8537);
or U8650 (N_8650,N_8593,N_8552);
xnor U8651 (N_8651,N_8527,N_8529);
or U8652 (N_8652,N_8599,N_8583);
nand U8653 (N_8653,N_8520,N_8549);
and U8654 (N_8654,N_8536,N_8565);
and U8655 (N_8655,N_8591,N_8592);
or U8656 (N_8656,N_8573,N_8595);
nor U8657 (N_8657,N_8580,N_8548);
nand U8658 (N_8658,N_8543,N_8523);
nor U8659 (N_8659,N_8589,N_8593);
and U8660 (N_8660,N_8566,N_8522);
or U8661 (N_8661,N_8547,N_8522);
xor U8662 (N_8662,N_8524,N_8530);
xor U8663 (N_8663,N_8591,N_8513);
or U8664 (N_8664,N_8527,N_8558);
nand U8665 (N_8665,N_8510,N_8518);
nand U8666 (N_8666,N_8518,N_8534);
nand U8667 (N_8667,N_8565,N_8543);
nor U8668 (N_8668,N_8555,N_8507);
nor U8669 (N_8669,N_8560,N_8509);
and U8670 (N_8670,N_8510,N_8500);
nand U8671 (N_8671,N_8574,N_8590);
nor U8672 (N_8672,N_8526,N_8502);
xnor U8673 (N_8673,N_8537,N_8509);
nor U8674 (N_8674,N_8553,N_8568);
or U8675 (N_8675,N_8542,N_8570);
nand U8676 (N_8676,N_8506,N_8559);
nand U8677 (N_8677,N_8557,N_8534);
or U8678 (N_8678,N_8590,N_8576);
and U8679 (N_8679,N_8519,N_8591);
or U8680 (N_8680,N_8505,N_8511);
nand U8681 (N_8681,N_8587,N_8504);
nor U8682 (N_8682,N_8591,N_8564);
nand U8683 (N_8683,N_8571,N_8508);
or U8684 (N_8684,N_8545,N_8552);
and U8685 (N_8685,N_8568,N_8599);
nand U8686 (N_8686,N_8520,N_8506);
or U8687 (N_8687,N_8575,N_8595);
xnor U8688 (N_8688,N_8583,N_8537);
nand U8689 (N_8689,N_8514,N_8553);
nor U8690 (N_8690,N_8548,N_8551);
nand U8691 (N_8691,N_8529,N_8589);
nand U8692 (N_8692,N_8538,N_8594);
nor U8693 (N_8693,N_8530,N_8567);
and U8694 (N_8694,N_8575,N_8554);
or U8695 (N_8695,N_8562,N_8540);
and U8696 (N_8696,N_8517,N_8569);
nor U8697 (N_8697,N_8591,N_8521);
and U8698 (N_8698,N_8544,N_8516);
nand U8699 (N_8699,N_8536,N_8563);
and U8700 (N_8700,N_8624,N_8658);
nand U8701 (N_8701,N_8605,N_8687);
and U8702 (N_8702,N_8643,N_8669);
nor U8703 (N_8703,N_8609,N_8626);
nor U8704 (N_8704,N_8646,N_8617);
or U8705 (N_8705,N_8613,N_8610);
xor U8706 (N_8706,N_8695,N_8684);
and U8707 (N_8707,N_8686,N_8673);
nand U8708 (N_8708,N_8660,N_8619);
xnor U8709 (N_8709,N_8670,N_8645);
nand U8710 (N_8710,N_8635,N_8638);
or U8711 (N_8711,N_8625,N_8672);
nand U8712 (N_8712,N_8693,N_8655);
and U8713 (N_8713,N_8677,N_8696);
nor U8714 (N_8714,N_8620,N_8689);
xor U8715 (N_8715,N_8606,N_8639);
nand U8716 (N_8716,N_8649,N_8678);
or U8717 (N_8717,N_8634,N_8698);
and U8718 (N_8718,N_8682,N_8691);
xnor U8719 (N_8719,N_8623,N_8621);
or U8720 (N_8720,N_8602,N_8603);
or U8721 (N_8721,N_8601,N_8627);
and U8722 (N_8722,N_8600,N_8663);
nand U8723 (N_8723,N_8661,N_8612);
or U8724 (N_8724,N_8607,N_8630);
or U8725 (N_8725,N_8688,N_8671);
xor U8726 (N_8726,N_8641,N_8642);
nand U8727 (N_8727,N_8640,N_8685);
and U8728 (N_8728,N_8608,N_8679);
and U8729 (N_8729,N_8675,N_8694);
nand U8730 (N_8730,N_8680,N_8656);
or U8731 (N_8731,N_8631,N_8659);
xor U8732 (N_8732,N_8628,N_8653);
xor U8733 (N_8733,N_8681,N_8690);
xor U8734 (N_8734,N_8647,N_8637);
nor U8735 (N_8735,N_8654,N_8644);
nor U8736 (N_8736,N_8676,N_8611);
or U8737 (N_8737,N_8651,N_8662);
nand U8738 (N_8738,N_8666,N_8692);
or U8739 (N_8739,N_8697,N_8668);
and U8740 (N_8740,N_8683,N_8650);
or U8741 (N_8741,N_8604,N_8664);
xor U8742 (N_8742,N_8618,N_8648);
nand U8743 (N_8743,N_8699,N_8614);
or U8744 (N_8744,N_8667,N_8657);
xor U8745 (N_8745,N_8674,N_8632);
nand U8746 (N_8746,N_8622,N_8629);
or U8747 (N_8747,N_8665,N_8616);
or U8748 (N_8748,N_8615,N_8636);
nor U8749 (N_8749,N_8633,N_8652);
nand U8750 (N_8750,N_8638,N_8620);
nor U8751 (N_8751,N_8658,N_8611);
nand U8752 (N_8752,N_8640,N_8680);
and U8753 (N_8753,N_8656,N_8664);
nor U8754 (N_8754,N_8612,N_8644);
nor U8755 (N_8755,N_8612,N_8658);
nand U8756 (N_8756,N_8699,N_8637);
nor U8757 (N_8757,N_8641,N_8622);
or U8758 (N_8758,N_8677,N_8698);
xor U8759 (N_8759,N_8649,N_8690);
nand U8760 (N_8760,N_8695,N_8670);
and U8761 (N_8761,N_8689,N_8601);
xor U8762 (N_8762,N_8686,N_8643);
nand U8763 (N_8763,N_8665,N_8621);
nor U8764 (N_8764,N_8634,N_8606);
nor U8765 (N_8765,N_8689,N_8642);
and U8766 (N_8766,N_8620,N_8670);
and U8767 (N_8767,N_8675,N_8649);
nand U8768 (N_8768,N_8602,N_8664);
or U8769 (N_8769,N_8687,N_8610);
and U8770 (N_8770,N_8621,N_8629);
or U8771 (N_8771,N_8651,N_8611);
xor U8772 (N_8772,N_8638,N_8649);
or U8773 (N_8773,N_8650,N_8652);
nand U8774 (N_8774,N_8618,N_8610);
and U8775 (N_8775,N_8677,N_8647);
and U8776 (N_8776,N_8685,N_8681);
or U8777 (N_8777,N_8665,N_8692);
nand U8778 (N_8778,N_8666,N_8606);
nand U8779 (N_8779,N_8676,N_8682);
nand U8780 (N_8780,N_8639,N_8690);
or U8781 (N_8781,N_8649,N_8619);
nor U8782 (N_8782,N_8607,N_8671);
nand U8783 (N_8783,N_8619,N_8632);
nor U8784 (N_8784,N_8639,N_8685);
xor U8785 (N_8785,N_8608,N_8641);
xnor U8786 (N_8786,N_8605,N_8662);
nand U8787 (N_8787,N_8640,N_8659);
nor U8788 (N_8788,N_8684,N_8617);
xor U8789 (N_8789,N_8683,N_8696);
and U8790 (N_8790,N_8617,N_8639);
nor U8791 (N_8791,N_8608,N_8627);
nand U8792 (N_8792,N_8675,N_8665);
nand U8793 (N_8793,N_8638,N_8680);
xor U8794 (N_8794,N_8607,N_8650);
nor U8795 (N_8795,N_8622,N_8659);
nor U8796 (N_8796,N_8600,N_8673);
and U8797 (N_8797,N_8603,N_8619);
and U8798 (N_8798,N_8673,N_8627);
nand U8799 (N_8799,N_8685,N_8688);
nand U8800 (N_8800,N_8714,N_8745);
or U8801 (N_8801,N_8704,N_8749);
and U8802 (N_8802,N_8770,N_8732);
or U8803 (N_8803,N_8727,N_8701);
nand U8804 (N_8804,N_8739,N_8796);
nand U8805 (N_8805,N_8791,N_8767);
nor U8806 (N_8806,N_8740,N_8711);
or U8807 (N_8807,N_8724,N_8799);
or U8808 (N_8808,N_8720,N_8762);
and U8809 (N_8809,N_8725,N_8754);
nor U8810 (N_8810,N_8798,N_8723);
and U8811 (N_8811,N_8776,N_8763);
or U8812 (N_8812,N_8783,N_8730);
nand U8813 (N_8813,N_8717,N_8794);
or U8814 (N_8814,N_8786,N_8702);
or U8815 (N_8815,N_8769,N_8765);
nand U8816 (N_8816,N_8775,N_8759);
nor U8817 (N_8817,N_8751,N_8774);
xnor U8818 (N_8818,N_8710,N_8744);
nand U8819 (N_8819,N_8729,N_8721);
nor U8820 (N_8820,N_8758,N_8736);
or U8821 (N_8821,N_8748,N_8703);
and U8822 (N_8822,N_8764,N_8785);
nor U8823 (N_8823,N_8750,N_8789);
or U8824 (N_8824,N_8733,N_8792);
or U8825 (N_8825,N_8706,N_8793);
xnor U8826 (N_8826,N_8722,N_8777);
or U8827 (N_8827,N_8779,N_8780);
and U8828 (N_8828,N_8766,N_8708);
or U8829 (N_8829,N_8738,N_8757);
xor U8830 (N_8830,N_8797,N_8715);
or U8831 (N_8831,N_8705,N_8747);
or U8832 (N_8832,N_8795,N_8728);
and U8833 (N_8833,N_8719,N_8700);
or U8834 (N_8834,N_8746,N_8741);
xnor U8835 (N_8835,N_8753,N_8772);
xnor U8836 (N_8836,N_8755,N_8773);
xor U8837 (N_8837,N_8761,N_8718);
nor U8838 (N_8838,N_8742,N_8788);
xor U8839 (N_8839,N_8707,N_8713);
xnor U8840 (N_8840,N_8760,N_8709);
and U8841 (N_8841,N_8716,N_8734);
and U8842 (N_8842,N_8756,N_8726);
nand U8843 (N_8843,N_8781,N_8768);
nor U8844 (N_8844,N_8737,N_8787);
or U8845 (N_8845,N_8743,N_8771);
nand U8846 (N_8846,N_8731,N_8784);
xnor U8847 (N_8847,N_8752,N_8712);
and U8848 (N_8848,N_8790,N_8782);
nor U8849 (N_8849,N_8735,N_8778);
xor U8850 (N_8850,N_8788,N_8735);
xor U8851 (N_8851,N_8716,N_8782);
and U8852 (N_8852,N_8739,N_8794);
nand U8853 (N_8853,N_8743,N_8784);
nor U8854 (N_8854,N_8702,N_8782);
nand U8855 (N_8855,N_8780,N_8744);
or U8856 (N_8856,N_8784,N_8778);
xnor U8857 (N_8857,N_8773,N_8711);
xor U8858 (N_8858,N_8717,N_8725);
xor U8859 (N_8859,N_8762,N_8711);
or U8860 (N_8860,N_8781,N_8745);
and U8861 (N_8861,N_8771,N_8730);
xor U8862 (N_8862,N_8749,N_8732);
nand U8863 (N_8863,N_8780,N_8717);
and U8864 (N_8864,N_8747,N_8732);
nor U8865 (N_8865,N_8732,N_8714);
nand U8866 (N_8866,N_8723,N_8729);
nand U8867 (N_8867,N_8785,N_8741);
and U8868 (N_8868,N_8740,N_8774);
nand U8869 (N_8869,N_8731,N_8735);
or U8870 (N_8870,N_8791,N_8732);
nand U8871 (N_8871,N_8726,N_8732);
or U8872 (N_8872,N_8751,N_8779);
xnor U8873 (N_8873,N_8742,N_8795);
xor U8874 (N_8874,N_8767,N_8747);
and U8875 (N_8875,N_8763,N_8772);
xor U8876 (N_8876,N_8788,N_8702);
xor U8877 (N_8877,N_8709,N_8763);
and U8878 (N_8878,N_8728,N_8736);
nor U8879 (N_8879,N_8742,N_8768);
xnor U8880 (N_8880,N_8760,N_8729);
and U8881 (N_8881,N_8775,N_8794);
or U8882 (N_8882,N_8755,N_8736);
nor U8883 (N_8883,N_8771,N_8787);
and U8884 (N_8884,N_8753,N_8764);
and U8885 (N_8885,N_8705,N_8789);
nand U8886 (N_8886,N_8724,N_8712);
xnor U8887 (N_8887,N_8799,N_8782);
xor U8888 (N_8888,N_8738,N_8722);
nor U8889 (N_8889,N_8773,N_8795);
or U8890 (N_8890,N_8759,N_8796);
nand U8891 (N_8891,N_8705,N_8795);
nor U8892 (N_8892,N_8792,N_8791);
xnor U8893 (N_8893,N_8722,N_8730);
or U8894 (N_8894,N_8708,N_8759);
and U8895 (N_8895,N_8795,N_8743);
or U8896 (N_8896,N_8753,N_8773);
nand U8897 (N_8897,N_8755,N_8756);
nor U8898 (N_8898,N_8719,N_8746);
nand U8899 (N_8899,N_8781,N_8723);
nor U8900 (N_8900,N_8886,N_8845);
or U8901 (N_8901,N_8834,N_8896);
xor U8902 (N_8902,N_8872,N_8848);
nand U8903 (N_8903,N_8830,N_8895);
nor U8904 (N_8904,N_8889,N_8876);
and U8905 (N_8905,N_8861,N_8841);
or U8906 (N_8906,N_8835,N_8806);
nor U8907 (N_8907,N_8866,N_8825);
nor U8908 (N_8908,N_8898,N_8827);
nor U8909 (N_8909,N_8887,N_8838);
xor U8910 (N_8910,N_8839,N_8897);
xnor U8911 (N_8911,N_8885,N_8802);
or U8912 (N_8912,N_8891,N_8819);
nor U8913 (N_8913,N_8852,N_8853);
or U8914 (N_8914,N_8826,N_8844);
or U8915 (N_8915,N_8851,N_8808);
nand U8916 (N_8916,N_8831,N_8800);
nor U8917 (N_8917,N_8842,N_8888);
or U8918 (N_8918,N_8812,N_8874);
nand U8919 (N_8919,N_8815,N_8854);
nor U8920 (N_8920,N_8855,N_8871);
nor U8921 (N_8921,N_8884,N_8865);
nand U8922 (N_8922,N_8879,N_8864);
nor U8923 (N_8923,N_8804,N_8823);
or U8924 (N_8924,N_8881,N_8880);
nor U8925 (N_8925,N_8849,N_8846);
nor U8926 (N_8926,N_8833,N_8822);
and U8927 (N_8927,N_8890,N_8810);
and U8928 (N_8928,N_8878,N_8814);
or U8929 (N_8929,N_8816,N_8829);
xor U8930 (N_8930,N_8894,N_8807);
and U8931 (N_8931,N_8860,N_8862);
xnor U8932 (N_8932,N_8818,N_8824);
nor U8933 (N_8933,N_8821,N_8857);
xnor U8934 (N_8934,N_8803,N_8832);
and U8935 (N_8935,N_8869,N_8856);
nand U8936 (N_8936,N_8820,N_8875);
nor U8937 (N_8937,N_8813,N_8883);
xor U8938 (N_8938,N_8868,N_8859);
and U8939 (N_8939,N_8870,N_8899);
nand U8940 (N_8940,N_8828,N_8893);
nor U8941 (N_8941,N_8892,N_8817);
nor U8942 (N_8942,N_8836,N_8843);
and U8943 (N_8943,N_8858,N_8847);
nand U8944 (N_8944,N_8840,N_8882);
or U8945 (N_8945,N_8811,N_8867);
or U8946 (N_8946,N_8877,N_8801);
and U8947 (N_8947,N_8873,N_8809);
nor U8948 (N_8948,N_8863,N_8805);
nor U8949 (N_8949,N_8850,N_8837);
nor U8950 (N_8950,N_8852,N_8893);
nor U8951 (N_8951,N_8874,N_8846);
xor U8952 (N_8952,N_8861,N_8869);
and U8953 (N_8953,N_8847,N_8804);
xnor U8954 (N_8954,N_8840,N_8842);
and U8955 (N_8955,N_8875,N_8850);
xor U8956 (N_8956,N_8820,N_8871);
xor U8957 (N_8957,N_8827,N_8853);
xnor U8958 (N_8958,N_8830,N_8820);
and U8959 (N_8959,N_8879,N_8880);
xnor U8960 (N_8960,N_8821,N_8813);
nand U8961 (N_8961,N_8875,N_8893);
and U8962 (N_8962,N_8837,N_8806);
nor U8963 (N_8963,N_8837,N_8845);
and U8964 (N_8964,N_8846,N_8861);
xnor U8965 (N_8965,N_8856,N_8887);
nand U8966 (N_8966,N_8806,N_8803);
or U8967 (N_8967,N_8890,N_8871);
nand U8968 (N_8968,N_8823,N_8833);
and U8969 (N_8969,N_8830,N_8810);
nor U8970 (N_8970,N_8895,N_8806);
and U8971 (N_8971,N_8845,N_8878);
or U8972 (N_8972,N_8868,N_8846);
xor U8973 (N_8973,N_8872,N_8810);
or U8974 (N_8974,N_8823,N_8871);
nor U8975 (N_8975,N_8866,N_8826);
nor U8976 (N_8976,N_8808,N_8892);
or U8977 (N_8977,N_8801,N_8811);
xnor U8978 (N_8978,N_8837,N_8873);
xor U8979 (N_8979,N_8885,N_8834);
or U8980 (N_8980,N_8837,N_8844);
or U8981 (N_8981,N_8891,N_8845);
and U8982 (N_8982,N_8868,N_8804);
xor U8983 (N_8983,N_8859,N_8880);
nand U8984 (N_8984,N_8874,N_8865);
or U8985 (N_8985,N_8835,N_8829);
nor U8986 (N_8986,N_8802,N_8881);
xnor U8987 (N_8987,N_8814,N_8877);
nand U8988 (N_8988,N_8812,N_8823);
nor U8989 (N_8989,N_8837,N_8819);
nand U8990 (N_8990,N_8892,N_8895);
and U8991 (N_8991,N_8888,N_8803);
and U8992 (N_8992,N_8836,N_8881);
or U8993 (N_8993,N_8818,N_8897);
and U8994 (N_8994,N_8876,N_8845);
nor U8995 (N_8995,N_8848,N_8809);
or U8996 (N_8996,N_8846,N_8803);
or U8997 (N_8997,N_8899,N_8891);
or U8998 (N_8998,N_8805,N_8897);
nor U8999 (N_8999,N_8873,N_8851);
xnor U9000 (N_9000,N_8966,N_8902);
nor U9001 (N_9001,N_8976,N_8998);
or U9002 (N_9002,N_8923,N_8900);
or U9003 (N_9003,N_8920,N_8939);
or U9004 (N_9004,N_8994,N_8934);
nand U9005 (N_9005,N_8972,N_8922);
nand U9006 (N_9006,N_8944,N_8967);
nand U9007 (N_9007,N_8982,N_8925);
nand U9008 (N_9008,N_8995,N_8949);
and U9009 (N_9009,N_8942,N_8956);
nand U9010 (N_9010,N_8947,N_8987);
or U9011 (N_9011,N_8901,N_8971);
xnor U9012 (N_9012,N_8983,N_8926);
nand U9013 (N_9013,N_8990,N_8959);
or U9014 (N_9014,N_8958,N_8984);
and U9015 (N_9015,N_8940,N_8904);
and U9016 (N_9016,N_8906,N_8964);
or U9017 (N_9017,N_8917,N_8955);
nor U9018 (N_9018,N_8991,N_8933);
xor U9019 (N_9019,N_8919,N_8954);
or U9020 (N_9020,N_8907,N_8935);
xnor U9021 (N_9021,N_8932,N_8973);
nand U9022 (N_9022,N_8946,N_8938);
nor U9023 (N_9023,N_8969,N_8979);
nand U9024 (N_9024,N_8910,N_8911);
or U9025 (N_9025,N_8943,N_8929);
nand U9026 (N_9026,N_8980,N_8997);
nand U9027 (N_9027,N_8931,N_8915);
and U9028 (N_9028,N_8985,N_8965);
nand U9029 (N_9029,N_8970,N_8941);
or U9030 (N_9030,N_8981,N_8908);
nor U9031 (N_9031,N_8961,N_8993);
or U9032 (N_9032,N_8952,N_8937);
or U9033 (N_9033,N_8992,N_8916);
xnor U9034 (N_9034,N_8936,N_8930);
nand U9035 (N_9035,N_8962,N_8960);
and U9036 (N_9036,N_8988,N_8905);
xnor U9037 (N_9037,N_8968,N_8986);
and U9038 (N_9038,N_8975,N_8977);
xor U9039 (N_9039,N_8918,N_8963);
nor U9040 (N_9040,N_8951,N_8927);
nand U9041 (N_9041,N_8903,N_8974);
and U9042 (N_9042,N_8989,N_8978);
xnor U9043 (N_9043,N_8921,N_8928);
and U9044 (N_9044,N_8912,N_8953);
xnor U9045 (N_9045,N_8914,N_8913);
and U9046 (N_9046,N_8924,N_8957);
xor U9047 (N_9047,N_8950,N_8948);
nand U9048 (N_9048,N_8945,N_8909);
and U9049 (N_9049,N_8999,N_8996);
nor U9050 (N_9050,N_8982,N_8923);
xnor U9051 (N_9051,N_8973,N_8904);
or U9052 (N_9052,N_8990,N_8995);
nand U9053 (N_9053,N_8974,N_8985);
nor U9054 (N_9054,N_8956,N_8994);
nor U9055 (N_9055,N_8931,N_8957);
nor U9056 (N_9056,N_8962,N_8923);
and U9057 (N_9057,N_8941,N_8953);
nor U9058 (N_9058,N_8951,N_8903);
and U9059 (N_9059,N_8995,N_8916);
nor U9060 (N_9060,N_8972,N_8980);
xnor U9061 (N_9061,N_8968,N_8969);
or U9062 (N_9062,N_8991,N_8961);
nand U9063 (N_9063,N_8996,N_8914);
nand U9064 (N_9064,N_8964,N_8908);
xnor U9065 (N_9065,N_8970,N_8945);
xor U9066 (N_9066,N_8972,N_8973);
or U9067 (N_9067,N_8972,N_8996);
and U9068 (N_9068,N_8946,N_8900);
or U9069 (N_9069,N_8918,N_8976);
or U9070 (N_9070,N_8972,N_8984);
nand U9071 (N_9071,N_8972,N_8938);
xnor U9072 (N_9072,N_8943,N_8986);
nand U9073 (N_9073,N_8949,N_8978);
nor U9074 (N_9074,N_8932,N_8950);
nand U9075 (N_9075,N_8927,N_8942);
xnor U9076 (N_9076,N_8960,N_8961);
nor U9077 (N_9077,N_8944,N_8971);
and U9078 (N_9078,N_8966,N_8903);
xnor U9079 (N_9079,N_8976,N_8965);
xnor U9080 (N_9080,N_8988,N_8904);
or U9081 (N_9081,N_8929,N_8979);
nor U9082 (N_9082,N_8910,N_8929);
nand U9083 (N_9083,N_8946,N_8973);
xor U9084 (N_9084,N_8960,N_8902);
nand U9085 (N_9085,N_8928,N_8955);
nor U9086 (N_9086,N_8976,N_8947);
nand U9087 (N_9087,N_8944,N_8908);
and U9088 (N_9088,N_8941,N_8918);
or U9089 (N_9089,N_8936,N_8995);
nor U9090 (N_9090,N_8934,N_8941);
xnor U9091 (N_9091,N_8969,N_8961);
nor U9092 (N_9092,N_8921,N_8945);
or U9093 (N_9093,N_8986,N_8993);
or U9094 (N_9094,N_8926,N_8915);
nand U9095 (N_9095,N_8975,N_8997);
nor U9096 (N_9096,N_8990,N_8938);
or U9097 (N_9097,N_8940,N_8987);
or U9098 (N_9098,N_8960,N_8947);
and U9099 (N_9099,N_8921,N_8956);
xor U9100 (N_9100,N_9084,N_9075);
and U9101 (N_9101,N_9062,N_9052);
nor U9102 (N_9102,N_9042,N_9040);
and U9103 (N_9103,N_9020,N_9011);
and U9104 (N_9104,N_9068,N_9070);
nor U9105 (N_9105,N_9045,N_9074);
and U9106 (N_9106,N_9021,N_9043);
nand U9107 (N_9107,N_9061,N_9099);
nor U9108 (N_9108,N_9051,N_9089);
or U9109 (N_9109,N_9044,N_9003);
nand U9110 (N_9110,N_9029,N_9034);
xnor U9111 (N_9111,N_9081,N_9080);
nor U9112 (N_9112,N_9049,N_9000);
xor U9113 (N_9113,N_9033,N_9063);
or U9114 (N_9114,N_9041,N_9028);
nor U9115 (N_9115,N_9024,N_9078);
nor U9116 (N_9116,N_9010,N_9058);
or U9117 (N_9117,N_9094,N_9006);
and U9118 (N_9118,N_9048,N_9086);
xor U9119 (N_9119,N_9064,N_9060);
nand U9120 (N_9120,N_9088,N_9018);
or U9121 (N_9121,N_9036,N_9039);
nor U9122 (N_9122,N_9056,N_9023);
and U9123 (N_9123,N_9093,N_9019);
nor U9124 (N_9124,N_9069,N_9053);
nand U9125 (N_9125,N_9085,N_9077);
nand U9126 (N_9126,N_9038,N_9082);
nor U9127 (N_9127,N_9013,N_9008);
and U9128 (N_9128,N_9050,N_9025);
or U9129 (N_9129,N_9097,N_9037);
nand U9130 (N_9130,N_9066,N_9059);
nor U9131 (N_9131,N_9007,N_9091);
and U9132 (N_9132,N_9079,N_9030);
or U9133 (N_9133,N_9031,N_9015);
and U9134 (N_9134,N_9046,N_9047);
and U9135 (N_9135,N_9009,N_9090);
xnor U9136 (N_9136,N_9001,N_9012);
or U9137 (N_9137,N_9022,N_9027);
xnor U9138 (N_9138,N_9095,N_9016);
or U9139 (N_9139,N_9073,N_9087);
and U9140 (N_9140,N_9017,N_9076);
nor U9141 (N_9141,N_9055,N_9092);
nand U9142 (N_9142,N_9065,N_9067);
or U9143 (N_9143,N_9014,N_9072);
nand U9144 (N_9144,N_9002,N_9035);
nand U9145 (N_9145,N_9054,N_9057);
xnor U9146 (N_9146,N_9026,N_9083);
nor U9147 (N_9147,N_9096,N_9032);
nand U9148 (N_9148,N_9005,N_9098);
nand U9149 (N_9149,N_9071,N_9004);
nand U9150 (N_9150,N_9019,N_9028);
or U9151 (N_9151,N_9004,N_9059);
nor U9152 (N_9152,N_9043,N_9086);
nor U9153 (N_9153,N_9070,N_9002);
nand U9154 (N_9154,N_9080,N_9010);
nor U9155 (N_9155,N_9058,N_9039);
nor U9156 (N_9156,N_9016,N_9009);
and U9157 (N_9157,N_9011,N_9059);
or U9158 (N_9158,N_9035,N_9012);
or U9159 (N_9159,N_9021,N_9034);
and U9160 (N_9160,N_9084,N_9021);
nor U9161 (N_9161,N_9009,N_9021);
or U9162 (N_9162,N_9023,N_9091);
xor U9163 (N_9163,N_9017,N_9056);
nor U9164 (N_9164,N_9041,N_9060);
and U9165 (N_9165,N_9071,N_9010);
xor U9166 (N_9166,N_9032,N_9038);
xor U9167 (N_9167,N_9047,N_9076);
and U9168 (N_9168,N_9042,N_9012);
nor U9169 (N_9169,N_9014,N_9004);
nor U9170 (N_9170,N_9004,N_9031);
nor U9171 (N_9171,N_9096,N_9012);
nor U9172 (N_9172,N_9075,N_9026);
or U9173 (N_9173,N_9082,N_9062);
nand U9174 (N_9174,N_9078,N_9034);
nand U9175 (N_9175,N_9040,N_9033);
or U9176 (N_9176,N_9026,N_9004);
xor U9177 (N_9177,N_9077,N_9018);
and U9178 (N_9178,N_9020,N_9092);
nor U9179 (N_9179,N_9048,N_9008);
and U9180 (N_9180,N_9084,N_9068);
nand U9181 (N_9181,N_9004,N_9065);
nand U9182 (N_9182,N_9030,N_9069);
or U9183 (N_9183,N_9065,N_9033);
and U9184 (N_9184,N_9002,N_9005);
xnor U9185 (N_9185,N_9040,N_9014);
and U9186 (N_9186,N_9035,N_9049);
and U9187 (N_9187,N_9075,N_9049);
or U9188 (N_9188,N_9073,N_9004);
xor U9189 (N_9189,N_9076,N_9064);
or U9190 (N_9190,N_9082,N_9092);
xnor U9191 (N_9191,N_9074,N_9022);
or U9192 (N_9192,N_9030,N_9066);
nor U9193 (N_9193,N_9009,N_9038);
and U9194 (N_9194,N_9082,N_9084);
nor U9195 (N_9195,N_9008,N_9097);
nand U9196 (N_9196,N_9065,N_9074);
xor U9197 (N_9197,N_9038,N_9004);
xor U9198 (N_9198,N_9066,N_9044);
nor U9199 (N_9199,N_9047,N_9064);
xor U9200 (N_9200,N_9114,N_9102);
xor U9201 (N_9201,N_9112,N_9119);
nor U9202 (N_9202,N_9121,N_9173);
or U9203 (N_9203,N_9171,N_9115);
nand U9204 (N_9204,N_9176,N_9174);
nand U9205 (N_9205,N_9191,N_9101);
nand U9206 (N_9206,N_9166,N_9188);
xor U9207 (N_9207,N_9165,N_9153);
nor U9208 (N_9208,N_9135,N_9162);
or U9209 (N_9209,N_9184,N_9120);
xnor U9210 (N_9210,N_9110,N_9199);
and U9211 (N_9211,N_9111,N_9168);
and U9212 (N_9212,N_9129,N_9170);
nor U9213 (N_9213,N_9124,N_9145);
and U9214 (N_9214,N_9118,N_9180);
or U9215 (N_9215,N_9142,N_9139);
nand U9216 (N_9216,N_9198,N_9152);
or U9217 (N_9217,N_9132,N_9144);
nor U9218 (N_9218,N_9181,N_9147);
nor U9219 (N_9219,N_9190,N_9109);
or U9220 (N_9220,N_9130,N_9137);
nand U9221 (N_9221,N_9106,N_9149);
and U9222 (N_9222,N_9146,N_9183);
nand U9223 (N_9223,N_9157,N_9116);
nand U9224 (N_9224,N_9134,N_9143);
and U9225 (N_9225,N_9136,N_9100);
xnor U9226 (N_9226,N_9103,N_9128);
and U9227 (N_9227,N_9107,N_9193);
xnor U9228 (N_9228,N_9178,N_9164);
and U9229 (N_9229,N_9108,N_9138);
and U9230 (N_9230,N_9185,N_9154);
and U9231 (N_9231,N_9127,N_9141);
and U9232 (N_9232,N_9187,N_9150);
nand U9233 (N_9233,N_9195,N_9159);
nor U9234 (N_9234,N_9104,N_9175);
nand U9235 (N_9235,N_9156,N_9123);
and U9236 (N_9236,N_9122,N_9169);
or U9237 (N_9237,N_9197,N_9179);
and U9238 (N_9238,N_9160,N_9167);
nor U9239 (N_9239,N_9192,N_9172);
and U9240 (N_9240,N_9194,N_9117);
and U9241 (N_9241,N_9189,N_9177);
xnor U9242 (N_9242,N_9161,N_9113);
and U9243 (N_9243,N_9163,N_9140);
and U9244 (N_9244,N_9182,N_9105);
xnor U9245 (N_9245,N_9125,N_9151);
or U9246 (N_9246,N_9186,N_9133);
xor U9247 (N_9247,N_9158,N_9131);
and U9248 (N_9248,N_9148,N_9196);
and U9249 (N_9249,N_9126,N_9155);
nor U9250 (N_9250,N_9196,N_9180);
nor U9251 (N_9251,N_9118,N_9170);
or U9252 (N_9252,N_9161,N_9196);
xnor U9253 (N_9253,N_9171,N_9173);
nand U9254 (N_9254,N_9114,N_9150);
nand U9255 (N_9255,N_9107,N_9172);
xnor U9256 (N_9256,N_9173,N_9197);
and U9257 (N_9257,N_9156,N_9152);
xnor U9258 (N_9258,N_9133,N_9103);
nand U9259 (N_9259,N_9142,N_9161);
nor U9260 (N_9260,N_9105,N_9191);
nand U9261 (N_9261,N_9160,N_9139);
nand U9262 (N_9262,N_9143,N_9154);
and U9263 (N_9263,N_9159,N_9133);
xnor U9264 (N_9264,N_9118,N_9134);
xor U9265 (N_9265,N_9183,N_9157);
nand U9266 (N_9266,N_9183,N_9126);
xnor U9267 (N_9267,N_9104,N_9178);
nor U9268 (N_9268,N_9162,N_9195);
or U9269 (N_9269,N_9120,N_9178);
nor U9270 (N_9270,N_9182,N_9180);
nand U9271 (N_9271,N_9157,N_9104);
nor U9272 (N_9272,N_9136,N_9194);
nand U9273 (N_9273,N_9114,N_9167);
nor U9274 (N_9274,N_9145,N_9112);
or U9275 (N_9275,N_9155,N_9144);
xor U9276 (N_9276,N_9158,N_9120);
nor U9277 (N_9277,N_9142,N_9188);
xor U9278 (N_9278,N_9104,N_9144);
nor U9279 (N_9279,N_9183,N_9133);
xor U9280 (N_9280,N_9147,N_9182);
xnor U9281 (N_9281,N_9161,N_9198);
or U9282 (N_9282,N_9147,N_9178);
nor U9283 (N_9283,N_9144,N_9159);
or U9284 (N_9284,N_9169,N_9142);
nand U9285 (N_9285,N_9144,N_9145);
nand U9286 (N_9286,N_9128,N_9143);
xor U9287 (N_9287,N_9173,N_9158);
or U9288 (N_9288,N_9187,N_9137);
or U9289 (N_9289,N_9119,N_9169);
xor U9290 (N_9290,N_9197,N_9108);
xnor U9291 (N_9291,N_9114,N_9198);
nand U9292 (N_9292,N_9164,N_9127);
nor U9293 (N_9293,N_9120,N_9170);
nand U9294 (N_9294,N_9173,N_9119);
and U9295 (N_9295,N_9137,N_9109);
or U9296 (N_9296,N_9127,N_9189);
nor U9297 (N_9297,N_9130,N_9165);
or U9298 (N_9298,N_9165,N_9118);
or U9299 (N_9299,N_9145,N_9108);
nor U9300 (N_9300,N_9292,N_9265);
and U9301 (N_9301,N_9212,N_9242);
nand U9302 (N_9302,N_9299,N_9203);
and U9303 (N_9303,N_9219,N_9298);
and U9304 (N_9304,N_9233,N_9209);
xor U9305 (N_9305,N_9249,N_9235);
or U9306 (N_9306,N_9200,N_9284);
or U9307 (N_9307,N_9218,N_9225);
nor U9308 (N_9308,N_9246,N_9217);
nand U9309 (N_9309,N_9254,N_9210);
nand U9310 (N_9310,N_9248,N_9285);
nand U9311 (N_9311,N_9228,N_9282);
and U9312 (N_9312,N_9216,N_9204);
nand U9313 (N_9313,N_9238,N_9229);
and U9314 (N_9314,N_9286,N_9258);
xnor U9315 (N_9315,N_9289,N_9205);
xor U9316 (N_9316,N_9240,N_9295);
and U9317 (N_9317,N_9237,N_9291);
xor U9318 (N_9318,N_9260,N_9234);
xor U9319 (N_9319,N_9226,N_9230);
and U9320 (N_9320,N_9250,N_9293);
or U9321 (N_9321,N_9243,N_9206);
and U9322 (N_9322,N_9208,N_9220);
nand U9323 (N_9323,N_9270,N_9257);
xor U9324 (N_9324,N_9278,N_9294);
or U9325 (N_9325,N_9268,N_9296);
xor U9326 (N_9326,N_9283,N_9244);
nand U9327 (N_9327,N_9251,N_9202);
nand U9328 (N_9328,N_9224,N_9274);
or U9329 (N_9329,N_9236,N_9247);
xnor U9330 (N_9330,N_9264,N_9266);
nand U9331 (N_9331,N_9241,N_9255);
xor U9332 (N_9332,N_9213,N_9245);
and U9333 (N_9333,N_9277,N_9207);
nand U9334 (N_9334,N_9276,N_9223);
or U9335 (N_9335,N_9252,N_9271);
xnor U9336 (N_9336,N_9231,N_9273);
and U9337 (N_9337,N_9201,N_9263);
or U9338 (N_9338,N_9227,N_9279);
nand U9339 (N_9339,N_9256,N_9215);
or U9340 (N_9340,N_9253,N_9211);
nor U9341 (N_9341,N_9269,N_9239);
or U9342 (N_9342,N_9272,N_9259);
xnor U9343 (N_9343,N_9262,N_9222);
nor U9344 (N_9344,N_9281,N_9297);
or U9345 (N_9345,N_9221,N_9287);
xor U9346 (N_9346,N_9232,N_9280);
nor U9347 (N_9347,N_9267,N_9290);
nand U9348 (N_9348,N_9275,N_9214);
nand U9349 (N_9349,N_9288,N_9261);
xor U9350 (N_9350,N_9246,N_9207);
nand U9351 (N_9351,N_9239,N_9291);
and U9352 (N_9352,N_9244,N_9225);
and U9353 (N_9353,N_9257,N_9275);
xor U9354 (N_9354,N_9216,N_9242);
nor U9355 (N_9355,N_9294,N_9285);
and U9356 (N_9356,N_9280,N_9264);
and U9357 (N_9357,N_9213,N_9211);
nor U9358 (N_9358,N_9259,N_9204);
xnor U9359 (N_9359,N_9230,N_9214);
or U9360 (N_9360,N_9259,N_9201);
or U9361 (N_9361,N_9270,N_9258);
nand U9362 (N_9362,N_9209,N_9279);
nand U9363 (N_9363,N_9263,N_9247);
nand U9364 (N_9364,N_9210,N_9229);
or U9365 (N_9365,N_9247,N_9286);
and U9366 (N_9366,N_9225,N_9295);
xnor U9367 (N_9367,N_9232,N_9262);
xnor U9368 (N_9368,N_9208,N_9266);
nand U9369 (N_9369,N_9271,N_9202);
nor U9370 (N_9370,N_9262,N_9248);
and U9371 (N_9371,N_9281,N_9225);
or U9372 (N_9372,N_9297,N_9268);
or U9373 (N_9373,N_9207,N_9242);
nand U9374 (N_9374,N_9227,N_9244);
or U9375 (N_9375,N_9259,N_9238);
nor U9376 (N_9376,N_9256,N_9242);
and U9377 (N_9377,N_9259,N_9236);
and U9378 (N_9378,N_9203,N_9259);
nand U9379 (N_9379,N_9223,N_9239);
or U9380 (N_9380,N_9211,N_9289);
xor U9381 (N_9381,N_9285,N_9282);
and U9382 (N_9382,N_9248,N_9224);
nand U9383 (N_9383,N_9227,N_9200);
xor U9384 (N_9384,N_9218,N_9238);
nand U9385 (N_9385,N_9208,N_9280);
and U9386 (N_9386,N_9277,N_9235);
nor U9387 (N_9387,N_9244,N_9218);
nand U9388 (N_9388,N_9245,N_9243);
and U9389 (N_9389,N_9227,N_9249);
and U9390 (N_9390,N_9243,N_9235);
or U9391 (N_9391,N_9227,N_9268);
nor U9392 (N_9392,N_9214,N_9244);
xor U9393 (N_9393,N_9295,N_9238);
and U9394 (N_9394,N_9235,N_9269);
xnor U9395 (N_9395,N_9232,N_9246);
xnor U9396 (N_9396,N_9220,N_9244);
and U9397 (N_9397,N_9267,N_9264);
and U9398 (N_9398,N_9259,N_9262);
nand U9399 (N_9399,N_9229,N_9261);
or U9400 (N_9400,N_9379,N_9399);
and U9401 (N_9401,N_9383,N_9307);
and U9402 (N_9402,N_9376,N_9365);
or U9403 (N_9403,N_9320,N_9380);
nand U9404 (N_9404,N_9315,N_9354);
nor U9405 (N_9405,N_9337,N_9369);
or U9406 (N_9406,N_9385,N_9318);
and U9407 (N_9407,N_9352,N_9311);
and U9408 (N_9408,N_9341,N_9346);
and U9409 (N_9409,N_9310,N_9325);
nand U9410 (N_9410,N_9340,N_9324);
nand U9411 (N_9411,N_9349,N_9394);
xnor U9412 (N_9412,N_9322,N_9359);
or U9413 (N_9413,N_9378,N_9330);
and U9414 (N_9414,N_9332,N_9309);
or U9415 (N_9415,N_9319,N_9398);
xnor U9416 (N_9416,N_9304,N_9356);
nand U9417 (N_9417,N_9377,N_9389);
or U9418 (N_9418,N_9338,N_9300);
or U9419 (N_9419,N_9312,N_9314);
or U9420 (N_9420,N_9348,N_9331);
xor U9421 (N_9421,N_9317,N_9328);
nor U9422 (N_9422,N_9327,N_9343);
nor U9423 (N_9423,N_9397,N_9388);
xor U9424 (N_9424,N_9382,N_9353);
and U9425 (N_9425,N_9390,N_9339);
and U9426 (N_9426,N_9321,N_9305);
and U9427 (N_9427,N_9386,N_9375);
nand U9428 (N_9428,N_9368,N_9393);
nand U9429 (N_9429,N_9374,N_9364);
nand U9430 (N_9430,N_9357,N_9335);
or U9431 (N_9431,N_9361,N_9345);
and U9432 (N_9432,N_9336,N_9381);
nor U9433 (N_9433,N_9363,N_9342);
xnor U9434 (N_9434,N_9306,N_9387);
or U9435 (N_9435,N_9395,N_9313);
nor U9436 (N_9436,N_9391,N_9371);
and U9437 (N_9437,N_9358,N_9329);
or U9438 (N_9438,N_9302,N_9362);
xor U9439 (N_9439,N_9370,N_9355);
nor U9440 (N_9440,N_9373,N_9372);
or U9441 (N_9441,N_9396,N_9316);
and U9442 (N_9442,N_9334,N_9303);
or U9443 (N_9443,N_9347,N_9384);
xor U9444 (N_9444,N_9323,N_9344);
xor U9445 (N_9445,N_9308,N_9392);
xor U9446 (N_9446,N_9326,N_9350);
xnor U9447 (N_9447,N_9367,N_9351);
and U9448 (N_9448,N_9366,N_9333);
or U9449 (N_9449,N_9360,N_9301);
nor U9450 (N_9450,N_9352,N_9307);
nand U9451 (N_9451,N_9393,N_9398);
xor U9452 (N_9452,N_9325,N_9318);
nor U9453 (N_9453,N_9304,N_9337);
nand U9454 (N_9454,N_9324,N_9321);
xnor U9455 (N_9455,N_9373,N_9302);
nor U9456 (N_9456,N_9387,N_9391);
nor U9457 (N_9457,N_9399,N_9335);
and U9458 (N_9458,N_9309,N_9345);
nor U9459 (N_9459,N_9312,N_9399);
or U9460 (N_9460,N_9332,N_9306);
or U9461 (N_9461,N_9339,N_9329);
nand U9462 (N_9462,N_9300,N_9346);
nor U9463 (N_9463,N_9393,N_9381);
and U9464 (N_9464,N_9379,N_9378);
nor U9465 (N_9465,N_9386,N_9378);
or U9466 (N_9466,N_9355,N_9335);
or U9467 (N_9467,N_9360,N_9399);
nor U9468 (N_9468,N_9335,N_9304);
xnor U9469 (N_9469,N_9344,N_9398);
nor U9470 (N_9470,N_9324,N_9329);
or U9471 (N_9471,N_9334,N_9387);
nor U9472 (N_9472,N_9393,N_9377);
and U9473 (N_9473,N_9350,N_9331);
nand U9474 (N_9474,N_9352,N_9314);
xnor U9475 (N_9475,N_9351,N_9328);
and U9476 (N_9476,N_9384,N_9399);
xor U9477 (N_9477,N_9318,N_9326);
and U9478 (N_9478,N_9346,N_9359);
nand U9479 (N_9479,N_9356,N_9345);
or U9480 (N_9480,N_9398,N_9366);
and U9481 (N_9481,N_9347,N_9321);
xnor U9482 (N_9482,N_9378,N_9312);
xnor U9483 (N_9483,N_9375,N_9326);
or U9484 (N_9484,N_9387,N_9392);
nand U9485 (N_9485,N_9382,N_9324);
nand U9486 (N_9486,N_9327,N_9377);
nor U9487 (N_9487,N_9325,N_9302);
nor U9488 (N_9488,N_9341,N_9308);
nand U9489 (N_9489,N_9365,N_9375);
nor U9490 (N_9490,N_9302,N_9353);
nor U9491 (N_9491,N_9312,N_9357);
nand U9492 (N_9492,N_9318,N_9309);
and U9493 (N_9493,N_9361,N_9350);
xnor U9494 (N_9494,N_9366,N_9341);
and U9495 (N_9495,N_9356,N_9373);
nor U9496 (N_9496,N_9328,N_9322);
nand U9497 (N_9497,N_9388,N_9322);
xnor U9498 (N_9498,N_9340,N_9372);
nor U9499 (N_9499,N_9320,N_9356);
and U9500 (N_9500,N_9402,N_9414);
and U9501 (N_9501,N_9413,N_9464);
and U9502 (N_9502,N_9417,N_9470);
and U9503 (N_9503,N_9404,N_9483);
nor U9504 (N_9504,N_9471,N_9479);
xor U9505 (N_9505,N_9496,N_9445);
nand U9506 (N_9506,N_9482,N_9453);
nor U9507 (N_9507,N_9447,N_9439);
xor U9508 (N_9508,N_9486,N_9450);
xor U9509 (N_9509,N_9499,N_9456);
xor U9510 (N_9510,N_9400,N_9493);
and U9511 (N_9511,N_9488,N_9425);
nor U9512 (N_9512,N_9476,N_9489);
xnor U9513 (N_9513,N_9465,N_9498);
xor U9514 (N_9514,N_9484,N_9431);
nand U9515 (N_9515,N_9408,N_9478);
or U9516 (N_9516,N_9481,N_9475);
nor U9517 (N_9517,N_9454,N_9474);
xor U9518 (N_9518,N_9419,N_9411);
and U9519 (N_9519,N_9415,N_9418);
and U9520 (N_9520,N_9492,N_9462);
nor U9521 (N_9521,N_9495,N_9448);
and U9522 (N_9522,N_9468,N_9491);
nand U9523 (N_9523,N_9463,N_9458);
xor U9524 (N_9524,N_9472,N_9436);
xor U9525 (N_9525,N_9438,N_9432);
xnor U9526 (N_9526,N_9426,N_9412);
xor U9527 (N_9527,N_9451,N_9455);
or U9528 (N_9528,N_9430,N_9424);
or U9529 (N_9529,N_9449,N_9490);
or U9530 (N_9530,N_9429,N_9443);
or U9531 (N_9531,N_9480,N_9441);
and U9532 (N_9532,N_9459,N_9497);
nor U9533 (N_9533,N_9467,N_9406);
xor U9534 (N_9534,N_9494,N_9444);
nor U9535 (N_9535,N_9416,N_9469);
nor U9536 (N_9536,N_9428,N_9446);
or U9537 (N_9537,N_9420,N_9422);
and U9538 (N_9538,N_9440,N_9421);
nor U9539 (N_9539,N_9405,N_9407);
or U9540 (N_9540,N_9403,N_9460);
nand U9541 (N_9541,N_9435,N_9487);
nand U9542 (N_9542,N_9434,N_9442);
nor U9543 (N_9543,N_9457,N_9410);
xor U9544 (N_9544,N_9433,N_9452);
nand U9545 (N_9545,N_9427,N_9466);
xor U9546 (N_9546,N_9423,N_9485);
or U9547 (N_9547,N_9461,N_9477);
or U9548 (N_9548,N_9409,N_9473);
nand U9549 (N_9549,N_9401,N_9437);
or U9550 (N_9550,N_9485,N_9440);
or U9551 (N_9551,N_9477,N_9429);
nor U9552 (N_9552,N_9466,N_9459);
or U9553 (N_9553,N_9456,N_9413);
xor U9554 (N_9554,N_9444,N_9417);
and U9555 (N_9555,N_9465,N_9427);
nand U9556 (N_9556,N_9448,N_9404);
nor U9557 (N_9557,N_9433,N_9489);
and U9558 (N_9558,N_9477,N_9463);
and U9559 (N_9559,N_9491,N_9429);
or U9560 (N_9560,N_9401,N_9476);
nor U9561 (N_9561,N_9450,N_9411);
or U9562 (N_9562,N_9481,N_9497);
nand U9563 (N_9563,N_9457,N_9479);
nand U9564 (N_9564,N_9495,N_9408);
nand U9565 (N_9565,N_9472,N_9493);
xnor U9566 (N_9566,N_9421,N_9414);
xor U9567 (N_9567,N_9495,N_9430);
xnor U9568 (N_9568,N_9416,N_9413);
and U9569 (N_9569,N_9443,N_9414);
xor U9570 (N_9570,N_9469,N_9475);
or U9571 (N_9571,N_9474,N_9427);
nor U9572 (N_9572,N_9454,N_9451);
and U9573 (N_9573,N_9431,N_9419);
nor U9574 (N_9574,N_9407,N_9438);
nor U9575 (N_9575,N_9490,N_9497);
or U9576 (N_9576,N_9408,N_9419);
xor U9577 (N_9577,N_9410,N_9482);
xnor U9578 (N_9578,N_9420,N_9448);
and U9579 (N_9579,N_9406,N_9431);
nor U9580 (N_9580,N_9408,N_9401);
nor U9581 (N_9581,N_9483,N_9444);
and U9582 (N_9582,N_9402,N_9405);
and U9583 (N_9583,N_9482,N_9441);
or U9584 (N_9584,N_9499,N_9421);
nand U9585 (N_9585,N_9461,N_9400);
or U9586 (N_9586,N_9462,N_9498);
xor U9587 (N_9587,N_9457,N_9402);
and U9588 (N_9588,N_9435,N_9403);
and U9589 (N_9589,N_9456,N_9480);
or U9590 (N_9590,N_9428,N_9466);
and U9591 (N_9591,N_9456,N_9491);
xor U9592 (N_9592,N_9459,N_9479);
or U9593 (N_9593,N_9412,N_9425);
or U9594 (N_9594,N_9419,N_9402);
xor U9595 (N_9595,N_9479,N_9477);
xnor U9596 (N_9596,N_9473,N_9427);
and U9597 (N_9597,N_9460,N_9457);
nand U9598 (N_9598,N_9406,N_9408);
xnor U9599 (N_9599,N_9411,N_9493);
nand U9600 (N_9600,N_9565,N_9581);
nand U9601 (N_9601,N_9599,N_9587);
nor U9602 (N_9602,N_9588,N_9585);
xor U9603 (N_9603,N_9522,N_9558);
nand U9604 (N_9604,N_9500,N_9556);
or U9605 (N_9605,N_9508,N_9507);
and U9606 (N_9606,N_9563,N_9503);
and U9607 (N_9607,N_9591,N_9578);
xnor U9608 (N_9608,N_9520,N_9559);
nand U9609 (N_9609,N_9574,N_9506);
or U9610 (N_9610,N_9577,N_9518);
nand U9611 (N_9611,N_9596,N_9521);
nand U9612 (N_9612,N_9555,N_9534);
or U9613 (N_9613,N_9502,N_9553);
and U9614 (N_9614,N_9523,N_9525);
nor U9615 (N_9615,N_9582,N_9593);
nor U9616 (N_9616,N_9547,N_9573);
xor U9617 (N_9617,N_9583,N_9514);
nand U9618 (N_9618,N_9528,N_9510);
and U9619 (N_9619,N_9570,N_9550);
and U9620 (N_9620,N_9575,N_9572);
nand U9621 (N_9621,N_9595,N_9540);
and U9622 (N_9622,N_9524,N_9576);
nand U9623 (N_9623,N_9566,N_9571);
nor U9624 (N_9624,N_9551,N_9594);
nor U9625 (N_9625,N_9526,N_9515);
or U9626 (N_9626,N_9568,N_9533);
xnor U9627 (N_9627,N_9519,N_9513);
nor U9628 (N_9628,N_9532,N_9501);
nor U9629 (N_9629,N_9561,N_9569);
xor U9630 (N_9630,N_9512,N_9579);
xnor U9631 (N_9631,N_9554,N_9516);
and U9632 (N_9632,N_9580,N_9505);
xor U9633 (N_9633,N_9504,N_9531);
or U9634 (N_9634,N_9557,N_9598);
and U9635 (N_9635,N_9592,N_9564);
and U9636 (N_9636,N_9545,N_9597);
nor U9637 (N_9637,N_9542,N_9539);
and U9638 (N_9638,N_9567,N_9544);
or U9639 (N_9639,N_9527,N_9530);
xnor U9640 (N_9640,N_9517,N_9589);
or U9641 (N_9641,N_9536,N_9546);
and U9642 (N_9642,N_9552,N_9535);
and U9643 (N_9643,N_9584,N_9538);
xor U9644 (N_9644,N_9562,N_9543);
or U9645 (N_9645,N_9529,N_9586);
xor U9646 (N_9646,N_9537,N_9560);
xor U9647 (N_9647,N_9511,N_9541);
xnor U9648 (N_9648,N_9590,N_9509);
xnor U9649 (N_9649,N_9549,N_9548);
and U9650 (N_9650,N_9505,N_9598);
xor U9651 (N_9651,N_9523,N_9502);
or U9652 (N_9652,N_9548,N_9543);
nand U9653 (N_9653,N_9554,N_9509);
and U9654 (N_9654,N_9540,N_9548);
xor U9655 (N_9655,N_9501,N_9533);
nor U9656 (N_9656,N_9509,N_9553);
nand U9657 (N_9657,N_9576,N_9542);
and U9658 (N_9658,N_9565,N_9558);
or U9659 (N_9659,N_9562,N_9520);
nand U9660 (N_9660,N_9552,N_9584);
xor U9661 (N_9661,N_9593,N_9560);
or U9662 (N_9662,N_9544,N_9552);
nor U9663 (N_9663,N_9564,N_9511);
nor U9664 (N_9664,N_9554,N_9504);
nor U9665 (N_9665,N_9563,N_9506);
nand U9666 (N_9666,N_9576,N_9564);
nand U9667 (N_9667,N_9509,N_9563);
nor U9668 (N_9668,N_9502,N_9585);
or U9669 (N_9669,N_9518,N_9591);
nor U9670 (N_9670,N_9535,N_9576);
and U9671 (N_9671,N_9501,N_9545);
nand U9672 (N_9672,N_9505,N_9577);
xor U9673 (N_9673,N_9522,N_9511);
nor U9674 (N_9674,N_9545,N_9564);
nand U9675 (N_9675,N_9599,N_9579);
nor U9676 (N_9676,N_9538,N_9594);
and U9677 (N_9677,N_9554,N_9581);
nor U9678 (N_9678,N_9540,N_9515);
nor U9679 (N_9679,N_9520,N_9547);
or U9680 (N_9680,N_9581,N_9536);
and U9681 (N_9681,N_9578,N_9529);
xnor U9682 (N_9682,N_9568,N_9585);
xor U9683 (N_9683,N_9598,N_9583);
nor U9684 (N_9684,N_9552,N_9571);
nor U9685 (N_9685,N_9547,N_9593);
and U9686 (N_9686,N_9561,N_9515);
nand U9687 (N_9687,N_9535,N_9558);
or U9688 (N_9688,N_9555,N_9544);
and U9689 (N_9689,N_9572,N_9515);
or U9690 (N_9690,N_9541,N_9573);
nand U9691 (N_9691,N_9528,N_9518);
nor U9692 (N_9692,N_9579,N_9591);
xor U9693 (N_9693,N_9596,N_9509);
and U9694 (N_9694,N_9519,N_9544);
and U9695 (N_9695,N_9599,N_9539);
nor U9696 (N_9696,N_9530,N_9511);
and U9697 (N_9697,N_9564,N_9597);
or U9698 (N_9698,N_9562,N_9538);
or U9699 (N_9699,N_9559,N_9543);
or U9700 (N_9700,N_9610,N_9685);
and U9701 (N_9701,N_9620,N_9622);
nor U9702 (N_9702,N_9631,N_9617);
and U9703 (N_9703,N_9657,N_9643);
nand U9704 (N_9704,N_9698,N_9673);
nand U9705 (N_9705,N_9665,N_9683);
or U9706 (N_9706,N_9606,N_9681);
and U9707 (N_9707,N_9625,N_9613);
nor U9708 (N_9708,N_9654,N_9621);
xor U9709 (N_9709,N_9647,N_9603);
nor U9710 (N_9710,N_9605,N_9637);
nand U9711 (N_9711,N_9626,N_9680);
xor U9712 (N_9712,N_9693,N_9634);
and U9713 (N_9713,N_9633,N_9629);
xnor U9714 (N_9714,N_9669,N_9691);
nand U9715 (N_9715,N_9687,N_9678);
xor U9716 (N_9716,N_9661,N_9639);
or U9717 (N_9717,N_9659,N_9618);
and U9718 (N_9718,N_9686,N_9664);
or U9719 (N_9719,N_9676,N_9609);
xnor U9720 (N_9720,N_9635,N_9646);
xor U9721 (N_9721,N_9619,N_9640);
and U9722 (N_9722,N_9627,N_9696);
xnor U9723 (N_9723,N_9632,N_9690);
xor U9724 (N_9724,N_9674,N_9649);
xnor U9725 (N_9725,N_9630,N_9688);
nor U9726 (N_9726,N_9684,N_9670);
nor U9727 (N_9727,N_9600,N_9694);
and U9728 (N_9728,N_9650,N_9616);
and U9729 (N_9729,N_9602,N_9623);
or U9730 (N_9730,N_9667,N_9672);
nor U9731 (N_9731,N_9677,N_9607);
or U9732 (N_9732,N_9652,N_9601);
xor U9733 (N_9733,N_9663,N_9648);
nor U9734 (N_9734,N_9612,N_9692);
or U9735 (N_9735,N_9697,N_9644);
xor U9736 (N_9736,N_9614,N_9636);
and U9737 (N_9737,N_9608,N_9638);
nor U9738 (N_9738,N_9666,N_9611);
and U9739 (N_9739,N_9628,N_9651);
and U9740 (N_9740,N_9604,N_9682);
and U9741 (N_9741,N_9679,N_9641);
xnor U9742 (N_9742,N_9695,N_9699);
xor U9743 (N_9743,N_9655,N_9645);
nor U9744 (N_9744,N_9658,N_9660);
nor U9745 (N_9745,N_9671,N_9615);
or U9746 (N_9746,N_9624,N_9662);
or U9747 (N_9747,N_9656,N_9668);
and U9748 (N_9748,N_9689,N_9675);
xnor U9749 (N_9749,N_9653,N_9642);
nand U9750 (N_9750,N_9655,N_9695);
and U9751 (N_9751,N_9625,N_9605);
xnor U9752 (N_9752,N_9608,N_9630);
and U9753 (N_9753,N_9674,N_9645);
nand U9754 (N_9754,N_9637,N_9620);
and U9755 (N_9755,N_9663,N_9666);
or U9756 (N_9756,N_9630,N_9683);
nor U9757 (N_9757,N_9654,N_9628);
xnor U9758 (N_9758,N_9618,N_9603);
xor U9759 (N_9759,N_9686,N_9699);
or U9760 (N_9760,N_9694,N_9643);
nand U9761 (N_9761,N_9666,N_9606);
and U9762 (N_9762,N_9632,N_9686);
or U9763 (N_9763,N_9670,N_9696);
nand U9764 (N_9764,N_9611,N_9648);
xnor U9765 (N_9765,N_9605,N_9646);
nor U9766 (N_9766,N_9609,N_9673);
nand U9767 (N_9767,N_9612,N_9653);
nand U9768 (N_9768,N_9602,N_9692);
nor U9769 (N_9769,N_9658,N_9661);
xor U9770 (N_9770,N_9663,N_9685);
xor U9771 (N_9771,N_9638,N_9669);
nor U9772 (N_9772,N_9632,N_9660);
nor U9773 (N_9773,N_9681,N_9610);
and U9774 (N_9774,N_9675,N_9671);
or U9775 (N_9775,N_9604,N_9638);
nor U9776 (N_9776,N_9626,N_9683);
nor U9777 (N_9777,N_9602,N_9688);
or U9778 (N_9778,N_9613,N_9640);
xor U9779 (N_9779,N_9676,N_9635);
or U9780 (N_9780,N_9604,N_9643);
nand U9781 (N_9781,N_9633,N_9612);
and U9782 (N_9782,N_9601,N_9615);
nand U9783 (N_9783,N_9624,N_9600);
xor U9784 (N_9784,N_9674,N_9680);
or U9785 (N_9785,N_9675,N_9602);
or U9786 (N_9786,N_9629,N_9654);
xor U9787 (N_9787,N_9659,N_9674);
nand U9788 (N_9788,N_9642,N_9608);
or U9789 (N_9789,N_9629,N_9685);
or U9790 (N_9790,N_9618,N_9645);
nor U9791 (N_9791,N_9622,N_9665);
nand U9792 (N_9792,N_9669,N_9601);
nand U9793 (N_9793,N_9646,N_9629);
nand U9794 (N_9794,N_9601,N_9651);
nand U9795 (N_9795,N_9699,N_9635);
nand U9796 (N_9796,N_9601,N_9694);
and U9797 (N_9797,N_9629,N_9667);
or U9798 (N_9798,N_9696,N_9639);
xnor U9799 (N_9799,N_9660,N_9672);
and U9800 (N_9800,N_9706,N_9702);
xnor U9801 (N_9801,N_9776,N_9762);
nand U9802 (N_9802,N_9701,N_9715);
nand U9803 (N_9803,N_9716,N_9765);
and U9804 (N_9804,N_9763,N_9786);
or U9805 (N_9805,N_9769,N_9720);
nand U9806 (N_9806,N_9714,N_9760);
xnor U9807 (N_9807,N_9770,N_9792);
xnor U9808 (N_9808,N_9703,N_9736);
xor U9809 (N_9809,N_9781,N_9708);
nand U9810 (N_9810,N_9751,N_9700);
xor U9811 (N_9811,N_9791,N_9747);
nand U9812 (N_9812,N_9789,N_9795);
nor U9813 (N_9813,N_9712,N_9705);
xnor U9814 (N_9814,N_9798,N_9794);
and U9815 (N_9815,N_9777,N_9718);
or U9816 (N_9816,N_9757,N_9771);
nand U9817 (N_9817,N_9787,N_9758);
nand U9818 (N_9818,N_9704,N_9796);
or U9819 (N_9819,N_9741,N_9709);
or U9820 (N_9820,N_9735,N_9755);
and U9821 (N_9821,N_9730,N_9783);
and U9822 (N_9822,N_9797,N_9790);
or U9823 (N_9823,N_9775,N_9768);
nor U9824 (N_9824,N_9734,N_9784);
xnor U9825 (N_9825,N_9728,N_9724);
nor U9826 (N_9826,N_9764,N_9753);
and U9827 (N_9827,N_9749,N_9713);
or U9828 (N_9828,N_9788,N_9719);
or U9829 (N_9829,N_9723,N_9772);
nor U9830 (N_9830,N_9711,N_9766);
nor U9831 (N_9831,N_9742,N_9726);
nor U9832 (N_9832,N_9733,N_9738);
and U9833 (N_9833,N_9778,N_9756);
xnor U9834 (N_9834,N_9717,N_9767);
nor U9835 (N_9835,N_9785,N_9740);
and U9836 (N_9836,N_9731,N_9793);
xor U9837 (N_9837,N_9737,N_9729);
nor U9838 (N_9838,N_9725,N_9748);
or U9839 (N_9839,N_9710,N_9759);
and U9840 (N_9840,N_9739,N_9745);
or U9841 (N_9841,N_9761,N_9744);
xnor U9842 (N_9842,N_9754,N_9721);
or U9843 (N_9843,N_9746,N_9752);
or U9844 (N_9844,N_9732,N_9707);
nor U9845 (N_9845,N_9782,N_9773);
nor U9846 (N_9846,N_9743,N_9727);
xor U9847 (N_9847,N_9774,N_9780);
nor U9848 (N_9848,N_9722,N_9799);
and U9849 (N_9849,N_9779,N_9750);
nor U9850 (N_9850,N_9718,N_9749);
and U9851 (N_9851,N_9718,N_9720);
or U9852 (N_9852,N_9788,N_9722);
nor U9853 (N_9853,N_9740,N_9794);
and U9854 (N_9854,N_9726,N_9785);
nand U9855 (N_9855,N_9786,N_9711);
nand U9856 (N_9856,N_9790,N_9777);
or U9857 (N_9857,N_9797,N_9780);
nand U9858 (N_9858,N_9775,N_9750);
or U9859 (N_9859,N_9731,N_9747);
or U9860 (N_9860,N_9786,N_9719);
xor U9861 (N_9861,N_9713,N_9731);
nand U9862 (N_9862,N_9755,N_9714);
xnor U9863 (N_9863,N_9794,N_9736);
nor U9864 (N_9864,N_9715,N_9722);
nor U9865 (N_9865,N_9718,N_9715);
nor U9866 (N_9866,N_9711,N_9787);
and U9867 (N_9867,N_9715,N_9723);
nand U9868 (N_9868,N_9704,N_9719);
nor U9869 (N_9869,N_9788,N_9761);
and U9870 (N_9870,N_9708,N_9775);
nand U9871 (N_9871,N_9778,N_9764);
nand U9872 (N_9872,N_9790,N_9774);
or U9873 (N_9873,N_9716,N_9707);
nor U9874 (N_9874,N_9774,N_9742);
xor U9875 (N_9875,N_9753,N_9740);
or U9876 (N_9876,N_9741,N_9773);
or U9877 (N_9877,N_9742,N_9789);
xor U9878 (N_9878,N_9792,N_9725);
or U9879 (N_9879,N_9739,N_9791);
nand U9880 (N_9880,N_9705,N_9760);
or U9881 (N_9881,N_9701,N_9765);
and U9882 (N_9882,N_9768,N_9718);
nor U9883 (N_9883,N_9732,N_9725);
xor U9884 (N_9884,N_9709,N_9744);
nand U9885 (N_9885,N_9761,N_9763);
and U9886 (N_9886,N_9714,N_9717);
and U9887 (N_9887,N_9781,N_9770);
and U9888 (N_9888,N_9731,N_9788);
or U9889 (N_9889,N_9721,N_9744);
xnor U9890 (N_9890,N_9700,N_9721);
nand U9891 (N_9891,N_9712,N_9749);
and U9892 (N_9892,N_9707,N_9701);
and U9893 (N_9893,N_9751,N_9799);
nand U9894 (N_9894,N_9745,N_9725);
xor U9895 (N_9895,N_9788,N_9785);
xnor U9896 (N_9896,N_9722,N_9701);
or U9897 (N_9897,N_9719,N_9757);
xor U9898 (N_9898,N_9724,N_9770);
nand U9899 (N_9899,N_9778,N_9749);
xor U9900 (N_9900,N_9810,N_9896);
nand U9901 (N_9901,N_9831,N_9844);
or U9902 (N_9902,N_9805,N_9832);
and U9903 (N_9903,N_9811,N_9858);
nand U9904 (N_9904,N_9880,N_9800);
nor U9905 (N_9905,N_9809,N_9877);
nor U9906 (N_9906,N_9815,N_9887);
or U9907 (N_9907,N_9890,N_9873);
or U9908 (N_9908,N_9820,N_9885);
nor U9909 (N_9909,N_9860,N_9835);
and U9910 (N_9910,N_9892,N_9855);
nor U9911 (N_9911,N_9841,N_9891);
xnor U9912 (N_9912,N_9803,N_9812);
or U9913 (N_9913,N_9851,N_9898);
xnor U9914 (N_9914,N_9876,N_9854);
nand U9915 (N_9915,N_9813,N_9827);
nor U9916 (N_9916,N_9826,N_9837);
xor U9917 (N_9917,N_9853,N_9839);
and U9918 (N_9918,N_9869,N_9861);
nor U9919 (N_9919,N_9875,N_9878);
or U9920 (N_9920,N_9806,N_9823);
and U9921 (N_9921,N_9856,N_9804);
nor U9922 (N_9922,N_9845,N_9828);
nor U9923 (N_9923,N_9871,N_9849);
xor U9924 (N_9924,N_9888,N_9893);
nor U9925 (N_9925,N_9847,N_9870);
nor U9926 (N_9926,N_9801,N_9821);
nor U9927 (N_9927,N_9864,N_9894);
and U9928 (N_9928,N_9843,N_9868);
nor U9929 (N_9929,N_9859,N_9830);
nand U9930 (N_9930,N_9816,N_9895);
or U9931 (N_9931,N_9857,N_9824);
and U9932 (N_9932,N_9846,N_9886);
or U9933 (N_9933,N_9850,N_9819);
nand U9934 (N_9934,N_9833,N_9865);
nand U9935 (N_9935,N_9863,N_9882);
nor U9936 (N_9936,N_9818,N_9834);
and U9937 (N_9937,N_9829,N_9889);
nor U9938 (N_9938,N_9872,N_9807);
nand U9939 (N_9939,N_9802,N_9822);
nor U9940 (N_9940,N_9825,N_9866);
nand U9941 (N_9941,N_9881,N_9862);
or U9942 (N_9942,N_9842,N_9867);
xnor U9943 (N_9943,N_9884,N_9897);
and U9944 (N_9944,N_9814,N_9879);
nor U9945 (N_9945,N_9883,N_9836);
nand U9946 (N_9946,N_9808,N_9852);
and U9947 (N_9947,N_9840,N_9817);
or U9948 (N_9948,N_9838,N_9874);
xor U9949 (N_9949,N_9848,N_9899);
nand U9950 (N_9950,N_9843,N_9817);
and U9951 (N_9951,N_9839,N_9885);
nand U9952 (N_9952,N_9850,N_9815);
nor U9953 (N_9953,N_9838,N_9867);
or U9954 (N_9954,N_9831,N_9813);
nor U9955 (N_9955,N_9896,N_9826);
xnor U9956 (N_9956,N_9882,N_9821);
or U9957 (N_9957,N_9895,N_9852);
nor U9958 (N_9958,N_9888,N_9837);
nor U9959 (N_9959,N_9823,N_9856);
nand U9960 (N_9960,N_9827,N_9889);
or U9961 (N_9961,N_9844,N_9855);
xor U9962 (N_9962,N_9871,N_9859);
or U9963 (N_9963,N_9844,N_9803);
and U9964 (N_9964,N_9869,N_9847);
nand U9965 (N_9965,N_9846,N_9802);
or U9966 (N_9966,N_9871,N_9819);
nor U9967 (N_9967,N_9884,N_9869);
nand U9968 (N_9968,N_9872,N_9883);
xnor U9969 (N_9969,N_9807,N_9813);
nand U9970 (N_9970,N_9818,N_9857);
xor U9971 (N_9971,N_9839,N_9887);
xor U9972 (N_9972,N_9805,N_9801);
or U9973 (N_9973,N_9849,N_9858);
and U9974 (N_9974,N_9891,N_9877);
and U9975 (N_9975,N_9809,N_9843);
xor U9976 (N_9976,N_9819,N_9848);
xnor U9977 (N_9977,N_9816,N_9865);
xnor U9978 (N_9978,N_9882,N_9804);
xor U9979 (N_9979,N_9839,N_9807);
and U9980 (N_9980,N_9891,N_9802);
and U9981 (N_9981,N_9846,N_9862);
or U9982 (N_9982,N_9891,N_9871);
nand U9983 (N_9983,N_9862,N_9849);
xnor U9984 (N_9984,N_9801,N_9824);
nor U9985 (N_9985,N_9844,N_9883);
or U9986 (N_9986,N_9843,N_9838);
nor U9987 (N_9987,N_9835,N_9803);
and U9988 (N_9988,N_9873,N_9838);
nor U9989 (N_9989,N_9889,N_9896);
or U9990 (N_9990,N_9883,N_9870);
nand U9991 (N_9991,N_9814,N_9831);
or U9992 (N_9992,N_9872,N_9838);
nand U9993 (N_9993,N_9878,N_9860);
or U9994 (N_9994,N_9805,N_9882);
xnor U9995 (N_9995,N_9833,N_9867);
nor U9996 (N_9996,N_9866,N_9837);
xor U9997 (N_9997,N_9875,N_9895);
nand U9998 (N_9998,N_9803,N_9846);
or U9999 (N_9999,N_9883,N_9831);
nor UO_0 (O_0,N_9942,N_9965);
and UO_1 (O_1,N_9915,N_9906);
nor UO_2 (O_2,N_9931,N_9909);
nand UO_3 (O_3,N_9975,N_9968);
xor UO_4 (O_4,N_9980,N_9984);
nor UO_5 (O_5,N_9918,N_9916);
and UO_6 (O_6,N_9903,N_9920);
or UO_7 (O_7,N_9921,N_9993);
nand UO_8 (O_8,N_9914,N_9939);
xnor UO_9 (O_9,N_9979,N_9971);
nand UO_10 (O_10,N_9977,N_9901);
and UO_11 (O_11,N_9961,N_9923);
xor UO_12 (O_12,N_9996,N_9994);
or UO_13 (O_13,N_9933,N_9960);
and UO_14 (O_14,N_9982,N_9998);
xnor UO_15 (O_15,N_9951,N_9922);
and UO_16 (O_16,N_9997,N_9929);
or UO_17 (O_17,N_9970,N_9955);
or UO_18 (O_18,N_9944,N_9950);
xor UO_19 (O_19,N_9981,N_9983);
or UO_20 (O_20,N_9926,N_9917);
nor UO_21 (O_21,N_9969,N_9935);
nor UO_22 (O_22,N_9930,N_9947);
nand UO_23 (O_23,N_9928,N_9927);
nand UO_24 (O_24,N_9952,N_9966);
xor UO_25 (O_25,N_9940,N_9904);
nor UO_26 (O_26,N_9924,N_9938);
nor UO_27 (O_27,N_9934,N_9958);
xor UO_28 (O_28,N_9956,N_9954);
nand UO_29 (O_29,N_9973,N_9925);
xnor UO_30 (O_30,N_9919,N_9987);
or UO_31 (O_31,N_9963,N_9905);
and UO_32 (O_32,N_9949,N_9957);
xor UO_33 (O_33,N_9988,N_9912);
nand UO_34 (O_34,N_9999,N_9976);
nand UO_35 (O_35,N_9953,N_9907);
xor UO_36 (O_36,N_9941,N_9974);
or UO_37 (O_37,N_9972,N_9962);
xor UO_38 (O_38,N_9986,N_9989);
or UO_39 (O_39,N_9937,N_9995);
xnor UO_40 (O_40,N_9932,N_9908);
nand UO_41 (O_41,N_9913,N_9967);
xor UO_42 (O_42,N_9948,N_9945);
nand UO_43 (O_43,N_9992,N_9959);
nor UO_44 (O_44,N_9936,N_9900);
xnor UO_45 (O_45,N_9985,N_9943);
or UO_46 (O_46,N_9964,N_9910);
or UO_47 (O_47,N_9978,N_9911);
nor UO_48 (O_48,N_9991,N_9990);
nand UO_49 (O_49,N_9946,N_9902);
nor UO_50 (O_50,N_9942,N_9997);
nand UO_51 (O_51,N_9947,N_9958);
nor UO_52 (O_52,N_9940,N_9982);
or UO_53 (O_53,N_9954,N_9953);
or UO_54 (O_54,N_9933,N_9942);
nand UO_55 (O_55,N_9935,N_9966);
nand UO_56 (O_56,N_9958,N_9909);
nor UO_57 (O_57,N_9911,N_9983);
xor UO_58 (O_58,N_9976,N_9997);
or UO_59 (O_59,N_9936,N_9988);
nand UO_60 (O_60,N_9945,N_9962);
and UO_61 (O_61,N_9984,N_9983);
and UO_62 (O_62,N_9995,N_9941);
and UO_63 (O_63,N_9994,N_9922);
xnor UO_64 (O_64,N_9974,N_9967);
xnor UO_65 (O_65,N_9938,N_9949);
nand UO_66 (O_66,N_9932,N_9915);
and UO_67 (O_67,N_9954,N_9966);
or UO_68 (O_68,N_9952,N_9981);
nand UO_69 (O_69,N_9951,N_9934);
xnor UO_70 (O_70,N_9930,N_9941);
nor UO_71 (O_71,N_9904,N_9912);
nand UO_72 (O_72,N_9998,N_9919);
xnor UO_73 (O_73,N_9930,N_9966);
nand UO_74 (O_74,N_9952,N_9964);
or UO_75 (O_75,N_9962,N_9997);
nor UO_76 (O_76,N_9997,N_9901);
nor UO_77 (O_77,N_9940,N_9903);
nor UO_78 (O_78,N_9988,N_9946);
xor UO_79 (O_79,N_9995,N_9975);
xnor UO_80 (O_80,N_9949,N_9926);
and UO_81 (O_81,N_9923,N_9917);
nand UO_82 (O_82,N_9968,N_9907);
or UO_83 (O_83,N_9956,N_9929);
nor UO_84 (O_84,N_9920,N_9945);
nand UO_85 (O_85,N_9964,N_9946);
and UO_86 (O_86,N_9924,N_9952);
nor UO_87 (O_87,N_9906,N_9950);
or UO_88 (O_88,N_9971,N_9986);
nor UO_89 (O_89,N_9956,N_9937);
and UO_90 (O_90,N_9934,N_9902);
nor UO_91 (O_91,N_9910,N_9987);
nand UO_92 (O_92,N_9982,N_9964);
xnor UO_93 (O_93,N_9943,N_9971);
and UO_94 (O_94,N_9909,N_9927);
or UO_95 (O_95,N_9945,N_9931);
xor UO_96 (O_96,N_9934,N_9979);
xor UO_97 (O_97,N_9965,N_9982);
and UO_98 (O_98,N_9937,N_9994);
nand UO_99 (O_99,N_9906,N_9957);
nand UO_100 (O_100,N_9926,N_9916);
xor UO_101 (O_101,N_9927,N_9908);
and UO_102 (O_102,N_9979,N_9973);
nand UO_103 (O_103,N_9928,N_9965);
or UO_104 (O_104,N_9920,N_9958);
nor UO_105 (O_105,N_9900,N_9948);
and UO_106 (O_106,N_9995,N_9964);
xor UO_107 (O_107,N_9964,N_9948);
and UO_108 (O_108,N_9963,N_9935);
and UO_109 (O_109,N_9928,N_9959);
or UO_110 (O_110,N_9956,N_9905);
nor UO_111 (O_111,N_9909,N_9914);
or UO_112 (O_112,N_9997,N_9969);
and UO_113 (O_113,N_9971,N_9999);
or UO_114 (O_114,N_9904,N_9956);
and UO_115 (O_115,N_9927,N_9944);
nand UO_116 (O_116,N_9976,N_9985);
nor UO_117 (O_117,N_9902,N_9924);
or UO_118 (O_118,N_9930,N_9979);
nand UO_119 (O_119,N_9932,N_9937);
and UO_120 (O_120,N_9964,N_9963);
xnor UO_121 (O_121,N_9933,N_9902);
nor UO_122 (O_122,N_9988,N_9915);
xor UO_123 (O_123,N_9954,N_9980);
nor UO_124 (O_124,N_9905,N_9926);
nor UO_125 (O_125,N_9930,N_9901);
and UO_126 (O_126,N_9931,N_9975);
or UO_127 (O_127,N_9946,N_9905);
nor UO_128 (O_128,N_9904,N_9938);
nand UO_129 (O_129,N_9991,N_9986);
nor UO_130 (O_130,N_9962,N_9913);
or UO_131 (O_131,N_9955,N_9984);
nor UO_132 (O_132,N_9917,N_9990);
xor UO_133 (O_133,N_9959,N_9918);
or UO_134 (O_134,N_9921,N_9962);
or UO_135 (O_135,N_9979,N_9933);
xor UO_136 (O_136,N_9990,N_9905);
nand UO_137 (O_137,N_9908,N_9942);
xor UO_138 (O_138,N_9961,N_9985);
and UO_139 (O_139,N_9970,N_9904);
nor UO_140 (O_140,N_9923,N_9921);
xor UO_141 (O_141,N_9942,N_9981);
or UO_142 (O_142,N_9956,N_9917);
nand UO_143 (O_143,N_9904,N_9954);
nand UO_144 (O_144,N_9985,N_9975);
xnor UO_145 (O_145,N_9981,N_9951);
nand UO_146 (O_146,N_9958,N_9985);
and UO_147 (O_147,N_9914,N_9931);
or UO_148 (O_148,N_9961,N_9980);
nor UO_149 (O_149,N_9966,N_9932);
or UO_150 (O_150,N_9925,N_9929);
nand UO_151 (O_151,N_9959,N_9940);
or UO_152 (O_152,N_9906,N_9947);
xnor UO_153 (O_153,N_9998,N_9928);
nor UO_154 (O_154,N_9988,N_9965);
xnor UO_155 (O_155,N_9947,N_9997);
xnor UO_156 (O_156,N_9925,N_9926);
xor UO_157 (O_157,N_9951,N_9910);
xnor UO_158 (O_158,N_9992,N_9970);
or UO_159 (O_159,N_9924,N_9910);
nand UO_160 (O_160,N_9962,N_9949);
nor UO_161 (O_161,N_9959,N_9958);
nand UO_162 (O_162,N_9980,N_9938);
and UO_163 (O_163,N_9943,N_9953);
or UO_164 (O_164,N_9971,N_9921);
nand UO_165 (O_165,N_9974,N_9954);
and UO_166 (O_166,N_9916,N_9991);
and UO_167 (O_167,N_9982,N_9948);
and UO_168 (O_168,N_9905,N_9994);
and UO_169 (O_169,N_9929,N_9918);
or UO_170 (O_170,N_9990,N_9965);
xnor UO_171 (O_171,N_9953,N_9940);
or UO_172 (O_172,N_9983,N_9955);
and UO_173 (O_173,N_9944,N_9988);
xnor UO_174 (O_174,N_9916,N_9978);
xor UO_175 (O_175,N_9913,N_9964);
and UO_176 (O_176,N_9906,N_9916);
or UO_177 (O_177,N_9904,N_9910);
nor UO_178 (O_178,N_9936,N_9981);
nor UO_179 (O_179,N_9937,N_9900);
nor UO_180 (O_180,N_9950,N_9905);
nor UO_181 (O_181,N_9988,N_9955);
xnor UO_182 (O_182,N_9907,N_9960);
nand UO_183 (O_183,N_9975,N_9952);
and UO_184 (O_184,N_9989,N_9943);
and UO_185 (O_185,N_9929,N_9973);
nand UO_186 (O_186,N_9915,N_9939);
nor UO_187 (O_187,N_9961,N_9906);
and UO_188 (O_188,N_9984,N_9954);
or UO_189 (O_189,N_9953,N_9942);
nand UO_190 (O_190,N_9955,N_9998);
nor UO_191 (O_191,N_9960,N_9934);
nand UO_192 (O_192,N_9931,N_9906);
xor UO_193 (O_193,N_9927,N_9951);
xnor UO_194 (O_194,N_9971,N_9928);
nand UO_195 (O_195,N_9915,N_9920);
or UO_196 (O_196,N_9909,N_9956);
and UO_197 (O_197,N_9938,N_9906);
xnor UO_198 (O_198,N_9979,N_9957);
nand UO_199 (O_199,N_9963,N_9945);
xor UO_200 (O_200,N_9971,N_9982);
nand UO_201 (O_201,N_9924,N_9998);
nand UO_202 (O_202,N_9978,N_9921);
xor UO_203 (O_203,N_9966,N_9937);
xor UO_204 (O_204,N_9914,N_9950);
nor UO_205 (O_205,N_9983,N_9915);
nand UO_206 (O_206,N_9988,N_9992);
nand UO_207 (O_207,N_9996,N_9901);
nor UO_208 (O_208,N_9961,N_9929);
or UO_209 (O_209,N_9926,N_9959);
nand UO_210 (O_210,N_9905,N_9992);
nor UO_211 (O_211,N_9992,N_9922);
or UO_212 (O_212,N_9987,N_9995);
nor UO_213 (O_213,N_9966,N_9906);
nor UO_214 (O_214,N_9949,N_9922);
and UO_215 (O_215,N_9948,N_9975);
nor UO_216 (O_216,N_9955,N_9904);
nand UO_217 (O_217,N_9939,N_9952);
nor UO_218 (O_218,N_9920,N_9994);
xnor UO_219 (O_219,N_9943,N_9951);
nand UO_220 (O_220,N_9999,N_9945);
nor UO_221 (O_221,N_9914,N_9988);
and UO_222 (O_222,N_9996,N_9908);
and UO_223 (O_223,N_9959,N_9980);
or UO_224 (O_224,N_9989,N_9974);
or UO_225 (O_225,N_9979,N_9986);
or UO_226 (O_226,N_9994,N_9955);
or UO_227 (O_227,N_9945,N_9959);
nand UO_228 (O_228,N_9902,N_9978);
xnor UO_229 (O_229,N_9911,N_9913);
nand UO_230 (O_230,N_9920,N_9995);
nor UO_231 (O_231,N_9990,N_9902);
or UO_232 (O_232,N_9968,N_9914);
xnor UO_233 (O_233,N_9918,N_9995);
or UO_234 (O_234,N_9973,N_9912);
and UO_235 (O_235,N_9945,N_9980);
or UO_236 (O_236,N_9999,N_9924);
nor UO_237 (O_237,N_9902,N_9943);
or UO_238 (O_238,N_9960,N_9958);
xnor UO_239 (O_239,N_9919,N_9941);
nand UO_240 (O_240,N_9988,N_9958);
xor UO_241 (O_241,N_9944,N_9924);
nand UO_242 (O_242,N_9985,N_9928);
xnor UO_243 (O_243,N_9975,N_9960);
nor UO_244 (O_244,N_9984,N_9971);
and UO_245 (O_245,N_9956,N_9977);
or UO_246 (O_246,N_9985,N_9944);
nor UO_247 (O_247,N_9976,N_9974);
or UO_248 (O_248,N_9950,N_9928);
and UO_249 (O_249,N_9984,N_9966);
or UO_250 (O_250,N_9908,N_9959);
nor UO_251 (O_251,N_9977,N_9929);
and UO_252 (O_252,N_9974,N_9931);
or UO_253 (O_253,N_9901,N_9916);
xor UO_254 (O_254,N_9944,N_9923);
nand UO_255 (O_255,N_9975,N_9951);
and UO_256 (O_256,N_9970,N_9905);
and UO_257 (O_257,N_9941,N_9988);
and UO_258 (O_258,N_9920,N_9904);
or UO_259 (O_259,N_9954,N_9911);
and UO_260 (O_260,N_9944,N_9994);
and UO_261 (O_261,N_9930,N_9997);
nand UO_262 (O_262,N_9968,N_9998);
nand UO_263 (O_263,N_9902,N_9948);
or UO_264 (O_264,N_9952,N_9957);
xor UO_265 (O_265,N_9965,N_9926);
xor UO_266 (O_266,N_9980,N_9970);
nor UO_267 (O_267,N_9936,N_9963);
nor UO_268 (O_268,N_9960,N_9908);
xnor UO_269 (O_269,N_9987,N_9992);
nor UO_270 (O_270,N_9930,N_9971);
nor UO_271 (O_271,N_9920,N_9951);
and UO_272 (O_272,N_9985,N_9935);
or UO_273 (O_273,N_9911,N_9982);
xor UO_274 (O_274,N_9931,N_9956);
and UO_275 (O_275,N_9957,N_9983);
and UO_276 (O_276,N_9939,N_9959);
nand UO_277 (O_277,N_9907,N_9959);
xnor UO_278 (O_278,N_9925,N_9932);
nand UO_279 (O_279,N_9991,N_9909);
nor UO_280 (O_280,N_9997,N_9934);
xnor UO_281 (O_281,N_9911,N_9953);
xnor UO_282 (O_282,N_9950,N_9980);
nand UO_283 (O_283,N_9967,N_9912);
and UO_284 (O_284,N_9922,N_9903);
and UO_285 (O_285,N_9935,N_9956);
nor UO_286 (O_286,N_9969,N_9963);
or UO_287 (O_287,N_9933,N_9971);
or UO_288 (O_288,N_9993,N_9954);
or UO_289 (O_289,N_9907,N_9987);
and UO_290 (O_290,N_9923,N_9918);
nor UO_291 (O_291,N_9927,N_9987);
xor UO_292 (O_292,N_9975,N_9930);
nor UO_293 (O_293,N_9984,N_9981);
nand UO_294 (O_294,N_9927,N_9968);
or UO_295 (O_295,N_9944,N_9997);
and UO_296 (O_296,N_9905,N_9988);
xor UO_297 (O_297,N_9900,N_9978);
nor UO_298 (O_298,N_9935,N_9955);
or UO_299 (O_299,N_9949,N_9944);
and UO_300 (O_300,N_9906,N_9904);
nor UO_301 (O_301,N_9909,N_9911);
nor UO_302 (O_302,N_9997,N_9987);
and UO_303 (O_303,N_9997,N_9964);
xnor UO_304 (O_304,N_9958,N_9948);
xnor UO_305 (O_305,N_9942,N_9987);
or UO_306 (O_306,N_9983,N_9989);
nor UO_307 (O_307,N_9914,N_9943);
and UO_308 (O_308,N_9955,N_9964);
and UO_309 (O_309,N_9935,N_9930);
or UO_310 (O_310,N_9943,N_9922);
nor UO_311 (O_311,N_9921,N_9902);
and UO_312 (O_312,N_9944,N_9965);
nor UO_313 (O_313,N_9959,N_9929);
nand UO_314 (O_314,N_9992,N_9909);
nand UO_315 (O_315,N_9918,N_9919);
and UO_316 (O_316,N_9997,N_9985);
nor UO_317 (O_317,N_9982,N_9946);
and UO_318 (O_318,N_9961,N_9978);
xnor UO_319 (O_319,N_9999,N_9981);
xor UO_320 (O_320,N_9955,N_9985);
or UO_321 (O_321,N_9939,N_9944);
xnor UO_322 (O_322,N_9943,N_9950);
and UO_323 (O_323,N_9945,N_9995);
or UO_324 (O_324,N_9956,N_9974);
nand UO_325 (O_325,N_9936,N_9938);
nand UO_326 (O_326,N_9934,N_9909);
nand UO_327 (O_327,N_9976,N_9900);
xnor UO_328 (O_328,N_9908,N_9987);
nand UO_329 (O_329,N_9922,N_9967);
xnor UO_330 (O_330,N_9937,N_9993);
nor UO_331 (O_331,N_9902,N_9953);
and UO_332 (O_332,N_9930,N_9991);
xor UO_333 (O_333,N_9926,N_9975);
nand UO_334 (O_334,N_9928,N_9978);
xnor UO_335 (O_335,N_9964,N_9993);
nor UO_336 (O_336,N_9906,N_9984);
or UO_337 (O_337,N_9937,N_9933);
and UO_338 (O_338,N_9920,N_9962);
nor UO_339 (O_339,N_9991,N_9949);
nand UO_340 (O_340,N_9921,N_9975);
and UO_341 (O_341,N_9981,N_9994);
nand UO_342 (O_342,N_9910,N_9991);
or UO_343 (O_343,N_9958,N_9929);
and UO_344 (O_344,N_9932,N_9912);
nand UO_345 (O_345,N_9942,N_9928);
nor UO_346 (O_346,N_9926,N_9924);
nor UO_347 (O_347,N_9986,N_9975);
xor UO_348 (O_348,N_9994,N_9906);
and UO_349 (O_349,N_9999,N_9954);
and UO_350 (O_350,N_9996,N_9961);
nor UO_351 (O_351,N_9987,N_9921);
or UO_352 (O_352,N_9950,N_9999);
nand UO_353 (O_353,N_9937,N_9914);
nor UO_354 (O_354,N_9980,N_9916);
xor UO_355 (O_355,N_9971,N_9996);
xor UO_356 (O_356,N_9924,N_9937);
xor UO_357 (O_357,N_9920,N_9919);
or UO_358 (O_358,N_9924,N_9912);
nand UO_359 (O_359,N_9946,N_9924);
or UO_360 (O_360,N_9910,N_9919);
and UO_361 (O_361,N_9912,N_9902);
nor UO_362 (O_362,N_9974,N_9965);
or UO_363 (O_363,N_9920,N_9999);
and UO_364 (O_364,N_9973,N_9971);
and UO_365 (O_365,N_9942,N_9970);
and UO_366 (O_366,N_9928,N_9999);
nand UO_367 (O_367,N_9938,N_9934);
and UO_368 (O_368,N_9966,N_9959);
xor UO_369 (O_369,N_9977,N_9955);
nor UO_370 (O_370,N_9990,N_9939);
nand UO_371 (O_371,N_9988,N_9931);
nor UO_372 (O_372,N_9978,N_9925);
xnor UO_373 (O_373,N_9996,N_9922);
nand UO_374 (O_374,N_9944,N_9955);
or UO_375 (O_375,N_9947,N_9955);
nand UO_376 (O_376,N_9938,N_9905);
nand UO_377 (O_377,N_9946,N_9972);
and UO_378 (O_378,N_9972,N_9951);
nand UO_379 (O_379,N_9943,N_9991);
nor UO_380 (O_380,N_9983,N_9918);
nor UO_381 (O_381,N_9985,N_9917);
and UO_382 (O_382,N_9909,N_9955);
nor UO_383 (O_383,N_9921,N_9907);
nand UO_384 (O_384,N_9927,N_9958);
or UO_385 (O_385,N_9975,N_9961);
xor UO_386 (O_386,N_9956,N_9933);
nand UO_387 (O_387,N_9998,N_9977);
and UO_388 (O_388,N_9981,N_9964);
and UO_389 (O_389,N_9924,N_9931);
nand UO_390 (O_390,N_9991,N_9933);
nand UO_391 (O_391,N_9939,N_9927);
nand UO_392 (O_392,N_9913,N_9981);
and UO_393 (O_393,N_9914,N_9965);
and UO_394 (O_394,N_9963,N_9929);
nand UO_395 (O_395,N_9971,N_9903);
nand UO_396 (O_396,N_9960,N_9997);
xor UO_397 (O_397,N_9954,N_9948);
and UO_398 (O_398,N_9984,N_9913);
nor UO_399 (O_399,N_9915,N_9992);
or UO_400 (O_400,N_9987,N_9912);
nor UO_401 (O_401,N_9903,N_9992);
nor UO_402 (O_402,N_9976,N_9956);
and UO_403 (O_403,N_9991,N_9950);
nand UO_404 (O_404,N_9944,N_9982);
nand UO_405 (O_405,N_9982,N_9984);
and UO_406 (O_406,N_9939,N_9933);
xor UO_407 (O_407,N_9961,N_9900);
nand UO_408 (O_408,N_9924,N_9989);
xor UO_409 (O_409,N_9973,N_9900);
nor UO_410 (O_410,N_9914,N_9901);
xor UO_411 (O_411,N_9935,N_9942);
nand UO_412 (O_412,N_9987,N_9974);
or UO_413 (O_413,N_9933,N_9929);
nor UO_414 (O_414,N_9905,N_9969);
xnor UO_415 (O_415,N_9930,N_9915);
xor UO_416 (O_416,N_9972,N_9992);
and UO_417 (O_417,N_9907,N_9997);
and UO_418 (O_418,N_9971,N_9992);
nor UO_419 (O_419,N_9938,N_9951);
or UO_420 (O_420,N_9977,N_9991);
nand UO_421 (O_421,N_9927,N_9907);
nor UO_422 (O_422,N_9947,N_9987);
xor UO_423 (O_423,N_9983,N_9972);
and UO_424 (O_424,N_9922,N_9923);
or UO_425 (O_425,N_9957,N_9951);
xnor UO_426 (O_426,N_9901,N_9987);
or UO_427 (O_427,N_9992,N_9974);
xnor UO_428 (O_428,N_9969,N_9971);
or UO_429 (O_429,N_9941,N_9961);
xnor UO_430 (O_430,N_9904,N_9947);
xor UO_431 (O_431,N_9976,N_9931);
nand UO_432 (O_432,N_9931,N_9905);
nor UO_433 (O_433,N_9995,N_9954);
nand UO_434 (O_434,N_9930,N_9992);
nor UO_435 (O_435,N_9997,N_9980);
nand UO_436 (O_436,N_9903,N_9932);
and UO_437 (O_437,N_9989,N_9994);
and UO_438 (O_438,N_9971,N_9953);
xor UO_439 (O_439,N_9945,N_9918);
and UO_440 (O_440,N_9921,N_9982);
nor UO_441 (O_441,N_9932,N_9961);
xnor UO_442 (O_442,N_9973,N_9938);
xnor UO_443 (O_443,N_9913,N_9952);
or UO_444 (O_444,N_9988,N_9991);
xnor UO_445 (O_445,N_9915,N_9944);
nand UO_446 (O_446,N_9920,N_9987);
nand UO_447 (O_447,N_9997,N_9968);
nand UO_448 (O_448,N_9950,N_9941);
nor UO_449 (O_449,N_9903,N_9961);
xor UO_450 (O_450,N_9926,N_9941);
nand UO_451 (O_451,N_9986,N_9999);
nor UO_452 (O_452,N_9976,N_9906);
nor UO_453 (O_453,N_9979,N_9968);
or UO_454 (O_454,N_9960,N_9994);
nand UO_455 (O_455,N_9983,N_9917);
nor UO_456 (O_456,N_9949,N_9990);
xor UO_457 (O_457,N_9941,N_9929);
and UO_458 (O_458,N_9959,N_9969);
or UO_459 (O_459,N_9981,N_9929);
xnor UO_460 (O_460,N_9903,N_9908);
and UO_461 (O_461,N_9904,N_9949);
and UO_462 (O_462,N_9953,N_9926);
and UO_463 (O_463,N_9970,N_9964);
nor UO_464 (O_464,N_9930,N_9904);
and UO_465 (O_465,N_9930,N_9917);
nor UO_466 (O_466,N_9993,N_9931);
nor UO_467 (O_467,N_9970,N_9968);
nand UO_468 (O_468,N_9970,N_9930);
xor UO_469 (O_469,N_9919,N_9973);
and UO_470 (O_470,N_9912,N_9903);
nand UO_471 (O_471,N_9933,N_9911);
nand UO_472 (O_472,N_9935,N_9909);
xnor UO_473 (O_473,N_9999,N_9992);
nor UO_474 (O_474,N_9903,N_9999);
nor UO_475 (O_475,N_9910,N_9990);
and UO_476 (O_476,N_9972,N_9986);
nand UO_477 (O_477,N_9955,N_9946);
and UO_478 (O_478,N_9972,N_9909);
xor UO_479 (O_479,N_9932,N_9985);
and UO_480 (O_480,N_9990,N_9985);
nand UO_481 (O_481,N_9902,N_9988);
nand UO_482 (O_482,N_9981,N_9934);
xnor UO_483 (O_483,N_9954,N_9936);
and UO_484 (O_484,N_9902,N_9941);
nand UO_485 (O_485,N_9940,N_9976);
and UO_486 (O_486,N_9961,N_9910);
nand UO_487 (O_487,N_9956,N_9992);
and UO_488 (O_488,N_9932,N_9994);
nor UO_489 (O_489,N_9960,N_9979);
xor UO_490 (O_490,N_9928,N_9920);
nor UO_491 (O_491,N_9987,N_9961);
xnor UO_492 (O_492,N_9923,N_9992);
xnor UO_493 (O_493,N_9958,N_9924);
or UO_494 (O_494,N_9929,N_9917);
nor UO_495 (O_495,N_9926,N_9904);
nand UO_496 (O_496,N_9983,N_9937);
xnor UO_497 (O_497,N_9931,N_9907);
xor UO_498 (O_498,N_9988,N_9984);
xnor UO_499 (O_499,N_9982,N_9919);
or UO_500 (O_500,N_9957,N_9934);
or UO_501 (O_501,N_9921,N_9928);
nand UO_502 (O_502,N_9971,N_9913);
nand UO_503 (O_503,N_9901,N_9955);
nor UO_504 (O_504,N_9938,N_9921);
or UO_505 (O_505,N_9936,N_9994);
nor UO_506 (O_506,N_9986,N_9903);
xor UO_507 (O_507,N_9935,N_9983);
nor UO_508 (O_508,N_9946,N_9913);
xor UO_509 (O_509,N_9981,N_9973);
nand UO_510 (O_510,N_9933,N_9909);
nand UO_511 (O_511,N_9938,N_9991);
and UO_512 (O_512,N_9984,N_9991);
and UO_513 (O_513,N_9958,N_9978);
nand UO_514 (O_514,N_9925,N_9986);
nand UO_515 (O_515,N_9982,N_9914);
xnor UO_516 (O_516,N_9947,N_9945);
xor UO_517 (O_517,N_9928,N_9917);
or UO_518 (O_518,N_9957,N_9956);
nor UO_519 (O_519,N_9907,N_9985);
or UO_520 (O_520,N_9900,N_9993);
and UO_521 (O_521,N_9979,N_9980);
or UO_522 (O_522,N_9989,N_9952);
nor UO_523 (O_523,N_9901,N_9941);
or UO_524 (O_524,N_9984,N_9962);
nor UO_525 (O_525,N_9947,N_9932);
xor UO_526 (O_526,N_9952,N_9978);
nand UO_527 (O_527,N_9915,N_9978);
nand UO_528 (O_528,N_9997,N_9935);
and UO_529 (O_529,N_9963,N_9980);
and UO_530 (O_530,N_9963,N_9989);
xor UO_531 (O_531,N_9920,N_9980);
nand UO_532 (O_532,N_9901,N_9956);
or UO_533 (O_533,N_9939,N_9958);
nor UO_534 (O_534,N_9940,N_9991);
and UO_535 (O_535,N_9975,N_9953);
or UO_536 (O_536,N_9984,N_9908);
or UO_537 (O_537,N_9937,N_9991);
xor UO_538 (O_538,N_9944,N_9974);
xnor UO_539 (O_539,N_9975,N_9902);
or UO_540 (O_540,N_9943,N_9910);
nand UO_541 (O_541,N_9996,N_9931);
and UO_542 (O_542,N_9955,N_9902);
xnor UO_543 (O_543,N_9930,N_9946);
or UO_544 (O_544,N_9906,N_9986);
nor UO_545 (O_545,N_9943,N_9984);
and UO_546 (O_546,N_9941,N_9946);
or UO_547 (O_547,N_9982,N_9933);
or UO_548 (O_548,N_9956,N_9941);
nor UO_549 (O_549,N_9947,N_9909);
and UO_550 (O_550,N_9979,N_9913);
and UO_551 (O_551,N_9903,N_9959);
xnor UO_552 (O_552,N_9903,N_9924);
or UO_553 (O_553,N_9917,N_9999);
and UO_554 (O_554,N_9909,N_9941);
nand UO_555 (O_555,N_9927,N_9900);
xnor UO_556 (O_556,N_9904,N_9941);
nand UO_557 (O_557,N_9957,N_9901);
or UO_558 (O_558,N_9908,N_9905);
xnor UO_559 (O_559,N_9986,N_9998);
nand UO_560 (O_560,N_9989,N_9941);
xor UO_561 (O_561,N_9955,N_9930);
nand UO_562 (O_562,N_9943,N_9964);
nor UO_563 (O_563,N_9916,N_9946);
and UO_564 (O_564,N_9998,N_9943);
and UO_565 (O_565,N_9918,N_9965);
nand UO_566 (O_566,N_9901,N_9921);
or UO_567 (O_567,N_9920,N_9944);
nor UO_568 (O_568,N_9946,N_9908);
nor UO_569 (O_569,N_9903,N_9974);
nor UO_570 (O_570,N_9944,N_9999);
xor UO_571 (O_571,N_9903,N_9964);
or UO_572 (O_572,N_9996,N_9935);
xnor UO_573 (O_573,N_9911,N_9991);
nand UO_574 (O_574,N_9948,N_9946);
nor UO_575 (O_575,N_9981,N_9995);
nand UO_576 (O_576,N_9967,N_9955);
nor UO_577 (O_577,N_9963,N_9924);
nand UO_578 (O_578,N_9908,N_9998);
and UO_579 (O_579,N_9921,N_9930);
nand UO_580 (O_580,N_9912,N_9972);
xnor UO_581 (O_581,N_9966,N_9947);
nor UO_582 (O_582,N_9942,N_9922);
xor UO_583 (O_583,N_9953,N_9905);
nor UO_584 (O_584,N_9940,N_9916);
nand UO_585 (O_585,N_9932,N_9990);
or UO_586 (O_586,N_9950,N_9939);
or UO_587 (O_587,N_9962,N_9947);
nand UO_588 (O_588,N_9935,N_9964);
xor UO_589 (O_589,N_9951,N_9916);
or UO_590 (O_590,N_9982,N_9968);
or UO_591 (O_591,N_9926,N_9955);
nor UO_592 (O_592,N_9926,N_9943);
and UO_593 (O_593,N_9924,N_9933);
nand UO_594 (O_594,N_9958,N_9942);
or UO_595 (O_595,N_9991,N_9970);
nand UO_596 (O_596,N_9985,N_9942);
nand UO_597 (O_597,N_9949,N_9936);
and UO_598 (O_598,N_9988,N_9996);
xnor UO_599 (O_599,N_9946,N_9996);
and UO_600 (O_600,N_9947,N_9905);
or UO_601 (O_601,N_9993,N_9918);
xnor UO_602 (O_602,N_9945,N_9900);
or UO_603 (O_603,N_9985,N_9938);
and UO_604 (O_604,N_9981,N_9974);
nor UO_605 (O_605,N_9927,N_9962);
nor UO_606 (O_606,N_9953,N_9978);
or UO_607 (O_607,N_9912,N_9901);
xor UO_608 (O_608,N_9943,N_9930);
or UO_609 (O_609,N_9949,N_9987);
nand UO_610 (O_610,N_9911,N_9930);
xor UO_611 (O_611,N_9949,N_9947);
xnor UO_612 (O_612,N_9919,N_9923);
xor UO_613 (O_613,N_9996,N_9990);
or UO_614 (O_614,N_9986,N_9933);
nor UO_615 (O_615,N_9983,N_9996);
and UO_616 (O_616,N_9975,N_9958);
or UO_617 (O_617,N_9939,N_9960);
xnor UO_618 (O_618,N_9971,N_9922);
nand UO_619 (O_619,N_9947,N_9908);
and UO_620 (O_620,N_9905,N_9918);
nand UO_621 (O_621,N_9962,N_9942);
nand UO_622 (O_622,N_9996,N_9982);
or UO_623 (O_623,N_9961,N_9953);
and UO_624 (O_624,N_9915,N_9985);
xnor UO_625 (O_625,N_9903,N_9929);
nor UO_626 (O_626,N_9973,N_9990);
or UO_627 (O_627,N_9956,N_9908);
xor UO_628 (O_628,N_9999,N_9988);
xor UO_629 (O_629,N_9979,N_9953);
nand UO_630 (O_630,N_9968,N_9925);
xnor UO_631 (O_631,N_9915,N_9955);
nor UO_632 (O_632,N_9994,N_9943);
or UO_633 (O_633,N_9907,N_9989);
xor UO_634 (O_634,N_9907,N_9947);
nand UO_635 (O_635,N_9953,N_9935);
and UO_636 (O_636,N_9983,N_9995);
or UO_637 (O_637,N_9993,N_9971);
or UO_638 (O_638,N_9949,N_9929);
or UO_639 (O_639,N_9922,N_9939);
and UO_640 (O_640,N_9973,N_9977);
nor UO_641 (O_641,N_9904,N_9975);
and UO_642 (O_642,N_9919,N_9948);
and UO_643 (O_643,N_9926,N_9993);
and UO_644 (O_644,N_9937,N_9963);
nand UO_645 (O_645,N_9982,N_9994);
nand UO_646 (O_646,N_9963,N_9944);
xor UO_647 (O_647,N_9900,N_9966);
nor UO_648 (O_648,N_9981,N_9924);
or UO_649 (O_649,N_9936,N_9901);
nor UO_650 (O_650,N_9945,N_9992);
or UO_651 (O_651,N_9973,N_9902);
nand UO_652 (O_652,N_9935,N_9945);
or UO_653 (O_653,N_9973,N_9969);
and UO_654 (O_654,N_9986,N_9940);
nor UO_655 (O_655,N_9926,N_9910);
nor UO_656 (O_656,N_9907,N_9986);
and UO_657 (O_657,N_9958,N_9991);
xor UO_658 (O_658,N_9979,N_9948);
or UO_659 (O_659,N_9995,N_9926);
and UO_660 (O_660,N_9944,N_9937);
or UO_661 (O_661,N_9932,N_9962);
and UO_662 (O_662,N_9904,N_9945);
nand UO_663 (O_663,N_9979,N_9938);
or UO_664 (O_664,N_9946,N_9993);
or UO_665 (O_665,N_9929,N_9990);
xnor UO_666 (O_666,N_9909,N_9952);
or UO_667 (O_667,N_9973,N_9980);
and UO_668 (O_668,N_9977,N_9937);
and UO_669 (O_669,N_9945,N_9957);
nand UO_670 (O_670,N_9974,N_9935);
nand UO_671 (O_671,N_9977,N_9915);
nand UO_672 (O_672,N_9960,N_9944);
nand UO_673 (O_673,N_9989,N_9960);
or UO_674 (O_674,N_9983,N_9946);
or UO_675 (O_675,N_9946,N_9997);
nor UO_676 (O_676,N_9927,N_9931);
or UO_677 (O_677,N_9976,N_9909);
nor UO_678 (O_678,N_9947,N_9925);
xnor UO_679 (O_679,N_9902,N_9995);
and UO_680 (O_680,N_9977,N_9976);
or UO_681 (O_681,N_9983,N_9906);
xor UO_682 (O_682,N_9911,N_9975);
and UO_683 (O_683,N_9917,N_9980);
nor UO_684 (O_684,N_9960,N_9971);
nand UO_685 (O_685,N_9900,N_9935);
and UO_686 (O_686,N_9904,N_9917);
nand UO_687 (O_687,N_9901,N_9943);
xor UO_688 (O_688,N_9942,N_9927);
nor UO_689 (O_689,N_9908,N_9989);
and UO_690 (O_690,N_9997,N_9936);
xor UO_691 (O_691,N_9934,N_9929);
xnor UO_692 (O_692,N_9998,N_9969);
nor UO_693 (O_693,N_9910,N_9978);
and UO_694 (O_694,N_9934,N_9953);
nor UO_695 (O_695,N_9941,N_9925);
and UO_696 (O_696,N_9978,N_9931);
xor UO_697 (O_697,N_9930,N_9989);
and UO_698 (O_698,N_9911,N_9970);
nand UO_699 (O_699,N_9927,N_9956);
nand UO_700 (O_700,N_9953,N_9924);
nor UO_701 (O_701,N_9906,N_9929);
xnor UO_702 (O_702,N_9945,N_9988);
nand UO_703 (O_703,N_9912,N_9970);
and UO_704 (O_704,N_9930,N_9944);
and UO_705 (O_705,N_9950,N_9973);
nor UO_706 (O_706,N_9919,N_9957);
nor UO_707 (O_707,N_9924,N_9930);
and UO_708 (O_708,N_9956,N_9907);
xnor UO_709 (O_709,N_9972,N_9931);
and UO_710 (O_710,N_9985,N_9941);
nand UO_711 (O_711,N_9922,N_9975);
and UO_712 (O_712,N_9994,N_9913);
and UO_713 (O_713,N_9984,N_9945);
nand UO_714 (O_714,N_9973,N_9921);
and UO_715 (O_715,N_9956,N_9946);
nor UO_716 (O_716,N_9949,N_9964);
nor UO_717 (O_717,N_9957,N_9902);
nor UO_718 (O_718,N_9932,N_9924);
or UO_719 (O_719,N_9941,N_9951);
or UO_720 (O_720,N_9900,N_9979);
nor UO_721 (O_721,N_9909,N_9985);
nor UO_722 (O_722,N_9914,N_9933);
xor UO_723 (O_723,N_9902,N_9985);
and UO_724 (O_724,N_9944,N_9919);
xnor UO_725 (O_725,N_9926,N_9902);
nor UO_726 (O_726,N_9930,N_9995);
and UO_727 (O_727,N_9937,N_9903);
nand UO_728 (O_728,N_9908,N_9931);
nand UO_729 (O_729,N_9903,N_9931);
and UO_730 (O_730,N_9967,N_9900);
nand UO_731 (O_731,N_9956,N_9939);
nor UO_732 (O_732,N_9925,N_9922);
nor UO_733 (O_733,N_9949,N_9915);
or UO_734 (O_734,N_9909,N_9900);
or UO_735 (O_735,N_9941,N_9993);
nand UO_736 (O_736,N_9933,N_9900);
or UO_737 (O_737,N_9934,N_9900);
nor UO_738 (O_738,N_9915,N_9976);
nand UO_739 (O_739,N_9928,N_9991);
or UO_740 (O_740,N_9901,N_9954);
and UO_741 (O_741,N_9972,N_9963);
or UO_742 (O_742,N_9929,N_9983);
nor UO_743 (O_743,N_9942,N_9915);
and UO_744 (O_744,N_9917,N_9900);
and UO_745 (O_745,N_9931,N_9932);
nor UO_746 (O_746,N_9944,N_9931);
or UO_747 (O_747,N_9971,N_9906);
nand UO_748 (O_748,N_9980,N_9903);
xnor UO_749 (O_749,N_9936,N_9980);
xnor UO_750 (O_750,N_9969,N_9961);
nor UO_751 (O_751,N_9901,N_9920);
nor UO_752 (O_752,N_9989,N_9945);
or UO_753 (O_753,N_9961,N_9944);
and UO_754 (O_754,N_9974,N_9947);
nor UO_755 (O_755,N_9964,N_9998);
or UO_756 (O_756,N_9915,N_9968);
nand UO_757 (O_757,N_9978,N_9949);
xnor UO_758 (O_758,N_9954,N_9968);
and UO_759 (O_759,N_9990,N_9955);
or UO_760 (O_760,N_9981,N_9906);
nor UO_761 (O_761,N_9908,N_9976);
and UO_762 (O_762,N_9954,N_9918);
or UO_763 (O_763,N_9973,N_9966);
and UO_764 (O_764,N_9923,N_9962);
nor UO_765 (O_765,N_9967,N_9942);
or UO_766 (O_766,N_9923,N_9951);
nor UO_767 (O_767,N_9911,N_9965);
or UO_768 (O_768,N_9999,N_9998);
and UO_769 (O_769,N_9981,N_9910);
or UO_770 (O_770,N_9933,N_9990);
or UO_771 (O_771,N_9985,N_9981);
nand UO_772 (O_772,N_9975,N_9912);
or UO_773 (O_773,N_9989,N_9922);
or UO_774 (O_774,N_9947,N_9937);
or UO_775 (O_775,N_9986,N_9942);
nor UO_776 (O_776,N_9972,N_9993);
nand UO_777 (O_777,N_9908,N_9924);
xnor UO_778 (O_778,N_9945,N_9960);
and UO_779 (O_779,N_9975,N_9916);
and UO_780 (O_780,N_9939,N_9930);
or UO_781 (O_781,N_9952,N_9986);
xnor UO_782 (O_782,N_9929,N_9939);
nor UO_783 (O_783,N_9985,N_9908);
and UO_784 (O_784,N_9989,N_9915);
or UO_785 (O_785,N_9930,N_9926);
xor UO_786 (O_786,N_9997,N_9949);
nor UO_787 (O_787,N_9907,N_9935);
or UO_788 (O_788,N_9954,N_9943);
nor UO_789 (O_789,N_9974,N_9993);
xor UO_790 (O_790,N_9956,N_9958);
and UO_791 (O_791,N_9950,N_9945);
xor UO_792 (O_792,N_9918,N_9989);
or UO_793 (O_793,N_9902,N_9916);
and UO_794 (O_794,N_9927,N_9964);
nor UO_795 (O_795,N_9928,N_9903);
nor UO_796 (O_796,N_9928,N_9955);
xor UO_797 (O_797,N_9915,N_9903);
nor UO_798 (O_798,N_9995,N_9906);
and UO_799 (O_799,N_9918,N_9909);
xor UO_800 (O_800,N_9917,N_9943);
nor UO_801 (O_801,N_9906,N_9943);
and UO_802 (O_802,N_9921,N_9986);
and UO_803 (O_803,N_9910,N_9977);
xnor UO_804 (O_804,N_9921,N_9988);
or UO_805 (O_805,N_9994,N_9970);
nand UO_806 (O_806,N_9969,N_9907);
or UO_807 (O_807,N_9912,N_9969);
nand UO_808 (O_808,N_9974,N_9900);
nand UO_809 (O_809,N_9913,N_9938);
xor UO_810 (O_810,N_9903,N_9913);
nor UO_811 (O_811,N_9916,N_9939);
nor UO_812 (O_812,N_9970,N_9959);
and UO_813 (O_813,N_9932,N_9965);
nor UO_814 (O_814,N_9911,N_9972);
nor UO_815 (O_815,N_9983,N_9959);
and UO_816 (O_816,N_9901,N_9951);
nand UO_817 (O_817,N_9991,N_9999);
nand UO_818 (O_818,N_9981,N_9921);
nor UO_819 (O_819,N_9975,N_9993);
or UO_820 (O_820,N_9993,N_9920);
or UO_821 (O_821,N_9908,N_9970);
and UO_822 (O_822,N_9952,N_9917);
or UO_823 (O_823,N_9980,N_9949);
and UO_824 (O_824,N_9930,N_9954);
or UO_825 (O_825,N_9933,N_9928);
nand UO_826 (O_826,N_9972,N_9949);
or UO_827 (O_827,N_9980,N_9972);
nand UO_828 (O_828,N_9963,N_9942);
xor UO_829 (O_829,N_9902,N_9925);
or UO_830 (O_830,N_9927,N_9993);
nor UO_831 (O_831,N_9923,N_9908);
nor UO_832 (O_832,N_9977,N_9940);
nor UO_833 (O_833,N_9971,N_9949);
and UO_834 (O_834,N_9916,N_9955);
nor UO_835 (O_835,N_9911,N_9998);
xnor UO_836 (O_836,N_9964,N_9915);
or UO_837 (O_837,N_9965,N_9921);
or UO_838 (O_838,N_9935,N_9950);
and UO_839 (O_839,N_9995,N_9967);
or UO_840 (O_840,N_9948,N_9913);
nor UO_841 (O_841,N_9910,N_9936);
xor UO_842 (O_842,N_9966,N_9949);
and UO_843 (O_843,N_9974,N_9980);
or UO_844 (O_844,N_9923,N_9952);
xor UO_845 (O_845,N_9924,N_9945);
or UO_846 (O_846,N_9966,N_9908);
or UO_847 (O_847,N_9975,N_9939);
xnor UO_848 (O_848,N_9929,N_9901);
nand UO_849 (O_849,N_9921,N_9997);
xor UO_850 (O_850,N_9903,N_9902);
nand UO_851 (O_851,N_9987,N_9946);
nor UO_852 (O_852,N_9994,N_9963);
or UO_853 (O_853,N_9958,N_9941);
and UO_854 (O_854,N_9967,N_9951);
or UO_855 (O_855,N_9963,N_9932);
nand UO_856 (O_856,N_9965,N_9951);
nand UO_857 (O_857,N_9992,N_9949);
and UO_858 (O_858,N_9918,N_9927);
nand UO_859 (O_859,N_9980,N_9995);
nor UO_860 (O_860,N_9943,N_9911);
xnor UO_861 (O_861,N_9978,N_9939);
and UO_862 (O_862,N_9966,N_9960);
xnor UO_863 (O_863,N_9921,N_9984);
xor UO_864 (O_864,N_9986,N_9956);
and UO_865 (O_865,N_9945,N_9987);
or UO_866 (O_866,N_9901,N_9942);
and UO_867 (O_867,N_9970,N_9907);
xor UO_868 (O_868,N_9948,N_9939);
or UO_869 (O_869,N_9991,N_9969);
nor UO_870 (O_870,N_9944,N_9947);
xor UO_871 (O_871,N_9992,N_9947);
xnor UO_872 (O_872,N_9967,N_9965);
or UO_873 (O_873,N_9956,N_9940);
and UO_874 (O_874,N_9961,N_9957);
nand UO_875 (O_875,N_9915,N_9994);
nor UO_876 (O_876,N_9958,N_9902);
xnor UO_877 (O_877,N_9923,N_9940);
or UO_878 (O_878,N_9929,N_9927);
and UO_879 (O_879,N_9968,N_9957);
xor UO_880 (O_880,N_9912,N_9981);
xor UO_881 (O_881,N_9981,N_9904);
and UO_882 (O_882,N_9945,N_9922);
nor UO_883 (O_883,N_9953,N_9959);
nand UO_884 (O_884,N_9995,N_9997);
and UO_885 (O_885,N_9902,N_9951);
nor UO_886 (O_886,N_9930,N_9936);
nor UO_887 (O_887,N_9979,N_9921);
xor UO_888 (O_888,N_9918,N_9953);
nor UO_889 (O_889,N_9982,N_9992);
xnor UO_890 (O_890,N_9955,N_9949);
xor UO_891 (O_891,N_9913,N_9924);
or UO_892 (O_892,N_9961,N_9918);
nor UO_893 (O_893,N_9947,N_9900);
xnor UO_894 (O_894,N_9918,N_9942);
nand UO_895 (O_895,N_9994,N_9954);
xnor UO_896 (O_896,N_9969,N_9931);
and UO_897 (O_897,N_9900,N_9939);
nand UO_898 (O_898,N_9903,N_9966);
nand UO_899 (O_899,N_9925,N_9934);
and UO_900 (O_900,N_9963,N_9957);
nand UO_901 (O_901,N_9975,N_9914);
or UO_902 (O_902,N_9966,N_9992);
or UO_903 (O_903,N_9932,N_9919);
or UO_904 (O_904,N_9965,N_9927);
and UO_905 (O_905,N_9993,N_9988);
nand UO_906 (O_906,N_9998,N_9989);
or UO_907 (O_907,N_9980,N_9955);
and UO_908 (O_908,N_9976,N_9923);
and UO_909 (O_909,N_9954,N_9939);
nor UO_910 (O_910,N_9949,N_9996);
xor UO_911 (O_911,N_9990,N_9976);
xnor UO_912 (O_912,N_9998,N_9902);
and UO_913 (O_913,N_9969,N_9988);
or UO_914 (O_914,N_9905,N_9982);
and UO_915 (O_915,N_9923,N_9949);
or UO_916 (O_916,N_9947,N_9983);
xnor UO_917 (O_917,N_9994,N_9945);
nand UO_918 (O_918,N_9996,N_9906);
nor UO_919 (O_919,N_9960,N_9925);
and UO_920 (O_920,N_9933,N_9949);
xor UO_921 (O_921,N_9978,N_9984);
and UO_922 (O_922,N_9913,N_9958);
nor UO_923 (O_923,N_9931,N_9947);
or UO_924 (O_924,N_9930,N_9953);
nor UO_925 (O_925,N_9991,N_9944);
nand UO_926 (O_926,N_9940,N_9952);
or UO_927 (O_927,N_9966,N_9970);
nor UO_928 (O_928,N_9930,N_9933);
xnor UO_929 (O_929,N_9939,N_9974);
nand UO_930 (O_930,N_9916,N_9905);
nand UO_931 (O_931,N_9914,N_9981);
and UO_932 (O_932,N_9950,N_9923);
nor UO_933 (O_933,N_9924,N_9988);
or UO_934 (O_934,N_9984,N_9917);
or UO_935 (O_935,N_9948,N_9927);
xnor UO_936 (O_936,N_9990,N_9928);
and UO_937 (O_937,N_9952,N_9928);
nand UO_938 (O_938,N_9948,N_9995);
or UO_939 (O_939,N_9995,N_9903);
nand UO_940 (O_940,N_9907,N_9950);
and UO_941 (O_941,N_9978,N_9950);
xor UO_942 (O_942,N_9951,N_9961);
or UO_943 (O_943,N_9944,N_9918);
nor UO_944 (O_944,N_9942,N_9956);
and UO_945 (O_945,N_9918,N_9972);
nor UO_946 (O_946,N_9960,N_9996);
xnor UO_947 (O_947,N_9907,N_9948);
and UO_948 (O_948,N_9999,N_9911);
or UO_949 (O_949,N_9912,N_9925);
xor UO_950 (O_950,N_9942,N_9979);
nand UO_951 (O_951,N_9998,N_9933);
xor UO_952 (O_952,N_9984,N_9961);
xnor UO_953 (O_953,N_9994,N_9935);
nor UO_954 (O_954,N_9959,N_9909);
and UO_955 (O_955,N_9944,N_9969);
nor UO_956 (O_956,N_9932,N_9968);
or UO_957 (O_957,N_9918,N_9920);
xnor UO_958 (O_958,N_9912,N_9938);
nor UO_959 (O_959,N_9982,N_9939);
xnor UO_960 (O_960,N_9926,N_9918);
or UO_961 (O_961,N_9922,N_9974);
nor UO_962 (O_962,N_9918,N_9992);
and UO_963 (O_963,N_9912,N_9910);
nor UO_964 (O_964,N_9987,N_9959);
and UO_965 (O_965,N_9993,N_9924);
nand UO_966 (O_966,N_9919,N_9917);
or UO_967 (O_967,N_9902,N_9961);
and UO_968 (O_968,N_9965,N_9938);
nor UO_969 (O_969,N_9918,N_9982);
nand UO_970 (O_970,N_9977,N_9902);
nor UO_971 (O_971,N_9905,N_9996);
nand UO_972 (O_972,N_9920,N_9960);
nor UO_973 (O_973,N_9965,N_9958);
nor UO_974 (O_974,N_9963,N_9913);
and UO_975 (O_975,N_9928,N_9975);
nand UO_976 (O_976,N_9966,N_9950);
xnor UO_977 (O_977,N_9920,N_9933);
and UO_978 (O_978,N_9994,N_9946);
or UO_979 (O_979,N_9933,N_9972);
or UO_980 (O_980,N_9987,N_9963);
nand UO_981 (O_981,N_9964,N_9987);
xor UO_982 (O_982,N_9963,N_9908);
xor UO_983 (O_983,N_9911,N_9940);
nor UO_984 (O_984,N_9922,N_9930);
nand UO_985 (O_985,N_9968,N_9959);
nand UO_986 (O_986,N_9953,N_9951);
nor UO_987 (O_987,N_9965,N_9910);
nor UO_988 (O_988,N_9967,N_9924);
xor UO_989 (O_989,N_9975,N_9947);
xnor UO_990 (O_990,N_9968,N_9946);
and UO_991 (O_991,N_9951,N_9987);
and UO_992 (O_992,N_9913,N_9992);
or UO_993 (O_993,N_9997,N_9984);
or UO_994 (O_994,N_9956,N_9932);
or UO_995 (O_995,N_9971,N_9962);
nor UO_996 (O_996,N_9912,N_9907);
xnor UO_997 (O_997,N_9910,N_9980);
and UO_998 (O_998,N_9991,N_9961);
nor UO_999 (O_999,N_9951,N_9940);
nor UO_1000 (O_1000,N_9923,N_9927);
or UO_1001 (O_1001,N_9911,N_9931);
nor UO_1002 (O_1002,N_9981,N_9946);
xnor UO_1003 (O_1003,N_9995,N_9961);
nand UO_1004 (O_1004,N_9919,N_9922);
and UO_1005 (O_1005,N_9936,N_9953);
nor UO_1006 (O_1006,N_9957,N_9991);
and UO_1007 (O_1007,N_9939,N_9940);
xnor UO_1008 (O_1008,N_9980,N_9951);
xor UO_1009 (O_1009,N_9932,N_9921);
nand UO_1010 (O_1010,N_9935,N_9962);
nand UO_1011 (O_1011,N_9996,N_9913);
and UO_1012 (O_1012,N_9910,N_9949);
xor UO_1013 (O_1013,N_9994,N_9974);
nor UO_1014 (O_1014,N_9925,N_9935);
nor UO_1015 (O_1015,N_9944,N_9907);
and UO_1016 (O_1016,N_9954,N_9927);
and UO_1017 (O_1017,N_9922,N_9905);
nor UO_1018 (O_1018,N_9962,N_9988);
nand UO_1019 (O_1019,N_9991,N_9918);
nand UO_1020 (O_1020,N_9965,N_9975);
and UO_1021 (O_1021,N_9946,N_9945);
nor UO_1022 (O_1022,N_9998,N_9958);
nand UO_1023 (O_1023,N_9963,N_9901);
nand UO_1024 (O_1024,N_9937,N_9999);
nand UO_1025 (O_1025,N_9991,N_9974);
xor UO_1026 (O_1026,N_9961,N_9921);
or UO_1027 (O_1027,N_9950,N_9940);
xnor UO_1028 (O_1028,N_9984,N_9910);
and UO_1029 (O_1029,N_9976,N_9963);
and UO_1030 (O_1030,N_9912,N_9963);
nor UO_1031 (O_1031,N_9946,N_9927);
or UO_1032 (O_1032,N_9950,N_9953);
nand UO_1033 (O_1033,N_9954,N_9922);
or UO_1034 (O_1034,N_9908,N_9901);
and UO_1035 (O_1035,N_9977,N_9913);
xnor UO_1036 (O_1036,N_9902,N_9920);
or UO_1037 (O_1037,N_9988,N_9961);
xnor UO_1038 (O_1038,N_9972,N_9902);
nor UO_1039 (O_1039,N_9921,N_9911);
or UO_1040 (O_1040,N_9950,N_9934);
and UO_1041 (O_1041,N_9993,N_9957);
nor UO_1042 (O_1042,N_9962,N_9957);
nor UO_1043 (O_1043,N_9949,N_9945);
nand UO_1044 (O_1044,N_9929,N_9935);
or UO_1045 (O_1045,N_9911,N_9934);
xnor UO_1046 (O_1046,N_9911,N_9995);
and UO_1047 (O_1047,N_9967,N_9940);
nor UO_1048 (O_1048,N_9944,N_9925);
or UO_1049 (O_1049,N_9956,N_9913);
or UO_1050 (O_1050,N_9940,N_9942);
or UO_1051 (O_1051,N_9973,N_9920);
and UO_1052 (O_1052,N_9917,N_9993);
and UO_1053 (O_1053,N_9968,N_9909);
or UO_1054 (O_1054,N_9956,N_9959);
and UO_1055 (O_1055,N_9989,N_9976);
and UO_1056 (O_1056,N_9994,N_9959);
or UO_1057 (O_1057,N_9933,N_9950);
nand UO_1058 (O_1058,N_9912,N_9983);
nor UO_1059 (O_1059,N_9990,N_9979);
or UO_1060 (O_1060,N_9960,N_9940);
nand UO_1061 (O_1061,N_9925,N_9914);
and UO_1062 (O_1062,N_9931,N_9973);
nand UO_1063 (O_1063,N_9904,N_9985);
nor UO_1064 (O_1064,N_9908,N_9974);
nor UO_1065 (O_1065,N_9986,N_9911);
xnor UO_1066 (O_1066,N_9985,N_9910);
nor UO_1067 (O_1067,N_9959,N_9935);
nand UO_1068 (O_1068,N_9933,N_9959);
nor UO_1069 (O_1069,N_9967,N_9907);
or UO_1070 (O_1070,N_9902,N_9966);
and UO_1071 (O_1071,N_9914,N_9911);
or UO_1072 (O_1072,N_9925,N_9928);
or UO_1073 (O_1073,N_9990,N_9964);
or UO_1074 (O_1074,N_9923,N_9947);
nor UO_1075 (O_1075,N_9982,N_9980);
or UO_1076 (O_1076,N_9981,N_9902);
nor UO_1077 (O_1077,N_9955,N_9992);
and UO_1078 (O_1078,N_9944,N_9909);
and UO_1079 (O_1079,N_9925,N_9999);
xor UO_1080 (O_1080,N_9906,N_9992);
nor UO_1081 (O_1081,N_9945,N_9912);
and UO_1082 (O_1082,N_9989,N_9903);
xnor UO_1083 (O_1083,N_9944,N_9932);
and UO_1084 (O_1084,N_9959,N_9913);
or UO_1085 (O_1085,N_9931,N_9979);
or UO_1086 (O_1086,N_9975,N_9941);
or UO_1087 (O_1087,N_9934,N_9988);
and UO_1088 (O_1088,N_9917,N_9941);
nor UO_1089 (O_1089,N_9958,N_9996);
and UO_1090 (O_1090,N_9987,N_9968);
nand UO_1091 (O_1091,N_9992,N_9927);
nor UO_1092 (O_1092,N_9999,N_9943);
or UO_1093 (O_1093,N_9943,N_9990);
nor UO_1094 (O_1094,N_9980,N_9993);
or UO_1095 (O_1095,N_9917,N_9907);
or UO_1096 (O_1096,N_9970,N_9926);
and UO_1097 (O_1097,N_9999,N_9984);
or UO_1098 (O_1098,N_9923,N_9996);
nand UO_1099 (O_1099,N_9965,N_9980);
or UO_1100 (O_1100,N_9919,N_9992);
or UO_1101 (O_1101,N_9989,N_9980);
nor UO_1102 (O_1102,N_9904,N_9900);
xnor UO_1103 (O_1103,N_9924,N_9927);
or UO_1104 (O_1104,N_9987,N_9924);
nand UO_1105 (O_1105,N_9959,N_9993);
or UO_1106 (O_1106,N_9998,N_9912);
and UO_1107 (O_1107,N_9985,N_9999);
nor UO_1108 (O_1108,N_9965,N_9950);
xor UO_1109 (O_1109,N_9900,N_9913);
nor UO_1110 (O_1110,N_9954,N_9929);
nor UO_1111 (O_1111,N_9945,N_9906);
xor UO_1112 (O_1112,N_9958,N_9921);
nor UO_1113 (O_1113,N_9919,N_9989);
or UO_1114 (O_1114,N_9995,N_9968);
and UO_1115 (O_1115,N_9904,N_9946);
xor UO_1116 (O_1116,N_9901,N_9965);
or UO_1117 (O_1117,N_9990,N_9972);
nor UO_1118 (O_1118,N_9901,N_9961);
or UO_1119 (O_1119,N_9920,N_9917);
and UO_1120 (O_1120,N_9993,N_9928);
nor UO_1121 (O_1121,N_9927,N_9938);
or UO_1122 (O_1122,N_9952,N_9903);
nand UO_1123 (O_1123,N_9948,N_9973);
or UO_1124 (O_1124,N_9929,N_9960);
or UO_1125 (O_1125,N_9957,N_9931);
nand UO_1126 (O_1126,N_9906,N_9977);
nor UO_1127 (O_1127,N_9946,N_9914);
nor UO_1128 (O_1128,N_9951,N_9976);
xnor UO_1129 (O_1129,N_9936,N_9914);
or UO_1130 (O_1130,N_9973,N_9916);
nand UO_1131 (O_1131,N_9985,N_9916);
xor UO_1132 (O_1132,N_9923,N_9912);
or UO_1133 (O_1133,N_9933,N_9965);
xor UO_1134 (O_1134,N_9998,N_9932);
and UO_1135 (O_1135,N_9912,N_9952);
or UO_1136 (O_1136,N_9911,N_9973);
nor UO_1137 (O_1137,N_9907,N_9910);
and UO_1138 (O_1138,N_9906,N_9973);
nor UO_1139 (O_1139,N_9970,N_9939);
or UO_1140 (O_1140,N_9982,N_9956);
and UO_1141 (O_1141,N_9972,N_9953);
or UO_1142 (O_1142,N_9970,N_9931);
xor UO_1143 (O_1143,N_9941,N_9966);
nand UO_1144 (O_1144,N_9987,N_9930);
nand UO_1145 (O_1145,N_9925,N_9983);
nand UO_1146 (O_1146,N_9998,N_9993);
nand UO_1147 (O_1147,N_9995,N_9917);
nand UO_1148 (O_1148,N_9914,N_9915);
xor UO_1149 (O_1149,N_9987,N_9984);
and UO_1150 (O_1150,N_9922,N_9983);
xnor UO_1151 (O_1151,N_9932,N_9914);
and UO_1152 (O_1152,N_9934,N_9917);
xor UO_1153 (O_1153,N_9996,N_9942);
or UO_1154 (O_1154,N_9925,N_9945);
nor UO_1155 (O_1155,N_9966,N_9958);
and UO_1156 (O_1156,N_9926,N_9934);
and UO_1157 (O_1157,N_9905,N_9941);
xor UO_1158 (O_1158,N_9968,N_9926);
xor UO_1159 (O_1159,N_9900,N_9965);
or UO_1160 (O_1160,N_9970,N_9928);
nor UO_1161 (O_1161,N_9930,N_9974);
xor UO_1162 (O_1162,N_9926,N_9938);
and UO_1163 (O_1163,N_9995,N_9900);
nor UO_1164 (O_1164,N_9955,N_9939);
and UO_1165 (O_1165,N_9928,N_9940);
or UO_1166 (O_1166,N_9975,N_9917);
or UO_1167 (O_1167,N_9909,N_9936);
xnor UO_1168 (O_1168,N_9922,N_9901);
and UO_1169 (O_1169,N_9959,N_9995);
nor UO_1170 (O_1170,N_9919,N_9900);
nand UO_1171 (O_1171,N_9963,N_9941);
nor UO_1172 (O_1172,N_9968,N_9901);
and UO_1173 (O_1173,N_9950,N_9993);
and UO_1174 (O_1174,N_9939,N_9992);
or UO_1175 (O_1175,N_9949,N_9973);
nor UO_1176 (O_1176,N_9959,N_9954);
and UO_1177 (O_1177,N_9912,N_9959);
xnor UO_1178 (O_1178,N_9936,N_9928);
xnor UO_1179 (O_1179,N_9976,N_9983);
nand UO_1180 (O_1180,N_9962,N_9951);
nor UO_1181 (O_1181,N_9950,N_9971);
nor UO_1182 (O_1182,N_9980,N_9957);
nand UO_1183 (O_1183,N_9997,N_9922);
nand UO_1184 (O_1184,N_9913,N_9982);
or UO_1185 (O_1185,N_9997,N_9926);
nor UO_1186 (O_1186,N_9906,N_9962);
nand UO_1187 (O_1187,N_9923,N_9942);
nand UO_1188 (O_1188,N_9958,N_9976);
nand UO_1189 (O_1189,N_9970,N_9929);
or UO_1190 (O_1190,N_9987,N_9989);
and UO_1191 (O_1191,N_9993,N_9969);
xor UO_1192 (O_1192,N_9991,N_9942);
and UO_1193 (O_1193,N_9995,N_9933);
nor UO_1194 (O_1194,N_9940,N_9965);
or UO_1195 (O_1195,N_9947,N_9915);
or UO_1196 (O_1196,N_9931,N_9942);
or UO_1197 (O_1197,N_9995,N_9994);
or UO_1198 (O_1198,N_9989,N_9999);
or UO_1199 (O_1199,N_9935,N_9926);
nand UO_1200 (O_1200,N_9976,N_9970);
and UO_1201 (O_1201,N_9962,N_9953);
xor UO_1202 (O_1202,N_9933,N_9954);
or UO_1203 (O_1203,N_9919,N_9942);
or UO_1204 (O_1204,N_9923,N_9984);
and UO_1205 (O_1205,N_9914,N_9921);
nor UO_1206 (O_1206,N_9987,N_9990);
or UO_1207 (O_1207,N_9973,N_9961);
nor UO_1208 (O_1208,N_9937,N_9915);
and UO_1209 (O_1209,N_9965,N_9997);
and UO_1210 (O_1210,N_9901,N_9913);
or UO_1211 (O_1211,N_9909,N_9939);
nand UO_1212 (O_1212,N_9975,N_9994);
and UO_1213 (O_1213,N_9928,N_9995);
or UO_1214 (O_1214,N_9917,N_9939);
nand UO_1215 (O_1215,N_9974,N_9957);
nor UO_1216 (O_1216,N_9938,N_9966);
or UO_1217 (O_1217,N_9925,N_9919);
and UO_1218 (O_1218,N_9918,N_9994);
nor UO_1219 (O_1219,N_9928,N_9923);
or UO_1220 (O_1220,N_9936,N_9960);
or UO_1221 (O_1221,N_9933,N_9943);
nand UO_1222 (O_1222,N_9952,N_9936);
xnor UO_1223 (O_1223,N_9996,N_9962);
and UO_1224 (O_1224,N_9977,N_9970);
or UO_1225 (O_1225,N_9906,N_9990);
and UO_1226 (O_1226,N_9947,N_9982);
xnor UO_1227 (O_1227,N_9964,N_9938);
and UO_1228 (O_1228,N_9955,N_9923);
nand UO_1229 (O_1229,N_9994,N_9924);
nor UO_1230 (O_1230,N_9998,N_9939);
and UO_1231 (O_1231,N_9966,N_9936);
and UO_1232 (O_1232,N_9903,N_9990);
nand UO_1233 (O_1233,N_9950,N_9989);
and UO_1234 (O_1234,N_9926,N_9915);
and UO_1235 (O_1235,N_9959,N_9934);
nor UO_1236 (O_1236,N_9912,N_9965);
nand UO_1237 (O_1237,N_9974,N_9909);
nand UO_1238 (O_1238,N_9900,N_9938);
nand UO_1239 (O_1239,N_9930,N_9952);
and UO_1240 (O_1240,N_9922,N_9917);
nand UO_1241 (O_1241,N_9972,N_9919);
xnor UO_1242 (O_1242,N_9929,N_9907);
nor UO_1243 (O_1243,N_9969,N_9929);
nand UO_1244 (O_1244,N_9915,N_9974);
nor UO_1245 (O_1245,N_9998,N_9920);
nor UO_1246 (O_1246,N_9923,N_9978);
or UO_1247 (O_1247,N_9950,N_9903);
xnor UO_1248 (O_1248,N_9981,N_9944);
and UO_1249 (O_1249,N_9909,N_9943);
or UO_1250 (O_1250,N_9969,N_9924);
or UO_1251 (O_1251,N_9980,N_9904);
nor UO_1252 (O_1252,N_9922,N_9946);
or UO_1253 (O_1253,N_9984,N_9957);
or UO_1254 (O_1254,N_9965,N_9962);
or UO_1255 (O_1255,N_9975,N_9976);
nor UO_1256 (O_1256,N_9985,N_9973);
or UO_1257 (O_1257,N_9929,N_9905);
and UO_1258 (O_1258,N_9946,N_9923);
and UO_1259 (O_1259,N_9988,N_9900);
nor UO_1260 (O_1260,N_9955,N_9910);
or UO_1261 (O_1261,N_9909,N_9986);
and UO_1262 (O_1262,N_9907,N_9930);
nand UO_1263 (O_1263,N_9989,N_9935);
nor UO_1264 (O_1264,N_9991,N_9946);
and UO_1265 (O_1265,N_9988,N_9928);
nor UO_1266 (O_1266,N_9943,N_9949);
or UO_1267 (O_1267,N_9947,N_9968);
or UO_1268 (O_1268,N_9979,N_9951);
xor UO_1269 (O_1269,N_9931,N_9919);
nand UO_1270 (O_1270,N_9959,N_9996);
xnor UO_1271 (O_1271,N_9954,N_9909);
nand UO_1272 (O_1272,N_9941,N_9981);
nor UO_1273 (O_1273,N_9915,N_9954);
nor UO_1274 (O_1274,N_9991,N_9978);
xnor UO_1275 (O_1275,N_9996,N_9940);
nand UO_1276 (O_1276,N_9926,N_9976);
nand UO_1277 (O_1277,N_9910,N_9979);
and UO_1278 (O_1278,N_9974,N_9997);
and UO_1279 (O_1279,N_9990,N_9907);
or UO_1280 (O_1280,N_9933,N_9970);
and UO_1281 (O_1281,N_9964,N_9996);
or UO_1282 (O_1282,N_9909,N_9932);
xor UO_1283 (O_1283,N_9921,N_9967);
and UO_1284 (O_1284,N_9955,N_9997);
nor UO_1285 (O_1285,N_9906,N_9946);
or UO_1286 (O_1286,N_9947,N_9988);
or UO_1287 (O_1287,N_9935,N_9903);
nand UO_1288 (O_1288,N_9928,N_9964);
xor UO_1289 (O_1289,N_9959,N_9960);
nor UO_1290 (O_1290,N_9929,N_9987);
nor UO_1291 (O_1291,N_9972,N_9910);
or UO_1292 (O_1292,N_9952,N_9949);
or UO_1293 (O_1293,N_9969,N_9925);
xor UO_1294 (O_1294,N_9992,N_9934);
nand UO_1295 (O_1295,N_9904,N_9901);
nor UO_1296 (O_1296,N_9983,N_9982);
and UO_1297 (O_1297,N_9916,N_9999);
or UO_1298 (O_1298,N_9935,N_9980);
nor UO_1299 (O_1299,N_9920,N_9927);
nor UO_1300 (O_1300,N_9983,N_9939);
and UO_1301 (O_1301,N_9983,N_9909);
nor UO_1302 (O_1302,N_9974,N_9986);
nand UO_1303 (O_1303,N_9947,N_9973);
or UO_1304 (O_1304,N_9975,N_9944);
or UO_1305 (O_1305,N_9985,N_9947);
nor UO_1306 (O_1306,N_9913,N_9972);
and UO_1307 (O_1307,N_9981,N_9953);
xnor UO_1308 (O_1308,N_9930,N_9940);
nor UO_1309 (O_1309,N_9957,N_9964);
nand UO_1310 (O_1310,N_9935,N_9998);
xnor UO_1311 (O_1311,N_9915,N_9971);
and UO_1312 (O_1312,N_9951,N_9939);
and UO_1313 (O_1313,N_9911,N_9981);
nand UO_1314 (O_1314,N_9957,N_9967);
or UO_1315 (O_1315,N_9968,N_9923);
and UO_1316 (O_1316,N_9997,N_9981);
nand UO_1317 (O_1317,N_9917,N_9931);
xnor UO_1318 (O_1318,N_9988,N_9951);
nand UO_1319 (O_1319,N_9931,N_9998);
nor UO_1320 (O_1320,N_9911,N_9968);
or UO_1321 (O_1321,N_9976,N_9988);
nor UO_1322 (O_1322,N_9997,N_9911);
or UO_1323 (O_1323,N_9980,N_9940);
and UO_1324 (O_1324,N_9938,N_9937);
nor UO_1325 (O_1325,N_9971,N_9925);
or UO_1326 (O_1326,N_9987,N_9923);
nand UO_1327 (O_1327,N_9967,N_9916);
or UO_1328 (O_1328,N_9938,N_9978);
xnor UO_1329 (O_1329,N_9959,N_9971);
or UO_1330 (O_1330,N_9911,N_9984);
or UO_1331 (O_1331,N_9927,N_9963);
xnor UO_1332 (O_1332,N_9948,N_9934);
xnor UO_1333 (O_1333,N_9977,N_9941);
or UO_1334 (O_1334,N_9942,N_9907);
and UO_1335 (O_1335,N_9987,N_9950);
or UO_1336 (O_1336,N_9941,N_9923);
and UO_1337 (O_1337,N_9950,N_9997);
nand UO_1338 (O_1338,N_9959,N_9955);
or UO_1339 (O_1339,N_9920,N_9947);
xor UO_1340 (O_1340,N_9914,N_9974);
nand UO_1341 (O_1341,N_9937,N_9911);
or UO_1342 (O_1342,N_9909,N_9937);
and UO_1343 (O_1343,N_9923,N_9975);
xor UO_1344 (O_1344,N_9969,N_9940);
nor UO_1345 (O_1345,N_9994,N_9926);
nor UO_1346 (O_1346,N_9966,N_9923);
nand UO_1347 (O_1347,N_9925,N_9980);
and UO_1348 (O_1348,N_9987,N_9916);
nor UO_1349 (O_1349,N_9989,N_9923);
and UO_1350 (O_1350,N_9964,N_9958);
nor UO_1351 (O_1351,N_9996,N_9993);
xor UO_1352 (O_1352,N_9959,N_9972);
nand UO_1353 (O_1353,N_9905,N_9987);
xnor UO_1354 (O_1354,N_9919,N_9968);
nand UO_1355 (O_1355,N_9983,N_9966);
xor UO_1356 (O_1356,N_9917,N_9936);
and UO_1357 (O_1357,N_9999,N_9907);
or UO_1358 (O_1358,N_9981,N_9940);
xnor UO_1359 (O_1359,N_9980,N_9900);
nor UO_1360 (O_1360,N_9928,N_9960);
or UO_1361 (O_1361,N_9962,N_9946);
and UO_1362 (O_1362,N_9969,N_9985);
nand UO_1363 (O_1363,N_9995,N_9952);
nor UO_1364 (O_1364,N_9910,N_9937);
nand UO_1365 (O_1365,N_9924,N_9919);
and UO_1366 (O_1366,N_9950,N_9949);
nor UO_1367 (O_1367,N_9916,N_9907);
xor UO_1368 (O_1368,N_9940,N_9943);
or UO_1369 (O_1369,N_9995,N_9984);
and UO_1370 (O_1370,N_9953,N_9925);
nand UO_1371 (O_1371,N_9960,N_9912);
nand UO_1372 (O_1372,N_9920,N_9986);
and UO_1373 (O_1373,N_9987,N_9903);
nor UO_1374 (O_1374,N_9937,N_9946);
or UO_1375 (O_1375,N_9966,N_9953);
or UO_1376 (O_1376,N_9972,N_9958);
nand UO_1377 (O_1377,N_9926,N_9912);
xor UO_1378 (O_1378,N_9955,N_9903);
and UO_1379 (O_1379,N_9921,N_9917);
nand UO_1380 (O_1380,N_9975,N_9932);
nor UO_1381 (O_1381,N_9975,N_9997);
nor UO_1382 (O_1382,N_9951,N_9983);
and UO_1383 (O_1383,N_9964,N_9986);
xnor UO_1384 (O_1384,N_9961,N_9990);
nor UO_1385 (O_1385,N_9901,N_9946);
nand UO_1386 (O_1386,N_9915,N_9908);
or UO_1387 (O_1387,N_9919,N_9954);
xnor UO_1388 (O_1388,N_9962,N_9908);
nand UO_1389 (O_1389,N_9900,N_9921);
nor UO_1390 (O_1390,N_9958,N_9979);
xnor UO_1391 (O_1391,N_9973,N_9957);
xnor UO_1392 (O_1392,N_9930,N_9925);
and UO_1393 (O_1393,N_9922,N_9934);
and UO_1394 (O_1394,N_9927,N_9910);
or UO_1395 (O_1395,N_9960,N_9992);
xor UO_1396 (O_1396,N_9940,N_9992);
nor UO_1397 (O_1397,N_9938,N_9920);
nand UO_1398 (O_1398,N_9909,N_9949);
nand UO_1399 (O_1399,N_9954,N_9996);
xnor UO_1400 (O_1400,N_9977,N_9972);
or UO_1401 (O_1401,N_9982,N_9959);
nor UO_1402 (O_1402,N_9963,N_9965);
nor UO_1403 (O_1403,N_9923,N_9965);
nor UO_1404 (O_1404,N_9944,N_9967);
nor UO_1405 (O_1405,N_9937,N_9954);
nor UO_1406 (O_1406,N_9934,N_9923);
and UO_1407 (O_1407,N_9976,N_9938);
nor UO_1408 (O_1408,N_9983,N_9913);
nor UO_1409 (O_1409,N_9980,N_9942);
and UO_1410 (O_1410,N_9998,N_9949);
nand UO_1411 (O_1411,N_9916,N_9923);
and UO_1412 (O_1412,N_9917,N_9963);
and UO_1413 (O_1413,N_9908,N_9954);
or UO_1414 (O_1414,N_9946,N_9974);
and UO_1415 (O_1415,N_9910,N_9930);
or UO_1416 (O_1416,N_9996,N_9997);
or UO_1417 (O_1417,N_9948,N_9990);
xor UO_1418 (O_1418,N_9993,N_9912);
and UO_1419 (O_1419,N_9918,N_9949);
xnor UO_1420 (O_1420,N_9914,N_9922);
xnor UO_1421 (O_1421,N_9919,N_9913);
or UO_1422 (O_1422,N_9905,N_9979);
xor UO_1423 (O_1423,N_9912,N_9992);
or UO_1424 (O_1424,N_9958,N_9918);
xor UO_1425 (O_1425,N_9914,N_9998);
nor UO_1426 (O_1426,N_9929,N_9995);
xnor UO_1427 (O_1427,N_9931,N_9951);
nor UO_1428 (O_1428,N_9990,N_9908);
nand UO_1429 (O_1429,N_9936,N_9968);
nand UO_1430 (O_1430,N_9917,N_9945);
nor UO_1431 (O_1431,N_9919,N_9960);
xnor UO_1432 (O_1432,N_9919,N_9937);
and UO_1433 (O_1433,N_9936,N_9977);
and UO_1434 (O_1434,N_9908,N_9948);
nor UO_1435 (O_1435,N_9994,N_9957);
nor UO_1436 (O_1436,N_9985,N_9911);
xor UO_1437 (O_1437,N_9902,N_9901);
or UO_1438 (O_1438,N_9953,N_9923);
and UO_1439 (O_1439,N_9965,N_9973);
nor UO_1440 (O_1440,N_9982,N_9987);
xnor UO_1441 (O_1441,N_9935,N_9904);
nor UO_1442 (O_1442,N_9992,N_9980);
nand UO_1443 (O_1443,N_9990,N_9995);
xnor UO_1444 (O_1444,N_9999,N_9939);
nor UO_1445 (O_1445,N_9904,N_9905);
and UO_1446 (O_1446,N_9901,N_9940);
nand UO_1447 (O_1447,N_9914,N_9926);
nor UO_1448 (O_1448,N_9910,N_9906);
or UO_1449 (O_1449,N_9922,N_9920);
nor UO_1450 (O_1450,N_9911,N_9958);
or UO_1451 (O_1451,N_9982,N_9991);
nor UO_1452 (O_1452,N_9907,N_9904);
or UO_1453 (O_1453,N_9922,N_9927);
xnor UO_1454 (O_1454,N_9952,N_9920);
or UO_1455 (O_1455,N_9976,N_9962);
and UO_1456 (O_1456,N_9960,N_9901);
nand UO_1457 (O_1457,N_9958,N_9907);
and UO_1458 (O_1458,N_9967,N_9979);
and UO_1459 (O_1459,N_9925,N_9940);
and UO_1460 (O_1460,N_9967,N_9972);
nand UO_1461 (O_1461,N_9910,N_9914);
nor UO_1462 (O_1462,N_9949,N_9999);
nand UO_1463 (O_1463,N_9938,N_9981);
nand UO_1464 (O_1464,N_9962,N_9928);
and UO_1465 (O_1465,N_9910,N_9920);
nor UO_1466 (O_1466,N_9944,N_9970);
or UO_1467 (O_1467,N_9967,N_9968);
and UO_1468 (O_1468,N_9913,N_9945);
or UO_1469 (O_1469,N_9906,N_9928);
or UO_1470 (O_1470,N_9946,N_9940);
and UO_1471 (O_1471,N_9983,N_9980);
and UO_1472 (O_1472,N_9950,N_9921);
or UO_1473 (O_1473,N_9992,N_9928);
xnor UO_1474 (O_1474,N_9947,N_9984);
xor UO_1475 (O_1475,N_9938,N_9911);
nor UO_1476 (O_1476,N_9912,N_9936);
and UO_1477 (O_1477,N_9996,N_9977);
xor UO_1478 (O_1478,N_9904,N_9977);
or UO_1479 (O_1479,N_9957,N_9908);
xnor UO_1480 (O_1480,N_9941,N_9971);
and UO_1481 (O_1481,N_9906,N_9987);
and UO_1482 (O_1482,N_9905,N_9945);
nor UO_1483 (O_1483,N_9900,N_9928);
and UO_1484 (O_1484,N_9927,N_9937);
or UO_1485 (O_1485,N_9977,N_9932);
nand UO_1486 (O_1486,N_9970,N_9945);
nand UO_1487 (O_1487,N_9990,N_9963);
xor UO_1488 (O_1488,N_9937,N_9902);
or UO_1489 (O_1489,N_9917,N_9962);
or UO_1490 (O_1490,N_9924,N_9904);
and UO_1491 (O_1491,N_9972,N_9923);
and UO_1492 (O_1492,N_9925,N_9946);
and UO_1493 (O_1493,N_9935,N_9913);
xnor UO_1494 (O_1494,N_9985,N_9933);
nand UO_1495 (O_1495,N_9912,N_9943);
and UO_1496 (O_1496,N_9974,N_9943);
or UO_1497 (O_1497,N_9950,N_9925);
or UO_1498 (O_1498,N_9980,N_9911);
nand UO_1499 (O_1499,N_9901,N_9923);
endmodule