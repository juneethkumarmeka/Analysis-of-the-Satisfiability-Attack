module basic_500_3000_500_6_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_190,In_375);
nand U1 (N_1,In_297,In_196);
nand U2 (N_2,In_10,In_359);
xnor U3 (N_3,In_6,In_305);
or U4 (N_4,In_276,In_425);
nand U5 (N_5,In_420,In_2);
nor U6 (N_6,In_310,In_421);
nor U7 (N_7,In_149,In_368);
nand U8 (N_8,In_114,In_378);
nor U9 (N_9,In_266,In_488);
nor U10 (N_10,In_122,In_111);
and U11 (N_11,In_129,In_479);
or U12 (N_12,In_20,In_292);
nand U13 (N_13,In_239,In_75);
or U14 (N_14,In_456,In_74);
xor U15 (N_15,In_7,In_346);
or U16 (N_16,In_381,In_370);
and U17 (N_17,In_256,In_207);
or U18 (N_18,In_429,In_162);
or U19 (N_19,In_22,In_95);
and U20 (N_20,In_433,In_324);
nand U21 (N_21,In_315,In_244);
xor U22 (N_22,In_308,In_438);
nor U23 (N_23,In_358,In_430);
or U24 (N_24,In_351,In_423);
nor U25 (N_25,In_79,In_236);
and U26 (N_26,In_274,In_102);
nand U27 (N_27,In_462,In_180);
nor U28 (N_28,In_61,In_495);
nand U29 (N_29,In_167,In_32);
nand U30 (N_30,In_209,In_374);
xor U31 (N_31,In_412,In_316);
xnor U32 (N_32,In_178,In_352);
nand U33 (N_33,In_335,In_53);
and U34 (N_34,In_41,In_270);
or U35 (N_35,In_123,In_81);
and U36 (N_36,In_281,In_131);
nand U37 (N_37,In_338,In_451);
or U38 (N_38,In_249,In_257);
nand U39 (N_39,In_128,In_48);
or U40 (N_40,In_90,In_384);
nor U41 (N_41,In_379,In_110);
nor U42 (N_42,In_477,In_182);
and U43 (N_43,In_169,In_86);
xor U44 (N_44,In_271,In_23);
xnor U45 (N_45,In_461,In_464);
nor U46 (N_46,In_158,In_255);
xor U47 (N_47,In_107,In_192);
nor U48 (N_48,In_83,In_36);
nor U49 (N_49,In_466,In_9);
and U50 (N_50,In_126,In_240);
or U51 (N_51,In_414,In_141);
or U52 (N_52,In_91,In_206);
and U53 (N_53,In_64,In_350);
or U54 (N_54,In_71,In_406);
and U55 (N_55,In_150,In_94);
xor U56 (N_56,In_432,In_37);
nand U57 (N_57,In_313,In_428);
nand U58 (N_58,In_388,In_476);
nor U59 (N_59,In_460,In_13);
xnor U60 (N_60,In_69,In_265);
nor U61 (N_61,In_470,In_220);
nor U62 (N_62,In_417,In_398);
nand U63 (N_63,In_469,In_437);
or U64 (N_64,In_104,In_106);
and U65 (N_65,In_117,In_387);
nand U66 (N_66,In_263,In_161);
or U67 (N_67,In_260,In_302);
xor U68 (N_68,In_24,In_17);
nand U69 (N_69,In_134,In_364);
nand U70 (N_70,In_232,In_436);
xnor U71 (N_71,In_355,In_321);
or U72 (N_72,In_184,In_280);
xnor U73 (N_73,In_96,In_208);
or U74 (N_74,In_395,In_418);
or U75 (N_75,In_309,In_185);
xor U76 (N_76,In_253,In_314);
nor U77 (N_77,In_199,In_35);
xnor U78 (N_78,In_73,In_402);
nor U79 (N_79,In_77,In_229);
nand U80 (N_80,In_404,In_76);
xor U81 (N_81,In_39,In_454);
nor U82 (N_82,In_98,In_393);
and U83 (N_83,In_5,In_340);
and U84 (N_84,In_168,In_112);
and U85 (N_85,In_250,In_225);
or U86 (N_86,In_245,In_286);
xnor U87 (N_87,In_19,In_92);
and U88 (N_88,In_365,In_45);
and U89 (N_89,In_170,In_344);
xor U90 (N_90,In_109,In_85);
xnor U91 (N_91,In_130,In_363);
nand U92 (N_92,In_480,In_57);
xnor U93 (N_93,In_103,In_473);
nor U94 (N_94,In_67,In_441);
nor U95 (N_95,In_383,In_28);
nor U96 (N_96,In_258,In_427);
nor U97 (N_97,In_319,In_60);
and U98 (N_98,In_431,In_186);
and U99 (N_99,In_163,In_226);
and U100 (N_100,In_285,In_216);
nor U101 (N_101,In_219,In_367);
nor U102 (N_102,In_361,In_147);
and U103 (N_103,In_334,In_332);
xor U104 (N_104,In_237,In_457);
nor U105 (N_105,In_63,In_27);
nand U106 (N_106,In_300,In_459);
and U107 (N_107,In_52,In_50);
and U108 (N_108,In_354,In_419);
xnor U109 (N_109,In_204,In_333);
xnor U110 (N_110,In_18,In_157);
nand U111 (N_111,In_336,In_179);
xnor U112 (N_112,In_264,In_31);
nor U113 (N_113,In_408,In_312);
or U114 (N_114,In_44,In_291);
xor U115 (N_115,In_136,In_160);
nor U116 (N_116,In_55,In_467);
nand U117 (N_117,In_440,In_318);
nor U118 (N_118,In_254,In_413);
or U119 (N_119,In_0,In_499);
nand U120 (N_120,In_177,In_140);
nor U121 (N_121,In_210,In_108);
or U122 (N_122,In_485,In_194);
or U123 (N_123,In_261,In_371);
or U124 (N_124,In_386,In_174);
xor U125 (N_125,In_228,In_84);
nor U126 (N_126,In_450,In_498);
nand U127 (N_127,In_349,In_449);
and U128 (N_128,In_8,In_360);
nand U129 (N_129,In_215,In_127);
nor U130 (N_130,In_288,In_203);
nand U131 (N_131,In_175,In_353);
or U132 (N_132,In_320,In_49);
or U133 (N_133,In_357,In_12);
xor U134 (N_134,In_135,In_296);
and U135 (N_135,In_472,In_295);
nand U136 (N_136,In_325,In_101);
and U137 (N_137,In_471,In_483);
nor U138 (N_138,In_205,In_156);
nand U139 (N_139,In_15,In_234);
nor U140 (N_140,In_1,In_284);
nand U141 (N_141,In_176,In_330);
nor U142 (N_142,In_411,In_113);
or U143 (N_143,In_100,In_400);
nand U144 (N_144,In_191,In_410);
nor U145 (N_145,In_247,In_491);
nand U146 (N_146,In_202,In_443);
xor U147 (N_147,In_329,In_153);
xnor U148 (N_148,In_246,In_455);
nor U149 (N_149,In_405,In_391);
xnor U150 (N_150,In_293,In_372);
or U151 (N_151,In_14,In_54);
or U152 (N_152,In_231,In_154);
or U153 (N_153,In_120,In_42);
xnor U154 (N_154,In_166,In_307);
and U155 (N_155,In_3,In_382);
and U156 (N_156,In_34,In_87);
nor U157 (N_157,In_4,In_97);
or U158 (N_158,In_342,In_463);
or U159 (N_159,In_145,In_487);
xnor U160 (N_160,In_89,In_221);
and U161 (N_161,In_181,In_65);
nor U162 (N_162,In_416,In_287);
or U163 (N_163,In_279,In_58);
or U164 (N_164,In_377,In_21);
and U165 (N_165,In_392,In_442);
or U166 (N_166,In_366,In_139);
and U167 (N_167,In_424,In_277);
xnor U168 (N_168,In_327,In_435);
or U169 (N_169,In_146,In_230);
and U170 (N_170,In_290,In_482);
or U171 (N_171,In_214,In_278);
nand U172 (N_172,In_242,In_51);
or U173 (N_173,In_119,In_369);
or U174 (N_174,In_481,In_337);
or U175 (N_175,In_275,In_447);
xor U176 (N_176,In_345,In_243);
xor U177 (N_177,In_137,In_227);
nor U178 (N_178,In_489,In_118);
or U179 (N_179,In_494,In_397);
xnor U180 (N_180,In_43,In_198);
or U181 (N_181,In_62,In_282);
nor U182 (N_182,In_407,In_304);
and U183 (N_183,In_294,In_484);
xnor U184 (N_184,In_99,In_72);
or U185 (N_185,In_70,In_26);
or U186 (N_186,In_331,In_306);
or U187 (N_187,In_46,In_262);
xor U188 (N_188,In_415,In_496);
and U189 (N_189,In_200,In_389);
nor U190 (N_190,In_273,In_422);
xor U191 (N_191,In_434,In_268);
nor U192 (N_192,In_409,In_187);
and U193 (N_193,In_348,In_143);
and U194 (N_194,In_326,In_448);
xor U195 (N_195,In_188,In_401);
xor U196 (N_196,In_47,In_16);
or U197 (N_197,In_356,In_317);
xor U198 (N_198,In_486,In_144);
or U199 (N_199,In_197,In_248);
nand U200 (N_200,In_490,In_68);
nand U201 (N_201,In_465,In_165);
nand U202 (N_202,In_115,In_29);
xnor U203 (N_203,In_159,In_376);
or U204 (N_204,In_125,In_211);
nand U205 (N_205,In_155,In_458);
nor U206 (N_206,In_121,In_171);
nor U207 (N_207,In_218,In_173);
nor U208 (N_208,In_303,In_252);
nand U209 (N_209,In_347,In_475);
and U210 (N_210,In_56,In_238);
xor U211 (N_211,In_66,In_311);
xnor U212 (N_212,In_172,In_152);
and U213 (N_213,In_267,In_183);
nand U214 (N_214,In_133,In_224);
nor U215 (N_215,In_269,In_341);
or U216 (N_216,In_299,In_339);
nand U217 (N_217,In_439,In_343);
or U218 (N_218,In_493,In_11);
nand U219 (N_219,In_116,In_59);
and U220 (N_220,In_497,In_272);
nand U221 (N_221,In_373,In_138);
nand U222 (N_222,In_233,In_193);
and U223 (N_223,In_301,In_445);
xor U224 (N_224,In_88,In_124);
nand U225 (N_225,In_148,In_30);
or U226 (N_226,In_478,In_474);
and U227 (N_227,In_38,In_213);
nand U228 (N_228,In_394,In_328);
or U229 (N_229,In_468,In_399);
xnor U230 (N_230,In_385,In_452);
and U231 (N_231,In_80,In_362);
xor U232 (N_232,In_403,In_105);
and U233 (N_233,In_259,In_241);
xor U234 (N_234,In_323,In_298);
nand U235 (N_235,In_151,In_164);
nand U236 (N_236,In_289,In_78);
and U237 (N_237,In_251,In_25);
nand U238 (N_238,In_40,In_380);
or U239 (N_239,In_217,In_132);
nand U240 (N_240,In_235,In_33);
nor U241 (N_241,In_444,In_492);
nand U242 (N_242,In_142,In_390);
or U243 (N_243,In_93,In_322);
nand U244 (N_244,In_426,In_396);
xnor U245 (N_245,In_283,In_212);
nand U246 (N_246,In_82,In_222);
and U247 (N_247,In_195,In_453);
nand U248 (N_248,In_201,In_189);
xor U249 (N_249,In_446,In_223);
nor U250 (N_250,In_395,In_219);
nor U251 (N_251,In_218,In_125);
nor U252 (N_252,In_122,In_466);
xnor U253 (N_253,In_154,In_251);
nor U254 (N_254,In_300,In_479);
xor U255 (N_255,In_210,In_327);
nand U256 (N_256,In_287,In_20);
nor U257 (N_257,In_465,In_312);
nor U258 (N_258,In_75,In_223);
xor U259 (N_259,In_55,In_311);
nor U260 (N_260,In_352,In_165);
and U261 (N_261,In_145,In_277);
xnor U262 (N_262,In_111,In_269);
and U263 (N_263,In_159,In_499);
xnor U264 (N_264,In_317,In_72);
and U265 (N_265,In_205,In_418);
and U266 (N_266,In_491,In_19);
and U267 (N_267,In_49,In_236);
xor U268 (N_268,In_474,In_95);
nand U269 (N_269,In_47,In_258);
or U270 (N_270,In_215,In_74);
and U271 (N_271,In_316,In_45);
xnor U272 (N_272,In_375,In_425);
xnor U273 (N_273,In_216,In_278);
and U274 (N_274,In_250,In_453);
and U275 (N_275,In_356,In_235);
and U276 (N_276,In_138,In_437);
nor U277 (N_277,In_123,In_162);
nor U278 (N_278,In_340,In_144);
and U279 (N_279,In_471,In_319);
nor U280 (N_280,In_67,In_140);
nor U281 (N_281,In_443,In_136);
and U282 (N_282,In_94,In_319);
and U283 (N_283,In_71,In_460);
nor U284 (N_284,In_15,In_153);
and U285 (N_285,In_248,In_212);
nand U286 (N_286,In_279,In_79);
nand U287 (N_287,In_404,In_319);
and U288 (N_288,In_54,In_136);
or U289 (N_289,In_64,In_471);
or U290 (N_290,In_400,In_347);
or U291 (N_291,In_58,In_62);
nand U292 (N_292,In_373,In_123);
or U293 (N_293,In_210,In_476);
nor U294 (N_294,In_285,In_384);
nand U295 (N_295,In_11,In_204);
xnor U296 (N_296,In_494,In_283);
nand U297 (N_297,In_406,In_126);
nand U298 (N_298,In_395,In_96);
nand U299 (N_299,In_277,In_60);
xor U300 (N_300,In_410,In_90);
xor U301 (N_301,In_25,In_319);
and U302 (N_302,In_125,In_89);
or U303 (N_303,In_90,In_202);
or U304 (N_304,In_380,In_60);
and U305 (N_305,In_39,In_419);
nor U306 (N_306,In_346,In_118);
xor U307 (N_307,In_263,In_29);
xor U308 (N_308,In_299,In_443);
and U309 (N_309,In_378,In_487);
and U310 (N_310,In_205,In_340);
or U311 (N_311,In_148,In_315);
or U312 (N_312,In_236,In_344);
and U313 (N_313,In_140,In_464);
nor U314 (N_314,In_293,In_195);
nor U315 (N_315,In_206,In_420);
or U316 (N_316,In_364,In_315);
nand U317 (N_317,In_186,In_90);
and U318 (N_318,In_253,In_117);
xor U319 (N_319,In_90,In_244);
xor U320 (N_320,In_477,In_266);
xor U321 (N_321,In_468,In_116);
or U322 (N_322,In_437,In_209);
xor U323 (N_323,In_98,In_367);
xor U324 (N_324,In_57,In_55);
and U325 (N_325,In_296,In_273);
nor U326 (N_326,In_241,In_11);
nand U327 (N_327,In_106,In_499);
or U328 (N_328,In_21,In_160);
or U329 (N_329,In_482,In_130);
nor U330 (N_330,In_130,In_367);
and U331 (N_331,In_273,In_335);
nor U332 (N_332,In_441,In_281);
or U333 (N_333,In_472,In_201);
xnor U334 (N_334,In_386,In_467);
and U335 (N_335,In_37,In_155);
nand U336 (N_336,In_183,In_191);
and U337 (N_337,In_437,In_277);
nor U338 (N_338,In_212,In_347);
nor U339 (N_339,In_166,In_278);
xor U340 (N_340,In_208,In_284);
or U341 (N_341,In_367,In_247);
or U342 (N_342,In_318,In_290);
or U343 (N_343,In_266,In_379);
and U344 (N_344,In_182,In_163);
nand U345 (N_345,In_269,In_392);
or U346 (N_346,In_469,In_404);
or U347 (N_347,In_339,In_425);
xor U348 (N_348,In_419,In_308);
nand U349 (N_349,In_199,In_154);
or U350 (N_350,In_490,In_159);
nand U351 (N_351,In_326,In_471);
xor U352 (N_352,In_337,In_277);
or U353 (N_353,In_231,In_46);
and U354 (N_354,In_171,In_347);
nand U355 (N_355,In_63,In_47);
or U356 (N_356,In_128,In_84);
nand U357 (N_357,In_441,In_187);
and U358 (N_358,In_472,In_444);
or U359 (N_359,In_331,In_10);
and U360 (N_360,In_376,In_352);
xnor U361 (N_361,In_59,In_422);
and U362 (N_362,In_41,In_476);
nand U363 (N_363,In_427,In_142);
nor U364 (N_364,In_207,In_140);
xnor U365 (N_365,In_358,In_31);
or U366 (N_366,In_225,In_14);
or U367 (N_367,In_247,In_454);
nor U368 (N_368,In_131,In_332);
or U369 (N_369,In_199,In_60);
xor U370 (N_370,In_195,In_496);
nor U371 (N_371,In_178,In_59);
or U372 (N_372,In_496,In_405);
nand U373 (N_373,In_28,In_333);
xor U374 (N_374,In_60,In_374);
nor U375 (N_375,In_431,In_182);
or U376 (N_376,In_239,In_204);
or U377 (N_377,In_41,In_129);
nor U378 (N_378,In_417,In_28);
xnor U379 (N_379,In_358,In_352);
xor U380 (N_380,In_94,In_205);
nand U381 (N_381,In_66,In_104);
xnor U382 (N_382,In_197,In_91);
xor U383 (N_383,In_344,In_296);
nor U384 (N_384,In_307,In_21);
xnor U385 (N_385,In_331,In_93);
nor U386 (N_386,In_175,In_362);
xor U387 (N_387,In_216,In_310);
and U388 (N_388,In_452,In_37);
and U389 (N_389,In_221,In_145);
nand U390 (N_390,In_202,In_425);
and U391 (N_391,In_78,In_274);
or U392 (N_392,In_342,In_467);
nand U393 (N_393,In_426,In_196);
xor U394 (N_394,In_340,In_328);
and U395 (N_395,In_237,In_481);
or U396 (N_396,In_329,In_257);
or U397 (N_397,In_161,In_108);
and U398 (N_398,In_109,In_166);
nor U399 (N_399,In_381,In_496);
nand U400 (N_400,In_402,In_251);
and U401 (N_401,In_248,In_374);
xnor U402 (N_402,In_262,In_416);
or U403 (N_403,In_280,In_356);
and U404 (N_404,In_404,In_363);
and U405 (N_405,In_261,In_244);
xnor U406 (N_406,In_7,In_199);
and U407 (N_407,In_359,In_38);
nand U408 (N_408,In_177,In_226);
or U409 (N_409,In_457,In_81);
nand U410 (N_410,In_376,In_86);
nand U411 (N_411,In_189,In_39);
xnor U412 (N_412,In_397,In_252);
xnor U413 (N_413,In_374,In_473);
or U414 (N_414,In_184,In_495);
nor U415 (N_415,In_373,In_364);
and U416 (N_416,In_367,In_253);
nand U417 (N_417,In_176,In_419);
nand U418 (N_418,In_119,In_374);
or U419 (N_419,In_429,In_459);
nor U420 (N_420,In_450,In_427);
or U421 (N_421,In_395,In_3);
and U422 (N_422,In_436,In_454);
nand U423 (N_423,In_221,In_39);
and U424 (N_424,In_411,In_314);
nor U425 (N_425,In_222,In_156);
and U426 (N_426,In_253,In_183);
xnor U427 (N_427,In_389,In_134);
nor U428 (N_428,In_370,In_246);
nand U429 (N_429,In_155,In_113);
nand U430 (N_430,In_478,In_197);
and U431 (N_431,In_364,In_464);
nor U432 (N_432,In_206,In_487);
nand U433 (N_433,In_199,In_214);
and U434 (N_434,In_493,In_189);
nand U435 (N_435,In_2,In_169);
or U436 (N_436,In_442,In_213);
nand U437 (N_437,In_247,In_450);
or U438 (N_438,In_93,In_317);
nor U439 (N_439,In_310,In_244);
and U440 (N_440,In_392,In_322);
nand U441 (N_441,In_300,In_95);
and U442 (N_442,In_464,In_41);
xnor U443 (N_443,In_61,In_186);
and U444 (N_444,In_469,In_57);
and U445 (N_445,In_139,In_443);
xor U446 (N_446,In_116,In_348);
nand U447 (N_447,In_285,In_226);
nand U448 (N_448,In_365,In_430);
nand U449 (N_449,In_144,In_290);
xor U450 (N_450,In_119,In_231);
and U451 (N_451,In_46,In_348);
and U452 (N_452,In_320,In_223);
or U453 (N_453,In_130,In_274);
and U454 (N_454,In_228,In_401);
or U455 (N_455,In_201,In_123);
nand U456 (N_456,In_9,In_464);
xnor U457 (N_457,In_197,In_314);
nand U458 (N_458,In_342,In_480);
nor U459 (N_459,In_199,In_444);
or U460 (N_460,In_488,In_72);
nor U461 (N_461,In_263,In_316);
xnor U462 (N_462,In_267,In_480);
and U463 (N_463,In_212,In_112);
or U464 (N_464,In_458,In_397);
or U465 (N_465,In_322,In_468);
nor U466 (N_466,In_2,In_385);
or U467 (N_467,In_318,In_4);
nand U468 (N_468,In_57,In_373);
or U469 (N_469,In_51,In_14);
or U470 (N_470,In_267,In_146);
xnor U471 (N_471,In_261,In_347);
nor U472 (N_472,In_1,In_60);
nand U473 (N_473,In_385,In_243);
xnor U474 (N_474,In_136,In_65);
or U475 (N_475,In_158,In_295);
or U476 (N_476,In_103,In_193);
nor U477 (N_477,In_6,In_469);
or U478 (N_478,In_483,In_132);
nand U479 (N_479,In_484,In_389);
xnor U480 (N_480,In_316,In_387);
or U481 (N_481,In_177,In_481);
nand U482 (N_482,In_291,In_91);
and U483 (N_483,In_46,In_244);
nand U484 (N_484,In_363,In_72);
nor U485 (N_485,In_355,In_427);
or U486 (N_486,In_219,In_374);
nor U487 (N_487,In_354,In_70);
nand U488 (N_488,In_382,In_433);
or U489 (N_489,In_244,In_331);
and U490 (N_490,In_413,In_187);
nor U491 (N_491,In_299,In_67);
nand U492 (N_492,In_188,In_98);
nand U493 (N_493,In_226,In_101);
nand U494 (N_494,In_148,In_135);
xor U495 (N_495,In_200,In_61);
or U496 (N_496,In_316,In_34);
or U497 (N_497,In_389,In_182);
nor U498 (N_498,In_158,In_107);
or U499 (N_499,In_382,In_144);
xnor U500 (N_500,N_177,N_137);
or U501 (N_501,N_49,N_417);
nand U502 (N_502,N_243,N_469);
or U503 (N_503,N_377,N_165);
nand U504 (N_504,N_191,N_478);
nor U505 (N_505,N_351,N_363);
or U506 (N_506,N_322,N_2);
and U507 (N_507,N_483,N_34);
xnor U508 (N_508,N_442,N_43);
nor U509 (N_509,N_208,N_87);
nor U510 (N_510,N_11,N_79);
xor U511 (N_511,N_328,N_340);
nor U512 (N_512,N_314,N_124);
nor U513 (N_513,N_278,N_371);
nor U514 (N_514,N_212,N_323);
nor U515 (N_515,N_150,N_361);
nand U516 (N_516,N_65,N_309);
nand U517 (N_517,N_179,N_427);
or U518 (N_518,N_226,N_424);
nor U519 (N_519,N_345,N_160);
nand U520 (N_520,N_293,N_491);
and U521 (N_521,N_46,N_370);
and U522 (N_522,N_274,N_145);
nor U523 (N_523,N_285,N_105);
nand U524 (N_524,N_229,N_162);
nor U525 (N_525,N_471,N_227);
or U526 (N_526,N_462,N_142);
or U527 (N_527,N_288,N_214);
and U528 (N_528,N_44,N_178);
nor U529 (N_529,N_95,N_92);
nand U530 (N_530,N_331,N_453);
or U531 (N_531,N_460,N_433);
xor U532 (N_532,N_342,N_88);
and U533 (N_533,N_292,N_380);
or U534 (N_534,N_31,N_473);
nand U535 (N_535,N_441,N_174);
or U536 (N_536,N_76,N_385);
nor U537 (N_537,N_90,N_86);
nor U538 (N_538,N_176,N_402);
and U539 (N_539,N_121,N_362);
and U540 (N_540,N_480,N_72);
nand U541 (N_541,N_404,N_277);
nand U542 (N_542,N_476,N_415);
nor U543 (N_543,N_339,N_201);
nor U544 (N_544,N_194,N_24);
xnor U545 (N_545,N_263,N_437);
and U546 (N_546,N_461,N_467);
and U547 (N_547,N_470,N_167);
or U548 (N_548,N_390,N_5);
or U549 (N_549,N_329,N_446);
and U550 (N_550,N_439,N_42);
nand U551 (N_551,N_463,N_468);
and U552 (N_552,N_175,N_298);
xor U553 (N_553,N_225,N_33);
nor U554 (N_554,N_59,N_307);
and U555 (N_555,N_429,N_428);
nand U556 (N_556,N_399,N_364);
and U557 (N_557,N_130,N_222);
nor U558 (N_558,N_279,N_21);
xor U559 (N_559,N_154,N_400);
xnor U560 (N_560,N_382,N_305);
nand U561 (N_561,N_352,N_290);
nor U562 (N_562,N_356,N_324);
nor U563 (N_563,N_421,N_458);
nand U564 (N_564,N_37,N_66);
nor U565 (N_565,N_158,N_302);
xnor U566 (N_566,N_444,N_310);
nor U567 (N_567,N_268,N_258);
nand U568 (N_568,N_232,N_32);
or U569 (N_569,N_487,N_186);
or U570 (N_570,N_204,N_117);
and U571 (N_571,N_20,N_25);
nand U572 (N_572,N_109,N_239);
and U573 (N_573,N_347,N_112);
xnor U574 (N_574,N_113,N_29);
nand U575 (N_575,N_19,N_316);
xnor U576 (N_576,N_211,N_378);
or U577 (N_577,N_0,N_320);
or U578 (N_578,N_335,N_472);
nand U579 (N_579,N_182,N_271);
xnor U580 (N_580,N_57,N_251);
nor U581 (N_581,N_411,N_122);
or U582 (N_582,N_493,N_234);
xnor U583 (N_583,N_423,N_343);
xor U584 (N_584,N_485,N_389);
nand U585 (N_585,N_353,N_374);
nor U586 (N_586,N_17,N_63);
nand U587 (N_587,N_198,N_184);
and U588 (N_588,N_391,N_284);
or U589 (N_589,N_125,N_78);
and U590 (N_590,N_30,N_315);
and U591 (N_591,N_156,N_303);
nor U592 (N_592,N_357,N_187);
or U593 (N_593,N_242,N_200);
nand U594 (N_594,N_414,N_481);
nand U595 (N_595,N_344,N_143);
and U596 (N_596,N_321,N_236);
and U597 (N_597,N_252,N_383);
or U598 (N_598,N_368,N_101);
nor U599 (N_599,N_396,N_163);
nor U600 (N_600,N_71,N_70);
nand U601 (N_601,N_372,N_15);
and U602 (N_602,N_157,N_172);
or U603 (N_603,N_326,N_304);
nor U604 (N_604,N_98,N_448);
or U605 (N_605,N_35,N_373);
nor U606 (N_606,N_217,N_265);
or U607 (N_607,N_140,N_45);
and U608 (N_608,N_38,N_23);
nor U609 (N_609,N_492,N_419);
and U610 (N_610,N_40,N_431);
and U611 (N_611,N_151,N_132);
xor U612 (N_612,N_381,N_318);
or U613 (N_613,N_135,N_26);
nand U614 (N_614,N_349,N_202);
nor U615 (N_615,N_376,N_77);
and U616 (N_616,N_12,N_435);
or U617 (N_617,N_193,N_126);
or U618 (N_618,N_369,N_273);
xnor U619 (N_619,N_136,N_219);
xnor U620 (N_620,N_294,N_148);
and U621 (N_621,N_203,N_97);
nor U622 (N_622,N_41,N_188);
nand U623 (N_623,N_386,N_327);
or U624 (N_624,N_272,N_412);
or U625 (N_625,N_498,N_216);
and U626 (N_626,N_250,N_96);
xnor U627 (N_627,N_306,N_91);
nand U628 (N_628,N_133,N_459);
nor U629 (N_629,N_409,N_482);
or U630 (N_630,N_103,N_449);
nand U631 (N_631,N_300,N_262);
and U632 (N_632,N_489,N_287);
and U633 (N_633,N_276,N_183);
or U634 (N_634,N_289,N_281);
or U635 (N_635,N_248,N_367);
or U636 (N_636,N_210,N_260);
nand U637 (N_637,N_436,N_181);
nor U638 (N_638,N_333,N_106);
nand U639 (N_639,N_450,N_457);
nand U640 (N_640,N_283,N_416);
nor U641 (N_641,N_401,N_311);
and U642 (N_642,N_107,N_224);
nand U643 (N_643,N_440,N_240);
nand U644 (N_644,N_456,N_341);
nand U645 (N_645,N_169,N_313);
nand U646 (N_646,N_430,N_166);
or U647 (N_647,N_116,N_451);
and U648 (N_648,N_255,N_118);
and U649 (N_649,N_195,N_297);
nor U650 (N_650,N_330,N_479);
or U651 (N_651,N_64,N_379);
or U652 (N_652,N_308,N_149);
xor U653 (N_653,N_221,N_168);
and U654 (N_654,N_426,N_354);
xor U655 (N_655,N_68,N_319);
xnor U656 (N_656,N_244,N_3);
and U657 (N_657,N_388,N_6);
xnor U658 (N_658,N_54,N_397);
nor U659 (N_659,N_393,N_39);
nor U660 (N_660,N_185,N_408);
nand U661 (N_661,N_490,N_58);
xor U662 (N_662,N_334,N_53);
nor U663 (N_663,N_102,N_104);
nor U664 (N_664,N_83,N_13);
nor U665 (N_665,N_235,N_114);
nor U666 (N_666,N_443,N_259);
nand U667 (N_667,N_69,N_296);
xnor U668 (N_668,N_438,N_422);
or U669 (N_669,N_81,N_120);
nand U670 (N_670,N_218,N_407);
nor U671 (N_671,N_455,N_60);
or U672 (N_672,N_230,N_14);
nor U673 (N_673,N_360,N_199);
and U674 (N_674,N_223,N_161);
nand U675 (N_675,N_253,N_190);
or U676 (N_676,N_488,N_180);
nand U677 (N_677,N_261,N_466);
or U678 (N_678,N_358,N_475);
or U679 (N_679,N_61,N_445);
and U680 (N_680,N_220,N_134);
nand U681 (N_681,N_454,N_317);
xnor U682 (N_682,N_269,N_205);
xor U683 (N_683,N_67,N_85);
nor U684 (N_684,N_119,N_16);
xor U685 (N_685,N_425,N_7);
or U686 (N_686,N_375,N_171);
xor U687 (N_687,N_280,N_312);
xor U688 (N_688,N_275,N_256);
nand U689 (N_689,N_52,N_80);
nor U690 (N_690,N_432,N_93);
nor U691 (N_691,N_337,N_405);
and U692 (N_692,N_266,N_496);
nand U693 (N_693,N_153,N_325);
nand U694 (N_694,N_495,N_197);
and U695 (N_695,N_138,N_245);
xnor U696 (N_696,N_51,N_139);
xnor U697 (N_697,N_1,N_254);
xnor U698 (N_698,N_22,N_84);
nor U699 (N_699,N_247,N_420);
and U700 (N_700,N_332,N_62);
xnor U701 (N_701,N_50,N_147);
and U702 (N_702,N_27,N_155);
nand U703 (N_703,N_406,N_108);
and U704 (N_704,N_486,N_392);
nand U705 (N_705,N_9,N_173);
nor U706 (N_706,N_10,N_238);
nand U707 (N_707,N_301,N_56);
nand U708 (N_708,N_89,N_355);
xnor U709 (N_709,N_99,N_94);
nand U710 (N_710,N_336,N_249);
nor U711 (N_711,N_410,N_18);
xnor U712 (N_712,N_366,N_36);
nor U713 (N_713,N_128,N_127);
nor U714 (N_714,N_286,N_270);
or U715 (N_715,N_8,N_159);
nand U716 (N_716,N_233,N_164);
or U717 (N_717,N_291,N_189);
or U718 (N_718,N_47,N_494);
xor U719 (N_719,N_123,N_413);
and U720 (N_720,N_115,N_387);
or U721 (N_721,N_209,N_74);
nor U722 (N_722,N_231,N_246);
and U723 (N_723,N_338,N_477);
nor U724 (N_724,N_465,N_170);
nor U725 (N_725,N_257,N_131);
xnor U726 (N_726,N_144,N_73);
nand U727 (N_727,N_241,N_484);
and U728 (N_728,N_474,N_28);
nor U729 (N_729,N_152,N_206);
or U730 (N_730,N_237,N_348);
or U731 (N_731,N_82,N_213);
and U732 (N_732,N_100,N_264);
and U733 (N_733,N_499,N_228);
nand U734 (N_734,N_75,N_452);
xnor U735 (N_735,N_4,N_55);
nor U736 (N_736,N_282,N_359);
xnor U737 (N_737,N_111,N_464);
nand U738 (N_738,N_384,N_447);
nand U739 (N_739,N_192,N_299);
xnor U740 (N_740,N_110,N_196);
and U741 (N_741,N_395,N_207);
nor U742 (N_742,N_267,N_398);
and U743 (N_743,N_394,N_346);
or U744 (N_744,N_141,N_350);
xnor U745 (N_745,N_295,N_215);
or U746 (N_746,N_48,N_434);
nor U747 (N_747,N_403,N_365);
or U748 (N_748,N_418,N_497);
xnor U749 (N_749,N_146,N_129);
nor U750 (N_750,N_69,N_334);
nor U751 (N_751,N_76,N_362);
nand U752 (N_752,N_166,N_258);
nor U753 (N_753,N_147,N_497);
and U754 (N_754,N_370,N_75);
nor U755 (N_755,N_231,N_160);
xnor U756 (N_756,N_72,N_310);
nand U757 (N_757,N_201,N_117);
and U758 (N_758,N_431,N_139);
and U759 (N_759,N_153,N_101);
xnor U760 (N_760,N_326,N_331);
xor U761 (N_761,N_178,N_287);
or U762 (N_762,N_117,N_69);
nor U763 (N_763,N_363,N_42);
nor U764 (N_764,N_462,N_454);
or U765 (N_765,N_271,N_347);
nor U766 (N_766,N_335,N_455);
or U767 (N_767,N_262,N_37);
or U768 (N_768,N_319,N_217);
or U769 (N_769,N_404,N_103);
and U770 (N_770,N_472,N_374);
nand U771 (N_771,N_302,N_47);
nand U772 (N_772,N_44,N_273);
nand U773 (N_773,N_112,N_50);
or U774 (N_774,N_364,N_264);
nand U775 (N_775,N_340,N_142);
xor U776 (N_776,N_368,N_415);
nor U777 (N_777,N_139,N_183);
or U778 (N_778,N_134,N_332);
xor U779 (N_779,N_191,N_398);
and U780 (N_780,N_246,N_226);
nor U781 (N_781,N_23,N_2);
nor U782 (N_782,N_178,N_369);
nor U783 (N_783,N_465,N_236);
xor U784 (N_784,N_376,N_73);
nor U785 (N_785,N_492,N_350);
nand U786 (N_786,N_441,N_114);
and U787 (N_787,N_281,N_264);
nand U788 (N_788,N_116,N_70);
nand U789 (N_789,N_341,N_385);
xnor U790 (N_790,N_49,N_113);
and U791 (N_791,N_452,N_497);
nor U792 (N_792,N_20,N_400);
nor U793 (N_793,N_385,N_127);
nor U794 (N_794,N_134,N_384);
xnor U795 (N_795,N_369,N_171);
nand U796 (N_796,N_93,N_299);
nand U797 (N_797,N_382,N_2);
nand U798 (N_798,N_465,N_449);
and U799 (N_799,N_150,N_165);
nand U800 (N_800,N_48,N_311);
and U801 (N_801,N_185,N_149);
or U802 (N_802,N_306,N_253);
xor U803 (N_803,N_450,N_448);
or U804 (N_804,N_120,N_14);
xor U805 (N_805,N_379,N_53);
xor U806 (N_806,N_72,N_289);
nor U807 (N_807,N_444,N_24);
and U808 (N_808,N_140,N_350);
nor U809 (N_809,N_116,N_165);
and U810 (N_810,N_308,N_168);
or U811 (N_811,N_212,N_327);
nand U812 (N_812,N_267,N_181);
nand U813 (N_813,N_181,N_150);
and U814 (N_814,N_219,N_316);
nand U815 (N_815,N_121,N_135);
xnor U816 (N_816,N_186,N_387);
and U817 (N_817,N_444,N_179);
or U818 (N_818,N_290,N_71);
xnor U819 (N_819,N_379,N_286);
or U820 (N_820,N_36,N_158);
xnor U821 (N_821,N_439,N_80);
nor U822 (N_822,N_270,N_117);
xnor U823 (N_823,N_472,N_315);
nand U824 (N_824,N_224,N_37);
nand U825 (N_825,N_339,N_306);
nand U826 (N_826,N_180,N_177);
and U827 (N_827,N_204,N_339);
or U828 (N_828,N_342,N_196);
or U829 (N_829,N_164,N_158);
or U830 (N_830,N_45,N_385);
xnor U831 (N_831,N_287,N_148);
and U832 (N_832,N_205,N_100);
nor U833 (N_833,N_54,N_212);
nand U834 (N_834,N_397,N_87);
and U835 (N_835,N_352,N_238);
and U836 (N_836,N_202,N_77);
or U837 (N_837,N_282,N_160);
or U838 (N_838,N_149,N_215);
nor U839 (N_839,N_205,N_412);
nand U840 (N_840,N_136,N_77);
or U841 (N_841,N_376,N_223);
nor U842 (N_842,N_106,N_86);
xor U843 (N_843,N_191,N_366);
nor U844 (N_844,N_106,N_393);
xnor U845 (N_845,N_239,N_139);
nand U846 (N_846,N_483,N_98);
nor U847 (N_847,N_70,N_230);
nand U848 (N_848,N_210,N_456);
nor U849 (N_849,N_238,N_270);
xnor U850 (N_850,N_419,N_238);
xor U851 (N_851,N_155,N_24);
and U852 (N_852,N_320,N_453);
nor U853 (N_853,N_226,N_220);
xor U854 (N_854,N_450,N_386);
and U855 (N_855,N_374,N_157);
and U856 (N_856,N_318,N_379);
nand U857 (N_857,N_226,N_339);
xnor U858 (N_858,N_257,N_36);
xnor U859 (N_859,N_436,N_467);
nor U860 (N_860,N_296,N_374);
nor U861 (N_861,N_211,N_236);
or U862 (N_862,N_474,N_493);
and U863 (N_863,N_367,N_106);
and U864 (N_864,N_244,N_410);
or U865 (N_865,N_112,N_156);
and U866 (N_866,N_487,N_471);
xor U867 (N_867,N_258,N_450);
nand U868 (N_868,N_112,N_455);
and U869 (N_869,N_458,N_15);
nand U870 (N_870,N_328,N_179);
and U871 (N_871,N_387,N_455);
nand U872 (N_872,N_220,N_395);
nand U873 (N_873,N_94,N_220);
nor U874 (N_874,N_47,N_1);
xor U875 (N_875,N_339,N_316);
nand U876 (N_876,N_58,N_80);
nand U877 (N_877,N_363,N_208);
nor U878 (N_878,N_9,N_454);
and U879 (N_879,N_354,N_3);
and U880 (N_880,N_274,N_115);
nand U881 (N_881,N_102,N_240);
nand U882 (N_882,N_480,N_63);
or U883 (N_883,N_288,N_28);
xnor U884 (N_884,N_452,N_170);
and U885 (N_885,N_305,N_168);
nand U886 (N_886,N_80,N_275);
xor U887 (N_887,N_85,N_140);
nand U888 (N_888,N_279,N_122);
and U889 (N_889,N_462,N_166);
nor U890 (N_890,N_264,N_220);
nand U891 (N_891,N_351,N_382);
or U892 (N_892,N_281,N_151);
nor U893 (N_893,N_254,N_381);
nand U894 (N_894,N_384,N_312);
nand U895 (N_895,N_104,N_33);
nor U896 (N_896,N_68,N_417);
and U897 (N_897,N_462,N_317);
xnor U898 (N_898,N_293,N_288);
and U899 (N_899,N_70,N_15);
xor U900 (N_900,N_246,N_353);
or U901 (N_901,N_82,N_138);
nand U902 (N_902,N_134,N_464);
or U903 (N_903,N_316,N_119);
or U904 (N_904,N_380,N_88);
xnor U905 (N_905,N_224,N_113);
or U906 (N_906,N_416,N_90);
nor U907 (N_907,N_180,N_350);
or U908 (N_908,N_280,N_324);
nor U909 (N_909,N_404,N_58);
and U910 (N_910,N_496,N_465);
xor U911 (N_911,N_239,N_148);
nand U912 (N_912,N_67,N_347);
or U913 (N_913,N_271,N_137);
xnor U914 (N_914,N_450,N_123);
xor U915 (N_915,N_310,N_321);
nor U916 (N_916,N_330,N_442);
or U917 (N_917,N_8,N_79);
and U918 (N_918,N_51,N_119);
or U919 (N_919,N_388,N_325);
nand U920 (N_920,N_388,N_28);
xor U921 (N_921,N_304,N_123);
nor U922 (N_922,N_455,N_412);
or U923 (N_923,N_38,N_181);
or U924 (N_924,N_385,N_309);
xor U925 (N_925,N_372,N_383);
nand U926 (N_926,N_268,N_264);
and U927 (N_927,N_64,N_495);
xor U928 (N_928,N_410,N_42);
nand U929 (N_929,N_74,N_472);
nor U930 (N_930,N_464,N_35);
nand U931 (N_931,N_412,N_227);
or U932 (N_932,N_310,N_165);
or U933 (N_933,N_27,N_354);
nand U934 (N_934,N_5,N_212);
nor U935 (N_935,N_204,N_149);
or U936 (N_936,N_153,N_17);
xor U937 (N_937,N_232,N_392);
or U938 (N_938,N_230,N_191);
xnor U939 (N_939,N_386,N_64);
or U940 (N_940,N_156,N_400);
or U941 (N_941,N_361,N_430);
and U942 (N_942,N_355,N_34);
or U943 (N_943,N_38,N_107);
or U944 (N_944,N_85,N_218);
nand U945 (N_945,N_200,N_186);
nor U946 (N_946,N_343,N_60);
xor U947 (N_947,N_483,N_3);
nand U948 (N_948,N_229,N_68);
nor U949 (N_949,N_60,N_271);
and U950 (N_950,N_233,N_28);
nor U951 (N_951,N_104,N_350);
nor U952 (N_952,N_398,N_224);
nand U953 (N_953,N_228,N_161);
and U954 (N_954,N_55,N_102);
xor U955 (N_955,N_167,N_198);
and U956 (N_956,N_483,N_216);
and U957 (N_957,N_152,N_175);
nand U958 (N_958,N_40,N_72);
or U959 (N_959,N_389,N_427);
or U960 (N_960,N_74,N_395);
and U961 (N_961,N_293,N_499);
and U962 (N_962,N_352,N_38);
xnor U963 (N_963,N_133,N_489);
nand U964 (N_964,N_448,N_482);
or U965 (N_965,N_176,N_368);
nand U966 (N_966,N_471,N_317);
and U967 (N_967,N_383,N_285);
nor U968 (N_968,N_497,N_89);
xor U969 (N_969,N_260,N_395);
xor U970 (N_970,N_148,N_102);
nand U971 (N_971,N_177,N_381);
nor U972 (N_972,N_432,N_227);
nand U973 (N_973,N_477,N_358);
and U974 (N_974,N_288,N_179);
xor U975 (N_975,N_259,N_26);
nor U976 (N_976,N_147,N_103);
xor U977 (N_977,N_316,N_42);
and U978 (N_978,N_80,N_5);
xnor U979 (N_979,N_48,N_59);
nand U980 (N_980,N_472,N_483);
or U981 (N_981,N_33,N_442);
nor U982 (N_982,N_268,N_110);
nor U983 (N_983,N_447,N_279);
and U984 (N_984,N_46,N_395);
nand U985 (N_985,N_405,N_328);
or U986 (N_986,N_330,N_299);
and U987 (N_987,N_181,N_45);
nor U988 (N_988,N_369,N_283);
xor U989 (N_989,N_297,N_64);
nor U990 (N_990,N_135,N_441);
or U991 (N_991,N_147,N_106);
xor U992 (N_992,N_424,N_468);
nor U993 (N_993,N_448,N_65);
and U994 (N_994,N_137,N_305);
nand U995 (N_995,N_471,N_461);
and U996 (N_996,N_430,N_473);
or U997 (N_997,N_238,N_155);
and U998 (N_998,N_467,N_386);
nor U999 (N_999,N_402,N_423);
or U1000 (N_1000,N_774,N_911);
xor U1001 (N_1001,N_882,N_540);
nand U1002 (N_1002,N_574,N_703);
nor U1003 (N_1003,N_735,N_765);
and U1004 (N_1004,N_707,N_744);
or U1005 (N_1005,N_616,N_661);
xnor U1006 (N_1006,N_965,N_558);
xnor U1007 (N_1007,N_657,N_914);
xor U1008 (N_1008,N_821,N_983);
xor U1009 (N_1009,N_981,N_739);
nor U1010 (N_1010,N_581,N_811);
xor U1011 (N_1011,N_857,N_923);
xnor U1012 (N_1012,N_942,N_876);
and U1013 (N_1013,N_918,N_879);
nand U1014 (N_1014,N_763,N_659);
or U1015 (N_1015,N_837,N_963);
nand U1016 (N_1016,N_673,N_782);
xnor U1017 (N_1017,N_714,N_897);
nor U1018 (N_1018,N_937,N_621);
nor U1019 (N_1019,N_589,N_600);
and U1020 (N_1020,N_627,N_900);
and U1021 (N_1021,N_881,N_772);
or U1022 (N_1022,N_802,N_781);
or U1023 (N_1023,N_929,N_531);
and U1024 (N_1024,N_972,N_688);
and U1025 (N_1025,N_896,N_947);
and U1026 (N_1026,N_509,N_518);
nor U1027 (N_1027,N_526,N_788);
or U1028 (N_1028,N_685,N_928);
or U1029 (N_1029,N_532,N_738);
xnor U1030 (N_1030,N_804,N_751);
nor U1031 (N_1031,N_587,N_592);
nor U1032 (N_1032,N_962,N_873);
or U1033 (N_1033,N_836,N_579);
nor U1034 (N_1034,N_790,N_733);
xor U1035 (N_1035,N_718,N_550);
or U1036 (N_1036,N_976,N_995);
or U1037 (N_1037,N_800,N_986);
xnor U1038 (N_1038,N_954,N_604);
xnor U1039 (N_1039,N_985,N_868);
nor U1040 (N_1040,N_823,N_646);
nor U1041 (N_1041,N_538,N_553);
and U1042 (N_1042,N_867,N_708);
and U1043 (N_1043,N_737,N_694);
nor U1044 (N_1044,N_752,N_905);
nor U1045 (N_1045,N_885,N_731);
nor U1046 (N_1046,N_910,N_671);
nor U1047 (N_1047,N_945,N_520);
or U1048 (N_1048,N_617,N_826);
nor U1049 (N_1049,N_960,N_663);
or U1050 (N_1050,N_852,N_562);
nand U1051 (N_1051,N_555,N_794);
xor U1052 (N_1052,N_920,N_583);
xnor U1053 (N_1053,N_597,N_530);
and U1054 (N_1054,N_634,N_511);
xnor U1055 (N_1055,N_813,N_869);
xnor U1056 (N_1056,N_808,N_570);
xor U1057 (N_1057,N_931,N_761);
nand U1058 (N_1058,N_969,N_590);
or U1059 (N_1059,N_796,N_950);
and U1060 (N_1060,N_717,N_620);
and U1061 (N_1061,N_878,N_537);
and U1062 (N_1062,N_818,N_567);
or U1063 (N_1063,N_771,N_814);
or U1064 (N_1064,N_750,N_948);
xor U1065 (N_1065,N_599,N_510);
xnor U1066 (N_1066,N_596,N_809);
nor U1067 (N_1067,N_638,N_593);
nor U1068 (N_1068,N_877,N_670);
or U1069 (N_1069,N_952,N_640);
and U1070 (N_1070,N_647,N_594);
and U1071 (N_1071,N_668,N_702);
nand U1072 (N_1072,N_568,N_767);
nand U1073 (N_1073,N_777,N_979);
xor U1074 (N_1074,N_564,N_504);
nor U1075 (N_1075,N_618,N_854);
or U1076 (N_1076,N_660,N_633);
nor U1077 (N_1077,N_909,N_609);
or U1078 (N_1078,N_501,N_541);
xnor U1079 (N_1079,N_825,N_623);
nand U1080 (N_1080,N_643,N_619);
nand U1081 (N_1081,N_850,N_613);
xor U1082 (N_1082,N_999,N_833);
and U1083 (N_1083,N_791,N_552);
and U1084 (N_1084,N_803,N_631);
or U1085 (N_1085,N_667,N_921);
xor U1086 (N_1086,N_758,N_637);
nand U1087 (N_1087,N_806,N_687);
nor U1088 (N_1088,N_724,N_658);
nor U1089 (N_1089,N_817,N_628);
nor U1090 (N_1090,N_514,N_560);
nand U1091 (N_1091,N_513,N_603);
and U1092 (N_1092,N_644,N_539);
or U1093 (N_1093,N_700,N_901);
xor U1094 (N_1094,N_893,N_548);
and U1095 (N_1095,N_994,N_815);
xnor U1096 (N_1096,N_582,N_624);
and U1097 (N_1097,N_614,N_684);
or U1098 (N_1098,N_875,N_768);
nor U1099 (N_1099,N_528,N_743);
or U1100 (N_1100,N_917,N_515);
and U1101 (N_1101,N_899,N_545);
nor U1102 (N_1102,N_784,N_829);
or U1103 (N_1103,N_968,N_760);
nor U1104 (N_1104,N_536,N_561);
nand U1105 (N_1105,N_810,N_840);
or U1106 (N_1106,N_672,N_629);
and U1107 (N_1107,N_892,N_522);
nor U1108 (N_1108,N_874,N_753);
or U1109 (N_1109,N_778,N_748);
and U1110 (N_1110,N_828,N_697);
or U1111 (N_1111,N_819,N_862);
or U1112 (N_1112,N_723,N_853);
and U1113 (N_1113,N_535,N_502);
and U1114 (N_1114,N_525,N_542);
or U1115 (N_1115,N_679,N_680);
and U1116 (N_1116,N_681,N_891);
and U1117 (N_1117,N_576,N_678);
nand U1118 (N_1118,N_725,N_785);
nand U1119 (N_1119,N_615,N_636);
nor U1120 (N_1120,N_849,N_769);
nand U1121 (N_1121,N_984,N_523);
nor U1122 (N_1122,N_861,N_730);
or U1123 (N_1123,N_726,N_866);
or U1124 (N_1124,N_958,N_557);
nor U1125 (N_1125,N_653,N_927);
nand U1126 (N_1126,N_719,N_505);
nand U1127 (N_1127,N_706,N_851);
xor U1128 (N_1128,N_699,N_951);
nand U1129 (N_1129,N_773,N_512);
or U1130 (N_1130,N_898,N_895);
nor U1131 (N_1131,N_789,N_838);
nand U1132 (N_1132,N_569,N_605);
nor U1133 (N_1133,N_641,N_792);
nor U1134 (N_1134,N_872,N_871);
nor U1135 (N_1135,N_727,N_938);
xnor U1136 (N_1136,N_775,N_559);
xnor U1137 (N_1137,N_507,N_766);
or U1138 (N_1138,N_656,N_747);
nand U1139 (N_1139,N_575,N_683);
nand U1140 (N_1140,N_662,N_770);
nor U1141 (N_1141,N_830,N_695);
nand U1142 (N_1142,N_585,N_577);
nand U1143 (N_1143,N_722,N_588);
or U1144 (N_1144,N_630,N_648);
nor U1145 (N_1145,N_936,N_903);
nand U1146 (N_1146,N_529,N_941);
or U1147 (N_1147,N_692,N_906);
nor U1148 (N_1148,N_508,N_988);
and U1149 (N_1149,N_610,N_759);
nor U1150 (N_1150,N_991,N_676);
xnor U1151 (N_1151,N_940,N_915);
xnor U1152 (N_1152,N_930,N_908);
nor U1153 (N_1153,N_654,N_797);
xnor U1154 (N_1154,N_956,N_664);
and U1155 (N_1155,N_556,N_847);
xnor U1156 (N_1156,N_527,N_601);
and U1157 (N_1157,N_865,N_544);
and U1158 (N_1158,N_964,N_578);
and U1159 (N_1159,N_801,N_749);
or U1160 (N_1160,N_953,N_889);
or U1161 (N_1161,N_736,N_690);
and U1162 (N_1162,N_608,N_939);
nand U1163 (N_1163,N_632,N_798);
xnor U1164 (N_1164,N_543,N_689);
or U1165 (N_1165,N_966,N_902);
nor U1166 (N_1166,N_682,N_551);
xnor U1167 (N_1167,N_563,N_572);
or U1168 (N_1168,N_884,N_888);
nand U1169 (N_1169,N_715,N_669);
nand U1170 (N_1170,N_907,N_955);
nand U1171 (N_1171,N_500,N_844);
nor U1172 (N_1172,N_860,N_704);
nor U1173 (N_1173,N_977,N_916);
xor U1174 (N_1174,N_611,N_580);
or U1175 (N_1175,N_859,N_845);
nor U1176 (N_1176,N_649,N_586);
nand U1177 (N_1177,N_754,N_573);
or U1178 (N_1178,N_701,N_602);
xnor U1179 (N_1179,N_705,N_971);
and U1180 (N_1180,N_639,N_795);
or U1181 (N_1181,N_989,N_807);
nand U1182 (N_1182,N_645,N_742);
or U1183 (N_1183,N_606,N_932);
nand U1184 (N_1184,N_741,N_665);
xnor U1185 (N_1185,N_924,N_858);
xnor U1186 (N_1186,N_547,N_549);
xor U1187 (N_1187,N_831,N_696);
nor U1188 (N_1188,N_622,N_846);
or U1189 (N_1189,N_880,N_762);
or U1190 (N_1190,N_674,N_934);
and U1191 (N_1191,N_721,N_970);
xnor U1192 (N_1192,N_776,N_812);
or U1193 (N_1193,N_787,N_728);
and U1194 (N_1194,N_843,N_799);
nand U1195 (N_1195,N_793,N_841);
nand U1196 (N_1196,N_835,N_961);
nor U1197 (N_1197,N_516,N_975);
and U1198 (N_1198,N_650,N_677);
or U1199 (N_1199,N_863,N_651);
or U1200 (N_1200,N_534,N_805);
or U1201 (N_1201,N_978,N_584);
nor U1202 (N_1202,N_713,N_820);
xnor U1203 (N_1203,N_720,N_712);
and U1204 (N_1204,N_887,N_925);
nor U1205 (N_1205,N_710,N_993);
nand U1206 (N_1206,N_635,N_943);
xor U1207 (N_1207,N_959,N_894);
or U1208 (N_1208,N_834,N_565);
and U1209 (N_1209,N_982,N_946);
xnor U1210 (N_1210,N_729,N_595);
nor U1211 (N_1211,N_990,N_691);
nand U1212 (N_1212,N_693,N_933);
or U1213 (N_1213,N_944,N_827);
nor U1214 (N_1214,N_655,N_949);
xor U1215 (N_1215,N_842,N_612);
and U1216 (N_1216,N_716,N_913);
and U1217 (N_1217,N_524,N_554);
xor U1218 (N_1218,N_839,N_566);
nand U1219 (N_1219,N_686,N_957);
or U1220 (N_1220,N_732,N_864);
or U1221 (N_1221,N_591,N_832);
xnor U1222 (N_1222,N_519,N_625);
or U1223 (N_1223,N_997,N_571);
nand U1224 (N_1224,N_992,N_786);
xor U1225 (N_1225,N_974,N_607);
or U1226 (N_1226,N_848,N_890);
xor U1227 (N_1227,N_666,N_745);
xor U1228 (N_1228,N_919,N_746);
or U1229 (N_1229,N_756,N_517);
and U1230 (N_1230,N_740,N_870);
nor U1231 (N_1231,N_855,N_922);
or U1232 (N_1232,N_987,N_652);
nor U1233 (N_1233,N_711,N_816);
or U1234 (N_1234,N_886,N_967);
and U1235 (N_1235,N_503,N_675);
nand U1236 (N_1236,N_709,N_698);
and U1237 (N_1237,N_521,N_973);
nor U1238 (N_1238,N_734,N_912);
or U1239 (N_1239,N_626,N_926);
xnor U1240 (N_1240,N_642,N_904);
nand U1241 (N_1241,N_598,N_980);
xor U1242 (N_1242,N_779,N_764);
and U1243 (N_1243,N_755,N_783);
and U1244 (N_1244,N_822,N_533);
nand U1245 (N_1245,N_883,N_546);
nor U1246 (N_1246,N_996,N_824);
nand U1247 (N_1247,N_998,N_780);
and U1248 (N_1248,N_506,N_935);
nor U1249 (N_1249,N_856,N_757);
nand U1250 (N_1250,N_771,N_970);
xor U1251 (N_1251,N_764,N_897);
nor U1252 (N_1252,N_927,N_738);
nand U1253 (N_1253,N_666,N_782);
and U1254 (N_1254,N_554,N_541);
nand U1255 (N_1255,N_667,N_589);
or U1256 (N_1256,N_887,N_770);
and U1257 (N_1257,N_509,N_724);
nand U1258 (N_1258,N_548,N_731);
or U1259 (N_1259,N_971,N_562);
xnor U1260 (N_1260,N_528,N_527);
nor U1261 (N_1261,N_953,N_635);
or U1262 (N_1262,N_529,N_909);
and U1263 (N_1263,N_794,N_928);
xnor U1264 (N_1264,N_813,N_973);
xnor U1265 (N_1265,N_932,N_944);
or U1266 (N_1266,N_576,N_764);
and U1267 (N_1267,N_853,N_800);
or U1268 (N_1268,N_554,N_931);
xor U1269 (N_1269,N_903,N_695);
and U1270 (N_1270,N_551,N_919);
or U1271 (N_1271,N_556,N_904);
xnor U1272 (N_1272,N_958,N_983);
nor U1273 (N_1273,N_982,N_524);
xor U1274 (N_1274,N_818,N_751);
or U1275 (N_1275,N_974,N_656);
or U1276 (N_1276,N_554,N_688);
xor U1277 (N_1277,N_875,N_983);
or U1278 (N_1278,N_913,N_713);
and U1279 (N_1279,N_876,N_944);
or U1280 (N_1280,N_573,N_794);
or U1281 (N_1281,N_713,N_675);
and U1282 (N_1282,N_766,N_912);
nor U1283 (N_1283,N_818,N_951);
and U1284 (N_1284,N_634,N_628);
xor U1285 (N_1285,N_647,N_868);
nand U1286 (N_1286,N_678,N_864);
and U1287 (N_1287,N_517,N_761);
nand U1288 (N_1288,N_761,N_803);
nor U1289 (N_1289,N_967,N_561);
nor U1290 (N_1290,N_908,N_974);
nand U1291 (N_1291,N_572,N_671);
xor U1292 (N_1292,N_845,N_541);
xor U1293 (N_1293,N_501,N_704);
xor U1294 (N_1294,N_964,N_558);
or U1295 (N_1295,N_993,N_815);
xor U1296 (N_1296,N_541,N_534);
nand U1297 (N_1297,N_577,N_816);
xnor U1298 (N_1298,N_934,N_586);
nor U1299 (N_1299,N_680,N_592);
nor U1300 (N_1300,N_733,N_599);
and U1301 (N_1301,N_656,N_979);
nor U1302 (N_1302,N_976,N_765);
nand U1303 (N_1303,N_756,N_737);
or U1304 (N_1304,N_644,N_771);
and U1305 (N_1305,N_756,N_677);
and U1306 (N_1306,N_845,N_742);
nand U1307 (N_1307,N_623,N_893);
and U1308 (N_1308,N_819,N_769);
nor U1309 (N_1309,N_543,N_981);
xor U1310 (N_1310,N_944,N_727);
nand U1311 (N_1311,N_790,N_578);
xnor U1312 (N_1312,N_685,N_831);
xnor U1313 (N_1313,N_622,N_660);
nor U1314 (N_1314,N_742,N_981);
xnor U1315 (N_1315,N_925,N_787);
nand U1316 (N_1316,N_748,N_671);
nor U1317 (N_1317,N_892,N_653);
nand U1318 (N_1318,N_583,N_862);
and U1319 (N_1319,N_956,N_683);
and U1320 (N_1320,N_835,N_705);
nor U1321 (N_1321,N_802,N_846);
nand U1322 (N_1322,N_711,N_623);
nand U1323 (N_1323,N_998,N_867);
nor U1324 (N_1324,N_590,N_511);
and U1325 (N_1325,N_738,N_674);
xnor U1326 (N_1326,N_792,N_974);
nand U1327 (N_1327,N_983,N_769);
xor U1328 (N_1328,N_946,N_805);
nor U1329 (N_1329,N_628,N_962);
or U1330 (N_1330,N_545,N_705);
nor U1331 (N_1331,N_708,N_825);
xor U1332 (N_1332,N_689,N_841);
nand U1333 (N_1333,N_612,N_698);
nand U1334 (N_1334,N_932,N_598);
xor U1335 (N_1335,N_829,N_736);
or U1336 (N_1336,N_854,N_578);
and U1337 (N_1337,N_539,N_928);
nand U1338 (N_1338,N_579,N_504);
xor U1339 (N_1339,N_675,N_994);
nand U1340 (N_1340,N_730,N_859);
nand U1341 (N_1341,N_627,N_724);
nand U1342 (N_1342,N_998,N_725);
nand U1343 (N_1343,N_595,N_856);
xnor U1344 (N_1344,N_686,N_774);
and U1345 (N_1345,N_748,N_853);
nor U1346 (N_1346,N_876,N_615);
nand U1347 (N_1347,N_847,N_638);
and U1348 (N_1348,N_958,N_791);
or U1349 (N_1349,N_978,N_737);
and U1350 (N_1350,N_576,N_527);
or U1351 (N_1351,N_884,N_984);
and U1352 (N_1352,N_521,N_745);
nand U1353 (N_1353,N_727,N_556);
or U1354 (N_1354,N_586,N_551);
xnor U1355 (N_1355,N_894,N_722);
or U1356 (N_1356,N_712,N_577);
or U1357 (N_1357,N_700,N_873);
nand U1358 (N_1358,N_749,N_567);
and U1359 (N_1359,N_757,N_672);
nor U1360 (N_1360,N_775,N_908);
nand U1361 (N_1361,N_561,N_713);
or U1362 (N_1362,N_930,N_664);
or U1363 (N_1363,N_613,N_883);
xnor U1364 (N_1364,N_866,N_778);
and U1365 (N_1365,N_527,N_540);
xnor U1366 (N_1366,N_749,N_573);
nor U1367 (N_1367,N_949,N_686);
nand U1368 (N_1368,N_813,N_584);
nor U1369 (N_1369,N_827,N_617);
nand U1370 (N_1370,N_898,N_529);
nand U1371 (N_1371,N_985,N_811);
and U1372 (N_1372,N_781,N_986);
and U1373 (N_1373,N_701,N_507);
nor U1374 (N_1374,N_953,N_506);
or U1375 (N_1375,N_558,N_814);
nor U1376 (N_1376,N_679,N_737);
or U1377 (N_1377,N_916,N_531);
xnor U1378 (N_1378,N_544,N_521);
nand U1379 (N_1379,N_651,N_927);
xnor U1380 (N_1380,N_811,N_818);
xnor U1381 (N_1381,N_799,N_934);
and U1382 (N_1382,N_631,N_802);
nand U1383 (N_1383,N_754,N_905);
nor U1384 (N_1384,N_525,N_653);
nor U1385 (N_1385,N_949,N_863);
xnor U1386 (N_1386,N_833,N_821);
or U1387 (N_1387,N_732,N_692);
nand U1388 (N_1388,N_952,N_845);
nand U1389 (N_1389,N_736,N_846);
nor U1390 (N_1390,N_591,N_902);
or U1391 (N_1391,N_705,N_872);
nor U1392 (N_1392,N_965,N_813);
and U1393 (N_1393,N_659,N_616);
nand U1394 (N_1394,N_923,N_823);
nor U1395 (N_1395,N_641,N_652);
nor U1396 (N_1396,N_974,N_560);
nand U1397 (N_1397,N_942,N_982);
nand U1398 (N_1398,N_541,N_985);
and U1399 (N_1399,N_566,N_901);
or U1400 (N_1400,N_962,N_631);
xnor U1401 (N_1401,N_911,N_782);
and U1402 (N_1402,N_791,N_556);
nand U1403 (N_1403,N_562,N_948);
xnor U1404 (N_1404,N_819,N_628);
nand U1405 (N_1405,N_620,N_989);
xnor U1406 (N_1406,N_571,N_923);
xnor U1407 (N_1407,N_821,N_876);
nand U1408 (N_1408,N_856,N_677);
xor U1409 (N_1409,N_639,N_994);
nand U1410 (N_1410,N_674,N_576);
xor U1411 (N_1411,N_559,N_674);
nand U1412 (N_1412,N_774,N_872);
nand U1413 (N_1413,N_667,N_608);
nor U1414 (N_1414,N_772,N_579);
nor U1415 (N_1415,N_830,N_846);
nor U1416 (N_1416,N_527,N_590);
and U1417 (N_1417,N_645,N_793);
or U1418 (N_1418,N_656,N_918);
xnor U1419 (N_1419,N_576,N_540);
nor U1420 (N_1420,N_711,N_788);
and U1421 (N_1421,N_758,N_961);
nand U1422 (N_1422,N_523,N_825);
xnor U1423 (N_1423,N_767,N_662);
or U1424 (N_1424,N_931,N_894);
nor U1425 (N_1425,N_579,N_835);
nand U1426 (N_1426,N_561,N_564);
and U1427 (N_1427,N_536,N_966);
or U1428 (N_1428,N_950,N_516);
nor U1429 (N_1429,N_850,N_657);
and U1430 (N_1430,N_685,N_502);
or U1431 (N_1431,N_697,N_898);
or U1432 (N_1432,N_638,N_768);
or U1433 (N_1433,N_761,N_536);
or U1434 (N_1434,N_850,N_837);
xnor U1435 (N_1435,N_876,N_532);
nand U1436 (N_1436,N_691,N_690);
nor U1437 (N_1437,N_601,N_512);
nand U1438 (N_1438,N_998,N_832);
and U1439 (N_1439,N_502,N_766);
and U1440 (N_1440,N_697,N_511);
nor U1441 (N_1441,N_798,N_563);
and U1442 (N_1442,N_805,N_808);
or U1443 (N_1443,N_533,N_660);
nand U1444 (N_1444,N_614,N_631);
and U1445 (N_1445,N_975,N_935);
nor U1446 (N_1446,N_568,N_538);
xnor U1447 (N_1447,N_686,N_753);
nor U1448 (N_1448,N_669,N_514);
xor U1449 (N_1449,N_824,N_648);
or U1450 (N_1450,N_770,N_820);
xor U1451 (N_1451,N_767,N_814);
xor U1452 (N_1452,N_946,N_830);
nor U1453 (N_1453,N_591,N_904);
and U1454 (N_1454,N_591,N_522);
or U1455 (N_1455,N_737,N_943);
or U1456 (N_1456,N_979,N_913);
and U1457 (N_1457,N_541,N_511);
nor U1458 (N_1458,N_550,N_851);
nor U1459 (N_1459,N_596,N_623);
nor U1460 (N_1460,N_788,N_634);
xnor U1461 (N_1461,N_591,N_659);
nor U1462 (N_1462,N_936,N_649);
and U1463 (N_1463,N_921,N_862);
nand U1464 (N_1464,N_722,N_932);
nand U1465 (N_1465,N_628,N_514);
or U1466 (N_1466,N_735,N_745);
nor U1467 (N_1467,N_631,N_706);
nor U1468 (N_1468,N_606,N_870);
xnor U1469 (N_1469,N_728,N_689);
xor U1470 (N_1470,N_912,N_927);
and U1471 (N_1471,N_665,N_916);
nand U1472 (N_1472,N_909,N_522);
xor U1473 (N_1473,N_890,N_870);
or U1474 (N_1474,N_509,N_558);
nand U1475 (N_1475,N_633,N_585);
nor U1476 (N_1476,N_792,N_899);
xnor U1477 (N_1477,N_935,N_968);
nand U1478 (N_1478,N_891,N_911);
nand U1479 (N_1479,N_663,N_540);
nand U1480 (N_1480,N_826,N_839);
nand U1481 (N_1481,N_567,N_821);
xnor U1482 (N_1482,N_813,N_702);
and U1483 (N_1483,N_549,N_835);
or U1484 (N_1484,N_950,N_944);
xor U1485 (N_1485,N_837,N_769);
xnor U1486 (N_1486,N_706,N_531);
xnor U1487 (N_1487,N_732,N_542);
and U1488 (N_1488,N_873,N_963);
or U1489 (N_1489,N_684,N_631);
xor U1490 (N_1490,N_616,N_729);
nor U1491 (N_1491,N_522,N_928);
xnor U1492 (N_1492,N_506,N_721);
nor U1493 (N_1493,N_532,N_859);
or U1494 (N_1494,N_700,N_547);
nand U1495 (N_1495,N_790,N_716);
nor U1496 (N_1496,N_570,N_776);
and U1497 (N_1497,N_899,N_658);
or U1498 (N_1498,N_777,N_933);
or U1499 (N_1499,N_853,N_788);
or U1500 (N_1500,N_1387,N_1124);
nand U1501 (N_1501,N_1171,N_1095);
nor U1502 (N_1502,N_1212,N_1037);
nor U1503 (N_1503,N_1316,N_1254);
xor U1504 (N_1504,N_1275,N_1063);
nor U1505 (N_1505,N_1065,N_1202);
and U1506 (N_1506,N_1240,N_1201);
nor U1507 (N_1507,N_1468,N_1229);
nor U1508 (N_1508,N_1239,N_1173);
or U1509 (N_1509,N_1474,N_1439);
or U1510 (N_1510,N_1121,N_1047);
and U1511 (N_1511,N_1315,N_1114);
xor U1512 (N_1512,N_1139,N_1306);
or U1513 (N_1513,N_1347,N_1192);
and U1514 (N_1514,N_1409,N_1465);
and U1515 (N_1515,N_1206,N_1313);
xnor U1516 (N_1516,N_1492,N_1189);
nand U1517 (N_1517,N_1279,N_1251);
or U1518 (N_1518,N_1167,N_1432);
nand U1519 (N_1519,N_1450,N_1336);
and U1520 (N_1520,N_1400,N_1143);
or U1521 (N_1521,N_1112,N_1354);
nand U1522 (N_1522,N_1214,N_1339);
or U1523 (N_1523,N_1042,N_1494);
xor U1524 (N_1524,N_1046,N_1464);
nand U1525 (N_1525,N_1105,N_1496);
xor U1526 (N_1526,N_1406,N_1425);
nor U1527 (N_1527,N_1122,N_1358);
or U1528 (N_1528,N_1002,N_1490);
nor U1529 (N_1529,N_1493,N_1281);
nor U1530 (N_1530,N_1050,N_1376);
nand U1531 (N_1531,N_1237,N_1357);
and U1532 (N_1532,N_1225,N_1327);
nand U1533 (N_1533,N_1412,N_1467);
nor U1534 (N_1534,N_1325,N_1182);
or U1535 (N_1535,N_1260,N_1321);
or U1536 (N_1536,N_1482,N_1128);
nand U1537 (N_1537,N_1278,N_1476);
nor U1538 (N_1538,N_1394,N_1159);
xnor U1539 (N_1539,N_1458,N_1001);
and U1540 (N_1540,N_1401,N_1334);
xnor U1541 (N_1541,N_1269,N_1183);
nor U1542 (N_1542,N_1006,N_1030);
nand U1543 (N_1543,N_1391,N_1066);
or U1544 (N_1544,N_1135,N_1204);
xor U1545 (N_1545,N_1483,N_1031);
or U1546 (N_1546,N_1443,N_1198);
nor U1547 (N_1547,N_1351,N_1098);
nor U1548 (N_1548,N_1486,N_1452);
or U1549 (N_1549,N_1228,N_1314);
or U1550 (N_1550,N_1041,N_1057);
nand U1551 (N_1551,N_1287,N_1372);
and U1552 (N_1552,N_1404,N_1234);
or U1553 (N_1553,N_1180,N_1129);
xor U1554 (N_1554,N_1052,N_1329);
or U1555 (N_1555,N_1253,N_1389);
or U1556 (N_1556,N_1344,N_1120);
xnor U1557 (N_1557,N_1403,N_1119);
xor U1558 (N_1558,N_1428,N_1078);
or U1559 (N_1559,N_1282,N_1266);
nand U1560 (N_1560,N_1020,N_1353);
or U1561 (N_1561,N_1392,N_1323);
nand U1562 (N_1562,N_1166,N_1016);
nor U1563 (N_1563,N_1059,N_1398);
nor U1564 (N_1564,N_1164,N_1337);
nor U1565 (N_1565,N_1283,N_1322);
and U1566 (N_1566,N_1144,N_1142);
nand U1567 (N_1567,N_1362,N_1116);
xor U1568 (N_1568,N_1029,N_1489);
xor U1569 (N_1569,N_1331,N_1013);
nand U1570 (N_1570,N_1154,N_1036);
and U1571 (N_1571,N_1285,N_1436);
nor U1572 (N_1572,N_1365,N_1259);
nor U1573 (N_1573,N_1262,N_1025);
nor U1574 (N_1574,N_1093,N_1067);
or U1575 (N_1575,N_1149,N_1009);
and U1576 (N_1576,N_1466,N_1012);
or U1577 (N_1577,N_1430,N_1484);
and U1578 (N_1578,N_1084,N_1457);
and U1579 (N_1579,N_1364,N_1440);
nor U1580 (N_1580,N_1184,N_1221);
or U1581 (N_1581,N_1305,N_1360);
or U1582 (N_1582,N_1276,N_1309);
nand U1583 (N_1583,N_1200,N_1333);
nor U1584 (N_1584,N_1223,N_1127);
xnor U1585 (N_1585,N_1296,N_1190);
xnor U1586 (N_1586,N_1491,N_1199);
or U1587 (N_1587,N_1039,N_1289);
nand U1588 (N_1588,N_1277,N_1011);
nor U1589 (N_1589,N_1181,N_1367);
and U1590 (N_1590,N_1397,N_1242);
nor U1591 (N_1591,N_1021,N_1416);
xnor U1592 (N_1592,N_1312,N_1429);
xor U1593 (N_1593,N_1090,N_1076);
nand U1594 (N_1594,N_1462,N_1408);
and U1595 (N_1595,N_1447,N_1338);
and U1596 (N_1596,N_1384,N_1170);
and U1597 (N_1597,N_1442,N_1003);
nand U1598 (N_1598,N_1194,N_1040);
or U1599 (N_1599,N_1475,N_1455);
nor U1600 (N_1600,N_1133,N_1405);
or U1601 (N_1601,N_1160,N_1075);
or U1602 (N_1602,N_1158,N_1445);
nand U1603 (N_1603,N_1356,N_1091);
nor U1604 (N_1604,N_1058,N_1137);
and U1605 (N_1605,N_1410,N_1382);
xnor U1606 (N_1606,N_1377,N_1390);
nor U1607 (N_1607,N_1169,N_1026);
nand U1608 (N_1608,N_1318,N_1115);
nand U1609 (N_1609,N_1023,N_1472);
nor U1610 (N_1610,N_1271,N_1261);
nand U1611 (N_1611,N_1108,N_1136);
and U1612 (N_1612,N_1273,N_1043);
nor U1613 (N_1613,N_1498,N_1371);
nand U1614 (N_1614,N_1444,N_1488);
nor U1615 (N_1615,N_1479,N_1343);
xor U1616 (N_1616,N_1086,N_1307);
xnor U1617 (N_1617,N_1311,N_1195);
and U1618 (N_1618,N_1487,N_1165);
and U1619 (N_1619,N_1069,N_1256);
xnor U1620 (N_1620,N_1097,N_1288);
or U1621 (N_1621,N_1132,N_1064);
or U1622 (N_1622,N_1446,N_1080);
xor U1623 (N_1623,N_1035,N_1438);
or U1624 (N_1624,N_1082,N_1051);
xnor U1625 (N_1625,N_1216,N_1383);
xor U1626 (N_1626,N_1032,N_1375);
nor U1627 (N_1627,N_1434,N_1471);
nor U1628 (N_1628,N_1469,N_1196);
xnor U1629 (N_1629,N_1068,N_1272);
xor U1630 (N_1630,N_1074,N_1257);
nand U1631 (N_1631,N_1417,N_1176);
and U1632 (N_1632,N_1304,N_1268);
nor U1633 (N_1633,N_1060,N_1014);
xnor U1634 (N_1634,N_1109,N_1419);
nor U1635 (N_1635,N_1366,N_1219);
and U1636 (N_1636,N_1220,N_1478);
or U1637 (N_1637,N_1099,N_1056);
xor U1638 (N_1638,N_1348,N_1102);
and U1639 (N_1639,N_1328,N_1463);
nor U1640 (N_1640,N_1033,N_1399);
nor U1641 (N_1641,N_1470,N_1437);
nand U1642 (N_1642,N_1424,N_1270);
xnor U1643 (N_1643,N_1236,N_1103);
or U1644 (N_1644,N_1381,N_1081);
nand U1645 (N_1645,N_1146,N_1326);
nor U1646 (N_1646,N_1034,N_1320);
nor U1647 (N_1647,N_1015,N_1079);
and U1648 (N_1648,N_1459,N_1448);
and U1649 (N_1649,N_1227,N_1053);
and U1650 (N_1650,N_1495,N_1395);
nor U1651 (N_1651,N_1168,N_1100);
and U1652 (N_1652,N_1298,N_1427);
xnor U1653 (N_1653,N_1301,N_1264);
nand U1654 (N_1654,N_1054,N_1473);
nor U1655 (N_1655,N_1113,N_1238);
and U1656 (N_1656,N_1187,N_1265);
or U1657 (N_1657,N_1191,N_1477);
nor U1658 (N_1658,N_1232,N_1085);
or U1659 (N_1659,N_1017,N_1453);
xor U1660 (N_1660,N_1481,N_1130);
nand U1661 (N_1661,N_1454,N_1374);
nor U1662 (N_1662,N_1267,N_1396);
nor U1663 (N_1663,N_1352,N_1071);
and U1664 (N_1664,N_1241,N_1308);
or U1665 (N_1665,N_1300,N_1156);
xor U1666 (N_1666,N_1193,N_1197);
nand U1667 (N_1667,N_1456,N_1330);
and U1668 (N_1668,N_1140,N_1286);
or U1669 (N_1669,N_1000,N_1208);
and U1670 (N_1670,N_1292,N_1407);
nor U1671 (N_1671,N_1295,N_1072);
or U1672 (N_1672,N_1157,N_1361);
and U1673 (N_1673,N_1083,N_1061);
and U1674 (N_1674,N_1290,N_1317);
or U1675 (N_1675,N_1062,N_1185);
xor U1676 (N_1676,N_1028,N_1186);
or U1677 (N_1677,N_1215,N_1038);
and U1678 (N_1678,N_1096,N_1117);
xnor U1679 (N_1679,N_1415,N_1255);
xnor U1680 (N_1680,N_1153,N_1151);
xor U1681 (N_1681,N_1045,N_1008);
xor U1682 (N_1682,N_1480,N_1340);
or U1683 (N_1683,N_1303,N_1055);
xor U1684 (N_1684,N_1150,N_1049);
or U1685 (N_1685,N_1209,N_1379);
xnor U1686 (N_1686,N_1310,N_1299);
nand U1687 (N_1687,N_1134,N_1118);
nand U1688 (N_1688,N_1433,N_1104);
nand U1689 (N_1689,N_1422,N_1244);
and U1690 (N_1690,N_1205,N_1087);
and U1691 (N_1691,N_1175,N_1155);
nand U1692 (N_1692,N_1018,N_1423);
xor U1693 (N_1693,N_1152,N_1044);
xor U1694 (N_1694,N_1431,N_1111);
xnor U1695 (N_1695,N_1145,N_1421);
and U1696 (N_1696,N_1294,N_1073);
nand U1697 (N_1697,N_1126,N_1172);
and U1698 (N_1698,N_1094,N_1393);
xnor U1699 (N_1699,N_1386,N_1022);
xnor U1700 (N_1700,N_1345,N_1174);
xnor U1701 (N_1701,N_1178,N_1231);
xnor U1702 (N_1702,N_1162,N_1233);
nor U1703 (N_1703,N_1027,N_1217);
xnor U1704 (N_1704,N_1418,N_1131);
or U1705 (N_1705,N_1324,N_1385);
nand U1706 (N_1706,N_1188,N_1211);
or U1707 (N_1707,N_1005,N_1280);
and U1708 (N_1708,N_1248,N_1213);
xor U1709 (N_1709,N_1359,N_1293);
nand U1710 (N_1710,N_1092,N_1319);
nor U1711 (N_1711,N_1089,N_1125);
nand U1712 (N_1712,N_1380,N_1024);
xnor U1713 (N_1713,N_1441,N_1499);
nand U1714 (N_1714,N_1258,N_1284);
nor U1715 (N_1715,N_1250,N_1497);
and U1716 (N_1716,N_1451,N_1349);
and U1717 (N_1717,N_1246,N_1332);
nand U1718 (N_1718,N_1342,N_1048);
xnor U1719 (N_1719,N_1435,N_1010);
nand U1720 (N_1720,N_1235,N_1207);
and U1721 (N_1721,N_1110,N_1402);
nand U1722 (N_1722,N_1218,N_1004);
nand U1723 (N_1723,N_1230,N_1274);
nand U1724 (N_1724,N_1088,N_1247);
and U1725 (N_1725,N_1388,N_1226);
nand U1726 (N_1726,N_1368,N_1346);
xnor U1727 (N_1727,N_1138,N_1147);
nor U1728 (N_1728,N_1179,N_1414);
and U1729 (N_1729,N_1363,N_1252);
or U1730 (N_1730,N_1341,N_1460);
nand U1731 (N_1731,N_1161,N_1370);
and U1732 (N_1732,N_1413,N_1378);
and U1733 (N_1733,N_1302,N_1245);
nor U1734 (N_1734,N_1291,N_1373);
xor U1735 (N_1735,N_1177,N_1107);
nand U1736 (N_1736,N_1019,N_1070);
nand U1737 (N_1737,N_1203,N_1163);
and U1738 (N_1738,N_1420,N_1369);
nand U1739 (N_1739,N_1449,N_1106);
nor U1740 (N_1740,N_1355,N_1141);
nor U1741 (N_1741,N_1210,N_1243);
nand U1742 (N_1742,N_1148,N_1224);
nand U1743 (N_1743,N_1222,N_1123);
nor U1744 (N_1744,N_1411,N_1077);
nor U1745 (N_1745,N_1426,N_1335);
xor U1746 (N_1746,N_1350,N_1101);
and U1747 (N_1747,N_1007,N_1461);
xor U1748 (N_1748,N_1297,N_1249);
nand U1749 (N_1749,N_1263,N_1485);
and U1750 (N_1750,N_1303,N_1457);
and U1751 (N_1751,N_1421,N_1110);
and U1752 (N_1752,N_1269,N_1412);
and U1753 (N_1753,N_1413,N_1320);
xor U1754 (N_1754,N_1282,N_1345);
xnor U1755 (N_1755,N_1484,N_1006);
xnor U1756 (N_1756,N_1192,N_1012);
and U1757 (N_1757,N_1493,N_1319);
nand U1758 (N_1758,N_1085,N_1279);
and U1759 (N_1759,N_1294,N_1145);
nor U1760 (N_1760,N_1194,N_1264);
xnor U1761 (N_1761,N_1482,N_1087);
nor U1762 (N_1762,N_1497,N_1054);
nand U1763 (N_1763,N_1226,N_1380);
xnor U1764 (N_1764,N_1131,N_1250);
or U1765 (N_1765,N_1267,N_1206);
and U1766 (N_1766,N_1410,N_1220);
or U1767 (N_1767,N_1269,N_1249);
xor U1768 (N_1768,N_1237,N_1037);
nand U1769 (N_1769,N_1025,N_1180);
or U1770 (N_1770,N_1475,N_1188);
xnor U1771 (N_1771,N_1094,N_1485);
nor U1772 (N_1772,N_1099,N_1406);
nor U1773 (N_1773,N_1473,N_1301);
and U1774 (N_1774,N_1029,N_1258);
xnor U1775 (N_1775,N_1333,N_1443);
xor U1776 (N_1776,N_1064,N_1051);
and U1777 (N_1777,N_1352,N_1060);
xnor U1778 (N_1778,N_1006,N_1016);
or U1779 (N_1779,N_1218,N_1435);
nand U1780 (N_1780,N_1103,N_1109);
xnor U1781 (N_1781,N_1216,N_1172);
or U1782 (N_1782,N_1462,N_1197);
or U1783 (N_1783,N_1193,N_1257);
xor U1784 (N_1784,N_1046,N_1057);
nor U1785 (N_1785,N_1313,N_1175);
and U1786 (N_1786,N_1394,N_1020);
nor U1787 (N_1787,N_1431,N_1316);
nand U1788 (N_1788,N_1042,N_1420);
nand U1789 (N_1789,N_1222,N_1418);
xnor U1790 (N_1790,N_1090,N_1238);
nor U1791 (N_1791,N_1170,N_1032);
nor U1792 (N_1792,N_1167,N_1003);
nor U1793 (N_1793,N_1082,N_1081);
nand U1794 (N_1794,N_1220,N_1317);
nand U1795 (N_1795,N_1122,N_1056);
xor U1796 (N_1796,N_1390,N_1181);
or U1797 (N_1797,N_1057,N_1303);
nand U1798 (N_1798,N_1152,N_1248);
or U1799 (N_1799,N_1184,N_1116);
and U1800 (N_1800,N_1156,N_1014);
nor U1801 (N_1801,N_1277,N_1371);
xnor U1802 (N_1802,N_1342,N_1192);
nand U1803 (N_1803,N_1436,N_1197);
nand U1804 (N_1804,N_1247,N_1006);
xnor U1805 (N_1805,N_1363,N_1128);
or U1806 (N_1806,N_1025,N_1466);
xnor U1807 (N_1807,N_1387,N_1068);
or U1808 (N_1808,N_1479,N_1182);
xor U1809 (N_1809,N_1437,N_1375);
nor U1810 (N_1810,N_1019,N_1494);
nor U1811 (N_1811,N_1176,N_1394);
nor U1812 (N_1812,N_1390,N_1476);
nand U1813 (N_1813,N_1043,N_1433);
xor U1814 (N_1814,N_1238,N_1064);
or U1815 (N_1815,N_1406,N_1024);
and U1816 (N_1816,N_1285,N_1094);
xnor U1817 (N_1817,N_1435,N_1284);
and U1818 (N_1818,N_1488,N_1258);
or U1819 (N_1819,N_1441,N_1089);
nor U1820 (N_1820,N_1431,N_1193);
nor U1821 (N_1821,N_1472,N_1273);
or U1822 (N_1822,N_1097,N_1400);
xor U1823 (N_1823,N_1062,N_1453);
nand U1824 (N_1824,N_1274,N_1496);
and U1825 (N_1825,N_1462,N_1379);
and U1826 (N_1826,N_1428,N_1044);
or U1827 (N_1827,N_1331,N_1214);
nand U1828 (N_1828,N_1242,N_1393);
nor U1829 (N_1829,N_1353,N_1289);
and U1830 (N_1830,N_1356,N_1406);
xnor U1831 (N_1831,N_1068,N_1358);
and U1832 (N_1832,N_1404,N_1274);
or U1833 (N_1833,N_1407,N_1254);
xor U1834 (N_1834,N_1135,N_1256);
and U1835 (N_1835,N_1235,N_1404);
or U1836 (N_1836,N_1318,N_1468);
xor U1837 (N_1837,N_1401,N_1094);
xnor U1838 (N_1838,N_1401,N_1039);
nand U1839 (N_1839,N_1020,N_1410);
nor U1840 (N_1840,N_1099,N_1319);
nand U1841 (N_1841,N_1231,N_1445);
nand U1842 (N_1842,N_1064,N_1074);
and U1843 (N_1843,N_1023,N_1499);
xor U1844 (N_1844,N_1001,N_1492);
nor U1845 (N_1845,N_1483,N_1102);
and U1846 (N_1846,N_1087,N_1192);
and U1847 (N_1847,N_1122,N_1439);
nand U1848 (N_1848,N_1156,N_1414);
and U1849 (N_1849,N_1231,N_1080);
or U1850 (N_1850,N_1002,N_1183);
or U1851 (N_1851,N_1055,N_1233);
nand U1852 (N_1852,N_1231,N_1240);
nor U1853 (N_1853,N_1402,N_1089);
xor U1854 (N_1854,N_1184,N_1196);
nor U1855 (N_1855,N_1219,N_1426);
nand U1856 (N_1856,N_1305,N_1317);
and U1857 (N_1857,N_1076,N_1002);
and U1858 (N_1858,N_1207,N_1495);
nor U1859 (N_1859,N_1034,N_1167);
or U1860 (N_1860,N_1178,N_1471);
and U1861 (N_1861,N_1122,N_1029);
xnor U1862 (N_1862,N_1299,N_1230);
xor U1863 (N_1863,N_1279,N_1185);
xnor U1864 (N_1864,N_1323,N_1442);
or U1865 (N_1865,N_1074,N_1165);
nand U1866 (N_1866,N_1143,N_1330);
or U1867 (N_1867,N_1215,N_1432);
xor U1868 (N_1868,N_1224,N_1075);
nor U1869 (N_1869,N_1157,N_1167);
and U1870 (N_1870,N_1124,N_1284);
xor U1871 (N_1871,N_1241,N_1265);
xor U1872 (N_1872,N_1230,N_1448);
or U1873 (N_1873,N_1087,N_1093);
nor U1874 (N_1874,N_1148,N_1472);
nor U1875 (N_1875,N_1407,N_1125);
nor U1876 (N_1876,N_1256,N_1058);
nor U1877 (N_1877,N_1273,N_1269);
or U1878 (N_1878,N_1368,N_1201);
or U1879 (N_1879,N_1202,N_1217);
or U1880 (N_1880,N_1099,N_1384);
nor U1881 (N_1881,N_1079,N_1328);
nor U1882 (N_1882,N_1248,N_1471);
xor U1883 (N_1883,N_1300,N_1260);
or U1884 (N_1884,N_1482,N_1457);
and U1885 (N_1885,N_1106,N_1045);
and U1886 (N_1886,N_1430,N_1443);
xor U1887 (N_1887,N_1386,N_1174);
or U1888 (N_1888,N_1172,N_1102);
xor U1889 (N_1889,N_1038,N_1256);
and U1890 (N_1890,N_1305,N_1424);
and U1891 (N_1891,N_1480,N_1230);
nand U1892 (N_1892,N_1181,N_1199);
and U1893 (N_1893,N_1367,N_1001);
nor U1894 (N_1894,N_1117,N_1228);
and U1895 (N_1895,N_1455,N_1429);
nor U1896 (N_1896,N_1314,N_1276);
or U1897 (N_1897,N_1005,N_1234);
nand U1898 (N_1898,N_1332,N_1403);
or U1899 (N_1899,N_1420,N_1170);
nor U1900 (N_1900,N_1075,N_1191);
and U1901 (N_1901,N_1191,N_1171);
nand U1902 (N_1902,N_1030,N_1240);
nor U1903 (N_1903,N_1446,N_1059);
or U1904 (N_1904,N_1396,N_1306);
nor U1905 (N_1905,N_1028,N_1385);
and U1906 (N_1906,N_1012,N_1334);
xnor U1907 (N_1907,N_1256,N_1200);
xor U1908 (N_1908,N_1490,N_1324);
nor U1909 (N_1909,N_1019,N_1052);
and U1910 (N_1910,N_1152,N_1449);
or U1911 (N_1911,N_1227,N_1284);
nor U1912 (N_1912,N_1375,N_1373);
nor U1913 (N_1913,N_1243,N_1177);
or U1914 (N_1914,N_1297,N_1124);
nand U1915 (N_1915,N_1419,N_1374);
xor U1916 (N_1916,N_1361,N_1072);
nand U1917 (N_1917,N_1054,N_1348);
nand U1918 (N_1918,N_1256,N_1025);
or U1919 (N_1919,N_1120,N_1339);
nand U1920 (N_1920,N_1488,N_1000);
nand U1921 (N_1921,N_1375,N_1207);
nor U1922 (N_1922,N_1122,N_1232);
nor U1923 (N_1923,N_1195,N_1301);
and U1924 (N_1924,N_1089,N_1477);
or U1925 (N_1925,N_1104,N_1430);
xnor U1926 (N_1926,N_1376,N_1485);
or U1927 (N_1927,N_1019,N_1129);
nor U1928 (N_1928,N_1267,N_1363);
xor U1929 (N_1929,N_1029,N_1300);
nor U1930 (N_1930,N_1431,N_1058);
xor U1931 (N_1931,N_1306,N_1237);
and U1932 (N_1932,N_1445,N_1356);
and U1933 (N_1933,N_1430,N_1156);
or U1934 (N_1934,N_1356,N_1177);
or U1935 (N_1935,N_1019,N_1365);
nand U1936 (N_1936,N_1481,N_1300);
or U1937 (N_1937,N_1310,N_1335);
and U1938 (N_1938,N_1360,N_1317);
nor U1939 (N_1939,N_1230,N_1228);
or U1940 (N_1940,N_1207,N_1310);
nand U1941 (N_1941,N_1456,N_1061);
nor U1942 (N_1942,N_1474,N_1404);
nand U1943 (N_1943,N_1357,N_1311);
nand U1944 (N_1944,N_1478,N_1329);
xnor U1945 (N_1945,N_1040,N_1089);
nand U1946 (N_1946,N_1059,N_1378);
xnor U1947 (N_1947,N_1015,N_1393);
nand U1948 (N_1948,N_1277,N_1194);
xnor U1949 (N_1949,N_1458,N_1039);
nor U1950 (N_1950,N_1308,N_1025);
or U1951 (N_1951,N_1134,N_1231);
nand U1952 (N_1952,N_1287,N_1037);
nor U1953 (N_1953,N_1251,N_1027);
and U1954 (N_1954,N_1243,N_1145);
xor U1955 (N_1955,N_1127,N_1240);
or U1956 (N_1956,N_1279,N_1019);
xnor U1957 (N_1957,N_1401,N_1329);
and U1958 (N_1958,N_1176,N_1145);
nor U1959 (N_1959,N_1216,N_1106);
nand U1960 (N_1960,N_1006,N_1042);
or U1961 (N_1961,N_1263,N_1461);
nor U1962 (N_1962,N_1138,N_1201);
nand U1963 (N_1963,N_1367,N_1013);
nand U1964 (N_1964,N_1118,N_1244);
nand U1965 (N_1965,N_1092,N_1165);
and U1966 (N_1966,N_1167,N_1146);
xnor U1967 (N_1967,N_1427,N_1113);
nand U1968 (N_1968,N_1263,N_1446);
xnor U1969 (N_1969,N_1443,N_1376);
nand U1970 (N_1970,N_1392,N_1104);
or U1971 (N_1971,N_1365,N_1467);
or U1972 (N_1972,N_1130,N_1051);
nor U1973 (N_1973,N_1191,N_1131);
nand U1974 (N_1974,N_1245,N_1053);
xnor U1975 (N_1975,N_1494,N_1483);
or U1976 (N_1976,N_1187,N_1232);
xor U1977 (N_1977,N_1032,N_1069);
or U1978 (N_1978,N_1499,N_1203);
nand U1979 (N_1979,N_1105,N_1384);
and U1980 (N_1980,N_1404,N_1392);
nor U1981 (N_1981,N_1032,N_1001);
nand U1982 (N_1982,N_1192,N_1241);
nand U1983 (N_1983,N_1243,N_1294);
nand U1984 (N_1984,N_1191,N_1430);
nand U1985 (N_1985,N_1043,N_1229);
xor U1986 (N_1986,N_1299,N_1128);
xnor U1987 (N_1987,N_1197,N_1457);
nor U1988 (N_1988,N_1200,N_1304);
or U1989 (N_1989,N_1307,N_1167);
nor U1990 (N_1990,N_1068,N_1215);
nor U1991 (N_1991,N_1131,N_1287);
xnor U1992 (N_1992,N_1479,N_1413);
nor U1993 (N_1993,N_1471,N_1127);
or U1994 (N_1994,N_1120,N_1119);
and U1995 (N_1995,N_1480,N_1319);
nor U1996 (N_1996,N_1220,N_1088);
xnor U1997 (N_1997,N_1431,N_1209);
nand U1998 (N_1998,N_1444,N_1387);
nand U1999 (N_1999,N_1452,N_1331);
xnor U2000 (N_2000,N_1582,N_1820);
xnor U2001 (N_2001,N_1860,N_1887);
nor U2002 (N_2002,N_1973,N_1566);
nor U2003 (N_2003,N_1950,N_1971);
xor U2004 (N_2004,N_1801,N_1586);
nor U2005 (N_2005,N_1906,N_1931);
nor U2006 (N_2006,N_1507,N_1946);
xnor U2007 (N_2007,N_1880,N_1808);
or U2008 (N_2008,N_1972,N_1641);
nand U2009 (N_2009,N_1854,N_1825);
xor U2010 (N_2010,N_1750,N_1509);
xnor U2011 (N_2011,N_1814,N_1824);
or U2012 (N_2012,N_1954,N_1584);
nand U2013 (N_2013,N_1719,N_1995);
nor U2014 (N_2014,N_1903,N_1714);
or U2015 (N_2015,N_1742,N_1567);
or U2016 (N_2016,N_1646,N_1920);
or U2017 (N_2017,N_1941,N_1798);
and U2018 (N_2018,N_1796,N_1899);
and U2019 (N_2019,N_1767,N_1760);
nor U2020 (N_2020,N_1660,N_1749);
and U2021 (N_2021,N_1657,N_1709);
or U2022 (N_2022,N_1610,N_1565);
nor U2023 (N_2023,N_1807,N_1698);
nor U2024 (N_2024,N_1753,N_1501);
xnor U2025 (N_2025,N_1847,N_1851);
and U2026 (N_2026,N_1800,N_1844);
or U2027 (N_2027,N_1664,N_1790);
or U2028 (N_2028,N_1916,N_1774);
nor U2029 (N_2029,N_1997,N_1724);
and U2030 (N_2030,N_1683,N_1883);
xnor U2031 (N_2031,N_1738,N_1831);
and U2032 (N_2032,N_1817,N_1710);
nand U2033 (N_2033,N_1624,N_1529);
and U2034 (N_2034,N_1703,N_1687);
nand U2035 (N_2035,N_1615,N_1651);
or U2036 (N_2036,N_1856,N_1722);
xnor U2037 (N_2037,N_1556,N_1969);
and U2038 (N_2038,N_1948,N_1729);
or U2039 (N_2039,N_1794,N_1721);
xor U2040 (N_2040,N_1616,N_1546);
xor U2041 (N_2041,N_1563,N_1806);
nor U2042 (N_2042,N_1984,N_1761);
and U2043 (N_2043,N_1676,N_1868);
xor U2044 (N_2044,N_1743,N_1803);
and U2045 (N_2045,N_1999,N_1513);
and U2046 (N_2046,N_1974,N_1754);
xnor U2047 (N_2047,N_1508,N_1909);
or U2048 (N_2048,N_1980,N_1520);
and U2049 (N_2049,N_1572,N_1765);
or U2050 (N_2050,N_1895,N_1871);
and U2051 (N_2051,N_1611,N_1737);
and U2052 (N_2052,N_1758,N_1589);
and U2053 (N_2053,N_1823,N_1991);
or U2054 (N_2054,N_1500,N_1921);
nor U2055 (N_2055,N_1930,N_1989);
or U2056 (N_2056,N_1894,N_1560);
xnor U2057 (N_2057,N_1647,N_1911);
or U2058 (N_2058,N_1601,N_1620);
nand U2059 (N_2059,N_1769,N_1922);
nand U2060 (N_2060,N_1875,N_1975);
nor U2061 (N_2061,N_1658,N_1994);
xnor U2062 (N_2062,N_1608,N_1732);
nand U2063 (N_2063,N_1604,N_1955);
nor U2064 (N_2064,N_1650,N_1713);
or U2065 (N_2065,N_1862,N_1544);
and U2066 (N_2066,N_1970,N_1515);
or U2067 (N_2067,N_1639,N_1898);
and U2068 (N_2068,N_1943,N_1813);
or U2069 (N_2069,N_1848,N_1835);
or U2070 (N_2070,N_1771,N_1675);
nor U2071 (N_2071,N_1587,N_1693);
and U2072 (N_2072,N_1874,N_1688);
or U2073 (N_2073,N_1841,N_1932);
nand U2074 (N_2074,N_1910,N_1778);
or U2075 (N_2075,N_1524,N_1740);
nor U2076 (N_2076,N_1992,N_1878);
and U2077 (N_2077,N_1528,N_1779);
or U2078 (N_2078,N_1625,N_1592);
or U2079 (N_2079,N_1925,N_1745);
xnor U2080 (N_2080,N_1967,N_1671);
or U2081 (N_2081,N_1746,N_1668);
or U2082 (N_2082,N_1547,N_1701);
nand U2083 (N_2083,N_1907,N_1963);
or U2084 (N_2084,N_1747,N_1846);
nor U2085 (N_2085,N_1821,N_1559);
and U2086 (N_2086,N_1818,N_1748);
xnor U2087 (N_2087,N_1670,N_1892);
or U2088 (N_2088,N_1988,N_1542);
and U2089 (N_2089,N_1935,N_1540);
or U2090 (N_2090,N_1797,N_1780);
or U2091 (N_2091,N_1518,N_1558);
or U2092 (N_2092,N_1786,N_1934);
nor U2093 (N_2093,N_1811,N_1885);
or U2094 (N_2094,N_1622,N_1833);
or U2095 (N_2095,N_1543,N_1642);
or U2096 (N_2096,N_1663,N_1727);
and U2097 (N_2097,N_1531,N_1886);
or U2098 (N_2098,N_1768,N_1978);
or U2099 (N_2099,N_1926,N_1652);
xnor U2100 (N_2100,N_1773,N_1990);
and U2101 (N_2101,N_1876,N_1557);
and U2102 (N_2102,N_1606,N_1590);
and U2103 (N_2103,N_1828,N_1968);
or U2104 (N_2104,N_1549,N_1867);
nand U2105 (N_2105,N_1504,N_1511);
or U2106 (N_2106,N_1653,N_1661);
nor U2107 (N_2107,N_1982,N_1550);
or U2108 (N_2108,N_1901,N_1623);
nand U2109 (N_2109,N_1599,N_1686);
or U2110 (N_2110,N_1891,N_1865);
or U2111 (N_2111,N_1929,N_1609);
or U2112 (N_2112,N_1965,N_1918);
xor U2113 (N_2113,N_1619,N_1637);
xnor U2114 (N_2114,N_1585,N_1957);
nand U2115 (N_2115,N_1949,N_1977);
and U2116 (N_2116,N_1964,N_1861);
nor U2117 (N_2117,N_1857,N_1672);
or U2118 (N_2118,N_1993,N_1777);
and U2119 (N_2119,N_1681,N_1945);
xor U2120 (N_2120,N_1849,N_1845);
xor U2121 (N_2121,N_1612,N_1712);
or U2122 (N_2122,N_1602,N_1863);
nor U2123 (N_2123,N_1942,N_1522);
nand U2124 (N_2124,N_1532,N_1776);
or U2125 (N_2125,N_1897,N_1579);
or U2126 (N_2126,N_1725,N_1789);
and U2127 (N_2127,N_1649,N_1689);
or U2128 (N_2128,N_1766,N_1541);
xnor U2129 (N_2129,N_1512,N_1952);
xnor U2130 (N_2130,N_1503,N_1837);
nand U2131 (N_2131,N_1530,N_1506);
or U2132 (N_2132,N_1762,N_1928);
nor U2133 (N_2133,N_1537,N_1947);
nor U2134 (N_2134,N_1804,N_1636);
xnor U2135 (N_2135,N_1576,N_1545);
xor U2136 (N_2136,N_1730,N_1525);
and U2137 (N_2137,N_1877,N_1678);
nor U2138 (N_2138,N_1632,N_1843);
or U2139 (N_2139,N_1691,N_1872);
nand U2140 (N_2140,N_1527,N_1638);
xor U2141 (N_2141,N_1832,N_1613);
nor U2142 (N_2142,N_1764,N_1827);
nand U2143 (N_2143,N_1697,N_1781);
xor U2144 (N_2144,N_1505,N_1870);
nand U2145 (N_2145,N_1621,N_1961);
nand U2146 (N_2146,N_1659,N_1917);
and U2147 (N_2147,N_1979,N_1564);
nand U2148 (N_2148,N_1553,N_1890);
and U2149 (N_2149,N_1521,N_1893);
and U2150 (N_2150,N_1834,N_1793);
xnor U2151 (N_2151,N_1884,N_1702);
nor U2152 (N_2152,N_1900,N_1607);
and U2153 (N_2153,N_1645,N_1873);
or U2154 (N_2154,N_1662,N_1554);
nand U2155 (N_2155,N_1694,N_1783);
nor U2156 (N_2156,N_1933,N_1919);
nand U2157 (N_2157,N_1596,N_1573);
nand U2158 (N_2158,N_1631,N_1580);
nor U2159 (N_2159,N_1575,N_1655);
or U2160 (N_2160,N_1514,N_1718);
xnor U2161 (N_2161,N_1864,N_1998);
nor U2162 (N_2162,N_1588,N_1684);
xnor U2163 (N_2163,N_1838,N_1535);
nor U2164 (N_2164,N_1706,N_1654);
nor U2165 (N_2165,N_1815,N_1731);
nor U2166 (N_2166,N_1640,N_1716);
nand U2167 (N_2167,N_1809,N_1889);
xor U2168 (N_2168,N_1555,N_1836);
xnor U2169 (N_2169,N_1756,N_1959);
nor U2170 (N_2170,N_1577,N_1578);
nor U2171 (N_2171,N_1600,N_1858);
nand U2172 (N_2172,N_1533,N_1744);
and U2173 (N_2173,N_1648,N_1669);
and U2174 (N_2174,N_1759,N_1630);
and U2175 (N_2175,N_1635,N_1679);
and U2176 (N_2176,N_1723,N_1830);
nor U2177 (N_2177,N_1690,N_1734);
and U2178 (N_2178,N_1539,N_1569);
and U2179 (N_2179,N_1966,N_1674);
and U2180 (N_2180,N_1937,N_1666);
xnor U2181 (N_2181,N_1939,N_1643);
nand U2182 (N_2182,N_1728,N_1908);
or U2183 (N_2183,N_1822,N_1960);
or U2184 (N_2184,N_1976,N_1736);
or U2185 (N_2185,N_1685,N_1629);
or U2186 (N_2186,N_1574,N_1855);
nor U2187 (N_2187,N_1699,N_1850);
and U2188 (N_2188,N_1904,N_1516);
nand U2189 (N_2189,N_1819,N_1958);
xor U2190 (N_2190,N_1951,N_1953);
or U2191 (N_2191,N_1881,N_1791);
xor U2192 (N_2192,N_1677,N_1534);
nand U2193 (N_2193,N_1805,N_1705);
xnor U2194 (N_2194,N_1597,N_1812);
nor U2195 (N_2195,N_1626,N_1502);
xor U2196 (N_2196,N_1538,N_1715);
and U2197 (N_2197,N_1614,N_1869);
or U2198 (N_2198,N_1924,N_1548);
nand U2199 (N_2199,N_1888,N_1914);
or U2200 (N_2200,N_1755,N_1618);
and U2201 (N_2201,N_1519,N_1810);
nand U2202 (N_2202,N_1962,N_1839);
xor U2203 (N_2203,N_1644,N_1717);
nor U2204 (N_2204,N_1981,N_1634);
nand U2205 (N_2205,N_1936,N_1562);
or U2206 (N_2206,N_1859,N_1826);
nand U2207 (N_2207,N_1986,N_1726);
or U2208 (N_2208,N_1913,N_1656);
xnor U2209 (N_2209,N_1680,N_1673);
xnor U2210 (N_2210,N_1816,N_1763);
xnor U2211 (N_2211,N_1568,N_1739);
and U2212 (N_2212,N_1733,N_1741);
and U2213 (N_2213,N_1628,N_1517);
nand U2214 (N_2214,N_1912,N_1605);
nand U2215 (N_2215,N_1757,N_1696);
nor U2216 (N_2216,N_1775,N_1782);
and U2217 (N_2217,N_1720,N_1523);
nand U2218 (N_2218,N_1840,N_1787);
and U2219 (N_2219,N_1799,N_1591);
nand U2220 (N_2220,N_1594,N_1711);
nand U2221 (N_2221,N_1752,N_1692);
and U2222 (N_2222,N_1552,N_1940);
nand U2223 (N_2223,N_1583,N_1956);
or U2224 (N_2224,N_1938,N_1603);
nor U2225 (N_2225,N_1536,N_1923);
or U2226 (N_2226,N_1896,N_1829);
nor U2227 (N_2227,N_1561,N_1667);
nand U2228 (N_2228,N_1751,N_1551);
nand U2229 (N_2229,N_1784,N_1983);
xor U2230 (N_2230,N_1633,N_1802);
and U2231 (N_2231,N_1571,N_1772);
or U2232 (N_2232,N_1735,N_1879);
nor U2233 (N_2233,N_1570,N_1996);
nor U2234 (N_2234,N_1598,N_1593);
nand U2235 (N_2235,N_1792,N_1581);
or U2236 (N_2236,N_1595,N_1708);
or U2237 (N_2237,N_1617,N_1788);
nand U2238 (N_2238,N_1704,N_1902);
or U2239 (N_2239,N_1627,N_1927);
or U2240 (N_2240,N_1944,N_1905);
nand U2241 (N_2241,N_1707,N_1866);
and U2242 (N_2242,N_1985,N_1852);
or U2243 (N_2243,N_1853,N_1700);
xnor U2244 (N_2244,N_1665,N_1882);
or U2245 (N_2245,N_1526,N_1795);
or U2246 (N_2246,N_1695,N_1842);
nor U2247 (N_2247,N_1915,N_1785);
and U2248 (N_2248,N_1682,N_1510);
nor U2249 (N_2249,N_1987,N_1770);
xnor U2250 (N_2250,N_1643,N_1556);
nor U2251 (N_2251,N_1932,N_1944);
xor U2252 (N_2252,N_1559,N_1810);
xor U2253 (N_2253,N_1839,N_1951);
nand U2254 (N_2254,N_1508,N_1830);
or U2255 (N_2255,N_1773,N_1914);
and U2256 (N_2256,N_1776,N_1766);
nand U2257 (N_2257,N_1933,N_1744);
xor U2258 (N_2258,N_1661,N_1978);
nand U2259 (N_2259,N_1832,N_1806);
xor U2260 (N_2260,N_1706,N_1720);
nand U2261 (N_2261,N_1608,N_1678);
and U2262 (N_2262,N_1515,N_1509);
nand U2263 (N_2263,N_1742,N_1696);
nor U2264 (N_2264,N_1778,N_1847);
and U2265 (N_2265,N_1861,N_1527);
nor U2266 (N_2266,N_1533,N_1697);
xor U2267 (N_2267,N_1857,N_1956);
nand U2268 (N_2268,N_1880,N_1760);
nor U2269 (N_2269,N_1842,N_1616);
nor U2270 (N_2270,N_1630,N_1934);
nand U2271 (N_2271,N_1992,N_1933);
xnor U2272 (N_2272,N_1798,N_1838);
nor U2273 (N_2273,N_1698,N_1729);
and U2274 (N_2274,N_1995,N_1696);
nand U2275 (N_2275,N_1823,N_1818);
or U2276 (N_2276,N_1886,N_1742);
xor U2277 (N_2277,N_1580,N_1615);
nor U2278 (N_2278,N_1593,N_1552);
xnor U2279 (N_2279,N_1616,N_1950);
nand U2280 (N_2280,N_1538,N_1852);
xnor U2281 (N_2281,N_1818,N_1939);
nand U2282 (N_2282,N_1957,N_1553);
or U2283 (N_2283,N_1624,N_1650);
xnor U2284 (N_2284,N_1865,N_1795);
xor U2285 (N_2285,N_1698,N_1976);
xor U2286 (N_2286,N_1602,N_1569);
xnor U2287 (N_2287,N_1934,N_1614);
xor U2288 (N_2288,N_1924,N_1753);
and U2289 (N_2289,N_1953,N_1803);
and U2290 (N_2290,N_1591,N_1537);
or U2291 (N_2291,N_1583,N_1953);
nor U2292 (N_2292,N_1892,N_1753);
and U2293 (N_2293,N_1970,N_1937);
nand U2294 (N_2294,N_1912,N_1617);
xor U2295 (N_2295,N_1706,N_1773);
nand U2296 (N_2296,N_1617,N_1936);
and U2297 (N_2297,N_1791,N_1520);
nor U2298 (N_2298,N_1928,N_1785);
or U2299 (N_2299,N_1533,N_1546);
and U2300 (N_2300,N_1530,N_1522);
or U2301 (N_2301,N_1749,N_1715);
and U2302 (N_2302,N_1730,N_1755);
or U2303 (N_2303,N_1660,N_1545);
nor U2304 (N_2304,N_1759,N_1918);
and U2305 (N_2305,N_1884,N_1586);
xor U2306 (N_2306,N_1723,N_1970);
or U2307 (N_2307,N_1843,N_1748);
nand U2308 (N_2308,N_1726,N_1900);
xnor U2309 (N_2309,N_1583,N_1732);
nor U2310 (N_2310,N_1554,N_1915);
or U2311 (N_2311,N_1882,N_1692);
xor U2312 (N_2312,N_1980,N_1840);
or U2313 (N_2313,N_1644,N_1576);
nor U2314 (N_2314,N_1804,N_1872);
nor U2315 (N_2315,N_1885,N_1525);
or U2316 (N_2316,N_1852,N_1979);
nor U2317 (N_2317,N_1757,N_1615);
xor U2318 (N_2318,N_1504,N_1685);
or U2319 (N_2319,N_1727,N_1924);
nor U2320 (N_2320,N_1542,N_1812);
xnor U2321 (N_2321,N_1786,N_1989);
or U2322 (N_2322,N_1958,N_1521);
nor U2323 (N_2323,N_1657,N_1510);
nor U2324 (N_2324,N_1937,N_1829);
or U2325 (N_2325,N_1934,N_1889);
or U2326 (N_2326,N_1535,N_1805);
or U2327 (N_2327,N_1967,N_1943);
nor U2328 (N_2328,N_1540,N_1790);
or U2329 (N_2329,N_1536,N_1887);
nor U2330 (N_2330,N_1705,N_1767);
or U2331 (N_2331,N_1666,N_1516);
nor U2332 (N_2332,N_1506,N_1925);
nand U2333 (N_2333,N_1827,N_1951);
or U2334 (N_2334,N_1798,N_1840);
nand U2335 (N_2335,N_1698,N_1547);
or U2336 (N_2336,N_1943,N_1946);
and U2337 (N_2337,N_1919,N_1776);
nor U2338 (N_2338,N_1757,N_1815);
xnor U2339 (N_2339,N_1702,N_1576);
xnor U2340 (N_2340,N_1591,N_1980);
nor U2341 (N_2341,N_1794,N_1878);
nand U2342 (N_2342,N_1680,N_1866);
and U2343 (N_2343,N_1667,N_1967);
or U2344 (N_2344,N_1620,N_1671);
nand U2345 (N_2345,N_1785,N_1563);
nand U2346 (N_2346,N_1592,N_1867);
nand U2347 (N_2347,N_1667,N_1621);
nor U2348 (N_2348,N_1528,N_1839);
nand U2349 (N_2349,N_1666,N_1702);
xor U2350 (N_2350,N_1915,N_1815);
and U2351 (N_2351,N_1931,N_1648);
nor U2352 (N_2352,N_1564,N_1570);
nor U2353 (N_2353,N_1641,N_1811);
or U2354 (N_2354,N_1946,N_1760);
xor U2355 (N_2355,N_1971,N_1843);
nor U2356 (N_2356,N_1815,N_1636);
or U2357 (N_2357,N_1529,N_1562);
nor U2358 (N_2358,N_1669,N_1629);
nor U2359 (N_2359,N_1638,N_1832);
xnor U2360 (N_2360,N_1725,N_1620);
nand U2361 (N_2361,N_1669,N_1521);
nand U2362 (N_2362,N_1727,N_1672);
nor U2363 (N_2363,N_1595,N_1697);
and U2364 (N_2364,N_1782,N_1545);
nand U2365 (N_2365,N_1692,N_1661);
and U2366 (N_2366,N_1701,N_1994);
or U2367 (N_2367,N_1981,N_1550);
nand U2368 (N_2368,N_1714,N_1612);
or U2369 (N_2369,N_1641,N_1946);
xnor U2370 (N_2370,N_1754,N_1887);
and U2371 (N_2371,N_1832,N_1658);
xor U2372 (N_2372,N_1711,N_1502);
xnor U2373 (N_2373,N_1990,N_1516);
nor U2374 (N_2374,N_1903,N_1618);
nand U2375 (N_2375,N_1999,N_1757);
nand U2376 (N_2376,N_1831,N_1820);
and U2377 (N_2377,N_1708,N_1825);
or U2378 (N_2378,N_1761,N_1766);
nand U2379 (N_2379,N_1976,N_1934);
or U2380 (N_2380,N_1908,N_1648);
xor U2381 (N_2381,N_1960,N_1659);
xnor U2382 (N_2382,N_1500,N_1517);
nand U2383 (N_2383,N_1937,N_1922);
or U2384 (N_2384,N_1869,N_1535);
or U2385 (N_2385,N_1950,N_1834);
xor U2386 (N_2386,N_1611,N_1660);
xor U2387 (N_2387,N_1684,N_1941);
and U2388 (N_2388,N_1552,N_1537);
xnor U2389 (N_2389,N_1824,N_1719);
or U2390 (N_2390,N_1914,N_1552);
or U2391 (N_2391,N_1969,N_1733);
and U2392 (N_2392,N_1763,N_1866);
and U2393 (N_2393,N_1734,N_1730);
xnor U2394 (N_2394,N_1677,N_1556);
nand U2395 (N_2395,N_1879,N_1695);
xor U2396 (N_2396,N_1655,N_1542);
and U2397 (N_2397,N_1630,N_1528);
or U2398 (N_2398,N_1840,N_1887);
nor U2399 (N_2399,N_1796,N_1937);
and U2400 (N_2400,N_1510,N_1974);
and U2401 (N_2401,N_1872,N_1502);
xor U2402 (N_2402,N_1816,N_1627);
xnor U2403 (N_2403,N_1925,N_1733);
nor U2404 (N_2404,N_1676,N_1691);
and U2405 (N_2405,N_1727,N_1928);
xnor U2406 (N_2406,N_1929,N_1690);
xor U2407 (N_2407,N_1760,N_1553);
xor U2408 (N_2408,N_1661,N_1997);
nand U2409 (N_2409,N_1878,N_1994);
nand U2410 (N_2410,N_1925,N_1608);
and U2411 (N_2411,N_1666,N_1630);
xnor U2412 (N_2412,N_1732,N_1544);
or U2413 (N_2413,N_1712,N_1533);
and U2414 (N_2414,N_1705,N_1871);
nand U2415 (N_2415,N_1925,N_1511);
and U2416 (N_2416,N_1677,N_1669);
or U2417 (N_2417,N_1864,N_1771);
xnor U2418 (N_2418,N_1568,N_1740);
nand U2419 (N_2419,N_1933,N_1758);
nand U2420 (N_2420,N_1717,N_1500);
nor U2421 (N_2421,N_1967,N_1666);
nand U2422 (N_2422,N_1534,N_1800);
xor U2423 (N_2423,N_1516,N_1901);
xor U2424 (N_2424,N_1540,N_1611);
nand U2425 (N_2425,N_1850,N_1838);
xnor U2426 (N_2426,N_1899,N_1539);
xor U2427 (N_2427,N_1761,N_1928);
nor U2428 (N_2428,N_1617,N_1990);
or U2429 (N_2429,N_1807,N_1903);
xnor U2430 (N_2430,N_1738,N_1890);
xnor U2431 (N_2431,N_1935,N_1917);
or U2432 (N_2432,N_1523,N_1692);
nand U2433 (N_2433,N_1515,N_1565);
nor U2434 (N_2434,N_1835,N_1760);
xor U2435 (N_2435,N_1867,N_1747);
xnor U2436 (N_2436,N_1653,N_1584);
or U2437 (N_2437,N_1938,N_1656);
nand U2438 (N_2438,N_1525,N_1970);
xor U2439 (N_2439,N_1948,N_1993);
and U2440 (N_2440,N_1665,N_1630);
nor U2441 (N_2441,N_1903,N_1958);
or U2442 (N_2442,N_1613,N_1782);
xor U2443 (N_2443,N_1547,N_1827);
xor U2444 (N_2444,N_1807,N_1591);
and U2445 (N_2445,N_1557,N_1803);
nand U2446 (N_2446,N_1584,N_1556);
or U2447 (N_2447,N_1797,N_1852);
nand U2448 (N_2448,N_1927,N_1672);
or U2449 (N_2449,N_1567,N_1744);
nor U2450 (N_2450,N_1750,N_1824);
xnor U2451 (N_2451,N_1768,N_1786);
and U2452 (N_2452,N_1663,N_1595);
nor U2453 (N_2453,N_1708,N_1761);
and U2454 (N_2454,N_1516,N_1889);
nand U2455 (N_2455,N_1768,N_1657);
xnor U2456 (N_2456,N_1965,N_1997);
and U2457 (N_2457,N_1660,N_1731);
or U2458 (N_2458,N_1963,N_1622);
or U2459 (N_2459,N_1960,N_1990);
nand U2460 (N_2460,N_1570,N_1885);
nor U2461 (N_2461,N_1920,N_1767);
xnor U2462 (N_2462,N_1749,N_1795);
nor U2463 (N_2463,N_1589,N_1839);
and U2464 (N_2464,N_1573,N_1857);
nand U2465 (N_2465,N_1939,N_1794);
xnor U2466 (N_2466,N_1948,N_1881);
nand U2467 (N_2467,N_1878,N_1670);
xor U2468 (N_2468,N_1735,N_1722);
or U2469 (N_2469,N_1868,N_1517);
nor U2470 (N_2470,N_1772,N_1563);
or U2471 (N_2471,N_1866,N_1651);
nor U2472 (N_2472,N_1800,N_1937);
xnor U2473 (N_2473,N_1646,N_1865);
or U2474 (N_2474,N_1626,N_1753);
or U2475 (N_2475,N_1771,N_1539);
xor U2476 (N_2476,N_1980,N_1712);
or U2477 (N_2477,N_1765,N_1641);
xor U2478 (N_2478,N_1667,N_1935);
nor U2479 (N_2479,N_1875,N_1804);
nor U2480 (N_2480,N_1940,N_1611);
nor U2481 (N_2481,N_1939,N_1945);
nor U2482 (N_2482,N_1893,N_1792);
or U2483 (N_2483,N_1985,N_1769);
or U2484 (N_2484,N_1717,N_1522);
or U2485 (N_2485,N_1981,N_1833);
and U2486 (N_2486,N_1840,N_1720);
nand U2487 (N_2487,N_1883,N_1878);
nand U2488 (N_2488,N_1747,N_1754);
or U2489 (N_2489,N_1723,N_1905);
nand U2490 (N_2490,N_1759,N_1945);
or U2491 (N_2491,N_1750,N_1716);
xor U2492 (N_2492,N_1864,N_1873);
nand U2493 (N_2493,N_1901,N_1666);
xnor U2494 (N_2494,N_1976,N_1547);
or U2495 (N_2495,N_1621,N_1684);
or U2496 (N_2496,N_1654,N_1729);
or U2497 (N_2497,N_1876,N_1664);
nor U2498 (N_2498,N_1794,N_1889);
or U2499 (N_2499,N_1939,N_1912);
nand U2500 (N_2500,N_2318,N_2401);
or U2501 (N_2501,N_2387,N_2404);
nor U2502 (N_2502,N_2455,N_2268);
and U2503 (N_2503,N_2198,N_2237);
or U2504 (N_2504,N_2279,N_2476);
and U2505 (N_2505,N_2309,N_2248);
nor U2506 (N_2506,N_2283,N_2117);
or U2507 (N_2507,N_2008,N_2233);
or U2508 (N_2508,N_2157,N_2488);
nand U2509 (N_2509,N_2320,N_2332);
or U2510 (N_2510,N_2200,N_2411);
and U2511 (N_2511,N_2343,N_2124);
or U2512 (N_2512,N_2415,N_2354);
nor U2513 (N_2513,N_2060,N_2039);
and U2514 (N_2514,N_2175,N_2012);
and U2515 (N_2515,N_2095,N_2249);
and U2516 (N_2516,N_2254,N_2016);
nor U2517 (N_2517,N_2462,N_2451);
xor U2518 (N_2518,N_2286,N_2158);
and U2519 (N_2519,N_2435,N_2431);
or U2520 (N_2520,N_2085,N_2092);
or U2521 (N_2521,N_2033,N_2295);
nor U2522 (N_2522,N_2061,N_2099);
or U2523 (N_2523,N_2018,N_2024);
nand U2524 (N_2524,N_2135,N_2262);
nand U2525 (N_2525,N_2164,N_2166);
xnor U2526 (N_2526,N_2360,N_2465);
nand U2527 (N_2527,N_2251,N_2377);
or U2528 (N_2528,N_2376,N_2482);
and U2529 (N_2529,N_2110,N_2478);
nor U2530 (N_2530,N_2424,N_2289);
or U2531 (N_2531,N_2300,N_2074);
nor U2532 (N_2532,N_2456,N_2409);
or U2533 (N_2533,N_2473,N_2241);
and U2534 (N_2534,N_2052,N_2475);
and U2535 (N_2535,N_2336,N_2065);
nor U2536 (N_2536,N_2019,N_2304);
and U2537 (N_2537,N_2281,N_2073);
xnor U2538 (N_2538,N_2181,N_2162);
and U2539 (N_2539,N_2302,N_2408);
and U2540 (N_2540,N_2470,N_2407);
nand U2541 (N_2541,N_2458,N_2349);
or U2542 (N_2542,N_2252,N_2285);
and U2543 (N_2543,N_2063,N_2416);
xor U2544 (N_2544,N_2217,N_2463);
xnor U2545 (N_2545,N_2413,N_2297);
or U2546 (N_2546,N_2245,N_2059);
xnor U2547 (N_2547,N_2271,N_2007);
nor U2548 (N_2548,N_2139,N_2156);
xor U2549 (N_2549,N_2430,N_2194);
xor U2550 (N_2550,N_2179,N_2222);
xnor U2551 (N_2551,N_2352,N_2188);
or U2552 (N_2552,N_2098,N_2256);
nor U2553 (N_2553,N_2160,N_2134);
or U2554 (N_2554,N_2373,N_2312);
nor U2555 (N_2555,N_2153,N_2047);
nor U2556 (N_2556,N_2113,N_2428);
nand U2557 (N_2557,N_2357,N_2247);
and U2558 (N_2558,N_2288,N_2493);
nand U2559 (N_2559,N_2400,N_2174);
or U2560 (N_2560,N_2397,N_2319);
nor U2561 (N_2561,N_2005,N_2466);
nor U2562 (N_2562,N_2103,N_2266);
or U2563 (N_2563,N_2056,N_2468);
nand U2564 (N_2564,N_2064,N_2027);
and U2565 (N_2565,N_2253,N_2298);
xnor U2566 (N_2566,N_2452,N_2489);
and U2567 (N_2567,N_2322,N_2363);
nor U2568 (N_2568,N_2022,N_2031);
and U2569 (N_2569,N_2267,N_2136);
or U2570 (N_2570,N_2277,N_2205);
and U2571 (N_2571,N_2310,N_2333);
and U2572 (N_2572,N_2227,N_2111);
nor U2573 (N_2573,N_2076,N_2338);
nor U2574 (N_2574,N_2474,N_2161);
nand U2575 (N_2575,N_2138,N_2422);
or U2576 (N_2576,N_2044,N_2218);
nor U2577 (N_2577,N_2472,N_2183);
or U2578 (N_2578,N_2121,N_2429);
nand U2579 (N_2579,N_2128,N_2278);
nor U2580 (N_2580,N_2382,N_2030);
and U2581 (N_2581,N_2402,N_2447);
or U2582 (N_2582,N_2013,N_2096);
or U2583 (N_2583,N_2009,N_2045);
xor U2584 (N_2584,N_2214,N_2351);
nand U2585 (N_2585,N_2461,N_2480);
nor U2586 (N_2586,N_2077,N_2391);
or U2587 (N_2587,N_2058,N_2094);
or U2588 (N_2588,N_2341,N_2328);
or U2589 (N_2589,N_2444,N_2026);
nand U2590 (N_2590,N_2083,N_2107);
nand U2591 (N_2591,N_2151,N_2118);
nand U2592 (N_2592,N_2358,N_2051);
xor U2593 (N_2593,N_2119,N_2004);
and U2594 (N_2594,N_2287,N_2421);
nor U2595 (N_2595,N_2150,N_2196);
and U2596 (N_2596,N_2479,N_2152);
or U2597 (N_2597,N_2460,N_2317);
or U2598 (N_2598,N_2078,N_2362);
nor U2599 (N_2599,N_2316,N_2417);
or U2600 (N_2600,N_2326,N_2273);
xor U2601 (N_2601,N_2201,N_2055);
nor U2602 (N_2602,N_2323,N_2497);
nand U2603 (N_2603,N_2071,N_2220);
or U2604 (N_2604,N_2224,N_2142);
xnor U2605 (N_2605,N_2403,N_2471);
nand U2606 (N_2606,N_2192,N_2204);
and U2607 (N_2607,N_2356,N_2173);
nand U2608 (N_2608,N_2003,N_2330);
or U2609 (N_2609,N_2154,N_2399);
or U2610 (N_2610,N_2487,N_2315);
nand U2611 (N_2611,N_2305,N_2001);
nor U2612 (N_2612,N_2361,N_2017);
and U2613 (N_2613,N_2053,N_2091);
xnor U2614 (N_2614,N_2250,N_2388);
nand U2615 (N_2615,N_2086,N_2412);
xnor U2616 (N_2616,N_2477,N_2396);
nor U2617 (N_2617,N_2020,N_2427);
xor U2618 (N_2618,N_2195,N_2246);
and U2619 (N_2619,N_2042,N_2325);
or U2620 (N_2620,N_2108,N_2484);
nor U2621 (N_2621,N_2068,N_2303);
or U2622 (N_2622,N_2038,N_2155);
or U2623 (N_2623,N_2449,N_2420);
or U2624 (N_2624,N_2345,N_2442);
nor U2625 (N_2625,N_2378,N_2414);
nand U2626 (N_2626,N_2210,N_2359);
nand U2627 (N_2627,N_2106,N_2436);
and U2628 (N_2628,N_2331,N_2082);
and U2629 (N_2629,N_2184,N_2269);
xnor U2630 (N_2630,N_2219,N_2491);
and U2631 (N_2631,N_2127,N_2221);
or U2632 (N_2632,N_2425,N_2054);
or U2633 (N_2633,N_2386,N_2141);
nor U2634 (N_2634,N_2129,N_2228);
nor U2635 (N_2635,N_2464,N_2225);
nor U2636 (N_2636,N_2080,N_2132);
nor U2637 (N_2637,N_2393,N_2335);
nor U2638 (N_2638,N_2244,N_2314);
or U2639 (N_2639,N_2180,N_2259);
and U2640 (N_2640,N_2177,N_2353);
or U2641 (N_2641,N_2079,N_2105);
nor U2642 (N_2642,N_2120,N_2276);
nor U2643 (N_2643,N_2116,N_2000);
nor U2644 (N_2644,N_2454,N_2090);
xor U2645 (N_2645,N_2272,N_2239);
or U2646 (N_2646,N_2384,N_2087);
or U2647 (N_2647,N_2450,N_2236);
or U2648 (N_2648,N_2048,N_2440);
and U2649 (N_2649,N_2112,N_2035);
xnor U2650 (N_2650,N_2093,N_2370);
xnor U2651 (N_2651,N_2202,N_2122);
nand U2652 (N_2652,N_2002,N_2406);
nand U2653 (N_2653,N_2206,N_2226);
nand U2654 (N_2654,N_2131,N_2190);
nand U2655 (N_2655,N_2102,N_2235);
and U2656 (N_2656,N_2230,N_2028);
or U2657 (N_2657,N_2392,N_2213);
or U2658 (N_2658,N_2189,N_2037);
and U2659 (N_2659,N_2390,N_2398);
nand U2660 (N_2660,N_2496,N_2292);
nor U2661 (N_2661,N_2114,N_2197);
or U2662 (N_2662,N_2342,N_2263);
or U2663 (N_2663,N_2100,N_2495);
or U2664 (N_2664,N_2178,N_2344);
xor U2665 (N_2665,N_2258,N_2459);
nor U2666 (N_2666,N_2439,N_2232);
or U2667 (N_2667,N_2485,N_2294);
and U2668 (N_2668,N_2025,N_2355);
nand U2669 (N_2669,N_2010,N_2101);
xor U2670 (N_2670,N_2395,N_2216);
nor U2671 (N_2671,N_2275,N_2291);
xor U2672 (N_2672,N_2308,N_2149);
and U2673 (N_2673,N_2011,N_2270);
nand U2674 (N_2674,N_2032,N_2383);
or U2675 (N_2675,N_2115,N_2499);
nor U2676 (N_2676,N_2171,N_2394);
nor U2677 (N_2677,N_2062,N_2494);
xor U2678 (N_2678,N_2029,N_2257);
xnor U2679 (N_2679,N_2203,N_2324);
or U2680 (N_2680,N_2374,N_2321);
nand U2681 (N_2681,N_2015,N_2381);
nand U2682 (N_2682,N_2069,N_2147);
nor U2683 (N_2683,N_2209,N_2123);
and U2684 (N_2684,N_2170,N_2049);
xor U2685 (N_2685,N_2498,N_2438);
and U2686 (N_2686,N_2172,N_2492);
xor U2687 (N_2687,N_2176,N_2311);
and U2688 (N_2688,N_2337,N_2187);
nand U2689 (N_2689,N_2223,N_2293);
nor U2690 (N_2690,N_2169,N_2034);
xnor U2691 (N_2691,N_2334,N_2148);
xor U2692 (N_2692,N_2405,N_2261);
xor U2693 (N_2693,N_2453,N_2240);
xor U2694 (N_2694,N_2481,N_2264);
or U2695 (N_2695,N_2445,N_2014);
xnor U2696 (N_2696,N_2231,N_2075);
and U2697 (N_2697,N_2097,N_2089);
and U2698 (N_2698,N_2486,N_2284);
nand U2699 (N_2699,N_2299,N_2339);
or U2700 (N_2700,N_2307,N_2346);
nand U2701 (N_2701,N_2006,N_2457);
and U2702 (N_2702,N_2372,N_2469);
nand U2703 (N_2703,N_2347,N_2432);
nand U2704 (N_2704,N_2379,N_2242);
nand U2705 (N_2705,N_2081,N_2385);
xnor U2706 (N_2706,N_2490,N_2191);
nand U2707 (N_2707,N_2021,N_2369);
xnor U2708 (N_2708,N_2350,N_2296);
nand U2709 (N_2709,N_2234,N_2229);
or U2710 (N_2710,N_2274,N_2327);
nand U2711 (N_2711,N_2419,N_2133);
nand U2712 (N_2712,N_2426,N_2040);
xor U2713 (N_2713,N_2348,N_2441);
nand U2714 (N_2714,N_2104,N_2211);
nor U2715 (N_2715,N_2146,N_2329);
nand U2716 (N_2716,N_2313,N_2282);
xnor U2717 (N_2717,N_2036,N_2280);
and U2718 (N_2718,N_2088,N_2109);
nand U2719 (N_2719,N_2137,N_2389);
or U2720 (N_2720,N_2144,N_2367);
nand U2721 (N_2721,N_2290,N_2072);
nand U2722 (N_2722,N_2301,N_2043);
nand U2723 (N_2723,N_2306,N_2483);
nor U2724 (N_2724,N_2185,N_2410);
or U2725 (N_2725,N_2243,N_2165);
and U2726 (N_2726,N_2067,N_2041);
or U2727 (N_2727,N_2418,N_2380);
or U2728 (N_2728,N_2130,N_2050);
xor U2729 (N_2729,N_2265,N_2140);
nor U2730 (N_2730,N_2255,N_2365);
xnor U2731 (N_2731,N_2023,N_2145);
and U2732 (N_2732,N_2084,N_2168);
or U2733 (N_2733,N_2467,N_2238);
nor U2734 (N_2734,N_2375,N_2159);
or U2735 (N_2735,N_2434,N_2186);
xnor U2736 (N_2736,N_2046,N_2212);
nor U2737 (N_2737,N_2167,N_2143);
nor U2738 (N_2738,N_2125,N_2437);
and U2739 (N_2739,N_2364,N_2182);
or U2740 (N_2740,N_2126,N_2193);
nor U2741 (N_2741,N_2199,N_2433);
nand U2742 (N_2742,N_2208,N_2066);
nand U2743 (N_2743,N_2207,N_2215);
xnor U2744 (N_2744,N_2423,N_2340);
or U2745 (N_2745,N_2371,N_2260);
or U2746 (N_2746,N_2070,N_2057);
or U2747 (N_2747,N_2443,N_2448);
and U2748 (N_2748,N_2368,N_2366);
nor U2749 (N_2749,N_2446,N_2163);
nand U2750 (N_2750,N_2152,N_2384);
nor U2751 (N_2751,N_2083,N_2494);
xnor U2752 (N_2752,N_2120,N_2105);
xnor U2753 (N_2753,N_2383,N_2221);
xor U2754 (N_2754,N_2005,N_2155);
nor U2755 (N_2755,N_2090,N_2068);
and U2756 (N_2756,N_2019,N_2498);
xnor U2757 (N_2757,N_2388,N_2259);
nor U2758 (N_2758,N_2387,N_2111);
nand U2759 (N_2759,N_2440,N_2207);
and U2760 (N_2760,N_2162,N_2017);
or U2761 (N_2761,N_2488,N_2438);
xor U2762 (N_2762,N_2273,N_2014);
and U2763 (N_2763,N_2021,N_2413);
nor U2764 (N_2764,N_2009,N_2323);
xnor U2765 (N_2765,N_2444,N_2279);
or U2766 (N_2766,N_2339,N_2241);
or U2767 (N_2767,N_2140,N_2472);
xnor U2768 (N_2768,N_2470,N_2307);
or U2769 (N_2769,N_2086,N_2328);
and U2770 (N_2770,N_2477,N_2123);
and U2771 (N_2771,N_2205,N_2026);
and U2772 (N_2772,N_2232,N_2054);
or U2773 (N_2773,N_2356,N_2412);
and U2774 (N_2774,N_2147,N_2063);
and U2775 (N_2775,N_2460,N_2274);
or U2776 (N_2776,N_2454,N_2195);
xor U2777 (N_2777,N_2471,N_2486);
or U2778 (N_2778,N_2017,N_2426);
nand U2779 (N_2779,N_2110,N_2322);
xnor U2780 (N_2780,N_2304,N_2271);
xor U2781 (N_2781,N_2104,N_2086);
nand U2782 (N_2782,N_2220,N_2207);
xor U2783 (N_2783,N_2175,N_2468);
or U2784 (N_2784,N_2412,N_2444);
xor U2785 (N_2785,N_2004,N_2375);
or U2786 (N_2786,N_2197,N_2340);
xnor U2787 (N_2787,N_2343,N_2283);
and U2788 (N_2788,N_2239,N_2111);
nand U2789 (N_2789,N_2488,N_2258);
or U2790 (N_2790,N_2018,N_2457);
xor U2791 (N_2791,N_2363,N_2378);
nor U2792 (N_2792,N_2089,N_2369);
nand U2793 (N_2793,N_2179,N_2050);
nor U2794 (N_2794,N_2460,N_2026);
nand U2795 (N_2795,N_2345,N_2477);
nor U2796 (N_2796,N_2294,N_2443);
and U2797 (N_2797,N_2141,N_2229);
and U2798 (N_2798,N_2370,N_2273);
nand U2799 (N_2799,N_2078,N_2189);
xnor U2800 (N_2800,N_2472,N_2006);
and U2801 (N_2801,N_2382,N_2011);
and U2802 (N_2802,N_2041,N_2464);
xor U2803 (N_2803,N_2459,N_2337);
or U2804 (N_2804,N_2034,N_2106);
or U2805 (N_2805,N_2117,N_2060);
nor U2806 (N_2806,N_2107,N_2050);
nand U2807 (N_2807,N_2171,N_2121);
xnor U2808 (N_2808,N_2060,N_2183);
xnor U2809 (N_2809,N_2064,N_2353);
nand U2810 (N_2810,N_2466,N_2421);
nor U2811 (N_2811,N_2486,N_2060);
and U2812 (N_2812,N_2286,N_2395);
and U2813 (N_2813,N_2287,N_2032);
xor U2814 (N_2814,N_2000,N_2293);
nor U2815 (N_2815,N_2172,N_2320);
or U2816 (N_2816,N_2259,N_2165);
nor U2817 (N_2817,N_2196,N_2094);
and U2818 (N_2818,N_2261,N_2475);
and U2819 (N_2819,N_2127,N_2223);
or U2820 (N_2820,N_2431,N_2467);
xnor U2821 (N_2821,N_2074,N_2084);
nor U2822 (N_2822,N_2160,N_2227);
and U2823 (N_2823,N_2282,N_2452);
or U2824 (N_2824,N_2133,N_2134);
and U2825 (N_2825,N_2046,N_2313);
nand U2826 (N_2826,N_2233,N_2351);
xor U2827 (N_2827,N_2321,N_2006);
nor U2828 (N_2828,N_2030,N_2380);
or U2829 (N_2829,N_2323,N_2241);
nand U2830 (N_2830,N_2360,N_2452);
nor U2831 (N_2831,N_2199,N_2145);
xor U2832 (N_2832,N_2416,N_2186);
or U2833 (N_2833,N_2474,N_2012);
nor U2834 (N_2834,N_2208,N_2088);
or U2835 (N_2835,N_2319,N_2194);
or U2836 (N_2836,N_2002,N_2061);
nand U2837 (N_2837,N_2434,N_2420);
nand U2838 (N_2838,N_2179,N_2252);
nor U2839 (N_2839,N_2374,N_2171);
and U2840 (N_2840,N_2200,N_2211);
or U2841 (N_2841,N_2010,N_2216);
or U2842 (N_2842,N_2142,N_2117);
and U2843 (N_2843,N_2469,N_2365);
nand U2844 (N_2844,N_2310,N_2219);
nand U2845 (N_2845,N_2484,N_2257);
nand U2846 (N_2846,N_2266,N_2164);
nand U2847 (N_2847,N_2402,N_2219);
xor U2848 (N_2848,N_2320,N_2138);
nor U2849 (N_2849,N_2462,N_2126);
and U2850 (N_2850,N_2163,N_2084);
and U2851 (N_2851,N_2237,N_2420);
nand U2852 (N_2852,N_2260,N_2199);
nand U2853 (N_2853,N_2221,N_2157);
xnor U2854 (N_2854,N_2445,N_2156);
and U2855 (N_2855,N_2055,N_2461);
and U2856 (N_2856,N_2253,N_2301);
or U2857 (N_2857,N_2214,N_2376);
xor U2858 (N_2858,N_2351,N_2276);
nand U2859 (N_2859,N_2447,N_2360);
nand U2860 (N_2860,N_2003,N_2055);
xor U2861 (N_2861,N_2296,N_2164);
or U2862 (N_2862,N_2044,N_2064);
or U2863 (N_2863,N_2139,N_2402);
nand U2864 (N_2864,N_2378,N_2394);
xor U2865 (N_2865,N_2420,N_2011);
nand U2866 (N_2866,N_2062,N_2266);
xnor U2867 (N_2867,N_2458,N_2273);
nand U2868 (N_2868,N_2064,N_2159);
nor U2869 (N_2869,N_2049,N_2056);
nand U2870 (N_2870,N_2197,N_2076);
xor U2871 (N_2871,N_2075,N_2088);
nor U2872 (N_2872,N_2071,N_2162);
or U2873 (N_2873,N_2267,N_2406);
and U2874 (N_2874,N_2067,N_2312);
and U2875 (N_2875,N_2405,N_2338);
xnor U2876 (N_2876,N_2152,N_2032);
and U2877 (N_2877,N_2018,N_2296);
or U2878 (N_2878,N_2060,N_2119);
xnor U2879 (N_2879,N_2382,N_2448);
xor U2880 (N_2880,N_2139,N_2264);
nand U2881 (N_2881,N_2407,N_2496);
nor U2882 (N_2882,N_2343,N_2216);
xnor U2883 (N_2883,N_2458,N_2030);
nor U2884 (N_2884,N_2155,N_2347);
or U2885 (N_2885,N_2170,N_2015);
nor U2886 (N_2886,N_2346,N_2016);
and U2887 (N_2887,N_2124,N_2293);
nand U2888 (N_2888,N_2318,N_2333);
nor U2889 (N_2889,N_2241,N_2496);
and U2890 (N_2890,N_2226,N_2164);
and U2891 (N_2891,N_2425,N_2377);
or U2892 (N_2892,N_2473,N_2165);
nand U2893 (N_2893,N_2113,N_2372);
nor U2894 (N_2894,N_2390,N_2239);
nand U2895 (N_2895,N_2233,N_2129);
xor U2896 (N_2896,N_2362,N_2090);
nand U2897 (N_2897,N_2388,N_2026);
nand U2898 (N_2898,N_2486,N_2272);
or U2899 (N_2899,N_2407,N_2281);
nor U2900 (N_2900,N_2102,N_2316);
nor U2901 (N_2901,N_2483,N_2053);
nand U2902 (N_2902,N_2159,N_2024);
or U2903 (N_2903,N_2028,N_2356);
xnor U2904 (N_2904,N_2363,N_2362);
or U2905 (N_2905,N_2245,N_2166);
and U2906 (N_2906,N_2035,N_2262);
nand U2907 (N_2907,N_2065,N_2220);
nand U2908 (N_2908,N_2371,N_2173);
nand U2909 (N_2909,N_2101,N_2480);
and U2910 (N_2910,N_2403,N_2175);
nor U2911 (N_2911,N_2303,N_2291);
nor U2912 (N_2912,N_2349,N_2178);
or U2913 (N_2913,N_2466,N_2382);
or U2914 (N_2914,N_2304,N_2457);
or U2915 (N_2915,N_2190,N_2201);
nand U2916 (N_2916,N_2019,N_2319);
or U2917 (N_2917,N_2164,N_2019);
xnor U2918 (N_2918,N_2310,N_2265);
nand U2919 (N_2919,N_2304,N_2285);
and U2920 (N_2920,N_2231,N_2211);
nand U2921 (N_2921,N_2415,N_2018);
nand U2922 (N_2922,N_2119,N_2194);
nand U2923 (N_2923,N_2106,N_2459);
and U2924 (N_2924,N_2477,N_2302);
nand U2925 (N_2925,N_2350,N_2229);
nand U2926 (N_2926,N_2399,N_2345);
xnor U2927 (N_2927,N_2229,N_2118);
nor U2928 (N_2928,N_2254,N_2435);
nand U2929 (N_2929,N_2426,N_2103);
xnor U2930 (N_2930,N_2289,N_2462);
nand U2931 (N_2931,N_2230,N_2074);
or U2932 (N_2932,N_2278,N_2396);
xor U2933 (N_2933,N_2153,N_2477);
nor U2934 (N_2934,N_2221,N_2149);
or U2935 (N_2935,N_2432,N_2393);
nand U2936 (N_2936,N_2241,N_2402);
or U2937 (N_2937,N_2199,N_2219);
xnor U2938 (N_2938,N_2280,N_2450);
and U2939 (N_2939,N_2138,N_2404);
and U2940 (N_2940,N_2048,N_2304);
nand U2941 (N_2941,N_2113,N_2351);
xnor U2942 (N_2942,N_2421,N_2338);
nor U2943 (N_2943,N_2178,N_2290);
or U2944 (N_2944,N_2459,N_2297);
nor U2945 (N_2945,N_2161,N_2193);
xnor U2946 (N_2946,N_2430,N_2164);
nor U2947 (N_2947,N_2146,N_2036);
nor U2948 (N_2948,N_2120,N_2318);
and U2949 (N_2949,N_2480,N_2408);
and U2950 (N_2950,N_2211,N_2387);
or U2951 (N_2951,N_2209,N_2258);
or U2952 (N_2952,N_2316,N_2215);
nand U2953 (N_2953,N_2252,N_2005);
nor U2954 (N_2954,N_2106,N_2460);
nor U2955 (N_2955,N_2260,N_2354);
and U2956 (N_2956,N_2464,N_2449);
and U2957 (N_2957,N_2346,N_2436);
and U2958 (N_2958,N_2228,N_2115);
and U2959 (N_2959,N_2335,N_2033);
and U2960 (N_2960,N_2207,N_2199);
xnor U2961 (N_2961,N_2085,N_2044);
nor U2962 (N_2962,N_2255,N_2035);
nor U2963 (N_2963,N_2326,N_2164);
nand U2964 (N_2964,N_2347,N_2309);
xor U2965 (N_2965,N_2397,N_2250);
or U2966 (N_2966,N_2420,N_2023);
or U2967 (N_2967,N_2121,N_2116);
nand U2968 (N_2968,N_2485,N_2052);
xnor U2969 (N_2969,N_2251,N_2457);
or U2970 (N_2970,N_2204,N_2222);
nor U2971 (N_2971,N_2465,N_2060);
nor U2972 (N_2972,N_2179,N_2278);
and U2973 (N_2973,N_2126,N_2299);
and U2974 (N_2974,N_2326,N_2264);
or U2975 (N_2975,N_2270,N_2356);
nand U2976 (N_2976,N_2051,N_2210);
or U2977 (N_2977,N_2446,N_2391);
xnor U2978 (N_2978,N_2149,N_2281);
or U2979 (N_2979,N_2189,N_2326);
nand U2980 (N_2980,N_2060,N_2339);
xnor U2981 (N_2981,N_2094,N_2109);
xor U2982 (N_2982,N_2258,N_2210);
nor U2983 (N_2983,N_2452,N_2226);
nand U2984 (N_2984,N_2086,N_2124);
nor U2985 (N_2985,N_2120,N_2383);
and U2986 (N_2986,N_2289,N_2489);
xnor U2987 (N_2987,N_2104,N_2256);
and U2988 (N_2988,N_2149,N_2451);
nor U2989 (N_2989,N_2090,N_2482);
nand U2990 (N_2990,N_2303,N_2452);
nor U2991 (N_2991,N_2390,N_2314);
xnor U2992 (N_2992,N_2224,N_2033);
nand U2993 (N_2993,N_2269,N_2448);
or U2994 (N_2994,N_2060,N_2380);
xnor U2995 (N_2995,N_2057,N_2007);
xnor U2996 (N_2996,N_2069,N_2410);
xnor U2997 (N_2997,N_2376,N_2317);
xor U2998 (N_2998,N_2221,N_2485);
nand U2999 (N_2999,N_2172,N_2243);
or UO_0 (O_0,N_2585,N_2799);
or UO_1 (O_1,N_2755,N_2950);
nor UO_2 (O_2,N_2544,N_2648);
nand UO_3 (O_3,N_2660,N_2628);
xor UO_4 (O_4,N_2654,N_2980);
nor UO_5 (O_5,N_2719,N_2655);
or UO_6 (O_6,N_2578,N_2632);
nand UO_7 (O_7,N_2905,N_2598);
nand UO_8 (O_8,N_2785,N_2514);
nor UO_9 (O_9,N_2732,N_2965);
or UO_10 (O_10,N_2715,N_2646);
xor UO_11 (O_11,N_2503,N_2545);
or UO_12 (O_12,N_2706,N_2639);
and UO_13 (O_13,N_2582,N_2864);
xnor UO_14 (O_14,N_2767,N_2900);
xor UO_15 (O_15,N_2998,N_2721);
nor UO_16 (O_16,N_2635,N_2659);
nor UO_17 (O_17,N_2929,N_2768);
or UO_18 (O_18,N_2524,N_2580);
xnor UO_19 (O_19,N_2939,N_2849);
nor UO_20 (O_20,N_2695,N_2845);
nand UO_21 (O_21,N_2787,N_2831);
nor UO_22 (O_22,N_2948,N_2528);
or UO_23 (O_23,N_2525,N_2903);
and UO_24 (O_24,N_2570,N_2685);
or UO_25 (O_25,N_2969,N_2681);
and UO_26 (O_26,N_2772,N_2739);
xor UO_27 (O_27,N_2761,N_2677);
and UO_28 (O_28,N_2671,N_2815);
xnor UO_29 (O_29,N_2577,N_2724);
nor UO_30 (O_30,N_2579,N_2581);
nand UO_31 (O_31,N_2691,N_2723);
or UO_32 (O_32,N_2667,N_2968);
and UO_33 (O_33,N_2971,N_2593);
and UO_34 (O_34,N_2989,N_2559);
or UO_35 (O_35,N_2919,N_2633);
and UO_36 (O_36,N_2614,N_2918);
nand UO_37 (O_37,N_2658,N_2661);
and UO_38 (O_38,N_2981,N_2820);
or UO_39 (O_39,N_2777,N_2534);
nor UO_40 (O_40,N_2923,N_2573);
nand UO_41 (O_41,N_2729,N_2836);
nor UO_42 (O_42,N_2589,N_2835);
or UO_43 (O_43,N_2696,N_2862);
or UO_44 (O_44,N_2674,N_2773);
nor UO_45 (O_45,N_2676,N_2844);
xor UO_46 (O_46,N_2801,N_2941);
nor UO_47 (O_47,N_2857,N_2978);
xnor UO_48 (O_48,N_2507,N_2557);
xnor UO_49 (O_49,N_2657,N_2811);
or UO_50 (O_50,N_2853,N_2793);
nand UO_51 (O_51,N_2623,N_2642);
nor UO_52 (O_52,N_2631,N_2832);
nand UO_53 (O_53,N_2595,N_2610);
and UO_54 (O_54,N_2531,N_2523);
or UO_55 (O_55,N_2966,N_2871);
nand UO_56 (O_56,N_2925,N_2931);
or UO_57 (O_57,N_2613,N_2548);
nand UO_58 (O_58,N_2500,N_2526);
or UO_59 (O_59,N_2842,N_2553);
and UO_60 (O_60,N_2776,N_2899);
and UO_61 (O_61,N_2607,N_2775);
xor UO_62 (O_62,N_2795,N_2975);
nor UO_63 (O_63,N_2837,N_2973);
and UO_64 (O_64,N_2834,N_2764);
and UO_65 (O_65,N_2656,N_2673);
xor UO_66 (O_66,N_2621,N_2819);
or UO_67 (O_67,N_2904,N_2812);
nor UO_68 (O_68,N_2885,N_2560);
or UO_69 (O_69,N_2783,N_2850);
or UO_70 (O_70,N_2908,N_2569);
nor UO_71 (O_71,N_2596,N_2802);
and UO_72 (O_72,N_2826,N_2823);
and UO_73 (O_73,N_2940,N_2502);
xor UO_74 (O_74,N_2769,N_2562);
nor UO_75 (O_75,N_2599,N_2814);
or UO_76 (O_76,N_2513,N_2907);
nor UO_77 (O_77,N_2993,N_2917);
xnor UO_78 (O_78,N_2745,N_2554);
nand UO_79 (O_79,N_2716,N_2920);
nor UO_80 (O_80,N_2800,N_2587);
xnor UO_81 (O_81,N_2692,N_2780);
nor UO_82 (O_82,N_2540,N_2670);
or UO_83 (O_83,N_2572,N_2816);
and UO_84 (O_84,N_2895,N_2882);
and UO_85 (O_85,N_2731,N_2663);
nand UO_86 (O_86,N_2797,N_2898);
nand UO_87 (O_87,N_2703,N_2792);
xor UO_88 (O_88,N_2839,N_2722);
nor UO_89 (O_89,N_2924,N_2901);
nand UO_90 (O_90,N_2701,N_2851);
nor UO_91 (O_91,N_2699,N_2710);
and UO_92 (O_92,N_2763,N_2694);
xnor UO_93 (O_93,N_2956,N_2913);
nor UO_94 (O_94,N_2693,N_2597);
nor UO_95 (O_95,N_2563,N_2818);
and UO_96 (O_96,N_2571,N_2720);
nand UO_97 (O_97,N_2958,N_2912);
nor UO_98 (O_98,N_2652,N_2932);
xnor UO_99 (O_99,N_2927,N_2742);
xor UO_100 (O_100,N_2873,N_2986);
xnor UO_101 (O_101,N_2584,N_2515);
nor UO_102 (O_102,N_2840,N_2959);
and UO_103 (O_103,N_2627,N_2915);
and UO_104 (O_104,N_2888,N_2675);
xor UO_105 (O_105,N_2626,N_2946);
xnor UO_106 (O_106,N_2892,N_2561);
xnor UO_107 (O_107,N_2556,N_2957);
nand UO_108 (O_108,N_2592,N_2704);
nor UO_109 (O_109,N_2841,N_2821);
xnor UO_110 (O_110,N_2734,N_2700);
and UO_111 (O_111,N_2884,N_2872);
or UO_112 (O_112,N_2609,N_2537);
xor UO_113 (O_113,N_2756,N_2875);
and UO_114 (O_114,N_2879,N_2859);
xor UO_115 (O_115,N_2758,N_2991);
nor UO_116 (O_116,N_2615,N_2711);
nand UO_117 (O_117,N_2668,N_2977);
nor UO_118 (O_118,N_2605,N_2672);
nand UO_119 (O_119,N_2748,N_2770);
or UO_120 (O_120,N_2619,N_2687);
nor UO_121 (O_121,N_2805,N_2542);
and UO_122 (O_122,N_2603,N_2678);
xnor UO_123 (O_123,N_2921,N_2664);
and UO_124 (O_124,N_2911,N_2974);
nor UO_125 (O_125,N_2539,N_2535);
xnor UO_126 (O_126,N_2751,N_2527);
nand UO_127 (O_127,N_2789,N_2618);
xnor UO_128 (O_128,N_2830,N_2988);
nand UO_129 (O_129,N_2890,N_2521);
xor UO_130 (O_130,N_2897,N_2883);
xnor UO_131 (O_131,N_2590,N_2717);
and UO_132 (O_132,N_2854,N_2766);
xor UO_133 (O_133,N_2817,N_2788);
and UO_134 (O_134,N_2952,N_2602);
and UO_135 (O_135,N_2551,N_2804);
xor UO_136 (O_136,N_2983,N_2600);
nor UO_137 (O_137,N_2867,N_2987);
xor UO_138 (O_138,N_2807,N_2868);
nand UO_139 (O_139,N_2709,N_2650);
nand UO_140 (O_140,N_2738,N_2606);
xor UO_141 (O_141,N_2887,N_2848);
xnor UO_142 (O_142,N_2889,N_2586);
and UO_143 (O_143,N_2855,N_2982);
xor UO_144 (O_144,N_2749,N_2746);
nand UO_145 (O_145,N_2622,N_2612);
and UO_146 (O_146,N_2530,N_2881);
nand UO_147 (O_147,N_2798,N_2645);
nor UO_148 (O_148,N_2653,N_2962);
xor UO_149 (O_149,N_2926,N_2630);
and UO_150 (O_150,N_2778,N_2866);
nand UO_151 (O_151,N_2794,N_2647);
xor UO_152 (O_152,N_2999,N_2733);
or UO_153 (O_153,N_2679,N_2617);
xnor UO_154 (O_154,N_2935,N_2752);
xor UO_155 (O_155,N_2822,N_2992);
nor UO_156 (O_156,N_2979,N_2714);
and UO_157 (O_157,N_2552,N_2730);
nor UO_158 (O_158,N_2666,N_2519);
or UO_159 (O_159,N_2906,N_2786);
xnor UO_160 (O_160,N_2942,N_2643);
nand UO_161 (O_161,N_2533,N_2970);
nand UO_162 (O_162,N_2914,N_2833);
nor UO_163 (O_163,N_2928,N_2747);
nand UO_164 (O_164,N_2953,N_2985);
nor UO_165 (O_165,N_2930,N_2697);
nor UO_166 (O_166,N_2508,N_2856);
xnor UO_167 (O_167,N_2662,N_2624);
and UO_168 (O_168,N_2636,N_2689);
xnor UO_169 (O_169,N_2808,N_2543);
xnor UO_170 (O_170,N_2705,N_2790);
or UO_171 (O_171,N_2984,N_2594);
or UO_172 (O_172,N_2640,N_2753);
and UO_173 (O_173,N_2869,N_2810);
nor UO_174 (O_174,N_2634,N_2549);
xor UO_175 (O_175,N_2860,N_2760);
xnor UO_176 (O_176,N_2774,N_2847);
xor UO_177 (O_177,N_2852,N_2686);
xnor UO_178 (O_178,N_2954,N_2967);
xnor UO_179 (O_179,N_2809,N_2501);
xnor UO_180 (O_180,N_2737,N_2604);
xor UO_181 (O_181,N_2690,N_2964);
nand UO_182 (O_182,N_2997,N_2791);
nand UO_183 (O_183,N_2902,N_2891);
or UO_184 (O_184,N_2637,N_2726);
nor UO_185 (O_185,N_2963,N_2861);
nor UO_186 (O_186,N_2547,N_2916);
xor UO_187 (O_187,N_2558,N_2713);
nand UO_188 (O_188,N_2520,N_2894);
nor UO_189 (O_189,N_2909,N_2566);
xor UO_190 (O_190,N_2995,N_2516);
or UO_191 (O_191,N_2684,N_2910);
and UO_192 (O_192,N_2506,N_2575);
and UO_193 (O_193,N_2994,N_2990);
or UO_194 (O_194,N_2625,N_2517);
xor UO_195 (O_195,N_2877,N_2735);
or UO_196 (O_196,N_2943,N_2870);
nand UO_197 (O_197,N_2555,N_2806);
nand UO_198 (O_198,N_2649,N_2796);
or UO_199 (O_199,N_2951,N_2665);
xnor UO_200 (O_200,N_2608,N_2949);
nor UO_201 (O_201,N_2876,N_2736);
and UO_202 (O_202,N_2765,N_2880);
or UO_203 (O_203,N_2510,N_2996);
nor UO_204 (O_204,N_2504,N_2863);
nor UO_205 (O_205,N_2682,N_2583);
and UO_206 (O_206,N_2829,N_2698);
or UO_207 (O_207,N_2505,N_2743);
nand UO_208 (O_208,N_2874,N_2538);
or UO_209 (O_209,N_2550,N_2532);
and UO_210 (O_210,N_2638,N_2536);
nor UO_211 (O_211,N_2574,N_2803);
nor UO_212 (O_212,N_2824,N_2782);
xnor UO_213 (O_213,N_2683,N_2707);
nand UO_214 (O_214,N_2976,N_2757);
nand UO_215 (O_215,N_2759,N_2813);
or UO_216 (O_216,N_2838,N_2779);
nand UO_217 (O_217,N_2576,N_2955);
or UO_218 (O_218,N_2518,N_2893);
nor UO_219 (O_219,N_2568,N_2896);
nor UO_220 (O_220,N_2762,N_2827);
and UO_221 (O_221,N_2944,N_2740);
nand UO_222 (O_222,N_2522,N_2858);
and UO_223 (O_223,N_2616,N_2509);
and UO_224 (O_224,N_2727,N_2933);
nand UO_225 (O_225,N_2922,N_2529);
and UO_226 (O_226,N_2961,N_2972);
or UO_227 (O_227,N_2728,N_2754);
nand UO_228 (O_228,N_2865,N_2878);
and UO_229 (O_229,N_2937,N_2629);
nand UO_230 (O_230,N_2718,N_2947);
xnor UO_231 (O_231,N_2511,N_2644);
and UO_232 (O_232,N_2541,N_2591);
nand UO_233 (O_233,N_2771,N_2828);
or UO_234 (O_234,N_2708,N_2784);
nand UO_235 (O_235,N_2567,N_2688);
nand UO_236 (O_236,N_2669,N_2846);
xnor UO_237 (O_237,N_2741,N_2825);
nor UO_238 (O_238,N_2611,N_2744);
and UO_239 (O_239,N_2565,N_2564);
xor UO_240 (O_240,N_2512,N_2620);
nor UO_241 (O_241,N_2886,N_2651);
or UO_242 (O_242,N_2702,N_2938);
nand UO_243 (O_243,N_2960,N_2680);
or UO_244 (O_244,N_2945,N_2934);
xnor UO_245 (O_245,N_2750,N_2936);
or UO_246 (O_246,N_2725,N_2546);
and UO_247 (O_247,N_2781,N_2588);
nand UO_248 (O_248,N_2601,N_2712);
and UO_249 (O_249,N_2641,N_2843);
nor UO_250 (O_250,N_2840,N_2719);
nor UO_251 (O_251,N_2535,N_2670);
or UO_252 (O_252,N_2774,N_2502);
or UO_253 (O_253,N_2990,N_2548);
or UO_254 (O_254,N_2892,N_2841);
nor UO_255 (O_255,N_2648,N_2913);
and UO_256 (O_256,N_2695,N_2775);
nand UO_257 (O_257,N_2888,N_2698);
xnor UO_258 (O_258,N_2657,N_2926);
nor UO_259 (O_259,N_2506,N_2857);
xor UO_260 (O_260,N_2639,N_2901);
nand UO_261 (O_261,N_2975,N_2888);
or UO_262 (O_262,N_2684,N_2735);
and UO_263 (O_263,N_2510,N_2750);
and UO_264 (O_264,N_2748,N_2700);
nand UO_265 (O_265,N_2872,N_2610);
nand UO_266 (O_266,N_2990,N_2744);
and UO_267 (O_267,N_2514,N_2565);
or UO_268 (O_268,N_2539,N_2646);
and UO_269 (O_269,N_2904,N_2562);
xor UO_270 (O_270,N_2942,N_2561);
nor UO_271 (O_271,N_2871,N_2738);
xnor UO_272 (O_272,N_2589,N_2515);
xor UO_273 (O_273,N_2643,N_2522);
xor UO_274 (O_274,N_2969,N_2868);
or UO_275 (O_275,N_2947,N_2608);
or UO_276 (O_276,N_2600,N_2607);
and UO_277 (O_277,N_2823,N_2971);
xor UO_278 (O_278,N_2936,N_2717);
xnor UO_279 (O_279,N_2658,N_2529);
or UO_280 (O_280,N_2719,N_2935);
nand UO_281 (O_281,N_2615,N_2622);
and UO_282 (O_282,N_2950,N_2829);
and UO_283 (O_283,N_2574,N_2603);
nor UO_284 (O_284,N_2997,N_2934);
xor UO_285 (O_285,N_2606,N_2912);
and UO_286 (O_286,N_2703,N_2524);
or UO_287 (O_287,N_2710,N_2638);
nand UO_288 (O_288,N_2544,N_2682);
xnor UO_289 (O_289,N_2772,N_2546);
nor UO_290 (O_290,N_2749,N_2781);
nor UO_291 (O_291,N_2859,N_2736);
and UO_292 (O_292,N_2712,N_2952);
xnor UO_293 (O_293,N_2978,N_2874);
nor UO_294 (O_294,N_2512,N_2787);
nor UO_295 (O_295,N_2822,N_2886);
nor UO_296 (O_296,N_2841,N_2978);
nor UO_297 (O_297,N_2818,N_2756);
nand UO_298 (O_298,N_2667,N_2625);
and UO_299 (O_299,N_2592,N_2641);
nor UO_300 (O_300,N_2806,N_2531);
xnor UO_301 (O_301,N_2761,N_2762);
and UO_302 (O_302,N_2504,N_2970);
or UO_303 (O_303,N_2525,N_2593);
and UO_304 (O_304,N_2832,N_2780);
and UO_305 (O_305,N_2648,N_2571);
nand UO_306 (O_306,N_2841,N_2913);
nor UO_307 (O_307,N_2777,N_2947);
xor UO_308 (O_308,N_2808,N_2643);
or UO_309 (O_309,N_2647,N_2639);
xnor UO_310 (O_310,N_2653,N_2757);
or UO_311 (O_311,N_2960,N_2519);
nand UO_312 (O_312,N_2687,N_2616);
nand UO_313 (O_313,N_2688,N_2921);
or UO_314 (O_314,N_2675,N_2755);
nor UO_315 (O_315,N_2574,N_2835);
nand UO_316 (O_316,N_2634,N_2973);
nand UO_317 (O_317,N_2872,N_2788);
nand UO_318 (O_318,N_2587,N_2729);
xnor UO_319 (O_319,N_2747,N_2694);
and UO_320 (O_320,N_2726,N_2535);
xor UO_321 (O_321,N_2529,N_2597);
and UO_322 (O_322,N_2563,N_2989);
nand UO_323 (O_323,N_2581,N_2857);
and UO_324 (O_324,N_2809,N_2841);
nor UO_325 (O_325,N_2671,N_2854);
and UO_326 (O_326,N_2836,N_2981);
xor UO_327 (O_327,N_2939,N_2708);
nand UO_328 (O_328,N_2840,N_2862);
and UO_329 (O_329,N_2814,N_2956);
nand UO_330 (O_330,N_2681,N_2764);
and UO_331 (O_331,N_2876,N_2519);
xnor UO_332 (O_332,N_2641,N_2934);
nor UO_333 (O_333,N_2905,N_2664);
nand UO_334 (O_334,N_2680,N_2677);
nand UO_335 (O_335,N_2986,N_2928);
nor UO_336 (O_336,N_2964,N_2729);
nand UO_337 (O_337,N_2826,N_2642);
or UO_338 (O_338,N_2633,N_2566);
nor UO_339 (O_339,N_2679,N_2529);
and UO_340 (O_340,N_2669,N_2737);
nor UO_341 (O_341,N_2548,N_2917);
xor UO_342 (O_342,N_2950,N_2521);
or UO_343 (O_343,N_2502,N_2890);
xor UO_344 (O_344,N_2684,N_2650);
and UO_345 (O_345,N_2597,N_2565);
and UO_346 (O_346,N_2804,N_2714);
nand UO_347 (O_347,N_2896,N_2527);
nand UO_348 (O_348,N_2602,N_2647);
nand UO_349 (O_349,N_2698,N_2782);
or UO_350 (O_350,N_2804,N_2656);
nor UO_351 (O_351,N_2814,N_2853);
and UO_352 (O_352,N_2828,N_2955);
xnor UO_353 (O_353,N_2871,N_2758);
xor UO_354 (O_354,N_2909,N_2726);
or UO_355 (O_355,N_2704,N_2942);
xor UO_356 (O_356,N_2611,N_2721);
nor UO_357 (O_357,N_2791,N_2879);
xnor UO_358 (O_358,N_2916,N_2790);
nand UO_359 (O_359,N_2798,N_2734);
nor UO_360 (O_360,N_2830,N_2975);
and UO_361 (O_361,N_2900,N_2974);
xor UO_362 (O_362,N_2984,N_2743);
nand UO_363 (O_363,N_2607,N_2826);
xor UO_364 (O_364,N_2778,N_2800);
nand UO_365 (O_365,N_2594,N_2553);
xor UO_366 (O_366,N_2824,N_2967);
nand UO_367 (O_367,N_2838,N_2814);
nor UO_368 (O_368,N_2757,N_2545);
nand UO_369 (O_369,N_2935,N_2607);
and UO_370 (O_370,N_2503,N_2972);
xor UO_371 (O_371,N_2686,N_2679);
nor UO_372 (O_372,N_2563,N_2672);
nand UO_373 (O_373,N_2958,N_2938);
nand UO_374 (O_374,N_2547,N_2842);
or UO_375 (O_375,N_2755,N_2606);
nor UO_376 (O_376,N_2901,N_2852);
xnor UO_377 (O_377,N_2547,N_2871);
and UO_378 (O_378,N_2524,N_2776);
nand UO_379 (O_379,N_2803,N_2975);
nor UO_380 (O_380,N_2745,N_2803);
or UO_381 (O_381,N_2866,N_2857);
and UO_382 (O_382,N_2917,N_2980);
nand UO_383 (O_383,N_2662,N_2970);
nand UO_384 (O_384,N_2570,N_2980);
nand UO_385 (O_385,N_2985,N_2886);
and UO_386 (O_386,N_2925,N_2609);
nand UO_387 (O_387,N_2631,N_2593);
or UO_388 (O_388,N_2738,N_2821);
and UO_389 (O_389,N_2908,N_2957);
and UO_390 (O_390,N_2562,N_2603);
or UO_391 (O_391,N_2524,N_2759);
nand UO_392 (O_392,N_2881,N_2631);
and UO_393 (O_393,N_2812,N_2941);
nor UO_394 (O_394,N_2797,N_2607);
xor UO_395 (O_395,N_2690,N_2992);
and UO_396 (O_396,N_2806,N_2916);
and UO_397 (O_397,N_2771,N_2546);
xnor UO_398 (O_398,N_2678,N_2916);
xnor UO_399 (O_399,N_2700,N_2586);
nand UO_400 (O_400,N_2854,N_2672);
nor UO_401 (O_401,N_2660,N_2650);
and UO_402 (O_402,N_2863,N_2668);
nand UO_403 (O_403,N_2849,N_2914);
xor UO_404 (O_404,N_2743,N_2838);
and UO_405 (O_405,N_2698,N_2878);
nor UO_406 (O_406,N_2640,N_2557);
and UO_407 (O_407,N_2781,N_2815);
and UO_408 (O_408,N_2854,N_2802);
xor UO_409 (O_409,N_2664,N_2930);
and UO_410 (O_410,N_2638,N_2660);
nand UO_411 (O_411,N_2540,N_2535);
and UO_412 (O_412,N_2740,N_2867);
xnor UO_413 (O_413,N_2738,N_2782);
and UO_414 (O_414,N_2722,N_2768);
xor UO_415 (O_415,N_2967,N_2585);
or UO_416 (O_416,N_2817,N_2762);
nor UO_417 (O_417,N_2756,N_2771);
nand UO_418 (O_418,N_2835,N_2902);
or UO_419 (O_419,N_2858,N_2813);
or UO_420 (O_420,N_2619,N_2911);
xnor UO_421 (O_421,N_2918,N_2963);
or UO_422 (O_422,N_2659,N_2782);
nor UO_423 (O_423,N_2916,N_2973);
nor UO_424 (O_424,N_2980,N_2897);
nor UO_425 (O_425,N_2615,N_2682);
xnor UO_426 (O_426,N_2610,N_2966);
or UO_427 (O_427,N_2864,N_2554);
nor UO_428 (O_428,N_2780,N_2926);
and UO_429 (O_429,N_2559,N_2724);
nand UO_430 (O_430,N_2927,N_2905);
nand UO_431 (O_431,N_2553,N_2701);
xnor UO_432 (O_432,N_2960,N_2896);
nand UO_433 (O_433,N_2930,N_2958);
xor UO_434 (O_434,N_2997,N_2808);
xnor UO_435 (O_435,N_2500,N_2968);
and UO_436 (O_436,N_2660,N_2966);
nor UO_437 (O_437,N_2695,N_2559);
nand UO_438 (O_438,N_2718,N_2811);
and UO_439 (O_439,N_2950,N_2565);
or UO_440 (O_440,N_2695,N_2846);
and UO_441 (O_441,N_2638,N_2855);
nand UO_442 (O_442,N_2936,N_2837);
and UO_443 (O_443,N_2607,N_2894);
nand UO_444 (O_444,N_2938,N_2799);
nor UO_445 (O_445,N_2843,N_2942);
nand UO_446 (O_446,N_2543,N_2579);
nor UO_447 (O_447,N_2609,N_2708);
xnor UO_448 (O_448,N_2647,N_2856);
nand UO_449 (O_449,N_2866,N_2505);
xnor UO_450 (O_450,N_2573,N_2918);
xor UO_451 (O_451,N_2571,N_2598);
xnor UO_452 (O_452,N_2976,N_2875);
nand UO_453 (O_453,N_2723,N_2669);
xor UO_454 (O_454,N_2855,N_2952);
and UO_455 (O_455,N_2945,N_2610);
xnor UO_456 (O_456,N_2822,N_2637);
xor UO_457 (O_457,N_2749,N_2974);
or UO_458 (O_458,N_2715,N_2979);
or UO_459 (O_459,N_2842,N_2946);
and UO_460 (O_460,N_2564,N_2952);
xnor UO_461 (O_461,N_2549,N_2668);
nor UO_462 (O_462,N_2505,N_2620);
nor UO_463 (O_463,N_2623,N_2527);
and UO_464 (O_464,N_2730,N_2528);
nor UO_465 (O_465,N_2532,N_2955);
xnor UO_466 (O_466,N_2855,N_2854);
nor UO_467 (O_467,N_2630,N_2971);
xor UO_468 (O_468,N_2631,N_2877);
xor UO_469 (O_469,N_2711,N_2592);
or UO_470 (O_470,N_2551,N_2566);
xnor UO_471 (O_471,N_2732,N_2821);
nor UO_472 (O_472,N_2917,N_2730);
or UO_473 (O_473,N_2589,N_2556);
xor UO_474 (O_474,N_2615,N_2961);
nor UO_475 (O_475,N_2652,N_2647);
nand UO_476 (O_476,N_2899,N_2701);
and UO_477 (O_477,N_2801,N_2983);
xnor UO_478 (O_478,N_2808,N_2657);
nand UO_479 (O_479,N_2738,N_2772);
xor UO_480 (O_480,N_2961,N_2569);
xor UO_481 (O_481,N_2535,N_2859);
xnor UO_482 (O_482,N_2768,N_2866);
nor UO_483 (O_483,N_2521,N_2778);
xnor UO_484 (O_484,N_2544,N_2894);
and UO_485 (O_485,N_2733,N_2820);
or UO_486 (O_486,N_2572,N_2628);
and UO_487 (O_487,N_2605,N_2737);
nand UO_488 (O_488,N_2688,N_2620);
nor UO_489 (O_489,N_2900,N_2736);
and UO_490 (O_490,N_2530,N_2788);
xnor UO_491 (O_491,N_2697,N_2754);
xnor UO_492 (O_492,N_2873,N_2861);
or UO_493 (O_493,N_2928,N_2865);
xnor UO_494 (O_494,N_2506,N_2980);
or UO_495 (O_495,N_2826,N_2640);
nand UO_496 (O_496,N_2673,N_2636);
or UO_497 (O_497,N_2835,N_2685);
nor UO_498 (O_498,N_2869,N_2544);
xnor UO_499 (O_499,N_2580,N_2993);
endmodule