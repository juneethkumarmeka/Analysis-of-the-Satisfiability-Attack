module basic_1500_15000_2000_75_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_889,In_221);
nand U1 (N_1,In_456,In_915);
nor U2 (N_2,In_232,In_524);
xor U3 (N_3,In_114,In_1162);
nor U4 (N_4,In_1481,In_1129);
nor U5 (N_5,In_1107,In_240);
and U6 (N_6,In_795,In_7);
and U7 (N_7,In_296,In_1121);
or U8 (N_8,In_1390,In_1232);
xor U9 (N_9,In_257,In_554);
nand U10 (N_10,In_390,In_778);
and U11 (N_11,In_0,In_1013);
xnor U12 (N_12,In_1073,In_767);
xor U13 (N_13,In_991,In_1347);
and U14 (N_14,In_12,In_25);
or U15 (N_15,In_319,In_1180);
nand U16 (N_16,In_634,In_1152);
and U17 (N_17,In_1236,In_1366);
nor U18 (N_18,In_1295,In_1456);
nand U19 (N_19,In_1490,In_1382);
nand U20 (N_20,In_657,In_452);
nand U21 (N_21,In_1161,In_649);
or U22 (N_22,In_1171,In_1282);
or U23 (N_23,In_275,In_1402);
xor U24 (N_24,In_723,In_1483);
or U25 (N_25,In_1420,In_850);
nand U26 (N_26,In_17,In_336);
nand U27 (N_27,In_960,In_303);
and U28 (N_28,In_822,In_529);
and U29 (N_29,In_1406,In_220);
nand U30 (N_30,In_412,In_1423);
nor U31 (N_31,In_994,In_383);
or U32 (N_32,In_1351,In_971);
xnor U33 (N_33,In_414,In_483);
nand U34 (N_34,In_1218,In_1345);
nor U35 (N_35,In_1296,In_478);
or U36 (N_36,In_169,In_227);
and U37 (N_37,In_1316,In_274);
xor U38 (N_38,In_1197,In_980);
and U39 (N_39,In_92,In_345);
nor U40 (N_40,In_909,In_987);
or U41 (N_41,In_838,In_941);
nand U42 (N_42,In_37,In_477);
nor U43 (N_43,In_702,In_985);
nor U44 (N_44,In_103,In_1393);
nand U45 (N_45,In_497,In_156);
nand U46 (N_46,In_66,In_1480);
and U47 (N_47,In_918,In_1496);
and U48 (N_48,In_983,In_794);
nor U49 (N_49,In_727,In_392);
or U50 (N_50,In_661,In_1243);
and U51 (N_51,In_570,In_1082);
xnor U52 (N_52,In_893,In_13);
and U53 (N_53,In_609,In_141);
or U54 (N_54,In_1223,In_1207);
and U55 (N_55,In_1247,In_413);
nand U56 (N_56,In_736,In_871);
nand U57 (N_57,In_1168,In_1126);
xor U58 (N_58,In_83,In_1169);
and U59 (N_59,In_984,In_69);
nand U60 (N_60,In_803,In_445);
or U61 (N_61,In_434,In_544);
nand U62 (N_62,In_1115,In_117);
nor U63 (N_63,In_614,In_481);
nand U64 (N_64,In_466,In_552);
nor U65 (N_65,In_196,In_1220);
nor U66 (N_66,In_40,In_690);
and U67 (N_67,In_1014,In_792);
and U68 (N_68,In_1302,In_1128);
nand U69 (N_69,In_1454,In_317);
nand U70 (N_70,In_1445,In_449);
or U71 (N_71,In_407,In_1384);
nor U72 (N_72,In_1053,In_272);
xor U73 (N_73,In_438,In_753);
nor U74 (N_74,In_1084,In_31);
nor U75 (N_75,In_1422,In_642);
and U76 (N_76,In_1353,In_1159);
xnor U77 (N_77,In_122,In_853);
and U78 (N_78,In_1348,In_841);
and U79 (N_79,In_1387,In_1269);
nand U80 (N_80,In_836,In_1335);
or U81 (N_81,In_338,In_940);
or U82 (N_82,In_1015,In_835);
or U83 (N_83,In_808,In_1036);
nand U84 (N_84,In_1367,In_709);
and U85 (N_85,In_258,In_140);
and U86 (N_86,In_582,In_1);
and U87 (N_87,In_1333,In_996);
and U88 (N_88,In_694,In_115);
nand U89 (N_89,In_185,In_430);
nor U90 (N_90,In_1285,In_1432);
xnor U91 (N_91,In_273,In_16);
and U92 (N_92,In_998,In_1185);
nor U93 (N_93,In_1440,In_260);
xnor U94 (N_94,In_57,In_658);
xnor U95 (N_95,In_160,In_520);
and U96 (N_96,In_1192,In_953);
xnor U97 (N_97,In_1144,In_168);
nor U98 (N_98,In_837,In_701);
nor U99 (N_99,In_118,In_815);
or U100 (N_100,In_1000,In_300);
xnor U101 (N_101,In_1158,In_113);
nor U102 (N_102,In_1149,In_217);
nor U103 (N_103,In_558,In_1424);
xnor U104 (N_104,In_968,In_1239);
and U105 (N_105,In_359,In_228);
xnor U106 (N_106,In_1277,In_305);
nand U107 (N_107,In_1441,In_1140);
xor U108 (N_108,In_954,In_485);
nand U109 (N_109,In_239,In_1352);
xor U110 (N_110,In_385,In_900);
or U111 (N_111,In_1326,In_1256);
or U112 (N_112,In_71,In_1116);
or U113 (N_113,In_1461,In_436);
xor U114 (N_114,In_1446,In_656);
and U115 (N_115,In_395,In_139);
and U116 (N_116,In_503,In_11);
xnor U117 (N_117,In_1146,In_313);
or U118 (N_118,In_206,In_310);
nor U119 (N_119,In_1179,In_19);
nor U120 (N_120,In_358,In_493);
or U121 (N_121,In_1315,In_705);
or U122 (N_122,In_1125,In_665);
xnor U123 (N_123,In_574,In_138);
or U124 (N_124,In_732,In_107);
nand U125 (N_125,In_1381,In_1359);
nor U126 (N_126,In_919,In_1404);
and U127 (N_127,In_699,In_93);
or U128 (N_128,In_1221,In_958);
nor U129 (N_129,In_890,In_1078);
nand U130 (N_130,In_324,In_667);
nand U131 (N_131,In_112,In_687);
nor U132 (N_132,In_734,In_856);
and U133 (N_133,In_223,In_212);
and U134 (N_134,In_910,In_1368);
and U135 (N_135,In_1254,In_200);
nand U136 (N_136,In_1486,In_788);
nor U137 (N_137,In_1061,In_1273);
nor U138 (N_138,In_1211,In_1259);
xnor U139 (N_139,In_646,In_376);
and U140 (N_140,In_1485,In_1099);
xor U141 (N_141,In_510,In_110);
or U142 (N_142,In_207,In_301);
xnor U143 (N_143,In_278,In_1439);
or U144 (N_144,In_819,In_410);
or U145 (N_145,In_1244,In_583);
nand U146 (N_146,In_1322,In_451);
or U147 (N_147,In_823,In_879);
nand U148 (N_148,In_482,In_796);
and U149 (N_149,In_526,In_32);
xor U150 (N_150,In_427,In_86);
nor U151 (N_151,In_840,In_1190);
nor U152 (N_152,In_1091,In_572);
xnor U153 (N_153,In_981,In_525);
xnor U154 (N_154,In_1350,In_264);
nor U155 (N_155,In_997,In_952);
nand U156 (N_156,In_1012,In_1327);
nor U157 (N_157,In_678,In_589);
and U158 (N_158,In_63,In_1317);
xnor U159 (N_159,In_455,In_302);
or U160 (N_160,In_78,In_1085);
nand U161 (N_161,In_533,In_213);
or U162 (N_162,In_1045,In_719);
xor U163 (N_163,In_209,In_760);
and U164 (N_164,In_1066,In_462);
nor U165 (N_165,In_721,In_151);
and U166 (N_166,In_774,In_882);
nor U167 (N_167,In_95,In_77);
or U168 (N_168,In_1238,In_903);
xnor U169 (N_169,In_1249,In_577);
nand U170 (N_170,In_486,In_454);
and U171 (N_171,In_1070,In_628);
or U172 (N_172,In_1009,In_888);
nand U173 (N_173,In_624,In_193);
xor U174 (N_174,In_1139,In_235);
nand U175 (N_175,In_1134,In_770);
xnor U176 (N_176,In_361,In_153);
or U177 (N_177,In_172,In_1253);
or U178 (N_178,In_1438,In_867);
xor U179 (N_179,In_54,In_757);
nand U180 (N_180,In_431,In_584);
or U181 (N_181,In_1370,In_907);
or U182 (N_182,In_560,In_859);
or U183 (N_183,In_1203,In_1164);
nand U184 (N_184,In_873,In_1356);
nor U185 (N_185,In_892,In_204);
nand U186 (N_186,In_548,In_946);
and U187 (N_187,In_959,In_1160);
nor U188 (N_188,In_1414,In_322);
and U189 (N_189,In_1464,In_1064);
and U190 (N_190,In_601,In_1004);
xnor U191 (N_191,In_834,In_253);
or U192 (N_192,In_740,In_72);
xnor U193 (N_193,In_1191,In_722);
or U194 (N_194,In_546,In_52);
and U195 (N_195,In_1275,In_1148);
nand U196 (N_196,In_780,In_370);
xnor U197 (N_197,In_801,In_1418);
xnor U198 (N_198,In_1241,In_513);
and U199 (N_199,In_743,In_143);
nor U200 (N_200,In_96,In_844);
nand U201 (N_201,N_184,N_61);
xor U202 (N_202,N_60,In_147);
nand U203 (N_203,In_136,In_26);
nor U204 (N_204,N_139,In_1453);
xor U205 (N_205,In_1475,In_350);
nand U206 (N_206,In_606,In_651);
and U207 (N_207,In_304,In_748);
xor U208 (N_208,In_556,In_1437);
xor U209 (N_209,In_259,In_1339);
or U210 (N_210,In_371,In_30);
and U211 (N_211,In_327,In_905);
xor U212 (N_212,In_429,N_157);
nor U213 (N_213,In_1391,In_18);
and U214 (N_214,In_1154,In_579);
or U215 (N_215,In_1261,N_22);
nor U216 (N_216,In_1122,N_120);
nor U217 (N_217,In_632,N_144);
and U218 (N_218,In_564,In_962);
nand U219 (N_219,In_202,In_365);
and U220 (N_220,N_194,In_1386);
nor U221 (N_221,In_1330,N_169);
nor U222 (N_222,In_6,In_276);
or U223 (N_223,In_1195,In_1213);
nor U224 (N_224,In_1110,In_435);
and U225 (N_225,In_501,N_11);
nand U226 (N_226,In_682,In_403);
xnor U227 (N_227,In_1262,N_54);
nand U228 (N_228,In_80,N_148);
nand U229 (N_229,In_1305,N_133);
xnor U230 (N_230,In_192,In_250);
and U231 (N_231,In_1200,In_176);
and U232 (N_232,In_1398,In_1242);
nand U233 (N_233,N_197,In_1289);
and U234 (N_234,In_9,In_81);
or U235 (N_235,In_1205,In_314);
or U236 (N_236,In_783,In_364);
xor U237 (N_237,In_1369,In_693);
xnor U238 (N_238,In_588,In_440);
nor U239 (N_239,N_128,In_1246);
nand U240 (N_240,In_424,In_639);
xnor U241 (N_241,In_1032,In_189);
or U242 (N_242,N_163,In_963);
nor U243 (N_243,In_813,In_831);
xnor U244 (N_244,In_1362,In_75);
and U245 (N_245,In_1119,In_730);
nand U246 (N_246,In_1396,In_1355);
nor U247 (N_247,In_800,In_126);
or U248 (N_248,In_97,In_473);
and U249 (N_249,In_1380,In_495);
nand U250 (N_250,In_394,In_947);
and U251 (N_251,N_28,In_331);
nand U252 (N_252,N_109,In_1231);
or U253 (N_253,In_1312,In_928);
and U254 (N_254,N_69,In_236);
and U255 (N_255,In_1033,In_1199);
xor U256 (N_256,In_88,In_1271);
or U257 (N_257,In_1021,N_89);
xnor U258 (N_258,In_2,In_1095);
and U259 (N_259,N_114,In_1314);
nor U260 (N_260,In_166,N_134);
and U261 (N_261,In_862,In_1307);
or U262 (N_262,N_193,In_951);
xnor U263 (N_263,N_187,In_161);
nor U264 (N_264,In_620,In_567);
or U265 (N_265,In_1329,In_541);
xnor U266 (N_266,In_1344,In_1103);
nand U267 (N_267,In_1167,N_12);
or U268 (N_268,In_870,In_128);
or U269 (N_269,In_1166,In_186);
or U270 (N_270,In_1142,In_750);
nor U271 (N_271,In_388,In_746);
xor U272 (N_272,N_108,In_349);
xnor U273 (N_273,In_598,N_165);
xor U274 (N_274,N_150,In_664);
or U275 (N_275,In_599,In_377);
nand U276 (N_276,In_784,In_474);
or U277 (N_277,In_681,In_182);
nor U278 (N_278,In_712,In_608);
and U279 (N_279,N_145,In_726);
or U280 (N_280,In_1057,In_1034);
and U281 (N_281,In_179,N_124);
xor U282 (N_282,In_858,In_540);
and U283 (N_283,N_104,In_1338);
or U284 (N_284,In_1360,In_1092);
nand U285 (N_285,In_669,In_605);
xor U286 (N_286,In_84,In_293);
nor U287 (N_287,In_929,In_47);
xnor U288 (N_288,In_171,In_1052);
nand U289 (N_289,In_828,In_1008);
nor U290 (N_290,N_171,In_34);
and U291 (N_291,In_1044,In_1340);
and U292 (N_292,In_233,In_861);
nor U293 (N_293,In_308,In_1071);
or U294 (N_294,N_71,In_471);
nand U295 (N_295,In_1300,In_85);
nor U296 (N_296,In_676,In_165);
nor U297 (N_297,In_629,N_159);
or U298 (N_298,N_146,In_591);
nor U299 (N_299,In_1358,In_1299);
and U300 (N_300,In_469,In_864);
xor U301 (N_301,In_1448,In_417);
or U302 (N_302,N_107,In_1467);
or U303 (N_303,In_1006,In_1497);
nor U304 (N_304,In_863,In_728);
nor U305 (N_305,In_286,In_1026);
and U306 (N_306,In_1143,In_36);
nor U307 (N_307,In_1047,In_936);
nor U308 (N_308,N_195,In_1173);
and U309 (N_309,In_433,In_340);
or U310 (N_310,In_504,In_492);
nor U311 (N_311,In_362,In_1365);
and U312 (N_312,In_428,In_152);
nor U313 (N_313,N_5,In_74);
nor U314 (N_314,In_1002,In_98);
and U315 (N_315,In_1318,In_876);
xnor U316 (N_316,In_183,N_35);
xnor U317 (N_317,In_295,In_1007);
or U318 (N_318,In_1498,In_8);
nand U319 (N_319,In_851,In_1039);
nand U320 (N_320,In_1260,N_188);
or U321 (N_321,In_342,In_993);
nor U322 (N_322,In_398,In_937);
and U323 (N_323,In_706,N_95);
nand U324 (N_324,In_270,In_44);
nand U325 (N_325,N_176,In_966);
nor U326 (N_326,In_1240,N_179);
xor U327 (N_327,In_1194,In_1417);
or U328 (N_328,In_1489,In_1266);
and U329 (N_329,In_269,N_86);
nor U330 (N_330,In_886,In_1074);
xnor U331 (N_331,In_1463,In_1124);
or U332 (N_332,In_617,In_640);
xor U333 (N_333,In_593,In_729);
nand U334 (N_334,In_218,In_1263);
nor U335 (N_335,In_214,In_306);
xnor U336 (N_336,In_268,In_557);
nand U337 (N_337,In_814,In_982);
nand U338 (N_338,In_245,N_154);
nor U339 (N_339,In_852,In_224);
nand U340 (N_340,N_119,In_244);
or U341 (N_341,In_1482,In_976);
or U342 (N_342,In_562,In_880);
and U343 (N_343,N_115,In_150);
and U344 (N_344,In_46,In_1201);
and U345 (N_345,N_24,In_970);
and U346 (N_346,In_901,N_185);
and U347 (N_347,In_847,In_865);
xor U348 (N_348,In_580,In_333);
nand U349 (N_349,In_1250,In_839);
nor U350 (N_350,In_177,In_255);
xnor U351 (N_351,In_1287,In_881);
nand U352 (N_352,In_1206,In_511);
or U353 (N_353,In_1090,In_1258);
xnor U354 (N_354,N_170,In_924);
nor U355 (N_355,In_453,In_348);
xor U356 (N_356,In_1388,N_18);
and U357 (N_357,In_318,N_111);
nand U358 (N_358,In_789,N_110);
nor U359 (N_359,In_986,In_137);
or U360 (N_360,In_1443,In_120);
nor U361 (N_361,In_1077,In_1165);
or U362 (N_362,In_1229,N_47);
or U363 (N_363,In_1080,In_480);
nor U364 (N_364,N_125,In_1117);
nor U365 (N_365,In_432,In_1449);
xnor U366 (N_366,In_488,In_842);
and U367 (N_367,In_374,In_1476);
xnor U368 (N_368,N_68,In_779);
and U369 (N_369,In_369,In_1215);
nand U370 (N_370,In_1291,In_499);
or U371 (N_371,N_90,In_1109);
nand U372 (N_372,In_472,In_967);
nor U373 (N_373,In_1421,In_400);
and U374 (N_374,In_1293,In_521);
and U375 (N_375,In_1429,N_156);
xor U376 (N_376,In_849,In_555);
or U377 (N_377,In_360,In_536);
or U378 (N_378,In_500,In_1048);
and U379 (N_379,In_1474,In_505);
xor U380 (N_380,N_99,In_612);
xor U381 (N_381,In_515,In_1016);
nand U382 (N_382,In_116,In_1175);
nor U383 (N_383,In_1410,In_496);
or U384 (N_384,In_479,In_39);
nor U385 (N_385,In_149,N_30);
nand U386 (N_386,In_1172,In_1403);
or U387 (N_387,In_804,In_1471);
or U388 (N_388,In_53,In_1083);
nor U389 (N_389,In_1212,In_973);
nand U390 (N_390,In_595,In_906);
xor U391 (N_391,In_696,In_592);
nor U392 (N_392,N_27,In_697);
or U393 (N_393,In_1138,In_1466);
or U394 (N_394,In_222,In_124);
or U395 (N_395,In_761,In_1187);
or U396 (N_396,In_1428,In_597);
and U397 (N_397,In_1478,In_616);
xnor U398 (N_398,In_381,In_1184);
nand U399 (N_399,N_151,In_325);
xnor U400 (N_400,In_754,In_1460);
nand U401 (N_401,N_75,N_122);
nor U402 (N_402,N_64,N_208);
nand U403 (N_403,In_829,In_1176);
xor U404 (N_404,In_307,N_191);
and U405 (N_405,N_189,In_446);
or U406 (N_406,N_2,N_355);
and U407 (N_407,N_10,In_104);
nor U408 (N_408,In_1430,N_172);
nand U409 (N_409,In_191,N_392);
and U410 (N_410,N_186,N_379);
nor U411 (N_411,In_1136,In_1145);
and U412 (N_412,In_1286,In_633);
or U413 (N_413,In_76,In_568);
nor U414 (N_414,In_1216,In_777);
nor U415 (N_415,In_1068,N_97);
nand U416 (N_416,In_550,In_1208);
xnor U417 (N_417,In_547,In_27);
nor U418 (N_418,In_442,N_83);
or U419 (N_419,N_142,N_205);
xor U420 (N_420,In_912,In_242);
and U421 (N_421,In_1038,In_1086);
nor U422 (N_422,In_389,In_1063);
nand U423 (N_423,In_1059,N_235);
or U424 (N_424,In_463,In_448);
xor U425 (N_425,In_675,In_917);
nand U426 (N_426,In_1067,In_1188);
nor U427 (N_427,In_1412,In_460);
xnor U428 (N_428,In_802,N_129);
and U429 (N_429,In_630,In_421);
nand U430 (N_430,In_1493,In_1377);
nor U431 (N_431,In_194,In_1284);
or U432 (N_432,In_89,N_326);
and U433 (N_433,In_742,In_798);
nor U434 (N_434,In_1030,In_527);
and U435 (N_435,N_305,N_141);
and U436 (N_436,N_221,In_816);
or U437 (N_437,In_312,N_92);
nor U438 (N_438,In_101,In_1373);
nand U439 (N_439,In_315,In_523);
or U440 (N_440,N_256,In_1321);
nand U441 (N_441,N_297,N_267);
or U442 (N_442,In_957,In_91);
or U443 (N_443,In_1298,N_285);
and U444 (N_444,N_395,In_576);
and U445 (N_445,N_56,N_9);
xor U446 (N_446,In_238,N_166);
xnor U447 (N_447,In_1096,In_718);
and U448 (N_448,N_204,In_70);
nand U449 (N_449,N_102,N_106);
xnor U450 (N_450,In_1442,N_135);
and U451 (N_451,In_710,N_174);
and U452 (N_452,N_8,In_195);
nor U453 (N_453,N_351,N_230);
and U454 (N_454,In_1328,In_1405);
nor U455 (N_455,In_955,In_363);
xnor U456 (N_456,N_85,In_387);
or U457 (N_457,In_393,In_964);
xor U458 (N_458,In_1280,N_67);
and U459 (N_459,N_66,N_152);
nand U460 (N_460,N_335,In_1235);
xor U461 (N_461,In_1005,In_437);
nand U462 (N_462,In_755,N_39);
or U463 (N_463,In_354,In_372);
nor U464 (N_464,N_344,In_566);
xnor U465 (N_465,In_869,In_668);
or U466 (N_466,N_76,In_762);
xnor U467 (N_467,N_373,N_264);
nand U468 (N_468,In_1469,In_752);
nor U469 (N_469,In_956,N_367);
or U470 (N_470,In_1320,N_43);
nand U471 (N_471,In_163,In_711);
and U472 (N_472,In_356,In_677);
nor U473 (N_473,In_1342,N_295);
and U474 (N_474,In_375,In_447);
nor U475 (N_475,In_45,N_359);
or U476 (N_476,In_514,In_1267);
or U477 (N_477,In_1025,In_1306);
xnor U478 (N_478,In_787,In_974);
nand U479 (N_479,In_686,In_105);
xnor U480 (N_480,N_36,In_1290);
nand U481 (N_481,In_1450,In_1156);
and U482 (N_482,N_4,N_399);
or U483 (N_483,In_545,In_1094);
xor U484 (N_484,In_467,In_49);
nor U485 (N_485,In_704,In_1087);
nor U486 (N_486,N_240,N_319);
xnor U487 (N_487,N_57,In_1484);
nand U488 (N_488,N_350,In_1304);
nand U489 (N_489,In_1472,In_771);
nand U490 (N_490,In_248,In_923);
nor U491 (N_491,In_90,N_140);
nor U492 (N_492,N_182,N_370);
nand U493 (N_493,N_279,N_312);
nor U494 (N_494,In_226,In_507);
and U495 (N_495,N_127,N_173);
nor U496 (N_496,In_411,In_1399);
or U497 (N_497,In_1313,In_843);
xor U498 (N_498,N_250,N_183);
nor U499 (N_499,In_127,In_1120);
and U500 (N_500,In_498,In_1245);
xnor U501 (N_501,In_1270,In_781);
nand U502 (N_502,In_1076,In_190);
xnor U503 (N_503,In_1470,N_132);
nand U504 (N_504,In_58,In_625);
and U505 (N_505,N_210,In_875);
nor U506 (N_506,In_368,In_698);
nor U507 (N_507,N_271,N_322);
and U508 (N_508,N_32,In_216);
xnor U509 (N_509,In_3,N_374);
xor U510 (N_510,In_464,N_53);
nor U511 (N_511,In_321,N_88);
nand U512 (N_512,In_908,In_1444);
xnor U513 (N_513,In_807,In_1311);
and U514 (N_514,In_1042,N_263);
nand U515 (N_515,In_1363,In_280);
nand U516 (N_516,In_341,In_645);
and U517 (N_517,In_581,In_67);
xor U518 (N_518,In_399,N_383);
nand U519 (N_519,In_670,N_311);
and U520 (N_520,In_1431,N_254);
or U521 (N_521,In_284,In_1272);
xnor U522 (N_522,In_386,In_1452);
xnor U523 (N_523,In_1135,In_299);
or U524 (N_524,In_180,In_1319);
and U525 (N_525,In_33,In_878);
or U526 (N_526,N_51,N_357);
or U527 (N_527,In_1349,In_234);
or U528 (N_528,N_377,In_820);
xnor U529 (N_529,In_1037,In_181);
xor U530 (N_530,In_1357,N_313);
xnor U531 (N_531,In_692,In_1310);
nand U532 (N_532,In_465,In_1219);
xor U533 (N_533,In_607,In_159);
xor U534 (N_534,N_397,N_223);
and U535 (N_535,In_99,In_785);
xnor U536 (N_536,In_1354,In_62);
or U537 (N_537,N_298,In_637);
xor U538 (N_538,In_323,In_59);
or U539 (N_539,N_162,N_237);
nand U540 (N_540,In_100,In_211);
or U541 (N_541,N_274,In_231);
or U542 (N_542,In_703,N_323);
and U543 (N_543,In_573,In_1451);
or U544 (N_544,N_255,In_1459);
xor U545 (N_545,In_700,In_491);
or U546 (N_546,In_1447,N_136);
nand U547 (N_547,N_177,In_825);
xor U548 (N_548,In_1465,In_737);
or U549 (N_549,In_261,In_441);
xor U550 (N_550,In_426,In_82);
xor U551 (N_551,N_78,In_738);
or U552 (N_552,In_768,N_257);
nor U553 (N_553,In_811,In_895);
or U554 (N_554,In_855,N_218);
nand U555 (N_555,N_288,In_961);
or U556 (N_556,N_363,In_575);
and U557 (N_557,In_158,In_531);
xor U558 (N_558,N_345,In_346);
nor U559 (N_559,In_565,N_273);
and U560 (N_560,N_249,In_549);
nand U561 (N_561,In_1408,N_45);
nor U562 (N_562,In_1098,In_1274);
xnor U563 (N_563,In_23,In_635);
nand U564 (N_564,In_79,N_368);
xor U565 (N_565,In_857,In_713);
or U566 (N_566,In_751,In_1043);
xnor U567 (N_567,In_10,In_532);
xor U568 (N_568,In_334,In_600);
nand U569 (N_569,N_59,In_109);
nand U570 (N_570,In_590,In_157);
nor U571 (N_571,N_253,In_717);
or U572 (N_572,N_126,In_594);
nor U573 (N_573,N_283,N_16);
nand U574 (N_574,In_806,N_84);
or U575 (N_575,In_316,In_154);
or U576 (N_576,In_406,In_289);
xor U577 (N_577,In_1106,N_390);
and U578 (N_578,In_1458,In_263);
nor U579 (N_579,In_1494,In_1224);
xnor U580 (N_580,In_1325,N_277);
and U581 (N_581,In_123,In_1436);
nor U582 (N_582,In_285,In_174);
xor U583 (N_583,N_213,In_1276);
or U584 (N_584,In_1341,N_378);
nand U585 (N_585,In_458,N_34);
or U586 (N_586,In_1093,N_259);
xnor U587 (N_587,N_147,In_655);
nor U588 (N_588,In_643,N_396);
nor U589 (N_589,N_314,In_965);
xnor U590 (N_590,N_31,In_490);
or U591 (N_591,N_360,In_539);
or U592 (N_592,In_366,N_302);
or U593 (N_593,In_1100,N_382);
xnor U594 (N_594,N_116,In_378);
nand U595 (N_595,In_1113,In_1193);
xor U596 (N_596,In_1114,In_772);
nand U597 (N_597,N_398,In_1141);
nor U598 (N_598,In_237,N_318);
and U599 (N_599,In_764,In_683);
nand U600 (N_600,In_1376,N_217);
and U601 (N_601,N_252,N_155);
xnor U602 (N_602,N_599,N_384);
nand U603 (N_603,In_404,N_479);
nor U604 (N_604,N_499,In_1035);
or U605 (N_605,In_470,In_48);
nand U606 (N_606,In_262,N_468);
nand U607 (N_607,In_933,N_534);
and U608 (N_608,In_468,N_229);
and U609 (N_609,In_335,In_535);
nor U610 (N_610,In_311,N_541);
nand U611 (N_611,N_20,N_475);
and U612 (N_612,N_245,In_144);
nand U613 (N_613,N_375,In_517);
xor U614 (N_614,N_438,In_1281);
or U615 (N_615,In_1427,N_454);
and U616 (N_616,In_623,In_1031);
or U617 (N_617,N_436,N_327);
xor U618 (N_618,In_484,In_1089);
or U619 (N_619,N_540,In_872);
nor U620 (N_620,N_234,In_797);
or U621 (N_621,In_716,N_105);
and U622 (N_622,In_1255,In_949);
or U623 (N_623,In_543,N_0);
xnor U624 (N_624,In_1027,In_522);
nand U625 (N_625,N_505,In_587);
and U626 (N_626,N_167,N_1);
nand U627 (N_627,In_1337,N_516);
nor U628 (N_628,N_553,N_433);
or U629 (N_629,N_287,N_282);
nand U630 (N_630,In_1137,In_652);
xor U631 (N_631,N_356,In_845);
nor U632 (N_632,In_1046,N_521);
nor U633 (N_633,N_371,N_490);
or U634 (N_634,In_891,In_1392);
nor U635 (N_635,N_7,N_82);
nor U636 (N_636,N_19,In_1163);
nand U637 (N_637,In_644,N_492);
and U638 (N_638,In_439,In_1233);
or U639 (N_639,N_65,In_1374);
nand U640 (N_640,In_1029,In_418);
and U641 (N_641,N_457,In_135);
nand U642 (N_642,In_1416,N_201);
nand U643 (N_643,In_1248,In_1170);
or U644 (N_644,In_1477,In_1383);
nand U645 (N_645,In_569,N_278);
nor U646 (N_646,N_491,In_422);
and U647 (N_647,N_23,In_938);
nor U648 (N_648,In_41,In_1389);
nor U649 (N_649,In_178,N_206);
xor U650 (N_650,In_184,In_1151);
and U651 (N_651,N_353,In_902);
and U652 (N_652,N_50,In_1294);
nand U653 (N_653,In_450,In_1419);
and U654 (N_654,In_243,N_544);
nand U655 (N_655,N_198,In_1069);
and U656 (N_656,In_1495,In_148);
nor U657 (N_657,In_337,N_526);
or U658 (N_658,N_425,N_181);
or U659 (N_659,N_269,N_416);
and U660 (N_660,N_228,In_476);
xnor U661 (N_661,N_585,In_744);
and U662 (N_662,N_91,In_619);
nor U663 (N_663,In_1264,N_49);
xnor U664 (N_664,In_926,N_280);
xor U665 (N_665,In_1104,In_1433);
and U666 (N_666,In_765,In_833);
xor U667 (N_667,In_758,N_365);
xor U668 (N_668,In_1303,N_470);
nor U669 (N_669,In_1395,N_331);
or U670 (N_670,In_898,In_502);
nor U671 (N_671,N_552,N_41);
xnor U672 (N_672,N_480,N_261);
and U673 (N_673,N_484,N_533);
nand U674 (N_674,In_1177,N_440);
nand U675 (N_675,N_33,N_81);
or U676 (N_676,In_1371,N_419);
xor U677 (N_677,In_1018,In_1462);
and U678 (N_678,In_1055,N_512);
nand U679 (N_679,In_288,In_205);
nor U680 (N_680,In_408,In_883);
xor U681 (N_681,N_243,N_430);
nand U682 (N_682,In_805,In_65);
xor U683 (N_683,N_444,In_21);
nor U684 (N_684,N_477,N_199);
xnor U685 (N_685,In_534,N_214);
xnor U686 (N_686,In_1130,In_1309);
xor U687 (N_687,N_408,In_989);
nand U688 (N_688,N_414,In_265);
or U689 (N_689,In_230,N_281);
and U690 (N_690,N_284,N_301);
nand U691 (N_691,In_1332,N_117);
nor U692 (N_692,N_79,In_298);
xor U693 (N_693,N_448,In_1072);
xnor U694 (N_694,N_570,In_939);
and U695 (N_695,In_1060,N_538);
xor U696 (N_696,N_330,N_449);
xor U697 (N_697,N_112,N_515);
or U698 (N_698,In_615,In_1499);
nand U699 (N_699,In_509,N_346);
and U700 (N_700,In_1425,N_46);
nand U701 (N_701,In_660,In_817);
xor U702 (N_702,In_1331,N_303);
xnor U703 (N_703,N_153,In_162);
nor U704 (N_704,N_258,In_1108);
or U705 (N_705,In_846,In_932);
nand U706 (N_706,In_197,In_1283);
xnor U707 (N_707,N_545,N_77);
or U708 (N_708,In_1222,In_129);
nor U709 (N_709,In_247,N_577);
nor U710 (N_710,In_225,N_417);
or U711 (N_711,In_175,In_328);
xor U712 (N_712,N_386,In_489);
nand U713 (N_713,N_400,In_672);
nand U714 (N_714,In_329,In_405);
xnor U715 (N_715,N_458,In_516);
and U716 (N_716,N_260,N_123);
or U717 (N_717,N_537,N_452);
xnor U718 (N_718,In_343,In_707);
nor U719 (N_719,N_103,N_583);
nor U720 (N_720,N_591,In_519);
nand U721 (N_721,In_1375,N_336);
and U722 (N_722,In_830,In_1364);
nand U723 (N_723,In_680,In_1024);
and U724 (N_724,N_561,N_559);
and U725 (N_725,In_684,In_854);
or U726 (N_726,N_94,In_506);
xor U727 (N_727,N_29,N_211);
nand U728 (N_728,In_1292,In_945);
and U729 (N_729,In_641,In_401);
xor U730 (N_730,N_523,N_572);
xnor U731 (N_731,In_1401,N_415);
or U732 (N_732,In_1075,N_511);
xor U733 (N_733,N_525,N_426);
or U734 (N_734,N_332,N_37);
or U735 (N_735,N_238,In_708);
nand U736 (N_736,N_131,In_821);
or U737 (N_737,N_503,N_209);
xnor U738 (N_738,In_922,N_207);
nor U739 (N_739,N_481,In_782);
xor U740 (N_740,In_978,N_580);
xor U741 (N_741,N_558,N_588);
xor U742 (N_742,N_412,In_578);
or U743 (N_743,N_548,N_569);
nor U744 (N_744,In_419,N_268);
nor U745 (N_745,In_739,N_434);
or U746 (N_746,N_483,N_93);
nand U747 (N_747,In_131,N_573);
and U748 (N_748,N_293,N_501);
nor U749 (N_749,In_1230,N_216);
nand U750 (N_750,N_292,In_563);
or U751 (N_751,In_292,In_931);
or U752 (N_752,N_514,N_439);
xor U753 (N_753,In_24,N_233);
or U754 (N_754,In_1372,N_566);
nor U755 (N_755,In_673,N_366);
nand U756 (N_756,In_1010,In_1102);
xor U757 (N_757,In_28,N_413);
and U758 (N_758,In_108,In_930);
and U759 (N_759,N_455,In_596);
and U760 (N_760,In_290,In_1409);
or U761 (N_761,N_487,In_809);
nand U762 (N_762,N_354,N_507);
xnor U763 (N_763,N_539,In_1041);
or U764 (N_764,N_461,In_943);
nand U765 (N_765,In_1487,N_130);
xor U766 (N_766,N_175,N_178);
nand U767 (N_767,In_653,In_1001);
xnor U768 (N_768,In_1088,In_380);
nand U769 (N_769,In_602,N_478);
xnor U770 (N_770,In_894,In_1334);
and U771 (N_771,N_113,N_270);
nor U772 (N_772,N_560,N_405);
nand U773 (N_773,In_494,N_48);
xnor U774 (N_774,N_96,In_1336);
or U775 (N_775,N_328,In_848);
and U776 (N_776,N_462,N_486);
xor U777 (N_777,In_1278,In_256);
or U778 (N_778,In_942,In_130);
nand U779 (N_779,N_385,N_309);
nand U780 (N_780,N_465,In_528);
nand U781 (N_781,N_14,N_556);
nor U782 (N_782,N_421,In_125);
or U783 (N_783,In_155,N_496);
and U784 (N_784,N_504,In_561);
nor U785 (N_785,N_428,In_885);
xor U786 (N_786,N_272,In_648);
or U787 (N_787,N_576,In_384);
or U788 (N_788,N_321,In_827);
xnor U789 (N_789,In_990,In_688);
nor U790 (N_790,N_13,N_476);
and U791 (N_791,In_826,In_50);
and U792 (N_792,N_409,In_763);
nor U793 (N_793,In_1202,In_51);
or U794 (N_794,N_518,In_330);
and U795 (N_795,N_565,In_475);
nor U796 (N_796,In_925,N_225);
xnor U797 (N_797,N_192,N_510);
and U798 (N_798,In_94,In_1182);
nand U799 (N_799,In_87,N_361);
and U800 (N_800,In_1228,N_362);
and U801 (N_801,N_531,N_581);
xnor U802 (N_802,In_73,N_143);
nand U803 (N_803,In_35,In_1204);
and U804 (N_804,N_669,N_745);
or U805 (N_805,N_307,N_527);
or U806 (N_806,N_720,In_1118);
nand U807 (N_807,N_784,In_444);
or U808 (N_808,In_977,N_763);
nor U809 (N_809,N_393,N_695);
nand U810 (N_810,N_219,N_634);
nand U811 (N_811,N_604,N_632);
nand U812 (N_812,In_416,N_630);
xnor U813 (N_813,N_467,In_1097);
nand U814 (N_814,N_563,N_747);
or U815 (N_815,N_72,N_246);
nand U816 (N_816,N_160,N_495);
xor U817 (N_817,In_142,N_529);
or U818 (N_818,N_692,N_752);
and U819 (N_819,N_388,In_988);
and U820 (N_820,N_394,In_1050);
or U821 (N_821,N_691,In_1234);
and U822 (N_822,N_753,In_1225);
nor U823 (N_823,In_402,N_574);
xnor U824 (N_824,N_651,N_702);
nand U825 (N_825,In_170,N_762);
and U826 (N_826,In_1435,In_618);
nor U827 (N_827,N_584,N_38);
or U828 (N_828,In_1473,N_317);
and U829 (N_829,N_26,N_686);
and U830 (N_830,N_696,N_658);
nand U831 (N_831,In_210,In_1062);
nor U832 (N_832,N_427,N_769);
or U833 (N_833,N_422,In_914);
nor U834 (N_834,N_665,In_294);
xnor U835 (N_835,N_391,N_25);
xor U836 (N_836,N_754,In_695);
nor U837 (N_837,In_164,In_283);
or U838 (N_838,In_674,In_626);
xor U839 (N_839,In_1022,In_1237);
xor U840 (N_840,N_304,In_457);
xor U841 (N_841,In_904,N_704);
and U842 (N_842,N_622,N_795);
and U843 (N_843,In_61,In_15);
nand U844 (N_844,N_646,N_567);
or U845 (N_845,N_40,In_1426);
xnor U846 (N_846,N_601,In_42);
or U847 (N_847,In_339,In_396);
xnor U848 (N_848,N_625,N_594);
nor U849 (N_849,N_325,In_610);
or U850 (N_850,In_1003,N_589);
nand U851 (N_851,N_445,In_868);
xor U852 (N_852,In_999,N_509);
nor U853 (N_853,In_373,N_737);
nand U854 (N_854,In_1186,N_662);
xnor U855 (N_855,N_343,N_497);
nand U856 (N_856,N_15,N_653);
or U857 (N_857,N_535,In_252);
and U858 (N_858,N_532,In_585);
and U859 (N_859,N_755,N_485);
nand U860 (N_860,N_749,N_299);
nor U861 (N_861,N_793,In_735);
nand U862 (N_862,In_201,N_381);
nor U863 (N_863,N_618,N_215);
xnor U864 (N_864,In_1488,N_685);
or U865 (N_865,N_739,N_786);
and U866 (N_866,In_287,N_372);
and U867 (N_867,N_376,N_190);
nor U868 (N_868,N_649,N_517);
or U869 (N_869,In_650,In_282);
xor U870 (N_870,In_1051,In_382);
xor U871 (N_871,N_613,N_639);
and U872 (N_872,N_729,In_352);
and U873 (N_873,In_423,N_760);
xnor U874 (N_874,In_1268,N_451);
or U875 (N_875,N_659,In_1468);
nand U876 (N_876,In_1056,N_628);
nor U877 (N_877,N_798,In_1155);
nand U878 (N_878,N_672,N_698);
nor U879 (N_879,N_730,N_502);
nand U880 (N_880,N_44,In_1049);
or U881 (N_881,N_557,In_229);
or U882 (N_882,In_266,N_543);
and U883 (N_883,N_602,N_474);
xor U884 (N_884,In_866,In_1127);
and U885 (N_885,N_624,In_1198);
and U886 (N_886,N_62,N_52);
and U887 (N_887,In_791,N_524);
nor U888 (N_888,In_241,N_168);
nor U889 (N_889,N_726,In_1491);
or U890 (N_890,N_667,N_690);
or U891 (N_891,In_824,N_701);
and U892 (N_892,In_188,N_593);
or U893 (N_893,N_164,In_203);
nand U894 (N_894,In_1226,N_138);
nand U895 (N_895,In_1252,N_756);
nor U896 (N_896,In_199,In_367);
and U897 (N_897,In_759,In_685);
xnor U898 (N_898,In_1214,In_975);
nor U899 (N_899,N_21,In_198);
nor U900 (N_900,In_995,In_22);
xor U901 (N_901,In_1308,N_3);
nor U902 (N_902,N_609,N_645);
xor U903 (N_903,N_231,In_1153);
or U904 (N_904,N_498,In_1028);
and U905 (N_905,N_224,In_251);
and U906 (N_906,N_766,In_921);
nand U907 (N_907,N_450,N_513);
nand U908 (N_908,N_582,N_670);
nor U909 (N_909,In_132,N_247);
or U910 (N_910,N_663,N_797);
nor U911 (N_911,N_424,N_647);
nor U912 (N_912,In_1227,N_719);
nor U913 (N_913,N_680,In_320);
nor U914 (N_914,N_447,N_420);
nand U915 (N_915,N_773,In_1112);
xnor U916 (N_916,In_1011,N_364);
nor U917 (N_917,In_351,In_1196);
nand U918 (N_918,N_137,N_682);
nor U919 (N_919,N_488,N_767);
and U920 (N_920,In_790,N_725);
nor U921 (N_921,In_1147,N_347);
nand U922 (N_922,N_118,N_664);
nand U923 (N_923,N_222,N_708);
nand U924 (N_924,In_14,N_699);
nor U925 (N_925,In_173,N_275);
nor U926 (N_926,In_1181,N_642);
nand U927 (N_927,In_1040,In_271);
and U928 (N_928,N_500,N_87);
and U929 (N_929,In_415,N_432);
and U930 (N_930,In_355,N_743);
and U931 (N_931,In_1157,In_874);
xor U932 (N_932,N_387,N_693);
xnor U933 (N_933,N_638,N_380);
xnor U934 (N_934,In_1065,N_626);
nand U935 (N_935,In_326,In_775);
or U936 (N_936,In_1415,N_466);
nand U937 (N_937,In_133,N_443);
xnor U938 (N_938,N_748,In_972);
or U939 (N_939,N_677,N_758);
nor U940 (N_940,N_42,N_734);
and U941 (N_941,In_409,N_724);
or U942 (N_942,N_578,N_740);
and U943 (N_943,N_600,In_106);
and U944 (N_944,N_310,In_559);
nor U945 (N_945,N_341,N_348);
nand U946 (N_946,In_102,N_6);
nor U947 (N_947,In_397,N_671);
and U948 (N_948,N_528,In_944);
and U949 (N_949,N_291,N_536);
and U950 (N_950,N_333,N_792);
nor U951 (N_951,N_463,In_627);
xor U952 (N_952,N_411,In_38);
or U953 (N_953,In_1378,N_768);
nor U954 (N_954,In_20,N_621);
and U955 (N_955,In_1257,In_741);
or U956 (N_956,N_435,N_431);
xnor U957 (N_957,In_518,In_332);
or U958 (N_958,N_161,In_786);
or U959 (N_959,N_772,N_456);
or U960 (N_960,N_489,In_1123);
and U961 (N_961,N_575,N_741);
and U962 (N_962,N_633,N_493);
and U963 (N_963,In_1020,N_776);
xnor U964 (N_964,N_722,N_666);
nor U965 (N_965,N_407,In_1479);
nand U966 (N_966,N_339,N_551);
nand U967 (N_967,In_647,N_678);
or U968 (N_968,In_1019,N_751);
xor U969 (N_969,In_267,N_738);
and U970 (N_970,In_1210,N_595);
or U971 (N_971,In_663,In_215);
nand U972 (N_972,N_706,N_700);
nor U973 (N_973,N_648,In_799);
nand U974 (N_974,N_453,N_564);
and U975 (N_975,In_911,In_793);
xor U976 (N_976,N_554,In_29);
and U977 (N_977,N_661,N_239);
nand U978 (N_978,N_429,In_631);
nand U979 (N_979,In_279,In_979);
xnor U980 (N_980,N_614,In_508);
and U981 (N_981,N_471,In_916);
or U982 (N_982,N_349,N_286);
and U983 (N_983,In_1323,N_17);
nor U984 (N_984,N_338,In_1189);
nand U985 (N_985,N_640,N_679);
nor U986 (N_986,N_324,N_232);
xor U987 (N_987,In_571,N_568);
xnor U988 (N_988,In_208,In_773);
nor U989 (N_989,N_342,N_636);
nand U990 (N_990,N_494,In_1324);
nand U991 (N_991,In_1411,N_592);
or U992 (N_992,In_4,N_703);
and U993 (N_993,In_1407,N_464);
xnor U994 (N_994,N_759,In_638);
nor U995 (N_995,N_709,N_70);
and U996 (N_996,N_315,N_418);
nor U997 (N_997,N_58,In_551);
nand U998 (N_998,In_1217,N_617);
or U999 (N_999,N_389,In_530);
or U1000 (N_1000,N_248,In_745);
nor U1001 (N_1001,N_660,N_923);
or U1002 (N_1002,N_654,In_689);
and U1003 (N_1003,In_553,In_1379);
nor U1004 (N_1004,N_656,In_146);
nor U1005 (N_1005,N_864,N_300);
or U1006 (N_1006,N_802,In_43);
nor U1007 (N_1007,N_482,N_996);
or U1008 (N_1008,N_955,N_236);
nand U1009 (N_1009,N_868,In_1058);
or U1010 (N_1010,In_512,N_226);
nor U1011 (N_1011,N_637,N_635);
xnor U1012 (N_1012,N_863,N_839);
nand U1013 (N_1013,N_789,In_1132);
xor U1014 (N_1014,N_266,N_98);
nor U1015 (N_1015,In_812,N_982);
xnor U1016 (N_1016,N_780,N_823);
nor U1017 (N_1017,N_611,N_984);
or U1018 (N_1018,N_893,N_810);
nor U1019 (N_1019,N_675,N_831);
nor U1020 (N_1020,N_74,In_1361);
nand U1021 (N_1021,In_1081,In_604);
nand U1022 (N_1022,N_852,N_149);
nand U1023 (N_1023,N_808,In_1397);
xnor U1024 (N_1024,N_610,N_827);
xor U1025 (N_1025,N_121,In_254);
nor U1026 (N_1026,N_937,N_986);
xnor U1027 (N_1027,N_244,N_855);
nand U1028 (N_1028,N_681,N_555);
or U1029 (N_1029,N_460,N_712);
nor U1030 (N_1030,N_803,N_520);
nor U1031 (N_1031,N_951,In_1054);
or U1032 (N_1032,N_816,In_167);
and U1033 (N_1033,In_714,In_613);
xnor U1034 (N_1034,In_749,N_794);
or U1035 (N_1035,In_1111,N_579);
nand U1036 (N_1036,N_858,N_778);
or U1037 (N_1037,N_874,In_1413);
xnor U1038 (N_1038,N_926,N_807);
xor U1039 (N_1039,N_619,In_281);
and U1040 (N_1040,N_262,N_916);
or U1041 (N_1041,N_842,N_73);
and U1042 (N_1042,In_810,N_716);
nand U1043 (N_1043,N_841,N_731);
or U1044 (N_1044,N_861,N_775);
and U1045 (N_1045,N_590,N_811);
nor U1046 (N_1046,N_826,N_975);
nor U1047 (N_1047,N_779,N_306);
or U1048 (N_1048,N_974,N_804);
or U1049 (N_1049,N_608,N_612);
xor U1050 (N_1050,In_542,N_977);
nand U1051 (N_1051,N_220,In_950);
or U1052 (N_1052,In_715,N_900);
and U1053 (N_1053,N_907,N_933);
and U1054 (N_1054,N_369,In_935);
and U1055 (N_1055,N_866,N_833);
nand U1056 (N_1056,In_992,N_673);
and U1057 (N_1057,In_56,N_814);
xor U1058 (N_1058,N_717,N_251);
nor U1059 (N_1059,In_297,In_1209);
or U1060 (N_1060,In_1079,N_606);
or U1061 (N_1061,N_586,In_487);
or U1062 (N_1062,N_329,In_1301);
nand U1063 (N_1063,N_446,N_965);
or U1064 (N_1064,N_765,N_55);
nor U1065 (N_1065,In_145,N_846);
or U1066 (N_1066,N_914,In_621);
and U1067 (N_1067,In_246,N_870);
xor U1068 (N_1068,N_943,N_924);
and U1069 (N_1069,N_983,N_918);
and U1070 (N_1070,N_825,N_472);
nand U1071 (N_1071,In_897,N_781);
xnor U1072 (N_1072,N_687,N_787);
xnor U1073 (N_1073,N_100,In_1251);
nor U1074 (N_1074,N_340,N_735);
or U1075 (N_1075,N_655,N_853);
and U1076 (N_1076,In_111,N_812);
nand U1077 (N_1077,In_636,N_857);
or U1078 (N_1078,N_607,N_727);
nor U1079 (N_1079,N_801,N_886);
nor U1080 (N_1080,N_970,N_948);
and U1081 (N_1081,In_948,In_776);
nand U1082 (N_1082,N_828,N_742);
xnor U1083 (N_1083,N_979,In_5);
xnor U1084 (N_1084,N_844,N_202);
and U1085 (N_1085,In_1023,In_1131);
or U1086 (N_1086,N_158,In_920);
xnor U1087 (N_1087,In_1288,N_834);
or U1088 (N_1088,In_1297,N_873);
or U1089 (N_1089,N_961,N_597);
or U1090 (N_1090,N_650,N_888);
or U1091 (N_1091,In_68,N_316);
and U1092 (N_1092,In_353,N_837);
or U1093 (N_1093,N_308,In_1133);
nor U1094 (N_1094,N_889,In_309);
xor U1095 (N_1095,N_973,N_962);
and U1096 (N_1096,N_995,N_830);
nor U1097 (N_1097,N_713,N_849);
or U1098 (N_1098,In_896,N_915);
and U1099 (N_1099,N_936,In_277);
nor U1100 (N_1100,N_806,N_403);
or U1101 (N_1101,N_641,In_64);
xnor U1102 (N_1102,N_944,N_999);
xor U1103 (N_1103,N_930,N_880);
nand U1104 (N_1104,In_586,N_882);
or U1105 (N_1105,N_941,N_872);
or U1106 (N_1106,N_777,N_401);
and U1107 (N_1107,N_643,N_683);
nand U1108 (N_1108,In_459,N_337);
and U1109 (N_1109,N_697,N_832);
nor U1110 (N_1110,N_733,N_242);
or U1111 (N_1111,In_927,N_334);
xor U1112 (N_1112,In_832,N_410);
or U1113 (N_1113,N_241,N_200);
and U1114 (N_1114,N_785,N_969);
and U1115 (N_1115,N_901,In_691);
nor U1116 (N_1116,N_991,N_908);
or U1117 (N_1117,N_530,N_506);
or U1118 (N_1118,In_679,N_644);
nor U1119 (N_1119,N_459,N_714);
and U1120 (N_1120,N_912,N_437);
and U1121 (N_1121,N_820,In_1178);
nand U1122 (N_1122,In_1457,N_981);
and U1123 (N_1123,N_358,N_963);
nor U1124 (N_1124,In_1346,N_821);
or U1125 (N_1125,N_843,N_101);
nand U1126 (N_1126,N_985,N_902);
xnor U1127 (N_1127,In_887,N_603);
or U1128 (N_1128,N_796,N_788);
nand U1129 (N_1129,In_913,N_684);
nand U1130 (N_1130,In_121,N_519);
nor U1131 (N_1131,In_391,N_711);
xnor U1132 (N_1132,N_953,In_55);
or U1133 (N_1133,N_657,In_884);
nor U1134 (N_1134,N_265,N_652);
nand U1135 (N_1135,N_800,In_1279);
or U1136 (N_1136,N_919,N_542);
and U1137 (N_1137,N_867,N_694);
and U1138 (N_1138,N_971,N_942);
or U1139 (N_1139,N_771,N_910);
and U1140 (N_1140,N_992,N_728);
xnor U1141 (N_1141,N_423,In_1174);
xor U1142 (N_1142,N_770,N_813);
or U1143 (N_1143,N_668,N_764);
or U1144 (N_1144,N_976,N_894);
nor U1145 (N_1145,N_550,N_587);
xor U1146 (N_1146,N_856,N_851);
and U1147 (N_1147,In_818,N_967);
and U1148 (N_1148,N_718,N_885);
nand U1149 (N_1149,N_904,N_836);
nand U1150 (N_1150,N_883,N_897);
and U1151 (N_1151,In_622,N_508);
and U1152 (N_1152,N_895,N_674);
nor U1153 (N_1153,N_954,N_898);
and U1154 (N_1154,In_654,In_379);
and U1155 (N_1155,N_998,N_615);
nor U1156 (N_1156,N_546,In_291);
xor U1157 (N_1157,In_899,In_1101);
xnor U1158 (N_1158,N_989,N_783);
nor U1159 (N_1159,N_978,N_896);
nor U1160 (N_1160,In_119,N_473);
and U1161 (N_1161,N_881,In_1455);
nor U1162 (N_1162,In_1183,In_662);
nor U1163 (N_1163,N_790,N_913);
nor U1164 (N_1164,N_63,N_791);
and U1165 (N_1165,N_406,N_817);
or U1166 (N_1166,N_847,N_819);
xor U1167 (N_1167,In_1400,N_441);
and U1168 (N_1168,N_799,N_549);
nand U1169 (N_1169,N_917,N_736);
or U1170 (N_1170,In_347,N_929);
nor U1171 (N_1171,N_289,N_903);
nor U1172 (N_1172,N_865,N_877);
or U1173 (N_1173,N_899,N_835);
nand U1174 (N_1174,N_871,N_934);
nor U1175 (N_1175,N_988,N_878);
nor U1176 (N_1176,N_442,In_611);
and U1177 (N_1177,In_249,N_212);
nor U1178 (N_1178,In_443,N_547);
or U1179 (N_1179,In_877,N_469);
or U1180 (N_1180,N_715,N_627);
or U1181 (N_1181,N_822,N_320);
xnor U1182 (N_1182,N_688,N_957);
nor U1183 (N_1183,N_757,N_744);
and U1184 (N_1184,N_598,N_938);
or U1185 (N_1185,N_402,In_1150);
or U1186 (N_1186,N_939,N_838);
or U1187 (N_1187,N_921,N_805);
nor U1188 (N_1188,In_934,N_676);
nand U1189 (N_1189,N_905,In_1492);
and U1190 (N_1190,N_721,N_949);
nor U1191 (N_1191,N_940,N_352);
nand U1192 (N_1192,N_854,N_404);
nor U1193 (N_1193,N_884,N_968);
nor U1194 (N_1194,In_720,N_850);
nand U1195 (N_1195,In_969,N_840);
and U1196 (N_1196,N_928,In_1434);
xor U1197 (N_1197,N_887,N_997);
and U1198 (N_1198,In_420,N_750);
xor U1199 (N_1199,In_769,N_922);
and U1200 (N_1200,N_876,N_1024);
nand U1201 (N_1201,N_1082,N_1045);
xor U1202 (N_1202,N_1153,N_1081);
or U1203 (N_1203,N_1184,N_1112);
xor U1204 (N_1204,N_1018,N_705);
nand U1205 (N_1205,N_1102,N_1098);
or U1206 (N_1206,N_1079,N_1154);
nor U1207 (N_1207,N_890,N_932);
xor U1208 (N_1208,N_707,N_732);
xor U1209 (N_1209,N_1030,N_203);
xnor U1210 (N_1210,N_1063,N_1186);
and U1211 (N_1211,N_1100,N_1025);
nor U1212 (N_1212,N_1016,In_756);
or U1213 (N_1213,N_1124,N_1065);
and U1214 (N_1214,N_1048,In_1394);
nand U1215 (N_1215,N_1116,N_875);
and U1216 (N_1216,N_1057,In_666);
and U1217 (N_1217,N_1068,N_1128);
xnor U1218 (N_1218,N_1069,N_1193);
xor U1219 (N_1219,N_879,N_1113);
nand U1220 (N_1220,N_946,N_761);
or U1221 (N_1221,N_1046,N_1143);
nor U1222 (N_1222,N_1076,N_1126);
and U1223 (N_1223,N_1041,N_972);
xor U1224 (N_1224,N_1004,N_935);
xor U1225 (N_1225,In_134,N_1189);
and U1226 (N_1226,N_945,N_862);
nand U1227 (N_1227,N_1157,N_1129);
and U1228 (N_1228,N_596,N_950);
and U1229 (N_1229,N_1177,N_562);
nor U1230 (N_1230,In_733,N_1091);
and U1231 (N_1231,N_1147,N_1134);
nand U1232 (N_1232,N_809,N_631);
nor U1233 (N_1233,N_1096,In_671);
xnor U1234 (N_1234,N_1115,N_774);
and U1235 (N_1235,N_1121,N_1094);
nor U1236 (N_1236,N_1031,N_860);
xor U1237 (N_1237,In_187,N_605);
nor U1238 (N_1238,N_1060,N_1103);
or U1239 (N_1239,N_1095,N_1051);
or U1240 (N_1240,N_1119,N_1117);
xor U1241 (N_1241,N_1067,N_1050);
or U1242 (N_1242,N_1196,N_1118);
xnor U1243 (N_1243,N_1135,N_1173);
nor U1244 (N_1244,N_1192,N_1174);
xor U1245 (N_1245,N_1123,N_1182);
and U1246 (N_1246,N_1088,N_1009);
or U1247 (N_1247,N_1053,N_1062);
nand U1248 (N_1248,N_1089,In_725);
or U1249 (N_1249,N_522,N_1092);
nor U1250 (N_1250,N_1052,N_1183);
nor U1251 (N_1251,N_1109,N_723);
and U1252 (N_1252,N_1175,N_1132);
or U1253 (N_1253,N_1035,N_1167);
xnor U1254 (N_1254,N_1071,N_947);
or U1255 (N_1255,N_290,N_571);
and U1256 (N_1256,N_1011,N_1191);
or U1257 (N_1257,In_344,N_1038);
nand U1258 (N_1258,N_1101,N_958);
and U1259 (N_1259,N_920,N_1197);
nand U1260 (N_1260,In_357,N_1137);
or U1261 (N_1261,N_1074,N_1003);
nand U1262 (N_1262,N_1107,In_1343);
nand U1263 (N_1263,N_1164,N_960);
xnor U1264 (N_1264,In_425,N_1006);
nor U1265 (N_1265,N_1012,N_909);
nand U1266 (N_1266,In_1105,N_1169);
xnor U1267 (N_1267,N_980,N_1055);
nand U1268 (N_1268,N_1156,N_1138);
nor U1269 (N_1269,N_1015,N_294);
nand U1270 (N_1270,N_1127,In_1017);
nand U1271 (N_1271,N_1054,N_1176);
nand U1272 (N_1272,N_1028,In_659);
xor U1273 (N_1273,N_1066,N_1021);
or U1274 (N_1274,N_1111,N_1140);
and U1275 (N_1275,N_1078,In_860);
nor U1276 (N_1276,N_891,N_1027);
or U1277 (N_1277,N_1144,N_1032);
nor U1278 (N_1278,N_1000,N_1077);
xnor U1279 (N_1279,N_180,In_461);
and U1280 (N_1280,N_1148,N_990);
nor U1281 (N_1281,N_1160,N_1120);
and U1282 (N_1282,N_1141,In_1385);
or U1283 (N_1283,N_1014,N_1190);
nand U1284 (N_1284,N_1086,In_731);
nor U1285 (N_1285,N_1149,N_959);
and U1286 (N_1286,N_1162,N_623);
nand U1287 (N_1287,N_629,N_1151);
and U1288 (N_1288,N_746,N_815);
or U1289 (N_1289,N_1161,N_1179);
and U1290 (N_1290,N_1036,In_60);
or U1291 (N_1291,N_994,N_1072);
nand U1292 (N_1292,N_1010,N_1170);
or U1293 (N_1293,N_1125,N_964);
nand U1294 (N_1294,N_1007,N_1108);
nor U1295 (N_1295,N_1020,N_80);
nor U1296 (N_1296,N_1029,N_782);
xor U1297 (N_1297,N_196,In_747);
or U1298 (N_1298,N_1145,N_987);
and U1299 (N_1299,N_1188,N_1155);
and U1300 (N_1300,N_1139,N_1181);
nor U1301 (N_1301,N_818,N_1194);
nor U1302 (N_1302,N_925,N_1087);
nand U1303 (N_1303,In_1265,N_1198);
nor U1304 (N_1304,N_1013,N_1142);
nor U1305 (N_1305,N_927,N_1185);
or U1306 (N_1306,N_1168,N_1075);
or U1307 (N_1307,N_1008,N_1093);
or U1308 (N_1308,N_1039,N_1114);
or U1309 (N_1309,N_1084,N_1083);
nor U1310 (N_1310,N_1002,N_1059);
nor U1311 (N_1311,N_1049,N_1023);
nand U1312 (N_1312,N_1099,N_993);
nand U1313 (N_1313,N_931,N_1104);
xnor U1314 (N_1314,N_276,In_219);
or U1315 (N_1315,N_227,N_1005);
nor U1316 (N_1316,N_1165,N_1073);
and U1317 (N_1317,N_1034,N_1105);
nand U1318 (N_1318,N_1178,N_1056);
nor U1319 (N_1319,N_1131,N_1033);
or U1320 (N_1320,N_1150,N_1159);
and U1321 (N_1321,N_859,N_1042);
nand U1322 (N_1322,N_1152,In_766);
nor U1323 (N_1323,N_1058,In_724);
or U1324 (N_1324,N_1085,N_1136);
nor U1325 (N_1325,N_1061,N_1130);
nand U1326 (N_1326,N_1026,N_1195);
or U1327 (N_1327,In_537,N_1080);
nand U1328 (N_1328,N_869,N_616);
or U1329 (N_1329,N_1187,N_1106);
nand U1330 (N_1330,In_538,N_1047);
nand U1331 (N_1331,N_845,N_1022);
and U1332 (N_1332,N_911,N_1090);
nor U1333 (N_1333,N_1070,N_1163);
or U1334 (N_1334,N_1199,N_1146);
and U1335 (N_1335,N_966,N_1110);
xnor U1336 (N_1336,N_892,N_1043);
nand U1337 (N_1337,N_1064,N_1040);
and U1338 (N_1338,N_848,N_824);
xor U1339 (N_1339,N_1037,N_689);
nor U1340 (N_1340,N_1019,N_906);
or U1341 (N_1341,N_1133,N_1180);
xnor U1342 (N_1342,N_710,N_1001);
or U1343 (N_1343,N_1172,N_956);
and U1344 (N_1344,N_829,N_1158);
and U1345 (N_1345,N_1171,N_1122);
or U1346 (N_1346,In_603,N_296);
nor U1347 (N_1347,N_1166,N_620);
nand U1348 (N_1348,N_952,N_1097);
or U1349 (N_1349,N_1044,N_1017);
and U1350 (N_1350,N_1073,N_290);
xor U1351 (N_1351,N_1140,N_1036);
or U1352 (N_1352,N_1091,N_1076);
nor U1353 (N_1353,N_1145,N_1175);
or U1354 (N_1354,N_1017,N_1011);
nor U1355 (N_1355,N_1198,N_1070);
xnor U1356 (N_1356,N_809,N_1105);
nand U1357 (N_1357,N_959,N_1162);
and U1358 (N_1358,N_1137,N_1065);
nand U1359 (N_1359,N_1182,N_925);
xor U1360 (N_1360,N_993,N_1025);
and U1361 (N_1361,N_1115,N_180);
nor U1362 (N_1362,N_227,N_966);
or U1363 (N_1363,N_203,N_616);
xnor U1364 (N_1364,N_1040,N_562);
nand U1365 (N_1365,N_1108,N_1166);
nor U1366 (N_1366,N_1118,N_1182);
xor U1367 (N_1367,N_723,N_1137);
xnor U1368 (N_1368,N_710,N_1063);
xor U1369 (N_1369,N_987,N_956);
nor U1370 (N_1370,N_869,N_1009);
and U1371 (N_1371,N_1116,N_869);
or U1372 (N_1372,N_1033,N_1165);
nor U1373 (N_1373,N_1015,N_1095);
or U1374 (N_1374,In_60,N_1140);
or U1375 (N_1375,N_1144,N_1154);
and U1376 (N_1376,N_875,N_1015);
and U1377 (N_1377,N_809,N_1137);
and U1378 (N_1378,N_1184,N_1102);
and U1379 (N_1379,N_1118,N_1105);
xnor U1380 (N_1380,In_860,N_1024);
nor U1381 (N_1381,N_1173,N_1191);
and U1382 (N_1382,N_1164,N_227);
xnor U1383 (N_1383,N_1100,N_605);
nor U1384 (N_1384,N_1098,N_1190);
and U1385 (N_1385,N_1046,N_1097);
nand U1386 (N_1386,N_1034,N_1061);
xor U1387 (N_1387,N_1105,N_1079);
xnor U1388 (N_1388,N_596,N_1041);
or U1389 (N_1389,N_1120,N_946);
or U1390 (N_1390,N_1032,N_927);
xnor U1391 (N_1391,N_1112,N_1033);
nand U1392 (N_1392,N_1098,N_927);
and U1393 (N_1393,N_203,N_1128);
nor U1394 (N_1394,N_1106,N_990);
nor U1395 (N_1395,N_1163,N_1196);
nand U1396 (N_1396,N_1094,N_1031);
and U1397 (N_1397,N_1027,N_1112);
nor U1398 (N_1398,N_909,N_1180);
and U1399 (N_1399,In_425,N_1020);
or U1400 (N_1400,N_1391,N_1201);
or U1401 (N_1401,N_1350,N_1203);
xnor U1402 (N_1402,N_1340,N_1262);
xor U1403 (N_1403,N_1363,N_1247);
xor U1404 (N_1404,N_1343,N_1230);
or U1405 (N_1405,N_1258,N_1301);
nand U1406 (N_1406,N_1377,N_1282);
and U1407 (N_1407,N_1234,N_1392);
xnor U1408 (N_1408,N_1228,N_1227);
and U1409 (N_1409,N_1214,N_1366);
or U1410 (N_1410,N_1263,N_1371);
xor U1411 (N_1411,N_1370,N_1211);
xor U1412 (N_1412,N_1267,N_1202);
nor U1413 (N_1413,N_1305,N_1288);
xnor U1414 (N_1414,N_1224,N_1272);
xor U1415 (N_1415,N_1240,N_1386);
xor U1416 (N_1416,N_1244,N_1246);
and U1417 (N_1417,N_1342,N_1241);
nor U1418 (N_1418,N_1395,N_1261);
nand U1419 (N_1419,N_1379,N_1330);
and U1420 (N_1420,N_1205,N_1212);
nor U1421 (N_1421,N_1354,N_1289);
xor U1422 (N_1422,N_1285,N_1281);
nor U1423 (N_1423,N_1245,N_1249);
nor U1424 (N_1424,N_1336,N_1315);
or U1425 (N_1425,N_1274,N_1307);
and U1426 (N_1426,N_1259,N_1280);
xor U1427 (N_1427,N_1368,N_1365);
xnor U1428 (N_1428,N_1236,N_1328);
or U1429 (N_1429,N_1303,N_1251);
xnor U1430 (N_1430,N_1399,N_1325);
nand U1431 (N_1431,N_1313,N_1253);
and U1432 (N_1432,N_1300,N_1364);
or U1433 (N_1433,N_1398,N_1252);
nand U1434 (N_1434,N_1321,N_1260);
or U1435 (N_1435,N_1271,N_1359);
or U1436 (N_1436,N_1352,N_1332);
and U1437 (N_1437,N_1299,N_1273);
or U1438 (N_1438,N_1226,N_1223);
nor U1439 (N_1439,N_1238,N_1266);
nor U1440 (N_1440,N_1269,N_1207);
nand U1441 (N_1441,N_1292,N_1242);
nand U1442 (N_1442,N_1312,N_1200);
xnor U1443 (N_1443,N_1298,N_1372);
nand U1444 (N_1444,N_1382,N_1277);
and U1445 (N_1445,N_1326,N_1233);
nand U1446 (N_1446,N_1361,N_1357);
nand U1447 (N_1447,N_1302,N_1380);
and U1448 (N_1448,N_1390,N_1378);
nor U1449 (N_1449,N_1351,N_1250);
and U1450 (N_1450,N_1206,N_1295);
xnor U1451 (N_1451,N_1221,N_1344);
nand U1452 (N_1452,N_1338,N_1243);
nand U1453 (N_1453,N_1225,N_1358);
nand U1454 (N_1454,N_1264,N_1347);
or U1455 (N_1455,N_1323,N_1385);
nand U1456 (N_1456,N_1255,N_1345);
and U1457 (N_1457,N_1256,N_1387);
xnor U1458 (N_1458,N_1217,N_1215);
or U1459 (N_1459,N_1346,N_1283);
or U1460 (N_1460,N_1373,N_1209);
nor U1461 (N_1461,N_1254,N_1375);
or U1462 (N_1462,N_1213,N_1320);
nand U1463 (N_1463,N_1389,N_1396);
and U1464 (N_1464,N_1334,N_1327);
nor U1465 (N_1465,N_1367,N_1308);
and U1466 (N_1466,N_1268,N_1329);
or U1467 (N_1467,N_1237,N_1270);
nor U1468 (N_1468,N_1296,N_1388);
and U1469 (N_1469,N_1314,N_1278);
or U1470 (N_1470,N_1293,N_1349);
nand U1471 (N_1471,N_1204,N_1331);
nor U1472 (N_1472,N_1291,N_1222);
and U1473 (N_1473,N_1231,N_1290);
nand U1474 (N_1474,N_1265,N_1341);
nand U1475 (N_1475,N_1257,N_1279);
nand U1476 (N_1476,N_1319,N_1287);
nor U1477 (N_1477,N_1232,N_1369);
or U1478 (N_1478,N_1208,N_1318);
and U1479 (N_1479,N_1309,N_1284);
and U1480 (N_1480,N_1333,N_1220);
nor U1481 (N_1481,N_1337,N_1376);
or U1482 (N_1482,N_1239,N_1297);
or U1483 (N_1483,N_1384,N_1383);
nor U1484 (N_1484,N_1335,N_1355);
or U1485 (N_1485,N_1276,N_1294);
nand U1486 (N_1486,N_1304,N_1394);
and U1487 (N_1487,N_1229,N_1216);
xnor U1488 (N_1488,N_1322,N_1374);
or U1489 (N_1489,N_1353,N_1362);
and U1490 (N_1490,N_1348,N_1210);
or U1491 (N_1491,N_1324,N_1397);
nor U1492 (N_1492,N_1219,N_1235);
or U1493 (N_1493,N_1316,N_1393);
or U1494 (N_1494,N_1356,N_1310);
xnor U1495 (N_1495,N_1360,N_1218);
nor U1496 (N_1496,N_1317,N_1381);
xor U1497 (N_1497,N_1286,N_1275);
xnor U1498 (N_1498,N_1311,N_1248);
and U1499 (N_1499,N_1306,N_1339);
xor U1500 (N_1500,N_1393,N_1326);
or U1501 (N_1501,N_1342,N_1286);
nor U1502 (N_1502,N_1398,N_1271);
and U1503 (N_1503,N_1280,N_1309);
nand U1504 (N_1504,N_1252,N_1374);
nand U1505 (N_1505,N_1310,N_1297);
xor U1506 (N_1506,N_1350,N_1219);
nor U1507 (N_1507,N_1303,N_1372);
nor U1508 (N_1508,N_1384,N_1262);
nor U1509 (N_1509,N_1309,N_1354);
nor U1510 (N_1510,N_1367,N_1286);
nor U1511 (N_1511,N_1242,N_1328);
nand U1512 (N_1512,N_1340,N_1258);
or U1513 (N_1513,N_1270,N_1311);
nand U1514 (N_1514,N_1285,N_1303);
and U1515 (N_1515,N_1217,N_1213);
and U1516 (N_1516,N_1259,N_1217);
and U1517 (N_1517,N_1327,N_1206);
xnor U1518 (N_1518,N_1274,N_1215);
nand U1519 (N_1519,N_1280,N_1240);
nand U1520 (N_1520,N_1211,N_1338);
xnor U1521 (N_1521,N_1293,N_1220);
nor U1522 (N_1522,N_1337,N_1236);
nor U1523 (N_1523,N_1249,N_1256);
xor U1524 (N_1524,N_1320,N_1383);
nor U1525 (N_1525,N_1354,N_1270);
nor U1526 (N_1526,N_1307,N_1383);
nor U1527 (N_1527,N_1294,N_1242);
or U1528 (N_1528,N_1313,N_1222);
nor U1529 (N_1529,N_1268,N_1367);
or U1530 (N_1530,N_1356,N_1339);
or U1531 (N_1531,N_1203,N_1364);
xor U1532 (N_1532,N_1377,N_1300);
or U1533 (N_1533,N_1214,N_1240);
nand U1534 (N_1534,N_1228,N_1262);
or U1535 (N_1535,N_1219,N_1289);
xnor U1536 (N_1536,N_1398,N_1257);
nor U1537 (N_1537,N_1357,N_1355);
nand U1538 (N_1538,N_1343,N_1329);
or U1539 (N_1539,N_1229,N_1384);
or U1540 (N_1540,N_1355,N_1270);
nand U1541 (N_1541,N_1257,N_1387);
xor U1542 (N_1542,N_1374,N_1223);
or U1543 (N_1543,N_1233,N_1358);
xnor U1544 (N_1544,N_1351,N_1296);
and U1545 (N_1545,N_1333,N_1347);
nand U1546 (N_1546,N_1207,N_1376);
and U1547 (N_1547,N_1364,N_1378);
or U1548 (N_1548,N_1266,N_1321);
and U1549 (N_1549,N_1217,N_1389);
xor U1550 (N_1550,N_1314,N_1327);
nand U1551 (N_1551,N_1230,N_1268);
and U1552 (N_1552,N_1211,N_1368);
or U1553 (N_1553,N_1369,N_1389);
and U1554 (N_1554,N_1275,N_1365);
or U1555 (N_1555,N_1348,N_1369);
nor U1556 (N_1556,N_1370,N_1355);
and U1557 (N_1557,N_1388,N_1292);
nor U1558 (N_1558,N_1332,N_1308);
nand U1559 (N_1559,N_1296,N_1349);
or U1560 (N_1560,N_1340,N_1220);
nor U1561 (N_1561,N_1350,N_1254);
or U1562 (N_1562,N_1394,N_1219);
nor U1563 (N_1563,N_1282,N_1341);
nand U1564 (N_1564,N_1217,N_1398);
nand U1565 (N_1565,N_1212,N_1333);
or U1566 (N_1566,N_1311,N_1380);
and U1567 (N_1567,N_1234,N_1219);
nand U1568 (N_1568,N_1291,N_1391);
nor U1569 (N_1569,N_1349,N_1255);
xnor U1570 (N_1570,N_1384,N_1343);
and U1571 (N_1571,N_1349,N_1260);
nor U1572 (N_1572,N_1351,N_1207);
xor U1573 (N_1573,N_1209,N_1277);
nor U1574 (N_1574,N_1271,N_1308);
nor U1575 (N_1575,N_1366,N_1254);
or U1576 (N_1576,N_1277,N_1398);
and U1577 (N_1577,N_1368,N_1280);
and U1578 (N_1578,N_1217,N_1378);
and U1579 (N_1579,N_1303,N_1219);
xnor U1580 (N_1580,N_1279,N_1377);
nand U1581 (N_1581,N_1391,N_1304);
nor U1582 (N_1582,N_1368,N_1268);
or U1583 (N_1583,N_1269,N_1210);
xor U1584 (N_1584,N_1303,N_1393);
and U1585 (N_1585,N_1336,N_1327);
xnor U1586 (N_1586,N_1364,N_1338);
or U1587 (N_1587,N_1355,N_1393);
nand U1588 (N_1588,N_1293,N_1208);
and U1589 (N_1589,N_1342,N_1393);
nand U1590 (N_1590,N_1360,N_1213);
or U1591 (N_1591,N_1346,N_1354);
nand U1592 (N_1592,N_1289,N_1210);
nand U1593 (N_1593,N_1317,N_1351);
and U1594 (N_1594,N_1288,N_1281);
nor U1595 (N_1595,N_1293,N_1249);
nand U1596 (N_1596,N_1293,N_1355);
and U1597 (N_1597,N_1312,N_1247);
nand U1598 (N_1598,N_1358,N_1374);
or U1599 (N_1599,N_1350,N_1289);
nor U1600 (N_1600,N_1523,N_1544);
nor U1601 (N_1601,N_1541,N_1542);
or U1602 (N_1602,N_1483,N_1598);
or U1603 (N_1603,N_1529,N_1486);
or U1604 (N_1604,N_1467,N_1569);
and U1605 (N_1605,N_1531,N_1427);
xnor U1606 (N_1606,N_1548,N_1402);
and U1607 (N_1607,N_1491,N_1468);
or U1608 (N_1608,N_1530,N_1521);
nor U1609 (N_1609,N_1574,N_1538);
nand U1610 (N_1610,N_1442,N_1484);
and U1611 (N_1611,N_1553,N_1487);
nand U1612 (N_1612,N_1511,N_1455);
or U1613 (N_1613,N_1572,N_1517);
and U1614 (N_1614,N_1459,N_1573);
or U1615 (N_1615,N_1524,N_1565);
nand U1616 (N_1616,N_1460,N_1522);
xnor U1617 (N_1617,N_1528,N_1532);
xnor U1618 (N_1618,N_1571,N_1587);
nor U1619 (N_1619,N_1453,N_1477);
nor U1620 (N_1620,N_1594,N_1401);
and U1621 (N_1621,N_1406,N_1450);
or U1622 (N_1622,N_1443,N_1447);
or U1623 (N_1623,N_1539,N_1449);
xnor U1624 (N_1624,N_1514,N_1446);
xnor U1625 (N_1625,N_1589,N_1556);
and U1626 (N_1626,N_1465,N_1474);
and U1627 (N_1627,N_1489,N_1520);
and U1628 (N_1628,N_1502,N_1441);
nand U1629 (N_1629,N_1577,N_1552);
nor U1630 (N_1630,N_1567,N_1500);
or U1631 (N_1631,N_1526,N_1448);
nand U1632 (N_1632,N_1464,N_1423);
nor U1633 (N_1633,N_1504,N_1417);
nand U1634 (N_1634,N_1457,N_1512);
and U1635 (N_1635,N_1576,N_1579);
nand U1636 (N_1636,N_1431,N_1463);
nor U1637 (N_1637,N_1534,N_1586);
xnor U1638 (N_1638,N_1439,N_1596);
or U1639 (N_1639,N_1429,N_1516);
xnor U1640 (N_1640,N_1518,N_1543);
or U1641 (N_1641,N_1503,N_1490);
xor U1642 (N_1642,N_1471,N_1478);
nor U1643 (N_1643,N_1461,N_1582);
nand U1644 (N_1644,N_1481,N_1599);
nand U1645 (N_1645,N_1412,N_1563);
or U1646 (N_1646,N_1585,N_1506);
nor U1647 (N_1647,N_1421,N_1454);
nor U1648 (N_1648,N_1566,N_1422);
and U1649 (N_1649,N_1554,N_1400);
nand U1650 (N_1650,N_1475,N_1426);
and U1651 (N_1651,N_1535,N_1456);
xor U1652 (N_1652,N_1445,N_1411);
and U1653 (N_1653,N_1409,N_1434);
nand U1654 (N_1654,N_1419,N_1525);
nand U1655 (N_1655,N_1547,N_1536);
xnor U1656 (N_1656,N_1597,N_1537);
nor U1657 (N_1657,N_1432,N_1558);
or U1658 (N_1658,N_1591,N_1405);
and U1659 (N_1659,N_1435,N_1515);
and U1660 (N_1660,N_1404,N_1451);
xor U1661 (N_1661,N_1430,N_1551);
or U1662 (N_1662,N_1458,N_1414);
and U1663 (N_1663,N_1595,N_1438);
and U1664 (N_1664,N_1428,N_1424);
nand U1665 (N_1665,N_1472,N_1513);
nor U1666 (N_1666,N_1416,N_1479);
xnor U1667 (N_1667,N_1496,N_1470);
and U1668 (N_1668,N_1540,N_1592);
nand U1669 (N_1669,N_1546,N_1498);
and U1670 (N_1670,N_1418,N_1407);
and U1671 (N_1671,N_1462,N_1420);
xor U1672 (N_1672,N_1501,N_1482);
or U1673 (N_1673,N_1452,N_1555);
and U1674 (N_1674,N_1561,N_1485);
and U1675 (N_1675,N_1578,N_1497);
nand U1676 (N_1676,N_1593,N_1510);
or U1677 (N_1677,N_1410,N_1469);
xor U1678 (N_1678,N_1568,N_1492);
or U1679 (N_1679,N_1473,N_1527);
or U1680 (N_1680,N_1583,N_1476);
xor U1681 (N_1681,N_1557,N_1564);
xnor U1682 (N_1682,N_1425,N_1507);
or U1683 (N_1683,N_1570,N_1588);
xnor U1684 (N_1684,N_1575,N_1444);
or U1685 (N_1685,N_1580,N_1562);
xor U1686 (N_1686,N_1590,N_1509);
nand U1687 (N_1687,N_1440,N_1550);
or U1688 (N_1688,N_1494,N_1415);
xnor U1689 (N_1689,N_1437,N_1549);
and U1690 (N_1690,N_1560,N_1505);
or U1691 (N_1691,N_1436,N_1466);
nor U1692 (N_1692,N_1495,N_1559);
nand U1693 (N_1693,N_1584,N_1519);
or U1694 (N_1694,N_1581,N_1499);
or U1695 (N_1695,N_1413,N_1493);
and U1696 (N_1696,N_1533,N_1488);
xor U1697 (N_1697,N_1508,N_1433);
xor U1698 (N_1698,N_1545,N_1403);
nand U1699 (N_1699,N_1408,N_1480);
xor U1700 (N_1700,N_1495,N_1537);
and U1701 (N_1701,N_1527,N_1515);
and U1702 (N_1702,N_1410,N_1505);
and U1703 (N_1703,N_1472,N_1406);
nor U1704 (N_1704,N_1438,N_1522);
nor U1705 (N_1705,N_1596,N_1577);
or U1706 (N_1706,N_1570,N_1410);
nand U1707 (N_1707,N_1553,N_1555);
nor U1708 (N_1708,N_1477,N_1591);
and U1709 (N_1709,N_1500,N_1409);
nand U1710 (N_1710,N_1406,N_1489);
xor U1711 (N_1711,N_1573,N_1401);
and U1712 (N_1712,N_1474,N_1549);
xnor U1713 (N_1713,N_1459,N_1590);
nand U1714 (N_1714,N_1463,N_1486);
or U1715 (N_1715,N_1428,N_1495);
or U1716 (N_1716,N_1501,N_1504);
nand U1717 (N_1717,N_1421,N_1478);
xor U1718 (N_1718,N_1422,N_1486);
xnor U1719 (N_1719,N_1423,N_1425);
nand U1720 (N_1720,N_1457,N_1434);
or U1721 (N_1721,N_1436,N_1420);
and U1722 (N_1722,N_1595,N_1588);
or U1723 (N_1723,N_1564,N_1541);
or U1724 (N_1724,N_1597,N_1535);
or U1725 (N_1725,N_1519,N_1483);
nor U1726 (N_1726,N_1450,N_1508);
and U1727 (N_1727,N_1483,N_1482);
nand U1728 (N_1728,N_1492,N_1489);
nor U1729 (N_1729,N_1527,N_1506);
nor U1730 (N_1730,N_1589,N_1430);
xor U1731 (N_1731,N_1427,N_1566);
nand U1732 (N_1732,N_1480,N_1593);
or U1733 (N_1733,N_1415,N_1543);
and U1734 (N_1734,N_1516,N_1495);
nand U1735 (N_1735,N_1422,N_1473);
nor U1736 (N_1736,N_1532,N_1455);
xor U1737 (N_1737,N_1425,N_1430);
nor U1738 (N_1738,N_1573,N_1591);
nor U1739 (N_1739,N_1547,N_1523);
nand U1740 (N_1740,N_1526,N_1576);
and U1741 (N_1741,N_1403,N_1430);
nand U1742 (N_1742,N_1439,N_1564);
xor U1743 (N_1743,N_1421,N_1587);
xor U1744 (N_1744,N_1457,N_1502);
and U1745 (N_1745,N_1488,N_1431);
or U1746 (N_1746,N_1549,N_1571);
or U1747 (N_1747,N_1533,N_1431);
xnor U1748 (N_1748,N_1408,N_1429);
nor U1749 (N_1749,N_1571,N_1432);
nand U1750 (N_1750,N_1503,N_1451);
xor U1751 (N_1751,N_1577,N_1491);
nand U1752 (N_1752,N_1400,N_1538);
and U1753 (N_1753,N_1597,N_1551);
nor U1754 (N_1754,N_1572,N_1494);
nand U1755 (N_1755,N_1456,N_1421);
and U1756 (N_1756,N_1427,N_1568);
xor U1757 (N_1757,N_1552,N_1406);
and U1758 (N_1758,N_1474,N_1528);
xor U1759 (N_1759,N_1422,N_1479);
nor U1760 (N_1760,N_1574,N_1429);
or U1761 (N_1761,N_1424,N_1422);
nor U1762 (N_1762,N_1434,N_1469);
nor U1763 (N_1763,N_1422,N_1560);
or U1764 (N_1764,N_1557,N_1437);
xnor U1765 (N_1765,N_1534,N_1530);
or U1766 (N_1766,N_1401,N_1466);
or U1767 (N_1767,N_1454,N_1541);
and U1768 (N_1768,N_1525,N_1458);
nand U1769 (N_1769,N_1522,N_1598);
or U1770 (N_1770,N_1591,N_1434);
or U1771 (N_1771,N_1506,N_1517);
and U1772 (N_1772,N_1428,N_1555);
xnor U1773 (N_1773,N_1588,N_1479);
xor U1774 (N_1774,N_1435,N_1580);
or U1775 (N_1775,N_1444,N_1404);
or U1776 (N_1776,N_1446,N_1411);
nand U1777 (N_1777,N_1554,N_1587);
and U1778 (N_1778,N_1597,N_1447);
nor U1779 (N_1779,N_1534,N_1471);
nor U1780 (N_1780,N_1586,N_1541);
nor U1781 (N_1781,N_1518,N_1583);
nor U1782 (N_1782,N_1586,N_1558);
or U1783 (N_1783,N_1551,N_1439);
and U1784 (N_1784,N_1486,N_1541);
or U1785 (N_1785,N_1511,N_1439);
nand U1786 (N_1786,N_1445,N_1580);
or U1787 (N_1787,N_1511,N_1555);
and U1788 (N_1788,N_1403,N_1408);
xnor U1789 (N_1789,N_1456,N_1404);
or U1790 (N_1790,N_1506,N_1450);
nand U1791 (N_1791,N_1569,N_1590);
and U1792 (N_1792,N_1417,N_1409);
or U1793 (N_1793,N_1411,N_1578);
nor U1794 (N_1794,N_1599,N_1514);
nand U1795 (N_1795,N_1561,N_1576);
nor U1796 (N_1796,N_1417,N_1588);
and U1797 (N_1797,N_1589,N_1453);
nand U1798 (N_1798,N_1572,N_1406);
and U1799 (N_1799,N_1541,N_1538);
nor U1800 (N_1800,N_1694,N_1726);
and U1801 (N_1801,N_1670,N_1771);
or U1802 (N_1802,N_1776,N_1699);
nor U1803 (N_1803,N_1713,N_1666);
and U1804 (N_1804,N_1782,N_1787);
and U1805 (N_1805,N_1673,N_1675);
or U1806 (N_1806,N_1778,N_1646);
and U1807 (N_1807,N_1630,N_1679);
or U1808 (N_1808,N_1743,N_1680);
or U1809 (N_1809,N_1768,N_1634);
and U1810 (N_1810,N_1729,N_1616);
nand U1811 (N_1811,N_1732,N_1775);
and U1812 (N_1812,N_1760,N_1796);
xnor U1813 (N_1813,N_1629,N_1637);
xor U1814 (N_1814,N_1657,N_1693);
and U1815 (N_1815,N_1665,N_1749);
or U1816 (N_1816,N_1691,N_1725);
xor U1817 (N_1817,N_1790,N_1604);
xor U1818 (N_1818,N_1617,N_1669);
xnor U1819 (N_1819,N_1692,N_1689);
xor U1820 (N_1820,N_1767,N_1783);
or U1821 (N_1821,N_1607,N_1747);
nand U1822 (N_1822,N_1758,N_1764);
or U1823 (N_1823,N_1660,N_1626);
and U1824 (N_1824,N_1656,N_1750);
or U1825 (N_1825,N_1672,N_1707);
nor U1826 (N_1826,N_1754,N_1735);
xnor U1827 (N_1827,N_1623,N_1761);
or U1828 (N_1828,N_1678,N_1740);
xor U1829 (N_1829,N_1625,N_1662);
and U1830 (N_1830,N_1727,N_1636);
and U1831 (N_1831,N_1603,N_1702);
and U1832 (N_1832,N_1684,N_1635);
xor U1833 (N_1833,N_1716,N_1705);
xnor U1834 (N_1834,N_1601,N_1668);
and U1835 (N_1835,N_1661,N_1631);
and U1836 (N_1836,N_1714,N_1755);
nand U1837 (N_1837,N_1791,N_1773);
xor U1838 (N_1838,N_1730,N_1709);
nor U1839 (N_1839,N_1682,N_1650);
xnor U1840 (N_1840,N_1608,N_1639);
nor U1841 (N_1841,N_1769,N_1742);
nand U1842 (N_1842,N_1733,N_1721);
or U1843 (N_1843,N_1772,N_1664);
nand U1844 (N_1844,N_1677,N_1621);
xnor U1845 (N_1845,N_1703,N_1797);
nand U1846 (N_1846,N_1609,N_1793);
nand U1847 (N_1847,N_1741,N_1686);
or U1848 (N_1848,N_1606,N_1752);
nor U1849 (N_1849,N_1618,N_1799);
xnor U1850 (N_1850,N_1765,N_1676);
or U1851 (N_1851,N_1739,N_1622);
xnor U1852 (N_1852,N_1745,N_1792);
xor U1853 (N_1853,N_1614,N_1690);
xnor U1854 (N_1854,N_1640,N_1723);
nand U1855 (N_1855,N_1751,N_1720);
or U1856 (N_1856,N_1777,N_1789);
and U1857 (N_1857,N_1757,N_1704);
nand U1858 (N_1858,N_1645,N_1756);
and U1859 (N_1859,N_1762,N_1641);
xnor U1860 (N_1860,N_1780,N_1687);
and U1861 (N_1861,N_1651,N_1663);
and U1862 (N_1862,N_1770,N_1658);
or U1863 (N_1863,N_1697,N_1632);
or U1864 (N_1864,N_1708,N_1619);
nor U1865 (N_1865,N_1786,N_1712);
nand U1866 (N_1866,N_1642,N_1667);
nor U1867 (N_1867,N_1788,N_1633);
nor U1868 (N_1868,N_1798,N_1784);
nand U1869 (N_1869,N_1610,N_1647);
nand U1870 (N_1870,N_1794,N_1717);
xor U1871 (N_1871,N_1615,N_1718);
xor U1872 (N_1872,N_1711,N_1759);
and U1873 (N_1873,N_1649,N_1785);
and U1874 (N_1874,N_1605,N_1659);
nor U1875 (N_1875,N_1671,N_1681);
nand U1876 (N_1876,N_1753,N_1643);
nand U1877 (N_1877,N_1700,N_1600);
nor U1878 (N_1878,N_1644,N_1763);
xor U1879 (N_1879,N_1648,N_1620);
and U1880 (N_1880,N_1706,N_1628);
xnor U1881 (N_1881,N_1738,N_1654);
or U1882 (N_1882,N_1638,N_1624);
or U1883 (N_1883,N_1613,N_1724);
or U1884 (N_1884,N_1746,N_1652);
xor U1885 (N_1885,N_1731,N_1602);
nor U1886 (N_1886,N_1683,N_1779);
or U1887 (N_1887,N_1744,N_1696);
nand U1888 (N_1888,N_1715,N_1612);
nor U1889 (N_1889,N_1795,N_1698);
or U1890 (N_1890,N_1688,N_1781);
nor U1891 (N_1891,N_1627,N_1719);
nor U1892 (N_1892,N_1653,N_1611);
nand U1893 (N_1893,N_1734,N_1674);
xor U1894 (N_1894,N_1695,N_1710);
xnor U1895 (N_1895,N_1701,N_1728);
xor U1896 (N_1896,N_1748,N_1655);
nand U1897 (N_1897,N_1722,N_1737);
xor U1898 (N_1898,N_1736,N_1685);
nor U1899 (N_1899,N_1774,N_1766);
and U1900 (N_1900,N_1702,N_1723);
nand U1901 (N_1901,N_1655,N_1765);
or U1902 (N_1902,N_1752,N_1776);
nor U1903 (N_1903,N_1639,N_1706);
and U1904 (N_1904,N_1690,N_1670);
and U1905 (N_1905,N_1617,N_1709);
or U1906 (N_1906,N_1704,N_1749);
nand U1907 (N_1907,N_1747,N_1797);
or U1908 (N_1908,N_1649,N_1686);
xnor U1909 (N_1909,N_1623,N_1755);
and U1910 (N_1910,N_1738,N_1730);
nor U1911 (N_1911,N_1653,N_1702);
nand U1912 (N_1912,N_1700,N_1625);
nor U1913 (N_1913,N_1779,N_1675);
and U1914 (N_1914,N_1619,N_1685);
and U1915 (N_1915,N_1610,N_1694);
xor U1916 (N_1916,N_1710,N_1782);
xnor U1917 (N_1917,N_1753,N_1791);
xnor U1918 (N_1918,N_1700,N_1696);
and U1919 (N_1919,N_1688,N_1658);
xor U1920 (N_1920,N_1601,N_1741);
nand U1921 (N_1921,N_1664,N_1702);
nand U1922 (N_1922,N_1717,N_1662);
and U1923 (N_1923,N_1761,N_1795);
xnor U1924 (N_1924,N_1628,N_1649);
nor U1925 (N_1925,N_1785,N_1697);
nand U1926 (N_1926,N_1668,N_1670);
or U1927 (N_1927,N_1748,N_1732);
nand U1928 (N_1928,N_1734,N_1768);
xnor U1929 (N_1929,N_1659,N_1738);
nor U1930 (N_1930,N_1758,N_1736);
and U1931 (N_1931,N_1695,N_1601);
nand U1932 (N_1932,N_1712,N_1678);
nor U1933 (N_1933,N_1709,N_1755);
nor U1934 (N_1934,N_1663,N_1737);
xor U1935 (N_1935,N_1739,N_1649);
nand U1936 (N_1936,N_1723,N_1606);
nor U1937 (N_1937,N_1774,N_1625);
or U1938 (N_1938,N_1762,N_1771);
nand U1939 (N_1939,N_1704,N_1701);
nand U1940 (N_1940,N_1638,N_1712);
nand U1941 (N_1941,N_1761,N_1781);
nor U1942 (N_1942,N_1673,N_1658);
or U1943 (N_1943,N_1639,N_1744);
nand U1944 (N_1944,N_1622,N_1754);
nor U1945 (N_1945,N_1605,N_1749);
nor U1946 (N_1946,N_1620,N_1757);
and U1947 (N_1947,N_1604,N_1725);
nand U1948 (N_1948,N_1781,N_1696);
nand U1949 (N_1949,N_1719,N_1670);
or U1950 (N_1950,N_1741,N_1650);
and U1951 (N_1951,N_1752,N_1765);
nor U1952 (N_1952,N_1682,N_1716);
xnor U1953 (N_1953,N_1739,N_1724);
xnor U1954 (N_1954,N_1793,N_1752);
and U1955 (N_1955,N_1670,N_1790);
or U1956 (N_1956,N_1655,N_1710);
and U1957 (N_1957,N_1632,N_1757);
or U1958 (N_1958,N_1617,N_1661);
or U1959 (N_1959,N_1780,N_1672);
nand U1960 (N_1960,N_1746,N_1760);
nand U1961 (N_1961,N_1705,N_1616);
and U1962 (N_1962,N_1677,N_1640);
nand U1963 (N_1963,N_1663,N_1749);
nand U1964 (N_1964,N_1759,N_1619);
or U1965 (N_1965,N_1688,N_1656);
xor U1966 (N_1966,N_1607,N_1700);
xnor U1967 (N_1967,N_1757,N_1755);
xnor U1968 (N_1968,N_1664,N_1663);
or U1969 (N_1969,N_1634,N_1746);
and U1970 (N_1970,N_1637,N_1740);
nor U1971 (N_1971,N_1666,N_1754);
and U1972 (N_1972,N_1668,N_1694);
nand U1973 (N_1973,N_1696,N_1673);
and U1974 (N_1974,N_1695,N_1621);
nand U1975 (N_1975,N_1613,N_1774);
and U1976 (N_1976,N_1678,N_1668);
nand U1977 (N_1977,N_1644,N_1697);
and U1978 (N_1978,N_1631,N_1665);
and U1979 (N_1979,N_1797,N_1709);
and U1980 (N_1980,N_1791,N_1615);
nand U1981 (N_1981,N_1726,N_1799);
xnor U1982 (N_1982,N_1786,N_1757);
or U1983 (N_1983,N_1612,N_1770);
and U1984 (N_1984,N_1797,N_1711);
nor U1985 (N_1985,N_1731,N_1705);
nor U1986 (N_1986,N_1763,N_1762);
nor U1987 (N_1987,N_1775,N_1690);
and U1988 (N_1988,N_1762,N_1767);
nand U1989 (N_1989,N_1734,N_1756);
xor U1990 (N_1990,N_1666,N_1687);
or U1991 (N_1991,N_1778,N_1647);
nand U1992 (N_1992,N_1791,N_1717);
xor U1993 (N_1993,N_1612,N_1710);
xor U1994 (N_1994,N_1796,N_1719);
and U1995 (N_1995,N_1789,N_1621);
nand U1996 (N_1996,N_1739,N_1771);
or U1997 (N_1997,N_1604,N_1702);
or U1998 (N_1998,N_1765,N_1768);
nor U1999 (N_1999,N_1696,N_1619);
nor U2000 (N_2000,N_1928,N_1859);
nor U2001 (N_2001,N_1822,N_1906);
and U2002 (N_2002,N_1875,N_1827);
and U2003 (N_2003,N_1828,N_1903);
xor U2004 (N_2004,N_1963,N_1948);
and U2005 (N_2005,N_1933,N_1852);
nand U2006 (N_2006,N_1954,N_1939);
and U2007 (N_2007,N_1959,N_1934);
nor U2008 (N_2008,N_1802,N_1809);
xor U2009 (N_2009,N_1816,N_1805);
or U2010 (N_2010,N_1839,N_1890);
xor U2011 (N_2011,N_1814,N_1918);
nand U2012 (N_2012,N_1987,N_1873);
nor U2013 (N_2013,N_1872,N_1853);
xor U2014 (N_2014,N_1885,N_1833);
nand U2015 (N_2015,N_1800,N_1968);
nor U2016 (N_2016,N_1994,N_1941);
nor U2017 (N_2017,N_1920,N_1971);
or U2018 (N_2018,N_1949,N_1916);
nor U2019 (N_2019,N_1819,N_1868);
and U2020 (N_2020,N_1985,N_1865);
and U2021 (N_2021,N_1808,N_1983);
xnor U2022 (N_2022,N_1843,N_1857);
and U2023 (N_2023,N_1932,N_1989);
and U2024 (N_2024,N_1919,N_1811);
nand U2025 (N_2025,N_1862,N_1801);
nand U2026 (N_2026,N_1927,N_1915);
xnor U2027 (N_2027,N_1984,N_1810);
or U2028 (N_2028,N_1891,N_1883);
nand U2029 (N_2029,N_1898,N_1854);
nand U2030 (N_2030,N_1904,N_1829);
and U2031 (N_2031,N_1860,N_1943);
nor U2032 (N_2032,N_1978,N_1937);
and U2033 (N_2033,N_1869,N_1991);
xnor U2034 (N_2034,N_1961,N_1908);
nand U2035 (N_2035,N_1922,N_1823);
nor U2036 (N_2036,N_1965,N_1938);
xor U2037 (N_2037,N_1874,N_1900);
and U2038 (N_2038,N_1884,N_1967);
nand U2039 (N_2039,N_1804,N_1956);
nand U2040 (N_2040,N_1914,N_1861);
nor U2041 (N_2041,N_1806,N_1824);
xor U2042 (N_2042,N_1813,N_1913);
and U2043 (N_2043,N_1931,N_1996);
and U2044 (N_2044,N_1831,N_1911);
or U2045 (N_2045,N_1995,N_1988);
xor U2046 (N_2046,N_1969,N_1973);
nor U2047 (N_2047,N_1817,N_1935);
and U2048 (N_2048,N_1836,N_1998);
nand U2049 (N_2049,N_1909,N_1846);
nor U2050 (N_2050,N_1929,N_1835);
nand U2051 (N_2051,N_1979,N_1886);
nand U2052 (N_2052,N_1925,N_1924);
nand U2053 (N_2053,N_1851,N_1832);
or U2054 (N_2054,N_1975,N_1821);
and U2055 (N_2055,N_1964,N_1997);
nor U2056 (N_2056,N_1951,N_1876);
or U2057 (N_2057,N_1850,N_1858);
nand U2058 (N_2058,N_1901,N_1936);
nor U2059 (N_2059,N_1990,N_1818);
xnor U2060 (N_2060,N_1826,N_1878);
and U2061 (N_2061,N_1830,N_1897);
nor U2062 (N_2062,N_1892,N_1849);
or U2063 (N_2063,N_1864,N_1863);
and U2064 (N_2064,N_1820,N_1871);
nor U2065 (N_2065,N_1977,N_1970);
or U2066 (N_2066,N_1942,N_1837);
nand U2067 (N_2067,N_1986,N_1907);
nor U2068 (N_2068,N_1917,N_1807);
or U2069 (N_2069,N_1993,N_1894);
nand U2070 (N_2070,N_1887,N_1955);
or U2071 (N_2071,N_1882,N_1844);
xor U2072 (N_2072,N_1881,N_1910);
or U2073 (N_2073,N_1889,N_1856);
or U2074 (N_2074,N_1960,N_1962);
nor U2075 (N_2075,N_1855,N_1847);
nand U2076 (N_2076,N_1879,N_1966);
xor U2077 (N_2077,N_1866,N_1870);
nor U2078 (N_2078,N_1944,N_1999);
xor U2079 (N_2079,N_1930,N_1877);
xnor U2080 (N_2080,N_1921,N_1902);
xnor U2081 (N_2081,N_1815,N_1940);
or U2082 (N_2082,N_1957,N_1992);
nor U2083 (N_2083,N_1950,N_1845);
xnor U2084 (N_2084,N_1926,N_1947);
nand U2085 (N_2085,N_1980,N_1867);
nand U2086 (N_2086,N_1803,N_1972);
and U2087 (N_2087,N_1842,N_1953);
or U2088 (N_2088,N_1981,N_1899);
and U2089 (N_2089,N_1958,N_1976);
and U2090 (N_2090,N_1838,N_1923);
and U2091 (N_2091,N_1895,N_1952);
and U2092 (N_2092,N_1893,N_1912);
xnor U2093 (N_2093,N_1812,N_1982);
nand U2094 (N_2094,N_1974,N_1841);
or U2095 (N_2095,N_1840,N_1905);
nand U2096 (N_2096,N_1834,N_1946);
nor U2097 (N_2097,N_1825,N_1880);
nand U2098 (N_2098,N_1945,N_1848);
xnor U2099 (N_2099,N_1896,N_1888);
nor U2100 (N_2100,N_1829,N_1892);
and U2101 (N_2101,N_1895,N_1820);
and U2102 (N_2102,N_1965,N_1844);
nor U2103 (N_2103,N_1887,N_1837);
nor U2104 (N_2104,N_1811,N_1847);
and U2105 (N_2105,N_1857,N_1869);
and U2106 (N_2106,N_1968,N_1856);
nor U2107 (N_2107,N_1882,N_1854);
xor U2108 (N_2108,N_1981,N_1864);
and U2109 (N_2109,N_1994,N_1811);
or U2110 (N_2110,N_1865,N_1903);
or U2111 (N_2111,N_1902,N_1900);
nand U2112 (N_2112,N_1871,N_1961);
or U2113 (N_2113,N_1814,N_1821);
nand U2114 (N_2114,N_1968,N_1939);
nor U2115 (N_2115,N_1846,N_1961);
or U2116 (N_2116,N_1910,N_1841);
nand U2117 (N_2117,N_1986,N_1849);
and U2118 (N_2118,N_1904,N_1848);
or U2119 (N_2119,N_1806,N_1807);
nand U2120 (N_2120,N_1860,N_1922);
or U2121 (N_2121,N_1979,N_1805);
nand U2122 (N_2122,N_1902,N_1924);
and U2123 (N_2123,N_1814,N_1995);
and U2124 (N_2124,N_1894,N_1829);
and U2125 (N_2125,N_1982,N_1849);
xnor U2126 (N_2126,N_1835,N_1898);
xor U2127 (N_2127,N_1904,N_1927);
nor U2128 (N_2128,N_1932,N_1871);
xor U2129 (N_2129,N_1980,N_1821);
xor U2130 (N_2130,N_1835,N_1987);
nor U2131 (N_2131,N_1862,N_1904);
xor U2132 (N_2132,N_1908,N_1927);
nand U2133 (N_2133,N_1837,N_1920);
and U2134 (N_2134,N_1917,N_1938);
xnor U2135 (N_2135,N_1880,N_1877);
xor U2136 (N_2136,N_1999,N_1900);
or U2137 (N_2137,N_1882,N_1986);
nor U2138 (N_2138,N_1954,N_1895);
xnor U2139 (N_2139,N_1991,N_1919);
nand U2140 (N_2140,N_1947,N_1898);
nor U2141 (N_2141,N_1840,N_1952);
or U2142 (N_2142,N_1860,N_1908);
nor U2143 (N_2143,N_1922,N_1848);
nand U2144 (N_2144,N_1809,N_1907);
nand U2145 (N_2145,N_1928,N_1853);
and U2146 (N_2146,N_1926,N_1843);
and U2147 (N_2147,N_1993,N_1909);
and U2148 (N_2148,N_1967,N_1909);
nor U2149 (N_2149,N_1893,N_1837);
xnor U2150 (N_2150,N_1862,N_1803);
nand U2151 (N_2151,N_1841,N_1871);
and U2152 (N_2152,N_1875,N_1820);
nand U2153 (N_2153,N_1958,N_1893);
nor U2154 (N_2154,N_1903,N_1910);
and U2155 (N_2155,N_1848,N_1978);
nand U2156 (N_2156,N_1983,N_1838);
xnor U2157 (N_2157,N_1906,N_1940);
nand U2158 (N_2158,N_1942,N_1829);
nor U2159 (N_2159,N_1931,N_1899);
xnor U2160 (N_2160,N_1949,N_1998);
or U2161 (N_2161,N_1814,N_1888);
xor U2162 (N_2162,N_1811,N_1818);
nor U2163 (N_2163,N_1969,N_1805);
or U2164 (N_2164,N_1895,N_1885);
nor U2165 (N_2165,N_1967,N_1895);
nand U2166 (N_2166,N_1978,N_1896);
and U2167 (N_2167,N_1832,N_1984);
and U2168 (N_2168,N_1949,N_1959);
nor U2169 (N_2169,N_1908,N_1880);
nand U2170 (N_2170,N_1977,N_1876);
and U2171 (N_2171,N_1883,N_1823);
nor U2172 (N_2172,N_1894,N_1983);
nor U2173 (N_2173,N_1977,N_1836);
or U2174 (N_2174,N_1892,N_1934);
nor U2175 (N_2175,N_1985,N_1894);
and U2176 (N_2176,N_1882,N_1958);
nand U2177 (N_2177,N_1927,N_1901);
and U2178 (N_2178,N_1996,N_1944);
xor U2179 (N_2179,N_1894,N_1836);
xnor U2180 (N_2180,N_1968,N_1826);
and U2181 (N_2181,N_1970,N_1895);
nand U2182 (N_2182,N_1875,N_1837);
nand U2183 (N_2183,N_1836,N_1805);
nand U2184 (N_2184,N_1847,N_1986);
nor U2185 (N_2185,N_1963,N_1860);
nor U2186 (N_2186,N_1939,N_1870);
nand U2187 (N_2187,N_1888,N_1955);
xnor U2188 (N_2188,N_1930,N_1990);
nand U2189 (N_2189,N_1805,N_1833);
or U2190 (N_2190,N_1995,N_1808);
or U2191 (N_2191,N_1828,N_1969);
and U2192 (N_2192,N_1978,N_1818);
xnor U2193 (N_2193,N_1808,N_1812);
xor U2194 (N_2194,N_1965,N_1958);
or U2195 (N_2195,N_1923,N_1849);
nor U2196 (N_2196,N_1993,N_1825);
and U2197 (N_2197,N_1803,N_1982);
nand U2198 (N_2198,N_1820,N_1992);
nand U2199 (N_2199,N_1974,N_1955);
or U2200 (N_2200,N_2029,N_2124);
xor U2201 (N_2201,N_2183,N_2184);
or U2202 (N_2202,N_2120,N_2071);
xor U2203 (N_2203,N_2078,N_2160);
or U2204 (N_2204,N_2012,N_2043);
nor U2205 (N_2205,N_2158,N_2059);
nor U2206 (N_2206,N_2027,N_2005);
or U2207 (N_2207,N_2166,N_2190);
nand U2208 (N_2208,N_2168,N_2149);
and U2209 (N_2209,N_2000,N_2137);
or U2210 (N_2210,N_2019,N_2095);
and U2211 (N_2211,N_2172,N_2165);
and U2212 (N_2212,N_2135,N_2195);
nor U2213 (N_2213,N_2180,N_2018);
and U2214 (N_2214,N_2145,N_2098);
or U2215 (N_2215,N_2041,N_2131);
nor U2216 (N_2216,N_2020,N_2118);
nor U2217 (N_2217,N_2082,N_2117);
and U2218 (N_2218,N_2141,N_2067);
nor U2219 (N_2219,N_2154,N_2143);
and U2220 (N_2220,N_2077,N_2127);
and U2221 (N_2221,N_2147,N_2113);
xor U2222 (N_2222,N_2128,N_2001);
nand U2223 (N_2223,N_2044,N_2036);
nor U2224 (N_2224,N_2161,N_2133);
and U2225 (N_2225,N_2048,N_2104);
nor U2226 (N_2226,N_2076,N_2170);
nand U2227 (N_2227,N_2004,N_2159);
or U2228 (N_2228,N_2092,N_2070);
nor U2229 (N_2229,N_2016,N_2199);
or U2230 (N_2230,N_2189,N_2047);
and U2231 (N_2231,N_2148,N_2176);
xnor U2232 (N_2232,N_2032,N_2175);
nor U2233 (N_2233,N_2088,N_2009);
xor U2234 (N_2234,N_2139,N_2123);
nor U2235 (N_2235,N_2034,N_2063);
xor U2236 (N_2236,N_2052,N_2126);
and U2237 (N_2237,N_2191,N_2197);
xnor U2238 (N_2238,N_2023,N_2085);
or U2239 (N_2239,N_2013,N_2116);
and U2240 (N_2240,N_2039,N_2167);
nand U2241 (N_2241,N_2010,N_2015);
xnor U2242 (N_2242,N_2073,N_2130);
nor U2243 (N_2243,N_2090,N_2182);
nand U2244 (N_2244,N_2026,N_2134);
and U2245 (N_2245,N_2198,N_2142);
or U2246 (N_2246,N_2103,N_2038);
and U2247 (N_2247,N_2171,N_2062);
and U2248 (N_2248,N_2089,N_2025);
nor U2249 (N_2249,N_2028,N_2022);
nand U2250 (N_2250,N_2080,N_2006);
nor U2251 (N_2251,N_2030,N_2107);
nor U2252 (N_2252,N_2101,N_2066);
or U2253 (N_2253,N_2068,N_2136);
xor U2254 (N_2254,N_2188,N_2035);
or U2255 (N_2255,N_2040,N_2169);
or U2256 (N_2256,N_2065,N_2093);
and U2257 (N_2257,N_2164,N_2054);
and U2258 (N_2258,N_2109,N_2056);
and U2259 (N_2259,N_2129,N_2173);
or U2260 (N_2260,N_2181,N_2058);
nand U2261 (N_2261,N_2051,N_2187);
nor U2262 (N_2262,N_2053,N_2061);
nor U2263 (N_2263,N_2045,N_2091);
nor U2264 (N_2264,N_2152,N_2049);
xnor U2265 (N_2265,N_2096,N_2193);
xor U2266 (N_2266,N_2024,N_2074);
nor U2267 (N_2267,N_2122,N_2007);
and U2268 (N_2268,N_2194,N_2075);
or U2269 (N_2269,N_2146,N_2162);
and U2270 (N_2270,N_2121,N_2033);
and U2271 (N_2271,N_2153,N_2021);
nor U2272 (N_2272,N_2115,N_2108);
xnor U2273 (N_2273,N_2100,N_2112);
or U2274 (N_2274,N_2099,N_2125);
or U2275 (N_2275,N_2057,N_2196);
nor U2276 (N_2276,N_2046,N_2083);
xnor U2277 (N_2277,N_2132,N_2037);
and U2278 (N_2278,N_2177,N_2156);
nor U2279 (N_2279,N_2106,N_2151);
nand U2280 (N_2280,N_2185,N_2144);
nand U2281 (N_2281,N_2179,N_2111);
nor U2282 (N_2282,N_2069,N_2014);
nor U2283 (N_2283,N_2186,N_2105);
and U2284 (N_2284,N_2081,N_2119);
xnor U2285 (N_2285,N_2084,N_2174);
or U2286 (N_2286,N_2192,N_2114);
nor U2287 (N_2287,N_2138,N_2094);
and U2288 (N_2288,N_2008,N_2155);
or U2289 (N_2289,N_2060,N_2011);
and U2290 (N_2290,N_2087,N_2102);
xnor U2291 (N_2291,N_2140,N_2042);
nor U2292 (N_2292,N_2157,N_2086);
nor U2293 (N_2293,N_2002,N_2110);
and U2294 (N_2294,N_2055,N_2079);
or U2295 (N_2295,N_2031,N_2163);
nand U2296 (N_2296,N_2064,N_2003);
and U2297 (N_2297,N_2178,N_2017);
nor U2298 (N_2298,N_2097,N_2050);
or U2299 (N_2299,N_2072,N_2150);
nand U2300 (N_2300,N_2193,N_2035);
nand U2301 (N_2301,N_2179,N_2195);
nor U2302 (N_2302,N_2048,N_2020);
xnor U2303 (N_2303,N_2170,N_2066);
or U2304 (N_2304,N_2185,N_2101);
nor U2305 (N_2305,N_2198,N_2096);
nand U2306 (N_2306,N_2118,N_2016);
nand U2307 (N_2307,N_2110,N_2181);
nor U2308 (N_2308,N_2077,N_2152);
nand U2309 (N_2309,N_2056,N_2156);
and U2310 (N_2310,N_2167,N_2148);
xnor U2311 (N_2311,N_2176,N_2057);
nor U2312 (N_2312,N_2190,N_2176);
and U2313 (N_2313,N_2064,N_2108);
nand U2314 (N_2314,N_2087,N_2046);
and U2315 (N_2315,N_2161,N_2040);
or U2316 (N_2316,N_2051,N_2110);
xor U2317 (N_2317,N_2038,N_2102);
and U2318 (N_2318,N_2071,N_2139);
and U2319 (N_2319,N_2102,N_2176);
nor U2320 (N_2320,N_2195,N_2014);
or U2321 (N_2321,N_2087,N_2010);
nor U2322 (N_2322,N_2080,N_2077);
xor U2323 (N_2323,N_2141,N_2179);
and U2324 (N_2324,N_2115,N_2021);
xor U2325 (N_2325,N_2169,N_2130);
and U2326 (N_2326,N_2156,N_2090);
nor U2327 (N_2327,N_2065,N_2123);
xnor U2328 (N_2328,N_2019,N_2066);
or U2329 (N_2329,N_2040,N_2193);
xnor U2330 (N_2330,N_2152,N_2020);
and U2331 (N_2331,N_2089,N_2140);
nor U2332 (N_2332,N_2057,N_2101);
nor U2333 (N_2333,N_2115,N_2193);
and U2334 (N_2334,N_2100,N_2014);
nor U2335 (N_2335,N_2047,N_2146);
or U2336 (N_2336,N_2029,N_2011);
and U2337 (N_2337,N_2025,N_2022);
and U2338 (N_2338,N_2000,N_2144);
nand U2339 (N_2339,N_2080,N_2175);
and U2340 (N_2340,N_2056,N_2108);
and U2341 (N_2341,N_2050,N_2043);
xor U2342 (N_2342,N_2074,N_2092);
nand U2343 (N_2343,N_2005,N_2049);
nor U2344 (N_2344,N_2134,N_2136);
xor U2345 (N_2345,N_2003,N_2194);
or U2346 (N_2346,N_2126,N_2058);
xnor U2347 (N_2347,N_2142,N_2191);
or U2348 (N_2348,N_2177,N_2021);
nor U2349 (N_2349,N_2119,N_2044);
and U2350 (N_2350,N_2133,N_2148);
nor U2351 (N_2351,N_2123,N_2145);
xor U2352 (N_2352,N_2124,N_2024);
and U2353 (N_2353,N_2033,N_2004);
or U2354 (N_2354,N_2083,N_2010);
xnor U2355 (N_2355,N_2034,N_2020);
xor U2356 (N_2356,N_2138,N_2140);
or U2357 (N_2357,N_2115,N_2012);
and U2358 (N_2358,N_2113,N_2164);
and U2359 (N_2359,N_2038,N_2020);
xnor U2360 (N_2360,N_2091,N_2135);
or U2361 (N_2361,N_2197,N_2078);
nor U2362 (N_2362,N_2043,N_2030);
and U2363 (N_2363,N_2009,N_2033);
or U2364 (N_2364,N_2085,N_2026);
or U2365 (N_2365,N_2037,N_2156);
nor U2366 (N_2366,N_2117,N_2177);
nor U2367 (N_2367,N_2089,N_2003);
xor U2368 (N_2368,N_2159,N_2121);
nor U2369 (N_2369,N_2002,N_2073);
and U2370 (N_2370,N_2131,N_2171);
and U2371 (N_2371,N_2177,N_2070);
and U2372 (N_2372,N_2065,N_2074);
nand U2373 (N_2373,N_2156,N_2135);
and U2374 (N_2374,N_2030,N_2113);
or U2375 (N_2375,N_2184,N_2068);
nor U2376 (N_2376,N_2131,N_2199);
xnor U2377 (N_2377,N_2139,N_2061);
nor U2378 (N_2378,N_2163,N_2002);
nor U2379 (N_2379,N_2001,N_2193);
nor U2380 (N_2380,N_2168,N_2129);
xnor U2381 (N_2381,N_2088,N_2166);
or U2382 (N_2382,N_2160,N_2049);
nand U2383 (N_2383,N_2096,N_2045);
nand U2384 (N_2384,N_2118,N_2084);
nor U2385 (N_2385,N_2137,N_2095);
xor U2386 (N_2386,N_2161,N_2089);
xor U2387 (N_2387,N_2192,N_2174);
xnor U2388 (N_2388,N_2108,N_2159);
or U2389 (N_2389,N_2011,N_2046);
xnor U2390 (N_2390,N_2068,N_2027);
and U2391 (N_2391,N_2151,N_2035);
nand U2392 (N_2392,N_2024,N_2017);
or U2393 (N_2393,N_2105,N_2026);
or U2394 (N_2394,N_2017,N_2172);
or U2395 (N_2395,N_2065,N_2157);
or U2396 (N_2396,N_2125,N_2121);
or U2397 (N_2397,N_2058,N_2105);
xor U2398 (N_2398,N_2073,N_2077);
and U2399 (N_2399,N_2146,N_2155);
or U2400 (N_2400,N_2242,N_2229);
and U2401 (N_2401,N_2279,N_2281);
nor U2402 (N_2402,N_2297,N_2348);
or U2403 (N_2403,N_2303,N_2386);
or U2404 (N_2404,N_2390,N_2374);
xor U2405 (N_2405,N_2305,N_2313);
and U2406 (N_2406,N_2234,N_2333);
and U2407 (N_2407,N_2310,N_2252);
or U2408 (N_2408,N_2315,N_2209);
or U2409 (N_2409,N_2391,N_2253);
nand U2410 (N_2410,N_2328,N_2219);
xnor U2411 (N_2411,N_2384,N_2366);
or U2412 (N_2412,N_2357,N_2233);
and U2413 (N_2413,N_2228,N_2277);
nand U2414 (N_2414,N_2217,N_2284);
or U2415 (N_2415,N_2250,N_2389);
and U2416 (N_2416,N_2267,N_2353);
xnor U2417 (N_2417,N_2369,N_2396);
xnor U2418 (N_2418,N_2342,N_2240);
xnor U2419 (N_2419,N_2235,N_2225);
or U2420 (N_2420,N_2266,N_2370);
nor U2421 (N_2421,N_2356,N_2201);
nand U2422 (N_2422,N_2324,N_2330);
and U2423 (N_2423,N_2398,N_2245);
nor U2424 (N_2424,N_2377,N_2260);
xnor U2425 (N_2425,N_2285,N_2283);
nand U2426 (N_2426,N_2214,N_2208);
nor U2427 (N_2427,N_2382,N_2254);
nand U2428 (N_2428,N_2392,N_2215);
nand U2429 (N_2429,N_2367,N_2339);
nand U2430 (N_2430,N_2327,N_2336);
nor U2431 (N_2431,N_2272,N_2322);
xor U2432 (N_2432,N_2223,N_2202);
and U2433 (N_2433,N_2212,N_2273);
or U2434 (N_2434,N_2294,N_2221);
nor U2435 (N_2435,N_2372,N_2292);
or U2436 (N_2436,N_2352,N_2218);
xor U2437 (N_2437,N_2331,N_2231);
and U2438 (N_2438,N_2329,N_2230);
nand U2439 (N_2439,N_2319,N_2255);
and U2440 (N_2440,N_2290,N_2204);
nand U2441 (N_2441,N_2244,N_2317);
nand U2442 (N_2442,N_2347,N_2349);
nand U2443 (N_2443,N_2321,N_2371);
xor U2444 (N_2444,N_2270,N_2261);
and U2445 (N_2445,N_2318,N_2379);
and U2446 (N_2446,N_2278,N_2359);
xnor U2447 (N_2447,N_2335,N_2332);
nor U2448 (N_2448,N_2393,N_2309);
and U2449 (N_2449,N_2222,N_2334);
and U2450 (N_2450,N_2326,N_2205);
and U2451 (N_2451,N_2236,N_2320);
nor U2452 (N_2452,N_2210,N_2341);
and U2453 (N_2453,N_2307,N_2306);
nor U2454 (N_2454,N_2262,N_2376);
or U2455 (N_2455,N_2394,N_2368);
nand U2456 (N_2456,N_2375,N_2207);
xnor U2457 (N_2457,N_2314,N_2340);
or U2458 (N_2458,N_2289,N_2249);
nor U2459 (N_2459,N_2232,N_2247);
or U2460 (N_2460,N_2206,N_2256);
nand U2461 (N_2461,N_2346,N_2259);
nand U2462 (N_2462,N_2360,N_2387);
nand U2463 (N_2463,N_2216,N_2304);
nand U2464 (N_2464,N_2373,N_2263);
xor U2465 (N_2465,N_2343,N_2399);
nor U2466 (N_2466,N_2280,N_2395);
or U2467 (N_2467,N_2378,N_2226);
xnor U2468 (N_2468,N_2203,N_2323);
nand U2469 (N_2469,N_2337,N_2354);
nand U2470 (N_2470,N_2286,N_2388);
or U2471 (N_2471,N_2271,N_2344);
and U2472 (N_2472,N_2325,N_2264);
or U2473 (N_2473,N_2269,N_2213);
or U2474 (N_2474,N_2288,N_2351);
nand U2475 (N_2475,N_2363,N_2265);
nand U2476 (N_2476,N_2316,N_2211);
and U2477 (N_2477,N_2243,N_2302);
nor U2478 (N_2478,N_2380,N_2296);
xnor U2479 (N_2479,N_2287,N_2301);
nor U2480 (N_2480,N_2224,N_2350);
nor U2481 (N_2481,N_2275,N_2308);
nor U2482 (N_2482,N_2282,N_2362);
nor U2483 (N_2483,N_2298,N_2274);
nand U2484 (N_2484,N_2246,N_2311);
and U2485 (N_2485,N_2300,N_2358);
nor U2486 (N_2486,N_2248,N_2220);
xnor U2487 (N_2487,N_2237,N_2365);
nor U2488 (N_2488,N_2397,N_2361);
or U2489 (N_2489,N_2355,N_2338);
and U2490 (N_2490,N_2364,N_2381);
and U2491 (N_2491,N_2276,N_2241);
nor U2492 (N_2492,N_2385,N_2312);
xnor U2493 (N_2493,N_2345,N_2268);
nand U2494 (N_2494,N_2291,N_2200);
nand U2495 (N_2495,N_2258,N_2299);
or U2496 (N_2496,N_2251,N_2227);
xor U2497 (N_2497,N_2383,N_2293);
xnor U2498 (N_2498,N_2295,N_2238);
or U2499 (N_2499,N_2239,N_2257);
and U2500 (N_2500,N_2264,N_2371);
nand U2501 (N_2501,N_2308,N_2323);
xnor U2502 (N_2502,N_2240,N_2311);
nor U2503 (N_2503,N_2261,N_2314);
xor U2504 (N_2504,N_2383,N_2251);
nand U2505 (N_2505,N_2351,N_2367);
xor U2506 (N_2506,N_2329,N_2386);
nor U2507 (N_2507,N_2217,N_2306);
nand U2508 (N_2508,N_2231,N_2350);
nor U2509 (N_2509,N_2385,N_2370);
or U2510 (N_2510,N_2333,N_2236);
or U2511 (N_2511,N_2334,N_2227);
nor U2512 (N_2512,N_2269,N_2284);
nor U2513 (N_2513,N_2288,N_2251);
nor U2514 (N_2514,N_2305,N_2254);
or U2515 (N_2515,N_2396,N_2353);
nor U2516 (N_2516,N_2358,N_2375);
and U2517 (N_2517,N_2324,N_2340);
nand U2518 (N_2518,N_2352,N_2365);
nor U2519 (N_2519,N_2366,N_2334);
nand U2520 (N_2520,N_2321,N_2283);
nand U2521 (N_2521,N_2245,N_2276);
or U2522 (N_2522,N_2227,N_2356);
nand U2523 (N_2523,N_2266,N_2275);
xor U2524 (N_2524,N_2298,N_2275);
or U2525 (N_2525,N_2246,N_2258);
xnor U2526 (N_2526,N_2356,N_2392);
or U2527 (N_2527,N_2246,N_2299);
nor U2528 (N_2528,N_2232,N_2318);
and U2529 (N_2529,N_2276,N_2271);
nand U2530 (N_2530,N_2361,N_2375);
xor U2531 (N_2531,N_2353,N_2360);
xnor U2532 (N_2532,N_2357,N_2246);
or U2533 (N_2533,N_2234,N_2384);
or U2534 (N_2534,N_2377,N_2369);
or U2535 (N_2535,N_2235,N_2264);
or U2536 (N_2536,N_2301,N_2386);
xor U2537 (N_2537,N_2305,N_2292);
xor U2538 (N_2538,N_2327,N_2390);
nand U2539 (N_2539,N_2384,N_2357);
nor U2540 (N_2540,N_2339,N_2210);
xnor U2541 (N_2541,N_2382,N_2344);
nand U2542 (N_2542,N_2205,N_2381);
xnor U2543 (N_2543,N_2349,N_2343);
xnor U2544 (N_2544,N_2331,N_2376);
and U2545 (N_2545,N_2264,N_2381);
and U2546 (N_2546,N_2295,N_2244);
and U2547 (N_2547,N_2348,N_2369);
or U2548 (N_2548,N_2390,N_2241);
nor U2549 (N_2549,N_2366,N_2204);
or U2550 (N_2550,N_2360,N_2304);
nand U2551 (N_2551,N_2248,N_2305);
and U2552 (N_2552,N_2232,N_2352);
xnor U2553 (N_2553,N_2329,N_2367);
or U2554 (N_2554,N_2363,N_2278);
xnor U2555 (N_2555,N_2398,N_2261);
or U2556 (N_2556,N_2328,N_2322);
nand U2557 (N_2557,N_2292,N_2302);
or U2558 (N_2558,N_2379,N_2216);
xnor U2559 (N_2559,N_2389,N_2249);
nor U2560 (N_2560,N_2383,N_2310);
xor U2561 (N_2561,N_2399,N_2276);
and U2562 (N_2562,N_2391,N_2217);
nand U2563 (N_2563,N_2319,N_2250);
nor U2564 (N_2564,N_2239,N_2232);
and U2565 (N_2565,N_2353,N_2240);
nor U2566 (N_2566,N_2213,N_2380);
nand U2567 (N_2567,N_2277,N_2275);
nor U2568 (N_2568,N_2310,N_2392);
and U2569 (N_2569,N_2299,N_2307);
and U2570 (N_2570,N_2391,N_2382);
and U2571 (N_2571,N_2385,N_2301);
or U2572 (N_2572,N_2312,N_2249);
nand U2573 (N_2573,N_2213,N_2279);
xnor U2574 (N_2574,N_2212,N_2260);
and U2575 (N_2575,N_2237,N_2236);
nand U2576 (N_2576,N_2269,N_2341);
and U2577 (N_2577,N_2283,N_2326);
or U2578 (N_2578,N_2231,N_2389);
or U2579 (N_2579,N_2265,N_2304);
and U2580 (N_2580,N_2376,N_2302);
and U2581 (N_2581,N_2348,N_2267);
and U2582 (N_2582,N_2287,N_2296);
nor U2583 (N_2583,N_2316,N_2270);
nand U2584 (N_2584,N_2236,N_2274);
xor U2585 (N_2585,N_2392,N_2340);
nand U2586 (N_2586,N_2359,N_2370);
or U2587 (N_2587,N_2365,N_2322);
or U2588 (N_2588,N_2353,N_2225);
or U2589 (N_2589,N_2283,N_2234);
xor U2590 (N_2590,N_2247,N_2241);
and U2591 (N_2591,N_2235,N_2200);
nor U2592 (N_2592,N_2221,N_2370);
xnor U2593 (N_2593,N_2239,N_2336);
nand U2594 (N_2594,N_2322,N_2355);
nor U2595 (N_2595,N_2217,N_2258);
nor U2596 (N_2596,N_2392,N_2231);
nor U2597 (N_2597,N_2240,N_2233);
or U2598 (N_2598,N_2390,N_2283);
or U2599 (N_2599,N_2289,N_2266);
nand U2600 (N_2600,N_2489,N_2554);
nand U2601 (N_2601,N_2419,N_2481);
xnor U2602 (N_2602,N_2461,N_2404);
xnor U2603 (N_2603,N_2541,N_2584);
nor U2604 (N_2604,N_2587,N_2409);
or U2605 (N_2605,N_2508,N_2557);
xnor U2606 (N_2606,N_2411,N_2491);
xnor U2607 (N_2607,N_2414,N_2475);
xnor U2608 (N_2608,N_2438,N_2454);
and U2609 (N_2609,N_2552,N_2548);
xor U2610 (N_2610,N_2500,N_2518);
xnor U2611 (N_2611,N_2429,N_2553);
or U2612 (N_2612,N_2441,N_2527);
and U2613 (N_2613,N_2458,N_2580);
or U2614 (N_2614,N_2559,N_2456);
nor U2615 (N_2615,N_2550,N_2528);
and U2616 (N_2616,N_2540,N_2578);
nor U2617 (N_2617,N_2476,N_2569);
or U2618 (N_2618,N_2565,N_2446);
nand U2619 (N_2619,N_2581,N_2465);
xor U2620 (N_2620,N_2586,N_2591);
xor U2621 (N_2621,N_2537,N_2504);
or U2622 (N_2622,N_2472,N_2417);
nor U2623 (N_2623,N_2450,N_2597);
or U2624 (N_2624,N_2435,N_2480);
and U2625 (N_2625,N_2543,N_2596);
xor U2626 (N_2626,N_2524,N_2514);
nor U2627 (N_2627,N_2415,N_2471);
nor U2628 (N_2628,N_2583,N_2558);
nor U2629 (N_2629,N_2505,N_2462);
and U2630 (N_2630,N_2453,N_2468);
or U2631 (N_2631,N_2432,N_2466);
nor U2632 (N_2632,N_2460,N_2568);
nor U2633 (N_2633,N_2422,N_2592);
or U2634 (N_2634,N_2571,N_2562);
and U2635 (N_2635,N_2572,N_2521);
nand U2636 (N_2636,N_2436,N_2449);
xnor U2637 (N_2637,N_2561,N_2512);
xnor U2638 (N_2638,N_2551,N_2515);
nand U2639 (N_2639,N_2479,N_2503);
or U2640 (N_2640,N_2520,N_2511);
xnor U2641 (N_2641,N_2555,N_2522);
xor U2642 (N_2642,N_2443,N_2566);
nor U2643 (N_2643,N_2517,N_2542);
nand U2644 (N_2644,N_2532,N_2531);
or U2645 (N_2645,N_2485,N_2579);
xnor U2646 (N_2646,N_2513,N_2467);
nand U2647 (N_2647,N_2406,N_2423);
and U2648 (N_2648,N_2455,N_2473);
or U2649 (N_2649,N_2477,N_2405);
or U2650 (N_2650,N_2431,N_2442);
or U2651 (N_2651,N_2488,N_2594);
xor U2652 (N_2652,N_2538,N_2440);
nor U2653 (N_2653,N_2434,N_2530);
xor U2654 (N_2654,N_2501,N_2577);
or U2655 (N_2655,N_2563,N_2544);
nand U2656 (N_2656,N_2588,N_2483);
xnor U2657 (N_2657,N_2547,N_2556);
and U2658 (N_2658,N_2437,N_2595);
and U2659 (N_2659,N_2498,N_2421);
nor U2660 (N_2660,N_2516,N_2494);
xnor U2661 (N_2661,N_2576,N_2535);
or U2662 (N_2662,N_2448,N_2510);
xnor U2663 (N_2663,N_2523,N_2425);
nor U2664 (N_2664,N_2487,N_2447);
xnor U2665 (N_2665,N_2507,N_2567);
xor U2666 (N_2666,N_2590,N_2582);
and U2667 (N_2667,N_2493,N_2574);
xnor U2668 (N_2668,N_2402,N_2598);
nand U2669 (N_2669,N_2478,N_2457);
nor U2670 (N_2670,N_2539,N_2599);
or U2671 (N_2671,N_2420,N_2430);
nand U2672 (N_2672,N_2408,N_2412);
nand U2673 (N_2673,N_2573,N_2451);
nor U2674 (N_2674,N_2506,N_2496);
or U2675 (N_2675,N_2495,N_2546);
or U2676 (N_2676,N_2545,N_2464);
xnor U2677 (N_2677,N_2413,N_2490);
nor U2678 (N_2678,N_2492,N_2452);
xnor U2679 (N_2679,N_2593,N_2401);
nor U2680 (N_2680,N_2470,N_2526);
and U2681 (N_2681,N_2482,N_2560);
xor U2682 (N_2682,N_2410,N_2484);
nor U2683 (N_2683,N_2424,N_2529);
xnor U2684 (N_2684,N_2433,N_2426);
xor U2685 (N_2685,N_2445,N_2439);
and U2686 (N_2686,N_2416,N_2519);
xor U2687 (N_2687,N_2533,N_2463);
nor U2688 (N_2688,N_2497,N_2400);
nor U2689 (N_2689,N_2570,N_2407);
and U2690 (N_2690,N_2486,N_2509);
xor U2691 (N_2691,N_2403,N_2459);
nor U2692 (N_2692,N_2536,N_2564);
nand U2693 (N_2693,N_2444,N_2549);
nor U2694 (N_2694,N_2499,N_2575);
xnor U2695 (N_2695,N_2428,N_2427);
nor U2696 (N_2696,N_2525,N_2589);
nand U2697 (N_2697,N_2502,N_2585);
nand U2698 (N_2698,N_2534,N_2469);
or U2699 (N_2699,N_2474,N_2418);
nand U2700 (N_2700,N_2436,N_2527);
xor U2701 (N_2701,N_2589,N_2427);
nand U2702 (N_2702,N_2532,N_2465);
nor U2703 (N_2703,N_2575,N_2449);
nand U2704 (N_2704,N_2517,N_2505);
and U2705 (N_2705,N_2433,N_2596);
or U2706 (N_2706,N_2595,N_2403);
and U2707 (N_2707,N_2523,N_2570);
or U2708 (N_2708,N_2469,N_2448);
and U2709 (N_2709,N_2466,N_2444);
nor U2710 (N_2710,N_2528,N_2536);
or U2711 (N_2711,N_2499,N_2595);
and U2712 (N_2712,N_2597,N_2436);
or U2713 (N_2713,N_2517,N_2529);
or U2714 (N_2714,N_2428,N_2403);
and U2715 (N_2715,N_2446,N_2583);
and U2716 (N_2716,N_2593,N_2590);
xor U2717 (N_2717,N_2587,N_2588);
nor U2718 (N_2718,N_2557,N_2406);
or U2719 (N_2719,N_2534,N_2503);
and U2720 (N_2720,N_2400,N_2517);
xnor U2721 (N_2721,N_2487,N_2501);
or U2722 (N_2722,N_2430,N_2498);
or U2723 (N_2723,N_2430,N_2461);
nand U2724 (N_2724,N_2481,N_2435);
nor U2725 (N_2725,N_2585,N_2570);
and U2726 (N_2726,N_2565,N_2405);
and U2727 (N_2727,N_2501,N_2442);
nand U2728 (N_2728,N_2576,N_2483);
and U2729 (N_2729,N_2571,N_2560);
nand U2730 (N_2730,N_2565,N_2429);
nand U2731 (N_2731,N_2567,N_2552);
or U2732 (N_2732,N_2468,N_2438);
nand U2733 (N_2733,N_2478,N_2538);
xnor U2734 (N_2734,N_2400,N_2540);
or U2735 (N_2735,N_2569,N_2404);
xor U2736 (N_2736,N_2567,N_2514);
nor U2737 (N_2737,N_2436,N_2448);
nor U2738 (N_2738,N_2568,N_2592);
nor U2739 (N_2739,N_2507,N_2408);
or U2740 (N_2740,N_2530,N_2418);
xor U2741 (N_2741,N_2410,N_2427);
and U2742 (N_2742,N_2410,N_2446);
or U2743 (N_2743,N_2490,N_2431);
nand U2744 (N_2744,N_2510,N_2589);
xnor U2745 (N_2745,N_2525,N_2539);
or U2746 (N_2746,N_2582,N_2548);
or U2747 (N_2747,N_2500,N_2523);
xnor U2748 (N_2748,N_2521,N_2445);
xor U2749 (N_2749,N_2447,N_2404);
xor U2750 (N_2750,N_2433,N_2517);
or U2751 (N_2751,N_2555,N_2580);
nand U2752 (N_2752,N_2462,N_2464);
and U2753 (N_2753,N_2534,N_2565);
nor U2754 (N_2754,N_2405,N_2531);
xnor U2755 (N_2755,N_2414,N_2505);
nand U2756 (N_2756,N_2429,N_2566);
and U2757 (N_2757,N_2487,N_2536);
or U2758 (N_2758,N_2521,N_2543);
and U2759 (N_2759,N_2537,N_2591);
or U2760 (N_2760,N_2443,N_2420);
and U2761 (N_2761,N_2562,N_2461);
xnor U2762 (N_2762,N_2547,N_2595);
and U2763 (N_2763,N_2521,N_2517);
and U2764 (N_2764,N_2460,N_2589);
xnor U2765 (N_2765,N_2556,N_2581);
nand U2766 (N_2766,N_2482,N_2527);
nand U2767 (N_2767,N_2448,N_2577);
or U2768 (N_2768,N_2497,N_2465);
xor U2769 (N_2769,N_2573,N_2424);
or U2770 (N_2770,N_2502,N_2584);
or U2771 (N_2771,N_2525,N_2565);
or U2772 (N_2772,N_2502,N_2490);
or U2773 (N_2773,N_2489,N_2450);
nor U2774 (N_2774,N_2562,N_2558);
xor U2775 (N_2775,N_2426,N_2562);
nand U2776 (N_2776,N_2466,N_2469);
nor U2777 (N_2777,N_2438,N_2597);
or U2778 (N_2778,N_2572,N_2423);
xnor U2779 (N_2779,N_2583,N_2466);
or U2780 (N_2780,N_2590,N_2556);
nor U2781 (N_2781,N_2508,N_2433);
nor U2782 (N_2782,N_2442,N_2447);
or U2783 (N_2783,N_2592,N_2419);
nor U2784 (N_2784,N_2528,N_2537);
nand U2785 (N_2785,N_2564,N_2484);
xnor U2786 (N_2786,N_2535,N_2460);
nand U2787 (N_2787,N_2430,N_2432);
xor U2788 (N_2788,N_2472,N_2448);
and U2789 (N_2789,N_2574,N_2587);
nor U2790 (N_2790,N_2529,N_2582);
nor U2791 (N_2791,N_2485,N_2489);
nor U2792 (N_2792,N_2585,N_2510);
xor U2793 (N_2793,N_2417,N_2559);
and U2794 (N_2794,N_2590,N_2468);
or U2795 (N_2795,N_2493,N_2443);
and U2796 (N_2796,N_2538,N_2581);
and U2797 (N_2797,N_2469,N_2438);
or U2798 (N_2798,N_2443,N_2520);
and U2799 (N_2799,N_2480,N_2505);
or U2800 (N_2800,N_2654,N_2789);
or U2801 (N_2801,N_2703,N_2619);
and U2802 (N_2802,N_2651,N_2675);
xnor U2803 (N_2803,N_2667,N_2671);
xor U2804 (N_2804,N_2749,N_2732);
xnor U2805 (N_2805,N_2791,N_2645);
and U2806 (N_2806,N_2722,N_2674);
and U2807 (N_2807,N_2642,N_2699);
or U2808 (N_2808,N_2668,N_2603);
xor U2809 (N_2809,N_2765,N_2720);
or U2810 (N_2810,N_2794,N_2729);
or U2811 (N_2811,N_2751,N_2778);
xor U2812 (N_2812,N_2747,N_2723);
nand U2813 (N_2813,N_2679,N_2775);
xnor U2814 (N_2814,N_2786,N_2683);
nor U2815 (N_2815,N_2743,N_2680);
nor U2816 (N_2816,N_2664,N_2684);
or U2817 (N_2817,N_2735,N_2689);
xor U2818 (N_2818,N_2705,N_2643);
or U2819 (N_2819,N_2681,N_2741);
nand U2820 (N_2820,N_2677,N_2672);
nand U2821 (N_2821,N_2618,N_2781);
nor U2822 (N_2822,N_2727,N_2624);
or U2823 (N_2823,N_2607,N_2669);
nor U2824 (N_2824,N_2774,N_2780);
and U2825 (N_2825,N_2777,N_2627);
nand U2826 (N_2826,N_2754,N_2660);
nand U2827 (N_2827,N_2663,N_2620);
or U2828 (N_2828,N_2712,N_2628);
xnor U2829 (N_2829,N_2739,N_2752);
nor U2830 (N_2830,N_2695,N_2795);
or U2831 (N_2831,N_2636,N_2625);
xor U2832 (N_2832,N_2792,N_2767);
nand U2833 (N_2833,N_2616,N_2763);
or U2834 (N_2834,N_2662,N_2612);
and U2835 (N_2835,N_2733,N_2682);
or U2836 (N_2836,N_2773,N_2711);
xor U2837 (N_2837,N_2617,N_2764);
nor U2838 (N_2838,N_2641,N_2710);
xnor U2839 (N_2839,N_2782,N_2644);
nand U2840 (N_2840,N_2728,N_2796);
nand U2841 (N_2841,N_2713,N_2746);
and U2842 (N_2842,N_2633,N_2652);
nor U2843 (N_2843,N_2716,N_2647);
and U2844 (N_2844,N_2686,N_2707);
or U2845 (N_2845,N_2646,N_2772);
nor U2846 (N_2846,N_2629,N_2649);
and U2847 (N_2847,N_2788,N_2701);
xnor U2848 (N_2848,N_2717,N_2606);
nand U2849 (N_2849,N_2718,N_2631);
and U2850 (N_2850,N_2742,N_2687);
xor U2851 (N_2851,N_2638,N_2608);
xor U2852 (N_2852,N_2600,N_2704);
and U2853 (N_2853,N_2748,N_2700);
and U2854 (N_2854,N_2784,N_2771);
nor U2855 (N_2855,N_2670,N_2610);
nand U2856 (N_2856,N_2605,N_2760);
and U2857 (N_2857,N_2799,N_2637);
or U2858 (N_2858,N_2762,N_2696);
nor U2859 (N_2859,N_2693,N_2621);
or U2860 (N_2860,N_2691,N_2653);
nor U2861 (N_2861,N_2634,N_2657);
and U2862 (N_2862,N_2761,N_2736);
and U2863 (N_2863,N_2632,N_2787);
nor U2864 (N_2864,N_2744,N_2685);
xnor U2865 (N_2865,N_2726,N_2724);
nand U2866 (N_2866,N_2630,N_2656);
or U2867 (N_2867,N_2783,N_2655);
or U2868 (N_2868,N_2639,N_2769);
xnor U2869 (N_2869,N_2758,N_2715);
or U2870 (N_2870,N_2601,N_2740);
nand U2871 (N_2871,N_2658,N_2702);
and U2872 (N_2872,N_2759,N_2753);
nand U2873 (N_2873,N_2623,N_2650);
or U2874 (N_2874,N_2790,N_2798);
nand U2875 (N_2875,N_2725,N_2745);
or U2876 (N_2876,N_2738,N_2602);
or U2877 (N_2877,N_2708,N_2706);
nand U2878 (N_2878,N_2797,N_2666);
nand U2879 (N_2879,N_2750,N_2676);
or U2880 (N_2880,N_2770,N_2692);
and U2881 (N_2881,N_2766,N_2640);
or U2882 (N_2882,N_2698,N_2776);
and U2883 (N_2883,N_2756,N_2673);
nand U2884 (N_2884,N_2688,N_2678);
nand U2885 (N_2885,N_2614,N_2709);
nor U2886 (N_2886,N_2622,N_2659);
or U2887 (N_2887,N_2768,N_2721);
xnor U2888 (N_2888,N_2694,N_2731);
and U2889 (N_2889,N_2755,N_2615);
and U2890 (N_2890,N_2609,N_2613);
or U2891 (N_2891,N_2665,N_2785);
and U2892 (N_2892,N_2730,N_2757);
nand U2893 (N_2893,N_2635,N_2737);
xnor U2894 (N_2894,N_2648,N_2604);
nor U2895 (N_2895,N_2661,N_2793);
or U2896 (N_2896,N_2697,N_2719);
xor U2897 (N_2897,N_2626,N_2779);
or U2898 (N_2898,N_2714,N_2611);
or U2899 (N_2899,N_2690,N_2734);
and U2900 (N_2900,N_2648,N_2650);
or U2901 (N_2901,N_2618,N_2642);
and U2902 (N_2902,N_2794,N_2603);
nand U2903 (N_2903,N_2718,N_2713);
nor U2904 (N_2904,N_2797,N_2682);
xnor U2905 (N_2905,N_2720,N_2685);
nand U2906 (N_2906,N_2731,N_2687);
or U2907 (N_2907,N_2799,N_2783);
or U2908 (N_2908,N_2644,N_2619);
and U2909 (N_2909,N_2641,N_2755);
or U2910 (N_2910,N_2615,N_2746);
or U2911 (N_2911,N_2634,N_2602);
and U2912 (N_2912,N_2661,N_2612);
and U2913 (N_2913,N_2601,N_2727);
and U2914 (N_2914,N_2797,N_2625);
or U2915 (N_2915,N_2761,N_2701);
xor U2916 (N_2916,N_2653,N_2627);
and U2917 (N_2917,N_2694,N_2730);
or U2918 (N_2918,N_2793,N_2680);
nor U2919 (N_2919,N_2685,N_2716);
or U2920 (N_2920,N_2671,N_2646);
or U2921 (N_2921,N_2650,N_2760);
and U2922 (N_2922,N_2691,N_2612);
nand U2923 (N_2923,N_2717,N_2621);
or U2924 (N_2924,N_2785,N_2727);
nand U2925 (N_2925,N_2722,N_2690);
nand U2926 (N_2926,N_2666,N_2693);
and U2927 (N_2927,N_2729,N_2660);
and U2928 (N_2928,N_2714,N_2650);
nand U2929 (N_2929,N_2680,N_2677);
nand U2930 (N_2930,N_2656,N_2700);
nor U2931 (N_2931,N_2648,N_2694);
nand U2932 (N_2932,N_2794,N_2763);
or U2933 (N_2933,N_2748,N_2724);
nand U2934 (N_2934,N_2682,N_2655);
and U2935 (N_2935,N_2703,N_2697);
nor U2936 (N_2936,N_2601,N_2797);
and U2937 (N_2937,N_2694,N_2610);
or U2938 (N_2938,N_2705,N_2728);
xor U2939 (N_2939,N_2607,N_2708);
nor U2940 (N_2940,N_2728,N_2794);
nand U2941 (N_2941,N_2659,N_2776);
nor U2942 (N_2942,N_2770,N_2719);
and U2943 (N_2943,N_2609,N_2768);
xor U2944 (N_2944,N_2696,N_2726);
xnor U2945 (N_2945,N_2676,N_2658);
and U2946 (N_2946,N_2724,N_2643);
nor U2947 (N_2947,N_2669,N_2715);
and U2948 (N_2948,N_2641,N_2735);
nor U2949 (N_2949,N_2695,N_2759);
xor U2950 (N_2950,N_2700,N_2778);
xor U2951 (N_2951,N_2684,N_2737);
nor U2952 (N_2952,N_2739,N_2715);
xnor U2953 (N_2953,N_2741,N_2656);
nor U2954 (N_2954,N_2629,N_2605);
xor U2955 (N_2955,N_2767,N_2617);
nor U2956 (N_2956,N_2757,N_2688);
or U2957 (N_2957,N_2756,N_2603);
xor U2958 (N_2958,N_2696,N_2759);
xor U2959 (N_2959,N_2762,N_2746);
and U2960 (N_2960,N_2748,N_2782);
nor U2961 (N_2961,N_2744,N_2769);
nand U2962 (N_2962,N_2778,N_2706);
and U2963 (N_2963,N_2781,N_2697);
and U2964 (N_2964,N_2696,N_2655);
xnor U2965 (N_2965,N_2677,N_2756);
and U2966 (N_2966,N_2601,N_2781);
nand U2967 (N_2967,N_2777,N_2610);
or U2968 (N_2968,N_2623,N_2799);
xnor U2969 (N_2969,N_2666,N_2741);
and U2970 (N_2970,N_2723,N_2660);
nor U2971 (N_2971,N_2614,N_2673);
or U2972 (N_2972,N_2699,N_2724);
nor U2973 (N_2973,N_2788,N_2743);
xor U2974 (N_2974,N_2650,N_2787);
xor U2975 (N_2975,N_2709,N_2760);
xnor U2976 (N_2976,N_2601,N_2658);
nand U2977 (N_2977,N_2624,N_2641);
nor U2978 (N_2978,N_2797,N_2777);
nor U2979 (N_2979,N_2764,N_2696);
nor U2980 (N_2980,N_2765,N_2613);
or U2981 (N_2981,N_2688,N_2625);
or U2982 (N_2982,N_2632,N_2722);
nand U2983 (N_2983,N_2723,N_2629);
nand U2984 (N_2984,N_2766,N_2745);
nand U2985 (N_2985,N_2779,N_2676);
xor U2986 (N_2986,N_2654,N_2773);
or U2987 (N_2987,N_2673,N_2639);
and U2988 (N_2988,N_2716,N_2787);
nor U2989 (N_2989,N_2723,N_2700);
or U2990 (N_2990,N_2767,N_2672);
nand U2991 (N_2991,N_2690,N_2665);
nand U2992 (N_2992,N_2695,N_2665);
xor U2993 (N_2993,N_2748,N_2618);
nor U2994 (N_2994,N_2775,N_2764);
and U2995 (N_2995,N_2612,N_2626);
xor U2996 (N_2996,N_2711,N_2732);
or U2997 (N_2997,N_2725,N_2779);
nor U2998 (N_2998,N_2742,N_2712);
or U2999 (N_2999,N_2782,N_2672);
xor U3000 (N_3000,N_2821,N_2804);
nand U3001 (N_3001,N_2946,N_2928);
nand U3002 (N_3002,N_2919,N_2802);
nor U3003 (N_3003,N_2904,N_2973);
nand U3004 (N_3004,N_2996,N_2962);
nand U3005 (N_3005,N_2944,N_2922);
nor U3006 (N_3006,N_2947,N_2980);
nand U3007 (N_3007,N_2903,N_2851);
and U3008 (N_3008,N_2842,N_2881);
or U3009 (N_3009,N_2975,N_2987);
and U3010 (N_3010,N_2915,N_2895);
or U3011 (N_3011,N_2898,N_2989);
nand U3012 (N_3012,N_2817,N_2805);
or U3013 (N_3013,N_2809,N_2887);
nor U3014 (N_3014,N_2907,N_2905);
and U3015 (N_3015,N_2968,N_2844);
and U3016 (N_3016,N_2900,N_2872);
nor U3017 (N_3017,N_2998,N_2933);
and U3018 (N_3018,N_2825,N_2974);
nand U3019 (N_3019,N_2967,N_2826);
xor U3020 (N_3020,N_2934,N_2888);
and U3021 (N_3021,N_2880,N_2819);
or U3022 (N_3022,N_2840,N_2852);
xnor U3023 (N_3023,N_2927,N_2889);
nand U3024 (N_3024,N_2942,N_2836);
xor U3025 (N_3025,N_2866,N_2891);
xnor U3026 (N_3026,N_2961,N_2929);
nor U3027 (N_3027,N_2829,N_2976);
xnor U3028 (N_3028,N_2984,N_2909);
xor U3029 (N_3029,N_2988,N_2955);
and U3030 (N_3030,N_2878,N_2814);
or U3031 (N_3031,N_2867,N_2820);
nor U3032 (N_3032,N_2859,N_2913);
xnor U3033 (N_3033,N_2827,N_2876);
xor U3034 (N_3034,N_2992,N_2953);
or U3035 (N_3035,N_2812,N_2991);
xor U3036 (N_3036,N_2847,N_2983);
xnor U3037 (N_3037,N_2830,N_2849);
nor U3038 (N_3038,N_2808,N_2985);
and U3039 (N_3039,N_2969,N_2943);
or U3040 (N_3040,N_2924,N_2893);
and U3041 (N_3041,N_2885,N_2865);
and U3042 (N_3042,N_2853,N_2884);
xor U3043 (N_3043,N_2896,N_2917);
nor U3044 (N_3044,N_2910,N_2838);
nor U3045 (N_3045,N_2902,N_2939);
xor U3046 (N_3046,N_2930,N_2937);
nor U3047 (N_3047,N_2803,N_2828);
xnor U3048 (N_3048,N_2890,N_2824);
or U3049 (N_3049,N_2861,N_2897);
and U3050 (N_3050,N_2850,N_2858);
xor U3051 (N_3051,N_2877,N_2918);
or U3052 (N_3052,N_2822,N_2870);
and U3053 (N_3053,N_2823,N_2843);
or U3054 (N_3054,N_2835,N_2994);
and U3055 (N_3055,N_2874,N_2908);
or U3056 (N_3056,N_2920,N_2945);
xor U3057 (N_3057,N_2949,N_2837);
nand U3058 (N_3058,N_2818,N_2883);
nor U3059 (N_3059,N_2979,N_2990);
nand U3060 (N_3060,N_2834,N_2954);
nor U3061 (N_3061,N_2957,N_2906);
nor U3062 (N_3062,N_2894,N_2940);
or U3063 (N_3063,N_2882,N_2841);
and U3064 (N_3064,N_2916,N_2963);
xnor U3065 (N_3065,N_2854,N_2811);
and U3066 (N_3066,N_2923,N_2921);
and U3067 (N_3067,N_2952,N_2936);
and U3068 (N_3068,N_2958,N_2868);
and U3069 (N_3069,N_2999,N_2960);
nor U3070 (N_3070,N_2997,N_2875);
nor U3071 (N_3071,N_2869,N_2950);
nor U3072 (N_3072,N_2966,N_2807);
xor U3073 (N_3073,N_2879,N_2977);
nand U3074 (N_3074,N_2951,N_2982);
and U3075 (N_3075,N_2899,N_2948);
nor U3076 (N_3076,N_2970,N_2816);
nor U3077 (N_3077,N_2956,N_2932);
nand U3078 (N_3078,N_2855,N_2813);
nor U3079 (N_3079,N_2925,N_2965);
and U3080 (N_3080,N_2831,N_2862);
and U3081 (N_3081,N_2857,N_2860);
and U3082 (N_3082,N_2995,N_2901);
or U3083 (N_3083,N_2873,N_2832);
nor U3084 (N_3084,N_2846,N_2964);
nor U3085 (N_3085,N_2833,N_2935);
and U3086 (N_3086,N_2886,N_2871);
xor U3087 (N_3087,N_2911,N_2848);
or U3088 (N_3088,N_2864,N_2993);
nand U3089 (N_3089,N_2845,N_2931);
nor U3090 (N_3090,N_2972,N_2806);
nand U3091 (N_3091,N_2986,N_2801);
or U3092 (N_3092,N_2938,N_2978);
or U3093 (N_3093,N_2863,N_2815);
nor U3094 (N_3094,N_2981,N_2941);
xnor U3095 (N_3095,N_2839,N_2971);
and U3096 (N_3096,N_2800,N_2926);
nand U3097 (N_3097,N_2914,N_2912);
nand U3098 (N_3098,N_2892,N_2856);
xor U3099 (N_3099,N_2959,N_2810);
and U3100 (N_3100,N_2903,N_2924);
and U3101 (N_3101,N_2898,N_2829);
or U3102 (N_3102,N_2993,N_2909);
nor U3103 (N_3103,N_2955,N_2846);
or U3104 (N_3104,N_2892,N_2833);
nand U3105 (N_3105,N_2840,N_2937);
nand U3106 (N_3106,N_2984,N_2954);
nor U3107 (N_3107,N_2945,N_2997);
xnor U3108 (N_3108,N_2998,N_2849);
xnor U3109 (N_3109,N_2997,N_2811);
or U3110 (N_3110,N_2968,N_2916);
nand U3111 (N_3111,N_2899,N_2939);
xor U3112 (N_3112,N_2824,N_2866);
or U3113 (N_3113,N_2996,N_2800);
xor U3114 (N_3114,N_2914,N_2813);
nand U3115 (N_3115,N_2933,N_2813);
or U3116 (N_3116,N_2829,N_2980);
or U3117 (N_3117,N_2846,N_2909);
nor U3118 (N_3118,N_2825,N_2949);
nor U3119 (N_3119,N_2811,N_2960);
or U3120 (N_3120,N_2988,N_2934);
nand U3121 (N_3121,N_2860,N_2844);
nor U3122 (N_3122,N_2932,N_2925);
xnor U3123 (N_3123,N_2841,N_2924);
xor U3124 (N_3124,N_2917,N_2967);
nand U3125 (N_3125,N_2847,N_2915);
nor U3126 (N_3126,N_2947,N_2998);
nor U3127 (N_3127,N_2830,N_2887);
nor U3128 (N_3128,N_2976,N_2951);
and U3129 (N_3129,N_2967,N_2906);
xor U3130 (N_3130,N_2934,N_2937);
xor U3131 (N_3131,N_2804,N_2996);
and U3132 (N_3132,N_2966,N_2923);
nand U3133 (N_3133,N_2969,N_2823);
nand U3134 (N_3134,N_2899,N_2804);
and U3135 (N_3135,N_2957,N_2919);
nand U3136 (N_3136,N_2862,N_2828);
and U3137 (N_3137,N_2969,N_2959);
and U3138 (N_3138,N_2987,N_2807);
nor U3139 (N_3139,N_2819,N_2910);
nor U3140 (N_3140,N_2976,N_2991);
or U3141 (N_3141,N_2945,N_2862);
or U3142 (N_3142,N_2976,N_2882);
or U3143 (N_3143,N_2932,N_2886);
nand U3144 (N_3144,N_2947,N_2864);
or U3145 (N_3145,N_2935,N_2817);
or U3146 (N_3146,N_2949,N_2905);
xnor U3147 (N_3147,N_2864,N_2805);
or U3148 (N_3148,N_2904,N_2908);
xnor U3149 (N_3149,N_2946,N_2951);
or U3150 (N_3150,N_2874,N_2910);
and U3151 (N_3151,N_2840,N_2961);
and U3152 (N_3152,N_2919,N_2811);
nand U3153 (N_3153,N_2963,N_2999);
nor U3154 (N_3154,N_2825,N_2861);
and U3155 (N_3155,N_2897,N_2952);
or U3156 (N_3156,N_2970,N_2984);
nor U3157 (N_3157,N_2818,N_2974);
or U3158 (N_3158,N_2892,N_2830);
nor U3159 (N_3159,N_2816,N_2843);
nor U3160 (N_3160,N_2886,N_2942);
nor U3161 (N_3161,N_2997,N_2861);
xor U3162 (N_3162,N_2909,N_2879);
xnor U3163 (N_3163,N_2888,N_2964);
xor U3164 (N_3164,N_2915,N_2932);
nor U3165 (N_3165,N_2980,N_2881);
xor U3166 (N_3166,N_2847,N_2974);
nor U3167 (N_3167,N_2813,N_2994);
and U3168 (N_3168,N_2864,N_2833);
nand U3169 (N_3169,N_2876,N_2959);
nand U3170 (N_3170,N_2839,N_2899);
nand U3171 (N_3171,N_2880,N_2891);
and U3172 (N_3172,N_2852,N_2899);
or U3173 (N_3173,N_2828,N_2826);
and U3174 (N_3174,N_2841,N_2805);
nor U3175 (N_3175,N_2907,N_2939);
nor U3176 (N_3176,N_2990,N_2842);
nor U3177 (N_3177,N_2958,N_2803);
nor U3178 (N_3178,N_2826,N_2913);
or U3179 (N_3179,N_2888,N_2961);
nor U3180 (N_3180,N_2963,N_2951);
xnor U3181 (N_3181,N_2925,N_2943);
xnor U3182 (N_3182,N_2973,N_2985);
xnor U3183 (N_3183,N_2937,N_2939);
xnor U3184 (N_3184,N_2876,N_2801);
xnor U3185 (N_3185,N_2951,N_2972);
nand U3186 (N_3186,N_2826,N_2874);
or U3187 (N_3187,N_2865,N_2955);
or U3188 (N_3188,N_2839,N_2916);
nand U3189 (N_3189,N_2922,N_2930);
nor U3190 (N_3190,N_2999,N_2906);
nand U3191 (N_3191,N_2829,N_2950);
nor U3192 (N_3192,N_2858,N_2835);
and U3193 (N_3193,N_2965,N_2908);
nand U3194 (N_3194,N_2883,N_2891);
or U3195 (N_3195,N_2863,N_2884);
and U3196 (N_3196,N_2919,N_2825);
xor U3197 (N_3197,N_2804,N_2986);
xnor U3198 (N_3198,N_2976,N_2919);
and U3199 (N_3199,N_2887,N_2958);
xor U3200 (N_3200,N_3139,N_3063);
nor U3201 (N_3201,N_3110,N_3055);
nand U3202 (N_3202,N_3065,N_3004);
and U3203 (N_3203,N_3057,N_3198);
nand U3204 (N_3204,N_3126,N_3084);
or U3205 (N_3205,N_3144,N_3083);
or U3206 (N_3206,N_3094,N_3184);
or U3207 (N_3207,N_3115,N_3194);
nand U3208 (N_3208,N_3095,N_3145);
or U3209 (N_3209,N_3030,N_3005);
nor U3210 (N_3210,N_3120,N_3166);
nand U3211 (N_3211,N_3012,N_3069);
or U3212 (N_3212,N_3097,N_3066);
nand U3213 (N_3213,N_3013,N_3134);
or U3214 (N_3214,N_3190,N_3053);
xor U3215 (N_3215,N_3018,N_3046);
nor U3216 (N_3216,N_3143,N_3040);
xnor U3217 (N_3217,N_3150,N_3045);
nor U3218 (N_3218,N_3191,N_3182);
nand U3219 (N_3219,N_3161,N_3170);
xor U3220 (N_3220,N_3003,N_3148);
xnor U3221 (N_3221,N_3196,N_3147);
xor U3222 (N_3222,N_3071,N_3075);
nor U3223 (N_3223,N_3105,N_3060);
nand U3224 (N_3224,N_3033,N_3059);
or U3225 (N_3225,N_3101,N_3132);
xnor U3226 (N_3226,N_3099,N_3038);
and U3227 (N_3227,N_3189,N_3107);
nor U3228 (N_3228,N_3108,N_3141);
or U3229 (N_3229,N_3049,N_3006);
and U3230 (N_3230,N_3086,N_3017);
and U3231 (N_3231,N_3195,N_3015);
nand U3232 (N_3232,N_3137,N_3140);
or U3233 (N_3233,N_3167,N_3032);
nand U3234 (N_3234,N_3163,N_3106);
xnor U3235 (N_3235,N_3085,N_3173);
nor U3236 (N_3236,N_3149,N_3064);
xnor U3237 (N_3237,N_3061,N_3048);
nor U3238 (N_3238,N_3125,N_3178);
nor U3239 (N_3239,N_3118,N_3024);
nand U3240 (N_3240,N_3121,N_3042);
and U3241 (N_3241,N_3089,N_3010);
xor U3242 (N_3242,N_3181,N_3192);
nand U3243 (N_3243,N_3029,N_3093);
or U3244 (N_3244,N_3043,N_3112);
nand U3245 (N_3245,N_3183,N_3020);
and U3246 (N_3246,N_3025,N_3082);
or U3247 (N_3247,N_3026,N_3111);
nand U3248 (N_3248,N_3130,N_3186);
nand U3249 (N_3249,N_3138,N_3103);
and U3250 (N_3250,N_3171,N_3028);
and U3251 (N_3251,N_3176,N_3164);
nor U3252 (N_3252,N_3136,N_3152);
or U3253 (N_3253,N_3068,N_3062);
nor U3254 (N_3254,N_3039,N_3016);
and U3255 (N_3255,N_3096,N_3022);
xnor U3256 (N_3256,N_3188,N_3153);
nand U3257 (N_3257,N_3133,N_3021);
and U3258 (N_3258,N_3199,N_3169);
nand U3259 (N_3259,N_3142,N_3154);
or U3260 (N_3260,N_3113,N_3056);
nor U3261 (N_3261,N_3174,N_3014);
nand U3262 (N_3262,N_3011,N_3168);
nor U3263 (N_3263,N_3116,N_3102);
xnor U3264 (N_3264,N_3044,N_3135);
nor U3265 (N_3265,N_3009,N_3114);
xnor U3266 (N_3266,N_3129,N_3052);
or U3267 (N_3267,N_3160,N_3002);
nor U3268 (N_3268,N_3159,N_3104);
nor U3269 (N_3269,N_3180,N_3175);
xor U3270 (N_3270,N_3041,N_3054);
or U3271 (N_3271,N_3179,N_3151);
and U3272 (N_3272,N_3034,N_3008);
nand U3273 (N_3273,N_3070,N_3119);
or U3274 (N_3274,N_3127,N_3051);
nor U3275 (N_3275,N_3019,N_3100);
xnor U3276 (N_3276,N_3117,N_3162);
xnor U3277 (N_3277,N_3185,N_3023);
xnor U3278 (N_3278,N_3079,N_3078);
or U3279 (N_3279,N_3007,N_3158);
xor U3280 (N_3280,N_3155,N_3172);
and U3281 (N_3281,N_3000,N_3087);
xor U3282 (N_3282,N_3067,N_3073);
nor U3283 (N_3283,N_3035,N_3122);
nand U3284 (N_3284,N_3128,N_3131);
nor U3285 (N_3285,N_3074,N_3058);
nand U3286 (N_3286,N_3193,N_3090);
or U3287 (N_3287,N_3036,N_3177);
nand U3288 (N_3288,N_3091,N_3001);
nor U3289 (N_3289,N_3080,N_3027);
or U3290 (N_3290,N_3146,N_3088);
or U3291 (N_3291,N_3081,N_3077);
nand U3292 (N_3292,N_3092,N_3050);
nor U3293 (N_3293,N_3124,N_3197);
and U3294 (N_3294,N_3109,N_3047);
nor U3295 (N_3295,N_3123,N_3165);
and U3296 (N_3296,N_3156,N_3031);
nand U3297 (N_3297,N_3187,N_3157);
xnor U3298 (N_3298,N_3098,N_3072);
and U3299 (N_3299,N_3037,N_3076);
nor U3300 (N_3300,N_3112,N_3143);
or U3301 (N_3301,N_3141,N_3085);
or U3302 (N_3302,N_3133,N_3057);
nor U3303 (N_3303,N_3031,N_3198);
nand U3304 (N_3304,N_3008,N_3098);
and U3305 (N_3305,N_3141,N_3090);
nor U3306 (N_3306,N_3076,N_3150);
nand U3307 (N_3307,N_3131,N_3059);
and U3308 (N_3308,N_3131,N_3140);
and U3309 (N_3309,N_3140,N_3022);
or U3310 (N_3310,N_3011,N_3105);
and U3311 (N_3311,N_3091,N_3176);
nand U3312 (N_3312,N_3103,N_3185);
or U3313 (N_3313,N_3024,N_3137);
xor U3314 (N_3314,N_3179,N_3012);
and U3315 (N_3315,N_3182,N_3081);
or U3316 (N_3316,N_3178,N_3051);
or U3317 (N_3317,N_3083,N_3180);
xor U3318 (N_3318,N_3044,N_3195);
nand U3319 (N_3319,N_3199,N_3004);
or U3320 (N_3320,N_3179,N_3159);
or U3321 (N_3321,N_3020,N_3182);
nor U3322 (N_3322,N_3124,N_3091);
or U3323 (N_3323,N_3183,N_3111);
nand U3324 (N_3324,N_3014,N_3049);
and U3325 (N_3325,N_3023,N_3089);
nor U3326 (N_3326,N_3149,N_3016);
and U3327 (N_3327,N_3134,N_3045);
nand U3328 (N_3328,N_3032,N_3094);
or U3329 (N_3329,N_3159,N_3154);
xor U3330 (N_3330,N_3088,N_3116);
nand U3331 (N_3331,N_3022,N_3093);
nor U3332 (N_3332,N_3153,N_3040);
or U3333 (N_3333,N_3159,N_3043);
and U3334 (N_3334,N_3173,N_3026);
nor U3335 (N_3335,N_3134,N_3117);
and U3336 (N_3336,N_3040,N_3193);
xor U3337 (N_3337,N_3125,N_3182);
nand U3338 (N_3338,N_3012,N_3169);
or U3339 (N_3339,N_3094,N_3081);
or U3340 (N_3340,N_3070,N_3159);
nor U3341 (N_3341,N_3102,N_3051);
nor U3342 (N_3342,N_3162,N_3182);
or U3343 (N_3343,N_3155,N_3180);
nor U3344 (N_3344,N_3072,N_3170);
or U3345 (N_3345,N_3199,N_3011);
xnor U3346 (N_3346,N_3190,N_3073);
nor U3347 (N_3347,N_3106,N_3169);
and U3348 (N_3348,N_3149,N_3191);
xnor U3349 (N_3349,N_3021,N_3000);
nor U3350 (N_3350,N_3172,N_3039);
and U3351 (N_3351,N_3197,N_3060);
nand U3352 (N_3352,N_3043,N_3101);
and U3353 (N_3353,N_3184,N_3102);
nand U3354 (N_3354,N_3091,N_3098);
xor U3355 (N_3355,N_3193,N_3125);
and U3356 (N_3356,N_3153,N_3063);
and U3357 (N_3357,N_3010,N_3144);
nor U3358 (N_3358,N_3178,N_3162);
nand U3359 (N_3359,N_3016,N_3165);
and U3360 (N_3360,N_3199,N_3160);
xnor U3361 (N_3361,N_3002,N_3142);
and U3362 (N_3362,N_3167,N_3104);
or U3363 (N_3363,N_3075,N_3158);
nand U3364 (N_3364,N_3147,N_3154);
or U3365 (N_3365,N_3073,N_3157);
and U3366 (N_3366,N_3135,N_3115);
nor U3367 (N_3367,N_3070,N_3154);
and U3368 (N_3368,N_3112,N_3095);
or U3369 (N_3369,N_3116,N_3086);
or U3370 (N_3370,N_3099,N_3040);
or U3371 (N_3371,N_3094,N_3153);
and U3372 (N_3372,N_3122,N_3123);
or U3373 (N_3373,N_3133,N_3151);
nand U3374 (N_3374,N_3024,N_3104);
xnor U3375 (N_3375,N_3123,N_3097);
nor U3376 (N_3376,N_3035,N_3044);
xor U3377 (N_3377,N_3053,N_3130);
nand U3378 (N_3378,N_3159,N_3072);
nor U3379 (N_3379,N_3088,N_3147);
and U3380 (N_3380,N_3114,N_3122);
nor U3381 (N_3381,N_3192,N_3088);
xnor U3382 (N_3382,N_3135,N_3031);
xnor U3383 (N_3383,N_3091,N_3093);
and U3384 (N_3384,N_3142,N_3143);
and U3385 (N_3385,N_3091,N_3083);
nor U3386 (N_3386,N_3011,N_3131);
nor U3387 (N_3387,N_3112,N_3144);
xor U3388 (N_3388,N_3168,N_3137);
xor U3389 (N_3389,N_3006,N_3051);
nand U3390 (N_3390,N_3077,N_3066);
or U3391 (N_3391,N_3112,N_3150);
xor U3392 (N_3392,N_3112,N_3096);
xor U3393 (N_3393,N_3188,N_3113);
nor U3394 (N_3394,N_3025,N_3077);
nand U3395 (N_3395,N_3190,N_3011);
nor U3396 (N_3396,N_3191,N_3058);
and U3397 (N_3397,N_3045,N_3061);
or U3398 (N_3398,N_3047,N_3149);
xnor U3399 (N_3399,N_3060,N_3096);
nor U3400 (N_3400,N_3399,N_3289);
or U3401 (N_3401,N_3394,N_3298);
or U3402 (N_3402,N_3297,N_3328);
nor U3403 (N_3403,N_3398,N_3283);
or U3404 (N_3404,N_3301,N_3229);
nor U3405 (N_3405,N_3359,N_3288);
xnor U3406 (N_3406,N_3380,N_3210);
and U3407 (N_3407,N_3291,N_3296);
nand U3408 (N_3408,N_3323,N_3269);
nor U3409 (N_3409,N_3395,N_3276);
xor U3410 (N_3410,N_3389,N_3256);
or U3411 (N_3411,N_3260,N_3355);
nand U3412 (N_3412,N_3218,N_3209);
nor U3413 (N_3413,N_3384,N_3360);
and U3414 (N_3414,N_3266,N_3207);
or U3415 (N_3415,N_3300,N_3241);
xnor U3416 (N_3416,N_3373,N_3293);
and U3417 (N_3417,N_3315,N_3237);
xor U3418 (N_3418,N_3327,N_3273);
nor U3419 (N_3419,N_3324,N_3282);
xnor U3420 (N_3420,N_3208,N_3333);
or U3421 (N_3421,N_3294,N_3281);
and U3422 (N_3422,N_3284,N_3310);
nand U3423 (N_3423,N_3224,N_3236);
or U3424 (N_3424,N_3306,N_3357);
or U3425 (N_3425,N_3356,N_3215);
xor U3426 (N_3426,N_3325,N_3312);
nor U3427 (N_3427,N_3397,N_3279);
nor U3428 (N_3428,N_3319,N_3308);
or U3429 (N_3429,N_3219,N_3261);
and U3430 (N_3430,N_3352,N_3263);
nor U3431 (N_3431,N_3383,N_3204);
nand U3432 (N_3432,N_3311,N_3249);
nand U3433 (N_3433,N_3390,N_3363);
xor U3434 (N_3434,N_3347,N_3235);
and U3435 (N_3435,N_3332,N_3223);
xnor U3436 (N_3436,N_3232,N_3382);
nand U3437 (N_3437,N_3386,N_3330);
or U3438 (N_3438,N_3239,N_3372);
nand U3439 (N_3439,N_3346,N_3231);
nand U3440 (N_3440,N_3287,N_3268);
or U3441 (N_3441,N_3370,N_3216);
or U3442 (N_3442,N_3278,N_3248);
and U3443 (N_3443,N_3375,N_3320);
or U3444 (N_3444,N_3307,N_3392);
and U3445 (N_3445,N_3313,N_3343);
xor U3446 (N_3446,N_3362,N_3331);
and U3447 (N_3447,N_3227,N_3336);
nor U3448 (N_3448,N_3304,N_3212);
xor U3449 (N_3449,N_3234,N_3228);
or U3450 (N_3450,N_3337,N_3225);
nand U3451 (N_3451,N_3246,N_3230);
or U3452 (N_3452,N_3340,N_3366);
or U3453 (N_3453,N_3361,N_3271);
xnor U3454 (N_3454,N_3348,N_3240);
xnor U3455 (N_3455,N_3254,N_3316);
or U3456 (N_3456,N_3314,N_3290);
nand U3457 (N_3457,N_3201,N_3341);
or U3458 (N_3458,N_3322,N_3247);
xnor U3459 (N_3459,N_3303,N_3299);
nand U3460 (N_3460,N_3329,N_3335);
and U3461 (N_3461,N_3272,N_3326);
or U3462 (N_3462,N_3391,N_3213);
or U3463 (N_3463,N_3365,N_3345);
nor U3464 (N_3464,N_3262,N_3338);
and U3465 (N_3465,N_3385,N_3253);
nor U3466 (N_3466,N_3270,N_3233);
or U3467 (N_3467,N_3351,N_3358);
nand U3468 (N_3468,N_3377,N_3378);
xor U3469 (N_3469,N_3264,N_3396);
xnor U3470 (N_3470,N_3344,N_3221);
or U3471 (N_3471,N_3243,N_3214);
xnor U3472 (N_3472,N_3202,N_3203);
and U3473 (N_3473,N_3318,N_3244);
and U3474 (N_3474,N_3251,N_3286);
or U3475 (N_3475,N_3242,N_3302);
or U3476 (N_3476,N_3280,N_3376);
and U3477 (N_3477,N_3317,N_3220);
xor U3478 (N_3478,N_3374,N_3222);
nor U3479 (N_3479,N_3274,N_3259);
nand U3480 (N_3480,N_3250,N_3339);
nor U3481 (N_3481,N_3388,N_3381);
xor U3482 (N_3482,N_3368,N_3371);
nand U3483 (N_3483,N_3211,N_3217);
nor U3484 (N_3484,N_3354,N_3285);
or U3485 (N_3485,N_3353,N_3305);
nor U3486 (N_3486,N_3292,N_3200);
nor U3487 (N_3487,N_3252,N_3309);
nand U3488 (N_3488,N_3226,N_3379);
or U3489 (N_3489,N_3350,N_3295);
or U3490 (N_3490,N_3369,N_3342);
or U3491 (N_3491,N_3364,N_3267);
and U3492 (N_3492,N_3349,N_3387);
and U3493 (N_3493,N_3393,N_3238);
or U3494 (N_3494,N_3367,N_3245);
xor U3495 (N_3495,N_3275,N_3257);
xor U3496 (N_3496,N_3206,N_3277);
nor U3497 (N_3497,N_3205,N_3321);
and U3498 (N_3498,N_3265,N_3255);
nor U3499 (N_3499,N_3334,N_3258);
or U3500 (N_3500,N_3388,N_3259);
xor U3501 (N_3501,N_3302,N_3227);
or U3502 (N_3502,N_3280,N_3314);
and U3503 (N_3503,N_3308,N_3257);
xor U3504 (N_3504,N_3282,N_3218);
or U3505 (N_3505,N_3335,N_3271);
or U3506 (N_3506,N_3327,N_3306);
nand U3507 (N_3507,N_3260,N_3331);
nor U3508 (N_3508,N_3283,N_3345);
xnor U3509 (N_3509,N_3315,N_3343);
nor U3510 (N_3510,N_3295,N_3204);
nor U3511 (N_3511,N_3358,N_3220);
xor U3512 (N_3512,N_3294,N_3312);
nor U3513 (N_3513,N_3304,N_3250);
and U3514 (N_3514,N_3261,N_3280);
nand U3515 (N_3515,N_3369,N_3356);
xnor U3516 (N_3516,N_3376,N_3266);
xnor U3517 (N_3517,N_3348,N_3377);
and U3518 (N_3518,N_3276,N_3305);
xor U3519 (N_3519,N_3263,N_3333);
and U3520 (N_3520,N_3318,N_3316);
nand U3521 (N_3521,N_3213,N_3361);
xor U3522 (N_3522,N_3236,N_3275);
and U3523 (N_3523,N_3236,N_3348);
or U3524 (N_3524,N_3359,N_3376);
nor U3525 (N_3525,N_3274,N_3340);
nand U3526 (N_3526,N_3368,N_3310);
nor U3527 (N_3527,N_3279,N_3358);
nand U3528 (N_3528,N_3356,N_3216);
and U3529 (N_3529,N_3297,N_3269);
nand U3530 (N_3530,N_3254,N_3363);
or U3531 (N_3531,N_3245,N_3260);
xor U3532 (N_3532,N_3397,N_3242);
or U3533 (N_3533,N_3343,N_3399);
nor U3534 (N_3534,N_3320,N_3324);
and U3535 (N_3535,N_3263,N_3329);
and U3536 (N_3536,N_3313,N_3237);
nor U3537 (N_3537,N_3360,N_3383);
and U3538 (N_3538,N_3297,N_3216);
or U3539 (N_3539,N_3327,N_3229);
xor U3540 (N_3540,N_3207,N_3385);
or U3541 (N_3541,N_3220,N_3255);
nand U3542 (N_3542,N_3211,N_3283);
nor U3543 (N_3543,N_3344,N_3213);
xor U3544 (N_3544,N_3331,N_3241);
xor U3545 (N_3545,N_3347,N_3249);
nand U3546 (N_3546,N_3308,N_3341);
nor U3547 (N_3547,N_3258,N_3255);
nand U3548 (N_3548,N_3244,N_3371);
or U3549 (N_3549,N_3280,N_3342);
xor U3550 (N_3550,N_3297,N_3301);
nand U3551 (N_3551,N_3310,N_3369);
nor U3552 (N_3552,N_3246,N_3397);
and U3553 (N_3553,N_3272,N_3255);
nor U3554 (N_3554,N_3221,N_3305);
or U3555 (N_3555,N_3398,N_3245);
xnor U3556 (N_3556,N_3252,N_3206);
and U3557 (N_3557,N_3378,N_3208);
or U3558 (N_3558,N_3330,N_3230);
xor U3559 (N_3559,N_3357,N_3288);
or U3560 (N_3560,N_3308,N_3306);
or U3561 (N_3561,N_3364,N_3272);
nand U3562 (N_3562,N_3238,N_3281);
nand U3563 (N_3563,N_3339,N_3322);
nand U3564 (N_3564,N_3234,N_3311);
nor U3565 (N_3565,N_3253,N_3313);
xnor U3566 (N_3566,N_3330,N_3318);
nand U3567 (N_3567,N_3337,N_3255);
or U3568 (N_3568,N_3379,N_3311);
or U3569 (N_3569,N_3207,N_3367);
or U3570 (N_3570,N_3338,N_3365);
and U3571 (N_3571,N_3397,N_3214);
nand U3572 (N_3572,N_3346,N_3345);
nand U3573 (N_3573,N_3243,N_3358);
nand U3574 (N_3574,N_3206,N_3320);
nand U3575 (N_3575,N_3260,N_3347);
or U3576 (N_3576,N_3319,N_3221);
nand U3577 (N_3577,N_3240,N_3373);
xnor U3578 (N_3578,N_3395,N_3289);
nand U3579 (N_3579,N_3390,N_3304);
and U3580 (N_3580,N_3225,N_3235);
nor U3581 (N_3581,N_3233,N_3201);
nor U3582 (N_3582,N_3364,N_3329);
or U3583 (N_3583,N_3386,N_3366);
xnor U3584 (N_3584,N_3390,N_3344);
nor U3585 (N_3585,N_3385,N_3292);
or U3586 (N_3586,N_3280,N_3350);
nor U3587 (N_3587,N_3330,N_3346);
nor U3588 (N_3588,N_3249,N_3282);
or U3589 (N_3589,N_3290,N_3388);
and U3590 (N_3590,N_3299,N_3255);
and U3591 (N_3591,N_3373,N_3257);
nor U3592 (N_3592,N_3229,N_3386);
nand U3593 (N_3593,N_3325,N_3349);
nor U3594 (N_3594,N_3345,N_3337);
xnor U3595 (N_3595,N_3206,N_3282);
nand U3596 (N_3596,N_3330,N_3263);
nand U3597 (N_3597,N_3377,N_3336);
nor U3598 (N_3598,N_3396,N_3256);
or U3599 (N_3599,N_3293,N_3291);
and U3600 (N_3600,N_3553,N_3506);
nand U3601 (N_3601,N_3444,N_3571);
nor U3602 (N_3602,N_3466,N_3418);
xnor U3603 (N_3603,N_3591,N_3438);
or U3604 (N_3604,N_3523,N_3400);
or U3605 (N_3605,N_3423,N_3452);
nor U3606 (N_3606,N_3533,N_3589);
or U3607 (N_3607,N_3535,N_3541);
nor U3608 (N_3608,N_3585,N_3486);
xnor U3609 (N_3609,N_3515,N_3590);
nand U3610 (N_3610,N_3478,N_3410);
and U3611 (N_3611,N_3599,N_3443);
nand U3612 (N_3612,N_3419,N_3517);
or U3613 (N_3613,N_3538,N_3522);
nor U3614 (N_3614,N_3448,N_3406);
nor U3615 (N_3615,N_3567,N_3560);
xor U3616 (N_3616,N_3471,N_3507);
or U3617 (N_3617,N_3526,N_3453);
nor U3618 (N_3618,N_3436,N_3488);
and U3619 (N_3619,N_3430,N_3598);
xor U3620 (N_3620,N_3404,N_3451);
nand U3621 (N_3621,N_3556,N_3569);
xor U3622 (N_3622,N_3536,N_3501);
or U3623 (N_3623,N_3421,N_3498);
or U3624 (N_3624,N_3458,N_3477);
or U3625 (N_3625,N_3579,N_3532);
nand U3626 (N_3626,N_3414,N_3425);
xor U3627 (N_3627,N_3597,N_3409);
nor U3628 (N_3628,N_3485,N_3540);
and U3629 (N_3629,N_3516,N_3530);
and U3630 (N_3630,N_3461,N_3565);
nand U3631 (N_3631,N_3401,N_3415);
nand U3632 (N_3632,N_3519,N_3417);
nand U3633 (N_3633,N_3489,N_3482);
nor U3634 (N_3634,N_3480,N_3475);
and U3635 (N_3635,N_3426,N_3509);
nand U3636 (N_3636,N_3446,N_3572);
or U3637 (N_3637,N_3542,N_3462);
and U3638 (N_3638,N_3432,N_3441);
or U3639 (N_3639,N_3594,N_3576);
xnor U3640 (N_3640,N_3456,N_3412);
and U3641 (N_3641,N_3447,N_3586);
nand U3642 (N_3642,N_3468,N_3545);
nand U3643 (N_3643,N_3557,N_3513);
or U3644 (N_3644,N_3483,N_3543);
nand U3645 (N_3645,N_3550,N_3583);
and U3646 (N_3646,N_3472,N_3445);
nor U3647 (N_3647,N_3499,N_3424);
nor U3648 (N_3648,N_3484,N_3558);
nor U3649 (N_3649,N_3492,N_3577);
and U3650 (N_3650,N_3524,N_3405);
or U3651 (N_3651,N_3511,N_3407);
or U3652 (N_3652,N_3502,N_3470);
or U3653 (N_3653,N_3559,N_3491);
nand U3654 (N_3654,N_3433,N_3527);
nand U3655 (N_3655,N_3518,N_3463);
or U3656 (N_3656,N_3514,N_3587);
nand U3657 (N_3657,N_3460,N_3497);
nand U3658 (N_3658,N_3490,N_3549);
xnor U3659 (N_3659,N_3568,N_3493);
nand U3660 (N_3660,N_3544,N_3496);
or U3661 (N_3661,N_3429,N_3531);
nand U3662 (N_3662,N_3495,N_3582);
xor U3663 (N_3663,N_3563,N_3520);
nor U3664 (N_3664,N_3529,N_3505);
or U3665 (N_3665,N_3434,N_3442);
or U3666 (N_3666,N_3416,N_3469);
xnor U3667 (N_3667,N_3494,N_3413);
xor U3668 (N_3668,N_3573,N_3457);
nor U3669 (N_3669,N_3578,N_3454);
nand U3670 (N_3670,N_3566,N_3440);
nor U3671 (N_3671,N_3510,N_3439);
or U3672 (N_3672,N_3500,N_3588);
nor U3673 (N_3673,N_3593,N_3508);
nand U3674 (N_3674,N_3596,N_3403);
or U3675 (N_3675,N_3474,N_3479);
xor U3676 (N_3676,N_3562,N_3449);
or U3677 (N_3677,N_3408,N_3534);
or U3678 (N_3678,N_3525,N_3574);
nand U3679 (N_3679,N_3537,N_3547);
or U3680 (N_3680,N_3503,N_3551);
and U3681 (N_3681,N_3575,N_3592);
xor U3682 (N_3682,N_3459,N_3467);
xor U3683 (N_3683,N_3402,N_3554);
nor U3684 (N_3684,N_3555,N_3435);
nor U3685 (N_3685,N_3580,N_3422);
or U3686 (N_3686,N_3570,N_3564);
nor U3687 (N_3687,N_3428,N_3427);
and U3688 (N_3688,N_3411,N_3539);
xnor U3689 (N_3689,N_3512,N_3546);
or U3690 (N_3690,N_3548,N_3437);
and U3691 (N_3691,N_3420,N_3595);
xor U3692 (N_3692,N_3552,N_3528);
and U3693 (N_3693,N_3581,N_3476);
or U3694 (N_3694,N_3561,N_3450);
or U3695 (N_3695,N_3464,N_3431);
nor U3696 (N_3696,N_3504,N_3473);
nand U3697 (N_3697,N_3487,N_3465);
nand U3698 (N_3698,N_3481,N_3584);
or U3699 (N_3699,N_3521,N_3455);
nor U3700 (N_3700,N_3487,N_3548);
and U3701 (N_3701,N_3546,N_3465);
or U3702 (N_3702,N_3512,N_3526);
and U3703 (N_3703,N_3543,N_3495);
or U3704 (N_3704,N_3472,N_3414);
xnor U3705 (N_3705,N_3587,N_3410);
and U3706 (N_3706,N_3591,N_3475);
nand U3707 (N_3707,N_3418,N_3455);
nor U3708 (N_3708,N_3532,N_3491);
and U3709 (N_3709,N_3497,N_3570);
and U3710 (N_3710,N_3532,N_3493);
xnor U3711 (N_3711,N_3444,N_3585);
nand U3712 (N_3712,N_3442,N_3416);
nor U3713 (N_3713,N_3530,N_3549);
nand U3714 (N_3714,N_3570,N_3544);
or U3715 (N_3715,N_3455,N_3453);
nor U3716 (N_3716,N_3488,N_3573);
or U3717 (N_3717,N_3431,N_3581);
and U3718 (N_3718,N_3579,N_3466);
and U3719 (N_3719,N_3420,N_3471);
nand U3720 (N_3720,N_3578,N_3433);
or U3721 (N_3721,N_3514,N_3435);
nor U3722 (N_3722,N_3407,N_3476);
and U3723 (N_3723,N_3433,N_3526);
nand U3724 (N_3724,N_3439,N_3433);
nand U3725 (N_3725,N_3486,N_3420);
or U3726 (N_3726,N_3574,N_3483);
nand U3727 (N_3727,N_3552,N_3494);
xor U3728 (N_3728,N_3536,N_3564);
or U3729 (N_3729,N_3425,N_3434);
nor U3730 (N_3730,N_3570,N_3598);
and U3731 (N_3731,N_3541,N_3523);
or U3732 (N_3732,N_3421,N_3583);
and U3733 (N_3733,N_3424,N_3467);
xor U3734 (N_3734,N_3598,N_3476);
nand U3735 (N_3735,N_3552,N_3402);
nor U3736 (N_3736,N_3535,N_3598);
and U3737 (N_3737,N_3461,N_3462);
nand U3738 (N_3738,N_3524,N_3513);
and U3739 (N_3739,N_3546,N_3439);
xnor U3740 (N_3740,N_3416,N_3462);
or U3741 (N_3741,N_3513,N_3428);
and U3742 (N_3742,N_3485,N_3572);
and U3743 (N_3743,N_3488,N_3485);
or U3744 (N_3744,N_3555,N_3429);
or U3745 (N_3745,N_3415,N_3506);
nand U3746 (N_3746,N_3564,N_3466);
or U3747 (N_3747,N_3531,N_3448);
and U3748 (N_3748,N_3586,N_3585);
and U3749 (N_3749,N_3489,N_3496);
and U3750 (N_3750,N_3436,N_3581);
xnor U3751 (N_3751,N_3530,N_3492);
or U3752 (N_3752,N_3466,N_3518);
nor U3753 (N_3753,N_3500,N_3440);
nor U3754 (N_3754,N_3531,N_3431);
nor U3755 (N_3755,N_3576,N_3450);
xor U3756 (N_3756,N_3491,N_3471);
nand U3757 (N_3757,N_3552,N_3599);
nand U3758 (N_3758,N_3430,N_3566);
or U3759 (N_3759,N_3525,N_3415);
and U3760 (N_3760,N_3567,N_3516);
or U3761 (N_3761,N_3402,N_3427);
nor U3762 (N_3762,N_3445,N_3409);
and U3763 (N_3763,N_3402,N_3418);
or U3764 (N_3764,N_3594,N_3532);
xor U3765 (N_3765,N_3423,N_3556);
nor U3766 (N_3766,N_3534,N_3487);
nand U3767 (N_3767,N_3417,N_3465);
and U3768 (N_3768,N_3463,N_3534);
nand U3769 (N_3769,N_3412,N_3551);
or U3770 (N_3770,N_3540,N_3565);
nor U3771 (N_3771,N_3534,N_3581);
and U3772 (N_3772,N_3597,N_3421);
nand U3773 (N_3773,N_3561,N_3491);
nor U3774 (N_3774,N_3559,N_3572);
or U3775 (N_3775,N_3473,N_3496);
or U3776 (N_3776,N_3449,N_3443);
xor U3777 (N_3777,N_3429,N_3467);
or U3778 (N_3778,N_3533,N_3491);
and U3779 (N_3779,N_3498,N_3452);
nand U3780 (N_3780,N_3511,N_3512);
or U3781 (N_3781,N_3517,N_3493);
nand U3782 (N_3782,N_3422,N_3421);
and U3783 (N_3783,N_3583,N_3441);
nand U3784 (N_3784,N_3569,N_3510);
or U3785 (N_3785,N_3544,N_3504);
and U3786 (N_3786,N_3440,N_3505);
nand U3787 (N_3787,N_3438,N_3461);
or U3788 (N_3788,N_3558,N_3426);
nor U3789 (N_3789,N_3590,N_3495);
xnor U3790 (N_3790,N_3538,N_3577);
or U3791 (N_3791,N_3577,N_3409);
nor U3792 (N_3792,N_3574,N_3598);
nand U3793 (N_3793,N_3400,N_3453);
and U3794 (N_3794,N_3491,N_3451);
xnor U3795 (N_3795,N_3592,N_3474);
nor U3796 (N_3796,N_3424,N_3577);
and U3797 (N_3797,N_3432,N_3409);
nor U3798 (N_3798,N_3420,N_3513);
or U3799 (N_3799,N_3501,N_3596);
or U3800 (N_3800,N_3645,N_3790);
or U3801 (N_3801,N_3780,N_3743);
nand U3802 (N_3802,N_3707,N_3687);
or U3803 (N_3803,N_3644,N_3690);
xnor U3804 (N_3804,N_3651,N_3708);
nor U3805 (N_3805,N_3726,N_3677);
and U3806 (N_3806,N_3758,N_3731);
and U3807 (N_3807,N_3764,N_3717);
xor U3808 (N_3808,N_3608,N_3772);
xor U3809 (N_3809,N_3722,N_3665);
and U3810 (N_3810,N_3799,N_3694);
nand U3811 (N_3811,N_3692,N_3693);
nor U3812 (N_3812,N_3703,N_3617);
or U3813 (N_3813,N_3754,N_3634);
and U3814 (N_3814,N_3785,N_3727);
nand U3815 (N_3815,N_3770,N_3689);
or U3816 (N_3816,N_3710,N_3668);
nand U3817 (N_3817,N_3671,N_3709);
and U3818 (N_3818,N_3674,N_3776);
or U3819 (N_3819,N_3784,N_3788);
xor U3820 (N_3820,N_3612,N_3673);
xor U3821 (N_3821,N_3620,N_3734);
nor U3822 (N_3822,N_3649,N_3691);
and U3823 (N_3823,N_3713,N_3669);
or U3824 (N_3824,N_3626,N_3633);
xor U3825 (N_3825,N_3605,N_3656);
nand U3826 (N_3826,N_3721,N_3604);
nor U3827 (N_3827,N_3616,N_3643);
or U3828 (N_3828,N_3623,N_3789);
or U3829 (N_3829,N_3787,N_3768);
nand U3830 (N_3830,N_3744,N_3704);
nand U3831 (N_3831,N_3683,N_3684);
or U3832 (N_3832,N_3697,N_3615);
nand U3833 (N_3833,N_3682,N_3662);
or U3834 (N_3834,N_3747,N_3783);
and U3835 (N_3835,N_3796,N_3700);
xnor U3836 (N_3836,N_3628,N_3648);
and U3837 (N_3837,N_3609,N_3688);
xor U3838 (N_3838,N_3716,N_3658);
or U3839 (N_3839,N_3752,N_3733);
and U3840 (N_3840,N_3771,N_3793);
or U3841 (N_3841,N_3705,N_3757);
xor U3842 (N_3842,N_3745,N_3659);
or U3843 (N_3843,N_3753,N_3714);
nor U3844 (N_3844,N_3718,N_3611);
xnor U3845 (N_3845,N_3676,N_3715);
xor U3846 (N_3846,N_3756,N_3701);
nor U3847 (N_3847,N_3781,N_3746);
nand U3848 (N_3848,N_3640,N_3739);
xor U3849 (N_3849,N_3627,N_3748);
nand U3850 (N_3850,N_3765,N_3653);
and U3851 (N_3851,N_3660,N_3678);
nor U3852 (N_3852,N_3680,N_3650);
nand U3853 (N_3853,N_3794,N_3610);
xnor U3854 (N_3854,N_3760,N_3742);
nand U3855 (N_3855,N_3724,N_3670);
nor U3856 (N_3856,N_3630,N_3729);
or U3857 (N_3857,N_3773,N_3798);
or U3858 (N_3858,N_3774,N_3619);
nand U3859 (N_3859,N_3636,N_3767);
nor U3860 (N_3860,N_3663,N_3681);
or U3861 (N_3861,N_3763,N_3606);
or U3862 (N_3862,N_3738,N_3601);
nor U3863 (N_3863,N_3711,N_3762);
or U3864 (N_3864,N_3654,N_3624);
nand U3865 (N_3865,N_3631,N_3792);
xnor U3866 (N_3866,N_3741,N_3679);
xnor U3867 (N_3867,N_3666,N_3755);
nand U3868 (N_3868,N_3706,N_3702);
xnor U3869 (N_3869,N_3750,N_3795);
xor U3870 (N_3870,N_3646,N_3779);
xnor U3871 (N_3871,N_3775,N_3751);
nand U3872 (N_3872,N_3642,N_3652);
or U3873 (N_3873,N_3695,N_3667);
nand U3874 (N_3874,N_3712,N_3735);
nor U3875 (N_3875,N_3686,N_3699);
nor U3876 (N_3876,N_3737,N_3618);
nor U3877 (N_3877,N_3736,N_3664);
and U3878 (N_3878,N_3769,N_3791);
nand U3879 (N_3879,N_3625,N_3641);
and U3880 (N_3880,N_3614,N_3786);
nor U3881 (N_3881,N_3761,N_3725);
nand U3882 (N_3882,N_3766,N_3672);
xor U3883 (N_3883,N_3797,N_3639);
nor U3884 (N_3884,N_3603,N_3638);
xor U3885 (N_3885,N_3600,N_3635);
nand U3886 (N_3886,N_3622,N_3777);
nand U3887 (N_3887,N_3602,N_3728);
and U3888 (N_3888,N_3749,N_3607);
or U3889 (N_3889,N_3723,N_3698);
or U3890 (N_3890,N_3720,N_3661);
and U3891 (N_3891,N_3675,N_3782);
or U3892 (N_3892,N_3613,N_3696);
nand U3893 (N_3893,N_3719,N_3629);
nand U3894 (N_3894,N_3632,N_3730);
and U3895 (N_3895,N_3685,N_3732);
nand U3896 (N_3896,N_3655,N_3647);
nor U3897 (N_3897,N_3778,N_3657);
nand U3898 (N_3898,N_3759,N_3637);
or U3899 (N_3899,N_3621,N_3740);
nand U3900 (N_3900,N_3787,N_3670);
nand U3901 (N_3901,N_3639,N_3662);
or U3902 (N_3902,N_3676,N_3700);
or U3903 (N_3903,N_3679,N_3655);
and U3904 (N_3904,N_3679,N_3777);
nand U3905 (N_3905,N_3711,N_3749);
xor U3906 (N_3906,N_3797,N_3633);
xor U3907 (N_3907,N_3603,N_3797);
or U3908 (N_3908,N_3632,N_3789);
nor U3909 (N_3909,N_3688,N_3763);
and U3910 (N_3910,N_3724,N_3687);
nor U3911 (N_3911,N_3707,N_3616);
and U3912 (N_3912,N_3616,N_3703);
or U3913 (N_3913,N_3662,N_3607);
nand U3914 (N_3914,N_3658,N_3666);
xnor U3915 (N_3915,N_3793,N_3634);
or U3916 (N_3916,N_3760,N_3694);
or U3917 (N_3917,N_3656,N_3718);
nand U3918 (N_3918,N_3729,N_3615);
nor U3919 (N_3919,N_3688,N_3787);
and U3920 (N_3920,N_3771,N_3784);
and U3921 (N_3921,N_3617,N_3600);
and U3922 (N_3922,N_3629,N_3680);
nand U3923 (N_3923,N_3684,N_3795);
xor U3924 (N_3924,N_3614,N_3606);
or U3925 (N_3925,N_3716,N_3761);
or U3926 (N_3926,N_3649,N_3781);
nand U3927 (N_3927,N_3656,N_3692);
xor U3928 (N_3928,N_3737,N_3752);
nand U3929 (N_3929,N_3732,N_3659);
or U3930 (N_3930,N_3646,N_3704);
nand U3931 (N_3931,N_3626,N_3751);
or U3932 (N_3932,N_3775,N_3637);
and U3933 (N_3933,N_3722,N_3753);
and U3934 (N_3934,N_3722,N_3737);
and U3935 (N_3935,N_3676,N_3789);
nand U3936 (N_3936,N_3693,N_3785);
nor U3937 (N_3937,N_3637,N_3666);
or U3938 (N_3938,N_3654,N_3731);
or U3939 (N_3939,N_3705,N_3797);
nor U3940 (N_3940,N_3777,N_3697);
nor U3941 (N_3941,N_3678,N_3651);
and U3942 (N_3942,N_3656,N_3690);
and U3943 (N_3943,N_3677,N_3722);
nand U3944 (N_3944,N_3685,N_3724);
or U3945 (N_3945,N_3747,N_3698);
nor U3946 (N_3946,N_3793,N_3764);
or U3947 (N_3947,N_3628,N_3791);
nor U3948 (N_3948,N_3730,N_3772);
xnor U3949 (N_3949,N_3718,N_3629);
or U3950 (N_3950,N_3752,N_3668);
and U3951 (N_3951,N_3616,N_3640);
nor U3952 (N_3952,N_3760,N_3657);
and U3953 (N_3953,N_3759,N_3784);
xor U3954 (N_3954,N_3772,N_3642);
nand U3955 (N_3955,N_3672,N_3600);
xor U3956 (N_3956,N_3777,N_3621);
and U3957 (N_3957,N_3774,N_3643);
xnor U3958 (N_3958,N_3615,N_3684);
and U3959 (N_3959,N_3773,N_3674);
xor U3960 (N_3960,N_3742,N_3629);
nor U3961 (N_3961,N_3648,N_3682);
nor U3962 (N_3962,N_3771,N_3641);
and U3963 (N_3963,N_3773,N_3714);
nand U3964 (N_3964,N_3714,N_3622);
xor U3965 (N_3965,N_3730,N_3725);
and U3966 (N_3966,N_3776,N_3635);
nor U3967 (N_3967,N_3678,N_3736);
and U3968 (N_3968,N_3695,N_3679);
or U3969 (N_3969,N_3648,N_3785);
nor U3970 (N_3970,N_3758,N_3669);
nor U3971 (N_3971,N_3724,N_3723);
nand U3972 (N_3972,N_3635,N_3604);
or U3973 (N_3973,N_3769,N_3735);
or U3974 (N_3974,N_3798,N_3735);
nand U3975 (N_3975,N_3778,N_3736);
and U3976 (N_3976,N_3762,N_3743);
or U3977 (N_3977,N_3648,N_3755);
or U3978 (N_3978,N_3722,N_3635);
or U3979 (N_3979,N_3642,N_3630);
nor U3980 (N_3980,N_3759,N_3748);
xor U3981 (N_3981,N_3616,N_3729);
or U3982 (N_3982,N_3630,N_3684);
xnor U3983 (N_3983,N_3761,N_3728);
or U3984 (N_3984,N_3637,N_3714);
or U3985 (N_3985,N_3798,N_3674);
nand U3986 (N_3986,N_3765,N_3728);
nor U3987 (N_3987,N_3761,N_3665);
xor U3988 (N_3988,N_3648,N_3707);
or U3989 (N_3989,N_3663,N_3729);
xor U3990 (N_3990,N_3680,N_3691);
nor U3991 (N_3991,N_3668,N_3796);
nand U3992 (N_3992,N_3666,N_3799);
nor U3993 (N_3993,N_3612,N_3708);
nand U3994 (N_3994,N_3729,N_3769);
and U3995 (N_3995,N_3712,N_3626);
xnor U3996 (N_3996,N_3625,N_3796);
and U3997 (N_3997,N_3731,N_3679);
and U3998 (N_3998,N_3600,N_3756);
nor U3999 (N_3999,N_3612,N_3733);
xnor U4000 (N_4000,N_3959,N_3826);
and U4001 (N_4001,N_3939,N_3865);
nor U4002 (N_4002,N_3849,N_3946);
nand U4003 (N_4003,N_3975,N_3862);
xnor U4004 (N_4004,N_3875,N_3982);
or U4005 (N_4005,N_3868,N_3893);
nor U4006 (N_4006,N_3836,N_3910);
xnor U4007 (N_4007,N_3935,N_3859);
nor U4008 (N_4008,N_3858,N_3867);
or U4009 (N_4009,N_3976,N_3874);
and U4010 (N_4010,N_3914,N_3825);
or U4011 (N_4011,N_3827,N_3885);
nor U4012 (N_4012,N_3809,N_3969);
and U4013 (N_4013,N_3949,N_3991);
and U4014 (N_4014,N_3916,N_3842);
xor U4015 (N_4015,N_3936,N_3958);
nor U4016 (N_4016,N_3844,N_3947);
nor U4017 (N_4017,N_3845,N_3841);
xnor U4018 (N_4018,N_3920,N_3964);
xor U4019 (N_4019,N_3888,N_3981);
nand U4020 (N_4020,N_3919,N_3989);
or U4021 (N_4021,N_3987,N_3806);
xnor U4022 (N_4022,N_3924,N_3945);
nor U4023 (N_4023,N_3922,N_3904);
and U4024 (N_4024,N_3896,N_3837);
or U4025 (N_4025,N_3899,N_3866);
and U4026 (N_4026,N_3817,N_3968);
and U4027 (N_4027,N_3878,N_3953);
and U4028 (N_4028,N_3978,N_3800);
nand U4029 (N_4029,N_3801,N_3930);
xor U4030 (N_4030,N_3889,N_3909);
nor U4031 (N_4031,N_3852,N_3960);
or U4032 (N_4032,N_3913,N_3938);
or U4033 (N_4033,N_3966,N_3818);
xor U4034 (N_4034,N_3944,N_3985);
xor U4035 (N_4035,N_3876,N_3814);
nor U4036 (N_4036,N_3973,N_3847);
xnor U4037 (N_4037,N_3870,N_3871);
xnor U4038 (N_4038,N_3918,N_3912);
xnor U4039 (N_4039,N_3905,N_3895);
xnor U4040 (N_4040,N_3872,N_3940);
xor U4041 (N_4041,N_3816,N_3835);
nand U4042 (N_4042,N_3917,N_3911);
xnor U4043 (N_4043,N_3880,N_3831);
nor U4044 (N_4044,N_3863,N_3950);
nor U4045 (N_4045,N_3903,N_3840);
nor U4046 (N_4046,N_3990,N_3963);
and U4047 (N_4047,N_3829,N_3902);
nand U4048 (N_4048,N_3873,N_3853);
and U4049 (N_4049,N_3979,N_3972);
or U4050 (N_4050,N_3883,N_3951);
nand U4051 (N_4051,N_3851,N_3995);
nand U4052 (N_4052,N_3857,N_3846);
nand U4053 (N_4053,N_3815,N_3833);
and U4054 (N_4054,N_3998,N_3996);
nand U4055 (N_4055,N_3900,N_3906);
or U4056 (N_4056,N_3928,N_3999);
and U4057 (N_4057,N_3984,N_3802);
nand U4058 (N_4058,N_3881,N_3823);
and U4059 (N_4059,N_3892,N_3993);
nand U4060 (N_4060,N_3957,N_3901);
and U4061 (N_4061,N_3861,N_3933);
or U4062 (N_4062,N_3811,N_3855);
and U4063 (N_4063,N_3908,N_3890);
nor U4064 (N_4064,N_3838,N_3821);
nand U4065 (N_4065,N_3891,N_3992);
and U4066 (N_4066,N_3843,N_3971);
nor U4067 (N_4067,N_3923,N_3931);
nor U4068 (N_4068,N_3921,N_3967);
or U4069 (N_4069,N_3932,N_3970);
xnor U4070 (N_4070,N_3804,N_3864);
nand U4071 (N_4071,N_3884,N_3927);
or U4072 (N_4072,N_3819,N_3805);
xnor U4073 (N_4073,N_3988,N_3925);
xnor U4074 (N_4074,N_3848,N_3980);
or U4075 (N_4075,N_3850,N_3929);
or U4076 (N_4076,N_3937,N_3915);
nand U4077 (N_4077,N_3856,N_3997);
and U4078 (N_4078,N_3854,N_3820);
and U4079 (N_4079,N_3882,N_3948);
xor U4080 (N_4080,N_3822,N_3860);
nand U4081 (N_4081,N_3886,N_3828);
xor U4082 (N_4082,N_3994,N_3824);
nand U4083 (N_4083,N_3952,N_3808);
xor U4084 (N_4084,N_3956,N_3961);
xnor U4085 (N_4085,N_3955,N_3834);
nand U4086 (N_4086,N_3965,N_3897);
nand U4087 (N_4087,N_3877,N_3986);
or U4088 (N_4088,N_3830,N_3954);
and U4089 (N_4089,N_3813,N_3803);
and U4090 (N_4090,N_3894,N_3977);
xor U4091 (N_4091,N_3934,N_3941);
nand U4092 (N_4092,N_3839,N_3943);
and U4093 (N_4093,N_3962,N_3807);
and U4094 (N_4094,N_3983,N_3812);
and U4095 (N_4095,N_3974,N_3887);
xor U4096 (N_4096,N_3879,N_3926);
nand U4097 (N_4097,N_3942,N_3810);
or U4098 (N_4098,N_3832,N_3907);
nand U4099 (N_4099,N_3898,N_3869);
xnor U4100 (N_4100,N_3863,N_3852);
nand U4101 (N_4101,N_3887,N_3941);
or U4102 (N_4102,N_3829,N_3862);
and U4103 (N_4103,N_3806,N_3930);
nand U4104 (N_4104,N_3818,N_3926);
or U4105 (N_4105,N_3994,N_3807);
or U4106 (N_4106,N_3993,N_3974);
and U4107 (N_4107,N_3959,N_3900);
or U4108 (N_4108,N_3995,N_3963);
or U4109 (N_4109,N_3962,N_3950);
xnor U4110 (N_4110,N_3946,N_3981);
nand U4111 (N_4111,N_3805,N_3966);
nor U4112 (N_4112,N_3905,N_3854);
nor U4113 (N_4113,N_3800,N_3878);
nor U4114 (N_4114,N_3901,N_3893);
or U4115 (N_4115,N_3917,N_3884);
and U4116 (N_4116,N_3932,N_3917);
or U4117 (N_4117,N_3815,N_3943);
and U4118 (N_4118,N_3916,N_3908);
nor U4119 (N_4119,N_3922,N_3985);
nand U4120 (N_4120,N_3816,N_3973);
xor U4121 (N_4121,N_3917,N_3933);
nand U4122 (N_4122,N_3832,N_3978);
or U4123 (N_4123,N_3846,N_3964);
or U4124 (N_4124,N_3836,N_3824);
nand U4125 (N_4125,N_3992,N_3938);
xor U4126 (N_4126,N_3834,N_3949);
and U4127 (N_4127,N_3878,N_3810);
nand U4128 (N_4128,N_3999,N_3909);
nand U4129 (N_4129,N_3924,N_3905);
xor U4130 (N_4130,N_3898,N_3865);
nor U4131 (N_4131,N_3876,N_3898);
nand U4132 (N_4132,N_3842,N_3861);
or U4133 (N_4133,N_3986,N_3940);
or U4134 (N_4134,N_3882,N_3851);
and U4135 (N_4135,N_3996,N_3917);
nor U4136 (N_4136,N_3946,N_3826);
or U4137 (N_4137,N_3981,N_3860);
nor U4138 (N_4138,N_3906,N_3931);
xor U4139 (N_4139,N_3838,N_3848);
or U4140 (N_4140,N_3986,N_3807);
nand U4141 (N_4141,N_3906,N_3814);
or U4142 (N_4142,N_3926,N_3921);
xor U4143 (N_4143,N_3936,N_3904);
xnor U4144 (N_4144,N_3866,N_3812);
and U4145 (N_4145,N_3856,N_3916);
and U4146 (N_4146,N_3873,N_3982);
or U4147 (N_4147,N_3942,N_3987);
or U4148 (N_4148,N_3929,N_3841);
xnor U4149 (N_4149,N_3906,N_3895);
nor U4150 (N_4150,N_3833,N_3888);
nor U4151 (N_4151,N_3818,N_3804);
nor U4152 (N_4152,N_3838,N_3983);
and U4153 (N_4153,N_3914,N_3963);
nor U4154 (N_4154,N_3942,N_3821);
or U4155 (N_4155,N_3917,N_3967);
or U4156 (N_4156,N_3816,N_3981);
nor U4157 (N_4157,N_3913,N_3882);
nand U4158 (N_4158,N_3900,N_3961);
nand U4159 (N_4159,N_3957,N_3885);
nand U4160 (N_4160,N_3909,N_3854);
nand U4161 (N_4161,N_3864,N_3938);
or U4162 (N_4162,N_3986,N_3867);
and U4163 (N_4163,N_3999,N_3871);
or U4164 (N_4164,N_3850,N_3804);
nand U4165 (N_4165,N_3924,N_3853);
nand U4166 (N_4166,N_3987,N_3955);
xnor U4167 (N_4167,N_3974,N_3812);
and U4168 (N_4168,N_3955,N_3804);
nor U4169 (N_4169,N_3920,N_3840);
or U4170 (N_4170,N_3913,N_3905);
nor U4171 (N_4171,N_3971,N_3952);
and U4172 (N_4172,N_3820,N_3830);
nor U4173 (N_4173,N_3902,N_3936);
nor U4174 (N_4174,N_3912,N_3915);
nand U4175 (N_4175,N_3896,N_3941);
or U4176 (N_4176,N_3954,N_3862);
nand U4177 (N_4177,N_3906,N_3994);
xnor U4178 (N_4178,N_3833,N_3874);
nand U4179 (N_4179,N_3904,N_3848);
nand U4180 (N_4180,N_3821,N_3925);
nor U4181 (N_4181,N_3894,N_3827);
and U4182 (N_4182,N_3830,N_3872);
and U4183 (N_4183,N_3888,N_3870);
nor U4184 (N_4184,N_3936,N_3817);
nor U4185 (N_4185,N_3986,N_3908);
nor U4186 (N_4186,N_3906,N_3833);
or U4187 (N_4187,N_3849,N_3976);
or U4188 (N_4188,N_3877,N_3867);
xnor U4189 (N_4189,N_3864,N_3935);
nor U4190 (N_4190,N_3939,N_3886);
and U4191 (N_4191,N_3889,N_3848);
nand U4192 (N_4192,N_3836,N_3850);
xnor U4193 (N_4193,N_3925,N_3847);
xor U4194 (N_4194,N_3883,N_3808);
nand U4195 (N_4195,N_3944,N_3984);
nand U4196 (N_4196,N_3868,N_3978);
nor U4197 (N_4197,N_3855,N_3872);
and U4198 (N_4198,N_3886,N_3936);
or U4199 (N_4199,N_3933,N_3863);
nand U4200 (N_4200,N_4050,N_4067);
xnor U4201 (N_4201,N_4003,N_4103);
nor U4202 (N_4202,N_4146,N_4007);
xnor U4203 (N_4203,N_4099,N_4184);
nor U4204 (N_4204,N_4095,N_4046);
or U4205 (N_4205,N_4018,N_4144);
nor U4206 (N_4206,N_4166,N_4051);
or U4207 (N_4207,N_4000,N_4105);
nand U4208 (N_4208,N_4118,N_4048);
and U4209 (N_4209,N_4170,N_4187);
nor U4210 (N_4210,N_4196,N_4083);
and U4211 (N_4211,N_4194,N_4155);
or U4212 (N_4212,N_4060,N_4017);
nor U4213 (N_4213,N_4130,N_4025);
nand U4214 (N_4214,N_4181,N_4192);
or U4215 (N_4215,N_4016,N_4064);
or U4216 (N_4216,N_4027,N_4176);
or U4217 (N_4217,N_4162,N_4157);
nand U4218 (N_4218,N_4085,N_4120);
and U4219 (N_4219,N_4053,N_4113);
nand U4220 (N_4220,N_4056,N_4005);
and U4221 (N_4221,N_4164,N_4001);
nor U4222 (N_4222,N_4022,N_4014);
xnor U4223 (N_4223,N_4008,N_4147);
and U4224 (N_4224,N_4137,N_4075);
xor U4225 (N_4225,N_4133,N_4126);
or U4226 (N_4226,N_4026,N_4088);
xnor U4227 (N_4227,N_4115,N_4140);
xnor U4228 (N_4228,N_4078,N_4084);
and U4229 (N_4229,N_4044,N_4074);
and U4230 (N_4230,N_4108,N_4172);
or U4231 (N_4231,N_4106,N_4180);
and U4232 (N_4232,N_4093,N_4132);
nor U4233 (N_4233,N_4071,N_4136);
xnor U4234 (N_4234,N_4058,N_4021);
nand U4235 (N_4235,N_4042,N_4189);
xnor U4236 (N_4236,N_4109,N_4114);
and U4237 (N_4237,N_4143,N_4195);
nand U4238 (N_4238,N_4047,N_4043);
nor U4239 (N_4239,N_4160,N_4077);
and U4240 (N_4240,N_4198,N_4121);
xor U4241 (N_4241,N_4066,N_4020);
or U4242 (N_4242,N_4086,N_4135);
nand U4243 (N_4243,N_4029,N_4102);
nor U4244 (N_4244,N_4131,N_4117);
nand U4245 (N_4245,N_4129,N_4100);
and U4246 (N_4246,N_4023,N_4110);
nor U4247 (N_4247,N_4152,N_4142);
nand U4248 (N_4248,N_4069,N_4006);
xnor U4249 (N_4249,N_4057,N_4054);
xnor U4250 (N_4250,N_4171,N_4038);
nor U4251 (N_4251,N_4062,N_4168);
nand U4252 (N_4252,N_4197,N_4070);
nand U4253 (N_4253,N_4032,N_4141);
and U4254 (N_4254,N_4049,N_4175);
and U4255 (N_4255,N_4154,N_4098);
xor U4256 (N_4256,N_4024,N_4036);
and U4257 (N_4257,N_4188,N_4012);
or U4258 (N_4258,N_4041,N_4178);
xnor U4259 (N_4259,N_4191,N_4091);
and U4260 (N_4260,N_4149,N_4161);
and U4261 (N_4261,N_4080,N_4055);
and U4262 (N_4262,N_4011,N_4040);
xnor U4263 (N_4263,N_4186,N_4035);
xor U4264 (N_4264,N_4097,N_4165);
nand U4265 (N_4265,N_4123,N_4163);
nor U4266 (N_4266,N_4033,N_4090);
xnor U4267 (N_4267,N_4124,N_4079);
xor U4268 (N_4268,N_4094,N_4092);
nor U4269 (N_4269,N_4153,N_4045);
nor U4270 (N_4270,N_4019,N_4112);
and U4271 (N_4271,N_4111,N_4156);
or U4272 (N_4272,N_4125,N_4116);
and U4273 (N_4273,N_4076,N_4148);
nand U4274 (N_4274,N_4150,N_4139);
nand U4275 (N_4275,N_4096,N_4002);
xor U4276 (N_4276,N_4081,N_4031);
xor U4277 (N_4277,N_4199,N_4030);
and U4278 (N_4278,N_4028,N_4119);
nor U4279 (N_4279,N_4107,N_4159);
nor U4280 (N_4280,N_4061,N_4182);
xor U4281 (N_4281,N_4169,N_4009);
xnor U4282 (N_4282,N_4004,N_4138);
or U4283 (N_4283,N_4127,N_4151);
xor U4284 (N_4284,N_4059,N_4010);
or U4285 (N_4285,N_4183,N_4052);
nand U4286 (N_4286,N_4082,N_4037);
nand U4287 (N_4287,N_4134,N_4174);
or U4288 (N_4288,N_4177,N_4063);
or U4289 (N_4289,N_4089,N_4068);
xnor U4290 (N_4290,N_4122,N_4128);
xnor U4291 (N_4291,N_4013,N_4073);
nor U4292 (N_4292,N_4101,N_4034);
nand U4293 (N_4293,N_4104,N_4039);
or U4294 (N_4294,N_4072,N_4185);
xnor U4295 (N_4295,N_4158,N_4179);
and U4296 (N_4296,N_4087,N_4145);
xor U4297 (N_4297,N_4065,N_4193);
and U4298 (N_4298,N_4167,N_4015);
xor U4299 (N_4299,N_4173,N_4190);
and U4300 (N_4300,N_4165,N_4077);
and U4301 (N_4301,N_4148,N_4177);
or U4302 (N_4302,N_4096,N_4108);
and U4303 (N_4303,N_4026,N_4092);
nor U4304 (N_4304,N_4041,N_4004);
xnor U4305 (N_4305,N_4094,N_4080);
xor U4306 (N_4306,N_4173,N_4140);
or U4307 (N_4307,N_4012,N_4068);
xor U4308 (N_4308,N_4145,N_4012);
nor U4309 (N_4309,N_4029,N_4195);
nor U4310 (N_4310,N_4047,N_4108);
nor U4311 (N_4311,N_4092,N_4098);
nand U4312 (N_4312,N_4142,N_4192);
nand U4313 (N_4313,N_4197,N_4104);
and U4314 (N_4314,N_4005,N_4073);
and U4315 (N_4315,N_4038,N_4044);
nand U4316 (N_4316,N_4089,N_4069);
nor U4317 (N_4317,N_4011,N_4147);
and U4318 (N_4318,N_4155,N_4183);
nand U4319 (N_4319,N_4094,N_4154);
and U4320 (N_4320,N_4053,N_4111);
xor U4321 (N_4321,N_4166,N_4157);
xnor U4322 (N_4322,N_4115,N_4098);
nand U4323 (N_4323,N_4141,N_4026);
or U4324 (N_4324,N_4134,N_4021);
xnor U4325 (N_4325,N_4147,N_4009);
or U4326 (N_4326,N_4150,N_4186);
and U4327 (N_4327,N_4166,N_4104);
or U4328 (N_4328,N_4066,N_4187);
nor U4329 (N_4329,N_4068,N_4048);
nor U4330 (N_4330,N_4069,N_4054);
nand U4331 (N_4331,N_4125,N_4060);
and U4332 (N_4332,N_4087,N_4132);
xnor U4333 (N_4333,N_4095,N_4108);
xor U4334 (N_4334,N_4024,N_4011);
nor U4335 (N_4335,N_4051,N_4152);
and U4336 (N_4336,N_4109,N_4036);
or U4337 (N_4337,N_4005,N_4136);
nor U4338 (N_4338,N_4078,N_4027);
nor U4339 (N_4339,N_4156,N_4046);
or U4340 (N_4340,N_4074,N_4077);
or U4341 (N_4341,N_4101,N_4132);
xor U4342 (N_4342,N_4179,N_4008);
nor U4343 (N_4343,N_4167,N_4017);
and U4344 (N_4344,N_4127,N_4110);
and U4345 (N_4345,N_4085,N_4074);
nor U4346 (N_4346,N_4006,N_4126);
nand U4347 (N_4347,N_4131,N_4094);
xnor U4348 (N_4348,N_4076,N_4156);
xnor U4349 (N_4349,N_4079,N_4044);
and U4350 (N_4350,N_4147,N_4175);
nor U4351 (N_4351,N_4166,N_4184);
xor U4352 (N_4352,N_4036,N_4146);
nand U4353 (N_4353,N_4128,N_4139);
or U4354 (N_4354,N_4056,N_4167);
or U4355 (N_4355,N_4173,N_4063);
nor U4356 (N_4356,N_4098,N_4001);
nand U4357 (N_4357,N_4088,N_4183);
xor U4358 (N_4358,N_4089,N_4121);
nand U4359 (N_4359,N_4014,N_4088);
nor U4360 (N_4360,N_4103,N_4070);
or U4361 (N_4361,N_4129,N_4140);
xnor U4362 (N_4362,N_4141,N_4169);
nor U4363 (N_4363,N_4139,N_4176);
or U4364 (N_4364,N_4014,N_4015);
nor U4365 (N_4365,N_4117,N_4067);
and U4366 (N_4366,N_4111,N_4068);
or U4367 (N_4367,N_4185,N_4126);
xnor U4368 (N_4368,N_4130,N_4086);
xnor U4369 (N_4369,N_4067,N_4148);
nand U4370 (N_4370,N_4086,N_4171);
xnor U4371 (N_4371,N_4064,N_4134);
xnor U4372 (N_4372,N_4038,N_4130);
or U4373 (N_4373,N_4138,N_4141);
nand U4374 (N_4374,N_4179,N_4027);
and U4375 (N_4375,N_4094,N_4152);
nor U4376 (N_4376,N_4010,N_4006);
nand U4377 (N_4377,N_4176,N_4010);
or U4378 (N_4378,N_4084,N_4165);
xor U4379 (N_4379,N_4141,N_4181);
nand U4380 (N_4380,N_4126,N_4049);
or U4381 (N_4381,N_4082,N_4157);
and U4382 (N_4382,N_4075,N_4043);
or U4383 (N_4383,N_4045,N_4161);
nand U4384 (N_4384,N_4061,N_4175);
nor U4385 (N_4385,N_4024,N_4157);
and U4386 (N_4386,N_4134,N_4032);
xnor U4387 (N_4387,N_4145,N_4009);
and U4388 (N_4388,N_4133,N_4167);
or U4389 (N_4389,N_4002,N_4120);
nand U4390 (N_4390,N_4082,N_4137);
or U4391 (N_4391,N_4059,N_4068);
and U4392 (N_4392,N_4027,N_4165);
nand U4393 (N_4393,N_4102,N_4150);
xnor U4394 (N_4394,N_4165,N_4092);
nand U4395 (N_4395,N_4060,N_4112);
xor U4396 (N_4396,N_4135,N_4128);
nand U4397 (N_4397,N_4036,N_4187);
and U4398 (N_4398,N_4120,N_4040);
and U4399 (N_4399,N_4065,N_4136);
or U4400 (N_4400,N_4291,N_4337);
nor U4401 (N_4401,N_4287,N_4297);
nand U4402 (N_4402,N_4316,N_4217);
or U4403 (N_4403,N_4243,N_4300);
nand U4404 (N_4404,N_4391,N_4328);
and U4405 (N_4405,N_4336,N_4234);
or U4406 (N_4406,N_4314,N_4364);
nand U4407 (N_4407,N_4200,N_4263);
nand U4408 (N_4408,N_4371,N_4223);
nor U4409 (N_4409,N_4289,N_4239);
xnor U4410 (N_4410,N_4272,N_4228);
nor U4411 (N_4411,N_4224,N_4377);
xnor U4412 (N_4412,N_4214,N_4219);
nor U4413 (N_4413,N_4249,N_4344);
nor U4414 (N_4414,N_4346,N_4379);
xor U4415 (N_4415,N_4397,N_4309);
or U4416 (N_4416,N_4237,N_4203);
nand U4417 (N_4417,N_4395,N_4313);
or U4418 (N_4418,N_4247,N_4354);
xor U4419 (N_4419,N_4385,N_4343);
xnor U4420 (N_4420,N_4215,N_4329);
or U4421 (N_4421,N_4232,N_4295);
nand U4422 (N_4422,N_4251,N_4208);
nor U4423 (N_4423,N_4380,N_4281);
xor U4424 (N_4424,N_4386,N_4330);
xnor U4425 (N_4425,N_4393,N_4372);
nand U4426 (N_4426,N_4279,N_4242);
nor U4427 (N_4427,N_4335,N_4348);
nand U4428 (N_4428,N_4369,N_4227);
nor U4429 (N_4429,N_4288,N_4278);
and U4430 (N_4430,N_4229,N_4390);
xnor U4431 (N_4431,N_4218,N_4248);
nand U4432 (N_4432,N_4274,N_4366);
nor U4433 (N_4433,N_4210,N_4349);
nor U4434 (N_4434,N_4262,N_4374);
xor U4435 (N_4435,N_4353,N_4205);
nor U4436 (N_4436,N_4277,N_4238);
nand U4437 (N_4437,N_4352,N_4333);
nor U4438 (N_4438,N_4387,N_4368);
and U4439 (N_4439,N_4271,N_4202);
xnor U4440 (N_4440,N_4311,N_4254);
nor U4441 (N_4441,N_4222,N_4399);
nand U4442 (N_4442,N_4221,N_4357);
nand U4443 (N_4443,N_4304,N_4206);
and U4444 (N_4444,N_4308,N_4201);
and U4445 (N_4445,N_4240,N_4338);
xnor U4446 (N_4446,N_4323,N_4381);
and U4447 (N_4447,N_4356,N_4266);
or U4448 (N_4448,N_4216,N_4332);
nor U4449 (N_4449,N_4231,N_4236);
xor U4450 (N_4450,N_4261,N_4382);
nand U4451 (N_4451,N_4303,N_4334);
xor U4452 (N_4452,N_4244,N_4375);
or U4453 (N_4453,N_4358,N_4230);
nand U4454 (N_4454,N_4253,N_4355);
and U4455 (N_4455,N_4282,N_4267);
and U4456 (N_4456,N_4307,N_4235);
nor U4457 (N_4457,N_4299,N_4373);
or U4458 (N_4458,N_4270,N_4315);
and U4459 (N_4459,N_4305,N_4389);
or U4460 (N_4460,N_4384,N_4365);
xor U4461 (N_4461,N_4339,N_4285);
nor U4462 (N_4462,N_4204,N_4290);
and U4463 (N_4463,N_4225,N_4213);
nor U4464 (N_4464,N_4269,N_4245);
xor U4465 (N_4465,N_4293,N_4211);
and U4466 (N_4466,N_4345,N_4298);
and U4467 (N_4467,N_4360,N_4376);
and U4468 (N_4468,N_4246,N_4325);
nor U4469 (N_4469,N_4370,N_4321);
xor U4470 (N_4470,N_4260,N_4317);
and U4471 (N_4471,N_4284,N_4283);
nand U4472 (N_4472,N_4265,N_4341);
nor U4473 (N_4473,N_4212,N_4398);
or U4474 (N_4474,N_4351,N_4396);
or U4475 (N_4475,N_4226,N_4252);
and U4476 (N_4476,N_4320,N_4273);
nor U4477 (N_4477,N_4347,N_4319);
nand U4478 (N_4478,N_4367,N_4312);
xnor U4479 (N_4479,N_4340,N_4342);
and U4480 (N_4480,N_4363,N_4388);
nand U4481 (N_4481,N_4378,N_4233);
or U4482 (N_4482,N_4292,N_4302);
nor U4483 (N_4483,N_4359,N_4361);
xor U4484 (N_4484,N_4220,N_4392);
xnor U4485 (N_4485,N_4296,N_4275);
or U4486 (N_4486,N_4327,N_4350);
xnor U4487 (N_4487,N_4383,N_4209);
nand U4488 (N_4488,N_4250,N_4259);
or U4489 (N_4489,N_4286,N_4241);
and U4490 (N_4490,N_4310,N_4331);
and U4491 (N_4491,N_4264,N_4207);
or U4492 (N_4492,N_4362,N_4294);
nor U4493 (N_4493,N_4318,N_4258);
and U4494 (N_4494,N_4394,N_4268);
nand U4495 (N_4495,N_4257,N_4256);
nor U4496 (N_4496,N_4322,N_4255);
xnor U4497 (N_4497,N_4326,N_4306);
nor U4498 (N_4498,N_4276,N_4301);
and U4499 (N_4499,N_4280,N_4324);
nand U4500 (N_4500,N_4353,N_4365);
and U4501 (N_4501,N_4222,N_4317);
xor U4502 (N_4502,N_4231,N_4249);
or U4503 (N_4503,N_4302,N_4270);
and U4504 (N_4504,N_4293,N_4268);
nor U4505 (N_4505,N_4208,N_4351);
or U4506 (N_4506,N_4383,N_4333);
xnor U4507 (N_4507,N_4317,N_4202);
nor U4508 (N_4508,N_4346,N_4261);
or U4509 (N_4509,N_4372,N_4235);
or U4510 (N_4510,N_4253,N_4281);
nor U4511 (N_4511,N_4229,N_4249);
and U4512 (N_4512,N_4323,N_4275);
or U4513 (N_4513,N_4386,N_4255);
and U4514 (N_4514,N_4338,N_4245);
nand U4515 (N_4515,N_4392,N_4273);
and U4516 (N_4516,N_4215,N_4277);
nand U4517 (N_4517,N_4223,N_4332);
nand U4518 (N_4518,N_4313,N_4399);
nor U4519 (N_4519,N_4343,N_4313);
or U4520 (N_4520,N_4226,N_4219);
nand U4521 (N_4521,N_4368,N_4393);
xnor U4522 (N_4522,N_4338,N_4312);
nor U4523 (N_4523,N_4288,N_4352);
and U4524 (N_4524,N_4236,N_4212);
nor U4525 (N_4525,N_4379,N_4365);
nand U4526 (N_4526,N_4249,N_4202);
nor U4527 (N_4527,N_4336,N_4310);
nand U4528 (N_4528,N_4303,N_4266);
or U4529 (N_4529,N_4255,N_4257);
nand U4530 (N_4530,N_4261,N_4227);
nand U4531 (N_4531,N_4339,N_4324);
and U4532 (N_4532,N_4381,N_4351);
and U4533 (N_4533,N_4346,N_4270);
nand U4534 (N_4534,N_4396,N_4239);
or U4535 (N_4535,N_4273,N_4359);
nor U4536 (N_4536,N_4264,N_4366);
nand U4537 (N_4537,N_4319,N_4369);
and U4538 (N_4538,N_4243,N_4324);
or U4539 (N_4539,N_4381,N_4313);
nor U4540 (N_4540,N_4370,N_4352);
and U4541 (N_4541,N_4205,N_4253);
nor U4542 (N_4542,N_4341,N_4317);
nor U4543 (N_4543,N_4372,N_4250);
or U4544 (N_4544,N_4356,N_4371);
nor U4545 (N_4545,N_4231,N_4388);
and U4546 (N_4546,N_4216,N_4306);
and U4547 (N_4547,N_4383,N_4202);
and U4548 (N_4548,N_4378,N_4322);
nor U4549 (N_4549,N_4237,N_4232);
and U4550 (N_4550,N_4202,N_4297);
nand U4551 (N_4551,N_4282,N_4315);
and U4552 (N_4552,N_4231,N_4361);
nor U4553 (N_4553,N_4360,N_4298);
or U4554 (N_4554,N_4312,N_4217);
nand U4555 (N_4555,N_4365,N_4345);
nand U4556 (N_4556,N_4272,N_4381);
nand U4557 (N_4557,N_4336,N_4221);
nor U4558 (N_4558,N_4304,N_4236);
xor U4559 (N_4559,N_4221,N_4301);
nand U4560 (N_4560,N_4288,N_4343);
nor U4561 (N_4561,N_4359,N_4204);
nand U4562 (N_4562,N_4319,N_4360);
xor U4563 (N_4563,N_4291,N_4383);
nor U4564 (N_4564,N_4350,N_4264);
nor U4565 (N_4565,N_4233,N_4380);
xor U4566 (N_4566,N_4344,N_4325);
and U4567 (N_4567,N_4247,N_4290);
or U4568 (N_4568,N_4249,N_4320);
or U4569 (N_4569,N_4313,N_4231);
nand U4570 (N_4570,N_4377,N_4235);
nand U4571 (N_4571,N_4276,N_4225);
and U4572 (N_4572,N_4351,N_4278);
and U4573 (N_4573,N_4315,N_4264);
nand U4574 (N_4574,N_4337,N_4206);
or U4575 (N_4575,N_4200,N_4295);
xor U4576 (N_4576,N_4245,N_4397);
xor U4577 (N_4577,N_4253,N_4217);
or U4578 (N_4578,N_4322,N_4276);
nor U4579 (N_4579,N_4329,N_4295);
nand U4580 (N_4580,N_4236,N_4384);
or U4581 (N_4581,N_4307,N_4370);
and U4582 (N_4582,N_4317,N_4313);
nor U4583 (N_4583,N_4244,N_4279);
nor U4584 (N_4584,N_4250,N_4239);
nor U4585 (N_4585,N_4266,N_4375);
xor U4586 (N_4586,N_4379,N_4313);
nor U4587 (N_4587,N_4288,N_4301);
or U4588 (N_4588,N_4361,N_4316);
or U4589 (N_4589,N_4385,N_4227);
xor U4590 (N_4590,N_4211,N_4346);
nor U4591 (N_4591,N_4354,N_4397);
xnor U4592 (N_4592,N_4374,N_4322);
xnor U4593 (N_4593,N_4290,N_4210);
nand U4594 (N_4594,N_4355,N_4225);
nor U4595 (N_4595,N_4232,N_4329);
and U4596 (N_4596,N_4342,N_4300);
nor U4597 (N_4597,N_4304,N_4287);
or U4598 (N_4598,N_4291,N_4202);
xnor U4599 (N_4599,N_4263,N_4306);
nor U4600 (N_4600,N_4513,N_4477);
xor U4601 (N_4601,N_4573,N_4548);
or U4602 (N_4602,N_4499,N_4462);
or U4603 (N_4603,N_4459,N_4569);
and U4604 (N_4604,N_4501,N_4516);
or U4605 (N_4605,N_4409,N_4416);
nor U4606 (N_4606,N_4478,N_4420);
xnor U4607 (N_4607,N_4401,N_4560);
or U4608 (N_4608,N_4468,N_4567);
xor U4609 (N_4609,N_4551,N_4521);
xor U4610 (N_4610,N_4557,N_4599);
nand U4611 (N_4611,N_4490,N_4568);
xor U4612 (N_4612,N_4564,N_4469);
and U4613 (N_4613,N_4533,N_4503);
or U4614 (N_4614,N_4480,N_4570);
and U4615 (N_4615,N_4576,N_4437);
nor U4616 (N_4616,N_4473,N_4577);
or U4617 (N_4617,N_4565,N_4435);
and U4618 (N_4618,N_4422,N_4479);
nor U4619 (N_4619,N_4431,N_4474);
or U4620 (N_4620,N_4508,N_4586);
xor U4621 (N_4621,N_4593,N_4543);
nor U4622 (N_4622,N_4582,N_4465);
nor U4623 (N_4623,N_4550,N_4590);
xnor U4624 (N_4624,N_4408,N_4509);
nand U4625 (N_4625,N_4578,N_4587);
and U4626 (N_4626,N_4585,N_4574);
or U4627 (N_4627,N_4400,N_4522);
nand U4628 (N_4628,N_4546,N_4524);
and U4629 (N_4629,N_4453,N_4559);
nor U4630 (N_4630,N_4502,N_4447);
nand U4631 (N_4631,N_4506,N_4498);
or U4632 (N_4632,N_4417,N_4563);
nand U4633 (N_4633,N_4427,N_4597);
xor U4634 (N_4634,N_4491,N_4575);
xnor U4635 (N_4635,N_4412,N_4445);
and U4636 (N_4636,N_4429,N_4457);
nand U4637 (N_4637,N_4596,N_4413);
nand U4638 (N_4638,N_4443,N_4542);
or U4639 (N_4639,N_4484,N_4558);
nor U4640 (N_4640,N_4512,N_4483);
nand U4641 (N_4641,N_4486,N_4460);
nor U4642 (N_4642,N_4539,N_4554);
nor U4643 (N_4643,N_4519,N_4549);
or U4644 (N_4644,N_4482,N_4538);
xnor U4645 (N_4645,N_4467,N_4588);
xnor U4646 (N_4646,N_4406,N_4481);
nor U4647 (N_4647,N_4507,N_4494);
or U4648 (N_4648,N_4493,N_4535);
or U4649 (N_4649,N_4584,N_4544);
and U4650 (N_4650,N_4485,N_4451);
nor U4651 (N_4651,N_4531,N_4419);
xnor U4652 (N_4652,N_4556,N_4444);
and U4653 (N_4653,N_4511,N_4438);
xor U4654 (N_4654,N_4526,N_4488);
and U4655 (N_4655,N_4471,N_4500);
nand U4656 (N_4656,N_4475,N_4530);
xor U4657 (N_4657,N_4594,N_4532);
nor U4658 (N_4658,N_4515,N_4464);
or U4659 (N_4659,N_4425,N_4547);
or U4660 (N_4660,N_4452,N_4402);
or U4661 (N_4661,N_4518,N_4421);
nand U4662 (N_4662,N_4598,N_4514);
nand U4663 (N_4663,N_4495,N_4589);
nor U4664 (N_4664,N_4528,N_4449);
or U4665 (N_4665,N_4463,N_4487);
xor U4666 (N_4666,N_4553,N_4442);
or U4667 (N_4667,N_4537,N_4403);
or U4668 (N_4668,N_4579,N_4572);
or U4669 (N_4669,N_4434,N_4418);
or U4670 (N_4670,N_4433,N_4562);
nor U4671 (N_4671,N_4439,N_4424);
and U4672 (N_4672,N_4470,N_4517);
or U4673 (N_4673,N_4555,N_4428);
nand U4674 (N_4674,N_4405,N_4566);
and U4675 (N_4675,N_4497,N_4440);
nand U4676 (N_4676,N_4407,N_4461);
xor U4677 (N_4677,N_4545,N_4536);
nor U4678 (N_4678,N_4436,N_4561);
nand U4679 (N_4679,N_4446,N_4472);
or U4680 (N_4680,N_4534,N_4414);
nand U4681 (N_4681,N_4496,N_4591);
xnor U4682 (N_4682,N_4592,N_4450);
or U4683 (N_4683,N_4595,N_4458);
nor U4684 (N_4684,N_4476,N_4525);
or U4685 (N_4685,N_4510,N_4489);
and U4686 (N_4686,N_4571,N_4454);
nand U4687 (N_4687,N_4456,N_4527);
or U4688 (N_4688,N_4455,N_4541);
and U4689 (N_4689,N_4529,N_4426);
or U4690 (N_4690,N_4504,N_4583);
or U4691 (N_4691,N_4441,N_4505);
xor U4692 (N_4692,N_4466,N_4430);
nor U4693 (N_4693,N_4404,N_4432);
nand U4694 (N_4694,N_4581,N_4448);
xnor U4695 (N_4695,N_4410,N_4415);
xnor U4696 (N_4696,N_4540,N_4580);
and U4697 (N_4697,N_4423,N_4520);
or U4698 (N_4698,N_4411,N_4552);
or U4699 (N_4699,N_4492,N_4523);
and U4700 (N_4700,N_4526,N_4546);
and U4701 (N_4701,N_4412,N_4568);
xnor U4702 (N_4702,N_4592,N_4464);
nand U4703 (N_4703,N_4409,N_4452);
nor U4704 (N_4704,N_4539,N_4472);
nor U4705 (N_4705,N_4495,N_4410);
xor U4706 (N_4706,N_4432,N_4576);
and U4707 (N_4707,N_4533,N_4424);
or U4708 (N_4708,N_4417,N_4426);
or U4709 (N_4709,N_4419,N_4448);
xor U4710 (N_4710,N_4579,N_4491);
and U4711 (N_4711,N_4567,N_4452);
and U4712 (N_4712,N_4485,N_4531);
nor U4713 (N_4713,N_4513,N_4527);
nor U4714 (N_4714,N_4589,N_4418);
nor U4715 (N_4715,N_4483,N_4559);
or U4716 (N_4716,N_4578,N_4536);
and U4717 (N_4717,N_4548,N_4524);
and U4718 (N_4718,N_4575,N_4414);
xor U4719 (N_4719,N_4520,N_4405);
or U4720 (N_4720,N_4548,N_4481);
xnor U4721 (N_4721,N_4428,N_4412);
and U4722 (N_4722,N_4486,N_4527);
or U4723 (N_4723,N_4490,N_4517);
and U4724 (N_4724,N_4529,N_4482);
and U4725 (N_4725,N_4402,N_4465);
xnor U4726 (N_4726,N_4503,N_4455);
nand U4727 (N_4727,N_4464,N_4581);
nor U4728 (N_4728,N_4430,N_4564);
nand U4729 (N_4729,N_4481,N_4515);
xor U4730 (N_4730,N_4565,N_4554);
nand U4731 (N_4731,N_4542,N_4499);
xor U4732 (N_4732,N_4419,N_4538);
or U4733 (N_4733,N_4581,N_4403);
nand U4734 (N_4734,N_4591,N_4556);
or U4735 (N_4735,N_4547,N_4460);
nor U4736 (N_4736,N_4597,N_4552);
nand U4737 (N_4737,N_4555,N_4500);
nor U4738 (N_4738,N_4442,N_4584);
xor U4739 (N_4739,N_4544,N_4439);
nand U4740 (N_4740,N_4452,N_4550);
or U4741 (N_4741,N_4406,N_4447);
or U4742 (N_4742,N_4550,N_4530);
or U4743 (N_4743,N_4441,N_4539);
xor U4744 (N_4744,N_4536,N_4559);
xor U4745 (N_4745,N_4425,N_4497);
nor U4746 (N_4746,N_4528,N_4491);
or U4747 (N_4747,N_4501,N_4454);
nand U4748 (N_4748,N_4424,N_4427);
xnor U4749 (N_4749,N_4587,N_4575);
or U4750 (N_4750,N_4464,N_4500);
nand U4751 (N_4751,N_4587,N_4551);
xnor U4752 (N_4752,N_4454,N_4473);
or U4753 (N_4753,N_4469,N_4565);
or U4754 (N_4754,N_4498,N_4477);
nor U4755 (N_4755,N_4562,N_4469);
and U4756 (N_4756,N_4497,N_4462);
and U4757 (N_4757,N_4571,N_4562);
xnor U4758 (N_4758,N_4584,N_4564);
xor U4759 (N_4759,N_4479,N_4467);
nand U4760 (N_4760,N_4489,N_4548);
xor U4761 (N_4761,N_4510,N_4475);
nand U4762 (N_4762,N_4454,N_4433);
nand U4763 (N_4763,N_4443,N_4562);
and U4764 (N_4764,N_4530,N_4537);
or U4765 (N_4765,N_4511,N_4567);
and U4766 (N_4766,N_4435,N_4456);
xor U4767 (N_4767,N_4570,N_4599);
or U4768 (N_4768,N_4471,N_4444);
or U4769 (N_4769,N_4517,N_4498);
and U4770 (N_4770,N_4598,N_4460);
nand U4771 (N_4771,N_4482,N_4431);
xor U4772 (N_4772,N_4446,N_4429);
and U4773 (N_4773,N_4463,N_4533);
or U4774 (N_4774,N_4411,N_4473);
and U4775 (N_4775,N_4476,N_4498);
or U4776 (N_4776,N_4414,N_4525);
nor U4777 (N_4777,N_4454,N_4465);
nor U4778 (N_4778,N_4483,N_4445);
xor U4779 (N_4779,N_4508,N_4513);
or U4780 (N_4780,N_4482,N_4512);
nor U4781 (N_4781,N_4440,N_4488);
nor U4782 (N_4782,N_4546,N_4513);
and U4783 (N_4783,N_4550,N_4481);
xnor U4784 (N_4784,N_4532,N_4431);
nand U4785 (N_4785,N_4544,N_4460);
nand U4786 (N_4786,N_4401,N_4531);
nor U4787 (N_4787,N_4403,N_4486);
or U4788 (N_4788,N_4475,N_4595);
nor U4789 (N_4789,N_4421,N_4450);
and U4790 (N_4790,N_4558,N_4403);
nor U4791 (N_4791,N_4434,N_4407);
nor U4792 (N_4792,N_4445,N_4595);
and U4793 (N_4793,N_4443,N_4417);
nor U4794 (N_4794,N_4520,N_4559);
and U4795 (N_4795,N_4413,N_4471);
or U4796 (N_4796,N_4553,N_4422);
nor U4797 (N_4797,N_4414,N_4451);
nand U4798 (N_4798,N_4436,N_4559);
nand U4799 (N_4799,N_4590,N_4485);
xnor U4800 (N_4800,N_4635,N_4600);
or U4801 (N_4801,N_4719,N_4727);
and U4802 (N_4802,N_4690,N_4618);
or U4803 (N_4803,N_4636,N_4770);
nor U4804 (N_4804,N_4656,N_4699);
or U4805 (N_4805,N_4718,N_4627);
or U4806 (N_4806,N_4762,N_4711);
xor U4807 (N_4807,N_4693,N_4747);
xor U4808 (N_4808,N_4638,N_4685);
nor U4809 (N_4809,N_4725,N_4796);
nand U4810 (N_4810,N_4776,N_4767);
nand U4811 (N_4811,N_4722,N_4741);
nor U4812 (N_4812,N_4724,N_4705);
xnor U4813 (N_4813,N_4768,N_4620);
and U4814 (N_4814,N_4645,N_4717);
xor U4815 (N_4815,N_4630,N_4673);
or U4816 (N_4816,N_4723,N_4743);
or U4817 (N_4817,N_4646,N_4798);
and U4818 (N_4818,N_4737,N_4754);
nor U4819 (N_4819,N_4748,N_4613);
xor U4820 (N_4820,N_4708,N_4756);
nand U4821 (N_4821,N_4643,N_4652);
xor U4822 (N_4822,N_4650,N_4603);
nand U4823 (N_4823,N_4696,N_4639);
or U4824 (N_4824,N_4788,N_4772);
xnor U4825 (N_4825,N_4732,N_4609);
or U4826 (N_4826,N_4615,N_4612);
nor U4827 (N_4827,N_4780,N_4614);
xnor U4828 (N_4828,N_4771,N_4701);
nor U4829 (N_4829,N_4601,N_4628);
or U4830 (N_4830,N_4766,N_4700);
nor U4831 (N_4831,N_4640,N_4602);
xnor U4832 (N_4832,N_4605,N_4629);
xor U4833 (N_4833,N_4626,N_4774);
and U4834 (N_4834,N_4769,N_4649);
or U4835 (N_4835,N_4714,N_4675);
and U4836 (N_4836,N_4728,N_4784);
xor U4837 (N_4837,N_4757,N_4712);
nand U4838 (N_4838,N_4721,N_4687);
nor U4839 (N_4839,N_4773,N_4716);
or U4840 (N_4840,N_4647,N_4697);
and U4841 (N_4841,N_4642,N_4794);
and U4842 (N_4842,N_4790,N_4793);
xor U4843 (N_4843,N_4678,N_4688);
xor U4844 (N_4844,N_4703,N_4715);
xor U4845 (N_4845,N_4740,N_4755);
or U4846 (N_4846,N_4634,N_4765);
xnor U4847 (N_4847,N_4655,N_4707);
or U4848 (N_4848,N_4742,N_4709);
nand U4849 (N_4849,N_4761,N_4735);
nor U4850 (N_4850,N_4752,N_4713);
and U4851 (N_4851,N_4730,N_4698);
or U4852 (N_4852,N_4624,N_4654);
nand U4853 (N_4853,N_4676,N_4667);
xnor U4854 (N_4854,N_4720,N_4683);
xor U4855 (N_4855,N_4670,N_4669);
nand U4856 (N_4856,N_4674,N_4799);
xnor U4857 (N_4857,N_4759,N_4619);
xnor U4858 (N_4858,N_4651,N_4684);
nand U4859 (N_4859,N_4632,N_4750);
xnor U4860 (N_4860,N_4633,N_4734);
and U4861 (N_4861,N_4672,N_4631);
nand U4862 (N_4862,N_4795,N_4746);
nand U4863 (N_4863,N_4663,N_4691);
or U4864 (N_4864,N_4625,N_4616);
and U4865 (N_4865,N_4682,N_4787);
or U4866 (N_4866,N_4729,N_4610);
or U4867 (N_4867,N_4733,N_4775);
and U4868 (N_4868,N_4782,N_4786);
xor U4869 (N_4869,N_4753,N_4731);
or U4870 (N_4870,N_4738,N_4659);
or U4871 (N_4871,N_4710,N_4665);
nor U4872 (N_4872,N_4695,N_4764);
nor U4873 (N_4873,N_4604,N_4704);
xor U4874 (N_4874,N_4623,N_4657);
xor U4875 (N_4875,N_4744,N_4749);
or U4876 (N_4876,N_4781,N_4661);
xor U4877 (N_4877,N_4622,N_4689);
nand U4878 (N_4878,N_4664,N_4791);
nand U4879 (N_4879,N_4666,N_4637);
nand U4880 (N_4880,N_4658,N_4745);
nor U4881 (N_4881,N_4797,N_4789);
or U4882 (N_4882,N_4792,N_4668);
or U4883 (N_4883,N_4706,N_4778);
nand U4884 (N_4884,N_4763,N_4702);
nand U4885 (N_4885,N_4680,N_4779);
or U4886 (N_4886,N_4606,N_4681);
nor U4887 (N_4887,N_4644,N_4641);
nor U4888 (N_4888,N_4739,N_4671);
xor U4889 (N_4889,N_4648,N_4679);
xor U4890 (N_4890,N_4686,N_4758);
nand U4891 (N_4891,N_4607,N_4653);
nand U4892 (N_4892,N_4660,N_4662);
xor U4893 (N_4893,N_4611,N_4621);
and U4894 (N_4894,N_4736,N_4783);
nor U4895 (N_4895,N_4785,N_4751);
and U4896 (N_4896,N_4694,N_4608);
nand U4897 (N_4897,N_4617,N_4692);
nor U4898 (N_4898,N_4677,N_4760);
nand U4899 (N_4899,N_4777,N_4726);
nand U4900 (N_4900,N_4703,N_4753);
xor U4901 (N_4901,N_4783,N_4729);
xor U4902 (N_4902,N_4709,N_4633);
nor U4903 (N_4903,N_4778,N_4729);
nor U4904 (N_4904,N_4645,N_4626);
or U4905 (N_4905,N_4715,N_4629);
or U4906 (N_4906,N_4659,N_4746);
or U4907 (N_4907,N_4753,N_4722);
or U4908 (N_4908,N_4731,N_4652);
nor U4909 (N_4909,N_4704,N_4743);
and U4910 (N_4910,N_4704,N_4705);
xnor U4911 (N_4911,N_4620,N_4678);
nor U4912 (N_4912,N_4700,N_4693);
nand U4913 (N_4913,N_4656,N_4777);
nand U4914 (N_4914,N_4604,N_4713);
or U4915 (N_4915,N_4737,N_4728);
xnor U4916 (N_4916,N_4659,N_4688);
or U4917 (N_4917,N_4717,N_4609);
nand U4918 (N_4918,N_4714,N_4625);
nor U4919 (N_4919,N_4651,N_4753);
or U4920 (N_4920,N_4766,N_4676);
and U4921 (N_4921,N_4777,N_4732);
nor U4922 (N_4922,N_4755,N_4716);
xor U4923 (N_4923,N_4747,N_4737);
nor U4924 (N_4924,N_4721,N_4634);
nor U4925 (N_4925,N_4662,N_4764);
and U4926 (N_4926,N_4772,N_4770);
or U4927 (N_4927,N_4604,N_4655);
and U4928 (N_4928,N_4729,N_4690);
or U4929 (N_4929,N_4645,N_4622);
and U4930 (N_4930,N_4746,N_4708);
nand U4931 (N_4931,N_4767,N_4689);
and U4932 (N_4932,N_4792,N_4694);
and U4933 (N_4933,N_4615,N_4607);
or U4934 (N_4934,N_4706,N_4671);
nor U4935 (N_4935,N_4726,N_4692);
xor U4936 (N_4936,N_4618,N_4672);
nand U4937 (N_4937,N_4723,N_4750);
xor U4938 (N_4938,N_4769,N_4699);
xor U4939 (N_4939,N_4747,N_4687);
and U4940 (N_4940,N_4739,N_4634);
and U4941 (N_4941,N_4753,N_4603);
xor U4942 (N_4942,N_4624,N_4659);
and U4943 (N_4943,N_4705,N_4711);
nand U4944 (N_4944,N_4627,N_4726);
and U4945 (N_4945,N_4792,N_4644);
nor U4946 (N_4946,N_4703,N_4642);
nor U4947 (N_4947,N_4680,N_4769);
nand U4948 (N_4948,N_4648,N_4710);
nor U4949 (N_4949,N_4794,N_4781);
xnor U4950 (N_4950,N_4737,N_4733);
nand U4951 (N_4951,N_4607,N_4771);
nor U4952 (N_4952,N_4690,N_4771);
nand U4953 (N_4953,N_4640,N_4661);
or U4954 (N_4954,N_4736,N_4615);
nor U4955 (N_4955,N_4635,N_4609);
nand U4956 (N_4956,N_4786,N_4745);
xnor U4957 (N_4957,N_4677,N_4679);
or U4958 (N_4958,N_4768,N_4660);
or U4959 (N_4959,N_4646,N_4682);
and U4960 (N_4960,N_4669,N_4709);
xnor U4961 (N_4961,N_4740,N_4763);
and U4962 (N_4962,N_4742,N_4692);
and U4963 (N_4963,N_4670,N_4608);
and U4964 (N_4964,N_4697,N_4693);
nor U4965 (N_4965,N_4631,N_4662);
xor U4966 (N_4966,N_4683,N_4671);
nand U4967 (N_4967,N_4770,N_4752);
and U4968 (N_4968,N_4619,N_4612);
nor U4969 (N_4969,N_4720,N_4794);
nor U4970 (N_4970,N_4748,N_4686);
or U4971 (N_4971,N_4620,N_4660);
xor U4972 (N_4972,N_4690,N_4654);
xnor U4973 (N_4973,N_4764,N_4787);
nand U4974 (N_4974,N_4738,N_4653);
nor U4975 (N_4975,N_4653,N_4744);
or U4976 (N_4976,N_4772,N_4618);
xnor U4977 (N_4977,N_4600,N_4643);
xnor U4978 (N_4978,N_4723,N_4652);
nor U4979 (N_4979,N_4779,N_4759);
or U4980 (N_4980,N_4767,N_4683);
and U4981 (N_4981,N_4702,N_4619);
nand U4982 (N_4982,N_4659,N_4631);
or U4983 (N_4983,N_4739,N_4639);
xor U4984 (N_4984,N_4653,N_4614);
nor U4985 (N_4985,N_4704,N_4615);
nor U4986 (N_4986,N_4774,N_4777);
or U4987 (N_4987,N_4741,N_4798);
and U4988 (N_4988,N_4743,N_4738);
xnor U4989 (N_4989,N_4642,N_4780);
nand U4990 (N_4990,N_4717,N_4637);
nor U4991 (N_4991,N_4733,N_4645);
xnor U4992 (N_4992,N_4761,N_4784);
nor U4993 (N_4993,N_4769,N_4661);
nand U4994 (N_4994,N_4756,N_4622);
nand U4995 (N_4995,N_4618,N_4790);
and U4996 (N_4996,N_4714,N_4640);
or U4997 (N_4997,N_4690,N_4692);
nand U4998 (N_4998,N_4779,N_4619);
nor U4999 (N_4999,N_4758,N_4743);
and U5000 (N_5000,N_4953,N_4893);
nand U5001 (N_5001,N_4857,N_4907);
nor U5002 (N_5002,N_4887,N_4989);
and U5003 (N_5003,N_4910,N_4878);
and U5004 (N_5004,N_4902,N_4912);
xor U5005 (N_5005,N_4818,N_4832);
nand U5006 (N_5006,N_4801,N_4940);
or U5007 (N_5007,N_4838,N_4969);
nand U5008 (N_5008,N_4917,N_4964);
nand U5009 (N_5009,N_4949,N_4985);
and U5010 (N_5010,N_4869,N_4929);
nand U5011 (N_5011,N_4855,N_4837);
nor U5012 (N_5012,N_4924,N_4821);
or U5013 (N_5013,N_4871,N_4862);
nor U5014 (N_5014,N_4908,N_4941);
or U5015 (N_5015,N_4935,N_4930);
nor U5016 (N_5016,N_4840,N_4931);
and U5017 (N_5017,N_4959,N_4955);
and U5018 (N_5018,N_4879,N_4926);
nand U5019 (N_5019,N_4803,N_4997);
or U5020 (N_5020,N_4944,N_4901);
or U5021 (N_5021,N_4876,N_4916);
nand U5022 (N_5022,N_4937,N_4966);
xor U5023 (N_5023,N_4960,N_4865);
or U5024 (N_5024,N_4823,N_4962);
xor U5025 (N_5025,N_4813,N_4880);
nand U5026 (N_5026,N_4986,N_4973);
nand U5027 (N_5027,N_4928,N_4808);
or U5028 (N_5028,N_4829,N_4965);
nand U5029 (N_5029,N_4812,N_4906);
nand U5030 (N_5030,N_4806,N_4977);
xor U5031 (N_5031,N_4800,N_4830);
nand U5032 (N_5032,N_4927,N_4864);
xnor U5033 (N_5033,N_4888,N_4957);
or U5034 (N_5034,N_4811,N_4992);
and U5035 (N_5035,N_4822,N_4951);
xnor U5036 (N_5036,N_4947,N_4954);
and U5037 (N_5037,N_4886,N_4971);
or U5038 (N_5038,N_4885,N_4833);
or U5039 (N_5039,N_4820,N_4987);
or U5040 (N_5040,N_4828,N_4990);
nor U5041 (N_5041,N_4841,N_4807);
nor U5042 (N_5042,N_4817,N_4943);
nand U5043 (N_5043,N_4974,N_4972);
nor U5044 (N_5044,N_4827,N_4982);
and U5045 (N_5045,N_4881,N_4845);
or U5046 (N_5046,N_4850,N_4980);
xor U5047 (N_5047,N_4895,N_4810);
or U5048 (N_5048,N_4835,N_4995);
nor U5049 (N_5049,N_4853,N_4804);
nand U5050 (N_5050,N_4874,N_4814);
nor U5051 (N_5051,N_4922,N_4923);
xor U5052 (N_5052,N_4898,N_4856);
or U5053 (N_5053,N_4956,N_4999);
xnor U5054 (N_5054,N_4963,N_4860);
nand U5055 (N_5055,N_4915,N_4914);
and U5056 (N_5056,N_4897,N_4852);
xor U5057 (N_5057,N_4920,N_4900);
xnor U5058 (N_5058,N_4842,N_4933);
xor U5059 (N_5059,N_4936,N_4904);
nor U5060 (N_5060,N_4976,N_4945);
xnor U5061 (N_5061,N_4970,N_4934);
xor U5062 (N_5062,N_4925,N_4868);
and U5063 (N_5063,N_4996,N_4875);
nand U5064 (N_5064,N_4942,N_4844);
xor U5065 (N_5065,N_4873,N_4872);
and U5066 (N_5066,N_4913,N_4819);
nand U5067 (N_5067,N_4854,N_4883);
xnor U5068 (N_5068,N_4918,N_4805);
and U5069 (N_5069,N_4884,N_4892);
nand U5070 (N_5070,N_4834,N_4905);
and U5071 (N_5071,N_4858,N_4983);
nor U5072 (N_5072,N_4816,N_4968);
xor U5073 (N_5073,N_4846,N_4809);
nand U5074 (N_5074,N_4952,N_4899);
nand U5075 (N_5075,N_4851,N_4863);
or U5076 (N_5076,N_4975,N_4877);
or U5077 (N_5077,N_4998,N_4978);
xor U5078 (N_5078,N_4870,N_4866);
and U5079 (N_5079,N_4939,N_4938);
xor U5080 (N_5080,N_4802,N_4909);
nand U5081 (N_5081,N_4946,N_4831);
or U5082 (N_5082,N_4921,N_4948);
xnor U5083 (N_5083,N_4981,N_4979);
nand U5084 (N_5084,N_4889,N_4826);
and U5085 (N_5085,N_4911,N_4894);
xnor U5086 (N_5086,N_4836,N_4896);
nor U5087 (N_5087,N_4994,N_4839);
xor U5088 (N_5088,N_4967,N_4991);
xnor U5089 (N_5089,N_4824,N_4993);
nand U5090 (N_5090,N_4932,N_4849);
xnor U5091 (N_5091,N_4988,N_4815);
xnor U5092 (N_5092,N_4919,N_4950);
nor U5093 (N_5093,N_4891,N_4825);
or U5094 (N_5094,N_4958,N_4847);
nor U5095 (N_5095,N_4843,N_4984);
nand U5096 (N_5096,N_4861,N_4903);
xor U5097 (N_5097,N_4890,N_4882);
nor U5098 (N_5098,N_4867,N_4848);
nand U5099 (N_5099,N_4961,N_4859);
and U5100 (N_5100,N_4908,N_4958);
nor U5101 (N_5101,N_4906,N_4888);
nand U5102 (N_5102,N_4846,N_4858);
nor U5103 (N_5103,N_4932,N_4908);
xnor U5104 (N_5104,N_4804,N_4831);
and U5105 (N_5105,N_4893,N_4811);
xnor U5106 (N_5106,N_4971,N_4943);
and U5107 (N_5107,N_4895,N_4959);
or U5108 (N_5108,N_4820,N_4898);
or U5109 (N_5109,N_4978,N_4854);
or U5110 (N_5110,N_4908,N_4905);
nor U5111 (N_5111,N_4878,N_4906);
nand U5112 (N_5112,N_4928,N_4972);
and U5113 (N_5113,N_4987,N_4947);
or U5114 (N_5114,N_4848,N_4868);
xnor U5115 (N_5115,N_4806,N_4933);
nand U5116 (N_5116,N_4931,N_4809);
or U5117 (N_5117,N_4932,N_4991);
nand U5118 (N_5118,N_4931,N_4941);
nor U5119 (N_5119,N_4860,N_4902);
and U5120 (N_5120,N_4801,N_4896);
and U5121 (N_5121,N_4841,N_4853);
nor U5122 (N_5122,N_4951,N_4981);
nand U5123 (N_5123,N_4846,N_4895);
nand U5124 (N_5124,N_4842,N_4869);
nor U5125 (N_5125,N_4899,N_4908);
and U5126 (N_5126,N_4896,N_4887);
nand U5127 (N_5127,N_4951,N_4845);
xnor U5128 (N_5128,N_4853,N_4852);
or U5129 (N_5129,N_4865,N_4913);
and U5130 (N_5130,N_4979,N_4832);
xor U5131 (N_5131,N_4966,N_4957);
nor U5132 (N_5132,N_4954,N_4888);
nand U5133 (N_5133,N_4976,N_4824);
or U5134 (N_5134,N_4950,N_4839);
xor U5135 (N_5135,N_4847,N_4810);
xnor U5136 (N_5136,N_4922,N_4882);
xor U5137 (N_5137,N_4870,N_4910);
xnor U5138 (N_5138,N_4992,N_4939);
nor U5139 (N_5139,N_4956,N_4821);
nor U5140 (N_5140,N_4939,N_4891);
xor U5141 (N_5141,N_4988,N_4879);
nand U5142 (N_5142,N_4972,N_4927);
and U5143 (N_5143,N_4849,N_4836);
and U5144 (N_5144,N_4814,N_4934);
or U5145 (N_5145,N_4878,N_4956);
xor U5146 (N_5146,N_4899,N_4885);
xnor U5147 (N_5147,N_4982,N_4913);
or U5148 (N_5148,N_4870,N_4850);
nand U5149 (N_5149,N_4980,N_4998);
nor U5150 (N_5150,N_4874,N_4934);
nor U5151 (N_5151,N_4978,N_4945);
xnor U5152 (N_5152,N_4967,N_4979);
or U5153 (N_5153,N_4944,N_4874);
or U5154 (N_5154,N_4836,N_4926);
nor U5155 (N_5155,N_4828,N_4819);
or U5156 (N_5156,N_4883,N_4987);
nand U5157 (N_5157,N_4985,N_4892);
nor U5158 (N_5158,N_4908,N_4844);
nand U5159 (N_5159,N_4808,N_4958);
and U5160 (N_5160,N_4807,N_4842);
nand U5161 (N_5161,N_4905,N_4804);
and U5162 (N_5162,N_4857,N_4915);
or U5163 (N_5163,N_4816,N_4946);
and U5164 (N_5164,N_4843,N_4970);
nor U5165 (N_5165,N_4815,N_4824);
or U5166 (N_5166,N_4961,N_4842);
or U5167 (N_5167,N_4824,N_4877);
or U5168 (N_5168,N_4970,N_4873);
nor U5169 (N_5169,N_4828,N_4863);
and U5170 (N_5170,N_4941,N_4987);
nor U5171 (N_5171,N_4806,N_4805);
nor U5172 (N_5172,N_4924,N_4908);
or U5173 (N_5173,N_4999,N_4851);
xnor U5174 (N_5174,N_4812,N_4951);
and U5175 (N_5175,N_4992,N_4842);
xor U5176 (N_5176,N_4952,N_4943);
nor U5177 (N_5177,N_4921,N_4802);
and U5178 (N_5178,N_4996,N_4958);
nand U5179 (N_5179,N_4803,N_4844);
nand U5180 (N_5180,N_4915,N_4830);
and U5181 (N_5181,N_4828,N_4900);
nand U5182 (N_5182,N_4876,N_4846);
or U5183 (N_5183,N_4843,N_4830);
and U5184 (N_5184,N_4909,N_4873);
and U5185 (N_5185,N_4927,N_4973);
and U5186 (N_5186,N_4918,N_4972);
or U5187 (N_5187,N_4933,N_4901);
nor U5188 (N_5188,N_4955,N_4958);
nand U5189 (N_5189,N_4904,N_4920);
nand U5190 (N_5190,N_4811,N_4885);
or U5191 (N_5191,N_4864,N_4805);
nor U5192 (N_5192,N_4870,N_4803);
xnor U5193 (N_5193,N_4840,N_4933);
and U5194 (N_5194,N_4928,N_4852);
nand U5195 (N_5195,N_4952,N_4985);
or U5196 (N_5196,N_4993,N_4888);
nand U5197 (N_5197,N_4931,N_4885);
xnor U5198 (N_5198,N_4964,N_4860);
nor U5199 (N_5199,N_4961,N_4979);
xnor U5200 (N_5200,N_5026,N_5005);
nand U5201 (N_5201,N_5088,N_5012);
or U5202 (N_5202,N_5126,N_5024);
xor U5203 (N_5203,N_5098,N_5111);
xor U5204 (N_5204,N_5148,N_5171);
and U5205 (N_5205,N_5029,N_5145);
and U5206 (N_5206,N_5123,N_5032);
xnor U5207 (N_5207,N_5187,N_5020);
and U5208 (N_5208,N_5006,N_5066);
and U5209 (N_5209,N_5089,N_5146);
nand U5210 (N_5210,N_5159,N_5047);
and U5211 (N_5211,N_5114,N_5154);
nand U5212 (N_5212,N_5158,N_5097);
xnor U5213 (N_5213,N_5196,N_5186);
nor U5214 (N_5214,N_5194,N_5081);
nand U5215 (N_5215,N_5136,N_5071);
xnor U5216 (N_5216,N_5011,N_5049);
or U5217 (N_5217,N_5134,N_5162);
or U5218 (N_5218,N_5075,N_5058);
nand U5219 (N_5219,N_5142,N_5083);
nor U5220 (N_5220,N_5082,N_5040);
xnor U5221 (N_5221,N_5163,N_5110);
xor U5222 (N_5222,N_5055,N_5165);
and U5223 (N_5223,N_5008,N_5117);
and U5224 (N_5224,N_5156,N_5042);
or U5225 (N_5225,N_5067,N_5027);
xor U5226 (N_5226,N_5193,N_5072);
nor U5227 (N_5227,N_5153,N_5175);
nor U5228 (N_5228,N_5091,N_5016);
nand U5229 (N_5229,N_5178,N_5167);
nand U5230 (N_5230,N_5060,N_5090);
or U5231 (N_5231,N_5043,N_5144);
xnor U5232 (N_5232,N_5122,N_5003);
nand U5233 (N_5233,N_5100,N_5118);
and U5234 (N_5234,N_5061,N_5080);
nand U5235 (N_5235,N_5093,N_5199);
xnor U5236 (N_5236,N_5127,N_5069);
nand U5237 (N_5237,N_5197,N_5044);
nor U5238 (N_5238,N_5129,N_5056);
xor U5239 (N_5239,N_5119,N_5021);
and U5240 (N_5240,N_5076,N_5050);
xnor U5241 (N_5241,N_5007,N_5180);
xor U5242 (N_5242,N_5086,N_5065);
or U5243 (N_5243,N_5062,N_5130);
xor U5244 (N_5244,N_5189,N_5140);
nand U5245 (N_5245,N_5131,N_5137);
and U5246 (N_5246,N_5079,N_5157);
or U5247 (N_5247,N_5188,N_5172);
and U5248 (N_5248,N_5115,N_5033);
nand U5249 (N_5249,N_5169,N_5028);
and U5250 (N_5250,N_5143,N_5113);
xnor U5251 (N_5251,N_5063,N_5170);
nor U5252 (N_5252,N_5174,N_5035);
and U5253 (N_5253,N_5070,N_5077);
or U5254 (N_5254,N_5096,N_5101);
or U5255 (N_5255,N_5030,N_5051);
nor U5256 (N_5256,N_5017,N_5173);
xor U5257 (N_5257,N_5116,N_5135);
xor U5258 (N_5258,N_5022,N_5160);
or U5259 (N_5259,N_5181,N_5120);
and U5260 (N_5260,N_5023,N_5039);
and U5261 (N_5261,N_5191,N_5184);
and U5262 (N_5262,N_5068,N_5124);
or U5263 (N_5263,N_5045,N_5053);
or U5264 (N_5264,N_5106,N_5168);
or U5265 (N_5265,N_5064,N_5103);
and U5266 (N_5266,N_5176,N_5048);
xnor U5267 (N_5267,N_5152,N_5085);
and U5268 (N_5268,N_5092,N_5031);
nor U5269 (N_5269,N_5149,N_5182);
and U5270 (N_5270,N_5094,N_5059);
xnor U5271 (N_5271,N_5192,N_5179);
nor U5272 (N_5272,N_5037,N_5147);
nor U5273 (N_5273,N_5002,N_5001);
xor U5274 (N_5274,N_5010,N_5038);
or U5275 (N_5275,N_5133,N_5041);
nand U5276 (N_5276,N_5155,N_5015);
nor U5277 (N_5277,N_5084,N_5074);
nand U5278 (N_5278,N_5109,N_5107);
and U5279 (N_5279,N_5166,N_5190);
nor U5280 (N_5280,N_5102,N_5099);
and U5281 (N_5281,N_5141,N_5132);
xor U5282 (N_5282,N_5000,N_5087);
nor U5283 (N_5283,N_5177,N_5138);
or U5284 (N_5284,N_5161,N_5128);
nand U5285 (N_5285,N_5025,N_5054);
or U5286 (N_5286,N_5078,N_5073);
or U5287 (N_5287,N_5198,N_5004);
xor U5288 (N_5288,N_5108,N_5057);
and U5289 (N_5289,N_5009,N_5018);
and U5290 (N_5290,N_5139,N_5046);
and U5291 (N_5291,N_5164,N_5019);
and U5292 (N_5292,N_5185,N_5151);
xor U5293 (N_5293,N_5105,N_5014);
and U5294 (N_5294,N_5036,N_5150);
xnor U5295 (N_5295,N_5034,N_5121);
nor U5296 (N_5296,N_5052,N_5095);
nor U5297 (N_5297,N_5112,N_5125);
xor U5298 (N_5298,N_5104,N_5183);
and U5299 (N_5299,N_5013,N_5195);
nand U5300 (N_5300,N_5129,N_5186);
nor U5301 (N_5301,N_5162,N_5032);
xnor U5302 (N_5302,N_5014,N_5184);
xor U5303 (N_5303,N_5045,N_5055);
nor U5304 (N_5304,N_5030,N_5153);
or U5305 (N_5305,N_5077,N_5185);
nor U5306 (N_5306,N_5058,N_5009);
xor U5307 (N_5307,N_5019,N_5088);
and U5308 (N_5308,N_5056,N_5001);
nor U5309 (N_5309,N_5186,N_5141);
nand U5310 (N_5310,N_5039,N_5108);
nor U5311 (N_5311,N_5053,N_5029);
or U5312 (N_5312,N_5011,N_5127);
and U5313 (N_5313,N_5100,N_5099);
and U5314 (N_5314,N_5086,N_5187);
nor U5315 (N_5315,N_5009,N_5129);
and U5316 (N_5316,N_5049,N_5071);
and U5317 (N_5317,N_5050,N_5060);
xnor U5318 (N_5318,N_5192,N_5133);
or U5319 (N_5319,N_5158,N_5029);
nand U5320 (N_5320,N_5076,N_5034);
nor U5321 (N_5321,N_5150,N_5100);
nor U5322 (N_5322,N_5156,N_5088);
or U5323 (N_5323,N_5108,N_5032);
nand U5324 (N_5324,N_5104,N_5122);
xor U5325 (N_5325,N_5154,N_5030);
xnor U5326 (N_5326,N_5108,N_5157);
nand U5327 (N_5327,N_5184,N_5125);
nor U5328 (N_5328,N_5100,N_5190);
nor U5329 (N_5329,N_5188,N_5018);
xnor U5330 (N_5330,N_5116,N_5014);
or U5331 (N_5331,N_5065,N_5031);
xnor U5332 (N_5332,N_5061,N_5148);
or U5333 (N_5333,N_5069,N_5155);
xor U5334 (N_5334,N_5166,N_5045);
nand U5335 (N_5335,N_5074,N_5193);
nand U5336 (N_5336,N_5085,N_5167);
nand U5337 (N_5337,N_5199,N_5034);
xor U5338 (N_5338,N_5081,N_5111);
nor U5339 (N_5339,N_5094,N_5109);
xor U5340 (N_5340,N_5189,N_5115);
xnor U5341 (N_5341,N_5114,N_5081);
or U5342 (N_5342,N_5026,N_5189);
nor U5343 (N_5343,N_5007,N_5137);
xnor U5344 (N_5344,N_5162,N_5076);
or U5345 (N_5345,N_5135,N_5044);
or U5346 (N_5346,N_5090,N_5111);
and U5347 (N_5347,N_5112,N_5126);
and U5348 (N_5348,N_5076,N_5008);
or U5349 (N_5349,N_5185,N_5175);
nor U5350 (N_5350,N_5067,N_5129);
and U5351 (N_5351,N_5110,N_5075);
or U5352 (N_5352,N_5057,N_5162);
and U5353 (N_5353,N_5067,N_5181);
xor U5354 (N_5354,N_5161,N_5139);
or U5355 (N_5355,N_5108,N_5176);
nand U5356 (N_5356,N_5010,N_5028);
xnor U5357 (N_5357,N_5146,N_5111);
nor U5358 (N_5358,N_5136,N_5061);
nor U5359 (N_5359,N_5071,N_5081);
and U5360 (N_5360,N_5048,N_5077);
and U5361 (N_5361,N_5053,N_5136);
nand U5362 (N_5362,N_5099,N_5119);
or U5363 (N_5363,N_5067,N_5154);
nand U5364 (N_5364,N_5093,N_5098);
or U5365 (N_5365,N_5078,N_5048);
or U5366 (N_5366,N_5012,N_5177);
nand U5367 (N_5367,N_5036,N_5102);
or U5368 (N_5368,N_5169,N_5062);
and U5369 (N_5369,N_5180,N_5117);
and U5370 (N_5370,N_5169,N_5181);
and U5371 (N_5371,N_5178,N_5189);
and U5372 (N_5372,N_5129,N_5073);
xnor U5373 (N_5373,N_5048,N_5060);
xnor U5374 (N_5374,N_5059,N_5054);
nand U5375 (N_5375,N_5103,N_5065);
nand U5376 (N_5376,N_5190,N_5197);
xor U5377 (N_5377,N_5027,N_5189);
and U5378 (N_5378,N_5194,N_5062);
nand U5379 (N_5379,N_5002,N_5039);
nor U5380 (N_5380,N_5023,N_5146);
xnor U5381 (N_5381,N_5169,N_5117);
xor U5382 (N_5382,N_5164,N_5148);
and U5383 (N_5383,N_5195,N_5110);
and U5384 (N_5384,N_5054,N_5140);
nand U5385 (N_5385,N_5093,N_5013);
or U5386 (N_5386,N_5145,N_5136);
nor U5387 (N_5387,N_5149,N_5008);
nor U5388 (N_5388,N_5170,N_5094);
xor U5389 (N_5389,N_5128,N_5188);
or U5390 (N_5390,N_5066,N_5189);
nor U5391 (N_5391,N_5070,N_5109);
xnor U5392 (N_5392,N_5164,N_5126);
nand U5393 (N_5393,N_5101,N_5127);
nor U5394 (N_5394,N_5026,N_5146);
and U5395 (N_5395,N_5053,N_5014);
nand U5396 (N_5396,N_5116,N_5124);
xor U5397 (N_5397,N_5160,N_5076);
nor U5398 (N_5398,N_5092,N_5079);
xor U5399 (N_5399,N_5155,N_5001);
xnor U5400 (N_5400,N_5260,N_5374);
or U5401 (N_5401,N_5380,N_5350);
nor U5402 (N_5402,N_5268,N_5275);
nand U5403 (N_5403,N_5397,N_5384);
and U5404 (N_5404,N_5265,N_5230);
and U5405 (N_5405,N_5386,N_5359);
xnor U5406 (N_5406,N_5222,N_5269);
nand U5407 (N_5407,N_5321,N_5361);
nor U5408 (N_5408,N_5319,N_5231);
and U5409 (N_5409,N_5390,N_5335);
nor U5410 (N_5410,N_5342,N_5371);
nor U5411 (N_5411,N_5398,N_5360);
and U5412 (N_5412,N_5343,N_5340);
nand U5413 (N_5413,N_5225,N_5202);
nor U5414 (N_5414,N_5250,N_5239);
nand U5415 (N_5415,N_5259,N_5338);
and U5416 (N_5416,N_5216,N_5238);
or U5417 (N_5417,N_5292,N_5248);
nand U5418 (N_5418,N_5389,N_5363);
or U5419 (N_5419,N_5304,N_5305);
and U5420 (N_5420,N_5296,N_5328);
nor U5421 (N_5421,N_5249,N_5388);
nor U5422 (N_5422,N_5283,N_5278);
nor U5423 (N_5423,N_5209,N_5232);
and U5424 (N_5424,N_5309,N_5364);
xor U5425 (N_5425,N_5205,N_5226);
and U5426 (N_5426,N_5312,N_5351);
or U5427 (N_5427,N_5313,N_5208);
or U5428 (N_5428,N_5348,N_5333);
xor U5429 (N_5429,N_5323,N_5317);
nand U5430 (N_5430,N_5284,N_5293);
nor U5431 (N_5431,N_5372,N_5396);
or U5432 (N_5432,N_5233,N_5214);
xor U5433 (N_5433,N_5315,N_5266);
xor U5434 (N_5434,N_5382,N_5242);
nand U5435 (N_5435,N_5316,N_5310);
or U5436 (N_5436,N_5224,N_5279);
nor U5437 (N_5437,N_5287,N_5289);
and U5438 (N_5438,N_5339,N_5379);
nor U5439 (N_5439,N_5356,N_5277);
nand U5440 (N_5440,N_5353,N_5307);
nand U5441 (N_5441,N_5206,N_5299);
and U5442 (N_5442,N_5253,N_5294);
nand U5443 (N_5443,N_5377,N_5271);
nor U5444 (N_5444,N_5203,N_5282);
and U5445 (N_5445,N_5347,N_5220);
nand U5446 (N_5446,N_5276,N_5244);
xnor U5447 (N_5447,N_5327,N_5358);
and U5448 (N_5448,N_5332,N_5375);
nand U5449 (N_5449,N_5320,N_5236);
or U5450 (N_5450,N_5211,N_5223);
and U5451 (N_5451,N_5280,N_5345);
nand U5452 (N_5452,N_5393,N_5241);
or U5453 (N_5453,N_5235,N_5337);
nor U5454 (N_5454,N_5325,N_5263);
and U5455 (N_5455,N_5281,N_5395);
xnor U5456 (N_5456,N_5212,N_5267);
and U5457 (N_5457,N_5301,N_5258);
or U5458 (N_5458,N_5368,N_5246);
nor U5459 (N_5459,N_5392,N_5354);
xnor U5460 (N_5460,N_5257,N_5251);
nand U5461 (N_5461,N_5352,N_5385);
and U5462 (N_5462,N_5262,N_5272);
xor U5463 (N_5463,N_5245,N_5273);
or U5464 (N_5464,N_5391,N_5215);
nand U5465 (N_5465,N_5344,N_5213);
nor U5466 (N_5466,N_5228,N_5331);
nand U5467 (N_5467,N_5298,N_5218);
nor U5468 (N_5468,N_5314,N_5219);
or U5469 (N_5469,N_5297,N_5373);
xnor U5470 (N_5470,N_5394,N_5229);
nor U5471 (N_5471,N_5300,N_5200);
or U5472 (N_5472,N_5306,N_5210);
or U5473 (N_5473,N_5311,N_5274);
or U5474 (N_5474,N_5252,N_5201);
or U5475 (N_5475,N_5336,N_5378);
xnor U5476 (N_5476,N_5329,N_5288);
nor U5477 (N_5477,N_5308,N_5207);
xnor U5478 (N_5478,N_5341,N_5221);
or U5479 (N_5479,N_5318,N_5291);
or U5480 (N_5480,N_5234,N_5247);
and U5481 (N_5481,N_5330,N_5322);
xnor U5482 (N_5482,N_5302,N_5254);
xor U5483 (N_5483,N_5286,N_5237);
nor U5484 (N_5484,N_5387,N_5362);
and U5485 (N_5485,N_5217,N_5264);
nor U5486 (N_5486,N_5376,N_5256);
or U5487 (N_5487,N_5365,N_5204);
nand U5488 (N_5488,N_5370,N_5399);
nor U5489 (N_5489,N_5303,N_5381);
nor U5490 (N_5490,N_5357,N_5355);
nor U5491 (N_5491,N_5227,N_5243);
xor U5492 (N_5492,N_5366,N_5383);
nor U5493 (N_5493,N_5326,N_5295);
or U5494 (N_5494,N_5369,N_5290);
or U5495 (N_5495,N_5270,N_5349);
xnor U5496 (N_5496,N_5255,N_5324);
nor U5497 (N_5497,N_5334,N_5285);
or U5498 (N_5498,N_5346,N_5367);
nor U5499 (N_5499,N_5261,N_5240);
and U5500 (N_5500,N_5202,N_5319);
nor U5501 (N_5501,N_5341,N_5294);
or U5502 (N_5502,N_5209,N_5346);
nor U5503 (N_5503,N_5336,N_5334);
xor U5504 (N_5504,N_5294,N_5286);
and U5505 (N_5505,N_5331,N_5213);
or U5506 (N_5506,N_5257,N_5240);
and U5507 (N_5507,N_5373,N_5204);
and U5508 (N_5508,N_5344,N_5223);
xor U5509 (N_5509,N_5302,N_5275);
or U5510 (N_5510,N_5257,N_5303);
and U5511 (N_5511,N_5299,N_5347);
or U5512 (N_5512,N_5302,N_5238);
or U5513 (N_5513,N_5231,N_5236);
nor U5514 (N_5514,N_5379,N_5334);
nor U5515 (N_5515,N_5312,N_5284);
and U5516 (N_5516,N_5294,N_5399);
nor U5517 (N_5517,N_5238,N_5315);
nor U5518 (N_5518,N_5254,N_5320);
nor U5519 (N_5519,N_5393,N_5213);
xor U5520 (N_5520,N_5311,N_5355);
or U5521 (N_5521,N_5231,N_5287);
or U5522 (N_5522,N_5209,N_5396);
nor U5523 (N_5523,N_5242,N_5385);
and U5524 (N_5524,N_5243,N_5294);
and U5525 (N_5525,N_5311,N_5220);
nor U5526 (N_5526,N_5269,N_5260);
xor U5527 (N_5527,N_5341,N_5230);
and U5528 (N_5528,N_5271,N_5290);
xnor U5529 (N_5529,N_5362,N_5247);
xnor U5530 (N_5530,N_5294,N_5335);
xor U5531 (N_5531,N_5267,N_5350);
nor U5532 (N_5532,N_5319,N_5381);
nor U5533 (N_5533,N_5322,N_5344);
and U5534 (N_5534,N_5256,N_5302);
nor U5535 (N_5535,N_5247,N_5211);
xnor U5536 (N_5536,N_5280,N_5376);
and U5537 (N_5537,N_5278,N_5248);
and U5538 (N_5538,N_5282,N_5269);
nor U5539 (N_5539,N_5346,N_5325);
or U5540 (N_5540,N_5359,N_5321);
nor U5541 (N_5541,N_5210,N_5347);
xor U5542 (N_5542,N_5318,N_5261);
and U5543 (N_5543,N_5333,N_5391);
nand U5544 (N_5544,N_5319,N_5351);
xor U5545 (N_5545,N_5395,N_5300);
xor U5546 (N_5546,N_5393,N_5206);
nand U5547 (N_5547,N_5388,N_5390);
nor U5548 (N_5548,N_5308,N_5373);
or U5549 (N_5549,N_5370,N_5342);
nand U5550 (N_5550,N_5273,N_5334);
nand U5551 (N_5551,N_5248,N_5372);
nor U5552 (N_5552,N_5305,N_5264);
xnor U5553 (N_5553,N_5345,N_5347);
xnor U5554 (N_5554,N_5246,N_5336);
nand U5555 (N_5555,N_5385,N_5360);
xnor U5556 (N_5556,N_5288,N_5259);
nand U5557 (N_5557,N_5235,N_5202);
nor U5558 (N_5558,N_5224,N_5231);
nor U5559 (N_5559,N_5391,N_5352);
xor U5560 (N_5560,N_5390,N_5213);
xnor U5561 (N_5561,N_5234,N_5324);
and U5562 (N_5562,N_5378,N_5257);
or U5563 (N_5563,N_5353,N_5297);
and U5564 (N_5564,N_5394,N_5277);
nor U5565 (N_5565,N_5353,N_5316);
nor U5566 (N_5566,N_5330,N_5391);
and U5567 (N_5567,N_5356,N_5339);
nor U5568 (N_5568,N_5207,N_5321);
nor U5569 (N_5569,N_5294,N_5267);
xor U5570 (N_5570,N_5386,N_5338);
nand U5571 (N_5571,N_5215,N_5346);
nor U5572 (N_5572,N_5384,N_5291);
xor U5573 (N_5573,N_5283,N_5323);
and U5574 (N_5574,N_5246,N_5393);
nand U5575 (N_5575,N_5317,N_5310);
nand U5576 (N_5576,N_5305,N_5207);
or U5577 (N_5577,N_5355,N_5254);
and U5578 (N_5578,N_5321,N_5325);
nand U5579 (N_5579,N_5312,N_5286);
xnor U5580 (N_5580,N_5215,N_5350);
xnor U5581 (N_5581,N_5355,N_5244);
nand U5582 (N_5582,N_5252,N_5380);
and U5583 (N_5583,N_5246,N_5335);
or U5584 (N_5584,N_5362,N_5279);
xnor U5585 (N_5585,N_5335,N_5284);
nand U5586 (N_5586,N_5376,N_5207);
nor U5587 (N_5587,N_5242,N_5264);
xnor U5588 (N_5588,N_5291,N_5284);
nand U5589 (N_5589,N_5265,N_5256);
xor U5590 (N_5590,N_5396,N_5346);
nor U5591 (N_5591,N_5332,N_5279);
nand U5592 (N_5592,N_5284,N_5238);
or U5593 (N_5593,N_5343,N_5395);
xnor U5594 (N_5594,N_5289,N_5250);
nor U5595 (N_5595,N_5208,N_5229);
nor U5596 (N_5596,N_5363,N_5327);
nand U5597 (N_5597,N_5280,N_5299);
nor U5598 (N_5598,N_5312,N_5213);
nor U5599 (N_5599,N_5332,N_5291);
nor U5600 (N_5600,N_5570,N_5519);
xnor U5601 (N_5601,N_5430,N_5477);
or U5602 (N_5602,N_5539,N_5426);
nor U5603 (N_5603,N_5427,N_5450);
xor U5604 (N_5604,N_5428,N_5495);
and U5605 (N_5605,N_5599,N_5445);
xnor U5606 (N_5606,N_5520,N_5589);
xor U5607 (N_5607,N_5423,N_5444);
or U5608 (N_5608,N_5455,N_5437);
and U5609 (N_5609,N_5544,N_5530);
nand U5610 (N_5610,N_5541,N_5497);
nand U5611 (N_5611,N_5559,N_5419);
and U5612 (N_5612,N_5417,N_5583);
xnor U5613 (N_5613,N_5542,N_5564);
or U5614 (N_5614,N_5527,N_5479);
xnor U5615 (N_5615,N_5524,N_5441);
nand U5616 (N_5616,N_5503,N_5529);
nor U5617 (N_5617,N_5482,N_5490);
or U5618 (N_5618,N_5401,N_5443);
nor U5619 (N_5619,N_5573,N_5509);
and U5620 (N_5620,N_5436,N_5439);
or U5621 (N_5621,N_5594,N_5448);
nand U5622 (N_5622,N_5536,N_5484);
or U5623 (N_5623,N_5476,N_5410);
and U5624 (N_5624,N_5502,N_5449);
and U5625 (N_5625,N_5429,N_5596);
or U5626 (N_5626,N_5563,N_5560);
or U5627 (N_5627,N_5518,N_5404);
nor U5628 (N_5628,N_5505,N_5512);
nand U5629 (N_5629,N_5451,N_5470);
nor U5630 (N_5630,N_5584,N_5549);
and U5631 (N_5631,N_5442,N_5492);
or U5632 (N_5632,N_5532,N_5491);
nand U5633 (N_5633,N_5574,N_5597);
and U5634 (N_5634,N_5481,N_5551);
nor U5635 (N_5635,N_5561,N_5433);
and U5636 (N_5636,N_5538,N_5454);
nand U5637 (N_5637,N_5463,N_5587);
nor U5638 (N_5638,N_5489,N_5571);
nand U5639 (N_5639,N_5420,N_5461);
xnor U5640 (N_5640,N_5562,N_5456);
and U5641 (N_5641,N_5501,N_5438);
xnor U5642 (N_5642,N_5440,N_5507);
nand U5643 (N_5643,N_5468,N_5506);
nor U5644 (N_5644,N_5565,N_5431);
or U5645 (N_5645,N_5494,N_5554);
nand U5646 (N_5646,N_5557,N_5408);
nor U5647 (N_5647,N_5525,N_5471);
nor U5648 (N_5648,N_5446,N_5472);
xor U5649 (N_5649,N_5535,N_5550);
xnor U5650 (N_5650,N_5558,N_5407);
and U5651 (N_5651,N_5432,N_5511);
and U5652 (N_5652,N_5422,N_5434);
and U5653 (N_5653,N_5590,N_5547);
xnor U5654 (N_5654,N_5413,N_5435);
and U5655 (N_5655,N_5466,N_5460);
and U5656 (N_5656,N_5457,N_5510);
xor U5657 (N_5657,N_5415,N_5516);
xor U5658 (N_5658,N_5568,N_5425);
and U5659 (N_5659,N_5575,N_5580);
xor U5660 (N_5660,N_5552,N_5537);
or U5661 (N_5661,N_5412,N_5416);
or U5662 (N_5662,N_5486,N_5414);
nand U5663 (N_5663,N_5402,N_5540);
nor U5664 (N_5664,N_5500,N_5499);
or U5665 (N_5665,N_5504,N_5493);
nor U5666 (N_5666,N_5452,N_5548);
nand U5667 (N_5667,N_5588,N_5582);
nand U5668 (N_5668,N_5513,N_5483);
xnor U5669 (N_5669,N_5523,N_5487);
nand U5670 (N_5670,N_5534,N_5464);
nor U5671 (N_5671,N_5531,N_5555);
xor U5672 (N_5672,N_5598,N_5400);
nand U5673 (N_5673,N_5475,N_5403);
and U5674 (N_5674,N_5556,N_5453);
or U5675 (N_5675,N_5478,N_5480);
and U5676 (N_5676,N_5514,N_5474);
and U5677 (N_5677,N_5469,N_5496);
nor U5678 (N_5678,N_5517,N_5498);
nor U5679 (N_5679,N_5578,N_5577);
nand U5680 (N_5680,N_5508,N_5553);
nor U5681 (N_5681,N_5567,N_5488);
or U5682 (N_5682,N_5406,N_5515);
and U5683 (N_5683,N_5533,N_5421);
xor U5684 (N_5684,N_5592,N_5576);
or U5685 (N_5685,N_5546,N_5521);
and U5686 (N_5686,N_5526,N_5586);
xnor U5687 (N_5687,N_5595,N_5522);
nand U5688 (N_5688,N_5405,N_5409);
xor U5689 (N_5689,N_5581,N_5543);
and U5690 (N_5690,N_5593,N_5572);
xnor U5691 (N_5691,N_5459,N_5447);
nand U5692 (N_5692,N_5458,N_5424);
and U5693 (N_5693,N_5418,N_5566);
nand U5694 (N_5694,N_5528,N_5585);
and U5695 (N_5695,N_5485,N_5545);
nand U5696 (N_5696,N_5579,N_5467);
nor U5697 (N_5697,N_5411,N_5473);
xnor U5698 (N_5698,N_5465,N_5569);
and U5699 (N_5699,N_5591,N_5462);
and U5700 (N_5700,N_5498,N_5571);
or U5701 (N_5701,N_5481,N_5576);
and U5702 (N_5702,N_5518,N_5466);
nor U5703 (N_5703,N_5570,N_5400);
or U5704 (N_5704,N_5551,N_5465);
and U5705 (N_5705,N_5554,N_5503);
nor U5706 (N_5706,N_5430,N_5451);
and U5707 (N_5707,N_5515,N_5539);
xnor U5708 (N_5708,N_5519,N_5598);
and U5709 (N_5709,N_5450,N_5503);
nor U5710 (N_5710,N_5467,N_5543);
nor U5711 (N_5711,N_5598,N_5430);
nand U5712 (N_5712,N_5478,N_5407);
nor U5713 (N_5713,N_5555,N_5570);
xnor U5714 (N_5714,N_5558,N_5540);
xnor U5715 (N_5715,N_5507,N_5559);
nor U5716 (N_5716,N_5404,N_5570);
nand U5717 (N_5717,N_5400,N_5507);
xor U5718 (N_5718,N_5550,N_5505);
and U5719 (N_5719,N_5508,N_5426);
nor U5720 (N_5720,N_5505,N_5584);
nand U5721 (N_5721,N_5465,N_5451);
or U5722 (N_5722,N_5443,N_5412);
xor U5723 (N_5723,N_5568,N_5492);
xnor U5724 (N_5724,N_5407,N_5403);
and U5725 (N_5725,N_5455,N_5570);
nand U5726 (N_5726,N_5588,N_5488);
xnor U5727 (N_5727,N_5542,N_5451);
xnor U5728 (N_5728,N_5592,N_5420);
or U5729 (N_5729,N_5462,N_5565);
or U5730 (N_5730,N_5572,N_5569);
and U5731 (N_5731,N_5540,N_5428);
or U5732 (N_5732,N_5480,N_5412);
and U5733 (N_5733,N_5559,N_5556);
or U5734 (N_5734,N_5523,N_5499);
nand U5735 (N_5735,N_5549,N_5435);
nor U5736 (N_5736,N_5482,N_5597);
or U5737 (N_5737,N_5565,N_5437);
or U5738 (N_5738,N_5445,N_5539);
nor U5739 (N_5739,N_5456,N_5472);
nand U5740 (N_5740,N_5465,N_5594);
and U5741 (N_5741,N_5411,N_5565);
xor U5742 (N_5742,N_5585,N_5571);
and U5743 (N_5743,N_5458,N_5544);
and U5744 (N_5744,N_5422,N_5556);
nor U5745 (N_5745,N_5428,N_5574);
nand U5746 (N_5746,N_5400,N_5563);
xor U5747 (N_5747,N_5479,N_5568);
and U5748 (N_5748,N_5539,N_5495);
or U5749 (N_5749,N_5537,N_5520);
nand U5750 (N_5750,N_5505,N_5477);
xor U5751 (N_5751,N_5499,N_5473);
or U5752 (N_5752,N_5599,N_5538);
or U5753 (N_5753,N_5541,N_5412);
and U5754 (N_5754,N_5415,N_5433);
and U5755 (N_5755,N_5538,N_5528);
nand U5756 (N_5756,N_5409,N_5596);
nand U5757 (N_5757,N_5551,N_5506);
xor U5758 (N_5758,N_5403,N_5480);
xor U5759 (N_5759,N_5522,N_5518);
xnor U5760 (N_5760,N_5422,N_5574);
nand U5761 (N_5761,N_5523,N_5503);
nor U5762 (N_5762,N_5494,N_5511);
xor U5763 (N_5763,N_5551,N_5406);
nor U5764 (N_5764,N_5540,N_5492);
or U5765 (N_5765,N_5456,N_5458);
or U5766 (N_5766,N_5578,N_5433);
or U5767 (N_5767,N_5477,N_5441);
nand U5768 (N_5768,N_5481,N_5545);
and U5769 (N_5769,N_5462,N_5575);
or U5770 (N_5770,N_5505,N_5402);
xnor U5771 (N_5771,N_5449,N_5478);
nor U5772 (N_5772,N_5553,N_5455);
nor U5773 (N_5773,N_5436,N_5489);
and U5774 (N_5774,N_5442,N_5538);
and U5775 (N_5775,N_5526,N_5557);
and U5776 (N_5776,N_5433,N_5499);
or U5777 (N_5777,N_5465,N_5478);
nand U5778 (N_5778,N_5470,N_5583);
xor U5779 (N_5779,N_5522,N_5543);
or U5780 (N_5780,N_5457,N_5590);
xor U5781 (N_5781,N_5582,N_5590);
and U5782 (N_5782,N_5417,N_5442);
and U5783 (N_5783,N_5421,N_5466);
and U5784 (N_5784,N_5531,N_5566);
or U5785 (N_5785,N_5460,N_5598);
xor U5786 (N_5786,N_5471,N_5455);
nor U5787 (N_5787,N_5578,N_5425);
nand U5788 (N_5788,N_5420,N_5417);
or U5789 (N_5789,N_5495,N_5433);
and U5790 (N_5790,N_5422,N_5499);
nor U5791 (N_5791,N_5444,N_5422);
xnor U5792 (N_5792,N_5411,N_5475);
or U5793 (N_5793,N_5516,N_5530);
or U5794 (N_5794,N_5545,N_5422);
and U5795 (N_5795,N_5546,N_5580);
and U5796 (N_5796,N_5532,N_5550);
or U5797 (N_5797,N_5507,N_5439);
or U5798 (N_5798,N_5544,N_5489);
nor U5799 (N_5799,N_5416,N_5492);
or U5800 (N_5800,N_5755,N_5647);
nand U5801 (N_5801,N_5698,N_5736);
and U5802 (N_5802,N_5652,N_5786);
nand U5803 (N_5803,N_5721,N_5615);
nand U5804 (N_5804,N_5747,N_5669);
nor U5805 (N_5805,N_5785,N_5728);
or U5806 (N_5806,N_5600,N_5796);
xor U5807 (N_5807,N_5770,N_5625);
nand U5808 (N_5808,N_5663,N_5725);
nand U5809 (N_5809,N_5654,N_5776);
nand U5810 (N_5810,N_5639,N_5616);
nor U5811 (N_5811,N_5677,N_5749);
nor U5812 (N_5812,N_5607,N_5689);
nor U5813 (N_5813,N_5788,N_5738);
or U5814 (N_5814,N_5781,N_5762);
nor U5815 (N_5815,N_5711,N_5603);
nor U5816 (N_5816,N_5700,N_5727);
nand U5817 (N_5817,N_5658,N_5779);
nand U5818 (N_5818,N_5667,N_5623);
nor U5819 (N_5819,N_5719,N_5619);
xor U5820 (N_5820,N_5628,N_5685);
xnor U5821 (N_5821,N_5799,N_5774);
xor U5822 (N_5822,N_5634,N_5673);
nand U5823 (N_5823,N_5754,N_5742);
or U5824 (N_5824,N_5735,N_5641);
and U5825 (N_5825,N_5768,N_5712);
nor U5826 (N_5826,N_5691,N_5644);
or U5827 (N_5827,N_5761,N_5789);
xnor U5828 (N_5828,N_5764,N_5601);
or U5829 (N_5829,N_5696,N_5683);
nand U5830 (N_5830,N_5772,N_5737);
nand U5831 (N_5831,N_5649,N_5626);
or U5832 (N_5832,N_5688,N_5678);
xnor U5833 (N_5833,N_5775,N_5686);
or U5834 (N_5834,N_5769,N_5760);
xnor U5835 (N_5835,N_5617,N_5707);
or U5836 (N_5836,N_5795,N_5782);
nand U5837 (N_5837,N_5612,N_5726);
nor U5838 (N_5838,N_5733,N_5692);
and U5839 (N_5839,N_5713,N_5618);
nor U5840 (N_5840,N_5757,N_5620);
nor U5841 (N_5841,N_5773,N_5608);
or U5842 (N_5842,N_5629,N_5609);
xor U5843 (N_5843,N_5723,N_5767);
nor U5844 (N_5844,N_5633,N_5675);
nor U5845 (N_5845,N_5701,N_5604);
or U5846 (N_5846,N_5690,N_5792);
and U5847 (N_5847,N_5797,N_5714);
and U5848 (N_5848,N_5636,N_5602);
or U5849 (N_5849,N_5661,N_5752);
xor U5850 (N_5850,N_5610,N_5766);
nand U5851 (N_5851,N_5794,N_5680);
or U5852 (N_5852,N_5687,N_5648);
and U5853 (N_5853,N_5671,N_5672);
nor U5854 (N_5854,N_5638,N_5718);
nand U5855 (N_5855,N_5717,N_5756);
or U5856 (N_5856,N_5695,N_5732);
or U5857 (N_5857,N_5750,N_5708);
nand U5858 (N_5858,N_5622,N_5694);
xor U5859 (N_5859,N_5741,N_5758);
nor U5860 (N_5860,N_5621,N_5702);
nand U5861 (N_5861,N_5759,N_5783);
and U5862 (N_5862,N_5668,N_5630);
xnor U5863 (N_5863,N_5651,N_5715);
or U5864 (N_5864,N_5645,N_5640);
or U5865 (N_5865,N_5657,N_5676);
xor U5866 (N_5866,N_5653,N_5753);
or U5867 (N_5867,N_5611,N_5787);
and U5868 (N_5868,N_5720,N_5642);
and U5869 (N_5869,N_5693,N_5664);
and U5870 (N_5870,N_5703,N_5646);
or U5871 (N_5871,N_5709,N_5679);
and U5872 (N_5872,N_5793,N_5632);
and U5873 (N_5873,N_5697,N_5659);
nor U5874 (N_5874,N_5660,N_5729);
nand U5875 (N_5875,N_5627,N_5635);
and U5876 (N_5876,N_5684,N_5790);
nor U5877 (N_5877,N_5746,N_5656);
and U5878 (N_5878,N_5665,N_5699);
or U5879 (N_5879,N_5724,N_5722);
xnor U5880 (N_5880,N_5631,N_5798);
and U5881 (N_5881,N_5780,N_5734);
xor U5882 (N_5882,N_5710,N_5730);
nand U5883 (N_5883,N_5748,N_5771);
nand U5884 (N_5884,N_5655,N_5740);
and U5885 (N_5885,N_5682,N_5745);
nand U5886 (N_5886,N_5706,N_5643);
xnor U5887 (N_5887,N_5784,N_5739);
xnor U5888 (N_5888,N_5777,N_5791);
nor U5889 (N_5889,N_5778,N_5666);
nand U5890 (N_5890,N_5731,N_5705);
nand U5891 (N_5891,N_5662,N_5606);
and U5892 (N_5892,N_5613,N_5763);
or U5893 (N_5893,N_5614,N_5765);
and U5894 (N_5894,N_5751,N_5650);
and U5895 (N_5895,N_5605,N_5716);
or U5896 (N_5896,N_5637,N_5744);
and U5897 (N_5897,N_5743,N_5704);
nand U5898 (N_5898,N_5674,N_5681);
nor U5899 (N_5899,N_5624,N_5670);
xor U5900 (N_5900,N_5650,N_5720);
and U5901 (N_5901,N_5640,N_5675);
xnor U5902 (N_5902,N_5602,N_5772);
nor U5903 (N_5903,N_5686,N_5625);
nor U5904 (N_5904,N_5739,N_5608);
and U5905 (N_5905,N_5718,N_5783);
or U5906 (N_5906,N_5622,N_5759);
or U5907 (N_5907,N_5770,N_5731);
xnor U5908 (N_5908,N_5650,N_5603);
and U5909 (N_5909,N_5755,N_5697);
nand U5910 (N_5910,N_5658,N_5624);
or U5911 (N_5911,N_5778,N_5689);
xor U5912 (N_5912,N_5708,N_5612);
xor U5913 (N_5913,N_5684,N_5779);
or U5914 (N_5914,N_5632,N_5679);
xor U5915 (N_5915,N_5664,N_5635);
and U5916 (N_5916,N_5710,N_5691);
nor U5917 (N_5917,N_5646,N_5702);
xnor U5918 (N_5918,N_5631,N_5611);
and U5919 (N_5919,N_5685,N_5799);
nand U5920 (N_5920,N_5741,N_5777);
xor U5921 (N_5921,N_5610,N_5747);
or U5922 (N_5922,N_5626,N_5771);
and U5923 (N_5923,N_5786,N_5629);
nor U5924 (N_5924,N_5787,N_5669);
and U5925 (N_5925,N_5620,N_5790);
and U5926 (N_5926,N_5795,N_5640);
xor U5927 (N_5927,N_5703,N_5769);
xnor U5928 (N_5928,N_5779,N_5623);
and U5929 (N_5929,N_5607,N_5700);
nand U5930 (N_5930,N_5618,N_5660);
nand U5931 (N_5931,N_5693,N_5745);
or U5932 (N_5932,N_5750,N_5658);
or U5933 (N_5933,N_5685,N_5689);
and U5934 (N_5934,N_5790,N_5625);
nand U5935 (N_5935,N_5758,N_5786);
and U5936 (N_5936,N_5682,N_5798);
nand U5937 (N_5937,N_5613,N_5731);
and U5938 (N_5938,N_5690,N_5619);
and U5939 (N_5939,N_5622,N_5745);
nand U5940 (N_5940,N_5615,N_5641);
xnor U5941 (N_5941,N_5663,N_5696);
nor U5942 (N_5942,N_5602,N_5635);
xnor U5943 (N_5943,N_5719,N_5657);
nand U5944 (N_5944,N_5617,N_5630);
nor U5945 (N_5945,N_5726,N_5712);
or U5946 (N_5946,N_5707,N_5628);
and U5947 (N_5947,N_5724,N_5714);
and U5948 (N_5948,N_5721,N_5650);
or U5949 (N_5949,N_5627,N_5618);
and U5950 (N_5950,N_5659,N_5775);
and U5951 (N_5951,N_5752,N_5792);
nor U5952 (N_5952,N_5602,N_5703);
nor U5953 (N_5953,N_5767,N_5657);
xor U5954 (N_5954,N_5709,N_5767);
nand U5955 (N_5955,N_5706,N_5720);
and U5956 (N_5956,N_5634,N_5741);
or U5957 (N_5957,N_5643,N_5725);
or U5958 (N_5958,N_5668,N_5798);
nor U5959 (N_5959,N_5704,N_5602);
or U5960 (N_5960,N_5761,N_5640);
or U5961 (N_5961,N_5755,N_5796);
or U5962 (N_5962,N_5671,N_5782);
and U5963 (N_5963,N_5739,N_5793);
and U5964 (N_5964,N_5742,N_5671);
nor U5965 (N_5965,N_5751,N_5601);
nand U5966 (N_5966,N_5692,N_5741);
nand U5967 (N_5967,N_5687,N_5773);
nor U5968 (N_5968,N_5658,N_5722);
xor U5969 (N_5969,N_5775,N_5754);
or U5970 (N_5970,N_5641,N_5629);
nand U5971 (N_5971,N_5701,N_5776);
nand U5972 (N_5972,N_5759,N_5699);
nand U5973 (N_5973,N_5745,N_5776);
nand U5974 (N_5974,N_5720,N_5673);
xnor U5975 (N_5975,N_5637,N_5799);
or U5976 (N_5976,N_5713,N_5624);
and U5977 (N_5977,N_5602,N_5765);
or U5978 (N_5978,N_5686,N_5638);
or U5979 (N_5979,N_5782,N_5734);
or U5980 (N_5980,N_5685,N_5690);
and U5981 (N_5981,N_5634,N_5768);
or U5982 (N_5982,N_5625,N_5601);
or U5983 (N_5983,N_5643,N_5679);
xnor U5984 (N_5984,N_5719,N_5752);
and U5985 (N_5985,N_5745,N_5603);
nor U5986 (N_5986,N_5764,N_5744);
or U5987 (N_5987,N_5780,N_5698);
and U5988 (N_5988,N_5730,N_5764);
or U5989 (N_5989,N_5675,N_5758);
or U5990 (N_5990,N_5646,N_5734);
and U5991 (N_5991,N_5718,N_5609);
or U5992 (N_5992,N_5685,N_5674);
xnor U5993 (N_5993,N_5721,N_5670);
xor U5994 (N_5994,N_5660,N_5720);
xnor U5995 (N_5995,N_5661,N_5784);
xnor U5996 (N_5996,N_5688,N_5733);
and U5997 (N_5997,N_5651,N_5654);
and U5998 (N_5998,N_5765,N_5600);
xnor U5999 (N_5999,N_5775,N_5663);
nand U6000 (N_6000,N_5940,N_5831);
or U6001 (N_6001,N_5923,N_5873);
and U6002 (N_6002,N_5861,N_5841);
and U6003 (N_6003,N_5890,N_5889);
nand U6004 (N_6004,N_5826,N_5941);
or U6005 (N_6005,N_5833,N_5827);
nand U6006 (N_6006,N_5848,N_5982);
xor U6007 (N_6007,N_5807,N_5886);
or U6008 (N_6008,N_5955,N_5954);
and U6009 (N_6009,N_5881,N_5916);
xnor U6010 (N_6010,N_5930,N_5913);
xor U6011 (N_6011,N_5963,N_5868);
or U6012 (N_6012,N_5846,N_5839);
and U6013 (N_6013,N_5938,N_5858);
and U6014 (N_6014,N_5877,N_5864);
nand U6015 (N_6015,N_5885,N_5989);
and U6016 (N_6016,N_5897,N_5866);
and U6017 (N_6017,N_5957,N_5962);
nor U6018 (N_6018,N_5906,N_5842);
nand U6019 (N_6019,N_5949,N_5970);
or U6020 (N_6020,N_5870,N_5813);
and U6021 (N_6021,N_5820,N_5818);
nor U6022 (N_6022,N_5922,N_5974);
nand U6023 (N_6023,N_5952,N_5950);
and U6024 (N_6024,N_5956,N_5884);
or U6025 (N_6025,N_5903,N_5828);
nand U6026 (N_6026,N_5810,N_5898);
xor U6027 (N_6027,N_5953,N_5997);
xnor U6028 (N_6028,N_5915,N_5939);
nor U6029 (N_6029,N_5928,N_5863);
nand U6030 (N_6030,N_5800,N_5910);
xnor U6031 (N_6031,N_5925,N_5821);
nor U6032 (N_6032,N_5838,N_5936);
nand U6033 (N_6033,N_5811,N_5985);
and U6034 (N_6034,N_5917,N_5944);
xor U6035 (N_6035,N_5914,N_5934);
nor U6036 (N_6036,N_5933,N_5951);
or U6037 (N_6037,N_5869,N_5892);
and U6038 (N_6038,N_5887,N_5837);
xor U6039 (N_6039,N_5961,N_5968);
or U6040 (N_6040,N_5865,N_5999);
nor U6041 (N_6041,N_5882,N_5978);
or U6042 (N_6042,N_5876,N_5867);
and U6043 (N_6043,N_5819,N_5994);
nand U6044 (N_6044,N_5871,N_5981);
nor U6045 (N_6045,N_5891,N_5883);
and U6046 (N_6046,N_5998,N_5980);
xnor U6047 (N_6047,N_5942,N_5849);
nor U6048 (N_6048,N_5995,N_5878);
nor U6049 (N_6049,N_5836,N_5824);
xor U6050 (N_6050,N_5992,N_5948);
or U6051 (N_6051,N_5904,N_5975);
nor U6052 (N_6052,N_5815,N_5895);
or U6053 (N_6053,N_5894,N_5801);
xor U6054 (N_6054,N_5817,N_5911);
nand U6055 (N_6055,N_5830,N_5862);
xnor U6056 (N_6056,N_5937,N_5859);
nor U6057 (N_6057,N_5943,N_5996);
or U6058 (N_6058,N_5814,N_5805);
xor U6059 (N_6059,N_5947,N_5816);
nand U6060 (N_6060,N_5973,N_5977);
nor U6061 (N_6061,N_5823,N_5960);
xor U6062 (N_6062,N_5919,N_5929);
nor U6063 (N_6063,N_5843,N_5986);
and U6064 (N_6064,N_5804,N_5927);
xor U6065 (N_6065,N_5875,N_5988);
nor U6066 (N_6066,N_5912,N_5851);
or U6067 (N_6067,N_5893,N_5924);
nand U6068 (N_6068,N_5932,N_5931);
or U6069 (N_6069,N_5976,N_5806);
and U6070 (N_6070,N_5965,N_5822);
and U6071 (N_6071,N_5845,N_5874);
nor U6072 (N_6072,N_5901,N_5969);
or U6073 (N_6073,N_5850,N_5879);
xor U6074 (N_6074,N_5921,N_5802);
nor U6075 (N_6075,N_5918,N_5993);
and U6076 (N_6076,N_5909,N_5971);
and U6077 (N_6077,N_5959,N_5856);
or U6078 (N_6078,N_5987,N_5900);
xnor U6079 (N_6079,N_5854,N_5809);
and U6080 (N_6080,N_5902,N_5803);
nor U6081 (N_6081,N_5966,N_5972);
and U6082 (N_6082,N_5896,N_5853);
or U6083 (N_6083,N_5872,N_5899);
and U6084 (N_6084,N_5920,N_5825);
or U6085 (N_6085,N_5964,N_5983);
nand U6086 (N_6086,N_5967,N_5908);
nor U6087 (N_6087,N_5812,N_5880);
nor U6088 (N_6088,N_5888,N_5834);
nor U6089 (N_6089,N_5829,N_5946);
and U6090 (N_6090,N_5860,N_5840);
xnor U6091 (N_6091,N_5855,N_5852);
nand U6092 (N_6092,N_5905,N_5991);
nand U6093 (N_6093,N_5926,N_5945);
and U6094 (N_6094,N_5979,N_5857);
nor U6095 (N_6095,N_5935,N_5907);
nand U6096 (N_6096,N_5847,N_5832);
nor U6097 (N_6097,N_5835,N_5808);
or U6098 (N_6098,N_5958,N_5984);
xnor U6099 (N_6099,N_5844,N_5990);
or U6100 (N_6100,N_5937,N_5967);
xnor U6101 (N_6101,N_5811,N_5880);
xnor U6102 (N_6102,N_5923,N_5808);
and U6103 (N_6103,N_5990,N_5951);
and U6104 (N_6104,N_5919,N_5831);
or U6105 (N_6105,N_5954,N_5830);
and U6106 (N_6106,N_5910,N_5994);
nor U6107 (N_6107,N_5948,N_5966);
nand U6108 (N_6108,N_5982,N_5888);
xor U6109 (N_6109,N_5928,N_5976);
or U6110 (N_6110,N_5988,N_5826);
nor U6111 (N_6111,N_5940,N_5946);
or U6112 (N_6112,N_5934,N_5945);
or U6113 (N_6113,N_5805,N_5972);
and U6114 (N_6114,N_5840,N_5841);
nand U6115 (N_6115,N_5988,N_5923);
and U6116 (N_6116,N_5963,N_5874);
or U6117 (N_6117,N_5911,N_5805);
or U6118 (N_6118,N_5938,N_5842);
nand U6119 (N_6119,N_5981,N_5867);
nor U6120 (N_6120,N_5927,N_5954);
nand U6121 (N_6121,N_5866,N_5985);
or U6122 (N_6122,N_5836,N_5817);
nand U6123 (N_6123,N_5879,N_5978);
or U6124 (N_6124,N_5870,N_5800);
nor U6125 (N_6125,N_5932,N_5897);
or U6126 (N_6126,N_5924,N_5937);
and U6127 (N_6127,N_5909,N_5951);
or U6128 (N_6128,N_5894,N_5958);
and U6129 (N_6129,N_5856,N_5918);
nand U6130 (N_6130,N_5934,N_5801);
nor U6131 (N_6131,N_5936,N_5836);
nor U6132 (N_6132,N_5854,N_5936);
and U6133 (N_6133,N_5837,N_5957);
or U6134 (N_6134,N_5847,N_5823);
nand U6135 (N_6135,N_5917,N_5968);
nor U6136 (N_6136,N_5937,N_5977);
or U6137 (N_6137,N_5863,N_5851);
or U6138 (N_6138,N_5974,N_5829);
or U6139 (N_6139,N_5847,N_5900);
nor U6140 (N_6140,N_5827,N_5870);
or U6141 (N_6141,N_5901,N_5900);
nand U6142 (N_6142,N_5808,N_5841);
xor U6143 (N_6143,N_5867,N_5908);
nand U6144 (N_6144,N_5882,N_5814);
nand U6145 (N_6145,N_5899,N_5995);
or U6146 (N_6146,N_5936,N_5970);
xor U6147 (N_6147,N_5822,N_5801);
xnor U6148 (N_6148,N_5871,N_5913);
xnor U6149 (N_6149,N_5875,N_5914);
or U6150 (N_6150,N_5860,N_5938);
and U6151 (N_6151,N_5869,N_5956);
xor U6152 (N_6152,N_5936,N_5943);
nand U6153 (N_6153,N_5971,N_5858);
or U6154 (N_6154,N_5918,N_5998);
or U6155 (N_6155,N_5810,N_5822);
nand U6156 (N_6156,N_5921,N_5881);
xnor U6157 (N_6157,N_5857,N_5923);
xor U6158 (N_6158,N_5800,N_5979);
and U6159 (N_6159,N_5973,N_5972);
and U6160 (N_6160,N_5878,N_5812);
or U6161 (N_6161,N_5880,N_5959);
and U6162 (N_6162,N_5867,N_5849);
or U6163 (N_6163,N_5811,N_5834);
nor U6164 (N_6164,N_5985,N_5803);
nand U6165 (N_6165,N_5836,N_5955);
nor U6166 (N_6166,N_5805,N_5962);
nand U6167 (N_6167,N_5925,N_5808);
and U6168 (N_6168,N_5890,N_5960);
nor U6169 (N_6169,N_5887,N_5919);
xor U6170 (N_6170,N_5921,N_5854);
or U6171 (N_6171,N_5810,N_5983);
nand U6172 (N_6172,N_5982,N_5850);
xnor U6173 (N_6173,N_5812,N_5807);
or U6174 (N_6174,N_5889,N_5923);
or U6175 (N_6175,N_5878,N_5828);
and U6176 (N_6176,N_5944,N_5998);
xor U6177 (N_6177,N_5999,N_5866);
or U6178 (N_6178,N_5959,N_5987);
or U6179 (N_6179,N_5920,N_5950);
nor U6180 (N_6180,N_5913,N_5885);
or U6181 (N_6181,N_5816,N_5828);
xor U6182 (N_6182,N_5817,N_5969);
or U6183 (N_6183,N_5906,N_5805);
nand U6184 (N_6184,N_5819,N_5948);
nand U6185 (N_6185,N_5906,N_5858);
xnor U6186 (N_6186,N_5852,N_5848);
xnor U6187 (N_6187,N_5847,N_5805);
nand U6188 (N_6188,N_5879,N_5940);
nand U6189 (N_6189,N_5893,N_5968);
nand U6190 (N_6190,N_5999,N_5935);
nor U6191 (N_6191,N_5840,N_5888);
xnor U6192 (N_6192,N_5940,N_5884);
nand U6193 (N_6193,N_5807,N_5800);
and U6194 (N_6194,N_5896,N_5982);
nand U6195 (N_6195,N_5943,N_5864);
or U6196 (N_6196,N_5940,N_5804);
nor U6197 (N_6197,N_5823,N_5941);
or U6198 (N_6198,N_5957,N_5806);
nand U6199 (N_6199,N_5910,N_5816);
nand U6200 (N_6200,N_6101,N_6086);
nand U6201 (N_6201,N_6131,N_6051);
nor U6202 (N_6202,N_6088,N_6164);
xnor U6203 (N_6203,N_6083,N_6180);
xor U6204 (N_6204,N_6074,N_6040);
nand U6205 (N_6205,N_6011,N_6053);
nand U6206 (N_6206,N_6105,N_6046);
nor U6207 (N_6207,N_6031,N_6048);
nor U6208 (N_6208,N_6027,N_6050);
nand U6209 (N_6209,N_6084,N_6006);
nor U6210 (N_6210,N_6094,N_6103);
nand U6211 (N_6211,N_6179,N_6177);
nor U6212 (N_6212,N_6190,N_6115);
nor U6213 (N_6213,N_6157,N_6073);
or U6214 (N_6214,N_6199,N_6166);
and U6215 (N_6215,N_6021,N_6151);
and U6216 (N_6216,N_6186,N_6137);
nand U6217 (N_6217,N_6121,N_6041);
or U6218 (N_6218,N_6039,N_6120);
and U6219 (N_6219,N_6155,N_6150);
nor U6220 (N_6220,N_6197,N_6020);
and U6221 (N_6221,N_6173,N_6100);
and U6222 (N_6222,N_6152,N_6052);
and U6223 (N_6223,N_6172,N_6033);
xnor U6224 (N_6224,N_6154,N_6175);
or U6225 (N_6225,N_6176,N_6030);
nand U6226 (N_6226,N_6135,N_6159);
xnor U6227 (N_6227,N_6167,N_6072);
xor U6228 (N_6228,N_6097,N_6168);
nor U6229 (N_6229,N_6098,N_6127);
or U6230 (N_6230,N_6018,N_6194);
nand U6231 (N_6231,N_6079,N_6107);
or U6232 (N_6232,N_6080,N_6085);
nand U6233 (N_6233,N_6010,N_6095);
xor U6234 (N_6234,N_6140,N_6026);
xnor U6235 (N_6235,N_6111,N_6129);
nand U6236 (N_6236,N_6136,N_6062);
xor U6237 (N_6237,N_6161,N_6065);
or U6238 (N_6238,N_6185,N_6170);
or U6239 (N_6239,N_6071,N_6189);
nand U6240 (N_6240,N_6087,N_6195);
nand U6241 (N_6241,N_6004,N_6032);
nor U6242 (N_6242,N_6017,N_6188);
xnor U6243 (N_6243,N_6122,N_6109);
nand U6244 (N_6244,N_6163,N_6013);
and U6245 (N_6245,N_6093,N_6171);
nor U6246 (N_6246,N_6169,N_6058);
xor U6247 (N_6247,N_6144,N_6019);
nor U6248 (N_6248,N_6196,N_6090);
xnor U6249 (N_6249,N_6132,N_6067);
and U6250 (N_6250,N_6110,N_6156);
and U6251 (N_6251,N_6028,N_6012);
nand U6252 (N_6252,N_6038,N_6042);
nor U6253 (N_6253,N_6192,N_6008);
or U6254 (N_6254,N_6125,N_6060);
xnor U6255 (N_6255,N_6056,N_6148);
and U6256 (N_6256,N_6108,N_6066);
nor U6257 (N_6257,N_6162,N_6145);
and U6258 (N_6258,N_6191,N_6149);
nor U6259 (N_6259,N_6112,N_6153);
or U6260 (N_6260,N_6089,N_6118);
xor U6261 (N_6261,N_6104,N_6141);
or U6262 (N_6262,N_6000,N_6139);
nand U6263 (N_6263,N_6146,N_6055);
and U6264 (N_6264,N_6114,N_6025);
nor U6265 (N_6265,N_6193,N_6138);
nand U6266 (N_6266,N_6142,N_6143);
xnor U6267 (N_6267,N_6002,N_6081);
nor U6268 (N_6268,N_6061,N_6054);
xnor U6269 (N_6269,N_6178,N_6045);
nor U6270 (N_6270,N_6096,N_6016);
nand U6271 (N_6271,N_6198,N_6047);
nor U6272 (N_6272,N_6005,N_6126);
and U6273 (N_6273,N_6082,N_6187);
xnor U6274 (N_6274,N_6099,N_6124);
xor U6275 (N_6275,N_6119,N_6102);
nand U6276 (N_6276,N_6069,N_6147);
and U6277 (N_6277,N_6078,N_6014);
xnor U6278 (N_6278,N_6076,N_6117);
or U6279 (N_6279,N_6024,N_6009);
xnor U6280 (N_6280,N_6022,N_6075);
nand U6281 (N_6281,N_6184,N_6044);
xor U6282 (N_6282,N_6091,N_6023);
and U6283 (N_6283,N_6128,N_6160);
nor U6284 (N_6284,N_6029,N_6036);
nand U6285 (N_6285,N_6001,N_6130);
xor U6286 (N_6286,N_6106,N_6049);
xor U6287 (N_6287,N_6034,N_6113);
nor U6288 (N_6288,N_6174,N_6077);
nor U6289 (N_6289,N_6182,N_6059);
nor U6290 (N_6290,N_6123,N_6133);
xor U6291 (N_6291,N_6181,N_6134);
and U6292 (N_6292,N_6092,N_6165);
xor U6293 (N_6293,N_6064,N_6043);
and U6294 (N_6294,N_6007,N_6057);
xor U6295 (N_6295,N_6158,N_6070);
or U6296 (N_6296,N_6068,N_6063);
or U6297 (N_6297,N_6037,N_6003);
nor U6298 (N_6298,N_6015,N_6116);
or U6299 (N_6299,N_6035,N_6183);
nand U6300 (N_6300,N_6103,N_6042);
xnor U6301 (N_6301,N_6133,N_6189);
nor U6302 (N_6302,N_6196,N_6184);
or U6303 (N_6303,N_6052,N_6134);
xor U6304 (N_6304,N_6035,N_6003);
nand U6305 (N_6305,N_6140,N_6073);
xor U6306 (N_6306,N_6001,N_6038);
xnor U6307 (N_6307,N_6113,N_6015);
and U6308 (N_6308,N_6128,N_6136);
nand U6309 (N_6309,N_6198,N_6093);
nand U6310 (N_6310,N_6175,N_6166);
xnor U6311 (N_6311,N_6000,N_6190);
nand U6312 (N_6312,N_6028,N_6177);
nand U6313 (N_6313,N_6043,N_6146);
nor U6314 (N_6314,N_6081,N_6011);
nand U6315 (N_6315,N_6041,N_6192);
nand U6316 (N_6316,N_6102,N_6027);
nand U6317 (N_6317,N_6061,N_6119);
xnor U6318 (N_6318,N_6042,N_6174);
xor U6319 (N_6319,N_6097,N_6044);
or U6320 (N_6320,N_6012,N_6153);
xnor U6321 (N_6321,N_6177,N_6057);
nand U6322 (N_6322,N_6086,N_6051);
nand U6323 (N_6323,N_6054,N_6105);
and U6324 (N_6324,N_6054,N_6149);
and U6325 (N_6325,N_6052,N_6026);
xnor U6326 (N_6326,N_6092,N_6041);
and U6327 (N_6327,N_6113,N_6195);
and U6328 (N_6328,N_6075,N_6073);
and U6329 (N_6329,N_6115,N_6165);
nand U6330 (N_6330,N_6123,N_6038);
nand U6331 (N_6331,N_6007,N_6126);
or U6332 (N_6332,N_6178,N_6017);
or U6333 (N_6333,N_6028,N_6159);
xor U6334 (N_6334,N_6112,N_6058);
nor U6335 (N_6335,N_6049,N_6055);
nor U6336 (N_6336,N_6025,N_6088);
and U6337 (N_6337,N_6067,N_6138);
and U6338 (N_6338,N_6164,N_6002);
nor U6339 (N_6339,N_6164,N_6101);
nand U6340 (N_6340,N_6074,N_6037);
and U6341 (N_6341,N_6059,N_6095);
and U6342 (N_6342,N_6036,N_6198);
nand U6343 (N_6343,N_6144,N_6154);
nand U6344 (N_6344,N_6024,N_6172);
and U6345 (N_6345,N_6080,N_6188);
nor U6346 (N_6346,N_6000,N_6101);
nand U6347 (N_6347,N_6030,N_6167);
nor U6348 (N_6348,N_6094,N_6161);
xnor U6349 (N_6349,N_6113,N_6086);
and U6350 (N_6350,N_6117,N_6188);
xor U6351 (N_6351,N_6115,N_6035);
nor U6352 (N_6352,N_6196,N_6070);
xor U6353 (N_6353,N_6021,N_6067);
xor U6354 (N_6354,N_6189,N_6193);
xnor U6355 (N_6355,N_6003,N_6145);
nand U6356 (N_6356,N_6048,N_6055);
nor U6357 (N_6357,N_6174,N_6059);
and U6358 (N_6358,N_6031,N_6177);
or U6359 (N_6359,N_6153,N_6059);
xnor U6360 (N_6360,N_6186,N_6170);
nand U6361 (N_6361,N_6102,N_6167);
xor U6362 (N_6362,N_6032,N_6086);
xnor U6363 (N_6363,N_6047,N_6131);
or U6364 (N_6364,N_6126,N_6045);
xor U6365 (N_6365,N_6051,N_6111);
or U6366 (N_6366,N_6135,N_6150);
nand U6367 (N_6367,N_6138,N_6068);
or U6368 (N_6368,N_6182,N_6137);
and U6369 (N_6369,N_6148,N_6064);
nor U6370 (N_6370,N_6060,N_6015);
nand U6371 (N_6371,N_6177,N_6111);
or U6372 (N_6372,N_6119,N_6087);
nor U6373 (N_6373,N_6015,N_6025);
nand U6374 (N_6374,N_6073,N_6171);
and U6375 (N_6375,N_6165,N_6014);
xnor U6376 (N_6376,N_6199,N_6159);
and U6377 (N_6377,N_6082,N_6036);
nand U6378 (N_6378,N_6089,N_6093);
nor U6379 (N_6379,N_6036,N_6054);
nor U6380 (N_6380,N_6063,N_6142);
nor U6381 (N_6381,N_6074,N_6189);
xnor U6382 (N_6382,N_6139,N_6046);
or U6383 (N_6383,N_6047,N_6033);
xnor U6384 (N_6384,N_6053,N_6120);
and U6385 (N_6385,N_6019,N_6015);
or U6386 (N_6386,N_6064,N_6058);
and U6387 (N_6387,N_6149,N_6129);
nand U6388 (N_6388,N_6011,N_6045);
nand U6389 (N_6389,N_6197,N_6158);
nand U6390 (N_6390,N_6029,N_6102);
or U6391 (N_6391,N_6117,N_6194);
xor U6392 (N_6392,N_6154,N_6167);
or U6393 (N_6393,N_6126,N_6070);
or U6394 (N_6394,N_6197,N_6025);
and U6395 (N_6395,N_6054,N_6156);
nand U6396 (N_6396,N_6007,N_6027);
nor U6397 (N_6397,N_6056,N_6037);
xor U6398 (N_6398,N_6076,N_6069);
and U6399 (N_6399,N_6188,N_6094);
or U6400 (N_6400,N_6269,N_6230);
nor U6401 (N_6401,N_6262,N_6291);
nand U6402 (N_6402,N_6326,N_6212);
nor U6403 (N_6403,N_6229,N_6286);
or U6404 (N_6404,N_6203,N_6379);
or U6405 (N_6405,N_6318,N_6317);
nor U6406 (N_6406,N_6320,N_6348);
nand U6407 (N_6407,N_6282,N_6314);
or U6408 (N_6408,N_6332,N_6310);
nor U6409 (N_6409,N_6372,N_6353);
nand U6410 (N_6410,N_6341,N_6359);
nand U6411 (N_6411,N_6213,N_6329);
xnor U6412 (N_6412,N_6245,N_6254);
nor U6413 (N_6413,N_6392,N_6304);
nand U6414 (N_6414,N_6395,N_6370);
or U6415 (N_6415,N_6251,N_6390);
and U6416 (N_6416,N_6215,N_6330);
nor U6417 (N_6417,N_6323,N_6228);
xor U6418 (N_6418,N_6233,N_6253);
or U6419 (N_6419,N_6378,N_6319);
xnor U6420 (N_6420,N_6264,N_6327);
and U6421 (N_6421,N_6369,N_6394);
xnor U6422 (N_6422,N_6249,N_6287);
nand U6423 (N_6423,N_6289,N_6345);
nand U6424 (N_6424,N_6205,N_6288);
nor U6425 (N_6425,N_6223,N_6231);
and U6426 (N_6426,N_6204,N_6208);
xor U6427 (N_6427,N_6225,N_6259);
nand U6428 (N_6428,N_6239,N_6306);
and U6429 (N_6429,N_6297,N_6339);
and U6430 (N_6430,N_6383,N_6211);
xor U6431 (N_6431,N_6365,N_6373);
and U6432 (N_6432,N_6386,N_6385);
nor U6433 (N_6433,N_6387,N_6237);
or U6434 (N_6434,N_6350,N_6274);
nand U6435 (N_6435,N_6256,N_6375);
or U6436 (N_6436,N_6242,N_6235);
xnor U6437 (N_6437,N_6250,N_6312);
nor U6438 (N_6438,N_6311,N_6337);
xor U6439 (N_6439,N_6260,N_6305);
nand U6440 (N_6440,N_6263,N_6296);
nor U6441 (N_6441,N_6381,N_6295);
nor U6442 (N_6442,N_6328,N_6361);
and U6443 (N_6443,N_6255,N_6202);
xor U6444 (N_6444,N_6335,N_6331);
nand U6445 (N_6445,N_6380,N_6285);
nand U6446 (N_6446,N_6268,N_6338);
nor U6447 (N_6447,N_6397,N_6360);
nor U6448 (N_6448,N_6303,N_6316);
nor U6449 (N_6449,N_6384,N_6284);
and U6450 (N_6450,N_6398,N_6349);
and U6451 (N_6451,N_6218,N_6207);
and U6452 (N_6452,N_6399,N_6277);
and U6453 (N_6453,N_6283,N_6313);
and U6454 (N_6454,N_6325,N_6364);
xor U6455 (N_6455,N_6273,N_6377);
and U6456 (N_6456,N_6309,N_6240);
nand U6457 (N_6457,N_6324,N_6281);
xor U6458 (N_6458,N_6333,N_6376);
and U6459 (N_6459,N_6391,N_6389);
nor U6460 (N_6460,N_6272,N_6292);
or U6461 (N_6461,N_6347,N_6315);
nor U6462 (N_6462,N_6300,N_6200);
nand U6463 (N_6463,N_6265,N_6271);
or U6464 (N_6464,N_6371,N_6299);
nor U6465 (N_6465,N_6217,N_6206);
xnor U6466 (N_6466,N_6388,N_6201);
nor U6467 (N_6467,N_6368,N_6238);
or U6468 (N_6468,N_6294,N_6227);
and U6469 (N_6469,N_6234,N_6257);
and U6470 (N_6470,N_6221,N_6357);
nand U6471 (N_6471,N_6216,N_6355);
and U6472 (N_6472,N_6210,N_6363);
or U6473 (N_6473,N_6340,N_6366);
xnor U6474 (N_6474,N_6243,N_6367);
nand U6475 (N_6475,N_6301,N_6322);
or U6476 (N_6476,N_6354,N_6278);
and U6477 (N_6477,N_6280,N_6374);
and U6478 (N_6478,N_6334,N_6321);
nor U6479 (N_6479,N_6362,N_6252);
xor U6480 (N_6480,N_6356,N_6222);
xor U6481 (N_6481,N_6307,N_6352);
and U6482 (N_6482,N_6232,N_6258);
and U6483 (N_6483,N_6293,N_6248);
nand U6484 (N_6484,N_6351,N_6346);
and U6485 (N_6485,N_6290,N_6302);
or U6486 (N_6486,N_6214,N_6276);
xnor U6487 (N_6487,N_6358,N_6261);
nor U6488 (N_6488,N_6393,N_6336);
nor U6489 (N_6489,N_6241,N_6220);
xor U6490 (N_6490,N_6209,N_6267);
xnor U6491 (N_6491,N_6396,N_6270);
xor U6492 (N_6492,N_6246,N_6247);
nor U6493 (N_6493,N_6342,N_6244);
or U6494 (N_6494,N_6266,N_6308);
nor U6495 (N_6495,N_6382,N_6343);
nand U6496 (N_6496,N_6226,N_6224);
nor U6497 (N_6497,N_6236,N_6219);
xor U6498 (N_6498,N_6275,N_6298);
or U6499 (N_6499,N_6279,N_6344);
and U6500 (N_6500,N_6312,N_6202);
nand U6501 (N_6501,N_6219,N_6362);
and U6502 (N_6502,N_6386,N_6235);
nor U6503 (N_6503,N_6319,N_6383);
xnor U6504 (N_6504,N_6253,N_6381);
and U6505 (N_6505,N_6310,N_6292);
nand U6506 (N_6506,N_6239,N_6340);
nand U6507 (N_6507,N_6208,N_6380);
and U6508 (N_6508,N_6277,N_6296);
and U6509 (N_6509,N_6281,N_6289);
xor U6510 (N_6510,N_6376,N_6248);
nand U6511 (N_6511,N_6386,N_6275);
xor U6512 (N_6512,N_6332,N_6322);
xor U6513 (N_6513,N_6253,N_6226);
nand U6514 (N_6514,N_6254,N_6368);
or U6515 (N_6515,N_6222,N_6274);
xnor U6516 (N_6516,N_6240,N_6311);
and U6517 (N_6517,N_6328,N_6260);
or U6518 (N_6518,N_6288,N_6323);
nor U6519 (N_6519,N_6399,N_6219);
or U6520 (N_6520,N_6254,N_6352);
xor U6521 (N_6521,N_6246,N_6324);
nor U6522 (N_6522,N_6373,N_6262);
nand U6523 (N_6523,N_6349,N_6272);
xnor U6524 (N_6524,N_6256,N_6371);
or U6525 (N_6525,N_6242,N_6333);
nand U6526 (N_6526,N_6213,N_6231);
or U6527 (N_6527,N_6396,N_6373);
nand U6528 (N_6528,N_6352,N_6396);
xor U6529 (N_6529,N_6293,N_6331);
and U6530 (N_6530,N_6284,N_6376);
and U6531 (N_6531,N_6207,N_6296);
xnor U6532 (N_6532,N_6369,N_6236);
xnor U6533 (N_6533,N_6240,N_6333);
xor U6534 (N_6534,N_6271,N_6399);
xnor U6535 (N_6535,N_6390,N_6316);
or U6536 (N_6536,N_6296,N_6367);
nand U6537 (N_6537,N_6200,N_6389);
nor U6538 (N_6538,N_6231,N_6338);
xnor U6539 (N_6539,N_6237,N_6267);
and U6540 (N_6540,N_6287,N_6386);
and U6541 (N_6541,N_6295,N_6387);
nand U6542 (N_6542,N_6344,N_6302);
nand U6543 (N_6543,N_6327,N_6345);
and U6544 (N_6544,N_6338,N_6332);
or U6545 (N_6545,N_6333,N_6202);
and U6546 (N_6546,N_6218,N_6209);
nor U6547 (N_6547,N_6286,N_6311);
nor U6548 (N_6548,N_6278,N_6209);
xnor U6549 (N_6549,N_6370,N_6310);
and U6550 (N_6550,N_6371,N_6355);
xor U6551 (N_6551,N_6296,N_6257);
xor U6552 (N_6552,N_6205,N_6342);
xor U6553 (N_6553,N_6352,N_6257);
nor U6554 (N_6554,N_6393,N_6265);
and U6555 (N_6555,N_6289,N_6315);
and U6556 (N_6556,N_6347,N_6382);
or U6557 (N_6557,N_6201,N_6338);
or U6558 (N_6558,N_6360,N_6352);
xor U6559 (N_6559,N_6369,N_6293);
nor U6560 (N_6560,N_6323,N_6329);
nor U6561 (N_6561,N_6332,N_6312);
and U6562 (N_6562,N_6234,N_6232);
xor U6563 (N_6563,N_6305,N_6332);
xor U6564 (N_6564,N_6229,N_6248);
nand U6565 (N_6565,N_6369,N_6336);
nand U6566 (N_6566,N_6263,N_6254);
or U6567 (N_6567,N_6240,N_6296);
xnor U6568 (N_6568,N_6316,N_6315);
nor U6569 (N_6569,N_6245,N_6282);
nor U6570 (N_6570,N_6337,N_6365);
nand U6571 (N_6571,N_6325,N_6370);
nor U6572 (N_6572,N_6258,N_6312);
or U6573 (N_6573,N_6352,N_6377);
and U6574 (N_6574,N_6208,N_6265);
xor U6575 (N_6575,N_6329,N_6337);
and U6576 (N_6576,N_6370,N_6280);
or U6577 (N_6577,N_6303,N_6335);
nor U6578 (N_6578,N_6267,N_6379);
or U6579 (N_6579,N_6218,N_6354);
xor U6580 (N_6580,N_6245,N_6263);
and U6581 (N_6581,N_6395,N_6294);
or U6582 (N_6582,N_6385,N_6217);
nand U6583 (N_6583,N_6291,N_6272);
nand U6584 (N_6584,N_6339,N_6211);
or U6585 (N_6585,N_6382,N_6256);
xnor U6586 (N_6586,N_6360,N_6300);
or U6587 (N_6587,N_6387,N_6290);
or U6588 (N_6588,N_6336,N_6252);
nand U6589 (N_6589,N_6242,N_6296);
nand U6590 (N_6590,N_6379,N_6202);
xor U6591 (N_6591,N_6371,N_6264);
or U6592 (N_6592,N_6213,N_6360);
and U6593 (N_6593,N_6261,N_6380);
xor U6594 (N_6594,N_6373,N_6292);
or U6595 (N_6595,N_6303,N_6313);
nand U6596 (N_6596,N_6285,N_6298);
nor U6597 (N_6597,N_6376,N_6344);
or U6598 (N_6598,N_6373,N_6324);
xnor U6599 (N_6599,N_6290,N_6322);
or U6600 (N_6600,N_6502,N_6586);
and U6601 (N_6601,N_6430,N_6579);
or U6602 (N_6602,N_6420,N_6472);
or U6603 (N_6603,N_6530,N_6415);
or U6604 (N_6604,N_6436,N_6404);
nand U6605 (N_6605,N_6428,N_6573);
nand U6606 (N_6606,N_6401,N_6545);
and U6607 (N_6607,N_6521,N_6570);
or U6608 (N_6608,N_6537,N_6439);
and U6609 (N_6609,N_6477,N_6433);
xor U6610 (N_6610,N_6523,N_6540);
xor U6611 (N_6611,N_6510,N_6552);
nor U6612 (N_6612,N_6548,N_6435);
xnor U6613 (N_6613,N_6441,N_6514);
nor U6614 (N_6614,N_6487,N_6454);
xor U6615 (N_6615,N_6426,N_6598);
nand U6616 (N_6616,N_6453,N_6425);
xor U6617 (N_6617,N_6565,N_6566);
and U6618 (N_6618,N_6543,N_6507);
and U6619 (N_6619,N_6547,N_6538);
and U6620 (N_6620,N_6513,N_6468);
xnor U6621 (N_6621,N_6534,N_6488);
nor U6622 (N_6622,N_6446,N_6496);
or U6623 (N_6623,N_6531,N_6498);
and U6624 (N_6624,N_6527,N_6581);
nor U6625 (N_6625,N_6564,N_6495);
nand U6626 (N_6626,N_6485,N_6449);
or U6627 (N_6627,N_6535,N_6519);
or U6628 (N_6628,N_6549,N_6588);
xnor U6629 (N_6629,N_6451,N_6524);
nor U6630 (N_6630,N_6518,N_6445);
and U6631 (N_6631,N_6448,N_6438);
nor U6632 (N_6632,N_6529,N_6589);
nor U6633 (N_6633,N_6406,N_6422);
nor U6634 (N_6634,N_6458,N_6479);
and U6635 (N_6635,N_6580,N_6517);
or U6636 (N_6636,N_6432,N_6568);
nand U6637 (N_6637,N_6505,N_6596);
xnor U6638 (N_6638,N_6557,N_6442);
xnor U6639 (N_6639,N_6469,N_6533);
and U6640 (N_6640,N_6408,N_6417);
nand U6641 (N_6641,N_6594,N_6405);
nand U6642 (N_6642,N_6489,N_6452);
and U6643 (N_6643,N_6492,N_6554);
and U6644 (N_6644,N_6544,N_6486);
xor U6645 (N_6645,N_6463,N_6437);
nor U6646 (N_6646,N_6569,N_6550);
and U6647 (N_6647,N_6504,N_6567);
or U6648 (N_6648,N_6532,N_6466);
xnor U6649 (N_6649,N_6411,N_6528);
or U6650 (N_6650,N_6546,N_6423);
or U6651 (N_6651,N_6457,N_6525);
nand U6652 (N_6652,N_6440,N_6400);
and U6653 (N_6653,N_6402,N_6511);
xor U6654 (N_6654,N_6475,N_6575);
or U6655 (N_6655,N_6597,N_6459);
nor U6656 (N_6656,N_6585,N_6471);
xor U6657 (N_6657,N_6482,N_6414);
or U6658 (N_6658,N_6424,N_6558);
or U6659 (N_6659,N_6427,N_6590);
xnor U6660 (N_6660,N_6563,N_6499);
and U6661 (N_6661,N_6413,N_6431);
and U6662 (N_6662,N_6464,N_6576);
and U6663 (N_6663,N_6526,N_6478);
or U6664 (N_6664,N_6500,N_6541);
nand U6665 (N_6665,N_6416,N_6520);
and U6666 (N_6666,N_6516,N_6509);
or U6667 (N_6667,N_6562,N_6591);
nor U6668 (N_6668,N_6506,N_6595);
nand U6669 (N_6669,N_6462,N_6467);
nand U6670 (N_6670,N_6419,N_6456);
nand U6671 (N_6671,N_6403,N_6450);
xor U6672 (N_6672,N_6559,N_6560);
nor U6673 (N_6673,N_6539,N_6474);
xnor U6674 (N_6674,N_6536,N_6429);
xor U6675 (N_6675,N_6503,N_6501);
nand U6676 (N_6676,N_6571,N_6551);
or U6677 (N_6677,N_6484,N_6443);
nor U6678 (N_6678,N_6508,N_6542);
nand U6679 (N_6679,N_6483,N_6412);
xnor U6680 (N_6680,N_6512,N_6409);
nand U6681 (N_6681,N_6553,N_6447);
nand U6682 (N_6682,N_6444,N_6583);
xnor U6683 (N_6683,N_6480,N_6582);
nand U6684 (N_6684,N_6407,N_6556);
nor U6685 (N_6685,N_6476,N_6470);
nor U6686 (N_6686,N_6494,N_6578);
xor U6687 (N_6687,N_6497,N_6584);
or U6688 (N_6688,N_6561,N_6491);
xnor U6689 (N_6689,N_6455,N_6574);
xnor U6690 (N_6690,N_6493,N_6555);
or U6691 (N_6691,N_6490,N_6481);
or U6692 (N_6692,N_6572,N_6434);
or U6693 (N_6693,N_6460,N_6599);
or U6694 (N_6694,N_6593,N_6577);
nand U6695 (N_6695,N_6421,N_6461);
and U6696 (N_6696,N_6410,N_6592);
nand U6697 (N_6697,N_6473,N_6587);
and U6698 (N_6698,N_6515,N_6465);
or U6699 (N_6699,N_6418,N_6522);
and U6700 (N_6700,N_6475,N_6425);
xnor U6701 (N_6701,N_6579,N_6445);
xor U6702 (N_6702,N_6522,N_6583);
nor U6703 (N_6703,N_6540,N_6569);
xnor U6704 (N_6704,N_6444,N_6462);
nor U6705 (N_6705,N_6405,N_6597);
and U6706 (N_6706,N_6564,N_6412);
and U6707 (N_6707,N_6590,N_6525);
nor U6708 (N_6708,N_6539,N_6450);
and U6709 (N_6709,N_6501,N_6596);
and U6710 (N_6710,N_6523,N_6407);
or U6711 (N_6711,N_6466,N_6489);
or U6712 (N_6712,N_6405,N_6547);
nor U6713 (N_6713,N_6450,N_6576);
or U6714 (N_6714,N_6468,N_6487);
xnor U6715 (N_6715,N_6463,N_6465);
nand U6716 (N_6716,N_6582,N_6481);
or U6717 (N_6717,N_6554,N_6438);
and U6718 (N_6718,N_6491,N_6437);
nand U6719 (N_6719,N_6418,N_6461);
nor U6720 (N_6720,N_6559,N_6568);
and U6721 (N_6721,N_6488,N_6533);
nor U6722 (N_6722,N_6574,N_6514);
and U6723 (N_6723,N_6482,N_6412);
and U6724 (N_6724,N_6422,N_6476);
xor U6725 (N_6725,N_6570,N_6508);
nor U6726 (N_6726,N_6489,N_6424);
nand U6727 (N_6727,N_6559,N_6499);
nor U6728 (N_6728,N_6469,N_6405);
xnor U6729 (N_6729,N_6472,N_6587);
nor U6730 (N_6730,N_6456,N_6557);
or U6731 (N_6731,N_6516,N_6566);
and U6732 (N_6732,N_6508,N_6544);
and U6733 (N_6733,N_6401,N_6529);
nand U6734 (N_6734,N_6457,N_6558);
nor U6735 (N_6735,N_6400,N_6561);
nor U6736 (N_6736,N_6548,N_6577);
or U6737 (N_6737,N_6515,N_6568);
xor U6738 (N_6738,N_6405,N_6420);
and U6739 (N_6739,N_6469,N_6494);
and U6740 (N_6740,N_6408,N_6456);
and U6741 (N_6741,N_6523,N_6589);
nor U6742 (N_6742,N_6494,N_6414);
nand U6743 (N_6743,N_6497,N_6588);
xnor U6744 (N_6744,N_6533,N_6561);
nand U6745 (N_6745,N_6522,N_6566);
or U6746 (N_6746,N_6466,N_6517);
nand U6747 (N_6747,N_6573,N_6551);
xor U6748 (N_6748,N_6410,N_6598);
and U6749 (N_6749,N_6443,N_6440);
and U6750 (N_6750,N_6427,N_6401);
or U6751 (N_6751,N_6404,N_6523);
xnor U6752 (N_6752,N_6560,N_6502);
or U6753 (N_6753,N_6591,N_6563);
or U6754 (N_6754,N_6503,N_6414);
nor U6755 (N_6755,N_6410,N_6435);
and U6756 (N_6756,N_6566,N_6458);
or U6757 (N_6757,N_6532,N_6569);
and U6758 (N_6758,N_6514,N_6511);
or U6759 (N_6759,N_6471,N_6493);
and U6760 (N_6760,N_6580,N_6591);
nor U6761 (N_6761,N_6445,N_6438);
nor U6762 (N_6762,N_6424,N_6440);
nor U6763 (N_6763,N_6540,N_6537);
and U6764 (N_6764,N_6558,N_6551);
and U6765 (N_6765,N_6456,N_6484);
and U6766 (N_6766,N_6434,N_6447);
xor U6767 (N_6767,N_6482,N_6551);
or U6768 (N_6768,N_6570,N_6466);
nand U6769 (N_6769,N_6429,N_6425);
nand U6770 (N_6770,N_6590,N_6474);
or U6771 (N_6771,N_6593,N_6420);
xnor U6772 (N_6772,N_6520,N_6570);
and U6773 (N_6773,N_6517,N_6468);
or U6774 (N_6774,N_6481,N_6471);
or U6775 (N_6775,N_6493,N_6466);
and U6776 (N_6776,N_6499,N_6564);
and U6777 (N_6777,N_6567,N_6524);
nand U6778 (N_6778,N_6509,N_6464);
or U6779 (N_6779,N_6508,N_6521);
nor U6780 (N_6780,N_6424,N_6519);
or U6781 (N_6781,N_6403,N_6448);
nor U6782 (N_6782,N_6434,N_6522);
or U6783 (N_6783,N_6500,N_6555);
or U6784 (N_6784,N_6501,N_6574);
or U6785 (N_6785,N_6513,N_6439);
or U6786 (N_6786,N_6525,N_6553);
nand U6787 (N_6787,N_6423,N_6489);
nand U6788 (N_6788,N_6595,N_6432);
nor U6789 (N_6789,N_6487,N_6444);
nor U6790 (N_6790,N_6507,N_6471);
and U6791 (N_6791,N_6459,N_6454);
xnor U6792 (N_6792,N_6505,N_6430);
nor U6793 (N_6793,N_6493,N_6444);
and U6794 (N_6794,N_6592,N_6486);
or U6795 (N_6795,N_6441,N_6581);
and U6796 (N_6796,N_6457,N_6534);
or U6797 (N_6797,N_6511,N_6508);
xnor U6798 (N_6798,N_6434,N_6592);
nand U6799 (N_6799,N_6468,N_6511);
xor U6800 (N_6800,N_6702,N_6705);
nand U6801 (N_6801,N_6679,N_6650);
or U6802 (N_6802,N_6680,N_6669);
or U6803 (N_6803,N_6634,N_6636);
or U6804 (N_6804,N_6642,N_6731);
and U6805 (N_6805,N_6677,N_6749);
nand U6806 (N_6806,N_6689,N_6644);
nor U6807 (N_6807,N_6746,N_6715);
xnor U6808 (N_6808,N_6780,N_6791);
nand U6809 (N_6809,N_6739,N_6784);
and U6810 (N_6810,N_6700,N_6673);
nand U6811 (N_6811,N_6750,N_6652);
or U6812 (N_6812,N_6612,N_6733);
xor U6813 (N_6813,N_6633,N_6785);
nand U6814 (N_6814,N_6768,N_6628);
xor U6815 (N_6815,N_6719,N_6646);
xnor U6816 (N_6816,N_6706,N_6766);
and U6817 (N_6817,N_6714,N_6797);
nand U6818 (N_6818,N_6638,N_6683);
and U6819 (N_6819,N_6794,N_6615);
nand U6820 (N_6820,N_6657,N_6619);
nand U6821 (N_6821,N_6658,N_6606);
nand U6822 (N_6822,N_6748,N_6793);
xnor U6823 (N_6823,N_6608,N_6653);
nand U6824 (N_6824,N_6631,N_6602);
and U6825 (N_6825,N_6682,N_6774);
nand U6826 (N_6826,N_6639,N_6616);
and U6827 (N_6827,N_6693,N_6675);
nor U6828 (N_6828,N_6708,N_6681);
nand U6829 (N_6829,N_6713,N_6796);
and U6830 (N_6830,N_6778,N_6789);
nor U6831 (N_6831,N_6655,N_6729);
xor U6832 (N_6832,N_6697,N_6686);
nor U6833 (N_6833,N_6742,N_6699);
or U6834 (N_6834,N_6760,N_6643);
nand U6835 (N_6835,N_6757,N_6692);
nor U6836 (N_6836,N_6730,N_6776);
or U6837 (N_6837,N_6703,N_6745);
xnor U6838 (N_6838,N_6648,N_6779);
or U6839 (N_6839,N_6623,N_6663);
nor U6840 (N_6840,N_6754,N_6721);
or U6841 (N_6841,N_6605,N_6737);
or U6842 (N_6842,N_6747,N_6763);
nand U6843 (N_6843,N_6752,N_6620);
xor U6844 (N_6844,N_6764,N_6732);
and U6845 (N_6845,N_6711,N_6770);
xor U6846 (N_6846,N_6691,N_6662);
or U6847 (N_6847,N_6751,N_6775);
nand U6848 (N_6848,N_6649,N_6782);
nor U6849 (N_6849,N_6603,N_6790);
and U6850 (N_6850,N_6668,N_6607);
xor U6851 (N_6851,N_6672,N_6684);
and U6852 (N_6852,N_6661,N_6678);
or U6853 (N_6853,N_6736,N_6799);
nand U6854 (N_6854,N_6718,N_6629);
nand U6855 (N_6855,N_6722,N_6664);
nand U6856 (N_6856,N_6734,N_6647);
xor U6857 (N_6857,N_6630,N_6773);
nand U6858 (N_6858,N_6694,N_6792);
xnor U6859 (N_6859,N_6723,N_6618);
and U6860 (N_6860,N_6690,N_6676);
nor U6861 (N_6861,N_6667,N_6744);
xnor U6862 (N_6862,N_6753,N_6632);
nor U6863 (N_6863,N_6738,N_6614);
nor U6864 (N_6864,N_6709,N_6777);
nor U6865 (N_6865,N_6698,N_6670);
or U6866 (N_6866,N_6787,N_6610);
nand U6867 (N_6867,N_6666,N_6707);
and U6868 (N_6868,N_6601,N_6640);
or U6869 (N_6869,N_6767,N_6725);
nor U6870 (N_6870,N_6695,N_6617);
nor U6871 (N_6871,N_6637,N_6727);
nand U6872 (N_6872,N_6665,N_6624);
nor U6873 (N_6873,N_6635,N_6740);
or U6874 (N_6874,N_6735,N_6762);
xnor U6875 (N_6875,N_6685,N_6724);
or U6876 (N_6876,N_6626,N_6659);
nand U6877 (N_6877,N_6627,N_6651);
or U6878 (N_6878,N_6772,N_6716);
xor U6879 (N_6879,N_6717,N_6720);
nand U6880 (N_6880,N_6759,N_6728);
nor U6881 (N_6881,N_6743,N_6621);
or U6882 (N_6882,N_6795,N_6741);
nor U6883 (N_6883,N_6712,N_6604);
and U6884 (N_6884,N_6765,N_6611);
or U6885 (N_6885,N_6613,N_6755);
xnor U6886 (N_6886,N_6758,N_6783);
or U6887 (N_6887,N_6710,N_6645);
nor U6888 (N_6888,N_6701,N_6726);
xnor U6889 (N_6889,N_6654,N_6771);
and U6890 (N_6890,N_6671,N_6622);
nand U6891 (N_6891,N_6660,N_6788);
or U6892 (N_6892,N_6704,N_6625);
xor U6893 (N_6893,N_6786,N_6600);
or U6894 (N_6894,N_6656,N_6696);
and U6895 (N_6895,N_6674,N_6781);
nor U6896 (N_6896,N_6769,N_6761);
nor U6897 (N_6897,N_6688,N_6756);
and U6898 (N_6898,N_6798,N_6687);
or U6899 (N_6899,N_6609,N_6641);
or U6900 (N_6900,N_6667,N_6736);
nand U6901 (N_6901,N_6664,N_6799);
nand U6902 (N_6902,N_6614,N_6683);
xnor U6903 (N_6903,N_6786,N_6760);
nand U6904 (N_6904,N_6655,N_6686);
xor U6905 (N_6905,N_6669,N_6788);
nand U6906 (N_6906,N_6665,N_6695);
nor U6907 (N_6907,N_6618,N_6796);
nor U6908 (N_6908,N_6671,N_6674);
or U6909 (N_6909,N_6758,N_6673);
xnor U6910 (N_6910,N_6667,N_6730);
and U6911 (N_6911,N_6796,N_6667);
and U6912 (N_6912,N_6786,N_6708);
nor U6913 (N_6913,N_6687,N_6791);
or U6914 (N_6914,N_6671,N_6627);
and U6915 (N_6915,N_6732,N_6643);
nand U6916 (N_6916,N_6659,N_6668);
or U6917 (N_6917,N_6676,N_6757);
xor U6918 (N_6918,N_6636,N_6605);
nor U6919 (N_6919,N_6635,N_6717);
nor U6920 (N_6920,N_6741,N_6634);
xor U6921 (N_6921,N_6602,N_6630);
and U6922 (N_6922,N_6646,N_6685);
nand U6923 (N_6923,N_6649,N_6644);
xnor U6924 (N_6924,N_6606,N_6688);
or U6925 (N_6925,N_6751,N_6677);
and U6926 (N_6926,N_6647,N_6754);
nor U6927 (N_6927,N_6783,N_6616);
nand U6928 (N_6928,N_6654,N_6614);
and U6929 (N_6929,N_6754,N_6732);
nand U6930 (N_6930,N_6665,N_6760);
or U6931 (N_6931,N_6615,N_6732);
nor U6932 (N_6932,N_6679,N_6755);
or U6933 (N_6933,N_6771,N_6695);
and U6934 (N_6934,N_6744,N_6723);
and U6935 (N_6935,N_6624,N_6630);
or U6936 (N_6936,N_6791,N_6646);
or U6937 (N_6937,N_6619,N_6755);
nor U6938 (N_6938,N_6639,N_6621);
nand U6939 (N_6939,N_6620,N_6647);
nor U6940 (N_6940,N_6752,N_6740);
and U6941 (N_6941,N_6618,N_6661);
nor U6942 (N_6942,N_6680,N_6725);
nor U6943 (N_6943,N_6726,N_6755);
nor U6944 (N_6944,N_6632,N_6771);
nor U6945 (N_6945,N_6611,N_6639);
or U6946 (N_6946,N_6742,N_6616);
and U6947 (N_6947,N_6707,N_6749);
xnor U6948 (N_6948,N_6764,N_6751);
and U6949 (N_6949,N_6635,N_6648);
xor U6950 (N_6950,N_6623,N_6709);
or U6951 (N_6951,N_6617,N_6758);
xnor U6952 (N_6952,N_6625,N_6680);
xor U6953 (N_6953,N_6768,N_6618);
and U6954 (N_6954,N_6601,N_6679);
nand U6955 (N_6955,N_6740,N_6696);
nand U6956 (N_6956,N_6789,N_6772);
and U6957 (N_6957,N_6767,N_6648);
xnor U6958 (N_6958,N_6678,N_6613);
and U6959 (N_6959,N_6715,N_6769);
xnor U6960 (N_6960,N_6603,N_6610);
nand U6961 (N_6961,N_6753,N_6691);
nor U6962 (N_6962,N_6621,N_6649);
xnor U6963 (N_6963,N_6675,N_6737);
or U6964 (N_6964,N_6729,N_6726);
nor U6965 (N_6965,N_6683,N_6667);
and U6966 (N_6966,N_6659,N_6614);
nand U6967 (N_6967,N_6658,N_6795);
xnor U6968 (N_6968,N_6632,N_6685);
xor U6969 (N_6969,N_6627,N_6703);
and U6970 (N_6970,N_6727,N_6694);
nor U6971 (N_6971,N_6638,N_6667);
nor U6972 (N_6972,N_6739,N_6694);
nand U6973 (N_6973,N_6608,N_6612);
or U6974 (N_6974,N_6665,N_6620);
xnor U6975 (N_6975,N_6638,N_6793);
nor U6976 (N_6976,N_6690,N_6620);
xor U6977 (N_6977,N_6749,N_6658);
or U6978 (N_6978,N_6666,N_6737);
nor U6979 (N_6979,N_6647,N_6760);
or U6980 (N_6980,N_6634,N_6700);
or U6981 (N_6981,N_6701,N_6798);
nand U6982 (N_6982,N_6627,N_6657);
and U6983 (N_6983,N_6629,N_6633);
and U6984 (N_6984,N_6724,N_6609);
or U6985 (N_6985,N_6646,N_6683);
xnor U6986 (N_6986,N_6633,N_6713);
nor U6987 (N_6987,N_6786,N_6611);
nand U6988 (N_6988,N_6798,N_6752);
xnor U6989 (N_6989,N_6622,N_6758);
nor U6990 (N_6990,N_6693,N_6741);
nor U6991 (N_6991,N_6699,N_6673);
nor U6992 (N_6992,N_6740,N_6663);
xnor U6993 (N_6993,N_6640,N_6748);
nand U6994 (N_6994,N_6660,N_6675);
nand U6995 (N_6995,N_6757,N_6760);
nor U6996 (N_6996,N_6732,N_6793);
nand U6997 (N_6997,N_6712,N_6671);
nor U6998 (N_6998,N_6749,N_6778);
nor U6999 (N_6999,N_6747,N_6733);
and U7000 (N_7000,N_6821,N_6835);
or U7001 (N_7001,N_6808,N_6965);
and U7002 (N_7002,N_6879,N_6931);
nand U7003 (N_7003,N_6812,N_6809);
or U7004 (N_7004,N_6887,N_6924);
xor U7005 (N_7005,N_6846,N_6913);
xor U7006 (N_7006,N_6875,N_6828);
nor U7007 (N_7007,N_6992,N_6827);
xor U7008 (N_7008,N_6896,N_6807);
nand U7009 (N_7009,N_6991,N_6868);
and U7010 (N_7010,N_6825,N_6984);
and U7011 (N_7011,N_6970,N_6874);
xnor U7012 (N_7012,N_6982,N_6806);
xnor U7013 (N_7013,N_6902,N_6864);
nand U7014 (N_7014,N_6983,N_6901);
nor U7015 (N_7015,N_6976,N_6811);
or U7016 (N_7016,N_6939,N_6881);
and U7017 (N_7017,N_6973,N_6883);
and U7018 (N_7018,N_6941,N_6918);
nor U7019 (N_7019,N_6927,N_6969);
or U7020 (N_7020,N_6814,N_6859);
nor U7021 (N_7021,N_6888,N_6986);
and U7022 (N_7022,N_6886,N_6819);
or U7023 (N_7023,N_6999,N_6904);
xor U7024 (N_7024,N_6945,N_6925);
and U7025 (N_7025,N_6951,N_6805);
nor U7026 (N_7026,N_6958,N_6840);
and U7027 (N_7027,N_6909,N_6844);
and U7028 (N_7028,N_6975,N_6952);
or U7029 (N_7029,N_6802,N_6907);
nand U7030 (N_7030,N_6947,N_6877);
or U7031 (N_7031,N_6933,N_6943);
nor U7032 (N_7032,N_6987,N_6979);
nand U7033 (N_7033,N_6977,N_6855);
nor U7034 (N_7034,N_6826,N_6963);
xor U7035 (N_7035,N_6847,N_6856);
xor U7036 (N_7036,N_6823,N_6961);
or U7037 (N_7037,N_6900,N_6995);
nand U7038 (N_7038,N_6853,N_6833);
and U7039 (N_7039,N_6972,N_6928);
xor U7040 (N_7040,N_6930,N_6978);
or U7041 (N_7041,N_6955,N_6850);
nor U7042 (N_7042,N_6822,N_6895);
xor U7043 (N_7043,N_6842,N_6923);
or U7044 (N_7044,N_6870,N_6938);
nand U7045 (N_7045,N_6861,N_6843);
or U7046 (N_7046,N_6921,N_6820);
nor U7047 (N_7047,N_6839,N_6985);
nand U7048 (N_7048,N_6993,N_6932);
nor U7049 (N_7049,N_6981,N_6920);
and U7050 (N_7050,N_6989,N_6801);
nor U7051 (N_7051,N_6974,N_6967);
nand U7052 (N_7052,N_6890,N_6867);
nor U7053 (N_7053,N_6937,N_6836);
nand U7054 (N_7054,N_6954,N_6800);
nand U7055 (N_7055,N_6862,N_6953);
or U7056 (N_7056,N_6950,N_6813);
xnor U7057 (N_7057,N_6966,N_6815);
xor U7058 (N_7058,N_6916,N_6818);
or U7059 (N_7059,N_6948,N_6912);
nand U7060 (N_7060,N_6971,N_6857);
and U7061 (N_7061,N_6832,N_6949);
nor U7062 (N_7062,N_6891,N_6980);
nor U7063 (N_7063,N_6838,N_6851);
or U7064 (N_7064,N_6917,N_6880);
xnor U7065 (N_7065,N_6858,N_6914);
or U7066 (N_7066,N_6869,N_6968);
or U7067 (N_7067,N_6816,N_6804);
nor U7068 (N_7068,N_6942,N_6817);
xor U7069 (N_7069,N_6834,N_6898);
nor U7070 (N_7070,N_6926,N_6911);
or U7071 (N_7071,N_6882,N_6936);
or U7072 (N_7072,N_6860,N_6959);
xor U7073 (N_7073,N_6903,N_6824);
xor U7074 (N_7074,N_6849,N_6863);
or U7075 (N_7075,N_6946,N_6960);
xnor U7076 (N_7076,N_6866,N_6873);
xnor U7077 (N_7077,N_6871,N_6831);
or U7078 (N_7078,N_6906,N_6810);
and U7079 (N_7079,N_6910,N_6830);
xor U7080 (N_7080,N_6803,N_6878);
nand U7081 (N_7081,N_6905,N_6964);
xnor U7082 (N_7082,N_6929,N_6893);
or U7083 (N_7083,N_6884,N_6876);
nor U7084 (N_7084,N_6845,N_6872);
nand U7085 (N_7085,N_6988,N_6854);
xor U7086 (N_7086,N_6998,N_6919);
nor U7087 (N_7087,N_6897,N_6829);
nand U7088 (N_7088,N_6934,N_6837);
nor U7089 (N_7089,N_6996,N_6908);
nand U7090 (N_7090,N_6841,N_6994);
nand U7091 (N_7091,N_6894,N_6848);
nand U7092 (N_7092,N_6956,N_6962);
and U7093 (N_7093,N_6899,N_6892);
and U7094 (N_7094,N_6944,N_6957);
xor U7095 (N_7095,N_6990,N_6865);
and U7096 (N_7096,N_6935,N_6997);
xor U7097 (N_7097,N_6922,N_6915);
nor U7098 (N_7098,N_6885,N_6940);
or U7099 (N_7099,N_6852,N_6889);
nand U7100 (N_7100,N_6957,N_6808);
xor U7101 (N_7101,N_6960,N_6827);
and U7102 (N_7102,N_6888,N_6923);
and U7103 (N_7103,N_6812,N_6887);
xnor U7104 (N_7104,N_6861,N_6817);
nand U7105 (N_7105,N_6810,N_6894);
nor U7106 (N_7106,N_6913,N_6974);
or U7107 (N_7107,N_6897,N_6856);
and U7108 (N_7108,N_6907,N_6994);
nor U7109 (N_7109,N_6968,N_6878);
nor U7110 (N_7110,N_6865,N_6849);
nand U7111 (N_7111,N_6903,N_6835);
nand U7112 (N_7112,N_6813,N_6878);
nor U7113 (N_7113,N_6810,N_6922);
or U7114 (N_7114,N_6986,N_6910);
and U7115 (N_7115,N_6826,N_6822);
or U7116 (N_7116,N_6885,N_6897);
and U7117 (N_7117,N_6945,N_6868);
or U7118 (N_7118,N_6930,N_6948);
and U7119 (N_7119,N_6902,N_6933);
nor U7120 (N_7120,N_6819,N_6982);
and U7121 (N_7121,N_6956,N_6901);
and U7122 (N_7122,N_6831,N_6843);
or U7123 (N_7123,N_6943,N_6928);
nand U7124 (N_7124,N_6883,N_6947);
nand U7125 (N_7125,N_6810,N_6925);
and U7126 (N_7126,N_6804,N_6957);
xnor U7127 (N_7127,N_6922,N_6970);
and U7128 (N_7128,N_6902,N_6840);
nor U7129 (N_7129,N_6864,N_6887);
or U7130 (N_7130,N_6813,N_6998);
nor U7131 (N_7131,N_6894,N_6861);
xnor U7132 (N_7132,N_6978,N_6934);
or U7133 (N_7133,N_6853,N_6942);
and U7134 (N_7134,N_6957,N_6941);
and U7135 (N_7135,N_6927,N_6902);
and U7136 (N_7136,N_6948,N_6921);
nand U7137 (N_7137,N_6845,N_6871);
nand U7138 (N_7138,N_6819,N_6834);
nand U7139 (N_7139,N_6956,N_6938);
nor U7140 (N_7140,N_6961,N_6846);
and U7141 (N_7141,N_6873,N_6842);
nand U7142 (N_7142,N_6935,N_6936);
nand U7143 (N_7143,N_6958,N_6872);
or U7144 (N_7144,N_6800,N_6867);
or U7145 (N_7145,N_6804,N_6831);
or U7146 (N_7146,N_6881,N_6887);
nand U7147 (N_7147,N_6989,N_6928);
and U7148 (N_7148,N_6816,N_6900);
xnor U7149 (N_7149,N_6934,N_6950);
or U7150 (N_7150,N_6859,N_6930);
or U7151 (N_7151,N_6875,N_6832);
nand U7152 (N_7152,N_6881,N_6888);
and U7153 (N_7153,N_6817,N_6923);
and U7154 (N_7154,N_6825,N_6965);
xnor U7155 (N_7155,N_6849,N_6993);
and U7156 (N_7156,N_6904,N_6997);
nor U7157 (N_7157,N_6810,N_6800);
nand U7158 (N_7158,N_6854,N_6833);
or U7159 (N_7159,N_6995,N_6940);
nor U7160 (N_7160,N_6938,N_6809);
nor U7161 (N_7161,N_6946,N_6894);
and U7162 (N_7162,N_6886,N_6806);
xor U7163 (N_7163,N_6840,N_6976);
nand U7164 (N_7164,N_6982,N_6914);
nand U7165 (N_7165,N_6958,N_6837);
and U7166 (N_7166,N_6871,N_6813);
nor U7167 (N_7167,N_6995,N_6902);
and U7168 (N_7168,N_6818,N_6928);
xor U7169 (N_7169,N_6902,N_6890);
nor U7170 (N_7170,N_6807,N_6822);
xnor U7171 (N_7171,N_6979,N_6875);
nor U7172 (N_7172,N_6967,N_6982);
nor U7173 (N_7173,N_6976,N_6871);
xor U7174 (N_7174,N_6816,N_6853);
nor U7175 (N_7175,N_6832,N_6986);
nor U7176 (N_7176,N_6821,N_6869);
xnor U7177 (N_7177,N_6824,N_6810);
nor U7178 (N_7178,N_6873,N_6942);
xor U7179 (N_7179,N_6841,N_6889);
nand U7180 (N_7180,N_6972,N_6992);
and U7181 (N_7181,N_6939,N_6831);
or U7182 (N_7182,N_6854,N_6921);
and U7183 (N_7183,N_6954,N_6859);
or U7184 (N_7184,N_6964,N_6851);
or U7185 (N_7185,N_6821,N_6907);
nand U7186 (N_7186,N_6958,N_6893);
nand U7187 (N_7187,N_6902,N_6964);
and U7188 (N_7188,N_6906,N_6876);
and U7189 (N_7189,N_6979,N_6841);
nor U7190 (N_7190,N_6815,N_6887);
nor U7191 (N_7191,N_6826,N_6934);
nand U7192 (N_7192,N_6969,N_6827);
xor U7193 (N_7193,N_6967,N_6918);
xor U7194 (N_7194,N_6839,N_6819);
nor U7195 (N_7195,N_6852,N_6914);
nor U7196 (N_7196,N_6952,N_6996);
xnor U7197 (N_7197,N_6934,N_6888);
xnor U7198 (N_7198,N_6996,N_6947);
xor U7199 (N_7199,N_6974,N_6899);
nand U7200 (N_7200,N_7168,N_7122);
xnor U7201 (N_7201,N_7062,N_7053);
nor U7202 (N_7202,N_7070,N_7058);
nor U7203 (N_7203,N_7051,N_7159);
or U7204 (N_7204,N_7126,N_7130);
xor U7205 (N_7205,N_7115,N_7094);
nand U7206 (N_7206,N_7073,N_7014);
or U7207 (N_7207,N_7106,N_7108);
nor U7208 (N_7208,N_7135,N_7137);
nand U7209 (N_7209,N_7012,N_7023);
nor U7210 (N_7210,N_7161,N_7044);
or U7211 (N_7211,N_7133,N_7024);
or U7212 (N_7212,N_7020,N_7118);
or U7213 (N_7213,N_7072,N_7191);
xor U7214 (N_7214,N_7063,N_7178);
nand U7215 (N_7215,N_7165,N_7142);
and U7216 (N_7216,N_7117,N_7179);
nand U7217 (N_7217,N_7140,N_7113);
xnor U7218 (N_7218,N_7145,N_7158);
and U7219 (N_7219,N_7160,N_7138);
xnor U7220 (N_7220,N_7195,N_7190);
xnor U7221 (N_7221,N_7013,N_7010);
xor U7222 (N_7222,N_7171,N_7187);
nor U7223 (N_7223,N_7131,N_7186);
nor U7224 (N_7224,N_7156,N_7006);
xor U7225 (N_7225,N_7127,N_7128);
nand U7226 (N_7226,N_7180,N_7068);
nand U7227 (N_7227,N_7098,N_7121);
and U7228 (N_7228,N_7093,N_7005);
nand U7229 (N_7229,N_7055,N_7077);
nor U7230 (N_7230,N_7086,N_7147);
and U7231 (N_7231,N_7092,N_7041);
and U7232 (N_7232,N_7065,N_7054);
or U7233 (N_7233,N_7096,N_7114);
nor U7234 (N_7234,N_7066,N_7166);
nand U7235 (N_7235,N_7153,N_7148);
nand U7236 (N_7236,N_7132,N_7155);
or U7237 (N_7237,N_7002,N_7112);
nor U7238 (N_7238,N_7030,N_7034);
xor U7239 (N_7239,N_7083,N_7033);
xnor U7240 (N_7240,N_7087,N_7031);
nand U7241 (N_7241,N_7154,N_7004);
or U7242 (N_7242,N_7157,N_7037);
nor U7243 (N_7243,N_7175,N_7074);
nand U7244 (N_7244,N_7163,N_7109);
nor U7245 (N_7245,N_7018,N_7123);
nor U7246 (N_7246,N_7015,N_7176);
nand U7247 (N_7247,N_7001,N_7189);
and U7248 (N_7248,N_7043,N_7119);
xor U7249 (N_7249,N_7197,N_7177);
nor U7250 (N_7250,N_7011,N_7067);
xor U7251 (N_7251,N_7080,N_7144);
xor U7252 (N_7252,N_7100,N_7172);
or U7253 (N_7253,N_7017,N_7136);
and U7254 (N_7254,N_7170,N_7151);
and U7255 (N_7255,N_7110,N_7078);
or U7256 (N_7256,N_7082,N_7183);
and U7257 (N_7257,N_7125,N_7139);
xor U7258 (N_7258,N_7025,N_7009);
nor U7259 (N_7259,N_7076,N_7090);
and U7260 (N_7260,N_7103,N_7036);
xor U7261 (N_7261,N_7181,N_7129);
or U7262 (N_7262,N_7185,N_7134);
nor U7263 (N_7263,N_7003,N_7032);
and U7264 (N_7264,N_7173,N_7035);
nand U7265 (N_7265,N_7045,N_7102);
nor U7266 (N_7266,N_7146,N_7050);
xor U7267 (N_7267,N_7060,N_7056);
nand U7268 (N_7268,N_7016,N_7088);
xnor U7269 (N_7269,N_7059,N_7120);
nor U7270 (N_7270,N_7079,N_7040);
or U7271 (N_7271,N_7039,N_7174);
xor U7272 (N_7272,N_7107,N_7169);
nand U7273 (N_7273,N_7199,N_7000);
nand U7274 (N_7274,N_7021,N_7089);
nand U7275 (N_7275,N_7022,N_7061);
or U7276 (N_7276,N_7167,N_7194);
nor U7277 (N_7277,N_7105,N_7099);
and U7278 (N_7278,N_7198,N_7071);
nor U7279 (N_7279,N_7064,N_7184);
nand U7280 (N_7280,N_7046,N_7196);
or U7281 (N_7281,N_7095,N_7192);
and U7282 (N_7282,N_7019,N_7193);
xnor U7283 (N_7283,N_7097,N_7150);
or U7284 (N_7284,N_7162,N_7152);
nor U7285 (N_7285,N_7164,N_7052);
xnor U7286 (N_7286,N_7008,N_7091);
or U7287 (N_7287,N_7084,N_7026);
xor U7288 (N_7288,N_7182,N_7049);
and U7289 (N_7289,N_7042,N_7027);
xnor U7290 (N_7290,N_7069,N_7047);
or U7291 (N_7291,N_7188,N_7085);
xnor U7292 (N_7292,N_7104,N_7075);
nor U7293 (N_7293,N_7116,N_7028);
or U7294 (N_7294,N_7007,N_7101);
nand U7295 (N_7295,N_7111,N_7143);
and U7296 (N_7296,N_7048,N_7149);
or U7297 (N_7297,N_7081,N_7029);
or U7298 (N_7298,N_7057,N_7038);
or U7299 (N_7299,N_7141,N_7124);
nand U7300 (N_7300,N_7155,N_7103);
nand U7301 (N_7301,N_7008,N_7131);
xnor U7302 (N_7302,N_7068,N_7093);
and U7303 (N_7303,N_7046,N_7187);
nor U7304 (N_7304,N_7109,N_7002);
and U7305 (N_7305,N_7182,N_7133);
and U7306 (N_7306,N_7100,N_7076);
nor U7307 (N_7307,N_7047,N_7188);
and U7308 (N_7308,N_7082,N_7158);
nand U7309 (N_7309,N_7094,N_7082);
xnor U7310 (N_7310,N_7056,N_7035);
nor U7311 (N_7311,N_7165,N_7039);
nand U7312 (N_7312,N_7005,N_7015);
or U7313 (N_7313,N_7037,N_7020);
xnor U7314 (N_7314,N_7072,N_7157);
nand U7315 (N_7315,N_7096,N_7006);
xnor U7316 (N_7316,N_7007,N_7119);
nor U7317 (N_7317,N_7110,N_7137);
and U7318 (N_7318,N_7159,N_7047);
nor U7319 (N_7319,N_7048,N_7039);
or U7320 (N_7320,N_7007,N_7002);
or U7321 (N_7321,N_7142,N_7047);
nor U7322 (N_7322,N_7124,N_7096);
and U7323 (N_7323,N_7167,N_7094);
and U7324 (N_7324,N_7094,N_7145);
and U7325 (N_7325,N_7097,N_7076);
xor U7326 (N_7326,N_7042,N_7004);
or U7327 (N_7327,N_7066,N_7163);
or U7328 (N_7328,N_7005,N_7161);
and U7329 (N_7329,N_7023,N_7017);
and U7330 (N_7330,N_7140,N_7176);
nor U7331 (N_7331,N_7066,N_7110);
xor U7332 (N_7332,N_7051,N_7197);
and U7333 (N_7333,N_7157,N_7170);
nand U7334 (N_7334,N_7166,N_7082);
or U7335 (N_7335,N_7029,N_7067);
nor U7336 (N_7336,N_7103,N_7086);
xnor U7337 (N_7337,N_7062,N_7138);
or U7338 (N_7338,N_7125,N_7111);
nand U7339 (N_7339,N_7136,N_7187);
or U7340 (N_7340,N_7156,N_7022);
nor U7341 (N_7341,N_7181,N_7077);
nor U7342 (N_7342,N_7005,N_7171);
or U7343 (N_7343,N_7018,N_7059);
nand U7344 (N_7344,N_7185,N_7037);
nor U7345 (N_7345,N_7039,N_7079);
xor U7346 (N_7346,N_7116,N_7015);
xnor U7347 (N_7347,N_7149,N_7031);
nor U7348 (N_7348,N_7186,N_7192);
nand U7349 (N_7349,N_7035,N_7104);
xor U7350 (N_7350,N_7021,N_7114);
xor U7351 (N_7351,N_7091,N_7107);
xor U7352 (N_7352,N_7164,N_7129);
nand U7353 (N_7353,N_7054,N_7097);
and U7354 (N_7354,N_7188,N_7173);
xor U7355 (N_7355,N_7110,N_7029);
and U7356 (N_7356,N_7000,N_7143);
nor U7357 (N_7357,N_7047,N_7157);
nor U7358 (N_7358,N_7073,N_7082);
and U7359 (N_7359,N_7013,N_7150);
and U7360 (N_7360,N_7098,N_7040);
xnor U7361 (N_7361,N_7154,N_7137);
and U7362 (N_7362,N_7145,N_7012);
and U7363 (N_7363,N_7027,N_7083);
nand U7364 (N_7364,N_7094,N_7056);
xnor U7365 (N_7365,N_7166,N_7022);
nor U7366 (N_7366,N_7177,N_7133);
or U7367 (N_7367,N_7081,N_7054);
and U7368 (N_7368,N_7010,N_7012);
or U7369 (N_7369,N_7150,N_7023);
nand U7370 (N_7370,N_7167,N_7140);
xnor U7371 (N_7371,N_7068,N_7199);
and U7372 (N_7372,N_7151,N_7095);
or U7373 (N_7373,N_7034,N_7006);
nor U7374 (N_7374,N_7034,N_7058);
and U7375 (N_7375,N_7070,N_7078);
and U7376 (N_7376,N_7042,N_7005);
or U7377 (N_7377,N_7147,N_7159);
nor U7378 (N_7378,N_7145,N_7072);
or U7379 (N_7379,N_7147,N_7078);
nand U7380 (N_7380,N_7165,N_7182);
nand U7381 (N_7381,N_7194,N_7001);
nor U7382 (N_7382,N_7072,N_7084);
xnor U7383 (N_7383,N_7021,N_7093);
and U7384 (N_7384,N_7165,N_7107);
and U7385 (N_7385,N_7178,N_7066);
and U7386 (N_7386,N_7143,N_7106);
xnor U7387 (N_7387,N_7049,N_7100);
or U7388 (N_7388,N_7130,N_7012);
xnor U7389 (N_7389,N_7083,N_7001);
nand U7390 (N_7390,N_7040,N_7068);
and U7391 (N_7391,N_7051,N_7158);
xor U7392 (N_7392,N_7094,N_7162);
xnor U7393 (N_7393,N_7176,N_7096);
nor U7394 (N_7394,N_7103,N_7177);
nor U7395 (N_7395,N_7096,N_7140);
and U7396 (N_7396,N_7110,N_7179);
xor U7397 (N_7397,N_7139,N_7163);
and U7398 (N_7398,N_7015,N_7061);
and U7399 (N_7399,N_7169,N_7088);
and U7400 (N_7400,N_7244,N_7354);
or U7401 (N_7401,N_7395,N_7235);
nor U7402 (N_7402,N_7264,N_7392);
nand U7403 (N_7403,N_7359,N_7218);
xnor U7404 (N_7404,N_7257,N_7387);
or U7405 (N_7405,N_7315,N_7241);
or U7406 (N_7406,N_7310,N_7238);
xor U7407 (N_7407,N_7337,N_7249);
xor U7408 (N_7408,N_7302,N_7390);
and U7409 (N_7409,N_7393,N_7323);
or U7410 (N_7410,N_7230,N_7345);
xor U7411 (N_7411,N_7374,N_7263);
nand U7412 (N_7412,N_7367,N_7217);
and U7413 (N_7413,N_7386,N_7330);
xnor U7414 (N_7414,N_7294,N_7366);
or U7415 (N_7415,N_7360,N_7222);
or U7416 (N_7416,N_7388,N_7253);
or U7417 (N_7417,N_7389,N_7226);
and U7418 (N_7418,N_7240,N_7279);
and U7419 (N_7419,N_7258,N_7375);
or U7420 (N_7420,N_7364,N_7385);
or U7421 (N_7421,N_7382,N_7399);
nor U7422 (N_7422,N_7308,N_7334);
nand U7423 (N_7423,N_7358,N_7316);
nand U7424 (N_7424,N_7396,N_7321);
and U7425 (N_7425,N_7391,N_7259);
xnor U7426 (N_7426,N_7333,N_7381);
nor U7427 (N_7427,N_7261,N_7246);
xnor U7428 (N_7428,N_7232,N_7336);
xnor U7429 (N_7429,N_7312,N_7225);
or U7430 (N_7430,N_7346,N_7295);
nor U7431 (N_7431,N_7377,N_7309);
xor U7432 (N_7432,N_7280,N_7207);
nand U7433 (N_7433,N_7320,N_7229);
xnor U7434 (N_7434,N_7201,N_7324);
nand U7435 (N_7435,N_7234,N_7273);
or U7436 (N_7436,N_7384,N_7233);
nor U7437 (N_7437,N_7205,N_7340);
nand U7438 (N_7438,N_7210,N_7371);
nor U7439 (N_7439,N_7267,N_7221);
or U7440 (N_7440,N_7306,N_7304);
or U7441 (N_7441,N_7296,N_7228);
xnor U7442 (N_7442,N_7327,N_7204);
and U7443 (N_7443,N_7202,N_7300);
nand U7444 (N_7444,N_7219,N_7361);
xor U7445 (N_7445,N_7383,N_7332);
xnor U7446 (N_7446,N_7290,N_7292);
xnor U7447 (N_7447,N_7299,N_7255);
nand U7448 (N_7448,N_7365,N_7379);
nor U7449 (N_7449,N_7224,N_7339);
nand U7450 (N_7450,N_7293,N_7350);
nand U7451 (N_7451,N_7376,N_7301);
nor U7452 (N_7452,N_7322,N_7344);
xnor U7453 (N_7453,N_7239,N_7254);
or U7454 (N_7454,N_7227,N_7370);
nand U7455 (N_7455,N_7380,N_7352);
nor U7456 (N_7456,N_7343,N_7208);
xnor U7457 (N_7457,N_7398,N_7328);
nand U7458 (N_7458,N_7266,N_7285);
and U7459 (N_7459,N_7260,N_7338);
nand U7460 (N_7460,N_7215,N_7251);
xnor U7461 (N_7461,N_7209,N_7278);
or U7462 (N_7462,N_7265,N_7331);
xor U7463 (N_7463,N_7283,N_7319);
nor U7464 (N_7464,N_7270,N_7313);
nand U7465 (N_7465,N_7378,N_7372);
nand U7466 (N_7466,N_7348,N_7269);
xor U7467 (N_7467,N_7369,N_7281);
nand U7468 (N_7468,N_7200,N_7318);
and U7469 (N_7469,N_7213,N_7214);
nand U7470 (N_7470,N_7203,N_7357);
nor U7471 (N_7471,N_7262,N_7286);
nand U7472 (N_7472,N_7326,N_7250);
or U7473 (N_7473,N_7243,N_7274);
or U7474 (N_7474,N_7341,N_7272);
nand U7475 (N_7475,N_7291,N_7394);
nor U7476 (N_7476,N_7237,N_7353);
nand U7477 (N_7477,N_7342,N_7351);
or U7478 (N_7478,N_7317,N_7368);
nand U7479 (N_7479,N_7256,N_7271);
nand U7480 (N_7480,N_7268,N_7329);
or U7481 (N_7481,N_7275,N_7231);
and U7482 (N_7482,N_7277,N_7311);
or U7483 (N_7483,N_7248,N_7288);
or U7484 (N_7484,N_7289,N_7206);
or U7485 (N_7485,N_7363,N_7223);
nand U7486 (N_7486,N_7297,N_7247);
and U7487 (N_7487,N_7307,N_7356);
or U7488 (N_7488,N_7349,N_7236);
nand U7489 (N_7489,N_7220,N_7216);
and U7490 (N_7490,N_7245,N_7303);
nor U7491 (N_7491,N_7287,N_7347);
or U7492 (N_7492,N_7242,N_7252);
nand U7493 (N_7493,N_7335,N_7305);
nand U7494 (N_7494,N_7282,N_7211);
nand U7495 (N_7495,N_7298,N_7314);
or U7496 (N_7496,N_7276,N_7373);
xnor U7497 (N_7497,N_7325,N_7284);
xnor U7498 (N_7498,N_7362,N_7212);
and U7499 (N_7499,N_7355,N_7397);
nand U7500 (N_7500,N_7213,N_7269);
nand U7501 (N_7501,N_7387,N_7307);
nor U7502 (N_7502,N_7212,N_7305);
nor U7503 (N_7503,N_7349,N_7333);
xor U7504 (N_7504,N_7262,N_7381);
nor U7505 (N_7505,N_7201,N_7231);
and U7506 (N_7506,N_7240,N_7231);
or U7507 (N_7507,N_7289,N_7271);
xor U7508 (N_7508,N_7310,N_7222);
or U7509 (N_7509,N_7371,N_7301);
and U7510 (N_7510,N_7285,N_7261);
nand U7511 (N_7511,N_7303,N_7292);
or U7512 (N_7512,N_7233,N_7354);
nand U7513 (N_7513,N_7242,N_7285);
nand U7514 (N_7514,N_7365,N_7254);
nor U7515 (N_7515,N_7390,N_7267);
nor U7516 (N_7516,N_7313,N_7383);
nand U7517 (N_7517,N_7336,N_7383);
xnor U7518 (N_7518,N_7336,N_7253);
xnor U7519 (N_7519,N_7232,N_7267);
and U7520 (N_7520,N_7357,N_7337);
or U7521 (N_7521,N_7315,N_7394);
nand U7522 (N_7522,N_7398,N_7340);
or U7523 (N_7523,N_7216,N_7249);
nor U7524 (N_7524,N_7221,N_7322);
xnor U7525 (N_7525,N_7224,N_7323);
or U7526 (N_7526,N_7244,N_7300);
and U7527 (N_7527,N_7339,N_7229);
and U7528 (N_7528,N_7307,N_7351);
or U7529 (N_7529,N_7223,N_7386);
nor U7530 (N_7530,N_7365,N_7371);
nand U7531 (N_7531,N_7292,N_7205);
nor U7532 (N_7532,N_7385,N_7314);
or U7533 (N_7533,N_7245,N_7209);
or U7534 (N_7534,N_7243,N_7318);
nor U7535 (N_7535,N_7384,N_7302);
nor U7536 (N_7536,N_7287,N_7299);
and U7537 (N_7537,N_7325,N_7370);
xnor U7538 (N_7538,N_7343,N_7294);
and U7539 (N_7539,N_7229,N_7373);
nor U7540 (N_7540,N_7312,N_7308);
or U7541 (N_7541,N_7315,N_7247);
or U7542 (N_7542,N_7349,N_7363);
or U7543 (N_7543,N_7306,N_7236);
and U7544 (N_7544,N_7247,N_7203);
or U7545 (N_7545,N_7305,N_7223);
and U7546 (N_7546,N_7249,N_7394);
nand U7547 (N_7547,N_7300,N_7391);
xnor U7548 (N_7548,N_7395,N_7273);
or U7549 (N_7549,N_7222,N_7300);
xor U7550 (N_7550,N_7268,N_7256);
and U7551 (N_7551,N_7293,N_7273);
nand U7552 (N_7552,N_7230,N_7235);
xnor U7553 (N_7553,N_7347,N_7259);
nand U7554 (N_7554,N_7205,N_7244);
nand U7555 (N_7555,N_7393,N_7301);
or U7556 (N_7556,N_7239,N_7245);
xnor U7557 (N_7557,N_7313,N_7230);
xnor U7558 (N_7558,N_7341,N_7279);
or U7559 (N_7559,N_7212,N_7279);
nand U7560 (N_7560,N_7209,N_7255);
nor U7561 (N_7561,N_7308,N_7382);
or U7562 (N_7562,N_7374,N_7217);
nand U7563 (N_7563,N_7394,N_7352);
or U7564 (N_7564,N_7289,N_7335);
xnor U7565 (N_7565,N_7302,N_7238);
or U7566 (N_7566,N_7279,N_7306);
or U7567 (N_7567,N_7376,N_7263);
and U7568 (N_7568,N_7200,N_7265);
and U7569 (N_7569,N_7212,N_7284);
nor U7570 (N_7570,N_7218,N_7395);
or U7571 (N_7571,N_7200,N_7394);
xor U7572 (N_7572,N_7226,N_7354);
xnor U7573 (N_7573,N_7374,N_7264);
and U7574 (N_7574,N_7221,N_7223);
nor U7575 (N_7575,N_7252,N_7281);
and U7576 (N_7576,N_7265,N_7241);
xor U7577 (N_7577,N_7375,N_7248);
xnor U7578 (N_7578,N_7391,N_7212);
xor U7579 (N_7579,N_7302,N_7357);
nor U7580 (N_7580,N_7318,N_7206);
nor U7581 (N_7581,N_7231,N_7313);
nand U7582 (N_7582,N_7218,N_7235);
and U7583 (N_7583,N_7393,N_7276);
nand U7584 (N_7584,N_7312,N_7372);
nor U7585 (N_7585,N_7202,N_7383);
or U7586 (N_7586,N_7313,N_7368);
nor U7587 (N_7587,N_7235,N_7261);
nor U7588 (N_7588,N_7319,N_7383);
or U7589 (N_7589,N_7355,N_7298);
nor U7590 (N_7590,N_7250,N_7232);
and U7591 (N_7591,N_7391,N_7224);
nor U7592 (N_7592,N_7272,N_7207);
nand U7593 (N_7593,N_7278,N_7289);
or U7594 (N_7594,N_7373,N_7265);
nor U7595 (N_7595,N_7295,N_7329);
xor U7596 (N_7596,N_7346,N_7244);
nor U7597 (N_7597,N_7274,N_7261);
nor U7598 (N_7598,N_7389,N_7276);
nand U7599 (N_7599,N_7338,N_7227);
and U7600 (N_7600,N_7452,N_7443);
nor U7601 (N_7601,N_7591,N_7537);
nor U7602 (N_7602,N_7402,N_7500);
xor U7603 (N_7603,N_7413,N_7415);
xor U7604 (N_7604,N_7409,N_7521);
xor U7605 (N_7605,N_7585,N_7567);
xor U7606 (N_7606,N_7531,N_7554);
nor U7607 (N_7607,N_7529,N_7536);
xnor U7608 (N_7608,N_7575,N_7534);
nor U7609 (N_7609,N_7596,N_7514);
and U7610 (N_7610,N_7441,N_7459);
xor U7611 (N_7611,N_7455,N_7439);
and U7612 (N_7612,N_7578,N_7559);
nand U7613 (N_7613,N_7445,N_7449);
nor U7614 (N_7614,N_7466,N_7423);
or U7615 (N_7615,N_7507,N_7523);
or U7616 (N_7616,N_7418,N_7509);
and U7617 (N_7617,N_7577,N_7555);
xor U7618 (N_7618,N_7594,N_7457);
or U7619 (N_7619,N_7416,N_7518);
xnor U7620 (N_7620,N_7417,N_7505);
xor U7621 (N_7621,N_7580,N_7598);
and U7622 (N_7622,N_7513,N_7563);
and U7623 (N_7623,N_7428,N_7550);
xor U7624 (N_7624,N_7569,N_7498);
nand U7625 (N_7625,N_7545,N_7508);
nor U7626 (N_7626,N_7444,N_7502);
nor U7627 (N_7627,N_7453,N_7503);
and U7628 (N_7628,N_7404,N_7406);
nor U7629 (N_7629,N_7564,N_7481);
nand U7630 (N_7630,N_7494,N_7561);
and U7631 (N_7631,N_7541,N_7471);
nand U7632 (N_7632,N_7468,N_7442);
and U7633 (N_7633,N_7592,N_7462);
or U7634 (N_7634,N_7512,N_7519);
nor U7635 (N_7635,N_7425,N_7446);
nand U7636 (N_7636,N_7546,N_7422);
or U7637 (N_7637,N_7582,N_7581);
and U7638 (N_7638,N_7448,N_7562);
nor U7639 (N_7639,N_7478,N_7400);
or U7640 (N_7640,N_7405,N_7467);
and U7641 (N_7641,N_7408,N_7576);
xnor U7642 (N_7642,N_7574,N_7530);
nand U7643 (N_7643,N_7486,N_7515);
and U7644 (N_7644,N_7431,N_7407);
nor U7645 (N_7645,N_7590,N_7597);
xnor U7646 (N_7646,N_7589,N_7456);
nor U7647 (N_7647,N_7497,N_7470);
xor U7648 (N_7648,N_7482,N_7566);
and U7649 (N_7649,N_7461,N_7544);
xnor U7650 (N_7650,N_7477,N_7484);
or U7651 (N_7651,N_7480,N_7551);
or U7652 (N_7652,N_7464,N_7510);
nor U7653 (N_7653,N_7553,N_7401);
nor U7654 (N_7654,N_7543,N_7492);
or U7655 (N_7655,N_7473,N_7429);
or U7656 (N_7656,N_7463,N_7495);
nor U7657 (N_7657,N_7474,N_7556);
nand U7658 (N_7658,N_7447,N_7504);
nor U7659 (N_7659,N_7432,N_7465);
nand U7660 (N_7660,N_7565,N_7568);
xor U7661 (N_7661,N_7525,N_7437);
or U7662 (N_7662,N_7526,N_7420);
or U7663 (N_7663,N_7440,N_7522);
nor U7664 (N_7664,N_7532,N_7436);
or U7665 (N_7665,N_7524,N_7488);
and U7666 (N_7666,N_7493,N_7583);
nand U7667 (N_7667,N_7570,N_7511);
and U7668 (N_7668,N_7450,N_7454);
nor U7669 (N_7669,N_7485,N_7595);
xnor U7670 (N_7670,N_7419,N_7421);
and U7671 (N_7671,N_7472,N_7516);
xor U7672 (N_7672,N_7552,N_7560);
nand U7673 (N_7673,N_7538,N_7557);
xnor U7674 (N_7674,N_7540,N_7549);
and U7675 (N_7675,N_7547,N_7535);
xnor U7676 (N_7676,N_7533,N_7501);
nand U7677 (N_7677,N_7483,N_7435);
and U7678 (N_7678,N_7542,N_7586);
xor U7679 (N_7679,N_7411,N_7433);
nor U7680 (N_7680,N_7517,N_7460);
or U7681 (N_7681,N_7506,N_7475);
or U7682 (N_7682,N_7434,N_7599);
nor U7683 (N_7683,N_7438,N_7410);
xor U7684 (N_7684,N_7430,N_7572);
and U7685 (N_7685,N_7527,N_7412);
xor U7686 (N_7686,N_7579,N_7490);
nand U7687 (N_7687,N_7479,N_7520);
nor U7688 (N_7688,N_7593,N_7573);
and U7689 (N_7689,N_7528,N_7499);
nor U7690 (N_7690,N_7458,N_7587);
nor U7691 (N_7691,N_7489,N_7539);
and U7692 (N_7692,N_7548,N_7571);
or U7693 (N_7693,N_7469,N_7427);
nand U7694 (N_7694,N_7476,N_7403);
xor U7695 (N_7695,N_7558,N_7491);
and U7696 (N_7696,N_7424,N_7588);
or U7697 (N_7697,N_7487,N_7496);
or U7698 (N_7698,N_7584,N_7426);
and U7699 (N_7699,N_7451,N_7414);
and U7700 (N_7700,N_7480,N_7541);
nor U7701 (N_7701,N_7486,N_7559);
nor U7702 (N_7702,N_7473,N_7590);
or U7703 (N_7703,N_7432,N_7434);
nand U7704 (N_7704,N_7484,N_7482);
xnor U7705 (N_7705,N_7458,N_7596);
nor U7706 (N_7706,N_7402,N_7418);
nand U7707 (N_7707,N_7413,N_7496);
or U7708 (N_7708,N_7439,N_7597);
or U7709 (N_7709,N_7579,N_7466);
nor U7710 (N_7710,N_7425,N_7507);
nor U7711 (N_7711,N_7482,N_7429);
nand U7712 (N_7712,N_7486,N_7598);
nand U7713 (N_7713,N_7460,N_7467);
nor U7714 (N_7714,N_7444,N_7423);
xor U7715 (N_7715,N_7485,N_7435);
and U7716 (N_7716,N_7519,N_7593);
nand U7717 (N_7717,N_7535,N_7520);
and U7718 (N_7718,N_7596,N_7474);
xor U7719 (N_7719,N_7471,N_7491);
nand U7720 (N_7720,N_7490,N_7551);
xor U7721 (N_7721,N_7576,N_7587);
xnor U7722 (N_7722,N_7496,N_7545);
nor U7723 (N_7723,N_7523,N_7527);
and U7724 (N_7724,N_7555,N_7453);
nor U7725 (N_7725,N_7563,N_7471);
nor U7726 (N_7726,N_7404,N_7458);
nor U7727 (N_7727,N_7445,N_7544);
xnor U7728 (N_7728,N_7431,N_7418);
or U7729 (N_7729,N_7598,N_7474);
or U7730 (N_7730,N_7505,N_7490);
xor U7731 (N_7731,N_7419,N_7571);
or U7732 (N_7732,N_7496,N_7473);
or U7733 (N_7733,N_7493,N_7539);
xnor U7734 (N_7734,N_7429,N_7507);
nor U7735 (N_7735,N_7522,N_7504);
xor U7736 (N_7736,N_7446,N_7488);
xor U7737 (N_7737,N_7458,N_7452);
or U7738 (N_7738,N_7507,N_7446);
and U7739 (N_7739,N_7581,N_7506);
nor U7740 (N_7740,N_7526,N_7413);
and U7741 (N_7741,N_7401,N_7469);
nor U7742 (N_7742,N_7441,N_7466);
xnor U7743 (N_7743,N_7407,N_7439);
nor U7744 (N_7744,N_7507,N_7573);
nand U7745 (N_7745,N_7489,N_7528);
nand U7746 (N_7746,N_7473,N_7449);
or U7747 (N_7747,N_7557,N_7499);
and U7748 (N_7748,N_7537,N_7589);
nor U7749 (N_7749,N_7514,N_7405);
xor U7750 (N_7750,N_7410,N_7427);
nand U7751 (N_7751,N_7557,N_7425);
or U7752 (N_7752,N_7400,N_7463);
and U7753 (N_7753,N_7577,N_7478);
and U7754 (N_7754,N_7418,N_7410);
nand U7755 (N_7755,N_7529,N_7456);
xnor U7756 (N_7756,N_7429,N_7451);
or U7757 (N_7757,N_7587,N_7524);
xor U7758 (N_7758,N_7496,N_7481);
or U7759 (N_7759,N_7532,N_7512);
nand U7760 (N_7760,N_7416,N_7417);
nor U7761 (N_7761,N_7493,N_7401);
nor U7762 (N_7762,N_7433,N_7553);
xnor U7763 (N_7763,N_7552,N_7567);
or U7764 (N_7764,N_7530,N_7422);
and U7765 (N_7765,N_7493,N_7481);
or U7766 (N_7766,N_7492,N_7446);
or U7767 (N_7767,N_7429,N_7498);
nand U7768 (N_7768,N_7554,N_7518);
nor U7769 (N_7769,N_7424,N_7449);
and U7770 (N_7770,N_7480,N_7538);
nor U7771 (N_7771,N_7591,N_7487);
or U7772 (N_7772,N_7549,N_7401);
nand U7773 (N_7773,N_7443,N_7415);
and U7774 (N_7774,N_7498,N_7404);
or U7775 (N_7775,N_7558,N_7413);
xor U7776 (N_7776,N_7567,N_7590);
and U7777 (N_7777,N_7500,N_7415);
nor U7778 (N_7778,N_7535,N_7423);
nand U7779 (N_7779,N_7557,N_7582);
and U7780 (N_7780,N_7578,N_7589);
nor U7781 (N_7781,N_7532,N_7561);
or U7782 (N_7782,N_7492,N_7427);
nand U7783 (N_7783,N_7505,N_7481);
or U7784 (N_7784,N_7493,N_7497);
and U7785 (N_7785,N_7408,N_7596);
or U7786 (N_7786,N_7449,N_7597);
or U7787 (N_7787,N_7576,N_7462);
and U7788 (N_7788,N_7588,N_7460);
or U7789 (N_7789,N_7423,N_7537);
and U7790 (N_7790,N_7438,N_7559);
nand U7791 (N_7791,N_7422,N_7440);
xnor U7792 (N_7792,N_7411,N_7479);
or U7793 (N_7793,N_7482,N_7449);
nand U7794 (N_7794,N_7452,N_7585);
xor U7795 (N_7795,N_7404,N_7489);
nor U7796 (N_7796,N_7570,N_7452);
and U7797 (N_7797,N_7429,N_7436);
nand U7798 (N_7798,N_7475,N_7558);
xnor U7799 (N_7799,N_7511,N_7573);
xor U7800 (N_7800,N_7656,N_7747);
and U7801 (N_7801,N_7787,N_7777);
and U7802 (N_7802,N_7603,N_7616);
nor U7803 (N_7803,N_7760,N_7714);
xnor U7804 (N_7804,N_7732,N_7652);
and U7805 (N_7805,N_7734,N_7717);
and U7806 (N_7806,N_7793,N_7720);
xnor U7807 (N_7807,N_7698,N_7600);
nand U7808 (N_7808,N_7765,N_7790);
or U7809 (N_7809,N_7743,N_7664);
nor U7810 (N_7810,N_7620,N_7709);
and U7811 (N_7811,N_7657,N_7706);
or U7812 (N_7812,N_7677,N_7788);
or U7813 (N_7813,N_7633,N_7613);
or U7814 (N_7814,N_7624,N_7687);
xnor U7815 (N_7815,N_7769,N_7735);
nand U7816 (N_7816,N_7602,N_7666);
and U7817 (N_7817,N_7725,N_7642);
xnor U7818 (N_7818,N_7619,N_7679);
or U7819 (N_7819,N_7766,N_7775);
xnor U7820 (N_7820,N_7625,N_7730);
xor U7821 (N_7821,N_7739,N_7713);
or U7822 (N_7822,N_7688,N_7695);
or U7823 (N_7823,N_7712,N_7693);
xor U7824 (N_7824,N_7637,N_7771);
xnor U7825 (N_7825,N_7722,N_7605);
nand U7826 (N_7826,N_7680,N_7623);
and U7827 (N_7827,N_7697,N_7649);
nand U7828 (N_7828,N_7660,N_7736);
or U7829 (N_7829,N_7753,N_7745);
nor U7830 (N_7830,N_7641,N_7651);
nor U7831 (N_7831,N_7635,N_7715);
xnor U7832 (N_7832,N_7792,N_7797);
nand U7833 (N_7833,N_7675,N_7783);
nor U7834 (N_7834,N_7604,N_7690);
nand U7835 (N_7835,N_7789,N_7681);
and U7836 (N_7836,N_7757,N_7686);
nand U7837 (N_7837,N_7685,N_7670);
nor U7838 (N_7838,N_7723,N_7767);
or U7839 (N_7839,N_7663,N_7683);
or U7840 (N_7840,N_7755,N_7643);
nand U7841 (N_7841,N_7776,N_7778);
nand U7842 (N_7842,N_7606,N_7647);
or U7843 (N_7843,N_7627,N_7768);
nor U7844 (N_7844,N_7726,N_7758);
and U7845 (N_7845,N_7773,N_7785);
nand U7846 (N_7846,N_7678,N_7631);
nand U7847 (N_7847,N_7614,N_7781);
and U7848 (N_7848,N_7655,N_7696);
nor U7849 (N_7849,N_7622,N_7741);
nor U7850 (N_7850,N_7669,N_7774);
and U7851 (N_7851,N_7795,N_7634);
nor U7852 (N_7852,N_7721,N_7615);
nand U7853 (N_7853,N_7692,N_7780);
nand U7854 (N_7854,N_7610,N_7752);
and U7855 (N_7855,N_7798,N_7707);
nand U7856 (N_7856,N_7701,N_7728);
and U7857 (N_7857,N_7650,N_7719);
and U7858 (N_7858,N_7629,N_7645);
xnor U7859 (N_7859,N_7676,N_7756);
nor U7860 (N_7860,N_7628,N_7762);
xor U7861 (N_7861,N_7659,N_7746);
xor U7862 (N_7862,N_7749,N_7748);
nor U7863 (N_7863,N_7742,N_7638);
or U7864 (N_7864,N_7608,N_7729);
nor U7865 (N_7865,N_7761,N_7718);
and U7866 (N_7866,N_7711,N_7626);
nor U7867 (N_7867,N_7617,N_7727);
nor U7868 (N_7868,N_7779,N_7796);
or U7869 (N_7869,N_7764,N_7601);
nand U7870 (N_7870,N_7708,N_7673);
xor U7871 (N_7871,N_7674,N_7733);
nand U7872 (N_7872,N_7754,N_7699);
xor U7873 (N_7873,N_7700,N_7782);
nor U7874 (N_7874,N_7661,N_7731);
nor U7875 (N_7875,N_7646,N_7772);
or U7876 (N_7876,N_7770,N_7716);
xnor U7877 (N_7877,N_7702,N_7704);
or U7878 (N_7878,N_7612,N_7691);
and U7879 (N_7879,N_7607,N_7618);
nand U7880 (N_7880,N_7667,N_7671);
xnor U7881 (N_7881,N_7763,N_7644);
nand U7882 (N_7882,N_7759,N_7654);
nand U7883 (N_7883,N_7738,N_7662);
or U7884 (N_7884,N_7724,N_7630);
nand U7885 (N_7885,N_7640,N_7621);
xor U7886 (N_7886,N_7694,N_7786);
nor U7887 (N_7887,N_7658,N_7794);
xnor U7888 (N_7888,N_7653,N_7740);
xnor U7889 (N_7889,N_7648,N_7705);
xnor U7890 (N_7890,N_7784,N_7632);
nor U7891 (N_7891,N_7672,N_7684);
and U7892 (N_7892,N_7751,N_7611);
nand U7893 (N_7893,N_7737,N_7799);
nor U7894 (N_7894,N_7703,N_7791);
nand U7895 (N_7895,N_7750,N_7609);
nor U7896 (N_7896,N_7710,N_7744);
nand U7897 (N_7897,N_7639,N_7668);
or U7898 (N_7898,N_7682,N_7689);
or U7899 (N_7899,N_7665,N_7636);
nor U7900 (N_7900,N_7658,N_7656);
xnor U7901 (N_7901,N_7652,N_7745);
nor U7902 (N_7902,N_7629,N_7640);
nand U7903 (N_7903,N_7653,N_7703);
nor U7904 (N_7904,N_7650,N_7775);
nand U7905 (N_7905,N_7669,N_7727);
nand U7906 (N_7906,N_7798,N_7721);
nor U7907 (N_7907,N_7602,N_7693);
and U7908 (N_7908,N_7755,N_7709);
xnor U7909 (N_7909,N_7776,N_7656);
nand U7910 (N_7910,N_7663,N_7763);
and U7911 (N_7911,N_7728,N_7697);
nand U7912 (N_7912,N_7706,N_7671);
xor U7913 (N_7913,N_7736,N_7756);
xor U7914 (N_7914,N_7755,N_7741);
nor U7915 (N_7915,N_7798,N_7646);
and U7916 (N_7916,N_7681,N_7645);
and U7917 (N_7917,N_7735,N_7758);
xor U7918 (N_7918,N_7619,N_7645);
nor U7919 (N_7919,N_7635,N_7761);
xnor U7920 (N_7920,N_7713,N_7789);
or U7921 (N_7921,N_7689,N_7787);
nand U7922 (N_7922,N_7759,N_7668);
nand U7923 (N_7923,N_7785,N_7769);
nand U7924 (N_7924,N_7747,N_7671);
nor U7925 (N_7925,N_7785,N_7652);
and U7926 (N_7926,N_7608,N_7623);
nor U7927 (N_7927,N_7710,N_7787);
or U7928 (N_7928,N_7689,N_7760);
and U7929 (N_7929,N_7715,N_7716);
nand U7930 (N_7930,N_7767,N_7665);
xor U7931 (N_7931,N_7639,N_7756);
or U7932 (N_7932,N_7709,N_7676);
nor U7933 (N_7933,N_7791,N_7741);
nor U7934 (N_7934,N_7726,N_7698);
xor U7935 (N_7935,N_7689,N_7680);
and U7936 (N_7936,N_7780,N_7641);
and U7937 (N_7937,N_7788,N_7686);
or U7938 (N_7938,N_7702,N_7671);
or U7939 (N_7939,N_7796,N_7758);
nand U7940 (N_7940,N_7741,N_7770);
nand U7941 (N_7941,N_7620,N_7687);
nor U7942 (N_7942,N_7678,N_7666);
or U7943 (N_7943,N_7777,N_7601);
nand U7944 (N_7944,N_7742,N_7727);
and U7945 (N_7945,N_7724,N_7684);
xor U7946 (N_7946,N_7634,N_7651);
or U7947 (N_7947,N_7706,N_7658);
or U7948 (N_7948,N_7763,N_7719);
nor U7949 (N_7949,N_7700,N_7719);
or U7950 (N_7950,N_7777,N_7718);
or U7951 (N_7951,N_7786,N_7672);
nor U7952 (N_7952,N_7773,N_7685);
or U7953 (N_7953,N_7677,N_7682);
xnor U7954 (N_7954,N_7713,N_7776);
xnor U7955 (N_7955,N_7706,N_7719);
and U7956 (N_7956,N_7659,N_7785);
nand U7957 (N_7957,N_7729,N_7634);
xor U7958 (N_7958,N_7697,N_7735);
nand U7959 (N_7959,N_7780,N_7766);
nor U7960 (N_7960,N_7786,N_7724);
nand U7961 (N_7961,N_7604,N_7719);
nand U7962 (N_7962,N_7637,N_7792);
nor U7963 (N_7963,N_7719,N_7660);
or U7964 (N_7964,N_7625,N_7620);
and U7965 (N_7965,N_7794,N_7783);
and U7966 (N_7966,N_7612,N_7688);
xnor U7967 (N_7967,N_7751,N_7626);
xnor U7968 (N_7968,N_7748,N_7607);
xnor U7969 (N_7969,N_7752,N_7785);
nand U7970 (N_7970,N_7753,N_7608);
nor U7971 (N_7971,N_7648,N_7646);
nor U7972 (N_7972,N_7607,N_7741);
or U7973 (N_7973,N_7623,N_7731);
and U7974 (N_7974,N_7600,N_7756);
nor U7975 (N_7975,N_7738,N_7664);
and U7976 (N_7976,N_7710,N_7725);
and U7977 (N_7977,N_7613,N_7649);
nor U7978 (N_7978,N_7698,N_7742);
or U7979 (N_7979,N_7705,N_7686);
nand U7980 (N_7980,N_7709,N_7750);
or U7981 (N_7981,N_7723,N_7640);
or U7982 (N_7982,N_7774,N_7608);
nand U7983 (N_7983,N_7609,N_7603);
nor U7984 (N_7984,N_7675,N_7686);
nand U7985 (N_7985,N_7680,N_7760);
nor U7986 (N_7986,N_7686,N_7641);
or U7987 (N_7987,N_7699,N_7747);
xnor U7988 (N_7988,N_7712,N_7614);
nor U7989 (N_7989,N_7645,N_7648);
or U7990 (N_7990,N_7775,N_7713);
nand U7991 (N_7991,N_7688,N_7646);
xor U7992 (N_7992,N_7754,N_7677);
or U7993 (N_7993,N_7727,N_7674);
and U7994 (N_7994,N_7769,N_7739);
or U7995 (N_7995,N_7767,N_7601);
xor U7996 (N_7996,N_7779,N_7656);
nand U7997 (N_7997,N_7668,N_7769);
nand U7998 (N_7998,N_7771,N_7768);
or U7999 (N_7999,N_7612,N_7676);
nand U8000 (N_8000,N_7934,N_7954);
xor U8001 (N_8001,N_7864,N_7941);
and U8002 (N_8002,N_7863,N_7952);
and U8003 (N_8003,N_7838,N_7800);
nor U8004 (N_8004,N_7871,N_7873);
or U8005 (N_8005,N_7946,N_7916);
and U8006 (N_8006,N_7982,N_7928);
nor U8007 (N_8007,N_7883,N_7915);
or U8008 (N_8008,N_7936,N_7826);
or U8009 (N_8009,N_7847,N_7819);
nand U8010 (N_8010,N_7833,N_7917);
and U8011 (N_8011,N_7807,N_7905);
and U8012 (N_8012,N_7931,N_7832);
xor U8013 (N_8013,N_7879,N_7966);
nand U8014 (N_8014,N_7805,N_7890);
nand U8015 (N_8015,N_7978,N_7877);
nor U8016 (N_8016,N_7944,N_7835);
and U8017 (N_8017,N_7914,N_7850);
and U8018 (N_8018,N_7866,N_7821);
nand U8019 (N_8019,N_7911,N_7834);
xnor U8020 (N_8020,N_7989,N_7845);
nand U8021 (N_8021,N_7874,N_7906);
xnor U8022 (N_8022,N_7925,N_7912);
nand U8023 (N_8023,N_7910,N_7984);
and U8024 (N_8024,N_7967,N_7932);
nand U8025 (N_8025,N_7960,N_7981);
nand U8026 (N_8026,N_7888,N_7961);
nor U8027 (N_8027,N_7998,N_7843);
and U8028 (N_8028,N_7968,N_7976);
nand U8029 (N_8029,N_7803,N_7842);
nor U8030 (N_8030,N_7970,N_7852);
and U8031 (N_8031,N_7894,N_7959);
nand U8032 (N_8032,N_7898,N_7872);
nor U8033 (N_8033,N_7823,N_7858);
and U8034 (N_8034,N_7973,N_7991);
nand U8035 (N_8035,N_7812,N_7937);
nor U8036 (N_8036,N_7986,N_7861);
or U8037 (N_8037,N_7902,N_7837);
xnor U8038 (N_8038,N_7907,N_7948);
xnor U8039 (N_8039,N_7990,N_7810);
nand U8040 (N_8040,N_7816,N_7900);
or U8041 (N_8041,N_7909,N_7977);
xor U8042 (N_8042,N_7929,N_7997);
nand U8043 (N_8043,N_7891,N_7983);
or U8044 (N_8044,N_7942,N_7862);
nand U8045 (N_8045,N_7945,N_7995);
xor U8046 (N_8046,N_7950,N_7840);
and U8047 (N_8047,N_7848,N_7831);
and U8048 (N_8048,N_7867,N_7924);
nor U8049 (N_8049,N_7822,N_7806);
nor U8050 (N_8050,N_7996,N_7927);
or U8051 (N_8051,N_7811,N_7827);
and U8052 (N_8052,N_7951,N_7940);
or U8053 (N_8053,N_7971,N_7824);
nor U8054 (N_8054,N_7820,N_7884);
and U8055 (N_8055,N_7957,N_7969);
nor U8056 (N_8056,N_7809,N_7895);
nor U8057 (N_8057,N_7887,N_7930);
nor U8058 (N_8058,N_7980,N_7975);
xnor U8059 (N_8059,N_7920,N_7899);
xnor U8060 (N_8060,N_7869,N_7956);
xnor U8061 (N_8061,N_7965,N_7962);
nand U8062 (N_8062,N_7892,N_7904);
nand U8063 (N_8063,N_7938,N_7854);
xnor U8064 (N_8064,N_7829,N_7859);
or U8065 (N_8065,N_7881,N_7886);
nor U8066 (N_8066,N_7801,N_7933);
nor U8067 (N_8067,N_7878,N_7841);
and U8068 (N_8068,N_7919,N_7870);
nand U8069 (N_8069,N_7882,N_7923);
and U8070 (N_8070,N_7918,N_7849);
and U8071 (N_8071,N_7953,N_7813);
nand U8072 (N_8072,N_7943,N_7802);
and U8073 (N_8073,N_7893,N_7855);
and U8074 (N_8074,N_7901,N_7846);
nor U8075 (N_8075,N_7853,N_7851);
nand U8076 (N_8076,N_7828,N_7979);
or U8077 (N_8077,N_7921,N_7885);
nor U8078 (N_8078,N_7939,N_7908);
nor U8079 (N_8079,N_7804,N_7817);
and U8080 (N_8080,N_7857,N_7818);
and U8081 (N_8081,N_7815,N_7880);
nor U8082 (N_8082,N_7865,N_7897);
nor U8083 (N_8083,N_7839,N_7830);
xnor U8084 (N_8084,N_7985,N_7993);
and U8085 (N_8085,N_7987,N_7922);
and U8086 (N_8086,N_7964,N_7963);
nand U8087 (N_8087,N_7808,N_7935);
nor U8088 (N_8088,N_7994,N_7972);
or U8089 (N_8089,N_7949,N_7868);
and U8090 (N_8090,N_7896,N_7926);
xnor U8091 (N_8091,N_7955,N_7903);
or U8092 (N_8092,N_7999,N_7875);
nand U8093 (N_8093,N_7825,N_7836);
or U8094 (N_8094,N_7947,N_7844);
or U8095 (N_8095,N_7974,N_7860);
or U8096 (N_8096,N_7992,N_7988);
or U8097 (N_8097,N_7856,N_7876);
nor U8098 (N_8098,N_7889,N_7958);
nand U8099 (N_8099,N_7814,N_7913);
and U8100 (N_8100,N_7823,N_7953);
nand U8101 (N_8101,N_7964,N_7882);
nor U8102 (N_8102,N_7921,N_7880);
or U8103 (N_8103,N_7891,N_7843);
xnor U8104 (N_8104,N_7930,N_7909);
nand U8105 (N_8105,N_7930,N_7968);
nand U8106 (N_8106,N_7968,N_7959);
nor U8107 (N_8107,N_7830,N_7836);
nand U8108 (N_8108,N_7908,N_7816);
or U8109 (N_8109,N_7883,N_7840);
and U8110 (N_8110,N_7850,N_7939);
and U8111 (N_8111,N_7847,N_7817);
xor U8112 (N_8112,N_7891,N_7874);
or U8113 (N_8113,N_7901,N_7888);
nor U8114 (N_8114,N_7938,N_7932);
and U8115 (N_8115,N_7868,N_7942);
and U8116 (N_8116,N_7958,N_7924);
and U8117 (N_8117,N_7941,N_7885);
nor U8118 (N_8118,N_7847,N_7864);
nor U8119 (N_8119,N_7955,N_7803);
or U8120 (N_8120,N_7830,N_7898);
xor U8121 (N_8121,N_7836,N_7982);
or U8122 (N_8122,N_7848,N_7871);
nor U8123 (N_8123,N_7845,N_7944);
nand U8124 (N_8124,N_7944,N_7820);
xnor U8125 (N_8125,N_7885,N_7856);
nor U8126 (N_8126,N_7984,N_7969);
xnor U8127 (N_8127,N_7882,N_7906);
nand U8128 (N_8128,N_7803,N_7998);
xnor U8129 (N_8129,N_7861,N_7812);
nand U8130 (N_8130,N_7952,N_7843);
nand U8131 (N_8131,N_7937,N_7876);
or U8132 (N_8132,N_7844,N_7807);
nand U8133 (N_8133,N_7808,N_7977);
nand U8134 (N_8134,N_7814,N_7811);
xnor U8135 (N_8135,N_7911,N_7932);
xnor U8136 (N_8136,N_7840,N_7884);
or U8137 (N_8137,N_7889,N_7879);
nand U8138 (N_8138,N_7806,N_7988);
xnor U8139 (N_8139,N_7853,N_7888);
xnor U8140 (N_8140,N_7848,N_7951);
nand U8141 (N_8141,N_7890,N_7822);
nor U8142 (N_8142,N_7977,N_7907);
and U8143 (N_8143,N_7918,N_7873);
nand U8144 (N_8144,N_7877,N_7946);
xnor U8145 (N_8145,N_7806,N_7945);
or U8146 (N_8146,N_7829,N_7949);
xor U8147 (N_8147,N_7840,N_7961);
and U8148 (N_8148,N_7917,N_7877);
or U8149 (N_8149,N_7917,N_7818);
or U8150 (N_8150,N_7987,N_7995);
nand U8151 (N_8151,N_7943,N_7998);
nor U8152 (N_8152,N_7806,N_7858);
xor U8153 (N_8153,N_7929,N_7978);
nor U8154 (N_8154,N_7822,N_7920);
xnor U8155 (N_8155,N_7927,N_7811);
nor U8156 (N_8156,N_7982,N_7813);
nand U8157 (N_8157,N_7810,N_7842);
nand U8158 (N_8158,N_7984,N_7888);
xor U8159 (N_8159,N_7987,N_7806);
xnor U8160 (N_8160,N_7878,N_7860);
and U8161 (N_8161,N_7971,N_7907);
nand U8162 (N_8162,N_7913,N_7945);
and U8163 (N_8163,N_7830,N_7904);
and U8164 (N_8164,N_7818,N_7961);
or U8165 (N_8165,N_7982,N_7867);
nand U8166 (N_8166,N_7947,N_7977);
and U8167 (N_8167,N_7913,N_7904);
and U8168 (N_8168,N_7906,N_7982);
or U8169 (N_8169,N_7934,N_7959);
and U8170 (N_8170,N_7971,N_7811);
and U8171 (N_8171,N_7868,N_7826);
nand U8172 (N_8172,N_7952,N_7983);
nor U8173 (N_8173,N_7999,N_7829);
and U8174 (N_8174,N_7945,N_7922);
nor U8175 (N_8175,N_7920,N_7950);
xnor U8176 (N_8176,N_7850,N_7839);
nand U8177 (N_8177,N_7901,N_7928);
and U8178 (N_8178,N_7850,N_7924);
and U8179 (N_8179,N_7825,N_7971);
nor U8180 (N_8180,N_7920,N_7829);
or U8181 (N_8181,N_7870,N_7849);
or U8182 (N_8182,N_7825,N_7906);
nand U8183 (N_8183,N_7846,N_7881);
or U8184 (N_8184,N_7939,N_7887);
nand U8185 (N_8185,N_7952,N_7847);
or U8186 (N_8186,N_7959,N_7841);
nor U8187 (N_8187,N_7951,N_7894);
nor U8188 (N_8188,N_7979,N_7988);
or U8189 (N_8189,N_7995,N_7998);
or U8190 (N_8190,N_7855,N_7966);
and U8191 (N_8191,N_7977,N_7825);
nor U8192 (N_8192,N_7956,N_7950);
or U8193 (N_8193,N_7891,N_7913);
xnor U8194 (N_8194,N_7983,N_7926);
nor U8195 (N_8195,N_7995,N_7854);
or U8196 (N_8196,N_7889,N_7978);
xor U8197 (N_8197,N_7980,N_7881);
or U8198 (N_8198,N_7880,N_7878);
nand U8199 (N_8199,N_7990,N_7996);
nand U8200 (N_8200,N_8009,N_8160);
nor U8201 (N_8201,N_8034,N_8155);
and U8202 (N_8202,N_8041,N_8044);
or U8203 (N_8203,N_8111,N_8104);
xor U8204 (N_8204,N_8052,N_8136);
or U8205 (N_8205,N_8143,N_8144);
or U8206 (N_8206,N_8140,N_8168);
nor U8207 (N_8207,N_8188,N_8177);
nor U8208 (N_8208,N_8098,N_8071);
nand U8209 (N_8209,N_8054,N_8035);
nor U8210 (N_8210,N_8005,N_8036);
or U8211 (N_8211,N_8102,N_8132);
and U8212 (N_8212,N_8055,N_8003);
xor U8213 (N_8213,N_8158,N_8027);
nand U8214 (N_8214,N_8000,N_8148);
xnor U8215 (N_8215,N_8012,N_8196);
nor U8216 (N_8216,N_8002,N_8150);
nor U8217 (N_8217,N_8045,N_8024);
xor U8218 (N_8218,N_8163,N_8099);
nand U8219 (N_8219,N_8171,N_8047);
and U8220 (N_8220,N_8130,N_8128);
nand U8221 (N_8221,N_8011,N_8161);
nor U8222 (N_8222,N_8170,N_8137);
and U8223 (N_8223,N_8120,N_8029);
nor U8224 (N_8224,N_8076,N_8147);
and U8225 (N_8225,N_8008,N_8017);
nand U8226 (N_8226,N_8058,N_8095);
nand U8227 (N_8227,N_8084,N_8119);
nand U8228 (N_8228,N_8075,N_8097);
nand U8229 (N_8229,N_8125,N_8092);
nand U8230 (N_8230,N_8142,N_8192);
or U8231 (N_8231,N_8162,N_8100);
or U8232 (N_8232,N_8138,N_8069);
nand U8233 (N_8233,N_8073,N_8062);
xnor U8234 (N_8234,N_8060,N_8030);
nor U8235 (N_8235,N_8033,N_8023);
nand U8236 (N_8236,N_8079,N_8172);
nand U8237 (N_8237,N_8061,N_8039);
nor U8238 (N_8238,N_8127,N_8134);
nand U8239 (N_8239,N_8106,N_8078);
or U8240 (N_8240,N_8139,N_8156);
and U8241 (N_8241,N_8022,N_8121);
nor U8242 (N_8242,N_8031,N_8151);
xor U8243 (N_8243,N_8013,N_8080);
nor U8244 (N_8244,N_8059,N_8087);
or U8245 (N_8245,N_8187,N_8146);
and U8246 (N_8246,N_8016,N_8164);
xnor U8247 (N_8247,N_8042,N_8063);
xor U8248 (N_8248,N_8037,N_8107);
nand U8249 (N_8249,N_8105,N_8028);
and U8250 (N_8250,N_8149,N_8174);
nor U8251 (N_8251,N_8032,N_8116);
and U8252 (N_8252,N_8048,N_8064);
or U8253 (N_8253,N_8091,N_8072);
or U8254 (N_8254,N_8198,N_8129);
nor U8255 (N_8255,N_8179,N_8086);
and U8256 (N_8256,N_8083,N_8191);
nand U8257 (N_8257,N_8190,N_8176);
xor U8258 (N_8258,N_8004,N_8185);
nand U8259 (N_8259,N_8123,N_8109);
nor U8260 (N_8260,N_8199,N_8118);
and U8261 (N_8261,N_8089,N_8197);
or U8262 (N_8262,N_8001,N_8068);
or U8263 (N_8263,N_8050,N_8015);
or U8264 (N_8264,N_8154,N_8184);
or U8265 (N_8265,N_8153,N_8193);
and U8266 (N_8266,N_8026,N_8043);
nor U8267 (N_8267,N_8051,N_8018);
and U8268 (N_8268,N_8025,N_8152);
nand U8269 (N_8269,N_8124,N_8175);
nand U8270 (N_8270,N_8145,N_8066);
nand U8271 (N_8271,N_8194,N_8082);
nand U8272 (N_8272,N_8110,N_8096);
nand U8273 (N_8273,N_8114,N_8053);
and U8274 (N_8274,N_8189,N_8049);
nor U8275 (N_8275,N_8126,N_8108);
or U8276 (N_8276,N_8181,N_8157);
or U8277 (N_8277,N_8182,N_8113);
or U8278 (N_8278,N_8085,N_8103);
xnor U8279 (N_8279,N_8115,N_8159);
nor U8280 (N_8280,N_8094,N_8167);
and U8281 (N_8281,N_8117,N_8112);
nand U8282 (N_8282,N_8019,N_8122);
nor U8283 (N_8283,N_8131,N_8169);
and U8284 (N_8284,N_8195,N_8180);
xnor U8285 (N_8285,N_8046,N_8183);
or U8286 (N_8286,N_8038,N_8040);
and U8287 (N_8287,N_8007,N_8077);
and U8288 (N_8288,N_8081,N_8021);
xor U8289 (N_8289,N_8101,N_8088);
nor U8290 (N_8290,N_8173,N_8006);
nor U8291 (N_8291,N_8165,N_8010);
nand U8292 (N_8292,N_8020,N_8186);
xnor U8293 (N_8293,N_8133,N_8141);
nor U8294 (N_8294,N_8166,N_8135);
xnor U8295 (N_8295,N_8070,N_8067);
nor U8296 (N_8296,N_8178,N_8057);
nand U8297 (N_8297,N_8090,N_8056);
xnor U8298 (N_8298,N_8074,N_8093);
xnor U8299 (N_8299,N_8014,N_8065);
nor U8300 (N_8300,N_8089,N_8096);
and U8301 (N_8301,N_8111,N_8135);
nor U8302 (N_8302,N_8164,N_8094);
xor U8303 (N_8303,N_8007,N_8006);
and U8304 (N_8304,N_8073,N_8152);
nand U8305 (N_8305,N_8012,N_8144);
nor U8306 (N_8306,N_8182,N_8027);
xor U8307 (N_8307,N_8001,N_8181);
nand U8308 (N_8308,N_8104,N_8098);
or U8309 (N_8309,N_8100,N_8193);
nand U8310 (N_8310,N_8112,N_8087);
nor U8311 (N_8311,N_8018,N_8073);
or U8312 (N_8312,N_8066,N_8147);
or U8313 (N_8313,N_8125,N_8020);
or U8314 (N_8314,N_8122,N_8033);
nor U8315 (N_8315,N_8182,N_8001);
or U8316 (N_8316,N_8189,N_8013);
xor U8317 (N_8317,N_8161,N_8187);
or U8318 (N_8318,N_8078,N_8036);
xor U8319 (N_8319,N_8114,N_8043);
and U8320 (N_8320,N_8062,N_8038);
nor U8321 (N_8321,N_8172,N_8021);
nand U8322 (N_8322,N_8136,N_8062);
nor U8323 (N_8323,N_8188,N_8174);
or U8324 (N_8324,N_8013,N_8059);
and U8325 (N_8325,N_8057,N_8073);
xnor U8326 (N_8326,N_8145,N_8040);
or U8327 (N_8327,N_8075,N_8052);
and U8328 (N_8328,N_8087,N_8027);
or U8329 (N_8329,N_8168,N_8154);
nand U8330 (N_8330,N_8068,N_8022);
nor U8331 (N_8331,N_8083,N_8185);
nor U8332 (N_8332,N_8167,N_8123);
nand U8333 (N_8333,N_8087,N_8085);
and U8334 (N_8334,N_8006,N_8012);
and U8335 (N_8335,N_8175,N_8039);
or U8336 (N_8336,N_8087,N_8188);
xor U8337 (N_8337,N_8047,N_8055);
or U8338 (N_8338,N_8189,N_8128);
xor U8339 (N_8339,N_8182,N_8035);
or U8340 (N_8340,N_8078,N_8151);
nor U8341 (N_8341,N_8092,N_8066);
nor U8342 (N_8342,N_8180,N_8079);
xnor U8343 (N_8343,N_8036,N_8153);
nand U8344 (N_8344,N_8016,N_8168);
nor U8345 (N_8345,N_8194,N_8128);
nand U8346 (N_8346,N_8069,N_8001);
or U8347 (N_8347,N_8170,N_8103);
or U8348 (N_8348,N_8179,N_8070);
xor U8349 (N_8349,N_8129,N_8128);
or U8350 (N_8350,N_8186,N_8197);
or U8351 (N_8351,N_8006,N_8172);
nand U8352 (N_8352,N_8123,N_8099);
or U8353 (N_8353,N_8001,N_8085);
nand U8354 (N_8354,N_8014,N_8006);
xnor U8355 (N_8355,N_8075,N_8003);
nand U8356 (N_8356,N_8002,N_8034);
nand U8357 (N_8357,N_8003,N_8123);
xor U8358 (N_8358,N_8018,N_8099);
nor U8359 (N_8359,N_8075,N_8180);
xor U8360 (N_8360,N_8084,N_8192);
nand U8361 (N_8361,N_8158,N_8032);
or U8362 (N_8362,N_8187,N_8062);
nand U8363 (N_8363,N_8190,N_8001);
xnor U8364 (N_8364,N_8003,N_8186);
xor U8365 (N_8365,N_8168,N_8033);
nor U8366 (N_8366,N_8028,N_8146);
or U8367 (N_8367,N_8004,N_8115);
nor U8368 (N_8368,N_8157,N_8001);
or U8369 (N_8369,N_8099,N_8167);
or U8370 (N_8370,N_8047,N_8088);
and U8371 (N_8371,N_8096,N_8152);
and U8372 (N_8372,N_8165,N_8061);
or U8373 (N_8373,N_8174,N_8002);
xor U8374 (N_8374,N_8135,N_8160);
and U8375 (N_8375,N_8012,N_8182);
or U8376 (N_8376,N_8040,N_8039);
or U8377 (N_8377,N_8136,N_8032);
and U8378 (N_8378,N_8174,N_8014);
nand U8379 (N_8379,N_8168,N_8122);
and U8380 (N_8380,N_8036,N_8173);
nor U8381 (N_8381,N_8063,N_8046);
and U8382 (N_8382,N_8124,N_8037);
nand U8383 (N_8383,N_8146,N_8148);
or U8384 (N_8384,N_8006,N_8080);
xnor U8385 (N_8385,N_8171,N_8196);
and U8386 (N_8386,N_8143,N_8191);
and U8387 (N_8387,N_8009,N_8174);
nor U8388 (N_8388,N_8146,N_8002);
nor U8389 (N_8389,N_8026,N_8094);
or U8390 (N_8390,N_8143,N_8102);
nand U8391 (N_8391,N_8086,N_8009);
or U8392 (N_8392,N_8058,N_8059);
and U8393 (N_8393,N_8038,N_8155);
nand U8394 (N_8394,N_8102,N_8176);
nand U8395 (N_8395,N_8150,N_8089);
xor U8396 (N_8396,N_8086,N_8033);
and U8397 (N_8397,N_8048,N_8191);
xor U8398 (N_8398,N_8185,N_8157);
nand U8399 (N_8399,N_8078,N_8152);
xnor U8400 (N_8400,N_8229,N_8371);
xnor U8401 (N_8401,N_8227,N_8205);
and U8402 (N_8402,N_8266,N_8231);
xnor U8403 (N_8403,N_8260,N_8379);
xnor U8404 (N_8404,N_8233,N_8254);
xnor U8405 (N_8405,N_8362,N_8359);
nand U8406 (N_8406,N_8238,N_8208);
nor U8407 (N_8407,N_8226,N_8324);
nand U8408 (N_8408,N_8304,N_8329);
nand U8409 (N_8409,N_8396,N_8340);
and U8410 (N_8410,N_8213,N_8302);
or U8411 (N_8411,N_8272,N_8357);
and U8412 (N_8412,N_8292,N_8350);
nand U8413 (N_8413,N_8349,N_8286);
nor U8414 (N_8414,N_8248,N_8259);
xor U8415 (N_8415,N_8210,N_8202);
nand U8416 (N_8416,N_8337,N_8322);
or U8417 (N_8417,N_8207,N_8335);
xnor U8418 (N_8418,N_8280,N_8200);
nor U8419 (N_8419,N_8391,N_8386);
and U8420 (N_8420,N_8318,N_8282);
and U8421 (N_8421,N_8287,N_8263);
and U8422 (N_8422,N_8255,N_8392);
nor U8423 (N_8423,N_8369,N_8323);
xor U8424 (N_8424,N_8378,N_8373);
and U8425 (N_8425,N_8290,N_8399);
nand U8426 (N_8426,N_8261,N_8251);
xor U8427 (N_8427,N_8288,N_8285);
or U8428 (N_8428,N_8334,N_8345);
or U8429 (N_8429,N_8281,N_8367);
nor U8430 (N_8430,N_8348,N_8247);
or U8431 (N_8431,N_8344,N_8232);
and U8432 (N_8432,N_8388,N_8295);
nor U8433 (N_8433,N_8310,N_8242);
xor U8434 (N_8434,N_8253,N_8385);
nand U8435 (N_8435,N_8228,N_8355);
or U8436 (N_8436,N_8377,N_8339);
and U8437 (N_8437,N_8315,N_8278);
xor U8438 (N_8438,N_8244,N_8271);
and U8439 (N_8439,N_8296,N_8375);
nor U8440 (N_8440,N_8245,N_8330);
xnor U8441 (N_8441,N_8219,N_8372);
nor U8442 (N_8442,N_8390,N_8241);
nand U8443 (N_8443,N_8343,N_8217);
xnor U8444 (N_8444,N_8393,N_8230);
nor U8445 (N_8445,N_8294,N_8269);
or U8446 (N_8446,N_8325,N_8332);
and U8447 (N_8447,N_8289,N_8262);
and U8448 (N_8448,N_8270,N_8387);
and U8449 (N_8449,N_8316,N_8328);
nand U8450 (N_8450,N_8358,N_8374);
nand U8451 (N_8451,N_8353,N_8333);
and U8452 (N_8452,N_8303,N_8300);
nor U8453 (N_8453,N_8311,N_8309);
or U8454 (N_8454,N_8267,N_8236);
nand U8455 (N_8455,N_8275,N_8249);
xnor U8456 (N_8456,N_8346,N_8243);
nand U8457 (N_8457,N_8257,N_8203);
xor U8458 (N_8458,N_8368,N_8212);
nand U8459 (N_8459,N_8265,N_8327);
or U8460 (N_8460,N_8331,N_8273);
nor U8461 (N_8461,N_8321,N_8308);
and U8462 (N_8462,N_8234,N_8341);
nor U8463 (N_8463,N_8305,N_8398);
nand U8464 (N_8464,N_8363,N_8313);
or U8465 (N_8465,N_8376,N_8264);
xor U8466 (N_8466,N_8380,N_8209);
and U8467 (N_8467,N_8366,N_8220);
and U8468 (N_8468,N_8240,N_8314);
nand U8469 (N_8469,N_8383,N_8215);
and U8470 (N_8470,N_8206,N_8307);
nand U8471 (N_8471,N_8365,N_8291);
nor U8472 (N_8472,N_8252,N_8395);
and U8473 (N_8473,N_8283,N_8336);
nor U8474 (N_8474,N_8319,N_8394);
nand U8475 (N_8475,N_8360,N_8223);
and U8476 (N_8476,N_8312,N_8320);
nand U8477 (N_8477,N_8284,N_8246);
nand U8478 (N_8478,N_8381,N_8301);
nor U8479 (N_8479,N_8258,N_8298);
nand U8480 (N_8480,N_8224,N_8382);
and U8481 (N_8481,N_8352,N_8277);
or U8482 (N_8482,N_8221,N_8211);
or U8483 (N_8483,N_8347,N_8297);
and U8484 (N_8484,N_8239,N_8361);
and U8485 (N_8485,N_8204,N_8235);
nor U8486 (N_8486,N_8384,N_8256);
xnor U8487 (N_8487,N_8354,N_8299);
xnor U8488 (N_8488,N_8370,N_8364);
nand U8489 (N_8489,N_8250,N_8293);
nor U8490 (N_8490,N_8216,N_8389);
nor U8491 (N_8491,N_8201,N_8274);
or U8492 (N_8492,N_8351,N_8317);
and U8493 (N_8493,N_8222,N_8237);
nand U8494 (N_8494,N_8268,N_8342);
nor U8495 (N_8495,N_8218,N_8326);
and U8496 (N_8496,N_8306,N_8214);
nor U8497 (N_8497,N_8279,N_8225);
nor U8498 (N_8498,N_8397,N_8356);
nor U8499 (N_8499,N_8338,N_8276);
xor U8500 (N_8500,N_8280,N_8300);
and U8501 (N_8501,N_8281,N_8220);
or U8502 (N_8502,N_8383,N_8232);
nand U8503 (N_8503,N_8349,N_8351);
nor U8504 (N_8504,N_8255,N_8201);
nor U8505 (N_8505,N_8329,N_8221);
or U8506 (N_8506,N_8323,N_8346);
xnor U8507 (N_8507,N_8380,N_8292);
and U8508 (N_8508,N_8303,N_8261);
and U8509 (N_8509,N_8261,N_8355);
nor U8510 (N_8510,N_8375,N_8292);
nor U8511 (N_8511,N_8275,N_8279);
nor U8512 (N_8512,N_8228,N_8373);
and U8513 (N_8513,N_8257,N_8212);
nor U8514 (N_8514,N_8210,N_8288);
and U8515 (N_8515,N_8231,N_8313);
xor U8516 (N_8516,N_8388,N_8293);
or U8517 (N_8517,N_8210,N_8234);
or U8518 (N_8518,N_8309,N_8351);
or U8519 (N_8519,N_8231,N_8348);
or U8520 (N_8520,N_8238,N_8271);
and U8521 (N_8521,N_8245,N_8241);
nor U8522 (N_8522,N_8210,N_8299);
xnor U8523 (N_8523,N_8358,N_8269);
nor U8524 (N_8524,N_8295,N_8229);
nand U8525 (N_8525,N_8202,N_8245);
nand U8526 (N_8526,N_8398,N_8333);
nor U8527 (N_8527,N_8268,N_8275);
or U8528 (N_8528,N_8270,N_8259);
and U8529 (N_8529,N_8242,N_8314);
xor U8530 (N_8530,N_8315,N_8398);
xnor U8531 (N_8531,N_8239,N_8290);
nand U8532 (N_8532,N_8325,N_8246);
xor U8533 (N_8533,N_8341,N_8319);
or U8534 (N_8534,N_8345,N_8208);
and U8535 (N_8535,N_8343,N_8255);
nor U8536 (N_8536,N_8240,N_8322);
and U8537 (N_8537,N_8362,N_8246);
nand U8538 (N_8538,N_8239,N_8389);
nor U8539 (N_8539,N_8289,N_8381);
xor U8540 (N_8540,N_8214,N_8380);
xnor U8541 (N_8541,N_8297,N_8328);
nand U8542 (N_8542,N_8345,N_8386);
and U8543 (N_8543,N_8332,N_8245);
and U8544 (N_8544,N_8301,N_8210);
xnor U8545 (N_8545,N_8221,N_8270);
nand U8546 (N_8546,N_8252,N_8243);
nor U8547 (N_8547,N_8318,N_8267);
xnor U8548 (N_8548,N_8225,N_8222);
nor U8549 (N_8549,N_8351,N_8259);
xnor U8550 (N_8550,N_8370,N_8210);
or U8551 (N_8551,N_8380,N_8347);
nand U8552 (N_8552,N_8364,N_8316);
and U8553 (N_8553,N_8304,N_8395);
xnor U8554 (N_8554,N_8374,N_8373);
and U8555 (N_8555,N_8237,N_8302);
or U8556 (N_8556,N_8279,N_8361);
nand U8557 (N_8557,N_8375,N_8379);
and U8558 (N_8558,N_8310,N_8396);
nand U8559 (N_8559,N_8210,N_8330);
or U8560 (N_8560,N_8263,N_8320);
nor U8561 (N_8561,N_8365,N_8375);
and U8562 (N_8562,N_8240,N_8287);
xor U8563 (N_8563,N_8321,N_8201);
nand U8564 (N_8564,N_8284,N_8277);
xor U8565 (N_8565,N_8272,N_8313);
nand U8566 (N_8566,N_8248,N_8215);
xor U8567 (N_8567,N_8362,N_8317);
nor U8568 (N_8568,N_8375,N_8264);
or U8569 (N_8569,N_8381,N_8219);
nor U8570 (N_8570,N_8242,N_8286);
xor U8571 (N_8571,N_8379,N_8215);
nor U8572 (N_8572,N_8217,N_8262);
nor U8573 (N_8573,N_8219,N_8306);
nand U8574 (N_8574,N_8309,N_8231);
nand U8575 (N_8575,N_8399,N_8391);
or U8576 (N_8576,N_8299,N_8270);
xor U8577 (N_8577,N_8361,N_8280);
and U8578 (N_8578,N_8329,N_8349);
and U8579 (N_8579,N_8395,N_8384);
nor U8580 (N_8580,N_8257,N_8292);
nor U8581 (N_8581,N_8383,N_8384);
nand U8582 (N_8582,N_8320,N_8308);
xor U8583 (N_8583,N_8227,N_8291);
or U8584 (N_8584,N_8370,N_8300);
and U8585 (N_8585,N_8242,N_8381);
and U8586 (N_8586,N_8233,N_8244);
or U8587 (N_8587,N_8328,N_8218);
nand U8588 (N_8588,N_8336,N_8378);
and U8589 (N_8589,N_8327,N_8381);
or U8590 (N_8590,N_8218,N_8237);
xor U8591 (N_8591,N_8316,N_8266);
and U8592 (N_8592,N_8269,N_8324);
nor U8593 (N_8593,N_8394,N_8213);
or U8594 (N_8594,N_8228,N_8302);
and U8595 (N_8595,N_8277,N_8332);
nand U8596 (N_8596,N_8319,N_8255);
xnor U8597 (N_8597,N_8243,N_8309);
nor U8598 (N_8598,N_8338,N_8232);
xor U8599 (N_8599,N_8200,N_8263);
and U8600 (N_8600,N_8516,N_8478);
nor U8601 (N_8601,N_8472,N_8452);
and U8602 (N_8602,N_8495,N_8488);
xor U8603 (N_8603,N_8431,N_8499);
or U8604 (N_8604,N_8446,N_8465);
or U8605 (N_8605,N_8423,N_8419);
xnor U8606 (N_8606,N_8401,N_8480);
and U8607 (N_8607,N_8595,N_8521);
nand U8608 (N_8608,N_8556,N_8537);
and U8609 (N_8609,N_8425,N_8591);
and U8610 (N_8610,N_8466,N_8507);
xor U8611 (N_8611,N_8572,N_8497);
nor U8612 (N_8612,N_8503,N_8443);
xor U8613 (N_8613,N_8586,N_8546);
xnor U8614 (N_8614,N_8485,N_8405);
xor U8615 (N_8615,N_8592,N_8531);
and U8616 (N_8616,N_8581,N_8417);
xnor U8617 (N_8617,N_8512,N_8477);
nor U8618 (N_8618,N_8469,N_8434);
nand U8619 (N_8619,N_8534,N_8454);
nand U8620 (N_8620,N_8501,N_8471);
or U8621 (N_8621,N_8448,N_8492);
nand U8622 (N_8622,N_8447,N_8553);
nor U8623 (N_8623,N_8463,N_8475);
or U8624 (N_8624,N_8456,N_8580);
xor U8625 (N_8625,N_8544,N_8440);
xor U8626 (N_8626,N_8530,N_8517);
nand U8627 (N_8627,N_8514,N_8506);
nand U8628 (N_8628,N_8467,N_8543);
nor U8629 (N_8629,N_8594,N_8576);
and U8630 (N_8630,N_8528,N_8540);
nand U8631 (N_8631,N_8413,N_8461);
nor U8632 (N_8632,N_8569,N_8420);
or U8633 (N_8633,N_8529,N_8428);
nand U8634 (N_8634,N_8498,N_8402);
nor U8635 (N_8635,N_8574,N_8504);
nand U8636 (N_8636,N_8589,N_8438);
xnor U8637 (N_8637,N_8460,N_8563);
xnor U8638 (N_8638,N_8435,N_8411);
or U8639 (N_8639,N_8583,N_8483);
nand U8640 (N_8640,N_8552,N_8415);
and U8641 (N_8641,N_8468,N_8545);
nand U8642 (N_8642,N_8515,N_8558);
nor U8643 (N_8643,N_8513,N_8484);
xor U8644 (N_8644,N_8481,N_8532);
or U8645 (N_8645,N_8500,N_8561);
nand U8646 (N_8646,N_8567,N_8453);
nor U8647 (N_8647,N_8432,N_8464);
or U8648 (N_8648,N_8442,N_8598);
nand U8649 (N_8649,N_8439,N_8430);
nor U8650 (N_8650,N_8455,N_8409);
nor U8651 (N_8651,N_8496,N_8457);
nor U8652 (N_8652,N_8587,N_8489);
nand U8653 (N_8653,N_8565,N_8575);
and U8654 (N_8654,N_8406,N_8422);
or U8655 (N_8655,N_8538,N_8547);
nand U8656 (N_8656,N_8527,N_8570);
and U8657 (N_8657,N_8510,N_8427);
nand U8658 (N_8658,N_8559,N_8493);
or U8659 (N_8659,N_8424,N_8400);
or U8660 (N_8660,N_8541,N_8548);
nand U8661 (N_8661,N_8535,N_8444);
nor U8662 (N_8662,N_8542,N_8491);
or U8663 (N_8663,N_8584,N_8519);
xor U8664 (N_8664,N_8571,N_8482);
or U8665 (N_8665,N_8437,N_8486);
or U8666 (N_8666,N_8593,N_8459);
or U8667 (N_8667,N_8523,N_8585);
nor U8668 (N_8668,N_8550,N_8509);
or U8669 (N_8669,N_8410,N_8597);
or U8670 (N_8670,N_8533,N_8579);
nor U8671 (N_8671,N_8414,N_8450);
nand U8672 (N_8672,N_8577,N_8408);
or U8673 (N_8673,N_8557,N_8458);
nor U8674 (N_8674,N_8564,N_8596);
xnor U8675 (N_8675,N_8421,N_8573);
or U8676 (N_8676,N_8588,N_8433);
nor U8677 (N_8677,N_8490,N_8518);
or U8678 (N_8678,N_8555,N_8462);
and U8679 (N_8679,N_8474,N_8407);
xnor U8680 (N_8680,N_8520,N_8539);
xnor U8681 (N_8681,N_8599,N_8526);
and U8682 (N_8682,N_8429,N_8426);
or U8683 (N_8683,N_8404,N_8582);
xnor U8684 (N_8684,N_8502,N_8554);
xor U8685 (N_8685,N_8590,N_8470);
nor U8686 (N_8686,N_8473,N_8505);
and U8687 (N_8687,N_8525,N_8562);
nor U8688 (N_8688,N_8536,N_8479);
nand U8689 (N_8689,N_8451,N_8487);
or U8690 (N_8690,N_8578,N_8445);
xor U8691 (N_8691,N_8403,N_8568);
or U8692 (N_8692,N_8441,N_8449);
and U8693 (N_8693,N_8508,N_8511);
or U8694 (N_8694,N_8436,N_8476);
or U8695 (N_8695,N_8549,N_8560);
xnor U8696 (N_8696,N_8418,N_8494);
or U8697 (N_8697,N_8566,N_8551);
xnor U8698 (N_8698,N_8524,N_8522);
or U8699 (N_8699,N_8412,N_8416);
xnor U8700 (N_8700,N_8471,N_8569);
xnor U8701 (N_8701,N_8420,N_8465);
or U8702 (N_8702,N_8535,N_8590);
and U8703 (N_8703,N_8533,N_8564);
xor U8704 (N_8704,N_8571,N_8526);
or U8705 (N_8705,N_8480,N_8532);
or U8706 (N_8706,N_8487,N_8573);
or U8707 (N_8707,N_8556,N_8532);
xor U8708 (N_8708,N_8465,N_8480);
and U8709 (N_8709,N_8582,N_8597);
and U8710 (N_8710,N_8409,N_8502);
nor U8711 (N_8711,N_8424,N_8428);
nor U8712 (N_8712,N_8433,N_8422);
or U8713 (N_8713,N_8448,N_8534);
nand U8714 (N_8714,N_8453,N_8487);
and U8715 (N_8715,N_8514,N_8576);
nand U8716 (N_8716,N_8569,N_8461);
and U8717 (N_8717,N_8434,N_8436);
and U8718 (N_8718,N_8539,N_8436);
or U8719 (N_8719,N_8522,N_8511);
nand U8720 (N_8720,N_8483,N_8444);
nor U8721 (N_8721,N_8529,N_8412);
nor U8722 (N_8722,N_8426,N_8470);
nand U8723 (N_8723,N_8453,N_8583);
or U8724 (N_8724,N_8411,N_8431);
nand U8725 (N_8725,N_8564,N_8417);
or U8726 (N_8726,N_8440,N_8425);
nor U8727 (N_8727,N_8517,N_8541);
or U8728 (N_8728,N_8553,N_8506);
xor U8729 (N_8729,N_8420,N_8417);
nand U8730 (N_8730,N_8502,N_8466);
or U8731 (N_8731,N_8429,N_8473);
xnor U8732 (N_8732,N_8458,N_8485);
xor U8733 (N_8733,N_8569,N_8473);
xor U8734 (N_8734,N_8577,N_8505);
xor U8735 (N_8735,N_8479,N_8424);
xnor U8736 (N_8736,N_8538,N_8574);
nand U8737 (N_8737,N_8514,N_8475);
nand U8738 (N_8738,N_8413,N_8550);
nor U8739 (N_8739,N_8441,N_8422);
nor U8740 (N_8740,N_8494,N_8413);
nor U8741 (N_8741,N_8458,N_8472);
xor U8742 (N_8742,N_8478,N_8446);
or U8743 (N_8743,N_8507,N_8569);
nand U8744 (N_8744,N_8436,N_8506);
nor U8745 (N_8745,N_8593,N_8469);
xnor U8746 (N_8746,N_8407,N_8423);
xnor U8747 (N_8747,N_8514,N_8512);
and U8748 (N_8748,N_8471,N_8485);
xnor U8749 (N_8749,N_8515,N_8564);
xor U8750 (N_8750,N_8560,N_8559);
xor U8751 (N_8751,N_8598,N_8458);
or U8752 (N_8752,N_8487,N_8588);
xor U8753 (N_8753,N_8580,N_8449);
nand U8754 (N_8754,N_8566,N_8530);
nor U8755 (N_8755,N_8542,N_8552);
nor U8756 (N_8756,N_8472,N_8423);
and U8757 (N_8757,N_8438,N_8403);
nand U8758 (N_8758,N_8476,N_8557);
or U8759 (N_8759,N_8533,N_8476);
or U8760 (N_8760,N_8521,N_8570);
nand U8761 (N_8761,N_8574,N_8484);
and U8762 (N_8762,N_8521,N_8403);
nor U8763 (N_8763,N_8446,N_8445);
nor U8764 (N_8764,N_8557,N_8460);
nand U8765 (N_8765,N_8510,N_8483);
or U8766 (N_8766,N_8599,N_8460);
xnor U8767 (N_8767,N_8553,N_8492);
or U8768 (N_8768,N_8458,N_8586);
or U8769 (N_8769,N_8490,N_8574);
nor U8770 (N_8770,N_8539,N_8550);
and U8771 (N_8771,N_8529,N_8491);
nor U8772 (N_8772,N_8563,N_8465);
xor U8773 (N_8773,N_8484,N_8549);
or U8774 (N_8774,N_8463,N_8557);
or U8775 (N_8775,N_8405,N_8585);
xnor U8776 (N_8776,N_8485,N_8550);
nor U8777 (N_8777,N_8489,N_8548);
and U8778 (N_8778,N_8529,N_8465);
nand U8779 (N_8779,N_8580,N_8405);
nand U8780 (N_8780,N_8525,N_8588);
nand U8781 (N_8781,N_8549,N_8405);
nor U8782 (N_8782,N_8418,N_8468);
xor U8783 (N_8783,N_8518,N_8525);
xnor U8784 (N_8784,N_8470,N_8536);
xor U8785 (N_8785,N_8404,N_8457);
xnor U8786 (N_8786,N_8470,N_8427);
or U8787 (N_8787,N_8519,N_8530);
nor U8788 (N_8788,N_8402,N_8532);
xor U8789 (N_8789,N_8565,N_8400);
or U8790 (N_8790,N_8414,N_8453);
nand U8791 (N_8791,N_8576,N_8401);
and U8792 (N_8792,N_8437,N_8568);
or U8793 (N_8793,N_8538,N_8490);
nor U8794 (N_8794,N_8537,N_8521);
and U8795 (N_8795,N_8446,N_8544);
or U8796 (N_8796,N_8583,N_8411);
or U8797 (N_8797,N_8482,N_8551);
and U8798 (N_8798,N_8501,N_8526);
nor U8799 (N_8799,N_8431,N_8500);
and U8800 (N_8800,N_8638,N_8621);
nand U8801 (N_8801,N_8639,N_8791);
xor U8802 (N_8802,N_8793,N_8698);
nand U8803 (N_8803,N_8644,N_8661);
xor U8804 (N_8804,N_8646,N_8751);
and U8805 (N_8805,N_8641,N_8756);
xor U8806 (N_8806,N_8789,N_8712);
and U8807 (N_8807,N_8697,N_8777);
nand U8808 (N_8808,N_8784,N_8630);
nand U8809 (N_8809,N_8671,N_8734);
nand U8810 (N_8810,N_8695,N_8796);
nand U8811 (N_8811,N_8652,N_8729);
or U8812 (N_8812,N_8653,N_8607);
nor U8813 (N_8813,N_8669,N_8799);
xor U8814 (N_8814,N_8662,N_8676);
xnor U8815 (N_8815,N_8675,N_8629);
nor U8816 (N_8816,N_8634,N_8717);
nor U8817 (N_8817,N_8622,N_8776);
xor U8818 (N_8818,N_8680,N_8700);
and U8819 (N_8819,N_8772,N_8725);
nand U8820 (N_8820,N_8797,N_8612);
xnor U8821 (N_8821,N_8672,N_8625);
or U8822 (N_8822,N_8670,N_8703);
or U8823 (N_8823,N_8620,N_8699);
or U8824 (N_8824,N_8614,N_8771);
xnor U8825 (N_8825,N_8651,N_8754);
xor U8826 (N_8826,N_8761,N_8632);
xor U8827 (N_8827,N_8748,N_8604);
or U8828 (N_8828,N_8782,N_8721);
nor U8829 (N_8829,N_8613,N_8688);
nand U8830 (N_8830,N_8633,N_8763);
xnor U8831 (N_8831,N_8687,N_8684);
nand U8832 (N_8832,N_8656,N_8753);
nand U8833 (N_8833,N_8724,N_8606);
xor U8834 (N_8834,N_8664,N_8765);
nor U8835 (N_8835,N_8668,N_8611);
nand U8836 (N_8836,N_8677,N_8738);
nand U8837 (N_8837,N_8663,N_8655);
and U8838 (N_8838,N_8790,N_8746);
nand U8839 (N_8839,N_8658,N_8720);
or U8840 (N_8840,N_8723,N_8786);
or U8841 (N_8841,N_8750,N_8624);
nor U8842 (N_8842,N_8716,N_8749);
or U8843 (N_8843,N_8649,N_8673);
and U8844 (N_8844,N_8742,N_8602);
nor U8845 (N_8845,N_8645,N_8757);
xnor U8846 (N_8846,N_8618,N_8783);
and U8847 (N_8847,N_8706,N_8628);
or U8848 (N_8848,N_8713,N_8615);
and U8849 (N_8849,N_8758,N_8735);
or U8850 (N_8850,N_8635,N_8681);
nor U8851 (N_8851,N_8798,N_8623);
and U8852 (N_8852,N_8619,N_8631);
xor U8853 (N_8853,N_8601,N_8650);
nor U8854 (N_8854,N_8701,N_8794);
nor U8855 (N_8855,N_8636,N_8605);
xnor U8856 (N_8856,N_8743,N_8747);
and U8857 (N_8857,N_8792,N_8730);
and U8858 (N_8858,N_8707,N_8696);
or U8859 (N_8859,N_8767,N_8704);
or U8860 (N_8860,N_8764,N_8710);
xnor U8861 (N_8861,N_8711,N_8667);
nand U8862 (N_8862,N_8626,N_8637);
nor U8863 (N_8863,N_8768,N_8693);
nand U8864 (N_8864,N_8691,N_8654);
nor U8865 (N_8865,N_8708,N_8692);
xnor U8866 (N_8866,N_8719,N_8773);
nor U8867 (N_8867,N_8739,N_8787);
xnor U8868 (N_8868,N_8740,N_8705);
nor U8869 (N_8869,N_8745,N_8627);
and U8870 (N_8870,N_8659,N_8733);
xnor U8871 (N_8871,N_8788,N_8769);
nand U8872 (N_8872,N_8647,N_8648);
nor U8873 (N_8873,N_8690,N_8694);
and U8874 (N_8874,N_8674,N_8741);
and U8875 (N_8875,N_8744,N_8603);
nor U8876 (N_8876,N_8617,N_8755);
nand U8877 (N_8877,N_8774,N_8731);
nor U8878 (N_8878,N_8685,N_8775);
xor U8879 (N_8879,N_8683,N_8795);
nand U8880 (N_8880,N_8616,N_8781);
nand U8881 (N_8881,N_8665,N_8714);
and U8882 (N_8882,N_8760,N_8642);
nand U8883 (N_8883,N_8679,N_8766);
nand U8884 (N_8884,N_8689,N_8779);
xnor U8885 (N_8885,N_8732,N_8759);
xor U8886 (N_8886,N_8678,N_8718);
nand U8887 (N_8887,N_8715,N_8660);
xnor U8888 (N_8888,N_8722,N_8709);
or U8889 (N_8889,N_8643,N_8778);
and U8890 (N_8890,N_8682,N_8727);
and U8891 (N_8891,N_8728,N_8610);
xor U8892 (N_8892,N_8686,N_8726);
or U8893 (N_8893,N_8736,N_8785);
nor U8894 (N_8894,N_8600,N_8666);
xnor U8895 (N_8895,N_8762,N_8609);
xor U8896 (N_8896,N_8657,N_8702);
nand U8897 (N_8897,N_8780,N_8608);
nor U8898 (N_8898,N_8737,N_8640);
or U8899 (N_8899,N_8752,N_8770);
xnor U8900 (N_8900,N_8762,N_8656);
nand U8901 (N_8901,N_8778,N_8688);
and U8902 (N_8902,N_8740,N_8764);
nor U8903 (N_8903,N_8626,N_8765);
nor U8904 (N_8904,N_8752,N_8665);
nor U8905 (N_8905,N_8631,N_8755);
nand U8906 (N_8906,N_8718,N_8753);
or U8907 (N_8907,N_8650,N_8758);
nand U8908 (N_8908,N_8613,N_8699);
or U8909 (N_8909,N_8689,N_8707);
and U8910 (N_8910,N_8704,N_8694);
and U8911 (N_8911,N_8700,N_8772);
xor U8912 (N_8912,N_8672,N_8718);
or U8913 (N_8913,N_8663,N_8797);
and U8914 (N_8914,N_8646,N_8632);
xnor U8915 (N_8915,N_8696,N_8617);
or U8916 (N_8916,N_8699,N_8658);
and U8917 (N_8917,N_8737,N_8739);
and U8918 (N_8918,N_8676,N_8790);
nand U8919 (N_8919,N_8601,N_8764);
xnor U8920 (N_8920,N_8750,N_8751);
nor U8921 (N_8921,N_8731,N_8756);
or U8922 (N_8922,N_8670,N_8625);
xnor U8923 (N_8923,N_8669,N_8723);
and U8924 (N_8924,N_8679,N_8629);
nand U8925 (N_8925,N_8780,N_8638);
and U8926 (N_8926,N_8733,N_8601);
xnor U8927 (N_8927,N_8624,N_8796);
and U8928 (N_8928,N_8698,N_8690);
nand U8929 (N_8929,N_8692,N_8734);
xnor U8930 (N_8930,N_8782,N_8672);
nand U8931 (N_8931,N_8666,N_8665);
nor U8932 (N_8932,N_8635,N_8664);
and U8933 (N_8933,N_8621,N_8626);
xnor U8934 (N_8934,N_8707,N_8655);
nand U8935 (N_8935,N_8650,N_8610);
or U8936 (N_8936,N_8616,N_8642);
or U8937 (N_8937,N_8688,N_8726);
or U8938 (N_8938,N_8761,N_8771);
nor U8939 (N_8939,N_8661,N_8730);
xnor U8940 (N_8940,N_8744,N_8730);
xor U8941 (N_8941,N_8706,N_8784);
and U8942 (N_8942,N_8616,N_8758);
nand U8943 (N_8943,N_8681,N_8768);
and U8944 (N_8944,N_8612,N_8653);
xnor U8945 (N_8945,N_8684,N_8774);
or U8946 (N_8946,N_8781,N_8752);
or U8947 (N_8947,N_8761,N_8638);
xnor U8948 (N_8948,N_8609,N_8680);
or U8949 (N_8949,N_8637,N_8692);
and U8950 (N_8950,N_8632,N_8650);
xnor U8951 (N_8951,N_8737,N_8623);
xnor U8952 (N_8952,N_8676,N_8769);
or U8953 (N_8953,N_8729,N_8763);
and U8954 (N_8954,N_8718,N_8730);
nand U8955 (N_8955,N_8787,N_8667);
nor U8956 (N_8956,N_8773,N_8665);
nor U8957 (N_8957,N_8641,N_8725);
and U8958 (N_8958,N_8617,N_8621);
or U8959 (N_8959,N_8680,N_8767);
and U8960 (N_8960,N_8742,N_8634);
nor U8961 (N_8961,N_8761,N_8607);
nor U8962 (N_8962,N_8717,N_8747);
xor U8963 (N_8963,N_8685,N_8606);
or U8964 (N_8964,N_8682,N_8630);
xor U8965 (N_8965,N_8603,N_8752);
nand U8966 (N_8966,N_8740,N_8734);
or U8967 (N_8967,N_8632,N_8767);
and U8968 (N_8968,N_8779,N_8721);
nand U8969 (N_8969,N_8793,N_8762);
xor U8970 (N_8970,N_8691,N_8687);
and U8971 (N_8971,N_8648,N_8765);
or U8972 (N_8972,N_8751,N_8693);
xor U8973 (N_8973,N_8770,N_8649);
or U8974 (N_8974,N_8652,N_8666);
nand U8975 (N_8975,N_8719,N_8639);
xor U8976 (N_8976,N_8647,N_8732);
nor U8977 (N_8977,N_8626,N_8651);
and U8978 (N_8978,N_8682,N_8739);
and U8979 (N_8979,N_8719,N_8792);
or U8980 (N_8980,N_8767,N_8710);
and U8981 (N_8981,N_8767,N_8779);
nor U8982 (N_8982,N_8737,N_8630);
and U8983 (N_8983,N_8651,N_8793);
and U8984 (N_8984,N_8795,N_8688);
or U8985 (N_8985,N_8787,N_8733);
nand U8986 (N_8986,N_8628,N_8768);
or U8987 (N_8987,N_8724,N_8624);
and U8988 (N_8988,N_8735,N_8661);
or U8989 (N_8989,N_8733,N_8771);
xor U8990 (N_8990,N_8780,N_8692);
nand U8991 (N_8991,N_8694,N_8724);
xor U8992 (N_8992,N_8729,N_8635);
or U8993 (N_8993,N_8720,N_8619);
and U8994 (N_8994,N_8619,N_8660);
or U8995 (N_8995,N_8721,N_8603);
nand U8996 (N_8996,N_8692,N_8771);
xnor U8997 (N_8997,N_8600,N_8767);
and U8998 (N_8998,N_8670,N_8699);
and U8999 (N_8999,N_8727,N_8631);
nand U9000 (N_9000,N_8962,N_8905);
xor U9001 (N_9001,N_8838,N_8886);
or U9002 (N_9002,N_8880,N_8887);
xnor U9003 (N_9003,N_8981,N_8999);
and U9004 (N_9004,N_8970,N_8835);
xor U9005 (N_9005,N_8954,N_8992);
nor U9006 (N_9006,N_8995,N_8944);
xnor U9007 (N_9007,N_8934,N_8890);
xnor U9008 (N_9008,N_8878,N_8883);
and U9009 (N_9009,N_8881,N_8913);
nor U9010 (N_9010,N_8851,N_8917);
or U9011 (N_9011,N_8935,N_8839);
and U9012 (N_9012,N_8806,N_8870);
xnor U9013 (N_9013,N_8802,N_8943);
nand U9014 (N_9014,N_8859,N_8977);
or U9015 (N_9015,N_8831,N_8948);
or U9016 (N_9016,N_8902,N_8957);
nor U9017 (N_9017,N_8976,N_8847);
and U9018 (N_9018,N_8896,N_8939);
nor U9019 (N_9019,N_8958,N_8952);
xor U9020 (N_9020,N_8843,N_8991);
xor U9021 (N_9021,N_8900,N_8915);
nand U9022 (N_9022,N_8926,N_8894);
nand U9023 (N_9023,N_8908,N_8821);
nand U9024 (N_9024,N_8842,N_8959);
and U9025 (N_9025,N_8845,N_8929);
or U9026 (N_9026,N_8868,N_8918);
and U9027 (N_9027,N_8955,N_8882);
xor U9028 (N_9028,N_8893,N_8884);
or U9029 (N_9029,N_8849,N_8978);
and U9030 (N_9030,N_8996,N_8805);
nor U9031 (N_9031,N_8951,N_8993);
and U9032 (N_9032,N_8973,N_8897);
or U9033 (N_9033,N_8994,N_8830);
and U9034 (N_9034,N_8914,N_8850);
nand U9035 (N_9035,N_8815,N_8810);
nor U9036 (N_9036,N_8860,N_8803);
nor U9037 (N_9037,N_8809,N_8972);
and U9038 (N_9038,N_8931,N_8899);
nand U9039 (N_9039,N_8949,N_8875);
nor U9040 (N_9040,N_8820,N_8990);
nor U9041 (N_9041,N_8818,N_8930);
and U9042 (N_9042,N_8925,N_8819);
and U9043 (N_9043,N_8937,N_8927);
xnor U9044 (N_9044,N_8812,N_8832);
nor U9045 (N_9045,N_8855,N_8841);
nor U9046 (N_9046,N_8956,N_8857);
nand U9047 (N_9047,N_8828,N_8919);
or U9048 (N_9048,N_8848,N_8969);
nand U9049 (N_9049,N_8942,N_8910);
nand U9050 (N_9050,N_8984,N_8940);
nor U9051 (N_9051,N_8862,N_8861);
and U9052 (N_9052,N_8986,N_8968);
nor U9053 (N_9053,N_8824,N_8907);
and U9054 (N_9054,N_8936,N_8871);
nand U9055 (N_9055,N_8858,N_8980);
or U9056 (N_9056,N_8852,N_8898);
or U9057 (N_9057,N_8801,N_8998);
nor U9058 (N_9058,N_8891,N_8877);
xnor U9059 (N_9059,N_8854,N_8814);
and U9060 (N_9060,N_8879,N_8804);
xor U9061 (N_9061,N_8846,N_8950);
nor U9062 (N_9062,N_8833,N_8892);
or U9063 (N_9063,N_8924,N_8853);
xor U9064 (N_9064,N_8941,N_8953);
nand U9065 (N_9065,N_8921,N_8825);
xnor U9066 (N_9066,N_8922,N_8836);
nor U9067 (N_9067,N_8888,N_8933);
xnor U9068 (N_9068,N_8840,N_8997);
and U9069 (N_9069,N_8889,N_8982);
xnor U9070 (N_9070,N_8826,N_8965);
and U9071 (N_9071,N_8834,N_8966);
xor U9072 (N_9072,N_8963,N_8989);
nand U9073 (N_9073,N_8974,N_8817);
nand U9074 (N_9074,N_8863,N_8983);
and U9075 (N_9075,N_8979,N_8988);
nand U9076 (N_9076,N_8837,N_8909);
or U9077 (N_9077,N_8975,N_8923);
nand U9078 (N_9078,N_8987,N_8829);
and U9079 (N_9079,N_8822,N_8932);
nor U9080 (N_9080,N_8985,N_8844);
and U9081 (N_9081,N_8916,N_8945);
or U9082 (N_9082,N_8856,N_8971);
or U9083 (N_9083,N_8901,N_8960);
and U9084 (N_9084,N_8885,N_8869);
and U9085 (N_9085,N_8800,N_8906);
or U9086 (N_9086,N_8808,N_8827);
or U9087 (N_9087,N_8872,N_8816);
xnor U9088 (N_9088,N_8823,N_8920);
or U9089 (N_9089,N_8938,N_8964);
nand U9090 (N_9090,N_8967,N_8873);
xor U9091 (N_9091,N_8904,N_8928);
xnor U9092 (N_9092,N_8864,N_8903);
and U9093 (N_9093,N_8807,N_8947);
nand U9094 (N_9094,N_8911,N_8813);
xnor U9095 (N_9095,N_8866,N_8867);
nor U9096 (N_9096,N_8811,N_8865);
nand U9097 (N_9097,N_8912,N_8874);
and U9098 (N_9098,N_8946,N_8876);
or U9099 (N_9099,N_8961,N_8895);
or U9100 (N_9100,N_8823,N_8984);
xnor U9101 (N_9101,N_8952,N_8915);
nor U9102 (N_9102,N_8870,N_8973);
nor U9103 (N_9103,N_8974,N_8807);
xnor U9104 (N_9104,N_8900,N_8881);
nor U9105 (N_9105,N_8926,N_8863);
and U9106 (N_9106,N_8802,N_8936);
or U9107 (N_9107,N_8857,N_8842);
nand U9108 (N_9108,N_8962,N_8841);
and U9109 (N_9109,N_8869,N_8817);
or U9110 (N_9110,N_8885,N_8886);
nor U9111 (N_9111,N_8997,N_8964);
and U9112 (N_9112,N_8829,N_8909);
or U9113 (N_9113,N_8955,N_8852);
nand U9114 (N_9114,N_8807,N_8898);
or U9115 (N_9115,N_8842,N_8852);
nor U9116 (N_9116,N_8878,N_8927);
nand U9117 (N_9117,N_8909,N_8980);
or U9118 (N_9118,N_8933,N_8883);
xor U9119 (N_9119,N_8816,N_8810);
nand U9120 (N_9120,N_8851,N_8827);
or U9121 (N_9121,N_8910,N_8920);
or U9122 (N_9122,N_8904,N_8914);
nor U9123 (N_9123,N_8850,N_8902);
or U9124 (N_9124,N_8943,N_8902);
nand U9125 (N_9125,N_8811,N_8835);
nor U9126 (N_9126,N_8815,N_8946);
nor U9127 (N_9127,N_8866,N_8827);
xnor U9128 (N_9128,N_8897,N_8908);
or U9129 (N_9129,N_8896,N_8807);
or U9130 (N_9130,N_8956,N_8868);
nand U9131 (N_9131,N_8811,N_8898);
xor U9132 (N_9132,N_8809,N_8940);
nand U9133 (N_9133,N_8865,N_8889);
xor U9134 (N_9134,N_8950,N_8931);
or U9135 (N_9135,N_8809,N_8923);
and U9136 (N_9136,N_8963,N_8821);
or U9137 (N_9137,N_8994,N_8971);
xor U9138 (N_9138,N_8853,N_8902);
nor U9139 (N_9139,N_8948,N_8861);
xnor U9140 (N_9140,N_8916,N_8857);
xor U9141 (N_9141,N_8836,N_8842);
xor U9142 (N_9142,N_8831,N_8997);
xor U9143 (N_9143,N_8888,N_8821);
xnor U9144 (N_9144,N_8981,N_8920);
or U9145 (N_9145,N_8875,N_8905);
nand U9146 (N_9146,N_8958,N_8820);
and U9147 (N_9147,N_8879,N_8803);
nand U9148 (N_9148,N_8872,N_8992);
xor U9149 (N_9149,N_8954,N_8840);
xnor U9150 (N_9150,N_8829,N_8965);
nor U9151 (N_9151,N_8843,N_8982);
nor U9152 (N_9152,N_8880,N_8897);
nand U9153 (N_9153,N_8942,N_8930);
and U9154 (N_9154,N_8874,N_8851);
nor U9155 (N_9155,N_8890,N_8980);
nand U9156 (N_9156,N_8951,N_8813);
and U9157 (N_9157,N_8953,N_8990);
nor U9158 (N_9158,N_8950,N_8917);
or U9159 (N_9159,N_8966,N_8801);
xnor U9160 (N_9160,N_8890,N_8913);
xor U9161 (N_9161,N_8986,N_8881);
or U9162 (N_9162,N_8803,N_8935);
nand U9163 (N_9163,N_8851,N_8910);
nand U9164 (N_9164,N_8970,N_8888);
or U9165 (N_9165,N_8905,N_8868);
nand U9166 (N_9166,N_8889,N_8959);
and U9167 (N_9167,N_8851,N_8869);
xnor U9168 (N_9168,N_8824,N_8831);
nor U9169 (N_9169,N_8808,N_8854);
nand U9170 (N_9170,N_8931,N_8941);
nand U9171 (N_9171,N_8945,N_8882);
and U9172 (N_9172,N_8976,N_8946);
or U9173 (N_9173,N_8967,N_8936);
or U9174 (N_9174,N_8863,N_8932);
nor U9175 (N_9175,N_8807,N_8911);
nor U9176 (N_9176,N_8994,N_8862);
or U9177 (N_9177,N_8886,N_8865);
nor U9178 (N_9178,N_8842,N_8991);
nor U9179 (N_9179,N_8894,N_8961);
xnor U9180 (N_9180,N_8978,N_8806);
xnor U9181 (N_9181,N_8882,N_8826);
xnor U9182 (N_9182,N_8997,N_8807);
nand U9183 (N_9183,N_8893,N_8982);
or U9184 (N_9184,N_8956,N_8903);
nand U9185 (N_9185,N_8990,N_8869);
xor U9186 (N_9186,N_8822,N_8880);
and U9187 (N_9187,N_8883,N_8900);
or U9188 (N_9188,N_8899,N_8970);
xnor U9189 (N_9189,N_8916,N_8866);
or U9190 (N_9190,N_8840,N_8953);
nor U9191 (N_9191,N_8822,N_8966);
xor U9192 (N_9192,N_8940,N_8973);
and U9193 (N_9193,N_8959,N_8927);
nand U9194 (N_9194,N_8827,N_8837);
nor U9195 (N_9195,N_8911,N_8866);
nand U9196 (N_9196,N_8877,N_8961);
nand U9197 (N_9197,N_8837,N_8896);
nor U9198 (N_9198,N_8937,N_8849);
or U9199 (N_9199,N_8942,N_8884);
nand U9200 (N_9200,N_9018,N_9056);
nand U9201 (N_9201,N_9083,N_9059);
nor U9202 (N_9202,N_9051,N_9033);
nand U9203 (N_9203,N_9043,N_9188);
or U9204 (N_9204,N_9163,N_9032);
or U9205 (N_9205,N_9138,N_9076);
nand U9206 (N_9206,N_9180,N_9161);
nand U9207 (N_9207,N_9071,N_9149);
xor U9208 (N_9208,N_9072,N_9079);
nand U9209 (N_9209,N_9036,N_9114);
nand U9210 (N_9210,N_9034,N_9005);
nor U9211 (N_9211,N_9097,N_9062);
or U9212 (N_9212,N_9133,N_9102);
nor U9213 (N_9213,N_9131,N_9004);
or U9214 (N_9214,N_9027,N_9077);
xor U9215 (N_9215,N_9127,N_9195);
or U9216 (N_9216,N_9022,N_9153);
nand U9217 (N_9217,N_9098,N_9150);
nand U9218 (N_9218,N_9094,N_9189);
nor U9219 (N_9219,N_9158,N_9015);
or U9220 (N_9220,N_9060,N_9176);
xnor U9221 (N_9221,N_9115,N_9066);
xnor U9222 (N_9222,N_9081,N_9178);
nor U9223 (N_9223,N_9041,N_9106);
and U9224 (N_9224,N_9168,N_9135);
or U9225 (N_9225,N_9073,N_9017);
nand U9226 (N_9226,N_9055,N_9196);
xnor U9227 (N_9227,N_9112,N_9109);
and U9228 (N_9228,N_9101,N_9089);
nand U9229 (N_9229,N_9095,N_9031);
or U9230 (N_9230,N_9049,N_9105);
or U9231 (N_9231,N_9053,N_9169);
nand U9232 (N_9232,N_9046,N_9136);
nand U9233 (N_9233,N_9194,N_9019);
nor U9234 (N_9234,N_9035,N_9117);
or U9235 (N_9235,N_9086,N_9159);
nand U9236 (N_9236,N_9170,N_9093);
or U9237 (N_9237,N_9198,N_9167);
nor U9238 (N_9238,N_9122,N_9028);
or U9239 (N_9239,N_9099,N_9186);
nor U9240 (N_9240,N_9008,N_9160);
xor U9241 (N_9241,N_9087,N_9070);
xnor U9242 (N_9242,N_9184,N_9132);
or U9243 (N_9243,N_9152,N_9143);
nand U9244 (N_9244,N_9154,N_9045);
or U9245 (N_9245,N_9002,N_9107);
and U9246 (N_9246,N_9088,N_9185);
and U9247 (N_9247,N_9047,N_9048);
or U9248 (N_9248,N_9192,N_9108);
nor U9249 (N_9249,N_9040,N_9010);
xnor U9250 (N_9250,N_9074,N_9157);
nand U9251 (N_9251,N_9156,N_9110);
and U9252 (N_9252,N_9111,N_9164);
or U9253 (N_9253,N_9061,N_9068);
nand U9254 (N_9254,N_9006,N_9121);
and U9255 (N_9255,N_9120,N_9082);
nand U9256 (N_9256,N_9054,N_9003);
or U9257 (N_9257,N_9025,N_9011);
or U9258 (N_9258,N_9057,N_9029);
xnor U9259 (N_9259,N_9058,N_9050);
and U9260 (N_9260,N_9151,N_9030);
or U9261 (N_9261,N_9007,N_9137);
and U9262 (N_9262,N_9013,N_9012);
nor U9263 (N_9263,N_9139,N_9175);
nor U9264 (N_9264,N_9009,N_9144);
and U9265 (N_9265,N_9155,N_9125);
nor U9266 (N_9266,N_9199,N_9118);
and U9267 (N_9267,N_9140,N_9113);
nor U9268 (N_9268,N_9080,N_9119);
and U9269 (N_9269,N_9147,N_9044);
nor U9270 (N_9270,N_9166,N_9123);
nor U9271 (N_9271,N_9038,N_9000);
nand U9272 (N_9272,N_9171,N_9134);
and U9273 (N_9273,N_9177,N_9020);
nand U9274 (N_9274,N_9162,N_9037);
xor U9275 (N_9275,N_9001,N_9085);
nor U9276 (N_9276,N_9096,N_9078);
nand U9277 (N_9277,N_9067,N_9116);
nand U9278 (N_9278,N_9090,N_9126);
nand U9279 (N_9279,N_9069,N_9182);
or U9280 (N_9280,N_9141,N_9128);
nand U9281 (N_9281,N_9191,N_9024);
and U9282 (N_9282,N_9052,N_9174);
nor U9283 (N_9283,N_9065,N_9100);
xnor U9284 (N_9284,N_9084,N_9092);
and U9285 (N_9285,N_9091,N_9104);
nand U9286 (N_9286,N_9181,N_9190);
nand U9287 (N_9287,N_9179,N_9130);
nor U9288 (N_9288,N_9145,N_9187);
nor U9289 (N_9289,N_9064,N_9146);
or U9290 (N_9290,N_9142,N_9129);
xnor U9291 (N_9291,N_9021,N_9026);
nand U9292 (N_9292,N_9124,N_9197);
nand U9293 (N_9293,N_9014,N_9172);
and U9294 (N_9294,N_9039,N_9042);
or U9295 (N_9295,N_9103,N_9016);
xnor U9296 (N_9296,N_9075,N_9193);
or U9297 (N_9297,N_9173,N_9063);
and U9298 (N_9298,N_9023,N_9165);
or U9299 (N_9299,N_9183,N_9148);
and U9300 (N_9300,N_9163,N_9153);
xnor U9301 (N_9301,N_9005,N_9031);
xor U9302 (N_9302,N_9001,N_9100);
or U9303 (N_9303,N_9145,N_9040);
or U9304 (N_9304,N_9163,N_9012);
nand U9305 (N_9305,N_9013,N_9125);
nor U9306 (N_9306,N_9165,N_9186);
nand U9307 (N_9307,N_9106,N_9128);
or U9308 (N_9308,N_9195,N_9196);
xor U9309 (N_9309,N_9096,N_9040);
nand U9310 (N_9310,N_9086,N_9039);
or U9311 (N_9311,N_9100,N_9075);
nor U9312 (N_9312,N_9145,N_9025);
xor U9313 (N_9313,N_9118,N_9072);
nor U9314 (N_9314,N_9176,N_9077);
nand U9315 (N_9315,N_9024,N_9128);
and U9316 (N_9316,N_9195,N_9199);
and U9317 (N_9317,N_9138,N_9176);
or U9318 (N_9318,N_9139,N_9171);
or U9319 (N_9319,N_9006,N_9141);
and U9320 (N_9320,N_9177,N_9011);
and U9321 (N_9321,N_9178,N_9006);
or U9322 (N_9322,N_9138,N_9060);
nor U9323 (N_9323,N_9066,N_9022);
xnor U9324 (N_9324,N_9147,N_9177);
xor U9325 (N_9325,N_9104,N_9071);
or U9326 (N_9326,N_9134,N_9163);
xnor U9327 (N_9327,N_9146,N_9086);
nand U9328 (N_9328,N_9043,N_9166);
nor U9329 (N_9329,N_9183,N_9142);
nand U9330 (N_9330,N_9122,N_9016);
nand U9331 (N_9331,N_9133,N_9034);
nor U9332 (N_9332,N_9164,N_9003);
and U9333 (N_9333,N_9029,N_9113);
xor U9334 (N_9334,N_9100,N_9196);
xnor U9335 (N_9335,N_9196,N_9167);
nor U9336 (N_9336,N_9161,N_9111);
nand U9337 (N_9337,N_9023,N_9102);
or U9338 (N_9338,N_9006,N_9036);
nand U9339 (N_9339,N_9079,N_9101);
nor U9340 (N_9340,N_9059,N_9034);
nor U9341 (N_9341,N_9175,N_9117);
or U9342 (N_9342,N_9046,N_9062);
and U9343 (N_9343,N_9031,N_9071);
nand U9344 (N_9344,N_9046,N_9009);
nor U9345 (N_9345,N_9134,N_9061);
nand U9346 (N_9346,N_9095,N_9089);
and U9347 (N_9347,N_9042,N_9184);
nor U9348 (N_9348,N_9084,N_9145);
nand U9349 (N_9349,N_9183,N_9106);
nor U9350 (N_9350,N_9134,N_9092);
or U9351 (N_9351,N_9113,N_9124);
xnor U9352 (N_9352,N_9069,N_9044);
nand U9353 (N_9353,N_9176,N_9193);
nand U9354 (N_9354,N_9166,N_9145);
or U9355 (N_9355,N_9017,N_9071);
nand U9356 (N_9356,N_9078,N_9032);
and U9357 (N_9357,N_9175,N_9047);
xor U9358 (N_9358,N_9187,N_9127);
nor U9359 (N_9359,N_9193,N_9074);
nand U9360 (N_9360,N_9016,N_9128);
or U9361 (N_9361,N_9165,N_9108);
nand U9362 (N_9362,N_9073,N_9189);
nand U9363 (N_9363,N_9023,N_9018);
nor U9364 (N_9364,N_9184,N_9059);
or U9365 (N_9365,N_9102,N_9195);
xor U9366 (N_9366,N_9087,N_9139);
nor U9367 (N_9367,N_9031,N_9161);
nand U9368 (N_9368,N_9133,N_9008);
or U9369 (N_9369,N_9133,N_9058);
and U9370 (N_9370,N_9018,N_9180);
and U9371 (N_9371,N_9016,N_9106);
nand U9372 (N_9372,N_9118,N_9174);
or U9373 (N_9373,N_9092,N_9157);
nand U9374 (N_9374,N_9006,N_9037);
xor U9375 (N_9375,N_9131,N_9018);
nor U9376 (N_9376,N_9126,N_9133);
nand U9377 (N_9377,N_9129,N_9035);
xor U9378 (N_9378,N_9021,N_9000);
xnor U9379 (N_9379,N_9062,N_9069);
nor U9380 (N_9380,N_9188,N_9089);
or U9381 (N_9381,N_9190,N_9059);
or U9382 (N_9382,N_9098,N_9083);
and U9383 (N_9383,N_9070,N_9130);
nand U9384 (N_9384,N_9123,N_9164);
or U9385 (N_9385,N_9029,N_9047);
xor U9386 (N_9386,N_9003,N_9190);
and U9387 (N_9387,N_9005,N_9004);
or U9388 (N_9388,N_9130,N_9059);
or U9389 (N_9389,N_9094,N_9003);
xnor U9390 (N_9390,N_9151,N_9112);
nand U9391 (N_9391,N_9046,N_9053);
nand U9392 (N_9392,N_9082,N_9150);
and U9393 (N_9393,N_9166,N_9185);
nor U9394 (N_9394,N_9061,N_9075);
xor U9395 (N_9395,N_9132,N_9073);
nor U9396 (N_9396,N_9047,N_9094);
nand U9397 (N_9397,N_9072,N_9112);
xor U9398 (N_9398,N_9090,N_9111);
nand U9399 (N_9399,N_9023,N_9162);
and U9400 (N_9400,N_9339,N_9207);
nand U9401 (N_9401,N_9299,N_9292);
and U9402 (N_9402,N_9348,N_9282);
or U9403 (N_9403,N_9344,N_9235);
or U9404 (N_9404,N_9330,N_9377);
nand U9405 (N_9405,N_9390,N_9316);
or U9406 (N_9406,N_9386,N_9397);
nor U9407 (N_9407,N_9213,N_9347);
nand U9408 (N_9408,N_9322,N_9245);
or U9409 (N_9409,N_9206,N_9216);
or U9410 (N_9410,N_9358,N_9312);
or U9411 (N_9411,N_9369,N_9332);
or U9412 (N_9412,N_9258,N_9357);
nand U9413 (N_9413,N_9274,N_9266);
and U9414 (N_9414,N_9264,N_9331);
nor U9415 (N_9415,N_9210,N_9285);
xor U9416 (N_9416,N_9227,N_9387);
xnor U9417 (N_9417,N_9372,N_9342);
nor U9418 (N_9418,N_9222,N_9228);
nor U9419 (N_9419,N_9248,N_9305);
nand U9420 (N_9420,N_9336,N_9259);
nand U9421 (N_9421,N_9275,N_9204);
or U9422 (N_9422,N_9220,N_9229);
and U9423 (N_9423,N_9223,N_9252);
or U9424 (N_9424,N_9324,N_9205);
nor U9425 (N_9425,N_9380,N_9250);
or U9426 (N_9426,N_9329,N_9319);
or U9427 (N_9427,N_9277,N_9359);
or U9428 (N_9428,N_9366,N_9306);
xor U9429 (N_9429,N_9237,N_9289);
xor U9430 (N_9430,N_9238,N_9265);
xnor U9431 (N_9431,N_9374,N_9356);
nand U9432 (N_9432,N_9230,N_9364);
and U9433 (N_9433,N_9218,N_9307);
nand U9434 (N_9434,N_9212,N_9360);
or U9435 (N_9435,N_9224,N_9249);
and U9436 (N_9436,N_9368,N_9343);
nor U9437 (N_9437,N_9269,N_9239);
or U9438 (N_9438,N_9338,N_9236);
and U9439 (N_9439,N_9395,N_9202);
nor U9440 (N_9440,N_9389,N_9225);
or U9441 (N_9441,N_9349,N_9209);
or U9442 (N_9442,N_9291,N_9313);
and U9443 (N_9443,N_9333,N_9398);
or U9444 (N_9444,N_9276,N_9352);
nor U9445 (N_9445,N_9373,N_9328);
xnor U9446 (N_9446,N_9345,N_9355);
nand U9447 (N_9447,N_9382,N_9244);
nor U9448 (N_9448,N_9271,N_9262);
or U9449 (N_9449,N_9215,N_9351);
nor U9450 (N_9450,N_9391,N_9399);
nand U9451 (N_9451,N_9281,N_9214);
xor U9452 (N_9452,N_9273,N_9367);
and U9453 (N_9453,N_9318,N_9217);
xnor U9454 (N_9454,N_9354,N_9246);
or U9455 (N_9455,N_9392,N_9350);
xnor U9456 (N_9456,N_9303,N_9226);
nand U9457 (N_9457,N_9283,N_9396);
nor U9458 (N_9458,N_9286,N_9261);
nand U9459 (N_9459,N_9280,N_9363);
or U9460 (N_9460,N_9290,N_9201);
or U9461 (N_9461,N_9375,N_9256);
nand U9462 (N_9462,N_9384,N_9242);
xnor U9463 (N_9463,N_9231,N_9243);
or U9464 (N_9464,N_9300,N_9295);
nor U9465 (N_9465,N_9308,N_9340);
or U9466 (N_9466,N_9334,N_9388);
xnor U9467 (N_9467,N_9278,N_9309);
xor U9468 (N_9468,N_9211,N_9346);
or U9469 (N_9469,N_9203,N_9221);
nor U9470 (N_9470,N_9370,N_9341);
nor U9471 (N_9471,N_9267,N_9219);
and U9472 (N_9472,N_9379,N_9200);
xnor U9473 (N_9473,N_9335,N_9297);
and U9474 (N_9474,N_9257,N_9240);
or U9475 (N_9475,N_9287,N_9381);
xnor U9476 (N_9476,N_9361,N_9279);
or U9477 (N_9477,N_9365,N_9301);
and U9478 (N_9478,N_9323,N_9315);
xnor U9479 (N_9479,N_9270,N_9325);
xor U9480 (N_9480,N_9293,N_9394);
or U9481 (N_9481,N_9208,N_9310);
or U9482 (N_9482,N_9272,N_9327);
nand U9483 (N_9483,N_9260,N_9233);
and U9484 (N_9484,N_9296,N_9321);
nor U9485 (N_9485,N_9362,N_9284);
and U9486 (N_9486,N_9251,N_9320);
nor U9487 (N_9487,N_9268,N_9393);
or U9488 (N_9488,N_9254,N_9326);
xnor U9489 (N_9489,N_9255,N_9383);
nand U9490 (N_9490,N_9234,N_9241);
xnor U9491 (N_9491,N_9263,N_9288);
xor U9492 (N_9492,N_9314,N_9378);
or U9493 (N_9493,N_9298,N_9311);
and U9494 (N_9494,N_9302,N_9353);
and U9495 (N_9495,N_9376,N_9232);
and U9496 (N_9496,N_9294,N_9337);
and U9497 (N_9497,N_9385,N_9371);
nand U9498 (N_9498,N_9247,N_9253);
xnor U9499 (N_9499,N_9317,N_9304);
and U9500 (N_9500,N_9287,N_9221);
or U9501 (N_9501,N_9233,N_9358);
nor U9502 (N_9502,N_9284,N_9316);
nand U9503 (N_9503,N_9377,N_9270);
nor U9504 (N_9504,N_9256,N_9247);
or U9505 (N_9505,N_9223,N_9386);
or U9506 (N_9506,N_9350,N_9311);
nand U9507 (N_9507,N_9383,N_9388);
xnor U9508 (N_9508,N_9393,N_9308);
nand U9509 (N_9509,N_9299,N_9304);
xor U9510 (N_9510,N_9357,N_9237);
xnor U9511 (N_9511,N_9337,N_9311);
or U9512 (N_9512,N_9216,N_9237);
xnor U9513 (N_9513,N_9222,N_9307);
nand U9514 (N_9514,N_9291,N_9332);
and U9515 (N_9515,N_9200,N_9262);
nand U9516 (N_9516,N_9361,N_9308);
nand U9517 (N_9517,N_9216,N_9241);
nor U9518 (N_9518,N_9355,N_9260);
xnor U9519 (N_9519,N_9357,N_9251);
nand U9520 (N_9520,N_9314,N_9252);
nand U9521 (N_9521,N_9306,N_9217);
xnor U9522 (N_9522,N_9210,N_9208);
or U9523 (N_9523,N_9314,N_9276);
or U9524 (N_9524,N_9345,N_9230);
nor U9525 (N_9525,N_9354,N_9257);
nor U9526 (N_9526,N_9268,N_9271);
or U9527 (N_9527,N_9227,N_9237);
or U9528 (N_9528,N_9247,N_9379);
or U9529 (N_9529,N_9302,N_9233);
or U9530 (N_9530,N_9377,N_9212);
xor U9531 (N_9531,N_9366,N_9291);
xor U9532 (N_9532,N_9381,N_9351);
xnor U9533 (N_9533,N_9217,N_9368);
or U9534 (N_9534,N_9297,N_9325);
and U9535 (N_9535,N_9227,N_9207);
xor U9536 (N_9536,N_9275,N_9396);
and U9537 (N_9537,N_9318,N_9280);
or U9538 (N_9538,N_9285,N_9377);
xnor U9539 (N_9539,N_9335,N_9315);
and U9540 (N_9540,N_9281,N_9347);
and U9541 (N_9541,N_9207,N_9213);
nand U9542 (N_9542,N_9346,N_9247);
xor U9543 (N_9543,N_9286,N_9215);
nand U9544 (N_9544,N_9325,N_9356);
nor U9545 (N_9545,N_9356,N_9306);
or U9546 (N_9546,N_9232,N_9306);
or U9547 (N_9547,N_9261,N_9281);
and U9548 (N_9548,N_9293,N_9243);
xnor U9549 (N_9549,N_9295,N_9367);
and U9550 (N_9550,N_9282,N_9342);
nand U9551 (N_9551,N_9382,N_9389);
nand U9552 (N_9552,N_9210,N_9200);
and U9553 (N_9553,N_9373,N_9315);
xnor U9554 (N_9554,N_9226,N_9242);
nor U9555 (N_9555,N_9379,N_9392);
and U9556 (N_9556,N_9385,N_9230);
xor U9557 (N_9557,N_9240,N_9225);
or U9558 (N_9558,N_9254,N_9244);
xor U9559 (N_9559,N_9300,N_9315);
and U9560 (N_9560,N_9391,N_9288);
nand U9561 (N_9561,N_9311,N_9295);
and U9562 (N_9562,N_9210,N_9370);
xor U9563 (N_9563,N_9333,N_9225);
or U9564 (N_9564,N_9288,N_9243);
xor U9565 (N_9565,N_9388,N_9312);
nor U9566 (N_9566,N_9356,N_9389);
nor U9567 (N_9567,N_9234,N_9350);
nor U9568 (N_9568,N_9209,N_9216);
or U9569 (N_9569,N_9263,N_9391);
nand U9570 (N_9570,N_9201,N_9229);
nand U9571 (N_9571,N_9387,N_9330);
or U9572 (N_9572,N_9215,N_9314);
nand U9573 (N_9573,N_9331,N_9277);
nand U9574 (N_9574,N_9281,N_9265);
nand U9575 (N_9575,N_9364,N_9293);
and U9576 (N_9576,N_9338,N_9385);
and U9577 (N_9577,N_9267,N_9328);
nor U9578 (N_9578,N_9229,N_9296);
nor U9579 (N_9579,N_9288,N_9292);
xor U9580 (N_9580,N_9367,N_9223);
xor U9581 (N_9581,N_9254,N_9256);
and U9582 (N_9582,N_9271,N_9227);
or U9583 (N_9583,N_9328,N_9370);
nor U9584 (N_9584,N_9339,N_9206);
xnor U9585 (N_9585,N_9223,N_9333);
and U9586 (N_9586,N_9296,N_9399);
nor U9587 (N_9587,N_9240,N_9292);
nor U9588 (N_9588,N_9328,N_9376);
nand U9589 (N_9589,N_9390,N_9226);
nand U9590 (N_9590,N_9283,N_9344);
xnor U9591 (N_9591,N_9354,N_9328);
nor U9592 (N_9592,N_9305,N_9277);
nand U9593 (N_9593,N_9327,N_9265);
or U9594 (N_9594,N_9262,N_9385);
nand U9595 (N_9595,N_9321,N_9293);
or U9596 (N_9596,N_9210,N_9348);
nor U9597 (N_9597,N_9250,N_9394);
or U9598 (N_9598,N_9360,N_9359);
or U9599 (N_9599,N_9374,N_9344);
nand U9600 (N_9600,N_9509,N_9457);
nor U9601 (N_9601,N_9502,N_9456);
nand U9602 (N_9602,N_9407,N_9520);
nand U9603 (N_9603,N_9402,N_9555);
nor U9604 (N_9604,N_9417,N_9405);
xor U9605 (N_9605,N_9531,N_9472);
and U9606 (N_9606,N_9506,N_9533);
nor U9607 (N_9607,N_9521,N_9508);
or U9608 (N_9608,N_9418,N_9486);
nor U9609 (N_9609,N_9541,N_9538);
and U9610 (N_9610,N_9454,N_9503);
nand U9611 (N_9611,N_9567,N_9543);
nand U9612 (N_9612,N_9576,N_9469);
or U9613 (N_9613,N_9551,N_9411);
nand U9614 (N_9614,N_9451,N_9569);
xor U9615 (N_9615,N_9578,N_9568);
xnor U9616 (N_9616,N_9459,N_9462);
xnor U9617 (N_9617,N_9501,N_9545);
and U9618 (N_9618,N_9478,N_9516);
xor U9619 (N_9619,N_9484,N_9515);
and U9620 (N_9620,N_9575,N_9514);
xor U9621 (N_9621,N_9412,N_9585);
and U9622 (N_9622,N_9413,N_9445);
or U9623 (N_9623,N_9430,N_9554);
nand U9624 (N_9624,N_9439,N_9429);
and U9625 (N_9625,N_9489,N_9587);
nand U9626 (N_9626,N_9572,N_9561);
or U9627 (N_9627,N_9547,N_9530);
nand U9628 (N_9628,N_9477,N_9452);
nand U9629 (N_9629,N_9599,N_9577);
or U9630 (N_9630,N_9409,N_9450);
nand U9631 (N_9631,N_9434,N_9461);
nor U9632 (N_9632,N_9579,N_9422);
xor U9633 (N_9633,N_9475,N_9519);
nor U9634 (N_9634,N_9426,N_9565);
nand U9635 (N_9635,N_9574,N_9593);
and U9636 (N_9636,N_9562,N_9473);
xor U9637 (N_9637,N_9594,N_9573);
nor U9638 (N_9638,N_9586,N_9464);
xnor U9639 (N_9639,N_9490,N_9497);
nor U9640 (N_9640,N_9588,N_9589);
nand U9641 (N_9641,N_9527,N_9556);
and U9642 (N_9642,N_9458,N_9525);
and U9643 (N_9643,N_9485,N_9564);
nand U9644 (N_9644,N_9544,N_9592);
or U9645 (N_9645,N_9499,N_9535);
and U9646 (N_9646,N_9552,N_9548);
xnor U9647 (N_9647,N_9449,N_9518);
nand U9648 (N_9648,N_9460,N_9400);
nand U9649 (N_9649,N_9537,N_9546);
or U9650 (N_9650,N_9557,N_9491);
xor U9651 (N_9651,N_9500,N_9424);
nor U9652 (N_9652,N_9483,N_9421);
nand U9653 (N_9653,N_9474,N_9580);
xor U9654 (N_9654,N_9512,N_9529);
or U9655 (N_9655,N_9408,N_9549);
and U9656 (N_9656,N_9598,N_9528);
and U9657 (N_9657,N_9425,N_9570);
xor U9658 (N_9658,N_9480,N_9436);
nand U9659 (N_9659,N_9507,N_9584);
nand U9660 (N_9660,N_9414,N_9479);
nor U9661 (N_9661,N_9596,N_9540);
or U9662 (N_9662,N_9404,N_9420);
nand U9663 (N_9663,N_9582,N_9447);
or U9664 (N_9664,N_9453,N_9583);
or U9665 (N_9665,N_9435,N_9526);
xnor U9666 (N_9666,N_9558,N_9410);
nand U9667 (N_9667,N_9510,N_9496);
and U9668 (N_9668,N_9513,N_9446);
nor U9669 (N_9669,N_9517,N_9415);
or U9670 (N_9670,N_9443,N_9504);
nor U9671 (N_9671,N_9505,N_9494);
or U9672 (N_9672,N_9481,N_9523);
and U9673 (N_9673,N_9560,N_9539);
nand U9674 (N_9674,N_9444,N_9581);
nand U9675 (N_9675,N_9465,N_9559);
xor U9676 (N_9676,N_9448,N_9571);
nor U9677 (N_9677,N_9438,N_9522);
nor U9678 (N_9678,N_9597,N_9467);
nor U9679 (N_9679,N_9498,N_9416);
nand U9680 (N_9680,N_9401,N_9433);
nand U9681 (N_9681,N_9524,N_9553);
nor U9682 (N_9682,N_9488,N_9455);
xnor U9683 (N_9683,N_9428,N_9437);
nor U9684 (N_9684,N_9487,N_9482);
nor U9685 (N_9685,N_9595,N_9463);
and U9686 (N_9686,N_9440,N_9534);
nor U9687 (N_9687,N_9470,N_9532);
nor U9688 (N_9688,N_9550,N_9419);
nor U9689 (N_9689,N_9536,N_9442);
and U9690 (N_9690,N_9542,N_9423);
or U9691 (N_9691,N_9468,N_9591);
nand U9692 (N_9692,N_9403,N_9495);
and U9693 (N_9693,N_9432,N_9466);
nor U9694 (N_9694,N_9563,N_9441);
xor U9695 (N_9695,N_9590,N_9476);
or U9696 (N_9696,N_9493,N_9431);
and U9697 (N_9697,N_9566,N_9511);
nand U9698 (N_9698,N_9492,N_9406);
nor U9699 (N_9699,N_9471,N_9427);
or U9700 (N_9700,N_9534,N_9435);
xor U9701 (N_9701,N_9497,N_9499);
xnor U9702 (N_9702,N_9408,N_9523);
and U9703 (N_9703,N_9567,N_9503);
nor U9704 (N_9704,N_9584,N_9441);
and U9705 (N_9705,N_9491,N_9537);
and U9706 (N_9706,N_9470,N_9400);
nor U9707 (N_9707,N_9487,N_9457);
and U9708 (N_9708,N_9531,N_9424);
xnor U9709 (N_9709,N_9538,N_9591);
and U9710 (N_9710,N_9561,N_9447);
nand U9711 (N_9711,N_9558,N_9432);
nor U9712 (N_9712,N_9445,N_9549);
nand U9713 (N_9713,N_9542,N_9521);
and U9714 (N_9714,N_9434,N_9446);
and U9715 (N_9715,N_9410,N_9532);
nand U9716 (N_9716,N_9522,N_9511);
nor U9717 (N_9717,N_9488,N_9463);
nor U9718 (N_9718,N_9494,N_9578);
xnor U9719 (N_9719,N_9575,N_9460);
or U9720 (N_9720,N_9475,N_9442);
xnor U9721 (N_9721,N_9427,N_9582);
or U9722 (N_9722,N_9576,N_9504);
nand U9723 (N_9723,N_9451,N_9521);
xor U9724 (N_9724,N_9464,N_9512);
xor U9725 (N_9725,N_9583,N_9482);
xor U9726 (N_9726,N_9553,N_9476);
and U9727 (N_9727,N_9544,N_9570);
nand U9728 (N_9728,N_9441,N_9567);
or U9729 (N_9729,N_9586,N_9564);
nand U9730 (N_9730,N_9532,N_9515);
xnor U9731 (N_9731,N_9487,N_9468);
nor U9732 (N_9732,N_9462,N_9557);
nor U9733 (N_9733,N_9451,N_9453);
nand U9734 (N_9734,N_9405,N_9497);
and U9735 (N_9735,N_9417,N_9561);
or U9736 (N_9736,N_9432,N_9483);
nand U9737 (N_9737,N_9548,N_9466);
or U9738 (N_9738,N_9585,N_9510);
or U9739 (N_9739,N_9519,N_9582);
nor U9740 (N_9740,N_9571,N_9467);
or U9741 (N_9741,N_9576,N_9447);
xor U9742 (N_9742,N_9440,N_9497);
and U9743 (N_9743,N_9432,N_9486);
xor U9744 (N_9744,N_9477,N_9402);
or U9745 (N_9745,N_9591,N_9491);
xor U9746 (N_9746,N_9530,N_9517);
and U9747 (N_9747,N_9551,N_9474);
nand U9748 (N_9748,N_9514,N_9512);
nand U9749 (N_9749,N_9453,N_9447);
and U9750 (N_9750,N_9561,N_9480);
xnor U9751 (N_9751,N_9446,N_9472);
nand U9752 (N_9752,N_9414,N_9425);
and U9753 (N_9753,N_9583,N_9500);
and U9754 (N_9754,N_9541,N_9515);
or U9755 (N_9755,N_9445,N_9598);
nand U9756 (N_9756,N_9539,N_9401);
nor U9757 (N_9757,N_9440,N_9402);
or U9758 (N_9758,N_9526,N_9482);
xnor U9759 (N_9759,N_9506,N_9451);
nor U9760 (N_9760,N_9475,N_9414);
nand U9761 (N_9761,N_9425,N_9477);
nor U9762 (N_9762,N_9567,N_9502);
or U9763 (N_9763,N_9435,N_9494);
nand U9764 (N_9764,N_9519,N_9461);
xor U9765 (N_9765,N_9517,N_9426);
xnor U9766 (N_9766,N_9577,N_9561);
xnor U9767 (N_9767,N_9555,N_9462);
and U9768 (N_9768,N_9418,N_9465);
and U9769 (N_9769,N_9562,N_9456);
and U9770 (N_9770,N_9566,N_9555);
or U9771 (N_9771,N_9559,N_9562);
nand U9772 (N_9772,N_9527,N_9545);
xnor U9773 (N_9773,N_9403,N_9566);
and U9774 (N_9774,N_9575,N_9435);
xor U9775 (N_9775,N_9572,N_9425);
and U9776 (N_9776,N_9593,N_9562);
nand U9777 (N_9777,N_9404,N_9496);
nand U9778 (N_9778,N_9556,N_9473);
nand U9779 (N_9779,N_9443,N_9482);
nor U9780 (N_9780,N_9507,N_9559);
or U9781 (N_9781,N_9588,N_9568);
nor U9782 (N_9782,N_9459,N_9551);
and U9783 (N_9783,N_9402,N_9464);
nor U9784 (N_9784,N_9562,N_9461);
xnor U9785 (N_9785,N_9579,N_9586);
xor U9786 (N_9786,N_9426,N_9555);
or U9787 (N_9787,N_9405,N_9513);
xor U9788 (N_9788,N_9561,N_9555);
or U9789 (N_9789,N_9469,N_9495);
xnor U9790 (N_9790,N_9561,N_9537);
nand U9791 (N_9791,N_9445,N_9526);
and U9792 (N_9792,N_9406,N_9435);
nand U9793 (N_9793,N_9410,N_9545);
nand U9794 (N_9794,N_9563,N_9425);
or U9795 (N_9795,N_9527,N_9542);
nor U9796 (N_9796,N_9428,N_9458);
xor U9797 (N_9797,N_9460,N_9413);
nor U9798 (N_9798,N_9568,N_9569);
nor U9799 (N_9799,N_9416,N_9522);
or U9800 (N_9800,N_9795,N_9619);
nand U9801 (N_9801,N_9798,N_9664);
and U9802 (N_9802,N_9729,N_9735);
xnor U9803 (N_9803,N_9683,N_9726);
nand U9804 (N_9804,N_9780,N_9635);
or U9805 (N_9805,N_9738,N_9715);
xor U9806 (N_9806,N_9690,N_9713);
or U9807 (N_9807,N_9783,N_9751);
or U9808 (N_9808,N_9698,N_9608);
xor U9809 (N_9809,N_9772,N_9756);
nand U9810 (N_9810,N_9657,N_9719);
and U9811 (N_9811,N_9648,N_9606);
or U9812 (N_9812,N_9731,N_9760);
or U9813 (N_9813,N_9654,N_9642);
xor U9814 (N_9814,N_9623,N_9629);
or U9815 (N_9815,N_9644,N_9743);
nor U9816 (N_9816,N_9677,N_9655);
and U9817 (N_9817,N_9744,N_9651);
nor U9818 (N_9818,N_9781,N_9687);
and U9819 (N_9819,N_9730,N_9646);
nor U9820 (N_9820,N_9712,N_9706);
and U9821 (N_9821,N_9752,N_9609);
and U9822 (N_9822,N_9658,N_9645);
or U9823 (N_9823,N_9725,N_9675);
nor U9824 (N_9824,N_9691,N_9647);
nor U9825 (N_9825,N_9601,N_9748);
xnor U9826 (N_9826,N_9764,N_9750);
or U9827 (N_9827,N_9676,N_9742);
nand U9828 (N_9828,N_9758,N_9749);
nand U9829 (N_9829,N_9737,N_9768);
nor U9830 (N_9830,N_9704,N_9718);
nor U9831 (N_9831,N_9727,N_9785);
nand U9832 (N_9832,N_9659,N_9799);
nor U9833 (N_9833,N_9611,N_9714);
and U9834 (N_9834,N_9787,N_9782);
and U9835 (N_9835,N_9700,N_9757);
and U9836 (N_9836,N_9604,N_9733);
xor U9837 (N_9837,N_9784,N_9720);
nor U9838 (N_9838,N_9672,N_9600);
nand U9839 (N_9839,N_9716,N_9777);
or U9840 (N_9840,N_9797,N_9603);
or U9841 (N_9841,N_9724,N_9641);
or U9842 (N_9842,N_9634,N_9686);
nand U9843 (N_9843,N_9668,N_9650);
or U9844 (N_9844,N_9667,N_9674);
nand U9845 (N_9845,N_9638,N_9701);
and U9846 (N_9846,N_9736,N_9662);
nand U9847 (N_9847,N_9759,N_9660);
and U9848 (N_9848,N_9699,N_9734);
and U9849 (N_9849,N_9703,N_9633);
nand U9850 (N_9850,N_9707,N_9669);
or U9851 (N_9851,N_9637,N_9666);
nand U9852 (N_9852,N_9610,N_9754);
nand U9853 (N_9853,N_9702,N_9624);
or U9854 (N_9854,N_9747,N_9627);
xor U9855 (N_9855,N_9673,N_9670);
and U9856 (N_9856,N_9605,N_9717);
nor U9857 (N_9857,N_9786,N_9708);
xor U9858 (N_9858,N_9741,N_9792);
nor U9859 (N_9859,N_9639,N_9663);
or U9860 (N_9860,N_9649,N_9678);
or U9861 (N_9861,N_9761,N_9616);
xor U9862 (N_9862,N_9753,N_9684);
nor U9863 (N_9863,N_9788,N_9765);
xor U9864 (N_9864,N_9692,N_9607);
xor U9865 (N_9865,N_9705,N_9710);
or U9866 (N_9866,N_9770,N_9612);
or U9867 (N_9867,N_9653,N_9740);
or U9868 (N_9868,N_9656,N_9632);
xnor U9869 (N_9869,N_9694,N_9721);
xnor U9870 (N_9870,N_9680,N_9762);
and U9871 (N_9871,N_9789,N_9661);
nor U9872 (N_9872,N_9746,N_9679);
nand U9873 (N_9873,N_9688,N_9728);
nor U9874 (N_9874,N_9620,N_9630);
nor U9875 (N_9875,N_9755,N_9767);
nor U9876 (N_9876,N_9617,N_9793);
and U9877 (N_9877,N_9671,N_9775);
xor U9878 (N_9878,N_9602,N_9722);
nor U9879 (N_9879,N_9618,N_9640);
nor U9880 (N_9880,N_9774,N_9614);
or U9881 (N_9881,N_9732,N_9796);
and U9882 (N_9882,N_9696,N_9791);
and U9883 (N_9883,N_9665,N_9739);
nor U9884 (N_9884,N_9790,N_9622);
xor U9885 (N_9885,N_9745,N_9628);
nor U9886 (N_9886,N_9621,N_9723);
xor U9887 (N_9887,N_9681,N_9625);
and U9888 (N_9888,N_9776,N_9763);
xor U9889 (N_9889,N_9643,N_9695);
nand U9890 (N_9890,N_9652,N_9689);
nor U9891 (N_9891,N_9779,N_9771);
or U9892 (N_9892,N_9682,N_9615);
and U9893 (N_9893,N_9685,N_9778);
or U9894 (N_9894,N_9693,N_9794);
or U9895 (N_9895,N_9766,N_9613);
nand U9896 (N_9896,N_9709,N_9711);
or U9897 (N_9897,N_9636,N_9631);
xor U9898 (N_9898,N_9697,N_9769);
nor U9899 (N_9899,N_9773,N_9626);
and U9900 (N_9900,N_9763,N_9741);
and U9901 (N_9901,N_9698,N_9734);
xor U9902 (N_9902,N_9656,N_9698);
xor U9903 (N_9903,N_9690,N_9701);
and U9904 (N_9904,N_9613,N_9775);
nand U9905 (N_9905,N_9704,N_9629);
nand U9906 (N_9906,N_9757,N_9786);
xor U9907 (N_9907,N_9677,N_9718);
nor U9908 (N_9908,N_9764,N_9620);
nor U9909 (N_9909,N_9637,N_9748);
nand U9910 (N_9910,N_9729,N_9741);
nand U9911 (N_9911,N_9601,N_9608);
xor U9912 (N_9912,N_9619,N_9701);
nand U9913 (N_9913,N_9655,N_9711);
and U9914 (N_9914,N_9632,N_9636);
or U9915 (N_9915,N_9720,N_9666);
xnor U9916 (N_9916,N_9622,N_9733);
nor U9917 (N_9917,N_9757,N_9609);
xor U9918 (N_9918,N_9668,N_9706);
and U9919 (N_9919,N_9691,N_9615);
nor U9920 (N_9920,N_9668,N_9681);
or U9921 (N_9921,N_9601,N_9640);
nand U9922 (N_9922,N_9644,N_9671);
or U9923 (N_9923,N_9627,N_9718);
and U9924 (N_9924,N_9600,N_9793);
nand U9925 (N_9925,N_9765,N_9714);
nand U9926 (N_9926,N_9741,N_9758);
nor U9927 (N_9927,N_9719,N_9615);
nor U9928 (N_9928,N_9688,N_9776);
and U9929 (N_9929,N_9640,N_9725);
nand U9930 (N_9930,N_9662,N_9764);
nand U9931 (N_9931,N_9724,N_9672);
nor U9932 (N_9932,N_9660,N_9665);
xor U9933 (N_9933,N_9652,N_9683);
nand U9934 (N_9934,N_9791,N_9654);
xor U9935 (N_9935,N_9769,N_9676);
and U9936 (N_9936,N_9795,N_9609);
or U9937 (N_9937,N_9732,N_9729);
or U9938 (N_9938,N_9642,N_9675);
xnor U9939 (N_9939,N_9685,N_9790);
nand U9940 (N_9940,N_9790,N_9778);
or U9941 (N_9941,N_9728,N_9773);
xnor U9942 (N_9942,N_9765,N_9665);
nor U9943 (N_9943,N_9600,N_9771);
nand U9944 (N_9944,N_9698,N_9768);
nand U9945 (N_9945,N_9623,N_9718);
nor U9946 (N_9946,N_9635,N_9698);
and U9947 (N_9947,N_9790,N_9735);
and U9948 (N_9948,N_9733,N_9617);
nand U9949 (N_9949,N_9786,N_9667);
or U9950 (N_9950,N_9789,N_9606);
xnor U9951 (N_9951,N_9716,N_9738);
xnor U9952 (N_9952,N_9775,N_9790);
and U9953 (N_9953,N_9724,N_9719);
nor U9954 (N_9954,N_9789,N_9623);
xnor U9955 (N_9955,N_9633,N_9665);
and U9956 (N_9956,N_9692,N_9638);
and U9957 (N_9957,N_9757,N_9731);
nor U9958 (N_9958,N_9713,N_9767);
or U9959 (N_9959,N_9646,N_9708);
nor U9960 (N_9960,N_9735,N_9648);
xor U9961 (N_9961,N_9730,N_9763);
and U9962 (N_9962,N_9635,N_9654);
nand U9963 (N_9963,N_9613,N_9770);
xor U9964 (N_9964,N_9687,N_9782);
xor U9965 (N_9965,N_9737,N_9711);
xnor U9966 (N_9966,N_9625,N_9758);
nor U9967 (N_9967,N_9753,N_9666);
and U9968 (N_9968,N_9669,N_9688);
and U9969 (N_9969,N_9707,N_9677);
and U9970 (N_9970,N_9628,N_9732);
nand U9971 (N_9971,N_9612,N_9614);
nor U9972 (N_9972,N_9611,N_9710);
nor U9973 (N_9973,N_9757,N_9621);
nand U9974 (N_9974,N_9651,N_9715);
xnor U9975 (N_9975,N_9798,N_9791);
xor U9976 (N_9976,N_9603,N_9745);
or U9977 (N_9977,N_9776,N_9640);
or U9978 (N_9978,N_9637,N_9732);
nor U9979 (N_9979,N_9706,N_9620);
or U9980 (N_9980,N_9653,N_9706);
nor U9981 (N_9981,N_9750,N_9636);
nor U9982 (N_9982,N_9663,N_9761);
or U9983 (N_9983,N_9692,N_9627);
xor U9984 (N_9984,N_9604,N_9656);
or U9985 (N_9985,N_9708,N_9763);
nand U9986 (N_9986,N_9709,N_9790);
xnor U9987 (N_9987,N_9677,N_9722);
nand U9988 (N_9988,N_9796,N_9695);
nor U9989 (N_9989,N_9652,N_9732);
nor U9990 (N_9990,N_9680,N_9798);
nand U9991 (N_9991,N_9759,N_9798);
xor U9992 (N_9992,N_9729,N_9611);
nand U9993 (N_9993,N_9728,N_9636);
and U9994 (N_9994,N_9728,N_9615);
or U9995 (N_9995,N_9657,N_9680);
nor U9996 (N_9996,N_9664,N_9770);
nor U9997 (N_9997,N_9685,N_9762);
or U9998 (N_9998,N_9749,N_9611);
nand U9999 (N_9999,N_9762,N_9677);
nor U10000 (N_10000,N_9913,N_9961);
nor U10001 (N_10001,N_9959,N_9829);
nand U10002 (N_10002,N_9933,N_9910);
xnor U10003 (N_10003,N_9946,N_9917);
or U10004 (N_10004,N_9897,N_9845);
nor U10005 (N_10005,N_9958,N_9967);
nand U10006 (N_10006,N_9823,N_9812);
nand U10007 (N_10007,N_9867,N_9802);
xor U10008 (N_10008,N_9822,N_9847);
and U10009 (N_10009,N_9854,N_9944);
and U10010 (N_10010,N_9824,N_9973);
or U10011 (N_10011,N_9962,N_9887);
xor U10012 (N_10012,N_9989,N_9844);
nor U10013 (N_10013,N_9902,N_9996);
or U10014 (N_10014,N_9805,N_9850);
and U10015 (N_10015,N_9820,N_9950);
or U10016 (N_10016,N_9993,N_9932);
and U10017 (N_10017,N_9906,N_9825);
and U10018 (N_10018,N_9857,N_9992);
and U10019 (N_10019,N_9880,N_9927);
nand U10020 (N_10020,N_9954,N_9985);
nand U10021 (N_10021,N_9856,N_9835);
or U10022 (N_10022,N_9924,N_9849);
xnor U10023 (N_10023,N_9982,N_9843);
nor U10024 (N_10024,N_9876,N_9864);
xnor U10025 (N_10025,N_9907,N_9801);
and U10026 (N_10026,N_9863,N_9813);
xnor U10027 (N_10027,N_9833,N_9859);
nor U10028 (N_10028,N_9821,N_9804);
and U10029 (N_10029,N_9874,N_9817);
xor U10030 (N_10030,N_9869,N_9925);
nand U10031 (N_10031,N_9826,N_9838);
nand U10032 (N_10032,N_9896,N_9800);
or U10033 (N_10033,N_9828,N_9872);
or U10034 (N_10034,N_9885,N_9990);
and U10035 (N_10035,N_9977,N_9891);
nor U10036 (N_10036,N_9810,N_9834);
or U10037 (N_10037,N_9991,N_9939);
or U10038 (N_10038,N_9818,N_9928);
and U10039 (N_10039,N_9986,N_9968);
xor U10040 (N_10040,N_9807,N_9851);
xnor U10041 (N_10041,N_9949,N_9893);
or U10042 (N_10042,N_9918,N_9905);
and U10043 (N_10043,N_9846,N_9997);
and U10044 (N_10044,N_9920,N_9951);
or U10045 (N_10045,N_9900,N_9930);
and U10046 (N_10046,N_9979,N_9976);
nor U10047 (N_10047,N_9839,N_9811);
or U10048 (N_10048,N_9937,N_9981);
or U10049 (N_10049,N_9943,N_9965);
xnor U10050 (N_10050,N_9945,N_9929);
and U10051 (N_10051,N_9914,N_9858);
xnor U10052 (N_10052,N_9842,N_9878);
or U10053 (N_10053,N_9974,N_9888);
or U10054 (N_10054,N_9827,N_9879);
nor U10055 (N_10055,N_9971,N_9957);
nand U10056 (N_10056,N_9892,N_9916);
or U10057 (N_10057,N_9919,N_9923);
and U10058 (N_10058,N_9899,N_9983);
or U10059 (N_10059,N_9809,N_9941);
nor U10060 (N_10060,N_9832,N_9865);
nand U10061 (N_10061,N_9862,N_9921);
and U10062 (N_10062,N_9988,N_9963);
or U10063 (N_10063,N_9819,N_9815);
xnor U10064 (N_10064,N_9966,N_9912);
and U10065 (N_10065,N_9980,N_9938);
nor U10066 (N_10066,N_9908,N_9806);
and U10067 (N_10067,N_9909,N_9956);
xor U10068 (N_10068,N_9931,N_9873);
and U10069 (N_10069,N_9948,N_9868);
and U10070 (N_10070,N_9972,N_9934);
and U10071 (N_10071,N_9895,N_9884);
or U10072 (N_10072,N_9881,N_9875);
nand U10073 (N_10073,N_9853,N_9898);
nor U10074 (N_10074,N_9855,N_9890);
or U10075 (N_10075,N_9969,N_9830);
or U10076 (N_10076,N_9975,N_9964);
nor U10077 (N_10077,N_9882,N_9852);
xor U10078 (N_10078,N_9994,N_9970);
nand U10079 (N_10079,N_9952,N_9883);
nor U10080 (N_10080,N_9942,N_9841);
xor U10081 (N_10081,N_9936,N_9911);
and U10082 (N_10082,N_9894,N_9955);
and U10083 (N_10083,N_9886,N_9978);
nor U10084 (N_10084,N_9871,N_9960);
nor U10085 (N_10085,N_9935,N_9814);
and U10086 (N_10086,N_9998,N_9837);
nand U10087 (N_10087,N_9947,N_9870);
nor U10088 (N_10088,N_9803,N_9861);
nand U10089 (N_10089,N_9984,N_9901);
nand U10090 (N_10090,N_9860,N_9995);
and U10091 (N_10091,N_9848,N_9836);
xnor U10092 (N_10092,N_9904,N_9915);
xnor U10093 (N_10093,N_9808,N_9953);
and U10094 (N_10094,N_9840,N_9922);
nor U10095 (N_10095,N_9999,N_9926);
nor U10096 (N_10096,N_9903,N_9940);
and U10097 (N_10097,N_9816,N_9866);
or U10098 (N_10098,N_9987,N_9877);
nand U10099 (N_10099,N_9831,N_9889);
and U10100 (N_10100,N_9814,N_9911);
and U10101 (N_10101,N_9863,N_9897);
nand U10102 (N_10102,N_9871,N_9854);
xor U10103 (N_10103,N_9867,N_9959);
xnor U10104 (N_10104,N_9905,N_9912);
or U10105 (N_10105,N_9953,N_9892);
and U10106 (N_10106,N_9805,N_9905);
xnor U10107 (N_10107,N_9832,N_9989);
nor U10108 (N_10108,N_9808,N_9862);
nand U10109 (N_10109,N_9822,N_9821);
xor U10110 (N_10110,N_9808,N_9897);
nand U10111 (N_10111,N_9899,N_9868);
nor U10112 (N_10112,N_9949,N_9865);
nor U10113 (N_10113,N_9855,N_9869);
and U10114 (N_10114,N_9951,N_9875);
or U10115 (N_10115,N_9871,N_9967);
xnor U10116 (N_10116,N_9865,N_9909);
xnor U10117 (N_10117,N_9913,N_9858);
and U10118 (N_10118,N_9986,N_9864);
xor U10119 (N_10119,N_9915,N_9838);
nor U10120 (N_10120,N_9890,N_9943);
nand U10121 (N_10121,N_9877,N_9893);
nor U10122 (N_10122,N_9936,N_9927);
and U10123 (N_10123,N_9800,N_9929);
nor U10124 (N_10124,N_9800,N_9895);
and U10125 (N_10125,N_9892,N_9942);
nand U10126 (N_10126,N_9959,N_9860);
xnor U10127 (N_10127,N_9970,N_9977);
xor U10128 (N_10128,N_9914,N_9906);
or U10129 (N_10129,N_9984,N_9809);
and U10130 (N_10130,N_9988,N_9899);
nand U10131 (N_10131,N_9862,N_9856);
or U10132 (N_10132,N_9876,N_9860);
xor U10133 (N_10133,N_9825,N_9876);
and U10134 (N_10134,N_9836,N_9969);
or U10135 (N_10135,N_9907,N_9936);
nand U10136 (N_10136,N_9976,N_9814);
xor U10137 (N_10137,N_9995,N_9846);
nand U10138 (N_10138,N_9970,N_9895);
nor U10139 (N_10139,N_9872,N_9881);
or U10140 (N_10140,N_9828,N_9978);
or U10141 (N_10141,N_9822,N_9930);
nor U10142 (N_10142,N_9868,N_9965);
and U10143 (N_10143,N_9959,N_9957);
nor U10144 (N_10144,N_9842,N_9938);
nor U10145 (N_10145,N_9942,N_9872);
and U10146 (N_10146,N_9841,N_9983);
nand U10147 (N_10147,N_9986,N_9972);
nor U10148 (N_10148,N_9975,N_9978);
nor U10149 (N_10149,N_9876,N_9829);
xor U10150 (N_10150,N_9971,N_9989);
and U10151 (N_10151,N_9963,N_9853);
xnor U10152 (N_10152,N_9890,N_9882);
xnor U10153 (N_10153,N_9834,N_9875);
and U10154 (N_10154,N_9902,N_9930);
or U10155 (N_10155,N_9802,N_9992);
nor U10156 (N_10156,N_9878,N_9801);
nor U10157 (N_10157,N_9844,N_9920);
nor U10158 (N_10158,N_9920,N_9831);
or U10159 (N_10159,N_9997,N_9835);
and U10160 (N_10160,N_9933,N_9841);
nand U10161 (N_10161,N_9969,N_9880);
or U10162 (N_10162,N_9841,N_9830);
and U10163 (N_10163,N_9861,N_9898);
nand U10164 (N_10164,N_9877,N_9965);
nand U10165 (N_10165,N_9924,N_9847);
nor U10166 (N_10166,N_9866,N_9890);
and U10167 (N_10167,N_9842,N_9836);
or U10168 (N_10168,N_9991,N_9909);
and U10169 (N_10169,N_9837,N_9991);
and U10170 (N_10170,N_9846,N_9880);
xor U10171 (N_10171,N_9965,N_9878);
nor U10172 (N_10172,N_9863,N_9861);
xor U10173 (N_10173,N_9982,N_9801);
and U10174 (N_10174,N_9820,N_9969);
and U10175 (N_10175,N_9933,N_9977);
or U10176 (N_10176,N_9900,N_9884);
or U10177 (N_10177,N_9988,N_9835);
nor U10178 (N_10178,N_9849,N_9923);
nor U10179 (N_10179,N_9855,N_9984);
xnor U10180 (N_10180,N_9883,N_9897);
nor U10181 (N_10181,N_9952,N_9937);
or U10182 (N_10182,N_9893,N_9848);
xnor U10183 (N_10183,N_9872,N_9805);
xor U10184 (N_10184,N_9994,N_9974);
nand U10185 (N_10185,N_9971,N_9840);
xnor U10186 (N_10186,N_9805,N_9950);
xor U10187 (N_10187,N_9886,N_9931);
or U10188 (N_10188,N_9870,N_9978);
nand U10189 (N_10189,N_9915,N_9962);
nor U10190 (N_10190,N_9913,N_9830);
nand U10191 (N_10191,N_9970,N_9987);
xnor U10192 (N_10192,N_9878,N_9955);
nor U10193 (N_10193,N_9819,N_9973);
nor U10194 (N_10194,N_9934,N_9909);
or U10195 (N_10195,N_9894,N_9898);
nand U10196 (N_10196,N_9964,N_9930);
nor U10197 (N_10197,N_9876,N_9852);
nand U10198 (N_10198,N_9986,N_9996);
nor U10199 (N_10199,N_9828,N_9863);
xor U10200 (N_10200,N_10062,N_10195);
nor U10201 (N_10201,N_10045,N_10012);
or U10202 (N_10202,N_10050,N_10154);
nand U10203 (N_10203,N_10022,N_10165);
nand U10204 (N_10204,N_10097,N_10034);
xnor U10205 (N_10205,N_10115,N_10018);
nor U10206 (N_10206,N_10094,N_10085);
nand U10207 (N_10207,N_10046,N_10168);
and U10208 (N_10208,N_10116,N_10148);
xnor U10209 (N_10209,N_10127,N_10100);
nand U10210 (N_10210,N_10157,N_10003);
nor U10211 (N_10211,N_10030,N_10029);
and U10212 (N_10212,N_10074,N_10111);
xor U10213 (N_10213,N_10072,N_10130);
xor U10214 (N_10214,N_10042,N_10175);
nand U10215 (N_10215,N_10199,N_10019);
and U10216 (N_10216,N_10088,N_10119);
nor U10217 (N_10217,N_10176,N_10112);
nand U10218 (N_10218,N_10010,N_10169);
xor U10219 (N_10219,N_10193,N_10166);
or U10220 (N_10220,N_10044,N_10011);
nor U10221 (N_10221,N_10114,N_10006);
nor U10222 (N_10222,N_10126,N_10043);
and U10223 (N_10223,N_10180,N_10109);
xnor U10224 (N_10224,N_10086,N_10108);
nand U10225 (N_10225,N_10122,N_10078);
nand U10226 (N_10226,N_10136,N_10143);
nand U10227 (N_10227,N_10053,N_10016);
and U10228 (N_10228,N_10151,N_10039);
and U10229 (N_10229,N_10027,N_10170);
or U10230 (N_10230,N_10144,N_10020);
nor U10231 (N_10231,N_10129,N_10141);
nand U10232 (N_10232,N_10099,N_10061);
nand U10233 (N_10233,N_10041,N_10051);
nor U10234 (N_10234,N_10096,N_10083);
and U10235 (N_10235,N_10178,N_10118);
or U10236 (N_10236,N_10171,N_10007);
and U10237 (N_10237,N_10000,N_10159);
nor U10238 (N_10238,N_10002,N_10117);
nand U10239 (N_10239,N_10156,N_10190);
nor U10240 (N_10240,N_10080,N_10005);
xnor U10241 (N_10241,N_10052,N_10067);
and U10242 (N_10242,N_10155,N_10025);
and U10243 (N_10243,N_10132,N_10084);
nand U10244 (N_10244,N_10182,N_10128);
or U10245 (N_10245,N_10107,N_10037);
xnor U10246 (N_10246,N_10172,N_10149);
and U10247 (N_10247,N_10120,N_10070);
and U10248 (N_10248,N_10123,N_10137);
and U10249 (N_10249,N_10063,N_10160);
and U10250 (N_10250,N_10113,N_10060);
nor U10251 (N_10251,N_10140,N_10092);
xor U10252 (N_10252,N_10054,N_10163);
xor U10253 (N_10253,N_10057,N_10174);
nand U10254 (N_10254,N_10152,N_10153);
nor U10255 (N_10255,N_10075,N_10145);
nand U10256 (N_10256,N_10133,N_10077);
nor U10257 (N_10257,N_10104,N_10004);
xnor U10258 (N_10258,N_10031,N_10071);
and U10259 (N_10259,N_10049,N_10023);
and U10260 (N_10260,N_10150,N_10017);
nand U10261 (N_10261,N_10191,N_10142);
nand U10262 (N_10262,N_10135,N_10179);
or U10263 (N_10263,N_10095,N_10001);
xor U10264 (N_10264,N_10008,N_10105);
nand U10265 (N_10265,N_10093,N_10134);
nand U10266 (N_10266,N_10158,N_10181);
or U10267 (N_10267,N_10059,N_10032);
nand U10268 (N_10268,N_10089,N_10058);
xnor U10269 (N_10269,N_10103,N_10047);
and U10270 (N_10270,N_10079,N_10147);
nor U10271 (N_10271,N_10040,N_10087);
nor U10272 (N_10272,N_10066,N_10167);
or U10273 (N_10273,N_10125,N_10069);
and U10274 (N_10274,N_10186,N_10021);
and U10275 (N_10275,N_10161,N_10194);
or U10276 (N_10276,N_10121,N_10015);
nand U10277 (N_10277,N_10081,N_10068);
or U10278 (N_10278,N_10014,N_10173);
or U10279 (N_10279,N_10184,N_10091);
xnor U10280 (N_10280,N_10102,N_10183);
or U10281 (N_10281,N_10065,N_10038);
or U10282 (N_10282,N_10090,N_10187);
nor U10283 (N_10283,N_10131,N_10036);
nand U10284 (N_10284,N_10188,N_10138);
nor U10285 (N_10285,N_10177,N_10013);
or U10286 (N_10286,N_10189,N_10028);
xnor U10287 (N_10287,N_10196,N_10192);
and U10288 (N_10288,N_10076,N_10164);
nor U10289 (N_10289,N_10146,N_10024);
or U10290 (N_10290,N_10033,N_10035);
xnor U10291 (N_10291,N_10110,N_10056);
xor U10292 (N_10292,N_10197,N_10098);
and U10293 (N_10293,N_10064,N_10082);
nor U10294 (N_10294,N_10073,N_10198);
and U10295 (N_10295,N_10101,N_10185);
nor U10296 (N_10296,N_10124,N_10048);
xnor U10297 (N_10297,N_10106,N_10162);
and U10298 (N_10298,N_10139,N_10055);
or U10299 (N_10299,N_10026,N_10009);
and U10300 (N_10300,N_10083,N_10029);
nand U10301 (N_10301,N_10188,N_10082);
or U10302 (N_10302,N_10011,N_10092);
nand U10303 (N_10303,N_10003,N_10017);
nand U10304 (N_10304,N_10046,N_10063);
and U10305 (N_10305,N_10039,N_10077);
and U10306 (N_10306,N_10195,N_10084);
or U10307 (N_10307,N_10135,N_10172);
or U10308 (N_10308,N_10191,N_10075);
and U10309 (N_10309,N_10029,N_10129);
xor U10310 (N_10310,N_10012,N_10019);
or U10311 (N_10311,N_10025,N_10187);
nor U10312 (N_10312,N_10037,N_10083);
or U10313 (N_10313,N_10142,N_10043);
nor U10314 (N_10314,N_10134,N_10118);
nand U10315 (N_10315,N_10133,N_10003);
and U10316 (N_10316,N_10044,N_10131);
or U10317 (N_10317,N_10094,N_10112);
xnor U10318 (N_10318,N_10179,N_10046);
and U10319 (N_10319,N_10026,N_10085);
xnor U10320 (N_10320,N_10087,N_10181);
nand U10321 (N_10321,N_10176,N_10089);
nand U10322 (N_10322,N_10168,N_10054);
xor U10323 (N_10323,N_10117,N_10133);
nand U10324 (N_10324,N_10151,N_10009);
or U10325 (N_10325,N_10013,N_10066);
nor U10326 (N_10326,N_10025,N_10169);
nor U10327 (N_10327,N_10013,N_10114);
nand U10328 (N_10328,N_10099,N_10039);
xnor U10329 (N_10329,N_10042,N_10079);
and U10330 (N_10330,N_10003,N_10172);
nor U10331 (N_10331,N_10089,N_10025);
xor U10332 (N_10332,N_10146,N_10066);
xor U10333 (N_10333,N_10164,N_10044);
or U10334 (N_10334,N_10039,N_10182);
xor U10335 (N_10335,N_10170,N_10114);
or U10336 (N_10336,N_10150,N_10068);
or U10337 (N_10337,N_10076,N_10147);
and U10338 (N_10338,N_10146,N_10070);
nor U10339 (N_10339,N_10021,N_10047);
xor U10340 (N_10340,N_10051,N_10163);
nor U10341 (N_10341,N_10120,N_10141);
and U10342 (N_10342,N_10079,N_10002);
nand U10343 (N_10343,N_10083,N_10177);
nor U10344 (N_10344,N_10023,N_10130);
nand U10345 (N_10345,N_10038,N_10000);
and U10346 (N_10346,N_10121,N_10159);
nand U10347 (N_10347,N_10169,N_10072);
and U10348 (N_10348,N_10092,N_10045);
and U10349 (N_10349,N_10171,N_10181);
nor U10350 (N_10350,N_10136,N_10146);
or U10351 (N_10351,N_10086,N_10087);
xnor U10352 (N_10352,N_10181,N_10157);
xor U10353 (N_10353,N_10193,N_10001);
or U10354 (N_10354,N_10172,N_10173);
nor U10355 (N_10355,N_10086,N_10081);
nand U10356 (N_10356,N_10177,N_10173);
nor U10357 (N_10357,N_10156,N_10077);
xnor U10358 (N_10358,N_10120,N_10079);
and U10359 (N_10359,N_10168,N_10136);
nor U10360 (N_10360,N_10062,N_10070);
or U10361 (N_10361,N_10155,N_10040);
nor U10362 (N_10362,N_10066,N_10089);
and U10363 (N_10363,N_10042,N_10199);
xnor U10364 (N_10364,N_10116,N_10067);
and U10365 (N_10365,N_10057,N_10112);
and U10366 (N_10366,N_10164,N_10062);
and U10367 (N_10367,N_10084,N_10004);
nor U10368 (N_10368,N_10107,N_10022);
nor U10369 (N_10369,N_10085,N_10141);
nor U10370 (N_10370,N_10171,N_10070);
nand U10371 (N_10371,N_10041,N_10017);
nand U10372 (N_10372,N_10135,N_10187);
xnor U10373 (N_10373,N_10119,N_10170);
xor U10374 (N_10374,N_10044,N_10088);
nor U10375 (N_10375,N_10059,N_10045);
or U10376 (N_10376,N_10019,N_10059);
nand U10377 (N_10377,N_10027,N_10129);
xor U10378 (N_10378,N_10167,N_10033);
nand U10379 (N_10379,N_10064,N_10071);
or U10380 (N_10380,N_10014,N_10132);
nand U10381 (N_10381,N_10023,N_10005);
and U10382 (N_10382,N_10054,N_10108);
nor U10383 (N_10383,N_10000,N_10098);
or U10384 (N_10384,N_10029,N_10073);
xnor U10385 (N_10385,N_10109,N_10107);
nor U10386 (N_10386,N_10046,N_10008);
nand U10387 (N_10387,N_10136,N_10044);
and U10388 (N_10388,N_10026,N_10024);
nor U10389 (N_10389,N_10147,N_10196);
nand U10390 (N_10390,N_10038,N_10197);
or U10391 (N_10391,N_10135,N_10092);
xnor U10392 (N_10392,N_10085,N_10048);
nand U10393 (N_10393,N_10154,N_10169);
nor U10394 (N_10394,N_10092,N_10164);
or U10395 (N_10395,N_10173,N_10133);
nor U10396 (N_10396,N_10193,N_10070);
nor U10397 (N_10397,N_10011,N_10053);
or U10398 (N_10398,N_10198,N_10133);
nand U10399 (N_10399,N_10043,N_10049);
or U10400 (N_10400,N_10209,N_10230);
and U10401 (N_10401,N_10325,N_10212);
nor U10402 (N_10402,N_10345,N_10321);
xor U10403 (N_10403,N_10259,N_10221);
xor U10404 (N_10404,N_10295,N_10237);
nor U10405 (N_10405,N_10205,N_10225);
nor U10406 (N_10406,N_10231,N_10215);
xnor U10407 (N_10407,N_10355,N_10365);
or U10408 (N_10408,N_10396,N_10353);
nand U10409 (N_10409,N_10222,N_10398);
nor U10410 (N_10410,N_10323,N_10393);
xor U10411 (N_10411,N_10354,N_10287);
or U10412 (N_10412,N_10367,N_10236);
nor U10413 (N_10413,N_10256,N_10343);
nand U10414 (N_10414,N_10245,N_10272);
nand U10415 (N_10415,N_10238,N_10361);
nor U10416 (N_10416,N_10213,N_10313);
nor U10417 (N_10417,N_10327,N_10282);
xor U10418 (N_10418,N_10303,N_10244);
xor U10419 (N_10419,N_10386,N_10369);
and U10420 (N_10420,N_10219,N_10232);
xnor U10421 (N_10421,N_10218,N_10372);
nand U10422 (N_10422,N_10246,N_10376);
nor U10423 (N_10423,N_10357,N_10381);
or U10424 (N_10424,N_10336,N_10378);
nand U10425 (N_10425,N_10252,N_10302);
nor U10426 (N_10426,N_10203,N_10360);
nand U10427 (N_10427,N_10375,N_10342);
xor U10428 (N_10428,N_10242,N_10359);
and U10429 (N_10429,N_10391,N_10351);
nor U10430 (N_10430,N_10294,N_10285);
or U10431 (N_10431,N_10379,N_10208);
and U10432 (N_10432,N_10250,N_10216);
nor U10433 (N_10433,N_10362,N_10358);
or U10434 (N_10434,N_10317,N_10395);
nor U10435 (N_10435,N_10383,N_10331);
and U10436 (N_10436,N_10257,N_10234);
nor U10437 (N_10437,N_10322,N_10276);
or U10438 (N_10438,N_10266,N_10364);
nand U10439 (N_10439,N_10394,N_10271);
or U10440 (N_10440,N_10243,N_10201);
nor U10441 (N_10441,N_10377,N_10228);
nor U10442 (N_10442,N_10339,N_10350);
nand U10443 (N_10443,N_10348,N_10333);
nand U10444 (N_10444,N_10253,N_10286);
nand U10445 (N_10445,N_10263,N_10204);
and U10446 (N_10446,N_10278,N_10281);
nand U10447 (N_10447,N_10368,N_10399);
nor U10448 (N_10448,N_10206,N_10288);
and U10449 (N_10449,N_10308,N_10300);
nor U10450 (N_10450,N_10279,N_10289);
nand U10451 (N_10451,N_10283,N_10214);
or U10452 (N_10452,N_10249,N_10389);
nand U10453 (N_10453,N_10335,N_10385);
nor U10454 (N_10454,N_10258,N_10284);
and U10455 (N_10455,N_10247,N_10319);
xor U10456 (N_10456,N_10304,N_10223);
and U10457 (N_10457,N_10370,N_10312);
or U10458 (N_10458,N_10280,N_10380);
xnor U10459 (N_10459,N_10233,N_10324);
or U10460 (N_10460,N_10261,N_10207);
nand U10461 (N_10461,N_10305,N_10384);
nor U10462 (N_10462,N_10311,N_10291);
nand U10463 (N_10463,N_10292,N_10346);
xnor U10464 (N_10464,N_10307,N_10248);
or U10465 (N_10465,N_10224,N_10290);
or U10466 (N_10466,N_10217,N_10226);
xor U10467 (N_10467,N_10260,N_10382);
nor U10468 (N_10468,N_10297,N_10328);
and U10469 (N_10469,N_10314,N_10344);
xnor U10470 (N_10470,N_10241,N_10306);
or U10471 (N_10471,N_10274,N_10277);
or U10472 (N_10472,N_10338,N_10388);
nand U10473 (N_10473,N_10264,N_10262);
or U10474 (N_10474,N_10373,N_10347);
nor U10475 (N_10475,N_10363,N_10371);
and U10476 (N_10476,N_10267,N_10227);
or U10477 (N_10477,N_10268,N_10390);
xor U10478 (N_10478,N_10340,N_10310);
and U10479 (N_10479,N_10293,N_10273);
nor U10480 (N_10480,N_10254,N_10330);
xor U10481 (N_10481,N_10299,N_10269);
nand U10482 (N_10482,N_10397,N_10210);
xnor U10483 (N_10483,N_10309,N_10200);
nand U10484 (N_10484,N_10298,N_10265);
nand U10485 (N_10485,N_10320,N_10202);
and U10486 (N_10486,N_10270,N_10240);
nand U10487 (N_10487,N_10352,N_10334);
nand U10488 (N_10488,N_10220,N_10211);
xor U10489 (N_10489,N_10337,N_10349);
nand U10490 (N_10490,N_10235,N_10251);
or U10491 (N_10491,N_10332,N_10255);
xnor U10492 (N_10492,N_10326,N_10392);
nand U10493 (N_10493,N_10374,N_10329);
nor U10494 (N_10494,N_10275,N_10229);
nor U10495 (N_10495,N_10296,N_10316);
or U10496 (N_10496,N_10356,N_10366);
and U10497 (N_10497,N_10341,N_10387);
and U10498 (N_10498,N_10315,N_10318);
nor U10499 (N_10499,N_10301,N_10239);
and U10500 (N_10500,N_10285,N_10283);
nor U10501 (N_10501,N_10315,N_10237);
xnor U10502 (N_10502,N_10215,N_10226);
or U10503 (N_10503,N_10331,N_10210);
and U10504 (N_10504,N_10295,N_10282);
or U10505 (N_10505,N_10352,N_10203);
nand U10506 (N_10506,N_10281,N_10218);
nand U10507 (N_10507,N_10363,N_10362);
nand U10508 (N_10508,N_10347,N_10307);
or U10509 (N_10509,N_10341,N_10389);
and U10510 (N_10510,N_10235,N_10303);
and U10511 (N_10511,N_10366,N_10376);
nand U10512 (N_10512,N_10292,N_10338);
xor U10513 (N_10513,N_10295,N_10286);
or U10514 (N_10514,N_10251,N_10232);
nor U10515 (N_10515,N_10325,N_10380);
nor U10516 (N_10516,N_10371,N_10262);
and U10517 (N_10517,N_10380,N_10233);
xor U10518 (N_10518,N_10242,N_10378);
and U10519 (N_10519,N_10384,N_10262);
and U10520 (N_10520,N_10304,N_10373);
xnor U10521 (N_10521,N_10328,N_10350);
and U10522 (N_10522,N_10220,N_10366);
xnor U10523 (N_10523,N_10239,N_10322);
xnor U10524 (N_10524,N_10380,N_10398);
or U10525 (N_10525,N_10261,N_10343);
xnor U10526 (N_10526,N_10209,N_10258);
nand U10527 (N_10527,N_10338,N_10339);
or U10528 (N_10528,N_10335,N_10315);
xor U10529 (N_10529,N_10286,N_10246);
or U10530 (N_10530,N_10331,N_10391);
xnor U10531 (N_10531,N_10271,N_10349);
nor U10532 (N_10532,N_10368,N_10322);
xnor U10533 (N_10533,N_10347,N_10394);
or U10534 (N_10534,N_10274,N_10266);
nor U10535 (N_10535,N_10397,N_10223);
nand U10536 (N_10536,N_10312,N_10397);
or U10537 (N_10537,N_10247,N_10364);
xor U10538 (N_10538,N_10299,N_10274);
nor U10539 (N_10539,N_10287,N_10333);
or U10540 (N_10540,N_10337,N_10233);
nor U10541 (N_10541,N_10305,N_10216);
or U10542 (N_10542,N_10378,N_10296);
or U10543 (N_10543,N_10398,N_10281);
xnor U10544 (N_10544,N_10337,N_10368);
or U10545 (N_10545,N_10345,N_10352);
xnor U10546 (N_10546,N_10399,N_10221);
nand U10547 (N_10547,N_10375,N_10251);
nand U10548 (N_10548,N_10399,N_10333);
and U10549 (N_10549,N_10397,N_10221);
and U10550 (N_10550,N_10335,N_10330);
or U10551 (N_10551,N_10302,N_10319);
xor U10552 (N_10552,N_10303,N_10203);
or U10553 (N_10553,N_10373,N_10258);
nand U10554 (N_10554,N_10340,N_10351);
and U10555 (N_10555,N_10226,N_10382);
nor U10556 (N_10556,N_10329,N_10304);
nand U10557 (N_10557,N_10280,N_10318);
nand U10558 (N_10558,N_10361,N_10327);
nand U10559 (N_10559,N_10276,N_10321);
nand U10560 (N_10560,N_10326,N_10381);
or U10561 (N_10561,N_10352,N_10222);
and U10562 (N_10562,N_10302,N_10357);
nor U10563 (N_10563,N_10292,N_10383);
nor U10564 (N_10564,N_10250,N_10223);
nand U10565 (N_10565,N_10241,N_10208);
nand U10566 (N_10566,N_10223,N_10293);
nor U10567 (N_10567,N_10298,N_10290);
and U10568 (N_10568,N_10223,N_10339);
and U10569 (N_10569,N_10365,N_10350);
nand U10570 (N_10570,N_10209,N_10269);
and U10571 (N_10571,N_10262,N_10279);
xor U10572 (N_10572,N_10340,N_10381);
xor U10573 (N_10573,N_10364,N_10311);
and U10574 (N_10574,N_10363,N_10380);
and U10575 (N_10575,N_10398,N_10241);
and U10576 (N_10576,N_10267,N_10321);
xor U10577 (N_10577,N_10351,N_10323);
xor U10578 (N_10578,N_10332,N_10312);
nand U10579 (N_10579,N_10235,N_10305);
nand U10580 (N_10580,N_10343,N_10219);
nand U10581 (N_10581,N_10361,N_10249);
or U10582 (N_10582,N_10289,N_10219);
or U10583 (N_10583,N_10316,N_10399);
and U10584 (N_10584,N_10349,N_10390);
xor U10585 (N_10585,N_10315,N_10200);
xor U10586 (N_10586,N_10222,N_10319);
nand U10587 (N_10587,N_10273,N_10300);
and U10588 (N_10588,N_10329,N_10319);
or U10589 (N_10589,N_10257,N_10251);
and U10590 (N_10590,N_10399,N_10350);
nand U10591 (N_10591,N_10335,N_10275);
nand U10592 (N_10592,N_10239,N_10211);
nand U10593 (N_10593,N_10297,N_10289);
xnor U10594 (N_10594,N_10370,N_10395);
or U10595 (N_10595,N_10398,N_10253);
or U10596 (N_10596,N_10348,N_10393);
xnor U10597 (N_10597,N_10338,N_10345);
nand U10598 (N_10598,N_10294,N_10366);
or U10599 (N_10599,N_10206,N_10236);
nand U10600 (N_10600,N_10414,N_10544);
nor U10601 (N_10601,N_10549,N_10518);
nand U10602 (N_10602,N_10565,N_10526);
and U10603 (N_10603,N_10491,N_10409);
or U10604 (N_10604,N_10536,N_10511);
nor U10605 (N_10605,N_10467,N_10441);
and U10606 (N_10606,N_10478,N_10475);
xnor U10607 (N_10607,N_10578,N_10451);
nor U10608 (N_10608,N_10576,N_10408);
and U10609 (N_10609,N_10422,N_10462);
and U10610 (N_10610,N_10556,N_10548);
and U10611 (N_10611,N_10599,N_10551);
nor U10612 (N_10612,N_10501,N_10519);
nand U10613 (N_10613,N_10469,N_10427);
xor U10614 (N_10614,N_10428,N_10514);
nor U10615 (N_10615,N_10577,N_10579);
and U10616 (N_10616,N_10456,N_10468);
nand U10617 (N_10617,N_10572,N_10503);
xor U10618 (N_10618,N_10465,N_10477);
nor U10619 (N_10619,N_10403,N_10575);
nand U10620 (N_10620,N_10588,N_10535);
xnor U10621 (N_10621,N_10593,N_10582);
nor U10622 (N_10622,N_10480,N_10568);
nand U10623 (N_10623,N_10446,N_10569);
and U10624 (N_10624,N_10502,N_10532);
and U10625 (N_10625,N_10585,N_10564);
nand U10626 (N_10626,N_10589,N_10436);
xnor U10627 (N_10627,N_10424,N_10531);
and U10628 (N_10628,N_10471,N_10494);
nand U10629 (N_10629,N_10557,N_10506);
xor U10630 (N_10630,N_10473,N_10584);
nand U10631 (N_10631,N_10457,N_10405);
or U10632 (N_10632,N_10543,N_10410);
or U10633 (N_10633,N_10499,N_10521);
or U10634 (N_10634,N_10484,N_10455);
or U10635 (N_10635,N_10438,N_10534);
and U10636 (N_10636,N_10442,N_10592);
nand U10637 (N_10637,N_10450,N_10474);
xnor U10638 (N_10638,N_10476,N_10523);
and U10639 (N_10639,N_10597,N_10423);
nor U10640 (N_10640,N_10520,N_10472);
and U10641 (N_10641,N_10481,N_10524);
and U10642 (N_10642,N_10586,N_10482);
xor U10643 (N_10643,N_10583,N_10574);
xor U10644 (N_10644,N_10509,N_10561);
and U10645 (N_10645,N_10522,N_10433);
nor U10646 (N_10646,N_10538,N_10537);
or U10647 (N_10647,N_10464,N_10555);
and U10648 (N_10648,N_10541,N_10547);
xnor U10649 (N_10649,N_10412,N_10525);
nand U10650 (N_10650,N_10570,N_10401);
xor U10651 (N_10651,N_10552,N_10527);
or U10652 (N_10652,N_10516,N_10554);
and U10653 (N_10653,N_10454,N_10508);
xor U10654 (N_10654,N_10425,N_10447);
and U10655 (N_10655,N_10505,N_10594);
xnor U10656 (N_10656,N_10488,N_10545);
nor U10657 (N_10657,N_10449,N_10595);
or U10658 (N_10658,N_10483,N_10504);
or U10659 (N_10659,N_10453,N_10489);
nand U10660 (N_10660,N_10573,N_10513);
xnor U10661 (N_10661,N_10459,N_10406);
and U10662 (N_10662,N_10440,N_10400);
or U10663 (N_10663,N_10435,N_10486);
xor U10664 (N_10664,N_10418,N_10515);
and U10665 (N_10665,N_10439,N_10562);
nor U10666 (N_10666,N_10540,N_10493);
nand U10667 (N_10667,N_10415,N_10458);
or U10668 (N_10668,N_10533,N_10567);
and U10669 (N_10669,N_10563,N_10426);
nor U10670 (N_10670,N_10452,N_10479);
xor U10671 (N_10671,N_10580,N_10581);
nor U10672 (N_10672,N_10445,N_10528);
nor U10673 (N_10673,N_10550,N_10546);
or U10674 (N_10674,N_10432,N_10448);
or U10675 (N_10675,N_10413,N_10490);
or U10676 (N_10676,N_10431,N_10529);
or U10677 (N_10677,N_10539,N_10417);
and U10678 (N_10678,N_10510,N_10444);
nor U10679 (N_10679,N_10487,N_10558);
or U10680 (N_10680,N_10461,N_10485);
or U10681 (N_10681,N_10591,N_10596);
or U10682 (N_10682,N_10443,N_10530);
nor U10683 (N_10683,N_10460,N_10411);
or U10684 (N_10684,N_10497,N_10429);
or U10685 (N_10685,N_10566,N_10437);
or U10686 (N_10686,N_10498,N_10542);
nand U10687 (N_10687,N_10507,N_10421);
and U10688 (N_10688,N_10407,N_10430);
nor U10689 (N_10689,N_10553,N_10571);
nor U10690 (N_10690,N_10512,N_10560);
and U10691 (N_10691,N_10559,N_10587);
or U10692 (N_10692,N_10466,N_10463);
nand U10693 (N_10693,N_10434,N_10500);
nor U10694 (N_10694,N_10420,N_10402);
or U10695 (N_10695,N_10470,N_10590);
and U10696 (N_10696,N_10419,N_10492);
or U10697 (N_10697,N_10404,N_10517);
nor U10698 (N_10698,N_10495,N_10496);
or U10699 (N_10699,N_10598,N_10416);
and U10700 (N_10700,N_10513,N_10433);
xnor U10701 (N_10701,N_10523,N_10519);
or U10702 (N_10702,N_10461,N_10496);
nor U10703 (N_10703,N_10559,N_10518);
and U10704 (N_10704,N_10448,N_10597);
nor U10705 (N_10705,N_10413,N_10598);
and U10706 (N_10706,N_10458,N_10421);
nor U10707 (N_10707,N_10591,N_10504);
nand U10708 (N_10708,N_10580,N_10420);
and U10709 (N_10709,N_10531,N_10527);
xor U10710 (N_10710,N_10564,N_10404);
and U10711 (N_10711,N_10578,N_10479);
or U10712 (N_10712,N_10462,N_10541);
or U10713 (N_10713,N_10591,N_10530);
nor U10714 (N_10714,N_10560,N_10564);
nor U10715 (N_10715,N_10417,N_10503);
xor U10716 (N_10716,N_10473,N_10409);
xor U10717 (N_10717,N_10434,N_10448);
or U10718 (N_10718,N_10476,N_10574);
nand U10719 (N_10719,N_10474,N_10523);
and U10720 (N_10720,N_10544,N_10571);
or U10721 (N_10721,N_10417,N_10472);
nor U10722 (N_10722,N_10483,N_10415);
nor U10723 (N_10723,N_10499,N_10401);
xor U10724 (N_10724,N_10444,N_10477);
nor U10725 (N_10725,N_10506,N_10412);
nand U10726 (N_10726,N_10591,N_10413);
nand U10727 (N_10727,N_10540,N_10443);
nor U10728 (N_10728,N_10450,N_10593);
and U10729 (N_10729,N_10559,N_10413);
or U10730 (N_10730,N_10559,N_10491);
and U10731 (N_10731,N_10592,N_10464);
or U10732 (N_10732,N_10472,N_10490);
and U10733 (N_10733,N_10469,N_10518);
xnor U10734 (N_10734,N_10474,N_10506);
xor U10735 (N_10735,N_10447,N_10406);
xnor U10736 (N_10736,N_10522,N_10566);
or U10737 (N_10737,N_10459,N_10446);
nand U10738 (N_10738,N_10581,N_10407);
or U10739 (N_10739,N_10483,N_10486);
nor U10740 (N_10740,N_10541,N_10539);
xor U10741 (N_10741,N_10509,N_10444);
nand U10742 (N_10742,N_10479,N_10506);
or U10743 (N_10743,N_10566,N_10428);
nand U10744 (N_10744,N_10435,N_10448);
and U10745 (N_10745,N_10587,N_10532);
xnor U10746 (N_10746,N_10546,N_10483);
nor U10747 (N_10747,N_10579,N_10435);
xnor U10748 (N_10748,N_10420,N_10407);
nor U10749 (N_10749,N_10449,N_10459);
xnor U10750 (N_10750,N_10476,N_10532);
nor U10751 (N_10751,N_10487,N_10420);
or U10752 (N_10752,N_10461,N_10444);
or U10753 (N_10753,N_10566,N_10456);
nor U10754 (N_10754,N_10576,N_10418);
nor U10755 (N_10755,N_10524,N_10419);
nor U10756 (N_10756,N_10520,N_10426);
and U10757 (N_10757,N_10458,N_10504);
or U10758 (N_10758,N_10565,N_10552);
nor U10759 (N_10759,N_10506,N_10590);
or U10760 (N_10760,N_10456,N_10482);
xnor U10761 (N_10761,N_10532,N_10496);
xor U10762 (N_10762,N_10409,N_10516);
or U10763 (N_10763,N_10560,N_10450);
nor U10764 (N_10764,N_10419,N_10534);
xnor U10765 (N_10765,N_10466,N_10567);
nand U10766 (N_10766,N_10469,N_10583);
xor U10767 (N_10767,N_10493,N_10413);
and U10768 (N_10768,N_10479,N_10464);
and U10769 (N_10769,N_10458,N_10503);
or U10770 (N_10770,N_10537,N_10509);
nor U10771 (N_10771,N_10549,N_10520);
nor U10772 (N_10772,N_10594,N_10598);
nand U10773 (N_10773,N_10475,N_10507);
nor U10774 (N_10774,N_10404,N_10494);
xnor U10775 (N_10775,N_10417,N_10546);
and U10776 (N_10776,N_10451,N_10491);
or U10777 (N_10777,N_10476,N_10595);
or U10778 (N_10778,N_10558,N_10471);
or U10779 (N_10779,N_10444,N_10441);
nor U10780 (N_10780,N_10450,N_10576);
xnor U10781 (N_10781,N_10460,N_10409);
nor U10782 (N_10782,N_10451,N_10414);
nand U10783 (N_10783,N_10463,N_10596);
and U10784 (N_10784,N_10574,N_10512);
nor U10785 (N_10785,N_10527,N_10477);
nand U10786 (N_10786,N_10430,N_10591);
and U10787 (N_10787,N_10484,N_10483);
nand U10788 (N_10788,N_10510,N_10534);
and U10789 (N_10789,N_10509,N_10402);
nor U10790 (N_10790,N_10489,N_10596);
and U10791 (N_10791,N_10599,N_10547);
or U10792 (N_10792,N_10579,N_10443);
nor U10793 (N_10793,N_10591,N_10434);
and U10794 (N_10794,N_10511,N_10558);
xor U10795 (N_10795,N_10462,N_10444);
xnor U10796 (N_10796,N_10552,N_10495);
xnor U10797 (N_10797,N_10472,N_10426);
or U10798 (N_10798,N_10564,N_10587);
nor U10799 (N_10799,N_10449,N_10531);
nand U10800 (N_10800,N_10648,N_10621);
or U10801 (N_10801,N_10763,N_10649);
and U10802 (N_10802,N_10636,N_10720);
nand U10803 (N_10803,N_10654,N_10755);
xor U10804 (N_10804,N_10782,N_10790);
xnor U10805 (N_10805,N_10799,N_10667);
xnor U10806 (N_10806,N_10639,N_10634);
nor U10807 (N_10807,N_10664,N_10607);
and U10808 (N_10808,N_10663,N_10769);
or U10809 (N_10809,N_10736,N_10652);
or U10810 (N_10810,N_10624,N_10739);
xor U10811 (N_10811,N_10622,N_10767);
xor U10812 (N_10812,N_10601,N_10689);
and U10813 (N_10813,N_10789,N_10756);
nor U10814 (N_10814,N_10781,N_10614);
xor U10815 (N_10815,N_10647,N_10665);
nor U10816 (N_10816,N_10760,N_10686);
and U10817 (N_10817,N_10632,N_10656);
or U10818 (N_10818,N_10615,N_10796);
and U10819 (N_10819,N_10683,N_10707);
or U10820 (N_10820,N_10770,N_10694);
and U10821 (N_10821,N_10714,N_10741);
and U10822 (N_10822,N_10729,N_10630);
or U10823 (N_10823,N_10719,N_10602);
nor U10824 (N_10824,N_10780,N_10620);
and U10825 (N_10825,N_10783,N_10642);
or U10826 (N_10826,N_10618,N_10604);
nand U10827 (N_10827,N_10726,N_10681);
and U10828 (N_10828,N_10645,N_10635);
and U10829 (N_10829,N_10653,N_10606);
nor U10830 (N_10830,N_10679,N_10762);
or U10831 (N_10831,N_10629,N_10685);
nand U10832 (N_10832,N_10698,N_10625);
nor U10833 (N_10833,N_10740,N_10703);
nor U10834 (N_10834,N_10699,N_10777);
nand U10835 (N_10835,N_10724,N_10785);
xnor U10836 (N_10836,N_10786,N_10771);
or U10837 (N_10837,N_10603,N_10746);
xnor U10838 (N_10838,N_10678,N_10730);
xor U10839 (N_10839,N_10745,N_10731);
xnor U10840 (N_10840,N_10710,N_10791);
or U10841 (N_10841,N_10693,N_10706);
nor U10842 (N_10842,N_10761,N_10774);
xor U10843 (N_10843,N_10704,N_10670);
nand U10844 (N_10844,N_10705,N_10619);
xor U10845 (N_10845,N_10768,N_10687);
and U10846 (N_10846,N_10600,N_10795);
nand U10847 (N_10847,N_10675,N_10709);
nand U10848 (N_10848,N_10742,N_10697);
nor U10849 (N_10849,N_10669,N_10646);
or U10850 (N_10850,N_10626,N_10775);
and U10851 (N_10851,N_10691,N_10798);
and U10852 (N_10852,N_10793,N_10671);
xnor U10853 (N_10853,N_10715,N_10613);
and U10854 (N_10854,N_10721,N_10623);
or U10855 (N_10855,N_10688,N_10605);
or U10856 (N_10856,N_10711,N_10695);
nand U10857 (N_10857,N_10788,N_10757);
or U10858 (N_10858,N_10764,N_10734);
nand U10859 (N_10859,N_10696,N_10794);
nand U10860 (N_10860,N_10651,N_10743);
xnor U10861 (N_10861,N_10758,N_10751);
and U10862 (N_10862,N_10752,N_10753);
or U10863 (N_10863,N_10690,N_10778);
nand U10864 (N_10864,N_10672,N_10765);
or U10865 (N_10865,N_10633,N_10716);
or U10866 (N_10866,N_10792,N_10702);
or U10867 (N_10867,N_10713,N_10659);
and U10868 (N_10868,N_10617,N_10676);
or U10869 (N_10869,N_10735,N_10680);
and U10870 (N_10870,N_10668,N_10737);
nand U10871 (N_10871,N_10787,N_10784);
and U10872 (N_10872,N_10744,N_10684);
and U10873 (N_10873,N_10641,N_10738);
nand U10874 (N_10874,N_10666,N_10779);
nand U10875 (N_10875,N_10749,N_10748);
xor U10876 (N_10876,N_10658,N_10611);
nor U10877 (N_10877,N_10612,N_10660);
xor U10878 (N_10878,N_10727,N_10650);
xnor U10879 (N_10879,N_10723,N_10616);
and U10880 (N_10880,N_10725,N_10627);
nand U10881 (N_10881,N_10673,N_10733);
and U10882 (N_10882,N_10638,N_10608);
xnor U10883 (N_10883,N_10750,N_10797);
or U10884 (N_10884,N_10747,N_10657);
xor U10885 (N_10885,N_10766,N_10776);
nor U10886 (N_10886,N_10772,N_10692);
and U10887 (N_10887,N_10682,N_10759);
and U10888 (N_10888,N_10674,N_10662);
nor U10889 (N_10889,N_10728,N_10773);
xor U10890 (N_10890,N_10609,N_10712);
nor U10891 (N_10891,N_10718,N_10610);
or U10892 (N_10892,N_10708,N_10628);
nor U10893 (N_10893,N_10655,N_10661);
xor U10894 (N_10894,N_10754,N_10643);
xnor U10895 (N_10895,N_10640,N_10637);
and U10896 (N_10896,N_10717,N_10701);
nand U10897 (N_10897,N_10700,N_10732);
and U10898 (N_10898,N_10677,N_10644);
nand U10899 (N_10899,N_10722,N_10631);
or U10900 (N_10900,N_10730,N_10647);
and U10901 (N_10901,N_10665,N_10640);
nand U10902 (N_10902,N_10619,N_10662);
and U10903 (N_10903,N_10655,N_10751);
nor U10904 (N_10904,N_10726,N_10747);
xnor U10905 (N_10905,N_10602,N_10733);
nand U10906 (N_10906,N_10625,N_10714);
nand U10907 (N_10907,N_10799,N_10779);
and U10908 (N_10908,N_10751,N_10719);
nand U10909 (N_10909,N_10743,N_10676);
nor U10910 (N_10910,N_10744,N_10738);
xor U10911 (N_10911,N_10668,N_10641);
or U10912 (N_10912,N_10730,N_10791);
and U10913 (N_10913,N_10781,N_10752);
or U10914 (N_10914,N_10713,N_10605);
xnor U10915 (N_10915,N_10624,N_10795);
or U10916 (N_10916,N_10643,N_10603);
and U10917 (N_10917,N_10720,N_10689);
nor U10918 (N_10918,N_10644,N_10793);
nor U10919 (N_10919,N_10616,N_10620);
nand U10920 (N_10920,N_10612,N_10740);
and U10921 (N_10921,N_10647,N_10776);
and U10922 (N_10922,N_10760,N_10673);
and U10923 (N_10923,N_10740,N_10743);
and U10924 (N_10924,N_10604,N_10742);
or U10925 (N_10925,N_10751,N_10697);
and U10926 (N_10926,N_10650,N_10710);
and U10927 (N_10927,N_10668,N_10730);
xor U10928 (N_10928,N_10677,N_10719);
nand U10929 (N_10929,N_10773,N_10625);
or U10930 (N_10930,N_10702,N_10685);
nand U10931 (N_10931,N_10799,N_10778);
nand U10932 (N_10932,N_10686,N_10782);
nand U10933 (N_10933,N_10607,N_10682);
or U10934 (N_10934,N_10758,N_10719);
nand U10935 (N_10935,N_10641,N_10736);
nor U10936 (N_10936,N_10664,N_10718);
nand U10937 (N_10937,N_10689,N_10701);
or U10938 (N_10938,N_10642,N_10663);
nand U10939 (N_10939,N_10717,N_10776);
and U10940 (N_10940,N_10664,N_10637);
nand U10941 (N_10941,N_10715,N_10747);
or U10942 (N_10942,N_10612,N_10694);
nand U10943 (N_10943,N_10711,N_10787);
nor U10944 (N_10944,N_10649,N_10744);
nand U10945 (N_10945,N_10740,N_10728);
and U10946 (N_10946,N_10665,N_10760);
nand U10947 (N_10947,N_10737,N_10716);
and U10948 (N_10948,N_10771,N_10652);
nor U10949 (N_10949,N_10613,N_10738);
nor U10950 (N_10950,N_10704,N_10655);
or U10951 (N_10951,N_10775,N_10611);
or U10952 (N_10952,N_10705,N_10678);
nand U10953 (N_10953,N_10623,N_10617);
nand U10954 (N_10954,N_10651,N_10770);
nor U10955 (N_10955,N_10676,N_10609);
nand U10956 (N_10956,N_10778,N_10759);
or U10957 (N_10957,N_10694,N_10768);
nor U10958 (N_10958,N_10682,N_10742);
or U10959 (N_10959,N_10636,N_10647);
and U10960 (N_10960,N_10665,N_10776);
nor U10961 (N_10961,N_10781,N_10665);
xor U10962 (N_10962,N_10787,N_10691);
nor U10963 (N_10963,N_10768,N_10625);
nand U10964 (N_10964,N_10728,N_10779);
or U10965 (N_10965,N_10699,N_10792);
nand U10966 (N_10966,N_10674,N_10714);
xnor U10967 (N_10967,N_10641,N_10660);
or U10968 (N_10968,N_10683,N_10793);
nor U10969 (N_10969,N_10726,N_10686);
or U10970 (N_10970,N_10747,N_10696);
xnor U10971 (N_10971,N_10606,N_10648);
or U10972 (N_10972,N_10775,N_10606);
nor U10973 (N_10973,N_10728,N_10797);
nand U10974 (N_10974,N_10670,N_10610);
or U10975 (N_10975,N_10623,N_10680);
or U10976 (N_10976,N_10674,N_10687);
xnor U10977 (N_10977,N_10702,N_10660);
and U10978 (N_10978,N_10683,N_10709);
xor U10979 (N_10979,N_10797,N_10722);
and U10980 (N_10980,N_10691,N_10632);
and U10981 (N_10981,N_10638,N_10652);
xnor U10982 (N_10982,N_10769,N_10693);
or U10983 (N_10983,N_10662,N_10745);
nand U10984 (N_10984,N_10712,N_10741);
xor U10985 (N_10985,N_10786,N_10750);
xnor U10986 (N_10986,N_10694,N_10632);
nand U10987 (N_10987,N_10694,N_10731);
nor U10988 (N_10988,N_10615,N_10606);
nor U10989 (N_10989,N_10608,N_10785);
nor U10990 (N_10990,N_10690,N_10652);
nor U10991 (N_10991,N_10669,N_10793);
nor U10992 (N_10992,N_10693,N_10798);
nor U10993 (N_10993,N_10683,N_10686);
and U10994 (N_10994,N_10739,N_10606);
or U10995 (N_10995,N_10662,N_10786);
nor U10996 (N_10996,N_10777,N_10748);
nor U10997 (N_10997,N_10731,N_10643);
nand U10998 (N_10998,N_10771,N_10625);
nor U10999 (N_10999,N_10720,N_10700);
xor U11000 (N_11000,N_10968,N_10856);
or U11001 (N_11001,N_10916,N_10833);
nor U11002 (N_11002,N_10955,N_10852);
xor U11003 (N_11003,N_10969,N_10883);
xnor U11004 (N_11004,N_10962,N_10868);
or U11005 (N_11005,N_10972,N_10908);
xor U11006 (N_11006,N_10976,N_10815);
nand U11007 (N_11007,N_10836,N_10879);
xor U11008 (N_11008,N_10846,N_10959);
xnor U11009 (N_11009,N_10975,N_10826);
xnor U11010 (N_11010,N_10803,N_10907);
or U11011 (N_11011,N_10932,N_10889);
xnor U11012 (N_11012,N_10905,N_10811);
and U11013 (N_11013,N_10812,N_10813);
nor U11014 (N_11014,N_10954,N_10913);
xnor U11015 (N_11015,N_10985,N_10970);
nor U11016 (N_11016,N_10927,N_10983);
nand U11017 (N_11017,N_10900,N_10993);
and U11018 (N_11018,N_10922,N_10834);
and U11019 (N_11019,N_10958,N_10850);
and U11020 (N_11020,N_10861,N_10947);
nor U11021 (N_11021,N_10819,N_10810);
xnor U11022 (N_11022,N_10887,N_10857);
xnor U11023 (N_11023,N_10998,N_10831);
or U11024 (N_11024,N_10820,N_10816);
and U11025 (N_11025,N_10919,N_10891);
nand U11026 (N_11026,N_10862,N_10989);
xor U11027 (N_11027,N_10904,N_10839);
xor U11028 (N_11028,N_10953,N_10931);
nor U11029 (N_11029,N_10878,N_10841);
nand U11030 (N_11030,N_10934,N_10804);
xnor U11031 (N_11031,N_10869,N_10823);
or U11032 (N_11032,N_10801,N_10926);
nand U11033 (N_11033,N_10877,N_10882);
nand U11034 (N_11034,N_10873,N_10825);
xnor U11035 (N_11035,N_10988,N_10902);
and U11036 (N_11036,N_10832,N_10898);
xnor U11037 (N_11037,N_10928,N_10827);
or U11038 (N_11038,N_10888,N_10809);
nand U11039 (N_11039,N_10837,N_10940);
and U11040 (N_11040,N_10871,N_10829);
or U11041 (N_11041,N_10897,N_10890);
nand U11042 (N_11042,N_10893,N_10909);
nor U11043 (N_11043,N_10950,N_10875);
nand U11044 (N_11044,N_10964,N_10853);
or U11045 (N_11045,N_10876,N_10965);
or U11046 (N_11046,N_10963,N_10967);
or U11047 (N_11047,N_10937,N_10992);
nand U11048 (N_11048,N_10805,N_10982);
nor U11049 (N_11049,N_10866,N_10943);
or U11050 (N_11050,N_10817,N_10848);
and U11051 (N_11051,N_10977,N_10980);
or U11052 (N_11052,N_10966,N_10997);
or U11053 (N_11053,N_10995,N_10987);
nand U11054 (N_11054,N_10899,N_10859);
and U11055 (N_11055,N_10933,N_10822);
or U11056 (N_11056,N_10806,N_10984);
and U11057 (N_11057,N_10906,N_10874);
nor U11058 (N_11058,N_10894,N_10843);
nor U11059 (N_11059,N_10979,N_10821);
nor U11060 (N_11060,N_10924,N_10895);
nor U11061 (N_11061,N_10865,N_10814);
or U11062 (N_11062,N_10918,N_10855);
nor U11063 (N_11063,N_10981,N_10892);
nand U11064 (N_11064,N_10957,N_10946);
nor U11065 (N_11065,N_10941,N_10921);
and U11066 (N_11066,N_10863,N_10880);
and U11067 (N_11067,N_10807,N_10828);
xnor U11068 (N_11068,N_10870,N_10945);
and U11069 (N_11069,N_10949,N_10838);
nor U11070 (N_11070,N_10986,N_10936);
nor U11071 (N_11071,N_10978,N_10854);
and U11072 (N_11072,N_10800,N_10991);
xnor U11073 (N_11073,N_10917,N_10844);
xnor U11074 (N_11074,N_10942,N_10872);
or U11075 (N_11075,N_10849,N_10935);
xor U11076 (N_11076,N_10994,N_10990);
nand U11077 (N_11077,N_10802,N_10851);
xnor U11078 (N_11078,N_10910,N_10901);
and U11079 (N_11079,N_10920,N_10939);
xnor U11080 (N_11080,N_10858,N_10915);
and U11081 (N_11081,N_10835,N_10808);
and U11082 (N_11082,N_10911,N_10974);
and U11083 (N_11083,N_10929,N_10999);
nand U11084 (N_11084,N_10903,N_10971);
nand U11085 (N_11085,N_10847,N_10914);
nor U11086 (N_11086,N_10860,N_10818);
xor U11087 (N_11087,N_10824,N_10881);
and U11088 (N_11088,N_10896,N_10864);
nor U11089 (N_11089,N_10845,N_10867);
or U11090 (N_11090,N_10885,N_10830);
and U11091 (N_11091,N_10912,N_10842);
xnor U11092 (N_11092,N_10840,N_10884);
or U11093 (N_11093,N_10952,N_10951);
nand U11094 (N_11094,N_10973,N_10948);
or U11095 (N_11095,N_10961,N_10886);
or U11096 (N_11096,N_10956,N_10944);
and U11097 (N_11097,N_10925,N_10960);
and U11098 (N_11098,N_10923,N_10996);
or U11099 (N_11099,N_10938,N_10930);
and U11100 (N_11100,N_10840,N_10924);
nor U11101 (N_11101,N_10805,N_10809);
or U11102 (N_11102,N_10997,N_10818);
nor U11103 (N_11103,N_10978,N_10859);
or U11104 (N_11104,N_10825,N_10940);
xnor U11105 (N_11105,N_10922,N_10935);
and U11106 (N_11106,N_10959,N_10924);
nand U11107 (N_11107,N_10835,N_10972);
nor U11108 (N_11108,N_10861,N_10945);
or U11109 (N_11109,N_10847,N_10902);
or U11110 (N_11110,N_10968,N_10902);
xnor U11111 (N_11111,N_10952,N_10840);
and U11112 (N_11112,N_10954,N_10894);
or U11113 (N_11113,N_10946,N_10818);
nand U11114 (N_11114,N_10939,N_10941);
nand U11115 (N_11115,N_10817,N_10982);
and U11116 (N_11116,N_10901,N_10840);
xor U11117 (N_11117,N_10839,N_10870);
xor U11118 (N_11118,N_10990,N_10924);
nand U11119 (N_11119,N_10828,N_10986);
nor U11120 (N_11120,N_10809,N_10900);
xor U11121 (N_11121,N_10957,N_10898);
nor U11122 (N_11122,N_10972,N_10845);
xnor U11123 (N_11123,N_10992,N_10959);
xor U11124 (N_11124,N_10857,N_10965);
nand U11125 (N_11125,N_10928,N_10864);
xor U11126 (N_11126,N_10975,N_10964);
and U11127 (N_11127,N_10871,N_10830);
and U11128 (N_11128,N_10894,N_10888);
nand U11129 (N_11129,N_10959,N_10966);
nor U11130 (N_11130,N_10980,N_10846);
or U11131 (N_11131,N_10900,N_10810);
nand U11132 (N_11132,N_10858,N_10819);
xor U11133 (N_11133,N_10810,N_10922);
nor U11134 (N_11134,N_10852,N_10865);
xnor U11135 (N_11135,N_10837,N_10806);
xnor U11136 (N_11136,N_10830,N_10926);
nor U11137 (N_11137,N_10855,N_10857);
and U11138 (N_11138,N_10884,N_10934);
xnor U11139 (N_11139,N_10894,N_10837);
and U11140 (N_11140,N_10878,N_10882);
xor U11141 (N_11141,N_10964,N_10872);
and U11142 (N_11142,N_10830,N_10813);
nor U11143 (N_11143,N_10808,N_10954);
nor U11144 (N_11144,N_10845,N_10805);
xnor U11145 (N_11145,N_10910,N_10862);
and U11146 (N_11146,N_10910,N_10938);
nand U11147 (N_11147,N_10921,N_10906);
or U11148 (N_11148,N_10952,N_10876);
nor U11149 (N_11149,N_10889,N_10814);
xor U11150 (N_11150,N_10934,N_10855);
nand U11151 (N_11151,N_10832,N_10812);
or U11152 (N_11152,N_10855,N_10825);
or U11153 (N_11153,N_10888,N_10945);
and U11154 (N_11154,N_10855,N_10858);
xnor U11155 (N_11155,N_10852,N_10961);
nor U11156 (N_11156,N_10975,N_10892);
nand U11157 (N_11157,N_10998,N_10920);
or U11158 (N_11158,N_10838,N_10979);
or U11159 (N_11159,N_10844,N_10872);
and U11160 (N_11160,N_10923,N_10836);
nor U11161 (N_11161,N_10923,N_10934);
and U11162 (N_11162,N_10881,N_10952);
nor U11163 (N_11163,N_10835,N_10813);
nand U11164 (N_11164,N_10922,N_10973);
or U11165 (N_11165,N_10921,N_10820);
xnor U11166 (N_11166,N_10867,N_10941);
and U11167 (N_11167,N_10869,N_10984);
or U11168 (N_11168,N_10858,N_10824);
or U11169 (N_11169,N_10893,N_10912);
and U11170 (N_11170,N_10956,N_10827);
nor U11171 (N_11171,N_10954,N_10908);
nor U11172 (N_11172,N_10888,N_10908);
nor U11173 (N_11173,N_10800,N_10936);
and U11174 (N_11174,N_10805,N_10993);
xor U11175 (N_11175,N_10853,N_10936);
nand U11176 (N_11176,N_10834,N_10976);
nor U11177 (N_11177,N_10816,N_10926);
xor U11178 (N_11178,N_10960,N_10962);
nand U11179 (N_11179,N_10903,N_10991);
nor U11180 (N_11180,N_10886,N_10824);
and U11181 (N_11181,N_10824,N_10815);
nor U11182 (N_11182,N_10843,N_10871);
nand U11183 (N_11183,N_10966,N_10931);
and U11184 (N_11184,N_10937,N_10885);
nand U11185 (N_11185,N_10911,N_10816);
or U11186 (N_11186,N_10851,N_10927);
nand U11187 (N_11187,N_10857,N_10802);
and U11188 (N_11188,N_10928,N_10986);
nor U11189 (N_11189,N_10995,N_10930);
and U11190 (N_11190,N_10834,N_10890);
and U11191 (N_11191,N_10826,N_10878);
nor U11192 (N_11192,N_10826,N_10828);
nor U11193 (N_11193,N_10810,N_10905);
or U11194 (N_11194,N_10956,N_10934);
nor U11195 (N_11195,N_10949,N_10983);
or U11196 (N_11196,N_10804,N_10844);
nand U11197 (N_11197,N_10807,N_10979);
and U11198 (N_11198,N_10996,N_10861);
or U11199 (N_11199,N_10936,N_10909);
and U11200 (N_11200,N_11046,N_11105);
nand U11201 (N_11201,N_11072,N_11012);
nand U11202 (N_11202,N_11066,N_11097);
nor U11203 (N_11203,N_11170,N_11190);
nor U11204 (N_11204,N_11196,N_11060);
nand U11205 (N_11205,N_11133,N_11119);
or U11206 (N_11206,N_11031,N_11120);
or U11207 (N_11207,N_11109,N_11148);
nor U11208 (N_11208,N_11082,N_11050);
and U11209 (N_11209,N_11147,N_11161);
xor U11210 (N_11210,N_11079,N_11172);
and U11211 (N_11211,N_11156,N_11108);
nor U11212 (N_11212,N_11001,N_11113);
nor U11213 (N_11213,N_11026,N_11067);
xor U11214 (N_11214,N_11064,N_11122);
xor U11215 (N_11215,N_11013,N_11096);
nor U11216 (N_11216,N_11114,N_11007);
or U11217 (N_11217,N_11041,N_11140);
or U11218 (N_11218,N_11173,N_11033);
and U11219 (N_11219,N_11131,N_11044);
nand U11220 (N_11220,N_11132,N_11169);
nand U11221 (N_11221,N_11183,N_11090);
nand U11222 (N_11222,N_11154,N_11056);
nor U11223 (N_11223,N_11010,N_11102);
and U11224 (N_11224,N_11107,N_11143);
nand U11225 (N_11225,N_11163,N_11020);
nor U11226 (N_11226,N_11125,N_11029);
or U11227 (N_11227,N_11146,N_11098);
and U11228 (N_11228,N_11141,N_11115);
nor U11229 (N_11229,N_11152,N_11058);
or U11230 (N_11230,N_11074,N_11112);
or U11231 (N_11231,N_11037,N_11083);
and U11232 (N_11232,N_11008,N_11191);
xnor U11233 (N_11233,N_11022,N_11116);
and U11234 (N_11234,N_11179,N_11198);
or U11235 (N_11235,N_11065,N_11076);
nor U11236 (N_11236,N_11104,N_11166);
and U11237 (N_11237,N_11016,N_11021);
xor U11238 (N_11238,N_11099,N_11134);
or U11239 (N_11239,N_11075,N_11027);
or U11240 (N_11240,N_11175,N_11095);
nor U11241 (N_11241,N_11164,N_11078);
nor U11242 (N_11242,N_11128,N_11151);
nor U11243 (N_11243,N_11176,N_11047);
nor U11244 (N_11244,N_11073,N_11139);
nor U11245 (N_11245,N_11126,N_11145);
xnor U11246 (N_11246,N_11087,N_11071);
and U11247 (N_11247,N_11136,N_11070);
and U11248 (N_11248,N_11043,N_11086);
or U11249 (N_11249,N_11069,N_11182);
and U11250 (N_11250,N_11181,N_11180);
nand U11251 (N_11251,N_11063,N_11085);
or U11252 (N_11252,N_11003,N_11167);
and U11253 (N_11253,N_11129,N_11011);
and U11254 (N_11254,N_11130,N_11171);
nand U11255 (N_11255,N_11036,N_11138);
nand U11256 (N_11256,N_11195,N_11035);
nor U11257 (N_11257,N_11018,N_11121);
nor U11258 (N_11258,N_11054,N_11135);
and U11259 (N_11259,N_11077,N_11009);
and U11260 (N_11260,N_11059,N_11159);
or U11261 (N_11261,N_11045,N_11028);
nand U11262 (N_11262,N_11055,N_11194);
or U11263 (N_11263,N_11184,N_11149);
xnor U11264 (N_11264,N_11038,N_11053);
nor U11265 (N_11265,N_11144,N_11101);
or U11266 (N_11266,N_11158,N_11165);
xor U11267 (N_11267,N_11040,N_11186);
nor U11268 (N_11268,N_11049,N_11032);
nor U11269 (N_11269,N_11062,N_11091);
nor U11270 (N_11270,N_11189,N_11162);
or U11271 (N_11271,N_11005,N_11025);
and U11272 (N_11272,N_11006,N_11080);
xnor U11273 (N_11273,N_11034,N_11051);
nor U11274 (N_11274,N_11185,N_11002);
nand U11275 (N_11275,N_11153,N_11142);
or U11276 (N_11276,N_11081,N_11187);
nor U11277 (N_11277,N_11017,N_11199);
or U11278 (N_11278,N_11042,N_11024);
xor U11279 (N_11279,N_11160,N_11111);
xnor U11280 (N_11280,N_11094,N_11023);
or U11281 (N_11281,N_11174,N_11019);
and U11282 (N_11282,N_11177,N_11004);
nand U11283 (N_11283,N_11068,N_11197);
and U11284 (N_11284,N_11155,N_11124);
or U11285 (N_11285,N_11084,N_11015);
nor U11286 (N_11286,N_11117,N_11093);
and U11287 (N_11287,N_11123,N_11088);
nand U11288 (N_11288,N_11118,N_11188);
nand U11289 (N_11289,N_11061,N_11052);
or U11290 (N_11290,N_11000,N_11137);
and U11291 (N_11291,N_11193,N_11100);
and U11292 (N_11292,N_11178,N_11048);
and U11293 (N_11293,N_11103,N_11030);
and U11294 (N_11294,N_11168,N_11110);
xnor U11295 (N_11295,N_11150,N_11106);
and U11296 (N_11296,N_11039,N_11127);
or U11297 (N_11297,N_11089,N_11057);
nand U11298 (N_11298,N_11157,N_11192);
nand U11299 (N_11299,N_11014,N_11092);
and U11300 (N_11300,N_11086,N_11111);
or U11301 (N_11301,N_11075,N_11149);
xor U11302 (N_11302,N_11039,N_11125);
and U11303 (N_11303,N_11052,N_11152);
nor U11304 (N_11304,N_11027,N_11199);
and U11305 (N_11305,N_11189,N_11175);
nand U11306 (N_11306,N_11134,N_11115);
nand U11307 (N_11307,N_11076,N_11103);
xnor U11308 (N_11308,N_11152,N_11181);
xnor U11309 (N_11309,N_11098,N_11063);
or U11310 (N_11310,N_11097,N_11185);
xnor U11311 (N_11311,N_11087,N_11035);
nor U11312 (N_11312,N_11117,N_11111);
nand U11313 (N_11313,N_11024,N_11182);
nor U11314 (N_11314,N_11167,N_11196);
or U11315 (N_11315,N_11028,N_11027);
or U11316 (N_11316,N_11090,N_11117);
nor U11317 (N_11317,N_11168,N_11098);
xor U11318 (N_11318,N_11175,N_11132);
nor U11319 (N_11319,N_11028,N_11148);
xnor U11320 (N_11320,N_11175,N_11082);
and U11321 (N_11321,N_11091,N_11092);
and U11322 (N_11322,N_11131,N_11030);
nand U11323 (N_11323,N_11049,N_11072);
xor U11324 (N_11324,N_11089,N_11135);
and U11325 (N_11325,N_11073,N_11143);
nand U11326 (N_11326,N_11151,N_11060);
nand U11327 (N_11327,N_11191,N_11023);
and U11328 (N_11328,N_11188,N_11060);
and U11329 (N_11329,N_11159,N_11150);
nand U11330 (N_11330,N_11083,N_11006);
and U11331 (N_11331,N_11009,N_11155);
and U11332 (N_11332,N_11109,N_11180);
and U11333 (N_11333,N_11154,N_11116);
nand U11334 (N_11334,N_11103,N_11060);
xnor U11335 (N_11335,N_11070,N_11089);
and U11336 (N_11336,N_11068,N_11072);
xor U11337 (N_11337,N_11142,N_11036);
nand U11338 (N_11338,N_11056,N_11146);
or U11339 (N_11339,N_11096,N_11065);
and U11340 (N_11340,N_11079,N_11175);
nor U11341 (N_11341,N_11006,N_11035);
nor U11342 (N_11342,N_11062,N_11111);
xor U11343 (N_11343,N_11039,N_11090);
nand U11344 (N_11344,N_11059,N_11177);
or U11345 (N_11345,N_11021,N_11012);
nor U11346 (N_11346,N_11126,N_11080);
nor U11347 (N_11347,N_11157,N_11179);
nand U11348 (N_11348,N_11093,N_11033);
xnor U11349 (N_11349,N_11185,N_11159);
nor U11350 (N_11350,N_11128,N_11162);
xnor U11351 (N_11351,N_11081,N_11018);
xor U11352 (N_11352,N_11145,N_11180);
or U11353 (N_11353,N_11032,N_11128);
nand U11354 (N_11354,N_11096,N_11014);
or U11355 (N_11355,N_11121,N_11131);
nand U11356 (N_11356,N_11056,N_11199);
nand U11357 (N_11357,N_11088,N_11125);
nand U11358 (N_11358,N_11183,N_11193);
nor U11359 (N_11359,N_11195,N_11040);
and U11360 (N_11360,N_11012,N_11114);
nand U11361 (N_11361,N_11103,N_11017);
and U11362 (N_11362,N_11097,N_11088);
nand U11363 (N_11363,N_11165,N_11136);
nor U11364 (N_11364,N_11029,N_11081);
and U11365 (N_11365,N_11063,N_11190);
or U11366 (N_11366,N_11195,N_11016);
and U11367 (N_11367,N_11130,N_11199);
xor U11368 (N_11368,N_11017,N_11100);
nor U11369 (N_11369,N_11018,N_11053);
nor U11370 (N_11370,N_11032,N_11097);
nor U11371 (N_11371,N_11025,N_11029);
and U11372 (N_11372,N_11036,N_11155);
xnor U11373 (N_11373,N_11047,N_11003);
or U11374 (N_11374,N_11001,N_11196);
nor U11375 (N_11375,N_11173,N_11197);
xnor U11376 (N_11376,N_11163,N_11126);
xor U11377 (N_11377,N_11009,N_11195);
nor U11378 (N_11378,N_11161,N_11195);
or U11379 (N_11379,N_11068,N_11002);
nand U11380 (N_11380,N_11164,N_11058);
xnor U11381 (N_11381,N_11025,N_11173);
nand U11382 (N_11382,N_11198,N_11060);
nor U11383 (N_11383,N_11025,N_11001);
nand U11384 (N_11384,N_11131,N_11149);
or U11385 (N_11385,N_11164,N_11029);
and U11386 (N_11386,N_11120,N_11142);
and U11387 (N_11387,N_11145,N_11096);
xor U11388 (N_11388,N_11075,N_11145);
nor U11389 (N_11389,N_11017,N_11048);
or U11390 (N_11390,N_11185,N_11113);
nor U11391 (N_11391,N_11197,N_11119);
nand U11392 (N_11392,N_11106,N_11182);
and U11393 (N_11393,N_11137,N_11053);
or U11394 (N_11394,N_11045,N_11114);
or U11395 (N_11395,N_11007,N_11189);
or U11396 (N_11396,N_11001,N_11006);
xor U11397 (N_11397,N_11020,N_11001);
or U11398 (N_11398,N_11150,N_11085);
nor U11399 (N_11399,N_11185,N_11163);
nor U11400 (N_11400,N_11390,N_11247);
nor U11401 (N_11401,N_11269,N_11227);
and U11402 (N_11402,N_11329,N_11298);
nor U11403 (N_11403,N_11237,N_11249);
or U11404 (N_11404,N_11305,N_11394);
or U11405 (N_11405,N_11335,N_11371);
or U11406 (N_11406,N_11250,N_11261);
and U11407 (N_11407,N_11355,N_11318);
nor U11408 (N_11408,N_11339,N_11201);
or U11409 (N_11409,N_11274,N_11268);
or U11410 (N_11410,N_11324,N_11372);
xor U11411 (N_11411,N_11223,N_11235);
xnor U11412 (N_11412,N_11386,N_11234);
xor U11413 (N_11413,N_11203,N_11286);
xnor U11414 (N_11414,N_11230,N_11218);
nand U11415 (N_11415,N_11333,N_11285);
or U11416 (N_11416,N_11356,N_11266);
or U11417 (N_11417,N_11288,N_11352);
xor U11418 (N_11418,N_11273,N_11225);
and U11419 (N_11419,N_11381,N_11232);
xnor U11420 (N_11420,N_11308,N_11222);
and U11421 (N_11421,N_11342,N_11320);
nor U11422 (N_11422,N_11217,N_11349);
xor U11423 (N_11423,N_11360,N_11287);
xor U11424 (N_11424,N_11275,N_11303);
nand U11425 (N_11425,N_11351,N_11338);
or U11426 (N_11426,N_11361,N_11379);
nor U11427 (N_11427,N_11302,N_11296);
nor U11428 (N_11428,N_11359,N_11383);
nand U11429 (N_11429,N_11211,N_11300);
nor U11430 (N_11430,N_11253,N_11280);
and U11431 (N_11431,N_11378,N_11315);
nor U11432 (N_11432,N_11215,N_11376);
nor U11433 (N_11433,N_11325,N_11370);
or U11434 (N_11434,N_11243,N_11395);
nand U11435 (N_11435,N_11317,N_11233);
nor U11436 (N_11436,N_11219,N_11337);
or U11437 (N_11437,N_11343,N_11229);
or U11438 (N_11438,N_11348,N_11241);
and U11439 (N_11439,N_11251,N_11290);
xor U11440 (N_11440,N_11366,N_11231);
nand U11441 (N_11441,N_11397,N_11264);
xnor U11442 (N_11442,N_11369,N_11392);
or U11443 (N_11443,N_11239,N_11347);
and U11444 (N_11444,N_11293,N_11362);
nor U11445 (N_11445,N_11312,N_11399);
and U11446 (N_11446,N_11255,N_11216);
xnor U11447 (N_11447,N_11226,N_11322);
or U11448 (N_11448,N_11252,N_11240);
and U11449 (N_11449,N_11334,N_11353);
nor U11450 (N_11450,N_11221,N_11284);
nand U11451 (N_11451,N_11388,N_11295);
or U11452 (N_11452,N_11301,N_11262);
nor U11453 (N_11453,N_11246,N_11248);
or U11454 (N_11454,N_11354,N_11344);
nand U11455 (N_11455,N_11330,N_11224);
nor U11456 (N_11456,N_11238,N_11358);
nor U11457 (N_11457,N_11304,N_11297);
nand U11458 (N_11458,N_11220,N_11380);
or U11459 (N_11459,N_11377,N_11236);
and U11460 (N_11460,N_11382,N_11314);
and U11461 (N_11461,N_11294,N_11389);
or U11462 (N_11462,N_11259,N_11214);
nor U11463 (N_11463,N_11345,N_11385);
or U11464 (N_11464,N_11202,N_11260);
nor U11465 (N_11465,N_11357,N_11311);
nand U11466 (N_11466,N_11336,N_11244);
nor U11467 (N_11467,N_11391,N_11256);
nand U11468 (N_11468,N_11332,N_11207);
or U11469 (N_11469,N_11374,N_11331);
nand U11470 (N_11470,N_11254,N_11212);
nor U11471 (N_11471,N_11310,N_11364);
or U11472 (N_11472,N_11306,N_11209);
nor U11473 (N_11473,N_11245,N_11276);
or U11474 (N_11474,N_11291,N_11365);
and U11475 (N_11475,N_11319,N_11278);
xor U11476 (N_11476,N_11283,N_11375);
nor U11477 (N_11477,N_11208,N_11205);
or U11478 (N_11478,N_11263,N_11373);
nor U11479 (N_11479,N_11204,N_11398);
xnor U11480 (N_11480,N_11289,N_11340);
and U11481 (N_11481,N_11309,N_11270);
xnor U11482 (N_11482,N_11321,N_11299);
or U11483 (N_11483,N_11323,N_11242);
or U11484 (N_11484,N_11326,N_11396);
xnor U11485 (N_11485,N_11200,N_11292);
or U11486 (N_11486,N_11258,N_11350);
and U11487 (N_11487,N_11281,N_11327);
nand U11488 (N_11488,N_11346,N_11282);
xnor U11489 (N_11489,N_11228,N_11213);
and U11490 (N_11490,N_11363,N_11265);
or U11491 (N_11491,N_11341,N_11384);
or U11492 (N_11492,N_11267,N_11307);
or U11493 (N_11493,N_11328,N_11393);
nor U11494 (N_11494,N_11257,N_11271);
nor U11495 (N_11495,N_11313,N_11279);
and U11496 (N_11496,N_11277,N_11387);
nand U11497 (N_11497,N_11272,N_11210);
or U11498 (N_11498,N_11368,N_11367);
xnor U11499 (N_11499,N_11316,N_11206);
or U11500 (N_11500,N_11386,N_11350);
or U11501 (N_11501,N_11244,N_11360);
nand U11502 (N_11502,N_11328,N_11360);
and U11503 (N_11503,N_11394,N_11232);
and U11504 (N_11504,N_11298,N_11372);
or U11505 (N_11505,N_11266,N_11201);
nor U11506 (N_11506,N_11311,N_11305);
or U11507 (N_11507,N_11318,N_11227);
and U11508 (N_11508,N_11388,N_11348);
xnor U11509 (N_11509,N_11226,N_11380);
and U11510 (N_11510,N_11240,N_11271);
or U11511 (N_11511,N_11224,N_11229);
nor U11512 (N_11512,N_11365,N_11393);
or U11513 (N_11513,N_11236,N_11399);
nand U11514 (N_11514,N_11338,N_11254);
nand U11515 (N_11515,N_11262,N_11268);
or U11516 (N_11516,N_11328,N_11264);
xor U11517 (N_11517,N_11275,N_11221);
or U11518 (N_11518,N_11235,N_11341);
xnor U11519 (N_11519,N_11312,N_11245);
nor U11520 (N_11520,N_11338,N_11379);
nand U11521 (N_11521,N_11224,N_11273);
or U11522 (N_11522,N_11225,N_11286);
xor U11523 (N_11523,N_11314,N_11376);
xor U11524 (N_11524,N_11239,N_11344);
and U11525 (N_11525,N_11208,N_11320);
nand U11526 (N_11526,N_11201,N_11241);
nand U11527 (N_11527,N_11351,N_11205);
xnor U11528 (N_11528,N_11340,N_11324);
xnor U11529 (N_11529,N_11319,N_11285);
nor U11530 (N_11530,N_11250,N_11216);
or U11531 (N_11531,N_11287,N_11393);
nand U11532 (N_11532,N_11391,N_11244);
nor U11533 (N_11533,N_11336,N_11392);
nor U11534 (N_11534,N_11352,N_11339);
xor U11535 (N_11535,N_11204,N_11265);
or U11536 (N_11536,N_11235,N_11399);
and U11537 (N_11537,N_11266,N_11309);
nor U11538 (N_11538,N_11362,N_11245);
xor U11539 (N_11539,N_11244,N_11341);
and U11540 (N_11540,N_11215,N_11341);
nand U11541 (N_11541,N_11398,N_11241);
or U11542 (N_11542,N_11221,N_11218);
xnor U11543 (N_11543,N_11207,N_11305);
xor U11544 (N_11544,N_11285,N_11253);
and U11545 (N_11545,N_11300,N_11392);
and U11546 (N_11546,N_11313,N_11201);
nand U11547 (N_11547,N_11321,N_11210);
or U11548 (N_11548,N_11264,N_11213);
nor U11549 (N_11549,N_11282,N_11239);
nand U11550 (N_11550,N_11377,N_11279);
or U11551 (N_11551,N_11221,N_11332);
nor U11552 (N_11552,N_11380,N_11202);
xor U11553 (N_11553,N_11206,N_11271);
nand U11554 (N_11554,N_11210,N_11305);
and U11555 (N_11555,N_11226,N_11330);
xor U11556 (N_11556,N_11275,N_11268);
nand U11557 (N_11557,N_11337,N_11315);
nor U11558 (N_11558,N_11362,N_11399);
nor U11559 (N_11559,N_11227,N_11278);
and U11560 (N_11560,N_11352,N_11397);
and U11561 (N_11561,N_11225,N_11224);
and U11562 (N_11562,N_11240,N_11305);
and U11563 (N_11563,N_11297,N_11341);
nand U11564 (N_11564,N_11397,N_11217);
and U11565 (N_11565,N_11277,N_11221);
and U11566 (N_11566,N_11331,N_11248);
nand U11567 (N_11567,N_11379,N_11356);
and U11568 (N_11568,N_11376,N_11322);
nand U11569 (N_11569,N_11376,N_11213);
nand U11570 (N_11570,N_11201,N_11203);
xor U11571 (N_11571,N_11213,N_11398);
nor U11572 (N_11572,N_11207,N_11321);
or U11573 (N_11573,N_11376,N_11241);
nand U11574 (N_11574,N_11261,N_11237);
and U11575 (N_11575,N_11371,N_11235);
nand U11576 (N_11576,N_11200,N_11217);
nor U11577 (N_11577,N_11231,N_11211);
nor U11578 (N_11578,N_11253,N_11329);
xnor U11579 (N_11579,N_11327,N_11375);
nand U11580 (N_11580,N_11350,N_11274);
or U11581 (N_11581,N_11246,N_11205);
or U11582 (N_11582,N_11314,N_11270);
nand U11583 (N_11583,N_11306,N_11349);
and U11584 (N_11584,N_11309,N_11313);
nand U11585 (N_11585,N_11314,N_11282);
or U11586 (N_11586,N_11392,N_11202);
and U11587 (N_11587,N_11370,N_11329);
and U11588 (N_11588,N_11337,N_11261);
and U11589 (N_11589,N_11343,N_11258);
or U11590 (N_11590,N_11355,N_11240);
xor U11591 (N_11591,N_11233,N_11322);
or U11592 (N_11592,N_11205,N_11229);
or U11593 (N_11593,N_11387,N_11319);
and U11594 (N_11594,N_11274,N_11238);
or U11595 (N_11595,N_11398,N_11354);
xor U11596 (N_11596,N_11253,N_11232);
nand U11597 (N_11597,N_11240,N_11319);
nor U11598 (N_11598,N_11317,N_11386);
nor U11599 (N_11599,N_11296,N_11355);
nor U11600 (N_11600,N_11510,N_11404);
or U11601 (N_11601,N_11500,N_11573);
nor U11602 (N_11602,N_11555,N_11577);
or U11603 (N_11603,N_11584,N_11596);
nor U11604 (N_11604,N_11571,N_11436);
and U11605 (N_11605,N_11502,N_11589);
xnor U11606 (N_11606,N_11591,N_11492);
or U11607 (N_11607,N_11469,N_11578);
nor U11608 (N_11608,N_11564,N_11552);
and U11609 (N_11609,N_11495,N_11534);
nor U11610 (N_11610,N_11574,N_11576);
nor U11611 (N_11611,N_11529,N_11572);
or U11612 (N_11612,N_11496,N_11583);
nor U11613 (N_11613,N_11561,N_11411);
and U11614 (N_11614,N_11454,N_11517);
xnor U11615 (N_11615,N_11483,N_11493);
or U11616 (N_11616,N_11565,N_11462);
or U11617 (N_11617,N_11476,N_11523);
nand U11618 (N_11618,N_11417,N_11463);
and U11619 (N_11619,N_11410,N_11520);
xnor U11620 (N_11620,N_11482,N_11558);
xnor U11621 (N_11621,N_11557,N_11511);
and U11622 (N_11622,N_11414,N_11499);
xor U11623 (N_11623,N_11461,N_11536);
and U11624 (N_11624,N_11453,N_11560);
or U11625 (N_11625,N_11527,N_11441);
nor U11626 (N_11626,N_11575,N_11428);
xnor U11627 (N_11627,N_11467,N_11485);
nor U11628 (N_11628,N_11458,N_11559);
nand U11629 (N_11629,N_11531,N_11480);
nor U11630 (N_11630,N_11475,N_11468);
or U11631 (N_11631,N_11408,N_11400);
xor U11632 (N_11632,N_11440,N_11450);
or U11633 (N_11633,N_11568,N_11526);
nor U11634 (N_11634,N_11556,N_11540);
and U11635 (N_11635,N_11401,N_11473);
xnor U11636 (N_11636,N_11532,N_11409);
nand U11637 (N_11637,N_11595,N_11438);
or U11638 (N_11638,N_11491,N_11427);
nand U11639 (N_11639,N_11447,N_11490);
and U11640 (N_11640,N_11581,N_11506);
nand U11641 (N_11641,N_11539,N_11533);
xnor U11642 (N_11642,N_11449,N_11509);
nand U11643 (N_11643,N_11434,N_11407);
xnor U11644 (N_11644,N_11416,N_11466);
nor U11645 (N_11645,N_11516,N_11546);
xor U11646 (N_11646,N_11478,N_11471);
nor U11647 (N_11647,N_11422,N_11569);
or U11648 (N_11648,N_11456,N_11460);
and U11649 (N_11649,N_11553,N_11443);
nor U11650 (N_11650,N_11586,N_11412);
nand U11651 (N_11651,N_11518,N_11498);
nand U11652 (N_11652,N_11423,N_11594);
and U11653 (N_11653,N_11497,N_11489);
or U11654 (N_11654,N_11514,N_11579);
nor U11655 (N_11655,N_11508,N_11542);
xor U11656 (N_11656,N_11420,N_11425);
xnor U11657 (N_11657,N_11593,N_11437);
xnor U11658 (N_11658,N_11528,N_11544);
nand U11659 (N_11659,N_11598,N_11585);
nand U11660 (N_11660,N_11548,N_11525);
nand U11661 (N_11661,N_11426,N_11570);
nand U11662 (N_11662,N_11432,N_11457);
nand U11663 (N_11663,N_11562,N_11580);
nor U11664 (N_11664,N_11535,N_11477);
xnor U11665 (N_11665,N_11501,N_11418);
or U11666 (N_11666,N_11545,N_11530);
xor U11667 (N_11667,N_11592,N_11406);
and U11668 (N_11668,N_11435,N_11403);
xnor U11669 (N_11669,N_11547,N_11419);
or U11670 (N_11670,N_11582,N_11549);
xor U11671 (N_11671,N_11599,N_11504);
or U11672 (N_11672,N_11415,N_11446);
xor U11673 (N_11673,N_11474,N_11470);
nor U11674 (N_11674,N_11486,N_11421);
or U11675 (N_11675,N_11481,N_11543);
or U11676 (N_11676,N_11524,N_11551);
nand U11677 (N_11677,N_11472,N_11494);
or U11678 (N_11678,N_11430,N_11488);
nor U11679 (N_11679,N_11465,N_11484);
nor U11680 (N_11680,N_11505,N_11567);
xnor U11681 (N_11681,N_11541,N_11515);
xnor U11682 (N_11682,N_11431,N_11455);
nor U11683 (N_11683,N_11563,N_11445);
or U11684 (N_11684,N_11402,N_11424);
or U11685 (N_11685,N_11464,N_11439);
and U11686 (N_11686,N_11487,N_11590);
nand U11687 (N_11687,N_11451,N_11442);
and U11688 (N_11688,N_11513,N_11448);
and U11689 (N_11689,N_11519,N_11479);
and U11690 (N_11690,N_11512,N_11413);
and U11691 (N_11691,N_11429,N_11444);
nand U11692 (N_11692,N_11538,N_11459);
nand U11693 (N_11693,N_11537,N_11597);
and U11694 (N_11694,N_11550,N_11587);
nor U11695 (N_11695,N_11554,N_11588);
xnor U11696 (N_11696,N_11566,N_11433);
and U11697 (N_11697,N_11521,N_11405);
and U11698 (N_11698,N_11503,N_11507);
nand U11699 (N_11699,N_11452,N_11522);
nor U11700 (N_11700,N_11407,N_11451);
nand U11701 (N_11701,N_11523,N_11462);
or U11702 (N_11702,N_11513,N_11504);
nor U11703 (N_11703,N_11587,N_11506);
xnor U11704 (N_11704,N_11463,N_11401);
or U11705 (N_11705,N_11479,N_11523);
or U11706 (N_11706,N_11558,N_11443);
or U11707 (N_11707,N_11579,N_11524);
xnor U11708 (N_11708,N_11500,N_11551);
nor U11709 (N_11709,N_11475,N_11560);
and U11710 (N_11710,N_11469,N_11551);
and U11711 (N_11711,N_11510,N_11427);
and U11712 (N_11712,N_11524,N_11501);
nand U11713 (N_11713,N_11405,N_11586);
nand U11714 (N_11714,N_11432,N_11540);
nor U11715 (N_11715,N_11455,N_11428);
and U11716 (N_11716,N_11568,N_11595);
and U11717 (N_11717,N_11404,N_11437);
nor U11718 (N_11718,N_11447,N_11580);
and U11719 (N_11719,N_11411,N_11463);
and U11720 (N_11720,N_11522,N_11565);
nand U11721 (N_11721,N_11400,N_11403);
nand U11722 (N_11722,N_11402,N_11456);
nor U11723 (N_11723,N_11488,N_11542);
xor U11724 (N_11724,N_11518,N_11447);
or U11725 (N_11725,N_11596,N_11547);
or U11726 (N_11726,N_11440,N_11495);
or U11727 (N_11727,N_11574,N_11498);
xor U11728 (N_11728,N_11400,N_11429);
and U11729 (N_11729,N_11525,N_11594);
xnor U11730 (N_11730,N_11502,N_11538);
nor U11731 (N_11731,N_11546,N_11502);
nand U11732 (N_11732,N_11589,N_11427);
nor U11733 (N_11733,N_11497,N_11413);
xor U11734 (N_11734,N_11448,N_11549);
nand U11735 (N_11735,N_11438,N_11495);
or U11736 (N_11736,N_11443,N_11557);
or U11737 (N_11737,N_11459,N_11495);
or U11738 (N_11738,N_11505,N_11475);
xnor U11739 (N_11739,N_11568,N_11580);
nor U11740 (N_11740,N_11489,N_11520);
nand U11741 (N_11741,N_11485,N_11560);
nand U11742 (N_11742,N_11587,N_11485);
or U11743 (N_11743,N_11464,N_11462);
and U11744 (N_11744,N_11564,N_11549);
and U11745 (N_11745,N_11589,N_11443);
nor U11746 (N_11746,N_11461,N_11582);
xnor U11747 (N_11747,N_11455,N_11434);
and U11748 (N_11748,N_11508,N_11579);
and U11749 (N_11749,N_11534,N_11413);
or U11750 (N_11750,N_11590,N_11561);
and U11751 (N_11751,N_11506,N_11556);
xnor U11752 (N_11752,N_11511,N_11515);
nand U11753 (N_11753,N_11465,N_11542);
nor U11754 (N_11754,N_11467,N_11526);
or U11755 (N_11755,N_11490,N_11415);
and U11756 (N_11756,N_11599,N_11499);
nand U11757 (N_11757,N_11462,N_11456);
nand U11758 (N_11758,N_11469,N_11504);
and U11759 (N_11759,N_11584,N_11413);
and U11760 (N_11760,N_11517,N_11414);
nor U11761 (N_11761,N_11473,N_11468);
and U11762 (N_11762,N_11457,N_11552);
and U11763 (N_11763,N_11466,N_11480);
xor U11764 (N_11764,N_11412,N_11425);
and U11765 (N_11765,N_11406,N_11515);
and U11766 (N_11766,N_11583,N_11565);
nand U11767 (N_11767,N_11533,N_11519);
or U11768 (N_11768,N_11585,N_11443);
nand U11769 (N_11769,N_11540,N_11477);
nand U11770 (N_11770,N_11507,N_11515);
nand U11771 (N_11771,N_11517,N_11531);
or U11772 (N_11772,N_11422,N_11522);
xor U11773 (N_11773,N_11539,N_11441);
or U11774 (N_11774,N_11436,N_11570);
xnor U11775 (N_11775,N_11536,N_11533);
nor U11776 (N_11776,N_11478,N_11416);
xor U11777 (N_11777,N_11585,N_11469);
and U11778 (N_11778,N_11523,N_11427);
or U11779 (N_11779,N_11421,N_11414);
nor U11780 (N_11780,N_11517,N_11431);
nand U11781 (N_11781,N_11481,N_11535);
and U11782 (N_11782,N_11563,N_11418);
or U11783 (N_11783,N_11447,N_11534);
nand U11784 (N_11784,N_11424,N_11538);
or U11785 (N_11785,N_11509,N_11578);
or U11786 (N_11786,N_11517,N_11548);
xnor U11787 (N_11787,N_11592,N_11488);
xor U11788 (N_11788,N_11449,N_11552);
xnor U11789 (N_11789,N_11409,N_11480);
nand U11790 (N_11790,N_11588,N_11484);
and U11791 (N_11791,N_11577,N_11500);
nand U11792 (N_11792,N_11413,N_11446);
or U11793 (N_11793,N_11540,N_11521);
nor U11794 (N_11794,N_11545,N_11438);
and U11795 (N_11795,N_11402,N_11516);
nand U11796 (N_11796,N_11416,N_11436);
nor U11797 (N_11797,N_11420,N_11401);
xor U11798 (N_11798,N_11566,N_11419);
nand U11799 (N_11799,N_11400,N_11520);
and U11800 (N_11800,N_11732,N_11636);
xor U11801 (N_11801,N_11740,N_11794);
and U11802 (N_11802,N_11643,N_11731);
nor U11803 (N_11803,N_11669,N_11640);
nor U11804 (N_11804,N_11721,N_11602);
nand U11805 (N_11805,N_11775,N_11780);
xnor U11806 (N_11806,N_11662,N_11690);
nor U11807 (N_11807,N_11663,N_11699);
nand U11808 (N_11808,N_11729,N_11768);
or U11809 (N_11809,N_11645,N_11632);
or U11810 (N_11810,N_11601,N_11655);
or U11811 (N_11811,N_11620,N_11617);
and U11812 (N_11812,N_11724,N_11784);
and U11813 (N_11813,N_11675,N_11774);
xnor U11814 (N_11814,N_11603,N_11625);
or U11815 (N_11815,N_11702,N_11735);
or U11816 (N_11816,N_11641,N_11629);
xor U11817 (N_11817,N_11665,N_11667);
or U11818 (N_11818,N_11692,N_11738);
xnor U11819 (N_11819,N_11789,N_11756);
xnor U11820 (N_11820,N_11681,N_11711);
nor U11821 (N_11821,N_11718,N_11763);
or U11822 (N_11822,N_11705,N_11610);
and U11823 (N_11823,N_11634,N_11712);
nor U11824 (N_11824,N_11693,N_11747);
nand U11825 (N_11825,N_11781,N_11799);
xnor U11826 (N_11826,N_11605,N_11737);
xor U11827 (N_11827,N_11670,N_11743);
nand U11828 (N_11828,N_11791,N_11736);
xor U11829 (N_11829,N_11679,N_11638);
and U11830 (N_11830,N_11633,N_11770);
and U11831 (N_11831,N_11639,N_11748);
or U11832 (N_11832,N_11695,N_11691);
nand U11833 (N_11833,N_11710,N_11685);
and U11834 (N_11834,N_11726,N_11611);
nand U11835 (N_11835,N_11647,N_11683);
or U11836 (N_11836,N_11709,N_11618);
nand U11837 (N_11837,N_11708,N_11720);
nor U11838 (N_11838,N_11715,N_11642);
or U11839 (N_11839,N_11630,N_11751);
and U11840 (N_11840,N_11765,N_11779);
nand U11841 (N_11841,N_11761,N_11762);
xor U11842 (N_11842,N_11644,N_11628);
and U11843 (N_11843,N_11722,N_11795);
or U11844 (N_11844,N_11658,N_11772);
or U11845 (N_11845,N_11678,N_11788);
nor U11846 (N_11846,N_11608,N_11671);
nor U11847 (N_11847,N_11619,N_11688);
and U11848 (N_11848,N_11624,N_11745);
xnor U11849 (N_11849,N_11674,N_11696);
xnor U11850 (N_11850,N_11614,N_11622);
or U11851 (N_11851,N_11769,N_11787);
nor U11852 (N_11852,N_11616,N_11753);
and U11853 (N_11853,N_11777,N_11723);
nor U11854 (N_11854,N_11700,N_11697);
nor U11855 (N_11855,N_11713,N_11728);
xor U11856 (N_11856,N_11646,N_11612);
nor U11857 (N_11857,N_11661,N_11771);
and U11858 (N_11858,N_11786,N_11698);
xor U11859 (N_11859,N_11660,N_11652);
nand U11860 (N_11860,N_11676,N_11606);
nand U11861 (N_11861,N_11657,N_11600);
nand U11862 (N_11862,N_11649,N_11635);
nor U11863 (N_11863,N_11750,N_11785);
nand U11864 (N_11864,N_11659,N_11651);
or U11865 (N_11865,N_11607,N_11746);
nor U11866 (N_11866,N_11613,N_11648);
nor U11867 (N_11867,N_11776,N_11673);
nor U11868 (N_11868,N_11714,N_11672);
xor U11869 (N_11869,N_11796,N_11666);
xnor U11870 (N_11870,N_11668,N_11704);
nor U11871 (N_11871,N_11716,N_11621);
nand U11872 (N_11872,N_11783,N_11734);
nand U11873 (N_11873,N_11653,N_11752);
or U11874 (N_11874,N_11742,N_11627);
nor U11875 (N_11875,N_11754,N_11703);
xor U11876 (N_11876,N_11733,N_11717);
or U11877 (N_11877,N_11604,N_11727);
and U11878 (N_11878,N_11792,N_11626);
or U11879 (N_11879,N_11689,N_11782);
and U11880 (N_11880,N_11760,N_11631);
nor U11881 (N_11881,N_11790,N_11759);
xnor U11882 (N_11882,N_11719,N_11764);
nand U11883 (N_11883,N_11749,N_11687);
or U11884 (N_11884,N_11741,N_11637);
or U11885 (N_11885,N_11664,N_11730);
nor U11886 (N_11886,N_11757,N_11798);
or U11887 (N_11887,N_11684,N_11773);
nor U11888 (N_11888,N_11797,N_11758);
and U11889 (N_11889,N_11654,N_11755);
or U11890 (N_11890,N_11615,N_11623);
or U11891 (N_11891,N_11677,N_11766);
and U11892 (N_11892,N_11739,N_11707);
or U11893 (N_11893,N_11744,N_11682);
or U11894 (N_11894,N_11793,N_11706);
xor U11895 (N_11895,N_11767,N_11656);
or U11896 (N_11896,N_11680,N_11694);
nand U11897 (N_11897,N_11609,N_11686);
and U11898 (N_11898,N_11725,N_11650);
xnor U11899 (N_11899,N_11778,N_11701);
nand U11900 (N_11900,N_11686,N_11674);
nand U11901 (N_11901,N_11729,N_11798);
or U11902 (N_11902,N_11744,N_11720);
nor U11903 (N_11903,N_11724,N_11688);
nor U11904 (N_11904,N_11713,N_11771);
and U11905 (N_11905,N_11700,N_11667);
xor U11906 (N_11906,N_11669,N_11795);
xor U11907 (N_11907,N_11698,N_11615);
xnor U11908 (N_11908,N_11622,N_11709);
nor U11909 (N_11909,N_11628,N_11677);
xor U11910 (N_11910,N_11609,N_11764);
nand U11911 (N_11911,N_11642,N_11609);
or U11912 (N_11912,N_11741,N_11661);
xor U11913 (N_11913,N_11744,N_11752);
nor U11914 (N_11914,N_11690,N_11629);
and U11915 (N_11915,N_11719,N_11677);
nor U11916 (N_11916,N_11794,N_11643);
or U11917 (N_11917,N_11639,N_11707);
and U11918 (N_11918,N_11617,N_11619);
nand U11919 (N_11919,N_11754,N_11730);
and U11920 (N_11920,N_11748,N_11747);
and U11921 (N_11921,N_11675,N_11657);
or U11922 (N_11922,N_11764,N_11778);
nand U11923 (N_11923,N_11784,N_11743);
and U11924 (N_11924,N_11651,N_11641);
or U11925 (N_11925,N_11746,N_11748);
nand U11926 (N_11926,N_11706,N_11782);
nand U11927 (N_11927,N_11693,N_11659);
xnor U11928 (N_11928,N_11761,N_11603);
xnor U11929 (N_11929,N_11749,N_11618);
nor U11930 (N_11930,N_11609,N_11760);
nand U11931 (N_11931,N_11689,N_11704);
or U11932 (N_11932,N_11791,N_11730);
nor U11933 (N_11933,N_11612,N_11688);
xor U11934 (N_11934,N_11638,N_11747);
xnor U11935 (N_11935,N_11675,N_11641);
xor U11936 (N_11936,N_11797,N_11779);
and U11937 (N_11937,N_11601,N_11624);
nand U11938 (N_11938,N_11689,N_11624);
nor U11939 (N_11939,N_11692,N_11769);
and U11940 (N_11940,N_11600,N_11779);
or U11941 (N_11941,N_11771,N_11775);
xnor U11942 (N_11942,N_11604,N_11797);
nand U11943 (N_11943,N_11694,N_11688);
nor U11944 (N_11944,N_11668,N_11719);
or U11945 (N_11945,N_11719,N_11699);
or U11946 (N_11946,N_11728,N_11642);
nand U11947 (N_11947,N_11737,N_11620);
xor U11948 (N_11948,N_11652,N_11641);
xnor U11949 (N_11949,N_11672,N_11737);
or U11950 (N_11950,N_11613,N_11638);
nor U11951 (N_11951,N_11729,N_11695);
nand U11952 (N_11952,N_11669,N_11723);
xor U11953 (N_11953,N_11754,N_11775);
or U11954 (N_11954,N_11783,N_11673);
nand U11955 (N_11955,N_11657,N_11756);
nand U11956 (N_11956,N_11783,N_11787);
nor U11957 (N_11957,N_11678,N_11765);
or U11958 (N_11958,N_11767,N_11625);
and U11959 (N_11959,N_11705,N_11758);
nor U11960 (N_11960,N_11726,N_11691);
and U11961 (N_11961,N_11671,N_11782);
nand U11962 (N_11962,N_11753,N_11638);
and U11963 (N_11963,N_11612,N_11625);
nand U11964 (N_11964,N_11763,N_11703);
and U11965 (N_11965,N_11671,N_11625);
nor U11966 (N_11966,N_11661,N_11731);
xnor U11967 (N_11967,N_11695,N_11636);
nand U11968 (N_11968,N_11747,N_11639);
xor U11969 (N_11969,N_11672,N_11613);
nor U11970 (N_11970,N_11643,N_11785);
xnor U11971 (N_11971,N_11627,N_11797);
and U11972 (N_11972,N_11731,N_11748);
nand U11973 (N_11973,N_11774,N_11621);
xor U11974 (N_11974,N_11767,N_11672);
nand U11975 (N_11975,N_11724,N_11757);
or U11976 (N_11976,N_11735,N_11637);
nor U11977 (N_11977,N_11789,N_11766);
nor U11978 (N_11978,N_11638,N_11666);
xor U11979 (N_11979,N_11728,N_11656);
nand U11980 (N_11980,N_11719,N_11636);
nor U11981 (N_11981,N_11615,N_11738);
or U11982 (N_11982,N_11607,N_11749);
xor U11983 (N_11983,N_11759,N_11716);
nor U11984 (N_11984,N_11698,N_11757);
nand U11985 (N_11985,N_11629,N_11618);
nor U11986 (N_11986,N_11724,N_11789);
and U11987 (N_11987,N_11654,N_11605);
and U11988 (N_11988,N_11704,N_11776);
xnor U11989 (N_11989,N_11711,N_11689);
or U11990 (N_11990,N_11761,N_11750);
nor U11991 (N_11991,N_11690,N_11781);
nor U11992 (N_11992,N_11723,N_11736);
and U11993 (N_11993,N_11627,N_11729);
xor U11994 (N_11994,N_11714,N_11646);
nand U11995 (N_11995,N_11629,N_11631);
and U11996 (N_11996,N_11749,N_11609);
nand U11997 (N_11997,N_11777,N_11665);
nand U11998 (N_11998,N_11662,N_11648);
xor U11999 (N_11999,N_11778,N_11727);
nand U12000 (N_12000,N_11809,N_11832);
xor U12001 (N_12001,N_11892,N_11982);
nand U12002 (N_12002,N_11918,N_11998);
or U12003 (N_12003,N_11807,N_11837);
xnor U12004 (N_12004,N_11945,N_11886);
xor U12005 (N_12005,N_11845,N_11992);
and U12006 (N_12006,N_11802,N_11975);
or U12007 (N_12007,N_11880,N_11820);
nor U12008 (N_12008,N_11958,N_11804);
xor U12009 (N_12009,N_11859,N_11936);
and U12010 (N_12010,N_11872,N_11888);
nand U12011 (N_12011,N_11821,N_11986);
nor U12012 (N_12012,N_11874,N_11969);
and U12013 (N_12013,N_11949,N_11974);
and U12014 (N_12014,N_11956,N_11900);
nand U12015 (N_12015,N_11873,N_11884);
nor U12016 (N_12016,N_11805,N_11984);
or U12017 (N_12017,N_11950,N_11916);
or U12018 (N_12018,N_11833,N_11902);
and U12019 (N_12019,N_11964,N_11875);
and U12020 (N_12020,N_11919,N_11861);
and U12021 (N_12021,N_11843,N_11862);
xnor U12022 (N_12022,N_11838,N_11959);
or U12023 (N_12023,N_11860,N_11823);
nand U12024 (N_12024,N_11868,N_11924);
or U12025 (N_12025,N_11944,N_11907);
xor U12026 (N_12026,N_11895,N_11997);
nor U12027 (N_12027,N_11827,N_11896);
xor U12028 (N_12028,N_11881,N_11968);
nor U12029 (N_12029,N_11988,N_11800);
or U12030 (N_12030,N_11824,N_11803);
nand U12031 (N_12031,N_11852,N_11898);
xor U12032 (N_12032,N_11871,N_11962);
nand U12033 (N_12033,N_11911,N_11932);
xor U12034 (N_12034,N_11951,N_11921);
xor U12035 (N_12035,N_11811,N_11922);
xor U12036 (N_12036,N_11990,N_11857);
or U12037 (N_12037,N_11994,N_11897);
xor U12038 (N_12038,N_11858,N_11923);
xor U12039 (N_12039,N_11905,N_11926);
nand U12040 (N_12040,N_11835,N_11870);
and U12041 (N_12041,N_11995,N_11848);
or U12042 (N_12042,N_11899,N_11903);
nor U12043 (N_12043,N_11825,N_11985);
and U12044 (N_12044,N_11839,N_11993);
nand U12045 (N_12045,N_11864,N_11925);
or U12046 (N_12046,N_11830,N_11882);
nor U12047 (N_12047,N_11836,N_11894);
or U12048 (N_12048,N_11928,N_11834);
and U12049 (N_12049,N_11915,N_11978);
nor U12050 (N_12050,N_11912,N_11970);
or U12051 (N_12051,N_11806,N_11815);
nor U12052 (N_12052,N_11885,N_11935);
nor U12053 (N_12053,N_11849,N_11810);
and U12054 (N_12054,N_11981,N_11801);
nor U12055 (N_12055,N_11889,N_11939);
or U12056 (N_12056,N_11818,N_11842);
xnor U12057 (N_12057,N_11909,N_11967);
and U12058 (N_12058,N_11855,N_11817);
nand U12059 (N_12059,N_11943,N_11937);
xnor U12060 (N_12060,N_11901,N_11828);
and U12061 (N_12061,N_11841,N_11850);
or U12062 (N_12062,N_11883,N_11996);
or U12063 (N_12063,N_11819,N_11844);
nand U12064 (N_12064,N_11966,N_11863);
nand U12065 (N_12065,N_11856,N_11976);
and U12066 (N_12066,N_11846,N_11877);
or U12067 (N_12067,N_11973,N_11991);
xnor U12068 (N_12068,N_11808,N_11961);
xor U12069 (N_12069,N_11965,N_11865);
nor U12070 (N_12070,N_11980,N_11904);
or U12071 (N_12071,N_11917,N_11987);
and U12072 (N_12072,N_11953,N_11826);
nor U12073 (N_12073,N_11948,N_11829);
or U12074 (N_12074,N_11879,N_11814);
and U12075 (N_12075,N_11914,N_11866);
or U12076 (N_12076,N_11929,N_11977);
nor U12077 (N_12077,N_11938,N_11831);
nand U12078 (N_12078,N_11983,N_11954);
and U12079 (N_12079,N_11906,N_11851);
nor U12080 (N_12080,N_11979,N_11816);
and U12081 (N_12081,N_11854,N_11908);
and U12082 (N_12082,N_11920,N_11890);
xnor U12083 (N_12083,N_11989,N_11927);
xnor U12084 (N_12084,N_11930,N_11878);
nand U12085 (N_12085,N_11840,N_11853);
nor U12086 (N_12086,N_11957,N_11999);
and U12087 (N_12087,N_11941,N_11891);
or U12088 (N_12088,N_11946,N_11933);
nor U12089 (N_12089,N_11972,N_11822);
xnor U12090 (N_12090,N_11971,N_11960);
nand U12091 (N_12091,N_11940,N_11867);
or U12092 (N_12092,N_11913,N_11931);
nand U12093 (N_12093,N_11942,N_11952);
nor U12094 (N_12094,N_11869,N_11876);
xor U12095 (N_12095,N_11813,N_11847);
and U12096 (N_12096,N_11812,N_11963);
nand U12097 (N_12097,N_11887,N_11947);
xor U12098 (N_12098,N_11934,N_11910);
nand U12099 (N_12099,N_11893,N_11955);
nand U12100 (N_12100,N_11829,N_11862);
nor U12101 (N_12101,N_11874,N_11863);
or U12102 (N_12102,N_11940,N_11988);
nand U12103 (N_12103,N_11855,N_11807);
or U12104 (N_12104,N_11958,N_11828);
or U12105 (N_12105,N_11863,N_11826);
and U12106 (N_12106,N_11893,N_11984);
nand U12107 (N_12107,N_11849,N_11949);
or U12108 (N_12108,N_11959,N_11932);
xnor U12109 (N_12109,N_11920,N_11823);
nor U12110 (N_12110,N_11997,N_11902);
nor U12111 (N_12111,N_11859,N_11896);
nand U12112 (N_12112,N_11802,N_11850);
nor U12113 (N_12113,N_11965,N_11905);
nand U12114 (N_12114,N_11903,N_11807);
or U12115 (N_12115,N_11834,N_11818);
xnor U12116 (N_12116,N_11874,N_11935);
and U12117 (N_12117,N_11900,N_11844);
nand U12118 (N_12118,N_11987,N_11976);
or U12119 (N_12119,N_11850,N_11921);
or U12120 (N_12120,N_11888,N_11927);
nor U12121 (N_12121,N_11827,N_11834);
nand U12122 (N_12122,N_11974,N_11972);
xor U12123 (N_12123,N_11962,N_11925);
and U12124 (N_12124,N_11824,N_11984);
and U12125 (N_12125,N_11948,N_11864);
or U12126 (N_12126,N_11887,N_11886);
xnor U12127 (N_12127,N_11873,N_11847);
nand U12128 (N_12128,N_11894,N_11872);
and U12129 (N_12129,N_11831,N_11839);
or U12130 (N_12130,N_11872,N_11916);
nor U12131 (N_12131,N_11811,N_11809);
and U12132 (N_12132,N_11926,N_11909);
nand U12133 (N_12133,N_11844,N_11805);
nand U12134 (N_12134,N_11804,N_11975);
xnor U12135 (N_12135,N_11881,N_11811);
xor U12136 (N_12136,N_11865,N_11902);
or U12137 (N_12137,N_11894,N_11843);
and U12138 (N_12138,N_11817,N_11852);
or U12139 (N_12139,N_11939,N_11903);
xor U12140 (N_12140,N_11858,N_11839);
nor U12141 (N_12141,N_11911,N_11969);
or U12142 (N_12142,N_11820,N_11872);
and U12143 (N_12143,N_11973,N_11893);
nand U12144 (N_12144,N_11906,N_11985);
nor U12145 (N_12145,N_11881,N_11852);
nand U12146 (N_12146,N_11908,N_11960);
xnor U12147 (N_12147,N_11981,N_11989);
xnor U12148 (N_12148,N_11816,N_11872);
and U12149 (N_12149,N_11911,N_11995);
xor U12150 (N_12150,N_11994,N_11881);
nor U12151 (N_12151,N_11980,N_11836);
nand U12152 (N_12152,N_11914,N_11863);
xnor U12153 (N_12153,N_11898,N_11958);
nor U12154 (N_12154,N_11807,N_11810);
nand U12155 (N_12155,N_11927,N_11911);
or U12156 (N_12156,N_11854,N_11829);
nand U12157 (N_12157,N_11967,N_11852);
xnor U12158 (N_12158,N_11836,N_11860);
nor U12159 (N_12159,N_11819,N_11880);
nor U12160 (N_12160,N_11887,N_11819);
xor U12161 (N_12161,N_11975,N_11873);
nand U12162 (N_12162,N_11852,N_11840);
nand U12163 (N_12163,N_11824,N_11817);
and U12164 (N_12164,N_11897,N_11949);
xor U12165 (N_12165,N_11830,N_11979);
xnor U12166 (N_12166,N_11955,N_11877);
and U12167 (N_12167,N_11857,N_11855);
xor U12168 (N_12168,N_11910,N_11899);
nor U12169 (N_12169,N_11923,N_11953);
nor U12170 (N_12170,N_11837,N_11927);
or U12171 (N_12171,N_11999,N_11804);
xnor U12172 (N_12172,N_11868,N_11899);
xnor U12173 (N_12173,N_11905,N_11988);
nor U12174 (N_12174,N_11838,N_11944);
xnor U12175 (N_12175,N_11930,N_11967);
or U12176 (N_12176,N_11959,N_11829);
xor U12177 (N_12177,N_11964,N_11938);
nor U12178 (N_12178,N_11841,N_11855);
nand U12179 (N_12179,N_11862,N_11940);
and U12180 (N_12180,N_11925,N_11960);
or U12181 (N_12181,N_11862,N_11966);
xor U12182 (N_12182,N_11909,N_11990);
and U12183 (N_12183,N_11986,N_11989);
nor U12184 (N_12184,N_11810,N_11898);
and U12185 (N_12185,N_11891,N_11842);
xnor U12186 (N_12186,N_11914,N_11838);
nor U12187 (N_12187,N_11937,N_11835);
nand U12188 (N_12188,N_11939,N_11845);
nor U12189 (N_12189,N_11800,N_11874);
nand U12190 (N_12190,N_11861,N_11915);
xnor U12191 (N_12191,N_11883,N_11866);
nand U12192 (N_12192,N_11850,N_11886);
and U12193 (N_12193,N_11873,N_11943);
nor U12194 (N_12194,N_11917,N_11804);
nand U12195 (N_12195,N_11976,N_11963);
nor U12196 (N_12196,N_11813,N_11953);
nor U12197 (N_12197,N_11859,N_11845);
xor U12198 (N_12198,N_11883,N_11983);
nor U12199 (N_12199,N_11964,N_11992);
nor U12200 (N_12200,N_12026,N_12137);
nand U12201 (N_12201,N_12078,N_12128);
nor U12202 (N_12202,N_12073,N_12036);
and U12203 (N_12203,N_12127,N_12142);
and U12204 (N_12204,N_12063,N_12027);
or U12205 (N_12205,N_12153,N_12151);
nor U12206 (N_12206,N_12170,N_12131);
nor U12207 (N_12207,N_12108,N_12017);
nor U12208 (N_12208,N_12177,N_12143);
nor U12209 (N_12209,N_12080,N_12109);
xnor U12210 (N_12210,N_12051,N_12185);
xor U12211 (N_12211,N_12165,N_12147);
and U12212 (N_12212,N_12001,N_12172);
and U12213 (N_12213,N_12098,N_12112);
or U12214 (N_12214,N_12083,N_12015);
or U12215 (N_12215,N_12032,N_12114);
nand U12216 (N_12216,N_12130,N_12039);
or U12217 (N_12217,N_12184,N_12159);
xnor U12218 (N_12218,N_12124,N_12093);
or U12219 (N_12219,N_12067,N_12181);
and U12220 (N_12220,N_12022,N_12104);
nand U12221 (N_12221,N_12038,N_12190);
or U12222 (N_12222,N_12117,N_12050);
xnor U12223 (N_12223,N_12187,N_12090);
and U12224 (N_12224,N_12033,N_12100);
nand U12225 (N_12225,N_12101,N_12122);
and U12226 (N_12226,N_12123,N_12049);
nor U12227 (N_12227,N_12168,N_12002);
nor U12228 (N_12228,N_12011,N_12003);
or U12229 (N_12229,N_12040,N_12047);
xnor U12230 (N_12230,N_12081,N_12118);
nor U12231 (N_12231,N_12059,N_12082);
and U12232 (N_12232,N_12126,N_12023);
or U12233 (N_12233,N_12057,N_12183);
or U12234 (N_12234,N_12044,N_12019);
and U12235 (N_12235,N_12097,N_12148);
nor U12236 (N_12236,N_12161,N_12070);
nand U12237 (N_12237,N_12155,N_12195);
nand U12238 (N_12238,N_12006,N_12046);
xor U12239 (N_12239,N_12007,N_12156);
nand U12240 (N_12240,N_12099,N_12062);
nor U12241 (N_12241,N_12145,N_12110);
xor U12242 (N_12242,N_12107,N_12029);
nand U12243 (N_12243,N_12095,N_12139);
and U12244 (N_12244,N_12077,N_12133);
and U12245 (N_12245,N_12000,N_12166);
xor U12246 (N_12246,N_12005,N_12125);
nor U12247 (N_12247,N_12103,N_12158);
and U12248 (N_12248,N_12088,N_12053);
nand U12249 (N_12249,N_12192,N_12171);
or U12250 (N_12250,N_12004,N_12068);
nand U12251 (N_12251,N_12174,N_12119);
nand U12252 (N_12252,N_12175,N_12064);
nand U12253 (N_12253,N_12169,N_12025);
nor U12254 (N_12254,N_12162,N_12037);
nand U12255 (N_12255,N_12196,N_12191);
nand U12256 (N_12256,N_12071,N_12105);
nand U12257 (N_12257,N_12009,N_12179);
xor U12258 (N_12258,N_12091,N_12018);
nand U12259 (N_12259,N_12136,N_12089);
nor U12260 (N_12260,N_12149,N_12035);
nand U12261 (N_12261,N_12146,N_12060);
nor U12262 (N_12262,N_12054,N_12092);
and U12263 (N_12263,N_12031,N_12048);
nand U12264 (N_12264,N_12042,N_12189);
nor U12265 (N_12265,N_12176,N_12024);
xnor U12266 (N_12266,N_12084,N_12198);
nand U12267 (N_12267,N_12069,N_12034);
and U12268 (N_12268,N_12020,N_12111);
nand U12269 (N_12269,N_12016,N_12074);
xor U12270 (N_12270,N_12058,N_12085);
and U12271 (N_12271,N_12193,N_12115);
nor U12272 (N_12272,N_12140,N_12132);
nor U12273 (N_12273,N_12056,N_12154);
nor U12274 (N_12274,N_12014,N_12144);
nor U12275 (N_12275,N_12141,N_12065);
and U12276 (N_12276,N_12045,N_12178);
nor U12277 (N_12277,N_12134,N_12157);
and U12278 (N_12278,N_12012,N_12066);
or U12279 (N_12279,N_12182,N_12180);
xor U12280 (N_12280,N_12055,N_12138);
xor U12281 (N_12281,N_12113,N_12129);
or U12282 (N_12282,N_12087,N_12102);
xor U12283 (N_12283,N_12173,N_12096);
nor U12284 (N_12284,N_12076,N_12010);
xnor U12285 (N_12285,N_12094,N_12152);
and U12286 (N_12286,N_12043,N_12106);
nor U12287 (N_12287,N_12021,N_12013);
nor U12288 (N_12288,N_12041,N_12061);
nand U12289 (N_12289,N_12163,N_12008);
or U12290 (N_12290,N_12121,N_12075);
nand U12291 (N_12291,N_12028,N_12120);
or U12292 (N_12292,N_12160,N_12086);
nand U12293 (N_12293,N_12194,N_12197);
nor U12294 (N_12294,N_12030,N_12188);
xnor U12295 (N_12295,N_12116,N_12135);
and U12296 (N_12296,N_12072,N_12150);
or U12297 (N_12297,N_12079,N_12052);
nand U12298 (N_12298,N_12199,N_12164);
xor U12299 (N_12299,N_12167,N_12186);
nor U12300 (N_12300,N_12089,N_12038);
and U12301 (N_12301,N_12108,N_12187);
and U12302 (N_12302,N_12191,N_12174);
nor U12303 (N_12303,N_12153,N_12146);
and U12304 (N_12304,N_12118,N_12088);
xor U12305 (N_12305,N_12032,N_12020);
nor U12306 (N_12306,N_12027,N_12150);
and U12307 (N_12307,N_12049,N_12154);
nand U12308 (N_12308,N_12073,N_12046);
and U12309 (N_12309,N_12091,N_12120);
xor U12310 (N_12310,N_12067,N_12017);
nor U12311 (N_12311,N_12131,N_12064);
nor U12312 (N_12312,N_12024,N_12109);
xor U12313 (N_12313,N_12153,N_12195);
nand U12314 (N_12314,N_12194,N_12041);
xnor U12315 (N_12315,N_12122,N_12049);
nand U12316 (N_12316,N_12122,N_12045);
nand U12317 (N_12317,N_12101,N_12111);
and U12318 (N_12318,N_12023,N_12162);
nand U12319 (N_12319,N_12005,N_12128);
and U12320 (N_12320,N_12198,N_12082);
xor U12321 (N_12321,N_12091,N_12054);
nand U12322 (N_12322,N_12174,N_12072);
and U12323 (N_12323,N_12117,N_12051);
and U12324 (N_12324,N_12092,N_12037);
nor U12325 (N_12325,N_12041,N_12187);
nand U12326 (N_12326,N_12010,N_12185);
nor U12327 (N_12327,N_12162,N_12051);
nor U12328 (N_12328,N_12198,N_12174);
and U12329 (N_12329,N_12038,N_12123);
or U12330 (N_12330,N_12073,N_12015);
nand U12331 (N_12331,N_12013,N_12158);
or U12332 (N_12332,N_12047,N_12136);
or U12333 (N_12333,N_12198,N_12043);
nand U12334 (N_12334,N_12037,N_12191);
xor U12335 (N_12335,N_12106,N_12038);
xnor U12336 (N_12336,N_12089,N_12146);
and U12337 (N_12337,N_12192,N_12021);
xor U12338 (N_12338,N_12032,N_12130);
and U12339 (N_12339,N_12062,N_12189);
nand U12340 (N_12340,N_12086,N_12097);
and U12341 (N_12341,N_12182,N_12015);
nor U12342 (N_12342,N_12059,N_12085);
nand U12343 (N_12343,N_12052,N_12108);
and U12344 (N_12344,N_12156,N_12028);
nand U12345 (N_12345,N_12121,N_12020);
and U12346 (N_12346,N_12195,N_12092);
xor U12347 (N_12347,N_12084,N_12155);
and U12348 (N_12348,N_12179,N_12151);
xnor U12349 (N_12349,N_12014,N_12104);
nand U12350 (N_12350,N_12077,N_12004);
nand U12351 (N_12351,N_12088,N_12179);
or U12352 (N_12352,N_12095,N_12014);
or U12353 (N_12353,N_12145,N_12029);
and U12354 (N_12354,N_12053,N_12135);
and U12355 (N_12355,N_12119,N_12008);
xor U12356 (N_12356,N_12091,N_12162);
or U12357 (N_12357,N_12094,N_12052);
or U12358 (N_12358,N_12147,N_12023);
or U12359 (N_12359,N_12105,N_12138);
or U12360 (N_12360,N_12074,N_12101);
nand U12361 (N_12361,N_12190,N_12092);
nand U12362 (N_12362,N_12016,N_12170);
xnor U12363 (N_12363,N_12050,N_12180);
or U12364 (N_12364,N_12059,N_12176);
or U12365 (N_12365,N_12132,N_12010);
xor U12366 (N_12366,N_12047,N_12182);
nand U12367 (N_12367,N_12108,N_12184);
nand U12368 (N_12368,N_12070,N_12140);
and U12369 (N_12369,N_12136,N_12198);
nand U12370 (N_12370,N_12064,N_12044);
nand U12371 (N_12371,N_12102,N_12062);
or U12372 (N_12372,N_12120,N_12033);
xnor U12373 (N_12373,N_12024,N_12110);
nor U12374 (N_12374,N_12122,N_12168);
nand U12375 (N_12375,N_12086,N_12081);
or U12376 (N_12376,N_12050,N_12002);
and U12377 (N_12377,N_12108,N_12178);
or U12378 (N_12378,N_12172,N_12198);
nand U12379 (N_12379,N_12087,N_12082);
nand U12380 (N_12380,N_12069,N_12116);
xnor U12381 (N_12381,N_12122,N_12104);
nand U12382 (N_12382,N_12172,N_12133);
nand U12383 (N_12383,N_12017,N_12176);
xor U12384 (N_12384,N_12069,N_12088);
or U12385 (N_12385,N_12179,N_12148);
nor U12386 (N_12386,N_12110,N_12041);
or U12387 (N_12387,N_12195,N_12192);
or U12388 (N_12388,N_12002,N_12031);
or U12389 (N_12389,N_12099,N_12079);
or U12390 (N_12390,N_12194,N_12001);
xor U12391 (N_12391,N_12138,N_12107);
and U12392 (N_12392,N_12033,N_12163);
nor U12393 (N_12393,N_12029,N_12191);
and U12394 (N_12394,N_12146,N_12167);
or U12395 (N_12395,N_12028,N_12049);
and U12396 (N_12396,N_12146,N_12164);
or U12397 (N_12397,N_12169,N_12051);
nor U12398 (N_12398,N_12152,N_12176);
xor U12399 (N_12399,N_12067,N_12087);
and U12400 (N_12400,N_12326,N_12254);
and U12401 (N_12401,N_12223,N_12300);
xnor U12402 (N_12402,N_12271,N_12243);
nand U12403 (N_12403,N_12328,N_12259);
xor U12404 (N_12404,N_12386,N_12322);
xnor U12405 (N_12405,N_12237,N_12276);
nor U12406 (N_12406,N_12380,N_12216);
or U12407 (N_12407,N_12288,N_12369);
nor U12408 (N_12408,N_12229,N_12284);
nor U12409 (N_12409,N_12338,N_12309);
or U12410 (N_12410,N_12367,N_12398);
xor U12411 (N_12411,N_12324,N_12252);
or U12412 (N_12412,N_12342,N_12205);
nand U12413 (N_12413,N_12262,N_12201);
nor U12414 (N_12414,N_12203,N_12347);
nand U12415 (N_12415,N_12366,N_12343);
xor U12416 (N_12416,N_12379,N_12282);
nand U12417 (N_12417,N_12332,N_12245);
and U12418 (N_12418,N_12202,N_12236);
nand U12419 (N_12419,N_12219,N_12283);
nor U12420 (N_12420,N_12306,N_12396);
and U12421 (N_12421,N_12323,N_12339);
or U12422 (N_12422,N_12215,N_12220);
nor U12423 (N_12423,N_12267,N_12305);
nor U12424 (N_12424,N_12240,N_12384);
nand U12425 (N_12425,N_12311,N_12315);
nand U12426 (N_12426,N_12387,N_12295);
nor U12427 (N_12427,N_12354,N_12381);
xnor U12428 (N_12428,N_12256,N_12310);
xnor U12429 (N_12429,N_12281,N_12210);
or U12430 (N_12430,N_12330,N_12360);
and U12431 (N_12431,N_12255,N_12388);
nor U12432 (N_12432,N_12248,N_12222);
and U12433 (N_12433,N_12209,N_12390);
or U12434 (N_12434,N_12226,N_12241);
and U12435 (N_12435,N_12320,N_12359);
nor U12436 (N_12436,N_12289,N_12280);
and U12437 (N_12437,N_12302,N_12346);
nand U12438 (N_12438,N_12331,N_12224);
nor U12439 (N_12439,N_12263,N_12301);
xor U12440 (N_12440,N_12232,N_12365);
nor U12441 (N_12441,N_12313,N_12362);
and U12442 (N_12442,N_12351,N_12333);
or U12443 (N_12443,N_12206,N_12389);
xor U12444 (N_12444,N_12239,N_12304);
or U12445 (N_12445,N_12308,N_12272);
nand U12446 (N_12446,N_12238,N_12350);
and U12447 (N_12447,N_12235,N_12277);
nor U12448 (N_12448,N_12361,N_12257);
and U12449 (N_12449,N_12368,N_12213);
nand U12450 (N_12450,N_12296,N_12358);
nand U12451 (N_12451,N_12261,N_12374);
or U12452 (N_12452,N_12352,N_12292);
or U12453 (N_12453,N_12251,N_12244);
xnor U12454 (N_12454,N_12378,N_12207);
or U12455 (N_12455,N_12253,N_12266);
or U12456 (N_12456,N_12246,N_12234);
and U12457 (N_12457,N_12392,N_12287);
nand U12458 (N_12458,N_12377,N_12357);
nand U12459 (N_12459,N_12335,N_12337);
xor U12460 (N_12460,N_12260,N_12395);
and U12461 (N_12461,N_12264,N_12307);
nand U12462 (N_12462,N_12364,N_12376);
and U12463 (N_12463,N_12285,N_12269);
nor U12464 (N_12464,N_12247,N_12228);
nor U12465 (N_12465,N_12312,N_12373);
nand U12466 (N_12466,N_12230,N_12317);
nor U12467 (N_12467,N_12316,N_12344);
and U12468 (N_12468,N_12231,N_12278);
or U12469 (N_12469,N_12341,N_12270);
nand U12470 (N_12470,N_12204,N_12297);
and U12471 (N_12471,N_12348,N_12200);
xnor U12472 (N_12472,N_12208,N_12273);
nand U12473 (N_12473,N_12274,N_12391);
nand U12474 (N_12474,N_12372,N_12314);
or U12475 (N_12475,N_12345,N_12293);
nand U12476 (N_12476,N_12250,N_12363);
xnor U12477 (N_12477,N_12242,N_12298);
or U12478 (N_12478,N_12290,N_12371);
and U12479 (N_12479,N_12353,N_12214);
nor U12480 (N_12480,N_12399,N_12385);
and U12481 (N_12481,N_12393,N_12318);
or U12482 (N_12482,N_12383,N_12258);
xor U12483 (N_12483,N_12268,N_12233);
or U12484 (N_12484,N_12394,N_12397);
or U12485 (N_12485,N_12356,N_12299);
nand U12486 (N_12486,N_12275,N_12286);
or U12487 (N_12487,N_12218,N_12355);
and U12488 (N_12488,N_12329,N_12334);
and U12489 (N_12489,N_12294,N_12321);
xor U12490 (N_12490,N_12336,N_12382);
and U12491 (N_12491,N_12325,N_12327);
nor U12492 (N_12492,N_12291,N_12370);
nor U12493 (N_12493,N_12303,N_12375);
xnor U12494 (N_12494,N_12227,N_12217);
nand U12495 (N_12495,N_12225,N_12319);
nor U12496 (N_12496,N_12265,N_12279);
nor U12497 (N_12497,N_12249,N_12212);
nor U12498 (N_12498,N_12221,N_12349);
xor U12499 (N_12499,N_12211,N_12340);
nand U12500 (N_12500,N_12376,N_12337);
nand U12501 (N_12501,N_12352,N_12377);
nor U12502 (N_12502,N_12298,N_12362);
nand U12503 (N_12503,N_12242,N_12394);
nor U12504 (N_12504,N_12217,N_12300);
nand U12505 (N_12505,N_12275,N_12294);
xor U12506 (N_12506,N_12265,N_12235);
or U12507 (N_12507,N_12386,N_12235);
nor U12508 (N_12508,N_12228,N_12304);
or U12509 (N_12509,N_12219,N_12273);
nand U12510 (N_12510,N_12352,N_12240);
and U12511 (N_12511,N_12345,N_12257);
xnor U12512 (N_12512,N_12284,N_12312);
and U12513 (N_12513,N_12272,N_12203);
xnor U12514 (N_12514,N_12396,N_12262);
and U12515 (N_12515,N_12204,N_12386);
nor U12516 (N_12516,N_12356,N_12215);
or U12517 (N_12517,N_12298,N_12392);
and U12518 (N_12518,N_12229,N_12240);
or U12519 (N_12519,N_12352,N_12329);
xor U12520 (N_12520,N_12362,N_12270);
or U12521 (N_12521,N_12336,N_12283);
xor U12522 (N_12522,N_12249,N_12279);
xnor U12523 (N_12523,N_12346,N_12395);
nand U12524 (N_12524,N_12334,N_12332);
nand U12525 (N_12525,N_12328,N_12345);
nor U12526 (N_12526,N_12212,N_12288);
and U12527 (N_12527,N_12351,N_12360);
nand U12528 (N_12528,N_12345,N_12310);
nand U12529 (N_12529,N_12324,N_12205);
and U12530 (N_12530,N_12298,N_12307);
nand U12531 (N_12531,N_12390,N_12353);
and U12532 (N_12532,N_12397,N_12271);
nor U12533 (N_12533,N_12341,N_12213);
or U12534 (N_12534,N_12226,N_12283);
and U12535 (N_12535,N_12240,N_12394);
nor U12536 (N_12536,N_12248,N_12296);
nand U12537 (N_12537,N_12225,N_12326);
or U12538 (N_12538,N_12229,N_12364);
or U12539 (N_12539,N_12362,N_12280);
nor U12540 (N_12540,N_12266,N_12343);
xor U12541 (N_12541,N_12328,N_12281);
and U12542 (N_12542,N_12235,N_12292);
nand U12543 (N_12543,N_12396,N_12370);
nor U12544 (N_12544,N_12281,N_12211);
nor U12545 (N_12545,N_12318,N_12343);
nor U12546 (N_12546,N_12361,N_12374);
and U12547 (N_12547,N_12259,N_12288);
nand U12548 (N_12548,N_12290,N_12277);
nand U12549 (N_12549,N_12388,N_12321);
nor U12550 (N_12550,N_12223,N_12211);
nor U12551 (N_12551,N_12254,N_12288);
xor U12552 (N_12552,N_12398,N_12345);
nand U12553 (N_12553,N_12333,N_12257);
xor U12554 (N_12554,N_12387,N_12364);
or U12555 (N_12555,N_12327,N_12239);
and U12556 (N_12556,N_12324,N_12267);
nor U12557 (N_12557,N_12386,N_12283);
xor U12558 (N_12558,N_12227,N_12232);
nor U12559 (N_12559,N_12243,N_12265);
nand U12560 (N_12560,N_12281,N_12218);
and U12561 (N_12561,N_12262,N_12351);
nand U12562 (N_12562,N_12359,N_12299);
nand U12563 (N_12563,N_12224,N_12300);
nand U12564 (N_12564,N_12241,N_12396);
xnor U12565 (N_12565,N_12282,N_12253);
or U12566 (N_12566,N_12259,N_12380);
xor U12567 (N_12567,N_12269,N_12373);
or U12568 (N_12568,N_12231,N_12232);
or U12569 (N_12569,N_12218,N_12245);
and U12570 (N_12570,N_12210,N_12234);
nand U12571 (N_12571,N_12242,N_12365);
xnor U12572 (N_12572,N_12353,N_12323);
nand U12573 (N_12573,N_12315,N_12372);
xnor U12574 (N_12574,N_12365,N_12293);
or U12575 (N_12575,N_12285,N_12339);
or U12576 (N_12576,N_12320,N_12314);
nand U12577 (N_12577,N_12240,N_12246);
and U12578 (N_12578,N_12265,N_12343);
nand U12579 (N_12579,N_12261,N_12362);
and U12580 (N_12580,N_12327,N_12397);
and U12581 (N_12581,N_12261,N_12226);
and U12582 (N_12582,N_12211,N_12336);
xnor U12583 (N_12583,N_12227,N_12299);
or U12584 (N_12584,N_12378,N_12355);
and U12585 (N_12585,N_12247,N_12271);
or U12586 (N_12586,N_12379,N_12338);
xnor U12587 (N_12587,N_12286,N_12269);
xor U12588 (N_12588,N_12242,N_12366);
nor U12589 (N_12589,N_12203,N_12354);
or U12590 (N_12590,N_12221,N_12243);
nor U12591 (N_12591,N_12273,N_12380);
nand U12592 (N_12592,N_12370,N_12262);
nor U12593 (N_12593,N_12337,N_12378);
xor U12594 (N_12594,N_12257,N_12312);
or U12595 (N_12595,N_12345,N_12277);
or U12596 (N_12596,N_12298,N_12308);
nor U12597 (N_12597,N_12342,N_12333);
nor U12598 (N_12598,N_12278,N_12369);
nand U12599 (N_12599,N_12293,N_12204);
and U12600 (N_12600,N_12585,N_12481);
xor U12601 (N_12601,N_12454,N_12434);
or U12602 (N_12602,N_12464,N_12428);
and U12603 (N_12603,N_12441,N_12506);
or U12604 (N_12604,N_12475,N_12442);
xnor U12605 (N_12605,N_12427,N_12509);
xor U12606 (N_12606,N_12548,N_12457);
nand U12607 (N_12607,N_12564,N_12486);
and U12608 (N_12608,N_12407,N_12408);
xnor U12609 (N_12609,N_12535,N_12440);
nand U12610 (N_12610,N_12581,N_12589);
xnor U12611 (N_12611,N_12461,N_12538);
xnor U12612 (N_12612,N_12404,N_12420);
nand U12613 (N_12613,N_12588,N_12551);
and U12614 (N_12614,N_12561,N_12455);
nor U12615 (N_12615,N_12433,N_12406);
nand U12616 (N_12616,N_12488,N_12549);
or U12617 (N_12617,N_12542,N_12492);
xnor U12618 (N_12618,N_12444,N_12487);
and U12619 (N_12619,N_12591,N_12559);
nor U12620 (N_12620,N_12527,N_12537);
nand U12621 (N_12621,N_12520,N_12523);
xor U12622 (N_12622,N_12554,N_12416);
or U12623 (N_12623,N_12522,N_12592);
and U12624 (N_12624,N_12584,N_12436);
and U12625 (N_12625,N_12458,N_12423);
xor U12626 (N_12626,N_12419,N_12400);
nand U12627 (N_12627,N_12518,N_12411);
nand U12628 (N_12628,N_12576,N_12401);
or U12629 (N_12629,N_12553,N_12550);
xnor U12630 (N_12630,N_12540,N_12573);
nand U12631 (N_12631,N_12410,N_12402);
nor U12632 (N_12632,N_12534,N_12519);
nor U12633 (N_12633,N_12571,N_12499);
nor U12634 (N_12634,N_12463,N_12504);
xnor U12635 (N_12635,N_12438,N_12414);
nor U12636 (N_12636,N_12474,N_12482);
or U12637 (N_12637,N_12493,N_12451);
and U12638 (N_12638,N_12417,N_12526);
xnor U12639 (N_12639,N_12439,N_12525);
nand U12640 (N_12640,N_12539,N_12483);
xor U12641 (N_12641,N_12524,N_12477);
and U12642 (N_12642,N_12543,N_12432);
nor U12643 (N_12643,N_12412,N_12479);
xnor U12644 (N_12644,N_12594,N_12536);
nor U12645 (N_12645,N_12500,N_12453);
and U12646 (N_12646,N_12430,N_12473);
or U12647 (N_12647,N_12590,N_12447);
nand U12648 (N_12648,N_12579,N_12470);
xnor U12649 (N_12649,N_12403,N_12495);
nor U12650 (N_12650,N_12545,N_12530);
nand U12651 (N_12651,N_12468,N_12514);
nand U12652 (N_12652,N_12478,N_12508);
or U12653 (N_12653,N_12547,N_12510);
and U12654 (N_12654,N_12556,N_12574);
or U12655 (N_12655,N_12489,N_12435);
xnor U12656 (N_12656,N_12512,N_12565);
nand U12657 (N_12657,N_12491,N_12422);
or U12658 (N_12658,N_12586,N_12572);
and U12659 (N_12659,N_12459,N_12560);
or U12660 (N_12660,N_12544,N_12443);
and U12661 (N_12661,N_12462,N_12421);
xnor U12662 (N_12662,N_12484,N_12452);
nand U12663 (N_12663,N_12431,N_12490);
and U12664 (N_12664,N_12532,N_12424);
nor U12665 (N_12665,N_12567,N_12563);
nand U12666 (N_12666,N_12541,N_12409);
nand U12667 (N_12667,N_12562,N_12558);
nand U12668 (N_12668,N_12566,N_12596);
nor U12669 (N_12669,N_12480,N_12568);
nor U12670 (N_12670,N_12476,N_12502);
nor U12671 (N_12671,N_12466,N_12528);
xnor U12672 (N_12672,N_12557,N_12533);
or U12673 (N_12673,N_12448,N_12583);
nand U12674 (N_12674,N_12555,N_12469);
xor U12675 (N_12675,N_12472,N_12552);
nor U12676 (N_12676,N_12513,N_12467);
xnor U12677 (N_12677,N_12456,N_12505);
nand U12678 (N_12678,N_12445,N_12587);
or U12679 (N_12679,N_12599,N_12415);
or U12680 (N_12680,N_12593,N_12531);
nor U12681 (N_12681,N_12570,N_12437);
nand U12682 (N_12682,N_12516,N_12511);
nor U12683 (N_12683,N_12575,N_12405);
or U12684 (N_12684,N_12496,N_12501);
nand U12685 (N_12685,N_12418,N_12521);
xor U12686 (N_12686,N_12598,N_12460);
and U12687 (N_12687,N_12582,N_12515);
nand U12688 (N_12688,N_12450,N_12503);
nand U12689 (N_12689,N_12471,N_12429);
nor U12690 (N_12690,N_12497,N_12507);
xor U12691 (N_12691,N_12580,N_12569);
nor U12692 (N_12692,N_12597,N_12529);
or U12693 (N_12693,N_12546,N_12577);
or U12694 (N_12694,N_12485,N_12498);
nand U12695 (N_12695,N_12446,N_12425);
xor U12696 (N_12696,N_12413,N_12578);
or U12697 (N_12697,N_12595,N_12517);
or U12698 (N_12698,N_12449,N_12426);
xnor U12699 (N_12699,N_12465,N_12494);
and U12700 (N_12700,N_12496,N_12517);
or U12701 (N_12701,N_12593,N_12568);
and U12702 (N_12702,N_12445,N_12447);
nor U12703 (N_12703,N_12500,N_12405);
nand U12704 (N_12704,N_12410,N_12473);
nand U12705 (N_12705,N_12452,N_12477);
nor U12706 (N_12706,N_12522,N_12544);
or U12707 (N_12707,N_12554,N_12411);
or U12708 (N_12708,N_12498,N_12459);
or U12709 (N_12709,N_12415,N_12524);
xor U12710 (N_12710,N_12504,N_12575);
nor U12711 (N_12711,N_12408,N_12428);
and U12712 (N_12712,N_12407,N_12593);
and U12713 (N_12713,N_12463,N_12514);
nand U12714 (N_12714,N_12494,N_12594);
and U12715 (N_12715,N_12441,N_12545);
nor U12716 (N_12716,N_12502,N_12410);
nand U12717 (N_12717,N_12534,N_12423);
nor U12718 (N_12718,N_12517,N_12509);
nand U12719 (N_12719,N_12502,N_12596);
nand U12720 (N_12720,N_12477,N_12484);
or U12721 (N_12721,N_12574,N_12510);
and U12722 (N_12722,N_12437,N_12587);
and U12723 (N_12723,N_12514,N_12543);
and U12724 (N_12724,N_12513,N_12437);
nor U12725 (N_12725,N_12529,N_12583);
and U12726 (N_12726,N_12563,N_12528);
nand U12727 (N_12727,N_12496,N_12586);
or U12728 (N_12728,N_12503,N_12523);
nand U12729 (N_12729,N_12406,N_12446);
nand U12730 (N_12730,N_12542,N_12419);
or U12731 (N_12731,N_12524,N_12551);
or U12732 (N_12732,N_12421,N_12488);
xor U12733 (N_12733,N_12542,N_12485);
or U12734 (N_12734,N_12430,N_12404);
or U12735 (N_12735,N_12425,N_12483);
nor U12736 (N_12736,N_12557,N_12407);
nand U12737 (N_12737,N_12598,N_12579);
nand U12738 (N_12738,N_12468,N_12484);
nand U12739 (N_12739,N_12408,N_12431);
and U12740 (N_12740,N_12434,N_12557);
and U12741 (N_12741,N_12480,N_12514);
nand U12742 (N_12742,N_12425,N_12502);
or U12743 (N_12743,N_12465,N_12450);
nand U12744 (N_12744,N_12412,N_12530);
and U12745 (N_12745,N_12501,N_12564);
or U12746 (N_12746,N_12525,N_12457);
and U12747 (N_12747,N_12567,N_12595);
and U12748 (N_12748,N_12453,N_12426);
nand U12749 (N_12749,N_12415,N_12440);
or U12750 (N_12750,N_12484,N_12479);
and U12751 (N_12751,N_12408,N_12443);
and U12752 (N_12752,N_12584,N_12535);
xnor U12753 (N_12753,N_12528,N_12425);
and U12754 (N_12754,N_12499,N_12545);
xnor U12755 (N_12755,N_12494,N_12583);
or U12756 (N_12756,N_12538,N_12531);
xor U12757 (N_12757,N_12549,N_12546);
xnor U12758 (N_12758,N_12566,N_12573);
and U12759 (N_12759,N_12457,N_12406);
nor U12760 (N_12760,N_12544,N_12584);
xnor U12761 (N_12761,N_12515,N_12432);
and U12762 (N_12762,N_12476,N_12587);
nand U12763 (N_12763,N_12574,N_12495);
xor U12764 (N_12764,N_12442,N_12422);
nor U12765 (N_12765,N_12422,N_12495);
nor U12766 (N_12766,N_12403,N_12439);
nand U12767 (N_12767,N_12454,N_12523);
xor U12768 (N_12768,N_12477,N_12474);
xor U12769 (N_12769,N_12570,N_12516);
nor U12770 (N_12770,N_12454,N_12561);
nor U12771 (N_12771,N_12450,N_12460);
nand U12772 (N_12772,N_12480,N_12401);
nand U12773 (N_12773,N_12577,N_12492);
nand U12774 (N_12774,N_12532,N_12459);
xor U12775 (N_12775,N_12455,N_12454);
nor U12776 (N_12776,N_12420,N_12406);
or U12777 (N_12777,N_12574,N_12461);
nand U12778 (N_12778,N_12551,N_12547);
and U12779 (N_12779,N_12545,N_12520);
xor U12780 (N_12780,N_12489,N_12553);
and U12781 (N_12781,N_12493,N_12563);
xor U12782 (N_12782,N_12492,N_12429);
xnor U12783 (N_12783,N_12559,N_12509);
xor U12784 (N_12784,N_12539,N_12587);
or U12785 (N_12785,N_12575,N_12417);
and U12786 (N_12786,N_12550,N_12502);
or U12787 (N_12787,N_12547,N_12447);
nor U12788 (N_12788,N_12410,N_12418);
nor U12789 (N_12789,N_12483,N_12480);
and U12790 (N_12790,N_12594,N_12435);
nand U12791 (N_12791,N_12522,N_12511);
and U12792 (N_12792,N_12554,N_12570);
nor U12793 (N_12793,N_12427,N_12521);
nand U12794 (N_12794,N_12466,N_12555);
and U12795 (N_12795,N_12585,N_12420);
nand U12796 (N_12796,N_12530,N_12402);
nand U12797 (N_12797,N_12414,N_12402);
and U12798 (N_12798,N_12505,N_12525);
nand U12799 (N_12799,N_12526,N_12487);
nand U12800 (N_12800,N_12662,N_12792);
or U12801 (N_12801,N_12796,N_12646);
nand U12802 (N_12802,N_12695,N_12610);
xor U12803 (N_12803,N_12617,N_12783);
and U12804 (N_12804,N_12734,N_12715);
nand U12805 (N_12805,N_12670,N_12723);
nor U12806 (N_12806,N_12779,N_12624);
nand U12807 (N_12807,N_12639,N_12743);
and U12808 (N_12808,N_12665,N_12600);
xnor U12809 (N_12809,N_12747,N_12766);
nand U12810 (N_12810,N_12674,N_12650);
or U12811 (N_12811,N_12793,N_12777);
or U12812 (N_12812,N_12709,N_12609);
or U12813 (N_12813,N_12745,N_12686);
xnor U12814 (N_12814,N_12703,N_12730);
and U12815 (N_12815,N_12611,N_12725);
or U12816 (N_12816,N_12672,N_12698);
xor U12817 (N_12817,N_12755,N_12739);
or U12818 (N_12818,N_12719,N_12735);
and U12819 (N_12819,N_12673,N_12706);
nor U12820 (N_12820,N_12760,N_12780);
nand U12821 (N_12821,N_12696,N_12605);
nor U12822 (N_12822,N_12632,N_12630);
xor U12823 (N_12823,N_12750,N_12797);
xor U12824 (N_12824,N_12620,N_12737);
or U12825 (N_12825,N_12789,N_12623);
or U12826 (N_12826,N_12705,N_12769);
and U12827 (N_12827,N_12713,N_12722);
nor U12828 (N_12828,N_12647,N_12661);
nand U12829 (N_12829,N_12613,N_12700);
nand U12830 (N_12830,N_12603,N_12699);
and U12831 (N_12831,N_12729,N_12710);
nor U12832 (N_12832,N_12704,N_12656);
nor U12833 (N_12833,N_12770,N_12631);
xnor U12834 (N_12834,N_12638,N_12741);
nor U12835 (N_12835,N_12680,N_12691);
nor U12836 (N_12836,N_12681,N_12726);
xnor U12837 (N_12837,N_12635,N_12763);
xnor U12838 (N_12838,N_12782,N_12761);
nor U12839 (N_12839,N_12659,N_12795);
or U12840 (N_12840,N_12702,N_12757);
nand U12841 (N_12841,N_12648,N_12798);
nand U12842 (N_12842,N_12727,N_12784);
nor U12843 (N_12843,N_12668,N_12759);
xnor U12844 (N_12844,N_12718,N_12604);
or U12845 (N_12845,N_12640,N_12787);
and U12846 (N_12846,N_12666,N_12627);
or U12847 (N_12847,N_12669,N_12733);
or U12848 (N_12848,N_12606,N_12751);
nand U12849 (N_12849,N_12621,N_12682);
nor U12850 (N_12850,N_12664,N_12643);
nor U12851 (N_12851,N_12628,N_12602);
or U12852 (N_12852,N_12771,N_12618);
nand U12853 (N_12853,N_12667,N_12636);
nand U12854 (N_12854,N_12714,N_12772);
or U12855 (N_12855,N_12615,N_12688);
and U12856 (N_12856,N_12622,N_12775);
and U12857 (N_12857,N_12685,N_12671);
nor U12858 (N_12858,N_12658,N_12708);
nand U12859 (N_12859,N_12758,N_12684);
and U12860 (N_12860,N_12768,N_12655);
or U12861 (N_12861,N_12689,N_12612);
nand U12862 (N_12862,N_12676,N_12675);
nor U12863 (N_12863,N_12711,N_12712);
nand U12864 (N_12864,N_12794,N_12791);
or U12865 (N_12865,N_12790,N_12778);
and U12866 (N_12866,N_12764,N_12641);
and U12867 (N_12867,N_12644,N_12781);
and U12868 (N_12868,N_12767,N_12788);
and U12869 (N_12869,N_12679,N_12785);
nand U12870 (N_12870,N_12690,N_12637);
nand U12871 (N_12871,N_12642,N_12732);
or U12872 (N_12872,N_12692,N_12724);
and U12873 (N_12873,N_12746,N_12749);
or U12874 (N_12874,N_12651,N_12765);
and U12875 (N_12875,N_12683,N_12614);
nand U12876 (N_12876,N_12716,N_12616);
xor U12877 (N_12877,N_12720,N_12657);
and U12878 (N_12878,N_12697,N_12707);
nand U12879 (N_12879,N_12754,N_12728);
xnor U12880 (N_12880,N_12626,N_12786);
nand U12881 (N_12881,N_12742,N_12694);
nand U12882 (N_12882,N_12677,N_12663);
nand U12883 (N_12883,N_12660,N_12753);
or U12884 (N_12884,N_12601,N_12721);
and U12885 (N_12885,N_12717,N_12645);
or U12886 (N_12886,N_12748,N_12774);
nor U12887 (N_12887,N_12625,N_12652);
or U12888 (N_12888,N_12653,N_12633);
xor U12889 (N_12889,N_12740,N_12744);
nand U12890 (N_12890,N_12649,N_12608);
nand U12891 (N_12891,N_12693,N_12619);
xor U12892 (N_12892,N_12752,N_12634);
or U12893 (N_12893,N_12776,N_12654);
and U12894 (N_12894,N_12731,N_12773);
nand U12895 (N_12895,N_12736,N_12799);
and U12896 (N_12896,N_12738,N_12678);
nor U12897 (N_12897,N_12762,N_12701);
nand U12898 (N_12898,N_12607,N_12629);
or U12899 (N_12899,N_12687,N_12756);
or U12900 (N_12900,N_12677,N_12657);
nand U12901 (N_12901,N_12683,N_12698);
xor U12902 (N_12902,N_12658,N_12682);
xnor U12903 (N_12903,N_12603,N_12623);
nor U12904 (N_12904,N_12743,N_12627);
xnor U12905 (N_12905,N_12704,N_12643);
or U12906 (N_12906,N_12673,N_12661);
nand U12907 (N_12907,N_12624,N_12691);
nand U12908 (N_12908,N_12631,N_12798);
nor U12909 (N_12909,N_12785,N_12692);
or U12910 (N_12910,N_12682,N_12753);
nor U12911 (N_12911,N_12774,N_12642);
nand U12912 (N_12912,N_12744,N_12730);
nand U12913 (N_12913,N_12648,N_12765);
xor U12914 (N_12914,N_12647,N_12794);
and U12915 (N_12915,N_12630,N_12612);
or U12916 (N_12916,N_12731,N_12600);
and U12917 (N_12917,N_12770,N_12642);
or U12918 (N_12918,N_12608,N_12742);
or U12919 (N_12919,N_12742,N_12662);
nor U12920 (N_12920,N_12774,N_12690);
and U12921 (N_12921,N_12654,N_12648);
and U12922 (N_12922,N_12751,N_12784);
xnor U12923 (N_12923,N_12651,N_12744);
nand U12924 (N_12924,N_12696,N_12721);
and U12925 (N_12925,N_12673,N_12760);
or U12926 (N_12926,N_12630,N_12795);
or U12927 (N_12927,N_12725,N_12785);
xnor U12928 (N_12928,N_12715,N_12603);
or U12929 (N_12929,N_12770,N_12720);
nor U12930 (N_12930,N_12711,N_12790);
and U12931 (N_12931,N_12787,N_12798);
xor U12932 (N_12932,N_12713,N_12689);
nor U12933 (N_12933,N_12707,N_12737);
nor U12934 (N_12934,N_12630,N_12799);
nor U12935 (N_12935,N_12736,N_12619);
and U12936 (N_12936,N_12631,N_12761);
and U12937 (N_12937,N_12649,N_12772);
nand U12938 (N_12938,N_12784,N_12732);
or U12939 (N_12939,N_12766,N_12664);
nor U12940 (N_12940,N_12765,N_12656);
nand U12941 (N_12941,N_12767,N_12608);
and U12942 (N_12942,N_12792,N_12673);
xor U12943 (N_12943,N_12789,N_12760);
and U12944 (N_12944,N_12750,N_12708);
nor U12945 (N_12945,N_12722,N_12682);
nor U12946 (N_12946,N_12782,N_12797);
nor U12947 (N_12947,N_12665,N_12693);
xor U12948 (N_12948,N_12618,N_12673);
nand U12949 (N_12949,N_12703,N_12755);
and U12950 (N_12950,N_12738,N_12743);
xnor U12951 (N_12951,N_12764,N_12633);
and U12952 (N_12952,N_12752,N_12791);
xor U12953 (N_12953,N_12633,N_12663);
or U12954 (N_12954,N_12759,N_12789);
nor U12955 (N_12955,N_12765,N_12618);
nand U12956 (N_12956,N_12605,N_12702);
or U12957 (N_12957,N_12704,N_12743);
or U12958 (N_12958,N_12777,N_12636);
nand U12959 (N_12959,N_12712,N_12647);
nand U12960 (N_12960,N_12771,N_12707);
nand U12961 (N_12961,N_12631,N_12628);
xnor U12962 (N_12962,N_12768,N_12784);
or U12963 (N_12963,N_12785,N_12783);
xor U12964 (N_12964,N_12758,N_12780);
or U12965 (N_12965,N_12772,N_12765);
nor U12966 (N_12966,N_12607,N_12755);
xnor U12967 (N_12967,N_12608,N_12799);
nor U12968 (N_12968,N_12778,N_12732);
nor U12969 (N_12969,N_12629,N_12783);
and U12970 (N_12970,N_12702,N_12671);
nor U12971 (N_12971,N_12794,N_12762);
xnor U12972 (N_12972,N_12672,N_12690);
nand U12973 (N_12973,N_12620,N_12632);
xor U12974 (N_12974,N_12763,N_12715);
or U12975 (N_12975,N_12733,N_12600);
or U12976 (N_12976,N_12711,N_12669);
nand U12977 (N_12977,N_12621,N_12613);
and U12978 (N_12978,N_12638,N_12628);
and U12979 (N_12979,N_12646,N_12639);
xnor U12980 (N_12980,N_12690,N_12728);
nor U12981 (N_12981,N_12634,N_12785);
nand U12982 (N_12982,N_12776,N_12607);
nor U12983 (N_12983,N_12794,N_12695);
nand U12984 (N_12984,N_12782,N_12685);
nand U12985 (N_12985,N_12698,N_12717);
nand U12986 (N_12986,N_12613,N_12612);
xor U12987 (N_12987,N_12601,N_12755);
nor U12988 (N_12988,N_12659,N_12611);
and U12989 (N_12989,N_12674,N_12763);
or U12990 (N_12990,N_12607,N_12692);
and U12991 (N_12991,N_12721,N_12748);
and U12992 (N_12992,N_12673,N_12662);
nand U12993 (N_12993,N_12792,N_12681);
or U12994 (N_12994,N_12602,N_12780);
nand U12995 (N_12995,N_12728,N_12609);
or U12996 (N_12996,N_12794,N_12660);
and U12997 (N_12997,N_12756,N_12797);
or U12998 (N_12998,N_12712,N_12668);
nand U12999 (N_12999,N_12613,N_12706);
and U13000 (N_13000,N_12880,N_12947);
and U13001 (N_13001,N_12966,N_12992);
or U13002 (N_13002,N_12924,N_12824);
xnor U13003 (N_13003,N_12934,N_12949);
nand U13004 (N_13004,N_12987,N_12856);
nand U13005 (N_13005,N_12877,N_12915);
nand U13006 (N_13006,N_12845,N_12883);
and U13007 (N_13007,N_12882,N_12878);
and U13008 (N_13008,N_12954,N_12933);
xnor U13009 (N_13009,N_12980,N_12831);
or U13010 (N_13010,N_12900,N_12993);
nand U13011 (N_13011,N_12998,N_12996);
or U13012 (N_13012,N_12836,N_12879);
nand U13013 (N_13013,N_12800,N_12846);
xnor U13014 (N_13014,N_12852,N_12837);
nand U13015 (N_13015,N_12827,N_12896);
or U13016 (N_13016,N_12973,N_12972);
nor U13017 (N_13017,N_12862,N_12854);
nor U13018 (N_13018,N_12943,N_12884);
nand U13019 (N_13019,N_12974,N_12811);
nor U13020 (N_13020,N_12893,N_12959);
xnor U13021 (N_13021,N_12995,N_12835);
nand U13022 (N_13022,N_12841,N_12940);
xor U13023 (N_13023,N_12855,N_12806);
and U13024 (N_13024,N_12988,N_12953);
xnor U13025 (N_13025,N_12812,N_12948);
nor U13026 (N_13026,N_12925,N_12999);
xor U13027 (N_13027,N_12919,N_12802);
nand U13028 (N_13028,N_12994,N_12826);
and U13029 (N_13029,N_12945,N_12901);
or U13030 (N_13030,N_12834,N_12931);
or U13031 (N_13031,N_12939,N_12898);
xnor U13032 (N_13032,N_12829,N_12905);
xor U13033 (N_13033,N_12981,N_12808);
xor U13034 (N_13034,N_12902,N_12894);
xor U13035 (N_13035,N_12935,N_12873);
xor U13036 (N_13036,N_12912,N_12911);
and U13037 (N_13037,N_12897,N_12985);
nor U13038 (N_13038,N_12967,N_12871);
or U13039 (N_13039,N_12864,N_12918);
and U13040 (N_13040,N_12929,N_12810);
xnor U13041 (N_13041,N_12916,N_12844);
or U13042 (N_13042,N_12840,N_12874);
nand U13043 (N_13043,N_12865,N_12869);
and U13044 (N_13044,N_12923,N_12984);
and U13045 (N_13045,N_12801,N_12930);
and U13046 (N_13046,N_12858,N_12842);
or U13047 (N_13047,N_12926,N_12809);
xor U13048 (N_13048,N_12885,N_12821);
and U13049 (N_13049,N_12965,N_12921);
and U13050 (N_13050,N_12991,N_12820);
nor U13051 (N_13051,N_12850,N_12927);
nor U13052 (N_13052,N_12803,N_12964);
or U13053 (N_13053,N_12853,N_12906);
xnor U13054 (N_13054,N_12956,N_12848);
and U13055 (N_13055,N_12822,N_12859);
xor U13056 (N_13056,N_12963,N_12867);
nor U13057 (N_13057,N_12932,N_12920);
or U13058 (N_13058,N_12895,N_12955);
and U13059 (N_13059,N_12909,N_12922);
nor U13060 (N_13060,N_12832,N_12818);
nor U13061 (N_13061,N_12899,N_12975);
or U13062 (N_13062,N_12870,N_12961);
nand U13063 (N_13063,N_12989,N_12969);
xor U13064 (N_13064,N_12807,N_12887);
and U13065 (N_13065,N_12971,N_12952);
nor U13066 (N_13066,N_12942,N_12891);
nand U13067 (N_13067,N_12866,N_12982);
or U13068 (N_13068,N_12825,N_12881);
or U13069 (N_13069,N_12908,N_12805);
xor U13070 (N_13070,N_12814,N_12946);
or U13071 (N_13071,N_12978,N_12983);
and U13072 (N_13072,N_12857,N_12913);
xor U13073 (N_13073,N_12819,N_12907);
or U13074 (N_13074,N_12828,N_12977);
and U13075 (N_13075,N_12888,N_12839);
or U13076 (N_13076,N_12970,N_12892);
nand U13077 (N_13077,N_12804,N_12950);
or U13078 (N_13078,N_12875,N_12860);
or U13079 (N_13079,N_12816,N_12889);
xnor U13080 (N_13080,N_12851,N_12968);
nand U13081 (N_13081,N_12928,N_12890);
nand U13082 (N_13082,N_12843,N_12847);
and U13083 (N_13083,N_12817,N_12815);
and U13084 (N_13084,N_12938,N_12979);
and U13085 (N_13085,N_12941,N_12951);
xnor U13086 (N_13086,N_12876,N_12838);
and U13087 (N_13087,N_12960,N_12997);
nand U13088 (N_13088,N_12910,N_12936);
xor U13089 (N_13089,N_12886,N_12833);
nor U13090 (N_13090,N_12990,N_12904);
nor U13091 (N_13091,N_12976,N_12917);
nand U13092 (N_13092,N_12872,N_12849);
nand U13093 (N_13093,N_12914,N_12962);
and U13094 (N_13094,N_12823,N_12813);
xnor U13095 (N_13095,N_12986,N_12937);
xnor U13096 (N_13096,N_12863,N_12830);
nor U13097 (N_13097,N_12944,N_12868);
nor U13098 (N_13098,N_12903,N_12958);
nand U13099 (N_13099,N_12861,N_12957);
xor U13100 (N_13100,N_12883,N_12996);
or U13101 (N_13101,N_12969,N_12999);
nand U13102 (N_13102,N_12869,N_12986);
xor U13103 (N_13103,N_12808,N_12950);
xnor U13104 (N_13104,N_12995,N_12963);
nor U13105 (N_13105,N_12939,N_12960);
xnor U13106 (N_13106,N_12941,N_12955);
and U13107 (N_13107,N_12932,N_12885);
nor U13108 (N_13108,N_12852,N_12918);
or U13109 (N_13109,N_12813,N_12933);
or U13110 (N_13110,N_12965,N_12833);
xnor U13111 (N_13111,N_12971,N_12983);
or U13112 (N_13112,N_12855,N_12847);
nor U13113 (N_13113,N_12811,N_12843);
xor U13114 (N_13114,N_12807,N_12894);
xor U13115 (N_13115,N_12972,N_12899);
nor U13116 (N_13116,N_12917,N_12942);
xnor U13117 (N_13117,N_12821,N_12931);
and U13118 (N_13118,N_12935,N_12884);
or U13119 (N_13119,N_12867,N_12825);
nand U13120 (N_13120,N_12838,N_12971);
nor U13121 (N_13121,N_12861,N_12835);
nor U13122 (N_13122,N_12941,N_12836);
or U13123 (N_13123,N_12941,N_12964);
xor U13124 (N_13124,N_12872,N_12848);
and U13125 (N_13125,N_12854,N_12964);
nor U13126 (N_13126,N_12999,N_12929);
nor U13127 (N_13127,N_12991,N_12953);
and U13128 (N_13128,N_12940,N_12922);
or U13129 (N_13129,N_12913,N_12992);
xnor U13130 (N_13130,N_12875,N_12812);
xor U13131 (N_13131,N_12927,N_12888);
or U13132 (N_13132,N_12814,N_12937);
xor U13133 (N_13133,N_12820,N_12875);
and U13134 (N_13134,N_12941,N_12965);
xnor U13135 (N_13135,N_12981,N_12803);
nand U13136 (N_13136,N_12866,N_12962);
xnor U13137 (N_13137,N_12844,N_12984);
and U13138 (N_13138,N_12982,N_12901);
nand U13139 (N_13139,N_12949,N_12962);
xnor U13140 (N_13140,N_12994,N_12910);
nor U13141 (N_13141,N_12843,N_12903);
or U13142 (N_13142,N_12927,N_12981);
or U13143 (N_13143,N_12981,N_12817);
xor U13144 (N_13144,N_12858,N_12912);
xor U13145 (N_13145,N_12926,N_12968);
nand U13146 (N_13146,N_12939,N_12881);
xnor U13147 (N_13147,N_12864,N_12952);
nand U13148 (N_13148,N_12805,N_12930);
nand U13149 (N_13149,N_12915,N_12917);
nor U13150 (N_13150,N_12808,N_12818);
and U13151 (N_13151,N_12998,N_12967);
or U13152 (N_13152,N_12941,N_12864);
or U13153 (N_13153,N_12984,N_12961);
and U13154 (N_13154,N_12826,N_12975);
or U13155 (N_13155,N_12894,N_12851);
nor U13156 (N_13156,N_12904,N_12873);
or U13157 (N_13157,N_12879,N_12866);
nor U13158 (N_13158,N_12941,N_12892);
nor U13159 (N_13159,N_12986,N_12835);
and U13160 (N_13160,N_12852,N_12863);
nand U13161 (N_13161,N_12975,N_12848);
nand U13162 (N_13162,N_12826,N_12977);
xnor U13163 (N_13163,N_12998,N_12828);
and U13164 (N_13164,N_12828,N_12965);
or U13165 (N_13165,N_12914,N_12811);
nor U13166 (N_13166,N_12852,N_12825);
xor U13167 (N_13167,N_12955,N_12894);
and U13168 (N_13168,N_12933,N_12849);
or U13169 (N_13169,N_12800,N_12996);
or U13170 (N_13170,N_12834,N_12820);
and U13171 (N_13171,N_12851,N_12971);
nor U13172 (N_13172,N_12844,N_12959);
nand U13173 (N_13173,N_12823,N_12827);
or U13174 (N_13174,N_12931,N_12896);
nand U13175 (N_13175,N_12803,N_12914);
or U13176 (N_13176,N_12899,N_12852);
or U13177 (N_13177,N_12963,N_12916);
nor U13178 (N_13178,N_12999,N_12872);
xor U13179 (N_13179,N_12810,N_12890);
and U13180 (N_13180,N_12910,N_12981);
or U13181 (N_13181,N_12965,N_12917);
or U13182 (N_13182,N_12823,N_12821);
nand U13183 (N_13183,N_12801,N_12803);
or U13184 (N_13184,N_12928,N_12974);
and U13185 (N_13185,N_12931,N_12873);
nand U13186 (N_13186,N_12968,N_12892);
xor U13187 (N_13187,N_12831,N_12810);
or U13188 (N_13188,N_12809,N_12994);
and U13189 (N_13189,N_12958,N_12848);
xnor U13190 (N_13190,N_12940,N_12872);
nand U13191 (N_13191,N_12918,N_12963);
and U13192 (N_13192,N_12973,N_12935);
nor U13193 (N_13193,N_12850,N_12900);
and U13194 (N_13194,N_12879,N_12960);
xor U13195 (N_13195,N_12946,N_12982);
xor U13196 (N_13196,N_12897,N_12878);
nand U13197 (N_13197,N_12846,N_12985);
xnor U13198 (N_13198,N_12963,N_12954);
or U13199 (N_13199,N_12963,N_12990);
or U13200 (N_13200,N_13186,N_13112);
xnor U13201 (N_13201,N_13180,N_13148);
nor U13202 (N_13202,N_13096,N_13028);
or U13203 (N_13203,N_13077,N_13059);
nor U13204 (N_13204,N_13197,N_13018);
nor U13205 (N_13205,N_13058,N_13139);
nor U13206 (N_13206,N_13183,N_13167);
or U13207 (N_13207,N_13142,N_13178);
or U13208 (N_13208,N_13128,N_13061);
nand U13209 (N_13209,N_13118,N_13045);
or U13210 (N_13210,N_13157,N_13029);
or U13211 (N_13211,N_13198,N_13038);
or U13212 (N_13212,N_13001,N_13084);
and U13213 (N_13213,N_13026,N_13199);
or U13214 (N_13214,N_13039,N_13016);
and U13215 (N_13215,N_13185,N_13133);
nand U13216 (N_13216,N_13085,N_13131);
xnor U13217 (N_13217,N_13187,N_13170);
xor U13218 (N_13218,N_13005,N_13093);
or U13219 (N_13219,N_13177,N_13068);
or U13220 (N_13220,N_13046,N_13071);
nand U13221 (N_13221,N_13136,N_13175);
or U13222 (N_13222,N_13168,N_13098);
or U13223 (N_13223,N_13044,N_13114);
or U13224 (N_13224,N_13036,N_13094);
xor U13225 (N_13225,N_13134,N_13022);
nand U13226 (N_13226,N_13060,N_13126);
or U13227 (N_13227,N_13057,N_13123);
xor U13228 (N_13228,N_13152,N_13158);
nor U13229 (N_13229,N_13056,N_13172);
nor U13230 (N_13230,N_13115,N_13006);
or U13231 (N_13231,N_13159,N_13109);
or U13232 (N_13232,N_13047,N_13055);
nand U13233 (N_13233,N_13135,N_13087);
or U13234 (N_13234,N_13020,N_13196);
nor U13235 (N_13235,N_13017,N_13064);
xor U13236 (N_13236,N_13014,N_13154);
nand U13237 (N_13237,N_13082,N_13081);
and U13238 (N_13238,N_13011,N_13153);
or U13239 (N_13239,N_13143,N_13145);
xnor U13240 (N_13240,N_13156,N_13176);
and U13241 (N_13241,N_13032,N_13065);
nand U13242 (N_13242,N_13138,N_13063);
nor U13243 (N_13243,N_13160,N_13141);
and U13244 (N_13244,N_13000,N_13174);
and U13245 (N_13245,N_13072,N_13151);
xnor U13246 (N_13246,N_13002,N_13019);
nor U13247 (N_13247,N_13182,N_13099);
nor U13248 (N_13248,N_13088,N_13091);
nand U13249 (N_13249,N_13035,N_13078);
and U13250 (N_13250,N_13147,N_13015);
xnor U13251 (N_13251,N_13116,N_13052);
xor U13252 (N_13252,N_13073,N_13010);
or U13253 (N_13253,N_13075,N_13054);
nand U13254 (N_13254,N_13106,N_13119);
xor U13255 (N_13255,N_13100,N_13130);
or U13256 (N_13256,N_13169,N_13129);
nor U13257 (N_13257,N_13149,N_13009);
nand U13258 (N_13258,N_13103,N_13101);
and U13259 (N_13259,N_13092,N_13097);
xnor U13260 (N_13260,N_13021,N_13121);
or U13261 (N_13261,N_13108,N_13188);
and U13262 (N_13262,N_13181,N_13003);
nor U13263 (N_13263,N_13086,N_13195);
and U13264 (N_13264,N_13074,N_13102);
nand U13265 (N_13265,N_13164,N_13166);
and U13266 (N_13266,N_13155,N_13132);
or U13267 (N_13267,N_13191,N_13194);
nor U13268 (N_13268,N_13111,N_13179);
or U13269 (N_13269,N_13049,N_13069);
and U13270 (N_13270,N_13033,N_13146);
nand U13271 (N_13271,N_13037,N_13189);
and U13272 (N_13272,N_13013,N_13004);
nor U13273 (N_13273,N_13062,N_13070);
nor U13274 (N_13274,N_13163,N_13083);
nand U13275 (N_13275,N_13023,N_13104);
nor U13276 (N_13276,N_13125,N_13090);
nor U13277 (N_13277,N_13161,N_13079);
and U13278 (N_13278,N_13105,N_13192);
nor U13279 (N_13279,N_13173,N_13171);
xnor U13280 (N_13280,N_13165,N_13050);
nor U13281 (N_13281,N_13190,N_13067);
nand U13282 (N_13282,N_13053,N_13008);
xor U13283 (N_13283,N_13041,N_13031);
or U13284 (N_13284,N_13124,N_13117);
nor U13285 (N_13285,N_13120,N_13080);
nor U13286 (N_13286,N_13150,N_13043);
xnor U13287 (N_13287,N_13113,N_13030);
and U13288 (N_13288,N_13076,N_13024);
and U13289 (N_13289,N_13127,N_13027);
and U13290 (N_13290,N_13122,N_13110);
xor U13291 (N_13291,N_13162,N_13042);
and U13292 (N_13292,N_13095,N_13089);
nor U13293 (N_13293,N_13140,N_13066);
xnor U13294 (N_13294,N_13144,N_13137);
or U13295 (N_13295,N_13184,N_13048);
xor U13296 (N_13296,N_13012,N_13051);
xor U13297 (N_13297,N_13007,N_13034);
nand U13298 (N_13298,N_13040,N_13193);
and U13299 (N_13299,N_13025,N_13107);
xnor U13300 (N_13300,N_13076,N_13194);
nor U13301 (N_13301,N_13038,N_13162);
and U13302 (N_13302,N_13167,N_13011);
nand U13303 (N_13303,N_13182,N_13002);
and U13304 (N_13304,N_13076,N_13086);
nand U13305 (N_13305,N_13145,N_13054);
nand U13306 (N_13306,N_13167,N_13191);
nand U13307 (N_13307,N_13050,N_13152);
nand U13308 (N_13308,N_13036,N_13101);
nand U13309 (N_13309,N_13068,N_13013);
and U13310 (N_13310,N_13007,N_13133);
and U13311 (N_13311,N_13050,N_13090);
or U13312 (N_13312,N_13077,N_13139);
xor U13313 (N_13313,N_13144,N_13085);
nand U13314 (N_13314,N_13027,N_13002);
nor U13315 (N_13315,N_13156,N_13092);
and U13316 (N_13316,N_13034,N_13073);
or U13317 (N_13317,N_13186,N_13089);
and U13318 (N_13318,N_13144,N_13045);
nand U13319 (N_13319,N_13165,N_13176);
and U13320 (N_13320,N_13093,N_13095);
and U13321 (N_13321,N_13111,N_13066);
nand U13322 (N_13322,N_13006,N_13058);
and U13323 (N_13323,N_13039,N_13060);
or U13324 (N_13324,N_13007,N_13103);
nand U13325 (N_13325,N_13058,N_13180);
nand U13326 (N_13326,N_13108,N_13091);
or U13327 (N_13327,N_13145,N_13152);
nor U13328 (N_13328,N_13190,N_13151);
nor U13329 (N_13329,N_13011,N_13137);
nand U13330 (N_13330,N_13164,N_13030);
nand U13331 (N_13331,N_13079,N_13056);
nand U13332 (N_13332,N_13169,N_13025);
xnor U13333 (N_13333,N_13032,N_13064);
and U13334 (N_13334,N_13026,N_13022);
xor U13335 (N_13335,N_13111,N_13184);
xnor U13336 (N_13336,N_13020,N_13007);
and U13337 (N_13337,N_13145,N_13105);
nand U13338 (N_13338,N_13010,N_13049);
xnor U13339 (N_13339,N_13180,N_13086);
nand U13340 (N_13340,N_13099,N_13057);
and U13341 (N_13341,N_13139,N_13123);
nand U13342 (N_13342,N_13053,N_13046);
nand U13343 (N_13343,N_13086,N_13079);
xor U13344 (N_13344,N_13102,N_13093);
nand U13345 (N_13345,N_13185,N_13003);
nand U13346 (N_13346,N_13060,N_13166);
nand U13347 (N_13347,N_13062,N_13130);
xor U13348 (N_13348,N_13001,N_13086);
and U13349 (N_13349,N_13039,N_13077);
nand U13350 (N_13350,N_13159,N_13125);
and U13351 (N_13351,N_13142,N_13143);
nor U13352 (N_13352,N_13155,N_13093);
nand U13353 (N_13353,N_13061,N_13039);
and U13354 (N_13354,N_13096,N_13158);
or U13355 (N_13355,N_13075,N_13112);
nand U13356 (N_13356,N_13091,N_13093);
xnor U13357 (N_13357,N_13176,N_13151);
nand U13358 (N_13358,N_13178,N_13090);
and U13359 (N_13359,N_13027,N_13138);
or U13360 (N_13360,N_13080,N_13032);
nand U13361 (N_13361,N_13083,N_13141);
xor U13362 (N_13362,N_13011,N_13179);
nor U13363 (N_13363,N_13195,N_13109);
or U13364 (N_13364,N_13046,N_13171);
nor U13365 (N_13365,N_13178,N_13168);
nor U13366 (N_13366,N_13123,N_13120);
or U13367 (N_13367,N_13078,N_13045);
nor U13368 (N_13368,N_13091,N_13101);
xnor U13369 (N_13369,N_13102,N_13103);
or U13370 (N_13370,N_13015,N_13181);
and U13371 (N_13371,N_13053,N_13030);
or U13372 (N_13372,N_13152,N_13111);
and U13373 (N_13373,N_13166,N_13059);
and U13374 (N_13374,N_13098,N_13174);
nand U13375 (N_13375,N_13047,N_13060);
and U13376 (N_13376,N_13063,N_13083);
and U13377 (N_13377,N_13134,N_13106);
and U13378 (N_13378,N_13077,N_13053);
and U13379 (N_13379,N_13164,N_13063);
and U13380 (N_13380,N_13123,N_13036);
and U13381 (N_13381,N_13180,N_13163);
and U13382 (N_13382,N_13064,N_13104);
xnor U13383 (N_13383,N_13093,N_13110);
xor U13384 (N_13384,N_13194,N_13183);
xor U13385 (N_13385,N_13004,N_13109);
xor U13386 (N_13386,N_13158,N_13197);
nand U13387 (N_13387,N_13116,N_13033);
or U13388 (N_13388,N_13081,N_13186);
or U13389 (N_13389,N_13053,N_13050);
or U13390 (N_13390,N_13190,N_13065);
nand U13391 (N_13391,N_13175,N_13003);
and U13392 (N_13392,N_13025,N_13019);
xnor U13393 (N_13393,N_13102,N_13006);
xor U13394 (N_13394,N_13186,N_13046);
xnor U13395 (N_13395,N_13098,N_13154);
or U13396 (N_13396,N_13020,N_13155);
or U13397 (N_13397,N_13071,N_13198);
nand U13398 (N_13398,N_13043,N_13031);
and U13399 (N_13399,N_13062,N_13152);
nand U13400 (N_13400,N_13389,N_13266);
and U13401 (N_13401,N_13205,N_13380);
nand U13402 (N_13402,N_13385,N_13375);
and U13403 (N_13403,N_13364,N_13356);
nor U13404 (N_13404,N_13298,N_13286);
nor U13405 (N_13405,N_13297,N_13365);
xnor U13406 (N_13406,N_13395,N_13273);
xnor U13407 (N_13407,N_13347,N_13235);
xor U13408 (N_13408,N_13346,N_13256);
or U13409 (N_13409,N_13315,N_13249);
xor U13410 (N_13410,N_13383,N_13329);
nor U13411 (N_13411,N_13338,N_13353);
xor U13412 (N_13412,N_13220,N_13306);
nor U13413 (N_13413,N_13251,N_13330);
xor U13414 (N_13414,N_13366,N_13291);
nor U13415 (N_13415,N_13336,N_13254);
xnor U13416 (N_13416,N_13340,N_13283);
or U13417 (N_13417,N_13326,N_13225);
or U13418 (N_13418,N_13374,N_13281);
nand U13419 (N_13419,N_13371,N_13320);
or U13420 (N_13420,N_13224,N_13222);
and U13421 (N_13421,N_13337,N_13305);
nand U13422 (N_13422,N_13233,N_13206);
or U13423 (N_13423,N_13323,N_13360);
nand U13424 (N_13424,N_13212,N_13332);
or U13425 (N_13425,N_13282,N_13357);
xnor U13426 (N_13426,N_13342,N_13341);
nand U13427 (N_13427,N_13334,N_13362);
nand U13428 (N_13428,N_13232,N_13200);
or U13429 (N_13429,N_13361,N_13317);
nand U13430 (N_13430,N_13269,N_13230);
or U13431 (N_13431,N_13234,N_13372);
nor U13432 (N_13432,N_13214,N_13302);
and U13433 (N_13433,N_13388,N_13208);
or U13434 (N_13434,N_13335,N_13275);
and U13435 (N_13435,N_13253,N_13271);
xnor U13436 (N_13436,N_13373,N_13384);
nor U13437 (N_13437,N_13240,N_13242);
xor U13438 (N_13438,N_13310,N_13252);
or U13439 (N_13439,N_13239,N_13348);
or U13440 (N_13440,N_13217,N_13327);
or U13441 (N_13441,N_13203,N_13278);
xor U13442 (N_13442,N_13370,N_13322);
and U13443 (N_13443,N_13243,N_13300);
nor U13444 (N_13444,N_13295,N_13277);
or U13445 (N_13445,N_13287,N_13210);
or U13446 (N_13446,N_13363,N_13241);
or U13447 (N_13447,N_13279,N_13316);
and U13448 (N_13448,N_13379,N_13226);
and U13449 (N_13449,N_13245,N_13309);
nand U13450 (N_13450,N_13301,N_13328);
xor U13451 (N_13451,N_13213,N_13285);
nor U13452 (N_13452,N_13274,N_13261);
and U13453 (N_13453,N_13223,N_13311);
xnor U13454 (N_13454,N_13263,N_13288);
xor U13455 (N_13455,N_13387,N_13321);
and U13456 (N_13456,N_13262,N_13207);
nand U13457 (N_13457,N_13238,N_13228);
nor U13458 (N_13458,N_13313,N_13378);
and U13459 (N_13459,N_13294,N_13381);
nand U13460 (N_13460,N_13382,N_13229);
or U13461 (N_13461,N_13276,N_13308);
or U13462 (N_13462,N_13358,N_13218);
or U13463 (N_13463,N_13202,N_13258);
xor U13464 (N_13464,N_13345,N_13244);
xor U13465 (N_13465,N_13349,N_13284);
nor U13466 (N_13466,N_13216,N_13369);
nand U13467 (N_13467,N_13394,N_13339);
or U13468 (N_13468,N_13270,N_13355);
and U13469 (N_13469,N_13221,N_13272);
or U13470 (N_13470,N_13376,N_13350);
xor U13471 (N_13471,N_13280,N_13391);
nand U13472 (N_13472,N_13259,N_13333);
nand U13473 (N_13473,N_13246,N_13307);
or U13474 (N_13474,N_13359,N_13292);
or U13475 (N_13475,N_13265,N_13377);
and U13476 (N_13476,N_13344,N_13397);
nor U13477 (N_13477,N_13215,N_13264);
or U13478 (N_13478,N_13318,N_13236);
or U13479 (N_13479,N_13260,N_13352);
xor U13480 (N_13480,N_13324,N_13290);
nor U13481 (N_13481,N_13392,N_13325);
xor U13482 (N_13482,N_13398,N_13201);
or U13483 (N_13483,N_13289,N_13331);
nand U13484 (N_13484,N_13250,N_13268);
xnor U13485 (N_13485,N_13396,N_13367);
nor U13486 (N_13486,N_13257,N_13303);
and U13487 (N_13487,N_13267,N_13319);
nor U13488 (N_13488,N_13390,N_13237);
nor U13489 (N_13489,N_13227,N_13304);
xor U13490 (N_13490,N_13393,N_13209);
or U13491 (N_13491,N_13368,N_13293);
or U13492 (N_13492,N_13296,N_13211);
and U13493 (N_13493,N_13386,N_13231);
or U13494 (N_13494,N_13248,N_13204);
or U13495 (N_13495,N_13312,N_13399);
xnor U13496 (N_13496,N_13219,N_13314);
nor U13497 (N_13497,N_13351,N_13343);
xor U13498 (N_13498,N_13299,N_13247);
or U13499 (N_13499,N_13255,N_13354);
nand U13500 (N_13500,N_13231,N_13303);
nand U13501 (N_13501,N_13356,N_13338);
nand U13502 (N_13502,N_13379,N_13377);
nand U13503 (N_13503,N_13361,N_13369);
or U13504 (N_13504,N_13274,N_13355);
nor U13505 (N_13505,N_13341,N_13344);
or U13506 (N_13506,N_13307,N_13264);
xnor U13507 (N_13507,N_13223,N_13236);
nand U13508 (N_13508,N_13218,N_13268);
nor U13509 (N_13509,N_13285,N_13315);
nor U13510 (N_13510,N_13352,N_13270);
nor U13511 (N_13511,N_13328,N_13283);
or U13512 (N_13512,N_13291,N_13274);
and U13513 (N_13513,N_13234,N_13290);
xnor U13514 (N_13514,N_13318,N_13275);
or U13515 (N_13515,N_13242,N_13266);
and U13516 (N_13516,N_13240,N_13360);
nor U13517 (N_13517,N_13253,N_13317);
nand U13518 (N_13518,N_13225,N_13268);
or U13519 (N_13519,N_13356,N_13316);
nor U13520 (N_13520,N_13297,N_13314);
and U13521 (N_13521,N_13355,N_13348);
nor U13522 (N_13522,N_13254,N_13217);
xor U13523 (N_13523,N_13223,N_13238);
nor U13524 (N_13524,N_13293,N_13262);
and U13525 (N_13525,N_13366,N_13322);
nor U13526 (N_13526,N_13347,N_13373);
nand U13527 (N_13527,N_13206,N_13310);
nand U13528 (N_13528,N_13255,N_13220);
nor U13529 (N_13529,N_13383,N_13327);
or U13530 (N_13530,N_13248,N_13342);
and U13531 (N_13531,N_13306,N_13363);
nor U13532 (N_13532,N_13317,N_13299);
xor U13533 (N_13533,N_13353,N_13246);
xnor U13534 (N_13534,N_13367,N_13246);
nor U13535 (N_13535,N_13251,N_13300);
and U13536 (N_13536,N_13275,N_13305);
nor U13537 (N_13537,N_13310,N_13303);
nor U13538 (N_13538,N_13329,N_13363);
nand U13539 (N_13539,N_13391,N_13275);
nand U13540 (N_13540,N_13227,N_13377);
nor U13541 (N_13541,N_13306,N_13341);
nand U13542 (N_13542,N_13317,N_13385);
nand U13543 (N_13543,N_13293,N_13220);
nand U13544 (N_13544,N_13215,N_13393);
and U13545 (N_13545,N_13375,N_13386);
nor U13546 (N_13546,N_13354,N_13270);
or U13547 (N_13547,N_13390,N_13368);
xnor U13548 (N_13548,N_13206,N_13229);
or U13549 (N_13549,N_13291,N_13375);
or U13550 (N_13550,N_13289,N_13349);
nand U13551 (N_13551,N_13207,N_13381);
and U13552 (N_13552,N_13247,N_13248);
nand U13553 (N_13553,N_13265,N_13231);
xnor U13554 (N_13554,N_13266,N_13293);
xnor U13555 (N_13555,N_13331,N_13386);
xnor U13556 (N_13556,N_13313,N_13264);
xnor U13557 (N_13557,N_13249,N_13356);
nor U13558 (N_13558,N_13268,N_13341);
xnor U13559 (N_13559,N_13298,N_13292);
nand U13560 (N_13560,N_13344,N_13294);
or U13561 (N_13561,N_13329,N_13330);
nor U13562 (N_13562,N_13222,N_13346);
nor U13563 (N_13563,N_13275,N_13384);
xnor U13564 (N_13564,N_13368,N_13381);
xnor U13565 (N_13565,N_13371,N_13398);
xnor U13566 (N_13566,N_13260,N_13373);
nor U13567 (N_13567,N_13309,N_13272);
nor U13568 (N_13568,N_13318,N_13242);
and U13569 (N_13569,N_13328,N_13229);
nor U13570 (N_13570,N_13255,N_13315);
nor U13571 (N_13571,N_13274,N_13374);
and U13572 (N_13572,N_13234,N_13257);
nor U13573 (N_13573,N_13374,N_13272);
and U13574 (N_13574,N_13307,N_13375);
or U13575 (N_13575,N_13286,N_13304);
and U13576 (N_13576,N_13215,N_13230);
nand U13577 (N_13577,N_13255,N_13392);
or U13578 (N_13578,N_13241,N_13398);
nand U13579 (N_13579,N_13393,N_13370);
nand U13580 (N_13580,N_13257,N_13243);
nand U13581 (N_13581,N_13339,N_13256);
nand U13582 (N_13582,N_13333,N_13238);
nand U13583 (N_13583,N_13252,N_13292);
and U13584 (N_13584,N_13304,N_13325);
nor U13585 (N_13585,N_13335,N_13295);
nand U13586 (N_13586,N_13338,N_13347);
xor U13587 (N_13587,N_13317,N_13282);
nand U13588 (N_13588,N_13368,N_13321);
or U13589 (N_13589,N_13294,N_13312);
and U13590 (N_13590,N_13380,N_13290);
xor U13591 (N_13591,N_13332,N_13254);
nor U13592 (N_13592,N_13296,N_13208);
nand U13593 (N_13593,N_13364,N_13345);
nor U13594 (N_13594,N_13384,N_13322);
xor U13595 (N_13595,N_13211,N_13278);
and U13596 (N_13596,N_13280,N_13373);
nand U13597 (N_13597,N_13205,N_13342);
or U13598 (N_13598,N_13212,N_13237);
or U13599 (N_13599,N_13217,N_13260);
and U13600 (N_13600,N_13426,N_13540);
or U13601 (N_13601,N_13462,N_13407);
nor U13602 (N_13602,N_13406,N_13457);
nand U13603 (N_13603,N_13423,N_13566);
nor U13604 (N_13604,N_13469,N_13508);
or U13605 (N_13605,N_13560,N_13484);
and U13606 (N_13606,N_13455,N_13551);
xnor U13607 (N_13607,N_13420,N_13465);
or U13608 (N_13608,N_13432,N_13539);
or U13609 (N_13609,N_13576,N_13449);
or U13610 (N_13610,N_13417,N_13403);
and U13611 (N_13611,N_13519,N_13439);
xnor U13612 (N_13612,N_13411,N_13541);
and U13613 (N_13613,N_13518,N_13435);
nor U13614 (N_13614,N_13582,N_13436);
nand U13615 (N_13615,N_13425,N_13450);
nor U13616 (N_13616,N_13486,N_13590);
xor U13617 (N_13617,N_13568,N_13485);
or U13618 (N_13618,N_13434,N_13599);
or U13619 (N_13619,N_13507,N_13563);
or U13620 (N_13620,N_13546,N_13448);
and U13621 (N_13621,N_13553,N_13452);
nand U13622 (N_13622,N_13467,N_13476);
and U13623 (N_13623,N_13475,N_13575);
or U13624 (N_13624,N_13556,N_13506);
nand U13625 (N_13625,N_13483,N_13550);
nor U13626 (N_13626,N_13480,N_13535);
and U13627 (N_13627,N_13427,N_13438);
nor U13628 (N_13628,N_13409,N_13586);
and U13629 (N_13629,N_13474,N_13444);
nand U13630 (N_13630,N_13443,N_13445);
or U13631 (N_13631,N_13595,N_13543);
or U13632 (N_13632,N_13456,N_13559);
xor U13633 (N_13633,N_13433,N_13574);
xnor U13634 (N_13634,N_13419,N_13501);
xnor U13635 (N_13635,N_13562,N_13527);
xnor U13636 (N_13636,N_13515,N_13497);
nor U13637 (N_13637,N_13454,N_13493);
xnor U13638 (N_13638,N_13473,N_13405);
and U13639 (N_13639,N_13555,N_13533);
xnor U13640 (N_13640,N_13402,N_13463);
and U13641 (N_13641,N_13458,N_13557);
nor U13642 (N_13642,N_13513,N_13565);
xnor U13643 (N_13643,N_13431,N_13468);
nor U13644 (N_13644,N_13482,N_13464);
xnor U13645 (N_13645,N_13428,N_13471);
nor U13646 (N_13646,N_13549,N_13552);
nand U13647 (N_13647,N_13472,N_13544);
nand U13648 (N_13648,N_13422,N_13459);
nand U13649 (N_13649,N_13524,N_13412);
nand U13650 (N_13650,N_13470,N_13564);
or U13651 (N_13651,N_13440,N_13492);
nor U13652 (N_13652,N_13487,N_13538);
and U13653 (N_13653,N_13578,N_13509);
nand U13654 (N_13654,N_13542,N_13490);
nor U13655 (N_13655,N_13525,N_13430);
or U13656 (N_13656,N_13548,N_13481);
or U13657 (N_13657,N_13584,N_13596);
or U13658 (N_13658,N_13598,N_13570);
xnor U13659 (N_13659,N_13529,N_13442);
or U13660 (N_13660,N_13400,N_13413);
or U13661 (N_13661,N_13429,N_13453);
and U13662 (N_13662,N_13536,N_13477);
and U13663 (N_13663,N_13478,N_13588);
and U13664 (N_13664,N_13534,N_13577);
nand U13665 (N_13665,N_13567,N_13510);
nand U13666 (N_13666,N_13441,N_13528);
xor U13667 (N_13667,N_13516,N_13530);
or U13668 (N_13668,N_13437,N_13414);
or U13669 (N_13669,N_13505,N_13573);
nand U13670 (N_13670,N_13594,N_13491);
and U13671 (N_13671,N_13495,N_13421);
and U13672 (N_13672,N_13494,N_13593);
nand U13673 (N_13673,N_13526,N_13583);
nand U13674 (N_13674,N_13514,N_13503);
xnor U13675 (N_13675,N_13554,N_13488);
or U13676 (N_13676,N_13460,N_13580);
xnor U13677 (N_13677,N_13451,N_13523);
nand U13678 (N_13678,N_13558,N_13498);
nor U13679 (N_13679,N_13489,N_13466);
and U13680 (N_13680,N_13410,N_13500);
and U13681 (N_13681,N_13585,N_13446);
xor U13682 (N_13682,N_13502,N_13537);
xor U13683 (N_13683,N_13447,N_13520);
nor U13684 (N_13684,N_13517,N_13511);
and U13685 (N_13685,N_13512,N_13592);
nor U13686 (N_13686,N_13521,N_13561);
nor U13687 (N_13687,N_13499,N_13532);
xor U13688 (N_13688,N_13531,N_13496);
nand U13689 (N_13689,N_13581,N_13404);
and U13690 (N_13690,N_13547,N_13571);
nand U13691 (N_13691,N_13572,N_13418);
nand U13692 (N_13692,N_13408,N_13401);
nor U13693 (N_13693,N_13587,N_13591);
nand U13694 (N_13694,N_13579,N_13597);
xor U13695 (N_13695,N_13569,N_13504);
nand U13696 (N_13696,N_13416,N_13589);
xnor U13697 (N_13697,N_13415,N_13479);
xor U13698 (N_13698,N_13424,N_13545);
nand U13699 (N_13699,N_13522,N_13461);
and U13700 (N_13700,N_13508,N_13440);
xor U13701 (N_13701,N_13579,N_13580);
nand U13702 (N_13702,N_13512,N_13417);
nand U13703 (N_13703,N_13544,N_13489);
xnor U13704 (N_13704,N_13452,N_13500);
nor U13705 (N_13705,N_13524,N_13447);
or U13706 (N_13706,N_13591,N_13595);
and U13707 (N_13707,N_13565,N_13453);
or U13708 (N_13708,N_13476,N_13569);
and U13709 (N_13709,N_13444,N_13490);
and U13710 (N_13710,N_13494,N_13493);
xor U13711 (N_13711,N_13533,N_13426);
nand U13712 (N_13712,N_13415,N_13496);
or U13713 (N_13713,N_13486,N_13459);
nor U13714 (N_13714,N_13433,N_13430);
nand U13715 (N_13715,N_13405,N_13440);
nor U13716 (N_13716,N_13511,N_13423);
and U13717 (N_13717,N_13489,N_13502);
and U13718 (N_13718,N_13567,N_13557);
and U13719 (N_13719,N_13571,N_13444);
nor U13720 (N_13720,N_13526,N_13538);
nand U13721 (N_13721,N_13598,N_13434);
xnor U13722 (N_13722,N_13434,N_13417);
or U13723 (N_13723,N_13431,N_13518);
or U13724 (N_13724,N_13474,N_13485);
nand U13725 (N_13725,N_13488,N_13538);
nor U13726 (N_13726,N_13520,N_13598);
and U13727 (N_13727,N_13449,N_13517);
and U13728 (N_13728,N_13436,N_13517);
and U13729 (N_13729,N_13409,N_13589);
and U13730 (N_13730,N_13481,N_13589);
nand U13731 (N_13731,N_13495,N_13528);
nor U13732 (N_13732,N_13422,N_13472);
or U13733 (N_13733,N_13522,N_13575);
or U13734 (N_13734,N_13471,N_13490);
nand U13735 (N_13735,N_13577,N_13401);
or U13736 (N_13736,N_13515,N_13557);
and U13737 (N_13737,N_13472,N_13534);
nor U13738 (N_13738,N_13460,N_13512);
or U13739 (N_13739,N_13427,N_13524);
nor U13740 (N_13740,N_13538,N_13476);
and U13741 (N_13741,N_13597,N_13404);
or U13742 (N_13742,N_13497,N_13537);
nand U13743 (N_13743,N_13592,N_13467);
xnor U13744 (N_13744,N_13524,N_13590);
or U13745 (N_13745,N_13503,N_13482);
nand U13746 (N_13746,N_13404,N_13583);
xor U13747 (N_13747,N_13418,N_13450);
or U13748 (N_13748,N_13566,N_13593);
and U13749 (N_13749,N_13400,N_13545);
xnor U13750 (N_13750,N_13583,N_13436);
or U13751 (N_13751,N_13423,N_13537);
nand U13752 (N_13752,N_13517,N_13476);
or U13753 (N_13753,N_13437,N_13400);
nand U13754 (N_13754,N_13509,N_13503);
or U13755 (N_13755,N_13490,N_13543);
xor U13756 (N_13756,N_13413,N_13491);
nor U13757 (N_13757,N_13401,N_13451);
or U13758 (N_13758,N_13503,N_13401);
nor U13759 (N_13759,N_13420,N_13407);
xor U13760 (N_13760,N_13465,N_13497);
nor U13761 (N_13761,N_13503,N_13468);
xnor U13762 (N_13762,N_13428,N_13488);
and U13763 (N_13763,N_13460,N_13585);
and U13764 (N_13764,N_13504,N_13408);
xnor U13765 (N_13765,N_13565,N_13548);
xor U13766 (N_13766,N_13567,N_13484);
nor U13767 (N_13767,N_13497,N_13407);
or U13768 (N_13768,N_13404,N_13525);
nand U13769 (N_13769,N_13520,N_13464);
nand U13770 (N_13770,N_13458,N_13498);
or U13771 (N_13771,N_13538,N_13491);
xor U13772 (N_13772,N_13421,N_13548);
nand U13773 (N_13773,N_13494,N_13428);
nor U13774 (N_13774,N_13410,N_13556);
nand U13775 (N_13775,N_13593,N_13500);
and U13776 (N_13776,N_13577,N_13465);
or U13777 (N_13777,N_13587,N_13562);
and U13778 (N_13778,N_13461,N_13501);
xnor U13779 (N_13779,N_13467,N_13513);
or U13780 (N_13780,N_13461,N_13594);
nand U13781 (N_13781,N_13593,N_13525);
and U13782 (N_13782,N_13487,N_13521);
or U13783 (N_13783,N_13594,N_13509);
nor U13784 (N_13784,N_13503,N_13504);
nand U13785 (N_13785,N_13581,N_13550);
nand U13786 (N_13786,N_13454,N_13485);
and U13787 (N_13787,N_13567,N_13480);
nor U13788 (N_13788,N_13453,N_13535);
nor U13789 (N_13789,N_13517,N_13589);
nor U13790 (N_13790,N_13403,N_13450);
nor U13791 (N_13791,N_13456,N_13439);
and U13792 (N_13792,N_13499,N_13554);
xnor U13793 (N_13793,N_13421,N_13508);
or U13794 (N_13794,N_13484,N_13508);
nor U13795 (N_13795,N_13511,N_13524);
or U13796 (N_13796,N_13527,N_13550);
xnor U13797 (N_13797,N_13427,N_13569);
and U13798 (N_13798,N_13518,N_13526);
nand U13799 (N_13799,N_13578,N_13436);
nand U13800 (N_13800,N_13704,N_13777);
nor U13801 (N_13801,N_13635,N_13765);
or U13802 (N_13802,N_13657,N_13698);
xnor U13803 (N_13803,N_13606,N_13676);
nor U13804 (N_13804,N_13643,N_13671);
nor U13805 (N_13805,N_13736,N_13677);
nand U13806 (N_13806,N_13672,N_13733);
xnor U13807 (N_13807,N_13625,N_13660);
xor U13808 (N_13808,N_13726,N_13706);
nor U13809 (N_13809,N_13737,N_13757);
xor U13810 (N_13810,N_13682,N_13772);
nor U13811 (N_13811,N_13797,N_13692);
nor U13812 (N_13812,N_13709,N_13716);
nor U13813 (N_13813,N_13755,N_13613);
and U13814 (N_13814,N_13652,N_13750);
xnor U13815 (N_13815,N_13633,N_13749);
or U13816 (N_13816,N_13669,N_13723);
and U13817 (N_13817,N_13738,N_13612);
or U13818 (N_13818,N_13729,N_13794);
xor U13819 (N_13819,N_13761,N_13654);
or U13820 (N_13820,N_13775,N_13668);
nand U13821 (N_13821,N_13773,N_13611);
nand U13822 (N_13822,N_13776,N_13646);
nand U13823 (N_13823,N_13665,N_13715);
or U13824 (N_13824,N_13604,N_13770);
nor U13825 (N_13825,N_13684,N_13741);
nand U13826 (N_13826,N_13624,N_13616);
nand U13827 (N_13827,N_13666,N_13710);
or U13828 (N_13828,N_13694,N_13688);
nor U13829 (N_13829,N_13728,N_13629);
or U13830 (N_13830,N_13658,N_13703);
nor U13831 (N_13831,N_13744,N_13673);
or U13832 (N_13832,N_13605,N_13720);
nand U13833 (N_13833,N_13628,N_13711);
nand U13834 (N_13834,N_13696,N_13674);
nand U13835 (N_13835,N_13695,N_13735);
and U13836 (N_13836,N_13642,N_13748);
or U13837 (N_13837,N_13799,N_13621);
or U13838 (N_13838,N_13719,N_13640);
nor U13839 (N_13839,N_13742,N_13662);
and U13840 (N_13840,N_13762,N_13753);
nor U13841 (N_13841,N_13795,N_13650);
xor U13842 (N_13842,N_13705,N_13732);
and U13843 (N_13843,N_13649,N_13789);
or U13844 (N_13844,N_13766,N_13631);
and U13845 (N_13845,N_13615,N_13619);
or U13846 (N_13846,N_13796,N_13790);
nor U13847 (N_13847,N_13675,N_13683);
nand U13848 (N_13848,N_13632,N_13697);
nand U13849 (N_13849,N_13756,N_13620);
or U13850 (N_13850,N_13627,N_13681);
or U13851 (N_13851,N_13764,N_13734);
or U13852 (N_13852,N_13693,N_13641);
or U13853 (N_13853,N_13745,N_13712);
xor U13854 (N_13854,N_13622,N_13661);
nor U13855 (N_13855,N_13717,N_13699);
nor U13856 (N_13856,N_13780,N_13768);
nor U13857 (N_13857,N_13609,N_13667);
nor U13858 (N_13858,N_13691,N_13779);
or U13859 (N_13859,N_13751,N_13689);
and U13860 (N_13860,N_13739,N_13767);
nor U13861 (N_13861,N_13663,N_13784);
xor U13862 (N_13862,N_13608,N_13690);
nand U13863 (N_13863,N_13792,N_13786);
nand U13864 (N_13864,N_13714,N_13758);
or U13865 (N_13865,N_13656,N_13602);
and U13866 (N_13866,N_13743,N_13630);
nor U13867 (N_13867,N_13788,N_13645);
xnor U13868 (N_13868,N_13702,N_13746);
or U13869 (N_13869,N_13724,N_13783);
nand U13870 (N_13870,N_13678,N_13721);
or U13871 (N_13871,N_13730,N_13626);
and U13872 (N_13872,N_13638,N_13680);
xnor U13873 (N_13873,N_13727,N_13774);
and U13874 (N_13874,N_13722,N_13718);
or U13875 (N_13875,N_13639,N_13603);
nor U13876 (N_13876,N_13644,N_13782);
and U13877 (N_13877,N_13617,N_13634);
xor U13878 (N_13878,N_13778,N_13686);
nand U13879 (N_13879,N_13600,N_13670);
or U13880 (N_13880,N_13781,N_13754);
nand U13881 (N_13881,N_13614,N_13679);
nor U13882 (N_13882,N_13648,N_13687);
or U13883 (N_13883,N_13601,N_13725);
and U13884 (N_13884,N_13700,N_13647);
nand U13885 (N_13885,N_13708,N_13793);
nor U13886 (N_13886,N_13747,N_13740);
and U13887 (N_13887,N_13623,N_13659);
nand U13888 (N_13888,N_13798,N_13787);
nand U13889 (N_13889,N_13760,N_13713);
nor U13890 (N_13890,N_13769,N_13685);
xnor U13891 (N_13891,N_13651,N_13763);
or U13892 (N_13892,N_13655,N_13637);
or U13893 (N_13893,N_13759,N_13771);
nand U13894 (N_13894,N_13636,N_13707);
nor U13895 (N_13895,N_13731,N_13752);
nand U13896 (N_13896,N_13653,N_13618);
and U13897 (N_13897,N_13785,N_13791);
and U13898 (N_13898,N_13701,N_13610);
or U13899 (N_13899,N_13607,N_13664);
nor U13900 (N_13900,N_13674,N_13743);
and U13901 (N_13901,N_13747,N_13663);
or U13902 (N_13902,N_13670,N_13784);
and U13903 (N_13903,N_13607,N_13622);
or U13904 (N_13904,N_13609,N_13707);
nand U13905 (N_13905,N_13778,N_13741);
and U13906 (N_13906,N_13713,N_13740);
nand U13907 (N_13907,N_13755,N_13730);
or U13908 (N_13908,N_13783,N_13658);
nor U13909 (N_13909,N_13694,N_13693);
and U13910 (N_13910,N_13639,N_13677);
and U13911 (N_13911,N_13619,N_13684);
and U13912 (N_13912,N_13692,N_13667);
and U13913 (N_13913,N_13774,N_13611);
xor U13914 (N_13914,N_13774,N_13778);
xnor U13915 (N_13915,N_13607,N_13763);
or U13916 (N_13916,N_13712,N_13752);
and U13917 (N_13917,N_13681,N_13775);
and U13918 (N_13918,N_13783,N_13741);
xor U13919 (N_13919,N_13738,N_13652);
nor U13920 (N_13920,N_13626,N_13672);
xor U13921 (N_13921,N_13639,N_13610);
or U13922 (N_13922,N_13777,N_13746);
nand U13923 (N_13923,N_13609,N_13647);
nand U13924 (N_13924,N_13688,N_13714);
or U13925 (N_13925,N_13758,N_13604);
or U13926 (N_13926,N_13761,N_13773);
and U13927 (N_13927,N_13694,N_13795);
and U13928 (N_13928,N_13706,N_13778);
nor U13929 (N_13929,N_13772,N_13650);
nand U13930 (N_13930,N_13617,N_13685);
xor U13931 (N_13931,N_13693,N_13760);
nand U13932 (N_13932,N_13674,N_13609);
or U13933 (N_13933,N_13772,N_13625);
or U13934 (N_13934,N_13679,N_13611);
xnor U13935 (N_13935,N_13764,N_13634);
nand U13936 (N_13936,N_13676,N_13698);
or U13937 (N_13937,N_13695,N_13792);
nand U13938 (N_13938,N_13621,N_13702);
xor U13939 (N_13939,N_13778,N_13609);
or U13940 (N_13940,N_13677,N_13641);
or U13941 (N_13941,N_13618,N_13623);
or U13942 (N_13942,N_13777,N_13751);
xor U13943 (N_13943,N_13618,N_13685);
or U13944 (N_13944,N_13711,N_13707);
nand U13945 (N_13945,N_13663,N_13745);
and U13946 (N_13946,N_13641,N_13780);
or U13947 (N_13947,N_13745,N_13610);
or U13948 (N_13948,N_13758,N_13713);
and U13949 (N_13949,N_13761,N_13727);
and U13950 (N_13950,N_13694,N_13766);
xnor U13951 (N_13951,N_13743,N_13702);
and U13952 (N_13952,N_13604,N_13630);
nor U13953 (N_13953,N_13750,N_13704);
nand U13954 (N_13954,N_13649,N_13761);
xnor U13955 (N_13955,N_13609,N_13689);
and U13956 (N_13956,N_13645,N_13674);
nand U13957 (N_13957,N_13703,N_13693);
xnor U13958 (N_13958,N_13719,N_13619);
nor U13959 (N_13959,N_13794,N_13683);
and U13960 (N_13960,N_13718,N_13744);
nor U13961 (N_13961,N_13738,N_13784);
xor U13962 (N_13962,N_13713,N_13685);
xor U13963 (N_13963,N_13667,N_13799);
nand U13964 (N_13964,N_13798,N_13797);
nand U13965 (N_13965,N_13692,N_13659);
nor U13966 (N_13966,N_13794,N_13651);
nor U13967 (N_13967,N_13637,N_13796);
xnor U13968 (N_13968,N_13633,N_13693);
xor U13969 (N_13969,N_13657,N_13764);
nor U13970 (N_13970,N_13631,N_13756);
and U13971 (N_13971,N_13713,N_13723);
or U13972 (N_13972,N_13719,N_13745);
xnor U13973 (N_13973,N_13754,N_13656);
nor U13974 (N_13974,N_13747,N_13760);
xor U13975 (N_13975,N_13657,N_13625);
or U13976 (N_13976,N_13675,N_13695);
nand U13977 (N_13977,N_13614,N_13735);
or U13978 (N_13978,N_13746,N_13622);
nand U13979 (N_13979,N_13618,N_13758);
xnor U13980 (N_13980,N_13798,N_13663);
or U13981 (N_13981,N_13627,N_13750);
nand U13982 (N_13982,N_13751,N_13613);
xor U13983 (N_13983,N_13778,N_13757);
and U13984 (N_13984,N_13643,N_13625);
or U13985 (N_13985,N_13761,N_13651);
xnor U13986 (N_13986,N_13649,N_13646);
xor U13987 (N_13987,N_13656,N_13732);
and U13988 (N_13988,N_13777,N_13680);
xor U13989 (N_13989,N_13698,N_13613);
nor U13990 (N_13990,N_13720,N_13692);
or U13991 (N_13991,N_13793,N_13628);
or U13992 (N_13992,N_13645,N_13619);
and U13993 (N_13993,N_13759,N_13765);
or U13994 (N_13994,N_13697,N_13630);
nor U13995 (N_13995,N_13727,N_13729);
and U13996 (N_13996,N_13638,N_13747);
and U13997 (N_13997,N_13730,N_13657);
nor U13998 (N_13998,N_13675,N_13752);
nor U13999 (N_13999,N_13641,N_13668);
nor U14000 (N_14000,N_13831,N_13919);
nor U14001 (N_14001,N_13838,N_13858);
nor U14002 (N_14002,N_13917,N_13886);
and U14003 (N_14003,N_13980,N_13907);
or U14004 (N_14004,N_13813,N_13811);
or U14005 (N_14005,N_13990,N_13939);
nand U14006 (N_14006,N_13969,N_13952);
xor U14007 (N_14007,N_13946,N_13815);
nor U14008 (N_14008,N_13947,N_13844);
nand U14009 (N_14009,N_13982,N_13817);
or U14010 (N_14010,N_13897,N_13809);
and U14011 (N_14011,N_13934,N_13900);
nor U14012 (N_14012,N_13810,N_13859);
xor U14013 (N_14013,N_13891,N_13972);
nor U14014 (N_14014,N_13940,N_13856);
xnor U14015 (N_14015,N_13819,N_13832);
nor U14016 (N_14016,N_13883,N_13868);
nor U14017 (N_14017,N_13916,N_13818);
and U14018 (N_14018,N_13910,N_13887);
nand U14019 (N_14019,N_13943,N_13894);
nor U14020 (N_14020,N_13816,N_13884);
or U14021 (N_14021,N_13889,N_13824);
or U14022 (N_14022,N_13927,N_13906);
xnor U14023 (N_14023,N_13834,N_13997);
nor U14024 (N_14024,N_13950,N_13803);
nor U14025 (N_14025,N_13800,N_13911);
and U14026 (N_14026,N_13971,N_13964);
nor U14027 (N_14027,N_13960,N_13843);
xnor U14028 (N_14028,N_13975,N_13874);
or U14029 (N_14029,N_13877,N_13853);
xor U14030 (N_14030,N_13862,N_13961);
and U14031 (N_14031,N_13954,N_13935);
xor U14032 (N_14032,N_13867,N_13991);
nor U14033 (N_14033,N_13904,N_13846);
nand U14034 (N_14034,N_13914,N_13881);
xnor U14035 (N_14035,N_13888,N_13852);
xor U14036 (N_14036,N_13979,N_13849);
nor U14037 (N_14037,N_13976,N_13989);
nand U14038 (N_14038,N_13802,N_13829);
and U14039 (N_14039,N_13841,N_13922);
nand U14040 (N_14040,N_13977,N_13835);
nor U14041 (N_14041,N_13915,N_13928);
nand U14042 (N_14042,N_13845,N_13833);
and U14043 (N_14043,N_13872,N_13828);
nor U14044 (N_14044,N_13854,N_13936);
xnor U14045 (N_14045,N_13903,N_13873);
xnor U14046 (N_14046,N_13806,N_13981);
nand U14047 (N_14047,N_13973,N_13805);
and U14048 (N_14048,N_13901,N_13925);
xnor U14049 (N_14049,N_13959,N_13893);
nand U14050 (N_14050,N_13974,N_13863);
nand U14051 (N_14051,N_13808,N_13836);
and U14052 (N_14052,N_13822,N_13878);
nor U14053 (N_14053,N_13942,N_13801);
xor U14054 (N_14054,N_13966,N_13908);
nor U14055 (N_14055,N_13992,N_13984);
and U14056 (N_14056,N_13957,N_13968);
nand U14057 (N_14057,N_13861,N_13865);
xnor U14058 (N_14058,N_13931,N_13876);
nor U14059 (N_14059,N_13820,N_13932);
nand U14060 (N_14060,N_13965,N_13839);
xor U14061 (N_14061,N_13967,N_13804);
and U14062 (N_14062,N_13999,N_13921);
nor U14063 (N_14063,N_13912,N_13909);
xnor U14064 (N_14064,N_13913,N_13923);
or U14065 (N_14065,N_13827,N_13821);
nor U14066 (N_14066,N_13869,N_13945);
xor U14067 (N_14067,N_13937,N_13896);
xnor U14068 (N_14068,N_13892,N_13951);
nand U14069 (N_14069,N_13875,N_13895);
or U14070 (N_14070,N_13864,N_13956);
or U14071 (N_14071,N_13985,N_13963);
nand U14072 (N_14072,N_13993,N_13851);
nand U14073 (N_14073,N_13899,N_13949);
nor U14074 (N_14074,N_13823,N_13944);
nor U14075 (N_14075,N_13826,N_13924);
or U14076 (N_14076,N_13890,N_13983);
xnor U14077 (N_14077,N_13918,N_13830);
nand U14078 (N_14078,N_13812,N_13840);
or U14079 (N_14079,N_13933,N_13842);
and U14080 (N_14080,N_13955,N_13871);
xor U14081 (N_14081,N_13948,N_13807);
nand U14082 (N_14082,N_13995,N_13885);
nand U14083 (N_14083,N_13880,N_13970);
or U14084 (N_14084,N_13958,N_13837);
xor U14085 (N_14085,N_13902,N_13905);
and U14086 (N_14086,N_13941,N_13847);
and U14087 (N_14087,N_13962,N_13994);
and U14088 (N_14088,N_13988,N_13920);
or U14089 (N_14089,N_13882,N_13879);
nand U14090 (N_14090,N_13898,N_13857);
and U14091 (N_14091,N_13926,N_13870);
nand U14092 (N_14092,N_13866,N_13998);
nor U14093 (N_14093,N_13987,N_13986);
or U14094 (N_14094,N_13978,N_13953);
or U14095 (N_14095,N_13848,N_13855);
and U14096 (N_14096,N_13860,N_13930);
or U14097 (N_14097,N_13929,N_13850);
xnor U14098 (N_14098,N_13996,N_13825);
xor U14099 (N_14099,N_13938,N_13814);
nor U14100 (N_14100,N_13866,N_13871);
or U14101 (N_14101,N_13905,N_13901);
or U14102 (N_14102,N_13801,N_13946);
or U14103 (N_14103,N_13863,N_13996);
nor U14104 (N_14104,N_13908,N_13840);
xnor U14105 (N_14105,N_13989,N_13826);
nand U14106 (N_14106,N_13976,N_13864);
nor U14107 (N_14107,N_13966,N_13951);
and U14108 (N_14108,N_13824,N_13983);
xnor U14109 (N_14109,N_13811,N_13841);
xnor U14110 (N_14110,N_13822,N_13970);
nor U14111 (N_14111,N_13976,N_13954);
xnor U14112 (N_14112,N_13940,N_13964);
nand U14113 (N_14113,N_13927,N_13913);
or U14114 (N_14114,N_13820,N_13968);
or U14115 (N_14115,N_13988,N_13838);
and U14116 (N_14116,N_13835,N_13957);
nor U14117 (N_14117,N_13835,N_13935);
nor U14118 (N_14118,N_13801,N_13852);
nor U14119 (N_14119,N_13828,N_13860);
nand U14120 (N_14120,N_13924,N_13921);
nor U14121 (N_14121,N_13811,N_13964);
or U14122 (N_14122,N_13899,N_13871);
xor U14123 (N_14123,N_13991,N_13987);
xnor U14124 (N_14124,N_13866,N_13816);
xnor U14125 (N_14125,N_13925,N_13801);
nand U14126 (N_14126,N_13936,N_13980);
and U14127 (N_14127,N_13982,N_13825);
and U14128 (N_14128,N_13904,N_13815);
and U14129 (N_14129,N_13875,N_13996);
nor U14130 (N_14130,N_13916,N_13844);
nor U14131 (N_14131,N_13833,N_13927);
xor U14132 (N_14132,N_13984,N_13965);
and U14133 (N_14133,N_13972,N_13994);
and U14134 (N_14134,N_13857,N_13854);
nand U14135 (N_14135,N_13804,N_13944);
xnor U14136 (N_14136,N_13946,N_13968);
nor U14137 (N_14137,N_13865,N_13979);
nand U14138 (N_14138,N_13993,N_13873);
nand U14139 (N_14139,N_13810,N_13989);
nor U14140 (N_14140,N_13896,N_13849);
xor U14141 (N_14141,N_13967,N_13801);
and U14142 (N_14142,N_13963,N_13982);
or U14143 (N_14143,N_13972,N_13883);
xnor U14144 (N_14144,N_13883,N_13953);
or U14145 (N_14145,N_13934,N_13814);
nor U14146 (N_14146,N_13972,N_13818);
xnor U14147 (N_14147,N_13890,N_13955);
or U14148 (N_14148,N_13855,N_13835);
nor U14149 (N_14149,N_13899,N_13900);
nand U14150 (N_14150,N_13955,N_13997);
nor U14151 (N_14151,N_13873,N_13802);
nand U14152 (N_14152,N_13861,N_13949);
nor U14153 (N_14153,N_13838,N_13804);
or U14154 (N_14154,N_13906,N_13875);
xnor U14155 (N_14155,N_13998,N_13841);
xnor U14156 (N_14156,N_13936,N_13844);
nor U14157 (N_14157,N_13849,N_13917);
nor U14158 (N_14158,N_13845,N_13971);
xor U14159 (N_14159,N_13861,N_13822);
nor U14160 (N_14160,N_13818,N_13969);
or U14161 (N_14161,N_13839,N_13858);
nand U14162 (N_14162,N_13936,N_13925);
and U14163 (N_14163,N_13827,N_13950);
xor U14164 (N_14164,N_13977,N_13828);
nor U14165 (N_14165,N_13848,N_13861);
xor U14166 (N_14166,N_13828,N_13859);
xnor U14167 (N_14167,N_13807,N_13990);
nand U14168 (N_14168,N_13924,N_13815);
or U14169 (N_14169,N_13811,N_13925);
nor U14170 (N_14170,N_13929,N_13895);
nand U14171 (N_14171,N_13831,N_13939);
xor U14172 (N_14172,N_13836,N_13917);
nor U14173 (N_14173,N_13980,N_13844);
or U14174 (N_14174,N_13965,N_13841);
and U14175 (N_14175,N_13869,N_13854);
xor U14176 (N_14176,N_13982,N_13849);
nand U14177 (N_14177,N_13824,N_13806);
nand U14178 (N_14178,N_13939,N_13855);
nand U14179 (N_14179,N_13847,N_13961);
nand U14180 (N_14180,N_13949,N_13902);
and U14181 (N_14181,N_13829,N_13887);
nand U14182 (N_14182,N_13886,N_13814);
and U14183 (N_14183,N_13846,N_13990);
xor U14184 (N_14184,N_13879,N_13820);
or U14185 (N_14185,N_13897,N_13896);
nand U14186 (N_14186,N_13894,N_13848);
and U14187 (N_14187,N_13852,N_13857);
nand U14188 (N_14188,N_13804,N_13991);
nand U14189 (N_14189,N_13881,N_13967);
xnor U14190 (N_14190,N_13964,N_13852);
xor U14191 (N_14191,N_13934,N_13811);
nor U14192 (N_14192,N_13964,N_13982);
nor U14193 (N_14193,N_13978,N_13936);
xor U14194 (N_14194,N_13804,N_13883);
nand U14195 (N_14195,N_13983,N_13822);
nand U14196 (N_14196,N_13988,N_13824);
nor U14197 (N_14197,N_13991,N_13915);
xnor U14198 (N_14198,N_13868,N_13984);
nand U14199 (N_14199,N_13954,N_13939);
and U14200 (N_14200,N_14013,N_14170);
or U14201 (N_14201,N_14183,N_14017);
nand U14202 (N_14202,N_14055,N_14035);
and U14203 (N_14203,N_14159,N_14168);
nand U14204 (N_14204,N_14020,N_14145);
and U14205 (N_14205,N_14027,N_14021);
xor U14206 (N_14206,N_14056,N_14063);
nand U14207 (N_14207,N_14028,N_14005);
nor U14208 (N_14208,N_14113,N_14196);
xor U14209 (N_14209,N_14184,N_14048);
and U14210 (N_14210,N_14133,N_14120);
nand U14211 (N_14211,N_14084,N_14167);
or U14212 (N_14212,N_14111,N_14066);
nor U14213 (N_14213,N_14092,N_14047);
and U14214 (N_14214,N_14004,N_14000);
xnor U14215 (N_14215,N_14036,N_14138);
nor U14216 (N_14216,N_14097,N_14175);
nor U14217 (N_14217,N_14131,N_14107);
nand U14218 (N_14218,N_14153,N_14038);
nand U14219 (N_14219,N_14192,N_14102);
xnor U14220 (N_14220,N_14143,N_14094);
and U14221 (N_14221,N_14037,N_14018);
nor U14222 (N_14222,N_14051,N_14144);
nor U14223 (N_14223,N_14098,N_14079);
xnor U14224 (N_14224,N_14198,N_14095);
nor U14225 (N_14225,N_14029,N_14067);
and U14226 (N_14226,N_14002,N_14185);
nor U14227 (N_14227,N_14059,N_14060);
and U14228 (N_14228,N_14009,N_14032);
and U14229 (N_14229,N_14135,N_14134);
or U14230 (N_14230,N_14065,N_14186);
and U14231 (N_14231,N_14165,N_14034);
and U14232 (N_14232,N_14177,N_14171);
xnor U14233 (N_14233,N_14157,N_14085);
nand U14234 (N_14234,N_14052,N_14054);
nand U14235 (N_14235,N_14126,N_14069);
and U14236 (N_14236,N_14078,N_14103);
nand U14237 (N_14237,N_14108,N_14033);
and U14238 (N_14238,N_14129,N_14043);
or U14239 (N_14239,N_14161,N_14166);
nor U14240 (N_14240,N_14091,N_14190);
nand U14241 (N_14241,N_14125,N_14011);
xor U14242 (N_14242,N_14119,N_14044);
nand U14243 (N_14243,N_14016,N_14140);
and U14244 (N_14244,N_14096,N_14172);
xnor U14245 (N_14245,N_14109,N_14188);
nor U14246 (N_14246,N_14176,N_14040);
xnor U14247 (N_14247,N_14019,N_14100);
xnor U14248 (N_14248,N_14124,N_14008);
and U14249 (N_14249,N_14083,N_14174);
and U14250 (N_14250,N_14121,N_14158);
and U14251 (N_14251,N_14187,N_14156);
nor U14252 (N_14252,N_14023,N_14073);
nor U14253 (N_14253,N_14071,N_14075);
and U14254 (N_14254,N_14058,N_14042);
or U14255 (N_14255,N_14025,N_14147);
and U14256 (N_14256,N_14137,N_14064);
and U14257 (N_14257,N_14076,N_14101);
xnor U14258 (N_14258,N_14041,N_14199);
or U14259 (N_14259,N_14169,N_14142);
and U14260 (N_14260,N_14088,N_14081);
or U14261 (N_14261,N_14118,N_14045);
nor U14262 (N_14262,N_14050,N_14164);
xor U14263 (N_14263,N_14180,N_14001);
nand U14264 (N_14264,N_14082,N_14115);
nand U14265 (N_14265,N_14105,N_14114);
nand U14266 (N_14266,N_14136,N_14179);
nor U14267 (N_14267,N_14139,N_14122);
and U14268 (N_14268,N_14012,N_14022);
or U14269 (N_14269,N_14062,N_14099);
xnor U14270 (N_14270,N_14003,N_14049);
xor U14271 (N_14271,N_14080,N_14104);
and U14272 (N_14272,N_14072,N_14191);
nand U14273 (N_14273,N_14024,N_14155);
and U14274 (N_14274,N_14146,N_14106);
and U14275 (N_14275,N_14128,N_14141);
or U14276 (N_14276,N_14015,N_14031);
xor U14277 (N_14277,N_14007,N_14160);
and U14278 (N_14278,N_14026,N_14061);
xnor U14279 (N_14279,N_14194,N_14182);
or U14280 (N_14280,N_14077,N_14086);
and U14281 (N_14281,N_14162,N_14068);
nand U14282 (N_14282,N_14014,N_14087);
nand U14283 (N_14283,N_14112,N_14150);
xnor U14284 (N_14284,N_14148,N_14181);
or U14285 (N_14285,N_14053,N_14030);
nand U14286 (N_14286,N_14116,N_14197);
or U14287 (N_14287,N_14110,N_14057);
xor U14288 (N_14288,N_14127,N_14152);
and U14289 (N_14289,N_14090,N_14151);
nand U14290 (N_14290,N_14010,N_14189);
nand U14291 (N_14291,N_14074,N_14070);
nand U14292 (N_14292,N_14154,N_14132);
or U14293 (N_14293,N_14178,N_14130);
xnor U14294 (N_14294,N_14089,N_14117);
nor U14295 (N_14295,N_14123,N_14195);
or U14296 (N_14296,N_14173,N_14193);
and U14297 (N_14297,N_14046,N_14039);
xor U14298 (N_14298,N_14149,N_14093);
or U14299 (N_14299,N_14163,N_14006);
nand U14300 (N_14300,N_14011,N_14157);
and U14301 (N_14301,N_14173,N_14019);
nand U14302 (N_14302,N_14137,N_14126);
nand U14303 (N_14303,N_14093,N_14069);
nor U14304 (N_14304,N_14144,N_14088);
nand U14305 (N_14305,N_14007,N_14194);
and U14306 (N_14306,N_14080,N_14158);
nor U14307 (N_14307,N_14045,N_14029);
nand U14308 (N_14308,N_14047,N_14043);
and U14309 (N_14309,N_14107,N_14125);
xnor U14310 (N_14310,N_14010,N_14005);
or U14311 (N_14311,N_14059,N_14075);
nand U14312 (N_14312,N_14094,N_14166);
xor U14313 (N_14313,N_14093,N_14132);
xnor U14314 (N_14314,N_14191,N_14042);
and U14315 (N_14315,N_14180,N_14052);
and U14316 (N_14316,N_14121,N_14148);
or U14317 (N_14317,N_14129,N_14016);
xor U14318 (N_14318,N_14118,N_14040);
or U14319 (N_14319,N_14014,N_14175);
nand U14320 (N_14320,N_14152,N_14051);
and U14321 (N_14321,N_14120,N_14094);
nand U14322 (N_14322,N_14070,N_14187);
nor U14323 (N_14323,N_14133,N_14043);
or U14324 (N_14324,N_14161,N_14095);
and U14325 (N_14325,N_14111,N_14022);
or U14326 (N_14326,N_14138,N_14109);
nor U14327 (N_14327,N_14050,N_14175);
nor U14328 (N_14328,N_14011,N_14117);
nor U14329 (N_14329,N_14093,N_14184);
or U14330 (N_14330,N_14181,N_14021);
nor U14331 (N_14331,N_14108,N_14073);
nand U14332 (N_14332,N_14023,N_14170);
and U14333 (N_14333,N_14057,N_14052);
or U14334 (N_14334,N_14054,N_14026);
nand U14335 (N_14335,N_14079,N_14119);
nor U14336 (N_14336,N_14194,N_14141);
xor U14337 (N_14337,N_14095,N_14185);
nor U14338 (N_14338,N_14065,N_14067);
and U14339 (N_14339,N_14053,N_14103);
nor U14340 (N_14340,N_14130,N_14105);
xnor U14341 (N_14341,N_14192,N_14014);
xnor U14342 (N_14342,N_14156,N_14140);
xnor U14343 (N_14343,N_14135,N_14153);
or U14344 (N_14344,N_14174,N_14002);
and U14345 (N_14345,N_14079,N_14040);
nor U14346 (N_14346,N_14088,N_14082);
nand U14347 (N_14347,N_14127,N_14131);
or U14348 (N_14348,N_14157,N_14112);
nor U14349 (N_14349,N_14123,N_14095);
or U14350 (N_14350,N_14105,N_14132);
or U14351 (N_14351,N_14189,N_14153);
or U14352 (N_14352,N_14101,N_14159);
xor U14353 (N_14353,N_14054,N_14160);
and U14354 (N_14354,N_14121,N_14124);
xnor U14355 (N_14355,N_14136,N_14073);
and U14356 (N_14356,N_14061,N_14054);
nand U14357 (N_14357,N_14190,N_14090);
nor U14358 (N_14358,N_14140,N_14065);
and U14359 (N_14359,N_14152,N_14194);
nor U14360 (N_14360,N_14127,N_14132);
nand U14361 (N_14361,N_14054,N_14014);
nor U14362 (N_14362,N_14077,N_14083);
nor U14363 (N_14363,N_14172,N_14001);
nand U14364 (N_14364,N_14043,N_14164);
nand U14365 (N_14365,N_14195,N_14172);
nor U14366 (N_14366,N_14058,N_14049);
nor U14367 (N_14367,N_14054,N_14008);
xor U14368 (N_14368,N_14009,N_14067);
xor U14369 (N_14369,N_14183,N_14149);
nand U14370 (N_14370,N_14129,N_14173);
nand U14371 (N_14371,N_14137,N_14059);
and U14372 (N_14372,N_14072,N_14097);
and U14373 (N_14373,N_14183,N_14143);
nor U14374 (N_14374,N_14172,N_14187);
nand U14375 (N_14375,N_14068,N_14073);
or U14376 (N_14376,N_14152,N_14101);
nand U14377 (N_14377,N_14091,N_14166);
nand U14378 (N_14378,N_14016,N_14010);
xnor U14379 (N_14379,N_14195,N_14107);
xnor U14380 (N_14380,N_14173,N_14045);
xnor U14381 (N_14381,N_14062,N_14179);
xnor U14382 (N_14382,N_14166,N_14008);
and U14383 (N_14383,N_14075,N_14112);
or U14384 (N_14384,N_14157,N_14174);
nor U14385 (N_14385,N_14093,N_14084);
xor U14386 (N_14386,N_14153,N_14118);
nor U14387 (N_14387,N_14085,N_14017);
and U14388 (N_14388,N_14042,N_14044);
and U14389 (N_14389,N_14003,N_14110);
xnor U14390 (N_14390,N_14095,N_14155);
nor U14391 (N_14391,N_14150,N_14059);
or U14392 (N_14392,N_14142,N_14023);
nor U14393 (N_14393,N_14054,N_14007);
and U14394 (N_14394,N_14038,N_14030);
xor U14395 (N_14395,N_14166,N_14099);
nor U14396 (N_14396,N_14156,N_14020);
xor U14397 (N_14397,N_14020,N_14106);
or U14398 (N_14398,N_14042,N_14080);
nand U14399 (N_14399,N_14181,N_14156);
and U14400 (N_14400,N_14398,N_14238);
nor U14401 (N_14401,N_14249,N_14384);
or U14402 (N_14402,N_14336,N_14232);
xor U14403 (N_14403,N_14389,N_14221);
nor U14404 (N_14404,N_14280,N_14343);
nand U14405 (N_14405,N_14335,N_14369);
nand U14406 (N_14406,N_14345,N_14203);
nand U14407 (N_14407,N_14394,N_14278);
and U14408 (N_14408,N_14388,N_14275);
and U14409 (N_14409,N_14269,N_14287);
xor U14410 (N_14410,N_14285,N_14252);
nor U14411 (N_14411,N_14248,N_14344);
xnor U14412 (N_14412,N_14319,N_14245);
and U14413 (N_14413,N_14205,N_14339);
nor U14414 (N_14414,N_14274,N_14347);
nand U14415 (N_14415,N_14380,N_14243);
and U14416 (N_14416,N_14210,N_14362);
and U14417 (N_14417,N_14244,N_14211);
nand U14418 (N_14418,N_14301,N_14229);
nand U14419 (N_14419,N_14355,N_14333);
nor U14420 (N_14420,N_14202,N_14324);
nor U14421 (N_14421,N_14207,N_14391);
or U14422 (N_14422,N_14363,N_14304);
or U14423 (N_14423,N_14354,N_14250);
nand U14424 (N_14424,N_14268,N_14214);
nor U14425 (N_14425,N_14235,N_14292);
or U14426 (N_14426,N_14382,N_14390);
nand U14427 (N_14427,N_14370,N_14314);
or U14428 (N_14428,N_14360,N_14321);
and U14429 (N_14429,N_14367,N_14399);
or U14430 (N_14430,N_14374,N_14266);
or U14431 (N_14431,N_14209,N_14378);
nor U14432 (N_14432,N_14247,N_14239);
and U14433 (N_14433,N_14386,N_14272);
or U14434 (N_14434,N_14200,N_14340);
nor U14435 (N_14435,N_14261,N_14297);
or U14436 (N_14436,N_14387,N_14338);
or U14437 (N_14437,N_14326,N_14392);
and U14438 (N_14438,N_14204,N_14227);
and U14439 (N_14439,N_14226,N_14309);
or U14440 (N_14440,N_14311,N_14352);
and U14441 (N_14441,N_14322,N_14222);
nand U14442 (N_14442,N_14383,N_14315);
nor U14443 (N_14443,N_14234,N_14351);
and U14444 (N_14444,N_14323,N_14296);
xor U14445 (N_14445,N_14299,N_14356);
nor U14446 (N_14446,N_14317,N_14371);
nand U14447 (N_14447,N_14341,N_14373);
nand U14448 (N_14448,N_14242,N_14290);
xor U14449 (N_14449,N_14320,N_14377);
or U14450 (N_14450,N_14372,N_14375);
nor U14451 (N_14451,N_14307,N_14313);
xor U14452 (N_14452,N_14286,N_14328);
and U14453 (N_14453,N_14293,N_14251);
and U14454 (N_14454,N_14306,N_14316);
or U14455 (N_14455,N_14302,N_14225);
or U14456 (N_14456,N_14218,N_14288);
nand U14457 (N_14457,N_14330,N_14279);
xor U14458 (N_14458,N_14258,N_14318);
or U14459 (N_14459,N_14254,N_14361);
xor U14460 (N_14460,N_14310,N_14271);
xor U14461 (N_14461,N_14282,N_14350);
nor U14462 (N_14462,N_14349,N_14256);
or U14463 (N_14463,N_14253,N_14327);
nor U14464 (N_14464,N_14283,N_14300);
and U14465 (N_14465,N_14368,N_14237);
nand U14466 (N_14466,N_14212,N_14263);
or U14467 (N_14467,N_14359,N_14284);
and U14468 (N_14468,N_14267,N_14334);
xnor U14469 (N_14469,N_14376,N_14303);
nor U14470 (N_14470,N_14312,N_14381);
nand U14471 (N_14471,N_14223,N_14230);
and U14472 (N_14472,N_14281,N_14255);
nand U14473 (N_14473,N_14291,N_14206);
nand U14474 (N_14474,N_14379,N_14216);
xor U14475 (N_14475,N_14366,N_14397);
nand U14476 (N_14476,N_14260,N_14241);
and U14477 (N_14477,N_14217,N_14357);
nand U14478 (N_14478,N_14273,N_14201);
and U14479 (N_14479,N_14358,N_14213);
or U14480 (N_14480,N_14215,N_14331);
xnor U14481 (N_14481,N_14220,N_14294);
and U14482 (N_14482,N_14264,N_14329);
nor U14483 (N_14483,N_14295,N_14393);
or U14484 (N_14484,N_14348,N_14240);
xor U14485 (N_14485,N_14395,N_14236);
and U14486 (N_14486,N_14298,N_14224);
and U14487 (N_14487,N_14308,N_14259);
or U14488 (N_14488,N_14228,N_14231);
and U14489 (N_14489,N_14305,N_14353);
and U14490 (N_14490,N_14332,N_14364);
nor U14491 (N_14491,N_14277,N_14219);
xnor U14492 (N_14492,N_14276,N_14346);
nor U14493 (N_14493,N_14337,N_14246);
xnor U14494 (N_14494,N_14262,N_14208);
and U14495 (N_14495,N_14365,N_14385);
and U14496 (N_14496,N_14289,N_14233);
and U14497 (N_14497,N_14396,N_14257);
xor U14498 (N_14498,N_14265,N_14325);
or U14499 (N_14499,N_14270,N_14342);
and U14500 (N_14500,N_14349,N_14264);
and U14501 (N_14501,N_14294,N_14279);
xnor U14502 (N_14502,N_14379,N_14291);
and U14503 (N_14503,N_14215,N_14288);
nand U14504 (N_14504,N_14282,N_14352);
nor U14505 (N_14505,N_14397,N_14377);
and U14506 (N_14506,N_14319,N_14373);
and U14507 (N_14507,N_14399,N_14200);
nand U14508 (N_14508,N_14375,N_14335);
xnor U14509 (N_14509,N_14369,N_14345);
xor U14510 (N_14510,N_14369,N_14259);
xor U14511 (N_14511,N_14200,N_14341);
and U14512 (N_14512,N_14388,N_14352);
xor U14513 (N_14513,N_14398,N_14302);
nand U14514 (N_14514,N_14289,N_14202);
xor U14515 (N_14515,N_14229,N_14308);
and U14516 (N_14516,N_14202,N_14208);
nand U14517 (N_14517,N_14339,N_14248);
and U14518 (N_14518,N_14301,N_14365);
or U14519 (N_14519,N_14233,N_14356);
nor U14520 (N_14520,N_14205,N_14346);
or U14521 (N_14521,N_14343,N_14203);
or U14522 (N_14522,N_14339,N_14329);
nand U14523 (N_14523,N_14261,N_14395);
nand U14524 (N_14524,N_14278,N_14272);
nor U14525 (N_14525,N_14335,N_14249);
xor U14526 (N_14526,N_14315,N_14201);
nor U14527 (N_14527,N_14275,N_14346);
or U14528 (N_14528,N_14234,N_14362);
or U14529 (N_14529,N_14218,N_14278);
nor U14530 (N_14530,N_14298,N_14374);
or U14531 (N_14531,N_14384,N_14301);
xnor U14532 (N_14532,N_14349,N_14359);
nor U14533 (N_14533,N_14388,N_14392);
xor U14534 (N_14534,N_14355,N_14291);
or U14535 (N_14535,N_14397,N_14350);
nand U14536 (N_14536,N_14226,N_14273);
xnor U14537 (N_14537,N_14348,N_14365);
nor U14538 (N_14538,N_14242,N_14219);
or U14539 (N_14539,N_14346,N_14396);
nor U14540 (N_14540,N_14209,N_14269);
xor U14541 (N_14541,N_14229,N_14281);
nor U14542 (N_14542,N_14277,N_14306);
nor U14543 (N_14543,N_14281,N_14283);
xnor U14544 (N_14544,N_14336,N_14297);
nand U14545 (N_14545,N_14225,N_14311);
and U14546 (N_14546,N_14322,N_14242);
or U14547 (N_14547,N_14274,N_14346);
and U14548 (N_14548,N_14345,N_14331);
nor U14549 (N_14549,N_14254,N_14387);
or U14550 (N_14550,N_14291,N_14223);
nand U14551 (N_14551,N_14294,N_14213);
and U14552 (N_14552,N_14395,N_14238);
and U14553 (N_14553,N_14202,N_14205);
nand U14554 (N_14554,N_14284,N_14220);
and U14555 (N_14555,N_14365,N_14346);
xnor U14556 (N_14556,N_14231,N_14395);
nand U14557 (N_14557,N_14338,N_14328);
and U14558 (N_14558,N_14248,N_14334);
or U14559 (N_14559,N_14246,N_14372);
and U14560 (N_14560,N_14356,N_14246);
nor U14561 (N_14561,N_14308,N_14340);
nor U14562 (N_14562,N_14357,N_14291);
or U14563 (N_14563,N_14210,N_14367);
nor U14564 (N_14564,N_14290,N_14211);
xnor U14565 (N_14565,N_14212,N_14276);
nor U14566 (N_14566,N_14329,N_14216);
nand U14567 (N_14567,N_14391,N_14282);
or U14568 (N_14568,N_14217,N_14263);
xnor U14569 (N_14569,N_14326,N_14228);
or U14570 (N_14570,N_14289,N_14321);
and U14571 (N_14571,N_14325,N_14226);
nor U14572 (N_14572,N_14281,N_14321);
xnor U14573 (N_14573,N_14327,N_14352);
xnor U14574 (N_14574,N_14255,N_14366);
or U14575 (N_14575,N_14320,N_14351);
xnor U14576 (N_14576,N_14384,N_14202);
nand U14577 (N_14577,N_14398,N_14290);
or U14578 (N_14578,N_14257,N_14306);
nand U14579 (N_14579,N_14351,N_14331);
xor U14580 (N_14580,N_14251,N_14207);
xnor U14581 (N_14581,N_14344,N_14327);
and U14582 (N_14582,N_14348,N_14302);
nor U14583 (N_14583,N_14254,N_14223);
and U14584 (N_14584,N_14396,N_14393);
xor U14585 (N_14585,N_14264,N_14353);
xor U14586 (N_14586,N_14274,N_14325);
or U14587 (N_14587,N_14367,N_14325);
and U14588 (N_14588,N_14307,N_14399);
xnor U14589 (N_14589,N_14362,N_14227);
nand U14590 (N_14590,N_14287,N_14319);
xnor U14591 (N_14591,N_14222,N_14373);
nor U14592 (N_14592,N_14207,N_14318);
nor U14593 (N_14593,N_14378,N_14225);
or U14594 (N_14594,N_14321,N_14237);
and U14595 (N_14595,N_14298,N_14371);
or U14596 (N_14596,N_14334,N_14359);
xor U14597 (N_14597,N_14272,N_14345);
and U14598 (N_14598,N_14248,N_14219);
nand U14599 (N_14599,N_14373,N_14265);
and U14600 (N_14600,N_14445,N_14403);
xor U14601 (N_14601,N_14569,N_14455);
and U14602 (N_14602,N_14593,N_14542);
or U14603 (N_14603,N_14410,N_14434);
nand U14604 (N_14604,N_14500,N_14591);
nor U14605 (N_14605,N_14432,N_14531);
nand U14606 (N_14606,N_14519,N_14448);
nor U14607 (N_14607,N_14541,N_14435);
or U14608 (N_14608,N_14442,N_14524);
nand U14609 (N_14609,N_14515,N_14518);
and U14610 (N_14610,N_14472,N_14585);
or U14611 (N_14611,N_14417,N_14439);
or U14612 (N_14612,N_14503,N_14488);
nor U14613 (N_14613,N_14550,N_14504);
nand U14614 (N_14614,N_14446,N_14592);
nor U14615 (N_14615,N_14582,N_14421);
xnor U14616 (N_14616,N_14482,N_14554);
xnor U14617 (N_14617,N_14574,N_14427);
nand U14618 (N_14618,N_14563,N_14538);
xnor U14619 (N_14619,N_14549,N_14493);
nor U14620 (N_14620,N_14419,N_14548);
or U14621 (N_14621,N_14426,N_14491);
or U14622 (N_14622,N_14573,N_14551);
or U14623 (N_14623,N_14539,N_14578);
nor U14624 (N_14624,N_14566,N_14570);
nand U14625 (N_14625,N_14490,N_14444);
or U14626 (N_14626,N_14559,N_14590);
and U14627 (N_14627,N_14537,N_14430);
and U14628 (N_14628,N_14479,N_14425);
or U14629 (N_14629,N_14599,N_14498);
or U14630 (N_14630,N_14489,N_14579);
nand U14631 (N_14631,N_14483,N_14407);
nand U14632 (N_14632,N_14527,N_14598);
xor U14633 (N_14633,N_14583,N_14495);
nand U14634 (N_14634,N_14438,N_14576);
or U14635 (N_14635,N_14433,N_14497);
xnor U14636 (N_14636,N_14440,N_14552);
nor U14637 (N_14637,N_14530,N_14521);
or U14638 (N_14638,N_14516,N_14466);
nand U14639 (N_14639,N_14454,N_14437);
nor U14640 (N_14640,N_14588,N_14581);
and U14641 (N_14641,N_14486,N_14547);
and U14642 (N_14642,N_14546,N_14406);
and U14643 (N_14643,N_14422,N_14414);
nand U14644 (N_14644,N_14464,N_14568);
or U14645 (N_14645,N_14544,N_14564);
or U14646 (N_14646,N_14533,N_14557);
xor U14647 (N_14647,N_14405,N_14526);
xnor U14648 (N_14648,N_14499,N_14441);
nand U14649 (N_14649,N_14453,N_14485);
nor U14650 (N_14650,N_14436,N_14484);
xor U14651 (N_14651,N_14477,N_14431);
nor U14652 (N_14652,N_14523,N_14561);
xnor U14653 (N_14653,N_14517,N_14451);
and U14654 (N_14654,N_14468,N_14412);
or U14655 (N_14655,N_14536,N_14589);
nor U14656 (N_14656,N_14528,N_14481);
xnor U14657 (N_14657,N_14507,N_14501);
or U14658 (N_14658,N_14467,N_14565);
nor U14659 (N_14659,N_14465,N_14404);
xnor U14660 (N_14660,N_14513,N_14562);
or U14661 (N_14661,N_14416,N_14461);
nand U14662 (N_14662,N_14543,N_14449);
or U14663 (N_14663,N_14408,N_14514);
xor U14664 (N_14664,N_14474,N_14476);
nand U14665 (N_14665,N_14558,N_14560);
or U14666 (N_14666,N_14460,N_14411);
nand U14667 (N_14667,N_14494,N_14597);
nand U14668 (N_14668,N_14525,N_14413);
and U14669 (N_14669,N_14458,N_14480);
and U14670 (N_14670,N_14402,N_14509);
or U14671 (N_14671,N_14492,N_14456);
nor U14672 (N_14672,N_14512,N_14545);
xor U14673 (N_14673,N_14534,N_14577);
nor U14674 (N_14674,N_14511,N_14556);
and U14675 (N_14675,N_14510,N_14478);
and U14676 (N_14676,N_14529,N_14409);
or U14677 (N_14677,N_14584,N_14400);
and U14678 (N_14678,N_14450,N_14487);
and U14679 (N_14679,N_14424,N_14575);
nand U14680 (N_14680,N_14555,N_14471);
nor U14681 (N_14681,N_14594,N_14580);
or U14682 (N_14682,N_14535,N_14506);
nand U14683 (N_14683,N_14447,N_14443);
nor U14684 (N_14684,N_14596,N_14572);
nand U14685 (N_14685,N_14553,N_14496);
xor U14686 (N_14686,N_14567,N_14420);
and U14687 (N_14687,N_14429,N_14571);
nand U14688 (N_14688,N_14502,N_14508);
nor U14689 (N_14689,N_14520,N_14463);
nand U14690 (N_14690,N_14505,N_14587);
nor U14691 (N_14691,N_14401,N_14532);
nor U14692 (N_14692,N_14586,N_14418);
nor U14693 (N_14693,N_14415,N_14473);
or U14694 (N_14694,N_14457,N_14462);
nand U14695 (N_14695,N_14540,N_14423);
nand U14696 (N_14696,N_14522,N_14428);
nor U14697 (N_14697,N_14452,N_14459);
nand U14698 (N_14698,N_14469,N_14595);
and U14699 (N_14699,N_14470,N_14475);
and U14700 (N_14700,N_14508,N_14443);
xor U14701 (N_14701,N_14556,N_14587);
or U14702 (N_14702,N_14527,N_14526);
or U14703 (N_14703,N_14407,N_14583);
nand U14704 (N_14704,N_14408,N_14422);
and U14705 (N_14705,N_14560,N_14547);
and U14706 (N_14706,N_14467,N_14546);
nand U14707 (N_14707,N_14543,N_14544);
nand U14708 (N_14708,N_14455,N_14540);
xor U14709 (N_14709,N_14445,N_14582);
xnor U14710 (N_14710,N_14416,N_14471);
nand U14711 (N_14711,N_14539,N_14551);
nand U14712 (N_14712,N_14456,N_14408);
and U14713 (N_14713,N_14403,N_14520);
nor U14714 (N_14714,N_14436,N_14594);
nor U14715 (N_14715,N_14544,N_14409);
or U14716 (N_14716,N_14445,N_14479);
nand U14717 (N_14717,N_14402,N_14412);
or U14718 (N_14718,N_14514,N_14419);
xor U14719 (N_14719,N_14430,N_14596);
nand U14720 (N_14720,N_14547,N_14419);
or U14721 (N_14721,N_14595,N_14459);
nor U14722 (N_14722,N_14497,N_14529);
nand U14723 (N_14723,N_14470,N_14455);
xor U14724 (N_14724,N_14492,N_14591);
xor U14725 (N_14725,N_14579,N_14481);
nor U14726 (N_14726,N_14468,N_14588);
nand U14727 (N_14727,N_14534,N_14471);
and U14728 (N_14728,N_14488,N_14534);
nand U14729 (N_14729,N_14585,N_14446);
nand U14730 (N_14730,N_14484,N_14551);
and U14731 (N_14731,N_14495,N_14556);
nor U14732 (N_14732,N_14549,N_14507);
xor U14733 (N_14733,N_14496,N_14544);
nand U14734 (N_14734,N_14415,N_14531);
xor U14735 (N_14735,N_14507,N_14590);
nand U14736 (N_14736,N_14566,N_14590);
nand U14737 (N_14737,N_14563,N_14421);
xnor U14738 (N_14738,N_14406,N_14503);
xnor U14739 (N_14739,N_14471,N_14539);
or U14740 (N_14740,N_14440,N_14578);
nor U14741 (N_14741,N_14429,N_14546);
nor U14742 (N_14742,N_14454,N_14426);
xnor U14743 (N_14743,N_14533,N_14543);
or U14744 (N_14744,N_14470,N_14558);
xor U14745 (N_14745,N_14527,N_14533);
nor U14746 (N_14746,N_14570,N_14437);
or U14747 (N_14747,N_14467,N_14460);
or U14748 (N_14748,N_14575,N_14516);
and U14749 (N_14749,N_14504,N_14581);
and U14750 (N_14750,N_14566,N_14578);
nor U14751 (N_14751,N_14417,N_14590);
xnor U14752 (N_14752,N_14527,N_14523);
nand U14753 (N_14753,N_14586,N_14507);
nand U14754 (N_14754,N_14569,N_14468);
nor U14755 (N_14755,N_14434,N_14541);
nor U14756 (N_14756,N_14598,N_14468);
and U14757 (N_14757,N_14503,N_14468);
or U14758 (N_14758,N_14449,N_14563);
xor U14759 (N_14759,N_14579,N_14567);
nor U14760 (N_14760,N_14419,N_14584);
and U14761 (N_14761,N_14499,N_14582);
nor U14762 (N_14762,N_14509,N_14544);
and U14763 (N_14763,N_14407,N_14481);
xnor U14764 (N_14764,N_14424,N_14510);
and U14765 (N_14765,N_14564,N_14494);
xnor U14766 (N_14766,N_14445,N_14599);
nand U14767 (N_14767,N_14453,N_14500);
or U14768 (N_14768,N_14489,N_14436);
xor U14769 (N_14769,N_14482,N_14479);
xnor U14770 (N_14770,N_14550,N_14493);
and U14771 (N_14771,N_14492,N_14407);
nand U14772 (N_14772,N_14554,N_14558);
nor U14773 (N_14773,N_14422,N_14465);
xor U14774 (N_14774,N_14545,N_14469);
and U14775 (N_14775,N_14475,N_14583);
nand U14776 (N_14776,N_14512,N_14412);
or U14777 (N_14777,N_14513,N_14535);
nor U14778 (N_14778,N_14429,N_14478);
or U14779 (N_14779,N_14476,N_14593);
or U14780 (N_14780,N_14483,N_14502);
or U14781 (N_14781,N_14522,N_14559);
and U14782 (N_14782,N_14436,N_14498);
nor U14783 (N_14783,N_14507,N_14444);
nor U14784 (N_14784,N_14598,N_14506);
nand U14785 (N_14785,N_14427,N_14552);
nand U14786 (N_14786,N_14553,N_14446);
xor U14787 (N_14787,N_14505,N_14547);
xor U14788 (N_14788,N_14488,N_14494);
or U14789 (N_14789,N_14437,N_14417);
or U14790 (N_14790,N_14431,N_14566);
nand U14791 (N_14791,N_14573,N_14488);
and U14792 (N_14792,N_14462,N_14561);
nand U14793 (N_14793,N_14502,N_14562);
nand U14794 (N_14794,N_14586,N_14466);
xnor U14795 (N_14795,N_14465,N_14492);
and U14796 (N_14796,N_14554,N_14524);
xor U14797 (N_14797,N_14425,N_14489);
xnor U14798 (N_14798,N_14401,N_14560);
xnor U14799 (N_14799,N_14593,N_14409);
nand U14800 (N_14800,N_14603,N_14651);
nand U14801 (N_14801,N_14797,N_14788);
or U14802 (N_14802,N_14778,N_14798);
and U14803 (N_14803,N_14764,N_14690);
nand U14804 (N_14804,N_14721,N_14691);
xnor U14805 (N_14805,N_14611,N_14645);
or U14806 (N_14806,N_14765,N_14633);
nand U14807 (N_14807,N_14720,N_14696);
and U14808 (N_14808,N_14644,N_14713);
nand U14809 (N_14809,N_14648,N_14607);
nand U14810 (N_14810,N_14716,N_14752);
or U14811 (N_14811,N_14799,N_14731);
nor U14812 (N_14812,N_14763,N_14640);
nor U14813 (N_14813,N_14717,N_14602);
nor U14814 (N_14814,N_14727,N_14733);
xnor U14815 (N_14815,N_14749,N_14624);
nor U14816 (N_14816,N_14695,N_14652);
nand U14817 (N_14817,N_14792,N_14747);
nor U14818 (N_14818,N_14739,N_14679);
xor U14819 (N_14819,N_14672,N_14693);
or U14820 (N_14820,N_14662,N_14785);
xor U14821 (N_14821,N_14671,N_14722);
xor U14822 (N_14822,N_14723,N_14639);
or U14823 (N_14823,N_14780,N_14726);
or U14824 (N_14824,N_14794,N_14653);
nand U14825 (N_14825,N_14708,N_14684);
nand U14826 (N_14826,N_14630,N_14753);
or U14827 (N_14827,N_14689,N_14600);
or U14828 (N_14828,N_14702,N_14744);
nand U14829 (N_14829,N_14626,N_14632);
nand U14830 (N_14830,N_14680,N_14758);
xnor U14831 (N_14831,N_14629,N_14748);
and U14832 (N_14832,N_14725,N_14701);
nor U14833 (N_14833,N_14649,N_14606);
or U14834 (N_14834,N_14766,N_14756);
and U14835 (N_14835,N_14688,N_14746);
or U14836 (N_14836,N_14789,N_14775);
or U14837 (N_14837,N_14609,N_14646);
or U14838 (N_14838,N_14667,N_14705);
and U14839 (N_14839,N_14767,N_14668);
xnor U14840 (N_14840,N_14715,N_14635);
nor U14841 (N_14841,N_14694,N_14620);
nor U14842 (N_14842,N_14642,N_14628);
xnor U14843 (N_14843,N_14745,N_14735);
xnor U14844 (N_14844,N_14757,N_14771);
nor U14845 (N_14845,N_14683,N_14795);
or U14846 (N_14846,N_14711,N_14777);
or U14847 (N_14847,N_14773,N_14664);
nand U14848 (N_14848,N_14768,N_14623);
or U14849 (N_14849,N_14654,N_14755);
nand U14850 (N_14850,N_14613,N_14732);
nor U14851 (N_14851,N_14660,N_14728);
xnor U14852 (N_14852,N_14610,N_14619);
nor U14853 (N_14853,N_14736,N_14659);
nand U14854 (N_14854,N_14784,N_14614);
xnor U14855 (N_14855,N_14783,N_14709);
xnor U14856 (N_14856,N_14699,N_14769);
or U14857 (N_14857,N_14776,N_14673);
nor U14858 (N_14858,N_14779,N_14786);
and U14859 (N_14859,N_14793,N_14665);
nor U14860 (N_14860,N_14605,N_14622);
xnor U14861 (N_14861,N_14751,N_14601);
nand U14862 (N_14862,N_14681,N_14730);
nor U14863 (N_14863,N_14650,N_14782);
and U14864 (N_14864,N_14750,N_14618);
nand U14865 (N_14865,N_14615,N_14700);
nor U14866 (N_14866,N_14737,N_14703);
xor U14867 (N_14867,N_14686,N_14641);
and U14868 (N_14868,N_14655,N_14608);
or U14869 (N_14869,N_14714,N_14678);
nor U14870 (N_14870,N_14656,N_14706);
and U14871 (N_14871,N_14616,N_14631);
or U14872 (N_14872,N_14621,N_14729);
nand U14873 (N_14873,N_14770,N_14761);
and U14874 (N_14874,N_14685,N_14774);
and U14875 (N_14875,N_14687,N_14676);
nand U14876 (N_14876,N_14719,N_14627);
xor U14877 (N_14877,N_14741,N_14787);
or U14878 (N_14878,N_14781,N_14604);
nand U14879 (N_14879,N_14638,N_14692);
nor U14880 (N_14880,N_14698,N_14617);
xnor U14881 (N_14881,N_14682,N_14669);
xor U14882 (N_14882,N_14704,N_14762);
xnor U14883 (N_14883,N_14675,N_14657);
or U14884 (N_14884,N_14634,N_14677);
nor U14885 (N_14885,N_14718,N_14712);
nor U14886 (N_14886,N_14637,N_14734);
nor U14887 (N_14887,N_14663,N_14724);
nor U14888 (N_14888,N_14661,N_14791);
xnor U14889 (N_14889,N_14636,N_14759);
xnor U14890 (N_14890,N_14772,N_14670);
and U14891 (N_14891,N_14697,N_14740);
or U14892 (N_14892,N_14796,N_14643);
and U14893 (N_14893,N_14738,N_14760);
and U14894 (N_14894,N_14742,N_14710);
and U14895 (N_14895,N_14666,N_14625);
nor U14896 (N_14896,N_14790,N_14743);
nor U14897 (N_14897,N_14612,N_14658);
and U14898 (N_14898,N_14674,N_14647);
nand U14899 (N_14899,N_14754,N_14707);
nand U14900 (N_14900,N_14699,N_14618);
xor U14901 (N_14901,N_14684,N_14603);
or U14902 (N_14902,N_14711,N_14752);
or U14903 (N_14903,N_14743,N_14735);
or U14904 (N_14904,N_14770,N_14694);
nand U14905 (N_14905,N_14765,N_14654);
and U14906 (N_14906,N_14607,N_14661);
nand U14907 (N_14907,N_14750,N_14670);
nand U14908 (N_14908,N_14606,N_14648);
nor U14909 (N_14909,N_14726,N_14711);
xor U14910 (N_14910,N_14681,N_14680);
or U14911 (N_14911,N_14726,N_14752);
and U14912 (N_14912,N_14690,N_14726);
xnor U14913 (N_14913,N_14743,N_14762);
nor U14914 (N_14914,N_14694,N_14652);
and U14915 (N_14915,N_14628,N_14721);
nor U14916 (N_14916,N_14765,N_14602);
and U14917 (N_14917,N_14774,N_14621);
and U14918 (N_14918,N_14799,N_14636);
and U14919 (N_14919,N_14798,N_14727);
nand U14920 (N_14920,N_14632,N_14722);
and U14921 (N_14921,N_14664,N_14640);
xor U14922 (N_14922,N_14657,N_14640);
nor U14923 (N_14923,N_14685,N_14745);
xor U14924 (N_14924,N_14772,N_14613);
nor U14925 (N_14925,N_14754,N_14693);
xnor U14926 (N_14926,N_14637,N_14728);
or U14927 (N_14927,N_14703,N_14651);
and U14928 (N_14928,N_14669,N_14676);
or U14929 (N_14929,N_14640,N_14795);
or U14930 (N_14930,N_14775,N_14799);
nand U14931 (N_14931,N_14628,N_14610);
nor U14932 (N_14932,N_14696,N_14750);
or U14933 (N_14933,N_14661,N_14615);
nand U14934 (N_14934,N_14729,N_14721);
and U14935 (N_14935,N_14698,N_14700);
nor U14936 (N_14936,N_14789,N_14790);
nor U14937 (N_14937,N_14717,N_14695);
nor U14938 (N_14938,N_14662,N_14625);
xor U14939 (N_14939,N_14698,N_14640);
nand U14940 (N_14940,N_14631,N_14618);
xnor U14941 (N_14941,N_14688,N_14768);
nor U14942 (N_14942,N_14735,N_14637);
or U14943 (N_14943,N_14608,N_14791);
xor U14944 (N_14944,N_14690,N_14776);
xnor U14945 (N_14945,N_14784,N_14697);
xnor U14946 (N_14946,N_14791,N_14688);
or U14947 (N_14947,N_14662,N_14644);
or U14948 (N_14948,N_14793,N_14746);
nor U14949 (N_14949,N_14658,N_14793);
and U14950 (N_14950,N_14699,N_14719);
nor U14951 (N_14951,N_14792,N_14615);
nand U14952 (N_14952,N_14736,N_14693);
or U14953 (N_14953,N_14703,N_14668);
and U14954 (N_14954,N_14666,N_14610);
xor U14955 (N_14955,N_14753,N_14780);
and U14956 (N_14956,N_14612,N_14701);
nand U14957 (N_14957,N_14737,N_14712);
nand U14958 (N_14958,N_14662,N_14694);
nand U14959 (N_14959,N_14696,N_14704);
nor U14960 (N_14960,N_14793,N_14603);
and U14961 (N_14961,N_14674,N_14681);
or U14962 (N_14962,N_14739,N_14754);
nor U14963 (N_14963,N_14762,N_14655);
nor U14964 (N_14964,N_14607,N_14730);
or U14965 (N_14965,N_14735,N_14725);
xor U14966 (N_14966,N_14646,N_14724);
nor U14967 (N_14967,N_14650,N_14768);
or U14968 (N_14968,N_14609,N_14629);
or U14969 (N_14969,N_14683,N_14720);
or U14970 (N_14970,N_14685,N_14740);
or U14971 (N_14971,N_14638,N_14609);
nand U14972 (N_14972,N_14653,N_14603);
nand U14973 (N_14973,N_14781,N_14605);
nor U14974 (N_14974,N_14767,N_14709);
xnor U14975 (N_14975,N_14699,N_14656);
nor U14976 (N_14976,N_14603,N_14631);
xor U14977 (N_14977,N_14720,N_14614);
xnor U14978 (N_14978,N_14719,N_14684);
nand U14979 (N_14979,N_14678,N_14755);
nand U14980 (N_14980,N_14781,N_14743);
nor U14981 (N_14981,N_14752,N_14724);
or U14982 (N_14982,N_14672,N_14799);
nand U14983 (N_14983,N_14652,N_14715);
nand U14984 (N_14984,N_14605,N_14644);
or U14985 (N_14985,N_14749,N_14686);
or U14986 (N_14986,N_14604,N_14613);
xor U14987 (N_14987,N_14772,N_14657);
xor U14988 (N_14988,N_14662,N_14602);
nor U14989 (N_14989,N_14674,N_14776);
nand U14990 (N_14990,N_14790,N_14648);
xnor U14991 (N_14991,N_14795,N_14674);
and U14992 (N_14992,N_14635,N_14753);
or U14993 (N_14993,N_14703,N_14774);
nor U14994 (N_14994,N_14615,N_14757);
or U14995 (N_14995,N_14647,N_14782);
or U14996 (N_14996,N_14669,N_14700);
and U14997 (N_14997,N_14723,N_14718);
or U14998 (N_14998,N_14689,N_14780);
and U14999 (N_14999,N_14691,N_14766);
nor UO_0 (O_0,N_14911,N_14959);
nand UO_1 (O_1,N_14892,N_14812);
and UO_2 (O_2,N_14997,N_14882);
xor UO_3 (O_3,N_14978,N_14855);
xnor UO_4 (O_4,N_14816,N_14998);
xor UO_5 (O_5,N_14826,N_14946);
and UO_6 (O_6,N_14952,N_14989);
xnor UO_7 (O_7,N_14831,N_14994);
nor UO_8 (O_8,N_14836,N_14935);
nor UO_9 (O_9,N_14981,N_14813);
and UO_10 (O_10,N_14907,N_14995);
or UO_11 (O_11,N_14969,N_14954);
nor UO_12 (O_12,N_14865,N_14992);
and UO_13 (O_13,N_14863,N_14829);
nand UO_14 (O_14,N_14948,N_14843);
and UO_15 (O_15,N_14828,N_14929);
nand UO_16 (O_16,N_14899,N_14854);
nand UO_17 (O_17,N_14990,N_14868);
nand UO_18 (O_18,N_14824,N_14887);
xor UO_19 (O_19,N_14877,N_14861);
xnor UO_20 (O_20,N_14934,N_14850);
or UO_21 (O_21,N_14926,N_14975);
or UO_22 (O_22,N_14920,N_14918);
and UO_23 (O_23,N_14962,N_14919);
xor UO_24 (O_24,N_14837,N_14869);
nand UO_25 (O_25,N_14840,N_14936);
nand UO_26 (O_26,N_14885,N_14809);
nand UO_27 (O_27,N_14993,N_14818);
nor UO_28 (O_28,N_14800,N_14910);
and UO_29 (O_29,N_14957,N_14866);
and UO_30 (O_30,N_14968,N_14880);
and UO_31 (O_31,N_14852,N_14808);
nor UO_32 (O_32,N_14950,N_14974);
and UO_33 (O_33,N_14937,N_14961);
or UO_34 (O_34,N_14921,N_14916);
or UO_35 (O_35,N_14943,N_14896);
xnor UO_36 (O_36,N_14847,N_14856);
or UO_37 (O_37,N_14908,N_14979);
or UO_38 (O_38,N_14871,N_14966);
nand UO_39 (O_39,N_14941,N_14985);
nor UO_40 (O_40,N_14940,N_14833);
xor UO_41 (O_41,N_14984,N_14853);
nor UO_42 (O_42,N_14886,N_14963);
nand UO_43 (O_43,N_14864,N_14889);
nor UO_44 (O_44,N_14900,N_14967);
xor UO_45 (O_45,N_14872,N_14817);
nand UO_46 (O_46,N_14841,N_14846);
nand UO_47 (O_47,N_14832,N_14814);
and UO_48 (O_48,N_14858,N_14913);
and UO_49 (O_49,N_14915,N_14905);
nor UO_50 (O_50,N_14901,N_14928);
nand UO_51 (O_51,N_14873,N_14803);
nor UO_52 (O_52,N_14965,N_14951);
and UO_53 (O_53,N_14857,N_14874);
and UO_54 (O_54,N_14890,N_14895);
nand UO_55 (O_55,N_14925,N_14848);
nor UO_56 (O_56,N_14870,N_14999);
nand UO_57 (O_57,N_14912,N_14906);
and UO_58 (O_58,N_14973,N_14932);
nand UO_59 (O_59,N_14835,N_14909);
nor UO_60 (O_60,N_14825,N_14986);
or UO_61 (O_61,N_14867,N_14839);
xnor UO_62 (O_62,N_14804,N_14842);
nor UO_63 (O_63,N_14922,N_14971);
or UO_64 (O_64,N_14914,N_14945);
and UO_65 (O_65,N_14888,N_14811);
xor UO_66 (O_66,N_14830,N_14947);
or UO_67 (O_67,N_14862,N_14875);
nand UO_68 (O_68,N_14976,N_14810);
nor UO_69 (O_69,N_14844,N_14958);
and UO_70 (O_70,N_14987,N_14884);
nor UO_71 (O_71,N_14822,N_14923);
nand UO_72 (O_72,N_14933,N_14893);
nand UO_73 (O_73,N_14819,N_14917);
and UO_74 (O_74,N_14838,N_14815);
and UO_75 (O_75,N_14845,N_14904);
nor UO_76 (O_76,N_14960,N_14964);
xor UO_77 (O_77,N_14805,N_14949);
or UO_78 (O_78,N_14860,N_14883);
nand UO_79 (O_79,N_14927,N_14807);
and UO_80 (O_80,N_14956,N_14879);
and UO_81 (O_81,N_14970,N_14938);
or UO_82 (O_82,N_14980,N_14903);
nand UO_83 (O_83,N_14823,N_14988);
xor UO_84 (O_84,N_14878,N_14942);
nand UO_85 (O_85,N_14894,N_14953);
or UO_86 (O_86,N_14996,N_14897);
nor UO_87 (O_87,N_14972,N_14806);
and UO_88 (O_88,N_14802,N_14898);
nand UO_89 (O_89,N_14827,N_14991);
nand UO_90 (O_90,N_14851,N_14801);
and UO_91 (O_91,N_14820,N_14876);
nor UO_92 (O_92,N_14931,N_14834);
or UO_93 (O_93,N_14891,N_14924);
and UO_94 (O_94,N_14821,N_14902);
or UO_95 (O_95,N_14977,N_14849);
or UO_96 (O_96,N_14939,N_14881);
or UO_97 (O_97,N_14859,N_14930);
xor UO_98 (O_98,N_14944,N_14982);
or UO_99 (O_99,N_14983,N_14955);
and UO_100 (O_100,N_14943,N_14907);
nand UO_101 (O_101,N_14951,N_14889);
nand UO_102 (O_102,N_14857,N_14980);
or UO_103 (O_103,N_14938,N_14903);
and UO_104 (O_104,N_14925,N_14906);
nor UO_105 (O_105,N_14861,N_14827);
xor UO_106 (O_106,N_14890,N_14942);
nor UO_107 (O_107,N_14876,N_14967);
xor UO_108 (O_108,N_14926,N_14956);
and UO_109 (O_109,N_14902,N_14826);
or UO_110 (O_110,N_14893,N_14802);
nand UO_111 (O_111,N_14925,N_14834);
nand UO_112 (O_112,N_14920,N_14999);
or UO_113 (O_113,N_14811,N_14917);
and UO_114 (O_114,N_14925,N_14833);
nand UO_115 (O_115,N_14951,N_14828);
or UO_116 (O_116,N_14926,N_14865);
and UO_117 (O_117,N_14803,N_14982);
xnor UO_118 (O_118,N_14931,N_14837);
and UO_119 (O_119,N_14867,N_14966);
or UO_120 (O_120,N_14885,N_14965);
xor UO_121 (O_121,N_14971,N_14925);
nand UO_122 (O_122,N_14998,N_14872);
nand UO_123 (O_123,N_14948,N_14962);
nor UO_124 (O_124,N_14962,N_14880);
nand UO_125 (O_125,N_14892,N_14846);
nand UO_126 (O_126,N_14870,N_14928);
and UO_127 (O_127,N_14997,N_14893);
and UO_128 (O_128,N_14834,N_14841);
and UO_129 (O_129,N_14818,N_14927);
xor UO_130 (O_130,N_14933,N_14886);
nand UO_131 (O_131,N_14835,N_14878);
and UO_132 (O_132,N_14843,N_14961);
or UO_133 (O_133,N_14825,N_14961);
or UO_134 (O_134,N_14858,N_14866);
nand UO_135 (O_135,N_14854,N_14882);
or UO_136 (O_136,N_14851,N_14866);
or UO_137 (O_137,N_14839,N_14917);
nor UO_138 (O_138,N_14945,N_14950);
and UO_139 (O_139,N_14860,N_14829);
nand UO_140 (O_140,N_14944,N_14861);
nand UO_141 (O_141,N_14802,N_14996);
nor UO_142 (O_142,N_14957,N_14945);
and UO_143 (O_143,N_14991,N_14861);
nor UO_144 (O_144,N_14990,N_14877);
and UO_145 (O_145,N_14927,N_14893);
nand UO_146 (O_146,N_14842,N_14900);
and UO_147 (O_147,N_14885,N_14997);
and UO_148 (O_148,N_14854,N_14917);
nand UO_149 (O_149,N_14960,N_14851);
nor UO_150 (O_150,N_14942,N_14884);
and UO_151 (O_151,N_14876,N_14809);
xor UO_152 (O_152,N_14939,N_14974);
and UO_153 (O_153,N_14986,N_14897);
nor UO_154 (O_154,N_14858,N_14969);
or UO_155 (O_155,N_14974,N_14843);
and UO_156 (O_156,N_14845,N_14888);
nor UO_157 (O_157,N_14828,N_14905);
nor UO_158 (O_158,N_14867,N_14942);
xnor UO_159 (O_159,N_14912,N_14922);
or UO_160 (O_160,N_14924,N_14875);
nand UO_161 (O_161,N_14899,N_14967);
and UO_162 (O_162,N_14990,N_14963);
and UO_163 (O_163,N_14851,N_14943);
or UO_164 (O_164,N_14912,N_14850);
xnor UO_165 (O_165,N_14966,N_14907);
or UO_166 (O_166,N_14862,N_14817);
or UO_167 (O_167,N_14910,N_14994);
nand UO_168 (O_168,N_14855,N_14905);
or UO_169 (O_169,N_14956,N_14960);
and UO_170 (O_170,N_14859,N_14835);
or UO_171 (O_171,N_14980,N_14820);
and UO_172 (O_172,N_14839,N_14883);
or UO_173 (O_173,N_14830,N_14822);
nor UO_174 (O_174,N_14993,N_14873);
and UO_175 (O_175,N_14976,N_14843);
nor UO_176 (O_176,N_14932,N_14966);
and UO_177 (O_177,N_14881,N_14858);
nor UO_178 (O_178,N_14914,N_14971);
and UO_179 (O_179,N_14959,N_14895);
nand UO_180 (O_180,N_14912,N_14962);
xnor UO_181 (O_181,N_14821,N_14945);
nor UO_182 (O_182,N_14892,N_14963);
nand UO_183 (O_183,N_14967,N_14991);
nor UO_184 (O_184,N_14999,N_14929);
nand UO_185 (O_185,N_14973,N_14809);
or UO_186 (O_186,N_14958,N_14893);
xor UO_187 (O_187,N_14927,N_14966);
nor UO_188 (O_188,N_14939,N_14836);
nor UO_189 (O_189,N_14819,N_14928);
or UO_190 (O_190,N_14922,N_14804);
or UO_191 (O_191,N_14920,N_14804);
or UO_192 (O_192,N_14969,N_14856);
or UO_193 (O_193,N_14842,N_14887);
nand UO_194 (O_194,N_14936,N_14827);
nor UO_195 (O_195,N_14867,N_14844);
and UO_196 (O_196,N_14860,N_14937);
xor UO_197 (O_197,N_14813,N_14898);
nor UO_198 (O_198,N_14861,N_14867);
xnor UO_199 (O_199,N_14999,N_14938);
nand UO_200 (O_200,N_14933,N_14841);
and UO_201 (O_201,N_14989,N_14904);
nand UO_202 (O_202,N_14909,N_14834);
xnor UO_203 (O_203,N_14884,N_14875);
nor UO_204 (O_204,N_14867,N_14893);
and UO_205 (O_205,N_14933,N_14906);
and UO_206 (O_206,N_14844,N_14864);
nand UO_207 (O_207,N_14969,N_14813);
xnor UO_208 (O_208,N_14802,N_14897);
or UO_209 (O_209,N_14819,N_14952);
or UO_210 (O_210,N_14862,N_14826);
or UO_211 (O_211,N_14882,N_14938);
nand UO_212 (O_212,N_14891,N_14907);
nor UO_213 (O_213,N_14892,N_14908);
xnor UO_214 (O_214,N_14833,N_14950);
xor UO_215 (O_215,N_14973,N_14840);
and UO_216 (O_216,N_14805,N_14925);
nor UO_217 (O_217,N_14903,N_14896);
and UO_218 (O_218,N_14824,N_14997);
nor UO_219 (O_219,N_14937,N_14810);
nor UO_220 (O_220,N_14854,N_14826);
and UO_221 (O_221,N_14825,N_14937);
nor UO_222 (O_222,N_14983,N_14909);
or UO_223 (O_223,N_14915,N_14864);
nand UO_224 (O_224,N_14943,N_14936);
or UO_225 (O_225,N_14908,N_14837);
and UO_226 (O_226,N_14873,N_14969);
nor UO_227 (O_227,N_14881,N_14859);
xnor UO_228 (O_228,N_14935,N_14881);
nor UO_229 (O_229,N_14996,N_14878);
nand UO_230 (O_230,N_14977,N_14902);
xnor UO_231 (O_231,N_14963,N_14890);
nor UO_232 (O_232,N_14878,N_14897);
and UO_233 (O_233,N_14930,N_14888);
xnor UO_234 (O_234,N_14842,N_14985);
nor UO_235 (O_235,N_14960,N_14856);
nand UO_236 (O_236,N_14824,N_14945);
or UO_237 (O_237,N_14974,N_14867);
nor UO_238 (O_238,N_14803,N_14922);
nand UO_239 (O_239,N_14865,N_14987);
or UO_240 (O_240,N_14986,N_14849);
and UO_241 (O_241,N_14974,N_14891);
or UO_242 (O_242,N_14943,N_14823);
or UO_243 (O_243,N_14885,N_14855);
xnor UO_244 (O_244,N_14935,N_14820);
nor UO_245 (O_245,N_14802,N_14980);
and UO_246 (O_246,N_14816,N_14973);
and UO_247 (O_247,N_14898,N_14922);
nor UO_248 (O_248,N_14835,N_14837);
nor UO_249 (O_249,N_14847,N_14958);
xor UO_250 (O_250,N_14841,N_14892);
xnor UO_251 (O_251,N_14967,N_14891);
or UO_252 (O_252,N_14837,N_14997);
and UO_253 (O_253,N_14825,N_14863);
or UO_254 (O_254,N_14861,N_14903);
nand UO_255 (O_255,N_14888,N_14866);
nor UO_256 (O_256,N_14807,N_14814);
or UO_257 (O_257,N_14822,N_14805);
nand UO_258 (O_258,N_14838,N_14809);
nand UO_259 (O_259,N_14967,N_14844);
or UO_260 (O_260,N_14887,N_14825);
nand UO_261 (O_261,N_14883,N_14897);
xor UO_262 (O_262,N_14894,N_14945);
nor UO_263 (O_263,N_14998,N_14900);
or UO_264 (O_264,N_14875,N_14991);
and UO_265 (O_265,N_14814,N_14911);
nand UO_266 (O_266,N_14833,N_14954);
xnor UO_267 (O_267,N_14836,N_14919);
and UO_268 (O_268,N_14948,N_14824);
nand UO_269 (O_269,N_14892,N_14870);
nor UO_270 (O_270,N_14948,N_14869);
nor UO_271 (O_271,N_14914,N_14976);
nor UO_272 (O_272,N_14939,N_14923);
xnor UO_273 (O_273,N_14876,N_14837);
nand UO_274 (O_274,N_14931,N_14845);
or UO_275 (O_275,N_14843,N_14969);
nor UO_276 (O_276,N_14888,N_14960);
and UO_277 (O_277,N_14911,N_14850);
nor UO_278 (O_278,N_14992,N_14818);
and UO_279 (O_279,N_14898,N_14845);
and UO_280 (O_280,N_14975,N_14801);
nor UO_281 (O_281,N_14848,N_14845);
nor UO_282 (O_282,N_14952,N_14872);
or UO_283 (O_283,N_14845,N_14843);
nand UO_284 (O_284,N_14941,N_14913);
or UO_285 (O_285,N_14990,N_14942);
nor UO_286 (O_286,N_14976,N_14801);
or UO_287 (O_287,N_14882,N_14971);
nand UO_288 (O_288,N_14839,N_14874);
xnor UO_289 (O_289,N_14967,N_14867);
and UO_290 (O_290,N_14937,N_14892);
and UO_291 (O_291,N_14810,N_14803);
and UO_292 (O_292,N_14861,N_14977);
nand UO_293 (O_293,N_14814,N_14861);
nand UO_294 (O_294,N_14831,N_14979);
xor UO_295 (O_295,N_14858,N_14997);
or UO_296 (O_296,N_14984,N_14915);
nand UO_297 (O_297,N_14874,N_14867);
xnor UO_298 (O_298,N_14861,N_14866);
nor UO_299 (O_299,N_14817,N_14926);
xnor UO_300 (O_300,N_14878,N_14819);
nand UO_301 (O_301,N_14857,N_14821);
xor UO_302 (O_302,N_14964,N_14999);
and UO_303 (O_303,N_14900,N_14884);
nand UO_304 (O_304,N_14940,N_14836);
xor UO_305 (O_305,N_14958,N_14968);
nand UO_306 (O_306,N_14835,N_14958);
and UO_307 (O_307,N_14831,N_14930);
xnor UO_308 (O_308,N_14859,N_14961);
xnor UO_309 (O_309,N_14899,N_14961);
xor UO_310 (O_310,N_14842,N_14846);
nor UO_311 (O_311,N_14916,N_14954);
xor UO_312 (O_312,N_14875,N_14987);
nor UO_313 (O_313,N_14850,N_14998);
or UO_314 (O_314,N_14836,N_14810);
nor UO_315 (O_315,N_14822,N_14835);
xnor UO_316 (O_316,N_14802,N_14816);
xnor UO_317 (O_317,N_14867,N_14815);
and UO_318 (O_318,N_14804,N_14988);
xor UO_319 (O_319,N_14962,N_14811);
nor UO_320 (O_320,N_14814,N_14831);
or UO_321 (O_321,N_14804,N_14909);
and UO_322 (O_322,N_14944,N_14805);
nor UO_323 (O_323,N_14948,N_14836);
nand UO_324 (O_324,N_14943,N_14802);
nor UO_325 (O_325,N_14959,N_14831);
nor UO_326 (O_326,N_14878,N_14958);
nand UO_327 (O_327,N_14963,N_14976);
or UO_328 (O_328,N_14827,N_14870);
and UO_329 (O_329,N_14835,N_14955);
xor UO_330 (O_330,N_14846,N_14824);
xor UO_331 (O_331,N_14912,N_14867);
xor UO_332 (O_332,N_14944,N_14836);
nor UO_333 (O_333,N_14803,N_14901);
and UO_334 (O_334,N_14841,N_14900);
nand UO_335 (O_335,N_14973,N_14996);
xnor UO_336 (O_336,N_14871,N_14981);
or UO_337 (O_337,N_14846,N_14957);
xnor UO_338 (O_338,N_14933,N_14936);
nor UO_339 (O_339,N_14872,N_14977);
nand UO_340 (O_340,N_14822,N_14916);
and UO_341 (O_341,N_14925,N_14958);
and UO_342 (O_342,N_14838,N_14875);
nor UO_343 (O_343,N_14842,N_14869);
and UO_344 (O_344,N_14934,N_14951);
or UO_345 (O_345,N_14808,N_14887);
or UO_346 (O_346,N_14829,N_14861);
and UO_347 (O_347,N_14877,N_14908);
xnor UO_348 (O_348,N_14890,N_14861);
xnor UO_349 (O_349,N_14888,N_14997);
nand UO_350 (O_350,N_14859,N_14942);
nand UO_351 (O_351,N_14981,N_14968);
nand UO_352 (O_352,N_14861,N_14874);
nand UO_353 (O_353,N_14948,N_14816);
or UO_354 (O_354,N_14845,N_14994);
nand UO_355 (O_355,N_14962,N_14872);
or UO_356 (O_356,N_14810,N_14878);
nor UO_357 (O_357,N_14982,N_14829);
or UO_358 (O_358,N_14827,N_14884);
nand UO_359 (O_359,N_14992,N_14981);
nand UO_360 (O_360,N_14830,N_14868);
and UO_361 (O_361,N_14949,N_14947);
xnor UO_362 (O_362,N_14823,N_14878);
or UO_363 (O_363,N_14862,N_14815);
nand UO_364 (O_364,N_14827,N_14830);
xor UO_365 (O_365,N_14995,N_14927);
or UO_366 (O_366,N_14957,N_14890);
or UO_367 (O_367,N_14929,N_14946);
xor UO_368 (O_368,N_14947,N_14870);
or UO_369 (O_369,N_14807,N_14943);
xor UO_370 (O_370,N_14844,N_14834);
and UO_371 (O_371,N_14885,N_14864);
nor UO_372 (O_372,N_14832,N_14851);
and UO_373 (O_373,N_14937,N_14847);
nor UO_374 (O_374,N_14845,N_14840);
nor UO_375 (O_375,N_14822,N_14938);
or UO_376 (O_376,N_14984,N_14897);
nor UO_377 (O_377,N_14990,N_14991);
or UO_378 (O_378,N_14996,N_14919);
nor UO_379 (O_379,N_14800,N_14881);
or UO_380 (O_380,N_14981,N_14927);
or UO_381 (O_381,N_14965,N_14925);
and UO_382 (O_382,N_14985,N_14809);
and UO_383 (O_383,N_14852,N_14995);
and UO_384 (O_384,N_14866,N_14825);
nand UO_385 (O_385,N_14870,N_14934);
and UO_386 (O_386,N_14870,N_14948);
or UO_387 (O_387,N_14962,N_14838);
nor UO_388 (O_388,N_14872,N_14921);
nand UO_389 (O_389,N_14991,N_14841);
nand UO_390 (O_390,N_14984,N_14903);
or UO_391 (O_391,N_14829,N_14804);
xnor UO_392 (O_392,N_14907,N_14974);
or UO_393 (O_393,N_14824,N_14943);
and UO_394 (O_394,N_14925,N_14895);
nand UO_395 (O_395,N_14841,N_14946);
nor UO_396 (O_396,N_14825,N_14844);
xnor UO_397 (O_397,N_14838,N_14989);
nand UO_398 (O_398,N_14836,N_14818);
nand UO_399 (O_399,N_14819,N_14908);
xor UO_400 (O_400,N_14825,N_14921);
or UO_401 (O_401,N_14931,N_14919);
nor UO_402 (O_402,N_14942,N_14921);
and UO_403 (O_403,N_14904,N_14891);
nand UO_404 (O_404,N_14945,N_14848);
and UO_405 (O_405,N_14844,N_14959);
xor UO_406 (O_406,N_14969,N_14838);
xor UO_407 (O_407,N_14840,N_14950);
and UO_408 (O_408,N_14968,N_14999);
xor UO_409 (O_409,N_14806,N_14988);
xnor UO_410 (O_410,N_14801,N_14875);
nand UO_411 (O_411,N_14830,N_14951);
xnor UO_412 (O_412,N_14968,N_14980);
nand UO_413 (O_413,N_14811,N_14891);
nand UO_414 (O_414,N_14879,N_14914);
xnor UO_415 (O_415,N_14932,N_14881);
and UO_416 (O_416,N_14831,N_14982);
and UO_417 (O_417,N_14993,N_14998);
or UO_418 (O_418,N_14939,N_14960);
nor UO_419 (O_419,N_14895,N_14909);
or UO_420 (O_420,N_14828,N_14837);
nor UO_421 (O_421,N_14807,N_14847);
and UO_422 (O_422,N_14881,N_14802);
nand UO_423 (O_423,N_14995,N_14936);
nand UO_424 (O_424,N_14985,N_14883);
xnor UO_425 (O_425,N_14820,N_14906);
and UO_426 (O_426,N_14926,N_14896);
nor UO_427 (O_427,N_14967,N_14869);
nor UO_428 (O_428,N_14974,N_14978);
or UO_429 (O_429,N_14891,N_14853);
nand UO_430 (O_430,N_14841,N_14825);
nand UO_431 (O_431,N_14977,N_14856);
nand UO_432 (O_432,N_14932,N_14997);
nor UO_433 (O_433,N_14928,N_14973);
or UO_434 (O_434,N_14950,N_14858);
and UO_435 (O_435,N_14978,N_14915);
nand UO_436 (O_436,N_14824,N_14996);
nand UO_437 (O_437,N_14811,N_14807);
or UO_438 (O_438,N_14873,N_14805);
and UO_439 (O_439,N_14997,N_14836);
and UO_440 (O_440,N_14876,N_14828);
or UO_441 (O_441,N_14962,N_14864);
xor UO_442 (O_442,N_14978,N_14919);
xor UO_443 (O_443,N_14910,N_14905);
nand UO_444 (O_444,N_14831,N_14901);
and UO_445 (O_445,N_14809,N_14888);
or UO_446 (O_446,N_14874,N_14956);
and UO_447 (O_447,N_14997,N_14941);
nor UO_448 (O_448,N_14890,N_14935);
or UO_449 (O_449,N_14956,N_14970);
or UO_450 (O_450,N_14825,N_14882);
and UO_451 (O_451,N_14915,N_14814);
and UO_452 (O_452,N_14804,N_14979);
xor UO_453 (O_453,N_14828,N_14989);
nor UO_454 (O_454,N_14961,N_14811);
nand UO_455 (O_455,N_14970,N_14916);
nor UO_456 (O_456,N_14835,N_14843);
and UO_457 (O_457,N_14902,N_14981);
or UO_458 (O_458,N_14800,N_14864);
or UO_459 (O_459,N_14801,N_14987);
nor UO_460 (O_460,N_14996,N_14909);
xnor UO_461 (O_461,N_14936,N_14808);
xor UO_462 (O_462,N_14812,N_14969);
or UO_463 (O_463,N_14919,N_14890);
and UO_464 (O_464,N_14807,N_14935);
and UO_465 (O_465,N_14895,N_14807);
nor UO_466 (O_466,N_14916,N_14844);
xor UO_467 (O_467,N_14981,N_14910);
nand UO_468 (O_468,N_14857,N_14961);
and UO_469 (O_469,N_14981,N_14864);
nand UO_470 (O_470,N_14979,N_14940);
nor UO_471 (O_471,N_14817,N_14832);
nor UO_472 (O_472,N_14886,N_14851);
or UO_473 (O_473,N_14999,N_14888);
nand UO_474 (O_474,N_14952,N_14843);
xnor UO_475 (O_475,N_14887,N_14959);
or UO_476 (O_476,N_14805,N_14887);
nand UO_477 (O_477,N_14953,N_14984);
nor UO_478 (O_478,N_14979,N_14841);
nand UO_479 (O_479,N_14917,N_14968);
xnor UO_480 (O_480,N_14893,N_14805);
xor UO_481 (O_481,N_14946,N_14837);
or UO_482 (O_482,N_14920,N_14842);
nand UO_483 (O_483,N_14893,N_14939);
xnor UO_484 (O_484,N_14922,N_14878);
nand UO_485 (O_485,N_14984,N_14816);
xnor UO_486 (O_486,N_14895,N_14967);
nand UO_487 (O_487,N_14927,N_14959);
xor UO_488 (O_488,N_14989,N_14915);
and UO_489 (O_489,N_14978,N_14801);
nor UO_490 (O_490,N_14846,N_14945);
xnor UO_491 (O_491,N_14990,N_14843);
and UO_492 (O_492,N_14914,N_14870);
xor UO_493 (O_493,N_14971,N_14823);
nor UO_494 (O_494,N_14946,N_14984);
and UO_495 (O_495,N_14949,N_14826);
nor UO_496 (O_496,N_14972,N_14884);
and UO_497 (O_497,N_14858,N_14956);
nand UO_498 (O_498,N_14858,N_14863);
nand UO_499 (O_499,N_14837,N_14892);
or UO_500 (O_500,N_14995,N_14910);
nand UO_501 (O_501,N_14961,N_14824);
or UO_502 (O_502,N_14993,N_14891);
or UO_503 (O_503,N_14921,N_14817);
nor UO_504 (O_504,N_14938,N_14863);
and UO_505 (O_505,N_14947,N_14896);
nand UO_506 (O_506,N_14893,N_14823);
xnor UO_507 (O_507,N_14942,N_14903);
or UO_508 (O_508,N_14914,N_14845);
or UO_509 (O_509,N_14844,N_14852);
nor UO_510 (O_510,N_14969,N_14916);
nand UO_511 (O_511,N_14867,N_14811);
xnor UO_512 (O_512,N_14887,N_14876);
xnor UO_513 (O_513,N_14991,N_14937);
xnor UO_514 (O_514,N_14934,N_14981);
nor UO_515 (O_515,N_14891,N_14822);
xor UO_516 (O_516,N_14810,N_14883);
nand UO_517 (O_517,N_14858,N_14979);
or UO_518 (O_518,N_14944,N_14830);
or UO_519 (O_519,N_14933,N_14972);
xor UO_520 (O_520,N_14987,N_14985);
xnor UO_521 (O_521,N_14953,N_14866);
and UO_522 (O_522,N_14979,N_14988);
and UO_523 (O_523,N_14996,N_14851);
nor UO_524 (O_524,N_14987,N_14956);
nor UO_525 (O_525,N_14874,N_14922);
or UO_526 (O_526,N_14966,N_14947);
xnor UO_527 (O_527,N_14849,N_14909);
and UO_528 (O_528,N_14978,N_14996);
or UO_529 (O_529,N_14889,N_14857);
nor UO_530 (O_530,N_14944,N_14967);
and UO_531 (O_531,N_14954,N_14979);
nand UO_532 (O_532,N_14827,N_14812);
nand UO_533 (O_533,N_14883,N_14885);
nand UO_534 (O_534,N_14924,N_14958);
nor UO_535 (O_535,N_14985,N_14956);
nor UO_536 (O_536,N_14970,N_14886);
nor UO_537 (O_537,N_14961,N_14822);
nand UO_538 (O_538,N_14920,N_14960);
xnor UO_539 (O_539,N_14826,N_14855);
or UO_540 (O_540,N_14846,N_14818);
nor UO_541 (O_541,N_14927,N_14963);
or UO_542 (O_542,N_14856,N_14898);
nand UO_543 (O_543,N_14816,N_14907);
and UO_544 (O_544,N_14992,N_14894);
nand UO_545 (O_545,N_14933,N_14842);
nor UO_546 (O_546,N_14922,N_14983);
xnor UO_547 (O_547,N_14828,N_14942);
or UO_548 (O_548,N_14854,N_14802);
xor UO_549 (O_549,N_14973,N_14813);
or UO_550 (O_550,N_14954,N_14843);
nand UO_551 (O_551,N_14837,N_14992);
nor UO_552 (O_552,N_14900,N_14960);
or UO_553 (O_553,N_14971,N_14965);
xnor UO_554 (O_554,N_14976,N_14919);
nand UO_555 (O_555,N_14851,N_14859);
or UO_556 (O_556,N_14969,N_14946);
and UO_557 (O_557,N_14997,N_14821);
xnor UO_558 (O_558,N_14813,N_14803);
or UO_559 (O_559,N_14968,N_14898);
or UO_560 (O_560,N_14978,N_14863);
or UO_561 (O_561,N_14854,N_14897);
or UO_562 (O_562,N_14990,N_14836);
and UO_563 (O_563,N_14984,N_14931);
or UO_564 (O_564,N_14859,N_14810);
nand UO_565 (O_565,N_14945,N_14868);
xor UO_566 (O_566,N_14979,N_14896);
nand UO_567 (O_567,N_14942,N_14938);
nor UO_568 (O_568,N_14825,N_14870);
and UO_569 (O_569,N_14974,N_14946);
xor UO_570 (O_570,N_14855,N_14823);
nand UO_571 (O_571,N_14968,N_14918);
nor UO_572 (O_572,N_14960,N_14936);
and UO_573 (O_573,N_14936,N_14922);
or UO_574 (O_574,N_14936,N_14898);
xnor UO_575 (O_575,N_14826,N_14915);
nor UO_576 (O_576,N_14840,N_14853);
nor UO_577 (O_577,N_14929,N_14867);
xor UO_578 (O_578,N_14960,N_14968);
or UO_579 (O_579,N_14965,N_14927);
or UO_580 (O_580,N_14902,N_14822);
and UO_581 (O_581,N_14989,N_14899);
or UO_582 (O_582,N_14806,N_14864);
nand UO_583 (O_583,N_14901,N_14808);
nand UO_584 (O_584,N_14891,N_14984);
and UO_585 (O_585,N_14970,N_14802);
xnor UO_586 (O_586,N_14909,N_14857);
nor UO_587 (O_587,N_14899,N_14864);
xor UO_588 (O_588,N_14911,N_14919);
and UO_589 (O_589,N_14884,N_14837);
nor UO_590 (O_590,N_14848,N_14832);
nand UO_591 (O_591,N_14838,N_14852);
and UO_592 (O_592,N_14906,N_14917);
xnor UO_593 (O_593,N_14957,N_14875);
nand UO_594 (O_594,N_14884,N_14835);
and UO_595 (O_595,N_14936,N_14925);
or UO_596 (O_596,N_14919,N_14865);
nor UO_597 (O_597,N_14996,N_14924);
and UO_598 (O_598,N_14953,N_14930);
xnor UO_599 (O_599,N_14996,N_14871);
nand UO_600 (O_600,N_14844,N_14804);
nor UO_601 (O_601,N_14821,N_14953);
nor UO_602 (O_602,N_14840,N_14986);
nor UO_603 (O_603,N_14887,N_14993);
or UO_604 (O_604,N_14846,N_14979);
xnor UO_605 (O_605,N_14816,N_14875);
xor UO_606 (O_606,N_14942,N_14977);
nand UO_607 (O_607,N_14879,N_14851);
nor UO_608 (O_608,N_14802,N_14876);
or UO_609 (O_609,N_14973,N_14855);
and UO_610 (O_610,N_14998,N_14857);
and UO_611 (O_611,N_14924,N_14925);
nand UO_612 (O_612,N_14981,N_14858);
or UO_613 (O_613,N_14822,N_14956);
or UO_614 (O_614,N_14951,N_14903);
xnor UO_615 (O_615,N_14970,N_14936);
and UO_616 (O_616,N_14814,N_14986);
nand UO_617 (O_617,N_14949,N_14914);
nand UO_618 (O_618,N_14957,N_14803);
nand UO_619 (O_619,N_14966,N_14979);
nand UO_620 (O_620,N_14901,N_14828);
and UO_621 (O_621,N_14906,N_14818);
or UO_622 (O_622,N_14956,N_14953);
nor UO_623 (O_623,N_14982,N_14964);
nor UO_624 (O_624,N_14813,N_14804);
xnor UO_625 (O_625,N_14961,N_14939);
and UO_626 (O_626,N_14872,N_14965);
nand UO_627 (O_627,N_14905,N_14888);
xnor UO_628 (O_628,N_14825,N_14859);
nor UO_629 (O_629,N_14925,N_14952);
xor UO_630 (O_630,N_14821,N_14977);
and UO_631 (O_631,N_14917,N_14979);
or UO_632 (O_632,N_14949,N_14812);
nand UO_633 (O_633,N_14993,N_14915);
or UO_634 (O_634,N_14929,N_14943);
xor UO_635 (O_635,N_14942,N_14905);
or UO_636 (O_636,N_14990,N_14968);
nand UO_637 (O_637,N_14975,N_14874);
and UO_638 (O_638,N_14873,N_14815);
and UO_639 (O_639,N_14906,N_14852);
or UO_640 (O_640,N_14906,N_14862);
xor UO_641 (O_641,N_14886,N_14812);
xor UO_642 (O_642,N_14846,N_14883);
nor UO_643 (O_643,N_14869,N_14924);
and UO_644 (O_644,N_14966,N_14860);
nand UO_645 (O_645,N_14871,N_14826);
and UO_646 (O_646,N_14981,N_14931);
nand UO_647 (O_647,N_14924,N_14975);
nor UO_648 (O_648,N_14809,N_14859);
xor UO_649 (O_649,N_14967,N_14856);
nor UO_650 (O_650,N_14966,N_14936);
nor UO_651 (O_651,N_14922,N_14864);
nand UO_652 (O_652,N_14802,N_14977);
and UO_653 (O_653,N_14921,N_14900);
xnor UO_654 (O_654,N_14975,N_14868);
or UO_655 (O_655,N_14931,N_14918);
or UO_656 (O_656,N_14874,N_14815);
xor UO_657 (O_657,N_14963,N_14949);
or UO_658 (O_658,N_14916,N_14814);
nor UO_659 (O_659,N_14940,N_14937);
nand UO_660 (O_660,N_14968,N_14951);
nor UO_661 (O_661,N_14914,N_14985);
or UO_662 (O_662,N_14867,N_14924);
and UO_663 (O_663,N_14888,N_14918);
and UO_664 (O_664,N_14986,N_14972);
and UO_665 (O_665,N_14837,N_14961);
or UO_666 (O_666,N_14922,N_14991);
or UO_667 (O_667,N_14994,N_14977);
nand UO_668 (O_668,N_14938,N_14894);
or UO_669 (O_669,N_14967,N_14855);
nor UO_670 (O_670,N_14802,N_14974);
xor UO_671 (O_671,N_14808,N_14810);
xor UO_672 (O_672,N_14953,N_14965);
and UO_673 (O_673,N_14890,N_14968);
nand UO_674 (O_674,N_14966,N_14858);
nand UO_675 (O_675,N_14839,N_14815);
or UO_676 (O_676,N_14975,N_14988);
nor UO_677 (O_677,N_14998,N_14896);
nor UO_678 (O_678,N_14941,N_14830);
nand UO_679 (O_679,N_14850,N_14971);
and UO_680 (O_680,N_14933,N_14894);
or UO_681 (O_681,N_14962,N_14863);
xor UO_682 (O_682,N_14821,N_14877);
and UO_683 (O_683,N_14872,N_14853);
xnor UO_684 (O_684,N_14987,N_14843);
or UO_685 (O_685,N_14809,N_14905);
nor UO_686 (O_686,N_14940,N_14882);
and UO_687 (O_687,N_14980,N_14836);
and UO_688 (O_688,N_14863,N_14852);
nor UO_689 (O_689,N_14957,N_14805);
xnor UO_690 (O_690,N_14996,N_14807);
or UO_691 (O_691,N_14939,N_14885);
nor UO_692 (O_692,N_14863,N_14952);
xor UO_693 (O_693,N_14987,N_14847);
and UO_694 (O_694,N_14823,N_14950);
nor UO_695 (O_695,N_14856,N_14976);
xor UO_696 (O_696,N_14846,N_14815);
nand UO_697 (O_697,N_14942,N_14968);
and UO_698 (O_698,N_14901,N_14804);
and UO_699 (O_699,N_14929,N_14957);
xnor UO_700 (O_700,N_14875,N_14829);
or UO_701 (O_701,N_14955,N_14917);
xnor UO_702 (O_702,N_14984,N_14989);
and UO_703 (O_703,N_14841,N_14891);
nand UO_704 (O_704,N_14819,N_14853);
xor UO_705 (O_705,N_14826,N_14896);
xnor UO_706 (O_706,N_14928,N_14820);
nor UO_707 (O_707,N_14906,N_14930);
and UO_708 (O_708,N_14818,N_14809);
nor UO_709 (O_709,N_14940,N_14958);
xor UO_710 (O_710,N_14945,N_14882);
xnor UO_711 (O_711,N_14975,N_14970);
and UO_712 (O_712,N_14839,N_14915);
nor UO_713 (O_713,N_14841,N_14867);
nand UO_714 (O_714,N_14863,N_14809);
xor UO_715 (O_715,N_14992,N_14810);
xnor UO_716 (O_716,N_14921,N_14839);
and UO_717 (O_717,N_14989,N_14872);
and UO_718 (O_718,N_14933,N_14815);
and UO_719 (O_719,N_14806,N_14921);
and UO_720 (O_720,N_14897,N_14927);
or UO_721 (O_721,N_14886,N_14900);
xor UO_722 (O_722,N_14975,N_14844);
and UO_723 (O_723,N_14836,N_14837);
xnor UO_724 (O_724,N_14865,N_14877);
and UO_725 (O_725,N_14856,N_14850);
and UO_726 (O_726,N_14813,N_14911);
xor UO_727 (O_727,N_14872,N_14873);
and UO_728 (O_728,N_14953,N_14814);
and UO_729 (O_729,N_14944,N_14953);
or UO_730 (O_730,N_14930,N_14811);
and UO_731 (O_731,N_14930,N_14970);
and UO_732 (O_732,N_14954,N_14914);
nor UO_733 (O_733,N_14950,N_14817);
xnor UO_734 (O_734,N_14842,N_14863);
xor UO_735 (O_735,N_14893,N_14840);
and UO_736 (O_736,N_14831,N_14974);
nand UO_737 (O_737,N_14833,N_14843);
and UO_738 (O_738,N_14918,N_14838);
or UO_739 (O_739,N_14978,N_14810);
nor UO_740 (O_740,N_14944,N_14986);
xor UO_741 (O_741,N_14894,N_14977);
nor UO_742 (O_742,N_14975,N_14805);
xor UO_743 (O_743,N_14858,N_14963);
nor UO_744 (O_744,N_14970,N_14895);
nor UO_745 (O_745,N_14959,N_14817);
nor UO_746 (O_746,N_14863,N_14972);
xnor UO_747 (O_747,N_14883,N_14968);
or UO_748 (O_748,N_14844,N_14838);
or UO_749 (O_749,N_14859,N_14857);
xnor UO_750 (O_750,N_14983,N_14836);
xor UO_751 (O_751,N_14816,N_14864);
or UO_752 (O_752,N_14869,N_14894);
nor UO_753 (O_753,N_14957,N_14824);
xnor UO_754 (O_754,N_14843,N_14886);
xor UO_755 (O_755,N_14986,N_14846);
or UO_756 (O_756,N_14994,N_14940);
nand UO_757 (O_757,N_14829,N_14876);
and UO_758 (O_758,N_14840,N_14908);
or UO_759 (O_759,N_14808,N_14879);
nor UO_760 (O_760,N_14883,N_14802);
nand UO_761 (O_761,N_14991,N_14883);
and UO_762 (O_762,N_14920,N_14970);
nand UO_763 (O_763,N_14818,N_14851);
and UO_764 (O_764,N_14880,N_14944);
or UO_765 (O_765,N_14965,N_14934);
nand UO_766 (O_766,N_14929,N_14897);
nand UO_767 (O_767,N_14932,N_14803);
nand UO_768 (O_768,N_14945,N_14855);
and UO_769 (O_769,N_14845,N_14821);
xor UO_770 (O_770,N_14830,N_14874);
nor UO_771 (O_771,N_14946,N_14964);
nor UO_772 (O_772,N_14873,N_14842);
or UO_773 (O_773,N_14862,N_14913);
and UO_774 (O_774,N_14835,N_14992);
and UO_775 (O_775,N_14869,N_14961);
xor UO_776 (O_776,N_14954,N_14862);
or UO_777 (O_777,N_14866,N_14973);
xor UO_778 (O_778,N_14999,N_14969);
or UO_779 (O_779,N_14867,N_14833);
and UO_780 (O_780,N_14994,N_14852);
and UO_781 (O_781,N_14913,N_14879);
and UO_782 (O_782,N_14910,N_14900);
and UO_783 (O_783,N_14945,N_14811);
xor UO_784 (O_784,N_14813,N_14987);
nand UO_785 (O_785,N_14826,N_14929);
nand UO_786 (O_786,N_14969,N_14928);
or UO_787 (O_787,N_14883,N_14906);
nor UO_788 (O_788,N_14953,N_14955);
nor UO_789 (O_789,N_14885,N_14950);
xnor UO_790 (O_790,N_14923,N_14973);
and UO_791 (O_791,N_14873,N_14987);
and UO_792 (O_792,N_14904,N_14986);
xnor UO_793 (O_793,N_14963,N_14936);
nor UO_794 (O_794,N_14927,N_14853);
nor UO_795 (O_795,N_14924,N_14805);
nor UO_796 (O_796,N_14979,N_14848);
or UO_797 (O_797,N_14856,N_14994);
nand UO_798 (O_798,N_14965,N_14933);
nor UO_799 (O_799,N_14892,N_14998);
nor UO_800 (O_800,N_14961,N_14988);
xor UO_801 (O_801,N_14836,N_14957);
or UO_802 (O_802,N_14838,N_14991);
xor UO_803 (O_803,N_14881,N_14951);
nand UO_804 (O_804,N_14991,N_14823);
nor UO_805 (O_805,N_14872,N_14842);
nor UO_806 (O_806,N_14973,N_14957);
or UO_807 (O_807,N_14956,N_14978);
or UO_808 (O_808,N_14960,N_14944);
nand UO_809 (O_809,N_14918,N_14889);
nor UO_810 (O_810,N_14926,N_14823);
nand UO_811 (O_811,N_14923,N_14989);
nand UO_812 (O_812,N_14978,N_14901);
nor UO_813 (O_813,N_14946,N_14909);
nand UO_814 (O_814,N_14876,N_14851);
xnor UO_815 (O_815,N_14849,N_14814);
xnor UO_816 (O_816,N_14856,N_14910);
or UO_817 (O_817,N_14827,N_14954);
nor UO_818 (O_818,N_14857,N_14871);
and UO_819 (O_819,N_14819,N_14854);
nor UO_820 (O_820,N_14860,N_14859);
and UO_821 (O_821,N_14877,N_14934);
and UO_822 (O_822,N_14805,N_14895);
and UO_823 (O_823,N_14849,N_14852);
and UO_824 (O_824,N_14867,N_14920);
nor UO_825 (O_825,N_14804,N_14801);
nand UO_826 (O_826,N_14934,N_14960);
nand UO_827 (O_827,N_14912,N_14882);
nand UO_828 (O_828,N_14951,N_14924);
nor UO_829 (O_829,N_14869,N_14943);
nor UO_830 (O_830,N_14923,N_14870);
nand UO_831 (O_831,N_14989,N_14907);
nand UO_832 (O_832,N_14907,N_14827);
or UO_833 (O_833,N_14826,N_14963);
and UO_834 (O_834,N_14974,N_14870);
nand UO_835 (O_835,N_14922,N_14931);
nor UO_836 (O_836,N_14971,N_14953);
xor UO_837 (O_837,N_14817,N_14981);
nand UO_838 (O_838,N_14861,N_14847);
xnor UO_839 (O_839,N_14913,N_14976);
and UO_840 (O_840,N_14801,N_14889);
or UO_841 (O_841,N_14878,N_14896);
nand UO_842 (O_842,N_14800,N_14823);
or UO_843 (O_843,N_14956,N_14996);
nor UO_844 (O_844,N_14954,N_14800);
nand UO_845 (O_845,N_14992,N_14884);
nand UO_846 (O_846,N_14865,N_14847);
xor UO_847 (O_847,N_14888,N_14836);
and UO_848 (O_848,N_14983,N_14961);
and UO_849 (O_849,N_14891,N_14844);
nor UO_850 (O_850,N_14920,N_14962);
or UO_851 (O_851,N_14911,N_14819);
or UO_852 (O_852,N_14936,N_14871);
xnor UO_853 (O_853,N_14845,N_14810);
and UO_854 (O_854,N_14809,N_14819);
and UO_855 (O_855,N_14951,N_14895);
nand UO_856 (O_856,N_14982,N_14854);
nor UO_857 (O_857,N_14931,N_14862);
or UO_858 (O_858,N_14804,N_14810);
nand UO_859 (O_859,N_14926,N_14917);
nor UO_860 (O_860,N_14884,N_14895);
or UO_861 (O_861,N_14978,N_14982);
and UO_862 (O_862,N_14805,N_14954);
nand UO_863 (O_863,N_14983,N_14875);
and UO_864 (O_864,N_14811,N_14846);
or UO_865 (O_865,N_14935,N_14985);
nand UO_866 (O_866,N_14849,N_14809);
and UO_867 (O_867,N_14935,N_14938);
xnor UO_868 (O_868,N_14901,N_14847);
and UO_869 (O_869,N_14963,N_14926);
nand UO_870 (O_870,N_14970,N_14971);
nand UO_871 (O_871,N_14910,N_14932);
or UO_872 (O_872,N_14839,N_14907);
xnor UO_873 (O_873,N_14816,N_14902);
and UO_874 (O_874,N_14899,N_14859);
xnor UO_875 (O_875,N_14812,N_14951);
and UO_876 (O_876,N_14848,N_14802);
nand UO_877 (O_877,N_14931,N_14913);
nand UO_878 (O_878,N_14977,N_14862);
nor UO_879 (O_879,N_14977,N_14944);
and UO_880 (O_880,N_14811,N_14983);
or UO_881 (O_881,N_14808,N_14970);
xnor UO_882 (O_882,N_14950,N_14826);
or UO_883 (O_883,N_14901,N_14915);
or UO_884 (O_884,N_14868,N_14874);
nor UO_885 (O_885,N_14974,N_14855);
or UO_886 (O_886,N_14839,N_14899);
nand UO_887 (O_887,N_14816,N_14858);
or UO_888 (O_888,N_14899,N_14921);
nor UO_889 (O_889,N_14887,N_14896);
or UO_890 (O_890,N_14859,N_14931);
nand UO_891 (O_891,N_14896,N_14941);
nand UO_892 (O_892,N_14823,N_14977);
xnor UO_893 (O_893,N_14984,N_14965);
or UO_894 (O_894,N_14911,N_14990);
or UO_895 (O_895,N_14934,N_14806);
nor UO_896 (O_896,N_14913,N_14800);
nand UO_897 (O_897,N_14943,N_14942);
or UO_898 (O_898,N_14900,N_14979);
and UO_899 (O_899,N_14981,N_14814);
xnor UO_900 (O_900,N_14948,N_14858);
nand UO_901 (O_901,N_14930,N_14868);
nor UO_902 (O_902,N_14809,N_14894);
nand UO_903 (O_903,N_14955,N_14916);
or UO_904 (O_904,N_14847,N_14804);
xor UO_905 (O_905,N_14852,N_14913);
nand UO_906 (O_906,N_14813,N_14993);
nor UO_907 (O_907,N_14939,N_14826);
and UO_908 (O_908,N_14816,N_14995);
nor UO_909 (O_909,N_14838,N_14950);
or UO_910 (O_910,N_14923,N_14832);
or UO_911 (O_911,N_14853,N_14867);
and UO_912 (O_912,N_14891,N_14826);
nand UO_913 (O_913,N_14850,N_14858);
nor UO_914 (O_914,N_14929,N_14808);
nand UO_915 (O_915,N_14848,N_14924);
nor UO_916 (O_916,N_14843,N_14873);
nor UO_917 (O_917,N_14862,N_14804);
nand UO_918 (O_918,N_14973,N_14900);
or UO_919 (O_919,N_14827,N_14942);
nor UO_920 (O_920,N_14822,N_14880);
and UO_921 (O_921,N_14825,N_14833);
and UO_922 (O_922,N_14820,N_14969);
xnor UO_923 (O_923,N_14933,N_14827);
xor UO_924 (O_924,N_14912,N_14837);
or UO_925 (O_925,N_14819,N_14863);
nand UO_926 (O_926,N_14829,N_14890);
nor UO_927 (O_927,N_14806,N_14837);
and UO_928 (O_928,N_14876,N_14865);
nor UO_929 (O_929,N_14830,N_14806);
nand UO_930 (O_930,N_14937,N_14844);
nor UO_931 (O_931,N_14825,N_14923);
nor UO_932 (O_932,N_14934,N_14993);
xnor UO_933 (O_933,N_14874,N_14921);
xor UO_934 (O_934,N_14903,N_14839);
nor UO_935 (O_935,N_14949,N_14845);
nand UO_936 (O_936,N_14970,N_14862);
xor UO_937 (O_937,N_14883,N_14986);
nand UO_938 (O_938,N_14925,N_14926);
nand UO_939 (O_939,N_14924,N_14938);
or UO_940 (O_940,N_14935,N_14872);
nand UO_941 (O_941,N_14998,N_14809);
or UO_942 (O_942,N_14902,N_14852);
nand UO_943 (O_943,N_14875,N_14888);
nor UO_944 (O_944,N_14818,N_14987);
or UO_945 (O_945,N_14969,N_14853);
or UO_946 (O_946,N_14860,N_14922);
and UO_947 (O_947,N_14879,N_14819);
nor UO_948 (O_948,N_14897,N_14959);
xnor UO_949 (O_949,N_14959,N_14870);
nor UO_950 (O_950,N_14975,N_14890);
and UO_951 (O_951,N_14830,N_14984);
and UO_952 (O_952,N_14909,N_14973);
nand UO_953 (O_953,N_14942,N_14965);
and UO_954 (O_954,N_14994,N_14808);
and UO_955 (O_955,N_14808,N_14838);
xor UO_956 (O_956,N_14959,N_14808);
and UO_957 (O_957,N_14807,N_14833);
nand UO_958 (O_958,N_14829,N_14824);
xor UO_959 (O_959,N_14964,N_14957);
nor UO_960 (O_960,N_14949,N_14894);
or UO_961 (O_961,N_14923,N_14819);
or UO_962 (O_962,N_14890,N_14903);
nand UO_963 (O_963,N_14884,N_14809);
nand UO_964 (O_964,N_14829,N_14897);
nand UO_965 (O_965,N_14899,N_14869);
xor UO_966 (O_966,N_14897,N_14954);
nand UO_967 (O_967,N_14813,N_14991);
nand UO_968 (O_968,N_14915,N_14906);
nor UO_969 (O_969,N_14834,N_14852);
and UO_970 (O_970,N_14849,N_14910);
or UO_971 (O_971,N_14823,N_14949);
nor UO_972 (O_972,N_14993,N_14987);
nor UO_973 (O_973,N_14880,N_14849);
and UO_974 (O_974,N_14808,N_14883);
xnor UO_975 (O_975,N_14831,N_14881);
and UO_976 (O_976,N_14956,N_14856);
nor UO_977 (O_977,N_14942,N_14800);
or UO_978 (O_978,N_14879,N_14935);
and UO_979 (O_979,N_14985,N_14950);
nor UO_980 (O_980,N_14802,N_14995);
or UO_981 (O_981,N_14827,N_14904);
nor UO_982 (O_982,N_14992,N_14929);
and UO_983 (O_983,N_14978,N_14864);
or UO_984 (O_984,N_14865,N_14881);
nand UO_985 (O_985,N_14829,N_14816);
and UO_986 (O_986,N_14989,N_14983);
nor UO_987 (O_987,N_14878,N_14917);
xnor UO_988 (O_988,N_14887,N_14968);
nand UO_989 (O_989,N_14938,N_14825);
xor UO_990 (O_990,N_14905,N_14931);
or UO_991 (O_991,N_14886,N_14946);
and UO_992 (O_992,N_14947,N_14946);
or UO_993 (O_993,N_14878,N_14936);
or UO_994 (O_994,N_14847,N_14919);
xor UO_995 (O_995,N_14982,N_14860);
and UO_996 (O_996,N_14874,N_14927);
xnor UO_997 (O_997,N_14908,N_14902);
and UO_998 (O_998,N_14941,N_14887);
and UO_999 (O_999,N_14925,N_14908);
xor UO_1000 (O_1000,N_14842,N_14912);
nand UO_1001 (O_1001,N_14947,N_14861);
xnor UO_1002 (O_1002,N_14986,N_14905);
xor UO_1003 (O_1003,N_14822,N_14907);
or UO_1004 (O_1004,N_14853,N_14924);
xor UO_1005 (O_1005,N_14944,N_14850);
and UO_1006 (O_1006,N_14943,N_14930);
nor UO_1007 (O_1007,N_14870,N_14955);
xnor UO_1008 (O_1008,N_14981,N_14843);
nor UO_1009 (O_1009,N_14875,N_14863);
nand UO_1010 (O_1010,N_14900,N_14936);
and UO_1011 (O_1011,N_14863,N_14995);
and UO_1012 (O_1012,N_14852,N_14997);
and UO_1013 (O_1013,N_14920,N_14956);
nand UO_1014 (O_1014,N_14974,N_14837);
or UO_1015 (O_1015,N_14886,N_14956);
nor UO_1016 (O_1016,N_14910,N_14830);
xnor UO_1017 (O_1017,N_14980,N_14996);
xnor UO_1018 (O_1018,N_14874,N_14948);
nand UO_1019 (O_1019,N_14836,N_14931);
or UO_1020 (O_1020,N_14968,N_14870);
xor UO_1021 (O_1021,N_14953,N_14962);
and UO_1022 (O_1022,N_14923,N_14975);
xnor UO_1023 (O_1023,N_14901,N_14895);
or UO_1024 (O_1024,N_14834,N_14903);
or UO_1025 (O_1025,N_14886,N_14842);
xor UO_1026 (O_1026,N_14846,N_14801);
nor UO_1027 (O_1027,N_14808,N_14850);
nand UO_1028 (O_1028,N_14904,N_14861);
or UO_1029 (O_1029,N_14937,N_14968);
xnor UO_1030 (O_1030,N_14871,N_14958);
or UO_1031 (O_1031,N_14881,N_14970);
nor UO_1032 (O_1032,N_14912,N_14991);
or UO_1033 (O_1033,N_14977,N_14889);
nand UO_1034 (O_1034,N_14842,N_14945);
nand UO_1035 (O_1035,N_14917,N_14882);
and UO_1036 (O_1036,N_14976,N_14845);
or UO_1037 (O_1037,N_14905,N_14940);
and UO_1038 (O_1038,N_14942,N_14925);
xor UO_1039 (O_1039,N_14854,N_14928);
and UO_1040 (O_1040,N_14885,N_14843);
nor UO_1041 (O_1041,N_14824,N_14932);
nor UO_1042 (O_1042,N_14890,N_14966);
xnor UO_1043 (O_1043,N_14814,N_14948);
nand UO_1044 (O_1044,N_14800,N_14834);
or UO_1045 (O_1045,N_14879,N_14989);
nor UO_1046 (O_1046,N_14864,N_14994);
nand UO_1047 (O_1047,N_14983,N_14812);
or UO_1048 (O_1048,N_14832,N_14888);
nand UO_1049 (O_1049,N_14951,N_14925);
and UO_1050 (O_1050,N_14944,N_14872);
or UO_1051 (O_1051,N_14822,N_14876);
nand UO_1052 (O_1052,N_14841,N_14938);
and UO_1053 (O_1053,N_14971,N_14921);
nand UO_1054 (O_1054,N_14902,N_14953);
and UO_1055 (O_1055,N_14996,N_14915);
and UO_1056 (O_1056,N_14897,N_14863);
or UO_1057 (O_1057,N_14990,N_14831);
nand UO_1058 (O_1058,N_14870,N_14818);
xor UO_1059 (O_1059,N_14967,N_14812);
nand UO_1060 (O_1060,N_14858,N_14835);
or UO_1061 (O_1061,N_14842,N_14976);
and UO_1062 (O_1062,N_14968,N_14924);
nand UO_1063 (O_1063,N_14984,N_14975);
or UO_1064 (O_1064,N_14988,N_14910);
or UO_1065 (O_1065,N_14801,N_14815);
xnor UO_1066 (O_1066,N_14842,N_14967);
and UO_1067 (O_1067,N_14990,N_14951);
and UO_1068 (O_1068,N_14817,N_14836);
nor UO_1069 (O_1069,N_14993,N_14898);
and UO_1070 (O_1070,N_14857,N_14945);
xor UO_1071 (O_1071,N_14888,N_14990);
nor UO_1072 (O_1072,N_14943,N_14898);
nor UO_1073 (O_1073,N_14823,N_14919);
or UO_1074 (O_1074,N_14982,N_14997);
nand UO_1075 (O_1075,N_14999,N_14836);
nand UO_1076 (O_1076,N_14919,N_14834);
or UO_1077 (O_1077,N_14830,N_14879);
or UO_1078 (O_1078,N_14918,N_14976);
nand UO_1079 (O_1079,N_14915,N_14853);
nand UO_1080 (O_1080,N_14839,N_14922);
xnor UO_1081 (O_1081,N_14839,N_14926);
and UO_1082 (O_1082,N_14889,N_14969);
nand UO_1083 (O_1083,N_14820,N_14948);
nor UO_1084 (O_1084,N_14927,N_14924);
nand UO_1085 (O_1085,N_14841,N_14916);
xor UO_1086 (O_1086,N_14812,N_14841);
nand UO_1087 (O_1087,N_14880,N_14834);
or UO_1088 (O_1088,N_14835,N_14907);
xor UO_1089 (O_1089,N_14887,N_14832);
or UO_1090 (O_1090,N_14962,N_14845);
xor UO_1091 (O_1091,N_14855,N_14989);
and UO_1092 (O_1092,N_14842,N_14831);
nand UO_1093 (O_1093,N_14886,N_14898);
or UO_1094 (O_1094,N_14992,N_14889);
nand UO_1095 (O_1095,N_14907,N_14958);
or UO_1096 (O_1096,N_14878,N_14993);
nor UO_1097 (O_1097,N_14862,N_14921);
nand UO_1098 (O_1098,N_14930,N_14855);
or UO_1099 (O_1099,N_14852,N_14928);
or UO_1100 (O_1100,N_14880,N_14961);
xnor UO_1101 (O_1101,N_14867,N_14808);
nor UO_1102 (O_1102,N_14825,N_14949);
nand UO_1103 (O_1103,N_14825,N_14908);
nand UO_1104 (O_1104,N_14849,N_14805);
and UO_1105 (O_1105,N_14953,N_14878);
or UO_1106 (O_1106,N_14855,N_14995);
and UO_1107 (O_1107,N_14934,N_14860);
nor UO_1108 (O_1108,N_14865,N_14864);
nor UO_1109 (O_1109,N_14943,N_14945);
xnor UO_1110 (O_1110,N_14880,N_14940);
and UO_1111 (O_1111,N_14863,N_14999);
or UO_1112 (O_1112,N_14985,N_14929);
and UO_1113 (O_1113,N_14889,N_14900);
and UO_1114 (O_1114,N_14827,N_14838);
or UO_1115 (O_1115,N_14987,N_14849);
nand UO_1116 (O_1116,N_14870,N_14839);
or UO_1117 (O_1117,N_14944,N_14975);
nand UO_1118 (O_1118,N_14959,N_14915);
and UO_1119 (O_1119,N_14809,N_14924);
nand UO_1120 (O_1120,N_14972,N_14848);
nand UO_1121 (O_1121,N_14919,N_14864);
xor UO_1122 (O_1122,N_14946,N_14953);
nand UO_1123 (O_1123,N_14928,N_14894);
nand UO_1124 (O_1124,N_14810,N_14920);
nor UO_1125 (O_1125,N_14820,N_14961);
nor UO_1126 (O_1126,N_14947,N_14940);
nand UO_1127 (O_1127,N_14994,N_14906);
nor UO_1128 (O_1128,N_14901,N_14913);
and UO_1129 (O_1129,N_14815,N_14869);
or UO_1130 (O_1130,N_14864,N_14959);
nor UO_1131 (O_1131,N_14929,N_14990);
xnor UO_1132 (O_1132,N_14873,N_14920);
or UO_1133 (O_1133,N_14869,N_14880);
nand UO_1134 (O_1134,N_14830,N_14979);
or UO_1135 (O_1135,N_14895,N_14855);
nor UO_1136 (O_1136,N_14814,N_14942);
nor UO_1137 (O_1137,N_14973,N_14845);
xor UO_1138 (O_1138,N_14850,N_14997);
and UO_1139 (O_1139,N_14883,N_14861);
nand UO_1140 (O_1140,N_14972,N_14918);
or UO_1141 (O_1141,N_14898,N_14902);
xor UO_1142 (O_1142,N_14987,N_14805);
or UO_1143 (O_1143,N_14854,N_14887);
xnor UO_1144 (O_1144,N_14918,N_14913);
xor UO_1145 (O_1145,N_14898,N_14938);
xor UO_1146 (O_1146,N_14929,N_14806);
and UO_1147 (O_1147,N_14890,N_14940);
or UO_1148 (O_1148,N_14955,N_14800);
xor UO_1149 (O_1149,N_14989,N_14875);
and UO_1150 (O_1150,N_14810,N_14814);
or UO_1151 (O_1151,N_14864,N_14985);
or UO_1152 (O_1152,N_14877,N_14815);
xor UO_1153 (O_1153,N_14855,N_14999);
or UO_1154 (O_1154,N_14847,N_14880);
xnor UO_1155 (O_1155,N_14949,N_14857);
nand UO_1156 (O_1156,N_14806,N_14902);
xor UO_1157 (O_1157,N_14851,N_14968);
and UO_1158 (O_1158,N_14925,N_14915);
and UO_1159 (O_1159,N_14892,N_14936);
nand UO_1160 (O_1160,N_14865,N_14929);
nor UO_1161 (O_1161,N_14954,N_14927);
or UO_1162 (O_1162,N_14954,N_14905);
and UO_1163 (O_1163,N_14813,N_14949);
and UO_1164 (O_1164,N_14859,N_14873);
nand UO_1165 (O_1165,N_14903,N_14966);
nand UO_1166 (O_1166,N_14815,N_14817);
nand UO_1167 (O_1167,N_14963,N_14967);
or UO_1168 (O_1168,N_14989,N_14962);
nor UO_1169 (O_1169,N_14921,N_14913);
and UO_1170 (O_1170,N_14931,N_14982);
or UO_1171 (O_1171,N_14837,N_14913);
xor UO_1172 (O_1172,N_14987,N_14887);
nand UO_1173 (O_1173,N_14914,N_14834);
or UO_1174 (O_1174,N_14889,N_14906);
xnor UO_1175 (O_1175,N_14847,N_14868);
nor UO_1176 (O_1176,N_14969,N_14834);
nor UO_1177 (O_1177,N_14922,N_14947);
nor UO_1178 (O_1178,N_14818,N_14804);
nand UO_1179 (O_1179,N_14935,N_14834);
nand UO_1180 (O_1180,N_14842,N_14880);
xor UO_1181 (O_1181,N_14977,N_14834);
nor UO_1182 (O_1182,N_14972,N_14829);
and UO_1183 (O_1183,N_14956,N_14836);
and UO_1184 (O_1184,N_14820,N_14809);
and UO_1185 (O_1185,N_14984,N_14972);
or UO_1186 (O_1186,N_14877,N_14839);
nor UO_1187 (O_1187,N_14981,N_14946);
xnor UO_1188 (O_1188,N_14862,N_14955);
xnor UO_1189 (O_1189,N_14955,N_14998);
and UO_1190 (O_1190,N_14941,N_14829);
nand UO_1191 (O_1191,N_14978,N_14979);
or UO_1192 (O_1192,N_14940,N_14819);
nor UO_1193 (O_1193,N_14876,N_14900);
or UO_1194 (O_1194,N_14904,N_14843);
nand UO_1195 (O_1195,N_14973,N_14939);
and UO_1196 (O_1196,N_14930,N_14968);
nor UO_1197 (O_1197,N_14866,N_14864);
xnor UO_1198 (O_1198,N_14969,N_14976);
nor UO_1199 (O_1199,N_14990,N_14899);
nand UO_1200 (O_1200,N_14979,N_14808);
nor UO_1201 (O_1201,N_14993,N_14920);
or UO_1202 (O_1202,N_14954,N_14821);
xor UO_1203 (O_1203,N_14979,N_14981);
nor UO_1204 (O_1204,N_14805,N_14865);
nand UO_1205 (O_1205,N_14874,N_14854);
xor UO_1206 (O_1206,N_14846,N_14937);
xnor UO_1207 (O_1207,N_14944,N_14801);
xor UO_1208 (O_1208,N_14910,N_14814);
nor UO_1209 (O_1209,N_14941,N_14904);
and UO_1210 (O_1210,N_14980,N_14901);
xor UO_1211 (O_1211,N_14943,N_14990);
nor UO_1212 (O_1212,N_14803,N_14962);
xor UO_1213 (O_1213,N_14872,N_14920);
or UO_1214 (O_1214,N_14811,N_14875);
or UO_1215 (O_1215,N_14922,N_14846);
nand UO_1216 (O_1216,N_14825,N_14899);
or UO_1217 (O_1217,N_14905,N_14813);
and UO_1218 (O_1218,N_14847,N_14973);
nand UO_1219 (O_1219,N_14995,N_14966);
nand UO_1220 (O_1220,N_14889,N_14805);
and UO_1221 (O_1221,N_14842,N_14995);
and UO_1222 (O_1222,N_14831,N_14894);
nand UO_1223 (O_1223,N_14874,N_14806);
xor UO_1224 (O_1224,N_14873,N_14949);
xor UO_1225 (O_1225,N_14909,N_14830);
or UO_1226 (O_1226,N_14858,N_14842);
xor UO_1227 (O_1227,N_14858,N_14882);
xor UO_1228 (O_1228,N_14807,N_14886);
xnor UO_1229 (O_1229,N_14989,N_14937);
xnor UO_1230 (O_1230,N_14998,N_14935);
and UO_1231 (O_1231,N_14895,N_14898);
nand UO_1232 (O_1232,N_14861,N_14995);
and UO_1233 (O_1233,N_14821,N_14967);
xnor UO_1234 (O_1234,N_14972,N_14946);
nand UO_1235 (O_1235,N_14930,N_14920);
or UO_1236 (O_1236,N_14921,N_14904);
nor UO_1237 (O_1237,N_14800,N_14861);
xnor UO_1238 (O_1238,N_14943,N_14966);
nand UO_1239 (O_1239,N_14983,N_14862);
nor UO_1240 (O_1240,N_14916,N_14942);
and UO_1241 (O_1241,N_14863,N_14955);
and UO_1242 (O_1242,N_14945,N_14962);
xor UO_1243 (O_1243,N_14846,N_14879);
or UO_1244 (O_1244,N_14910,N_14970);
nand UO_1245 (O_1245,N_14816,N_14889);
or UO_1246 (O_1246,N_14973,N_14877);
xnor UO_1247 (O_1247,N_14936,N_14814);
xor UO_1248 (O_1248,N_14843,N_14905);
and UO_1249 (O_1249,N_14986,N_14879);
nor UO_1250 (O_1250,N_14966,N_14928);
xor UO_1251 (O_1251,N_14961,N_14998);
and UO_1252 (O_1252,N_14893,N_14877);
or UO_1253 (O_1253,N_14867,N_14957);
or UO_1254 (O_1254,N_14949,N_14875);
xnor UO_1255 (O_1255,N_14892,N_14880);
nand UO_1256 (O_1256,N_14850,N_14885);
nor UO_1257 (O_1257,N_14894,N_14975);
and UO_1258 (O_1258,N_14929,N_14868);
or UO_1259 (O_1259,N_14863,N_14964);
nand UO_1260 (O_1260,N_14877,N_14919);
xor UO_1261 (O_1261,N_14873,N_14833);
xor UO_1262 (O_1262,N_14826,N_14965);
or UO_1263 (O_1263,N_14925,N_14861);
xor UO_1264 (O_1264,N_14939,N_14936);
nand UO_1265 (O_1265,N_14907,N_14922);
and UO_1266 (O_1266,N_14816,N_14993);
nor UO_1267 (O_1267,N_14994,N_14946);
nand UO_1268 (O_1268,N_14931,N_14860);
and UO_1269 (O_1269,N_14803,N_14890);
xor UO_1270 (O_1270,N_14997,N_14833);
nor UO_1271 (O_1271,N_14913,N_14828);
and UO_1272 (O_1272,N_14894,N_14902);
nor UO_1273 (O_1273,N_14912,N_14826);
and UO_1274 (O_1274,N_14920,N_14933);
nor UO_1275 (O_1275,N_14807,N_14998);
or UO_1276 (O_1276,N_14899,N_14843);
nand UO_1277 (O_1277,N_14949,N_14848);
nand UO_1278 (O_1278,N_14913,N_14816);
and UO_1279 (O_1279,N_14985,N_14873);
nand UO_1280 (O_1280,N_14828,N_14974);
nor UO_1281 (O_1281,N_14960,N_14970);
nor UO_1282 (O_1282,N_14915,N_14985);
nand UO_1283 (O_1283,N_14894,N_14976);
nand UO_1284 (O_1284,N_14933,N_14945);
nor UO_1285 (O_1285,N_14810,N_14842);
or UO_1286 (O_1286,N_14831,N_14801);
and UO_1287 (O_1287,N_14972,N_14834);
xor UO_1288 (O_1288,N_14948,N_14944);
and UO_1289 (O_1289,N_14928,N_14979);
nor UO_1290 (O_1290,N_14924,N_14871);
and UO_1291 (O_1291,N_14897,N_14833);
xor UO_1292 (O_1292,N_14949,N_14912);
nor UO_1293 (O_1293,N_14820,N_14858);
xnor UO_1294 (O_1294,N_14894,N_14916);
nand UO_1295 (O_1295,N_14921,N_14987);
nand UO_1296 (O_1296,N_14840,N_14977);
nand UO_1297 (O_1297,N_14966,N_14961);
and UO_1298 (O_1298,N_14900,N_14968);
nor UO_1299 (O_1299,N_14934,N_14999);
nor UO_1300 (O_1300,N_14869,N_14870);
nor UO_1301 (O_1301,N_14884,N_14990);
nor UO_1302 (O_1302,N_14975,N_14813);
xnor UO_1303 (O_1303,N_14810,N_14918);
and UO_1304 (O_1304,N_14834,N_14853);
xnor UO_1305 (O_1305,N_14969,N_14808);
or UO_1306 (O_1306,N_14999,N_14944);
or UO_1307 (O_1307,N_14957,N_14990);
xnor UO_1308 (O_1308,N_14869,N_14913);
and UO_1309 (O_1309,N_14990,N_14924);
nand UO_1310 (O_1310,N_14926,N_14813);
or UO_1311 (O_1311,N_14912,N_14840);
and UO_1312 (O_1312,N_14822,N_14878);
nor UO_1313 (O_1313,N_14921,N_14894);
nor UO_1314 (O_1314,N_14970,N_14953);
xor UO_1315 (O_1315,N_14858,N_14878);
and UO_1316 (O_1316,N_14985,N_14819);
xnor UO_1317 (O_1317,N_14808,N_14865);
and UO_1318 (O_1318,N_14945,N_14913);
and UO_1319 (O_1319,N_14952,N_14963);
and UO_1320 (O_1320,N_14928,N_14816);
nor UO_1321 (O_1321,N_14918,N_14934);
or UO_1322 (O_1322,N_14858,N_14805);
xor UO_1323 (O_1323,N_14947,N_14924);
xnor UO_1324 (O_1324,N_14871,N_14837);
or UO_1325 (O_1325,N_14927,N_14904);
and UO_1326 (O_1326,N_14861,N_14941);
nor UO_1327 (O_1327,N_14890,N_14918);
and UO_1328 (O_1328,N_14924,N_14970);
and UO_1329 (O_1329,N_14921,N_14923);
nand UO_1330 (O_1330,N_14965,N_14810);
and UO_1331 (O_1331,N_14863,N_14802);
or UO_1332 (O_1332,N_14944,N_14803);
and UO_1333 (O_1333,N_14861,N_14885);
xnor UO_1334 (O_1334,N_14929,N_14958);
nor UO_1335 (O_1335,N_14990,N_14940);
nand UO_1336 (O_1336,N_14991,N_14919);
nor UO_1337 (O_1337,N_14917,N_14901);
or UO_1338 (O_1338,N_14952,N_14805);
and UO_1339 (O_1339,N_14989,N_14993);
nand UO_1340 (O_1340,N_14944,N_14870);
and UO_1341 (O_1341,N_14995,N_14895);
nand UO_1342 (O_1342,N_14806,N_14930);
nor UO_1343 (O_1343,N_14986,N_14821);
and UO_1344 (O_1344,N_14963,N_14954);
or UO_1345 (O_1345,N_14950,N_14805);
nor UO_1346 (O_1346,N_14838,N_14841);
and UO_1347 (O_1347,N_14892,N_14988);
and UO_1348 (O_1348,N_14998,N_14813);
or UO_1349 (O_1349,N_14942,N_14970);
and UO_1350 (O_1350,N_14955,N_14807);
nand UO_1351 (O_1351,N_14879,N_14912);
or UO_1352 (O_1352,N_14997,N_14998);
or UO_1353 (O_1353,N_14860,N_14944);
nand UO_1354 (O_1354,N_14904,N_14961);
xor UO_1355 (O_1355,N_14920,N_14814);
xor UO_1356 (O_1356,N_14824,N_14896);
xor UO_1357 (O_1357,N_14886,N_14883);
nand UO_1358 (O_1358,N_14993,N_14988);
xnor UO_1359 (O_1359,N_14894,N_14829);
or UO_1360 (O_1360,N_14946,N_14834);
nand UO_1361 (O_1361,N_14826,N_14962);
or UO_1362 (O_1362,N_14854,N_14988);
and UO_1363 (O_1363,N_14887,N_14871);
xor UO_1364 (O_1364,N_14825,N_14985);
or UO_1365 (O_1365,N_14819,N_14962);
and UO_1366 (O_1366,N_14984,N_14810);
and UO_1367 (O_1367,N_14954,N_14810);
nand UO_1368 (O_1368,N_14970,N_14943);
or UO_1369 (O_1369,N_14857,N_14968);
nor UO_1370 (O_1370,N_14828,N_14804);
or UO_1371 (O_1371,N_14949,N_14931);
or UO_1372 (O_1372,N_14927,N_14907);
or UO_1373 (O_1373,N_14820,N_14827);
and UO_1374 (O_1374,N_14867,N_14854);
nor UO_1375 (O_1375,N_14981,N_14842);
nor UO_1376 (O_1376,N_14857,N_14947);
nand UO_1377 (O_1377,N_14914,N_14829);
nand UO_1378 (O_1378,N_14911,N_14805);
or UO_1379 (O_1379,N_14800,N_14990);
and UO_1380 (O_1380,N_14852,N_14935);
xnor UO_1381 (O_1381,N_14909,N_14845);
nand UO_1382 (O_1382,N_14883,N_14844);
or UO_1383 (O_1383,N_14848,N_14955);
nor UO_1384 (O_1384,N_14971,N_14876);
xnor UO_1385 (O_1385,N_14877,N_14944);
and UO_1386 (O_1386,N_14967,N_14851);
xor UO_1387 (O_1387,N_14844,N_14875);
xor UO_1388 (O_1388,N_14816,N_14905);
or UO_1389 (O_1389,N_14840,N_14881);
xnor UO_1390 (O_1390,N_14926,N_14961);
or UO_1391 (O_1391,N_14960,N_14986);
nor UO_1392 (O_1392,N_14868,N_14837);
and UO_1393 (O_1393,N_14894,N_14842);
nor UO_1394 (O_1394,N_14961,N_14962);
nor UO_1395 (O_1395,N_14839,N_14893);
xor UO_1396 (O_1396,N_14809,N_14837);
nor UO_1397 (O_1397,N_14853,N_14992);
and UO_1398 (O_1398,N_14970,N_14898);
and UO_1399 (O_1399,N_14831,N_14981);
and UO_1400 (O_1400,N_14825,N_14903);
or UO_1401 (O_1401,N_14911,N_14960);
nand UO_1402 (O_1402,N_14935,N_14991);
xor UO_1403 (O_1403,N_14955,N_14820);
nand UO_1404 (O_1404,N_14987,N_14989);
xor UO_1405 (O_1405,N_14987,N_14974);
nand UO_1406 (O_1406,N_14960,N_14902);
or UO_1407 (O_1407,N_14908,N_14878);
xnor UO_1408 (O_1408,N_14802,N_14910);
nor UO_1409 (O_1409,N_14841,N_14886);
nand UO_1410 (O_1410,N_14976,N_14865);
xnor UO_1411 (O_1411,N_14884,N_14870);
or UO_1412 (O_1412,N_14820,N_14993);
and UO_1413 (O_1413,N_14800,N_14829);
or UO_1414 (O_1414,N_14866,N_14988);
nor UO_1415 (O_1415,N_14902,N_14891);
nand UO_1416 (O_1416,N_14847,N_14823);
or UO_1417 (O_1417,N_14803,N_14882);
or UO_1418 (O_1418,N_14916,N_14804);
and UO_1419 (O_1419,N_14887,N_14829);
nor UO_1420 (O_1420,N_14885,N_14906);
nand UO_1421 (O_1421,N_14858,N_14973);
and UO_1422 (O_1422,N_14815,N_14875);
or UO_1423 (O_1423,N_14899,N_14904);
nor UO_1424 (O_1424,N_14955,N_14964);
nand UO_1425 (O_1425,N_14821,N_14911);
or UO_1426 (O_1426,N_14878,N_14840);
and UO_1427 (O_1427,N_14843,N_14831);
or UO_1428 (O_1428,N_14946,N_14870);
nor UO_1429 (O_1429,N_14849,N_14995);
nand UO_1430 (O_1430,N_14864,N_14916);
nor UO_1431 (O_1431,N_14940,N_14867);
or UO_1432 (O_1432,N_14812,N_14945);
nand UO_1433 (O_1433,N_14955,N_14973);
xnor UO_1434 (O_1434,N_14922,N_14943);
xnor UO_1435 (O_1435,N_14938,N_14854);
xnor UO_1436 (O_1436,N_14959,N_14902);
nor UO_1437 (O_1437,N_14892,N_14851);
nand UO_1438 (O_1438,N_14940,N_14840);
nand UO_1439 (O_1439,N_14942,N_14973);
and UO_1440 (O_1440,N_14922,N_14959);
nand UO_1441 (O_1441,N_14915,N_14980);
nor UO_1442 (O_1442,N_14936,N_14998);
or UO_1443 (O_1443,N_14804,N_14803);
or UO_1444 (O_1444,N_14806,N_14894);
nand UO_1445 (O_1445,N_14922,N_14979);
or UO_1446 (O_1446,N_14952,N_14919);
and UO_1447 (O_1447,N_14836,N_14880);
nor UO_1448 (O_1448,N_14831,N_14956);
xnor UO_1449 (O_1449,N_14834,N_14906);
and UO_1450 (O_1450,N_14953,N_14949);
nor UO_1451 (O_1451,N_14903,N_14868);
nand UO_1452 (O_1452,N_14929,N_14995);
xor UO_1453 (O_1453,N_14898,N_14931);
nand UO_1454 (O_1454,N_14982,N_14951);
and UO_1455 (O_1455,N_14912,N_14934);
nor UO_1456 (O_1456,N_14960,N_14981);
xor UO_1457 (O_1457,N_14829,N_14901);
or UO_1458 (O_1458,N_14845,N_14950);
nand UO_1459 (O_1459,N_14919,N_14826);
and UO_1460 (O_1460,N_14852,N_14921);
nand UO_1461 (O_1461,N_14870,N_14881);
xnor UO_1462 (O_1462,N_14888,N_14949);
nor UO_1463 (O_1463,N_14810,N_14980);
or UO_1464 (O_1464,N_14887,N_14986);
nor UO_1465 (O_1465,N_14832,N_14903);
nor UO_1466 (O_1466,N_14861,N_14852);
nand UO_1467 (O_1467,N_14975,N_14860);
nor UO_1468 (O_1468,N_14892,N_14924);
nor UO_1469 (O_1469,N_14980,N_14856);
nand UO_1470 (O_1470,N_14993,N_14870);
nor UO_1471 (O_1471,N_14810,N_14800);
nand UO_1472 (O_1472,N_14926,N_14870);
or UO_1473 (O_1473,N_14840,N_14814);
nor UO_1474 (O_1474,N_14816,N_14853);
xor UO_1475 (O_1475,N_14985,N_14952);
nand UO_1476 (O_1476,N_14805,N_14800);
nor UO_1477 (O_1477,N_14816,N_14857);
nand UO_1478 (O_1478,N_14971,N_14956);
and UO_1479 (O_1479,N_14825,N_14987);
nand UO_1480 (O_1480,N_14996,N_14864);
xnor UO_1481 (O_1481,N_14926,N_14821);
and UO_1482 (O_1482,N_14934,N_14864);
xor UO_1483 (O_1483,N_14954,N_14967);
nand UO_1484 (O_1484,N_14885,N_14936);
nand UO_1485 (O_1485,N_14805,N_14947);
and UO_1486 (O_1486,N_14999,N_14830);
and UO_1487 (O_1487,N_14964,N_14951);
xor UO_1488 (O_1488,N_14986,N_14982);
and UO_1489 (O_1489,N_14917,N_14821);
xnor UO_1490 (O_1490,N_14913,N_14977);
xnor UO_1491 (O_1491,N_14966,N_14985);
nor UO_1492 (O_1492,N_14828,N_14943);
xor UO_1493 (O_1493,N_14863,N_14919);
or UO_1494 (O_1494,N_14863,N_14951);
nor UO_1495 (O_1495,N_14835,N_14834);
and UO_1496 (O_1496,N_14877,N_14916);
or UO_1497 (O_1497,N_14870,N_14997);
or UO_1498 (O_1498,N_14808,N_14921);
nor UO_1499 (O_1499,N_14848,N_14834);
nand UO_1500 (O_1500,N_14985,N_14911);
and UO_1501 (O_1501,N_14879,N_14897);
nor UO_1502 (O_1502,N_14899,N_14826);
and UO_1503 (O_1503,N_14961,N_14986);
nand UO_1504 (O_1504,N_14924,N_14872);
nand UO_1505 (O_1505,N_14985,N_14909);
xor UO_1506 (O_1506,N_14846,N_14902);
or UO_1507 (O_1507,N_14947,N_14847);
nor UO_1508 (O_1508,N_14937,N_14859);
xnor UO_1509 (O_1509,N_14996,N_14877);
or UO_1510 (O_1510,N_14894,N_14820);
xor UO_1511 (O_1511,N_14804,N_14954);
xor UO_1512 (O_1512,N_14825,N_14978);
nand UO_1513 (O_1513,N_14950,N_14986);
xor UO_1514 (O_1514,N_14978,N_14850);
nand UO_1515 (O_1515,N_14995,N_14833);
nand UO_1516 (O_1516,N_14879,N_14817);
nor UO_1517 (O_1517,N_14893,N_14891);
nand UO_1518 (O_1518,N_14879,N_14924);
xnor UO_1519 (O_1519,N_14945,N_14880);
and UO_1520 (O_1520,N_14895,N_14900);
nand UO_1521 (O_1521,N_14805,N_14847);
or UO_1522 (O_1522,N_14888,N_14985);
xor UO_1523 (O_1523,N_14980,N_14977);
and UO_1524 (O_1524,N_14979,N_14944);
nand UO_1525 (O_1525,N_14919,N_14828);
nor UO_1526 (O_1526,N_14957,N_14938);
or UO_1527 (O_1527,N_14801,N_14951);
xnor UO_1528 (O_1528,N_14821,N_14912);
nor UO_1529 (O_1529,N_14982,N_14839);
xnor UO_1530 (O_1530,N_14838,N_14979);
nor UO_1531 (O_1531,N_14850,N_14842);
xor UO_1532 (O_1532,N_14916,N_14949);
or UO_1533 (O_1533,N_14882,N_14829);
or UO_1534 (O_1534,N_14877,N_14800);
nor UO_1535 (O_1535,N_14999,N_14815);
nand UO_1536 (O_1536,N_14987,N_14820);
or UO_1537 (O_1537,N_14802,N_14932);
or UO_1538 (O_1538,N_14857,N_14997);
xor UO_1539 (O_1539,N_14823,N_14838);
nor UO_1540 (O_1540,N_14854,N_14821);
and UO_1541 (O_1541,N_14920,N_14850);
nand UO_1542 (O_1542,N_14993,N_14837);
nand UO_1543 (O_1543,N_14812,N_14934);
xor UO_1544 (O_1544,N_14922,N_14848);
or UO_1545 (O_1545,N_14975,N_14937);
nand UO_1546 (O_1546,N_14901,N_14956);
xor UO_1547 (O_1547,N_14883,N_14845);
xnor UO_1548 (O_1548,N_14849,N_14960);
or UO_1549 (O_1549,N_14922,N_14950);
xnor UO_1550 (O_1550,N_14937,N_14984);
and UO_1551 (O_1551,N_14984,N_14968);
nor UO_1552 (O_1552,N_14936,N_14803);
nand UO_1553 (O_1553,N_14806,N_14808);
nand UO_1554 (O_1554,N_14985,N_14975);
nor UO_1555 (O_1555,N_14990,N_14866);
nor UO_1556 (O_1556,N_14978,N_14931);
or UO_1557 (O_1557,N_14918,N_14984);
nand UO_1558 (O_1558,N_14810,N_14844);
and UO_1559 (O_1559,N_14907,N_14931);
xor UO_1560 (O_1560,N_14844,N_14842);
or UO_1561 (O_1561,N_14893,N_14910);
or UO_1562 (O_1562,N_14994,N_14965);
nand UO_1563 (O_1563,N_14864,N_14821);
and UO_1564 (O_1564,N_14986,N_14895);
or UO_1565 (O_1565,N_14816,N_14871);
nor UO_1566 (O_1566,N_14935,N_14910);
nand UO_1567 (O_1567,N_14843,N_14811);
and UO_1568 (O_1568,N_14979,N_14945);
nand UO_1569 (O_1569,N_14887,N_14909);
nor UO_1570 (O_1570,N_14944,N_14829);
or UO_1571 (O_1571,N_14960,N_14985);
nand UO_1572 (O_1572,N_14884,N_14971);
or UO_1573 (O_1573,N_14985,N_14897);
nand UO_1574 (O_1574,N_14855,N_14890);
and UO_1575 (O_1575,N_14987,N_14919);
nand UO_1576 (O_1576,N_14802,N_14820);
and UO_1577 (O_1577,N_14870,N_14843);
nand UO_1578 (O_1578,N_14893,N_14947);
or UO_1579 (O_1579,N_14858,N_14903);
nor UO_1580 (O_1580,N_14856,N_14894);
xnor UO_1581 (O_1581,N_14825,N_14901);
and UO_1582 (O_1582,N_14930,N_14840);
or UO_1583 (O_1583,N_14837,N_14910);
and UO_1584 (O_1584,N_14988,N_14870);
or UO_1585 (O_1585,N_14927,N_14831);
xnor UO_1586 (O_1586,N_14826,N_14894);
or UO_1587 (O_1587,N_14998,N_14825);
and UO_1588 (O_1588,N_14889,N_14890);
or UO_1589 (O_1589,N_14929,N_14925);
and UO_1590 (O_1590,N_14847,N_14843);
and UO_1591 (O_1591,N_14941,N_14911);
nor UO_1592 (O_1592,N_14884,N_14879);
or UO_1593 (O_1593,N_14902,N_14827);
xor UO_1594 (O_1594,N_14992,N_14943);
or UO_1595 (O_1595,N_14933,N_14848);
and UO_1596 (O_1596,N_14807,N_14851);
or UO_1597 (O_1597,N_14891,N_14935);
or UO_1598 (O_1598,N_14920,N_14961);
and UO_1599 (O_1599,N_14849,N_14954);
nor UO_1600 (O_1600,N_14896,N_14883);
nand UO_1601 (O_1601,N_14950,N_14915);
nand UO_1602 (O_1602,N_14902,N_14899);
nor UO_1603 (O_1603,N_14996,N_14860);
nand UO_1604 (O_1604,N_14821,N_14918);
or UO_1605 (O_1605,N_14842,N_14925);
or UO_1606 (O_1606,N_14956,N_14826);
and UO_1607 (O_1607,N_14922,N_14859);
nand UO_1608 (O_1608,N_14978,N_14809);
nor UO_1609 (O_1609,N_14837,N_14867);
and UO_1610 (O_1610,N_14989,N_14886);
xnor UO_1611 (O_1611,N_14941,N_14982);
xnor UO_1612 (O_1612,N_14830,N_14849);
and UO_1613 (O_1613,N_14911,N_14803);
nor UO_1614 (O_1614,N_14967,N_14886);
xnor UO_1615 (O_1615,N_14840,N_14901);
nand UO_1616 (O_1616,N_14936,N_14916);
and UO_1617 (O_1617,N_14930,N_14853);
or UO_1618 (O_1618,N_14966,N_14837);
and UO_1619 (O_1619,N_14956,N_14852);
or UO_1620 (O_1620,N_14915,N_14873);
nor UO_1621 (O_1621,N_14829,N_14912);
nor UO_1622 (O_1622,N_14968,N_14995);
or UO_1623 (O_1623,N_14850,N_14905);
and UO_1624 (O_1624,N_14953,N_14842);
and UO_1625 (O_1625,N_14897,N_14803);
and UO_1626 (O_1626,N_14999,N_14832);
and UO_1627 (O_1627,N_14827,N_14926);
or UO_1628 (O_1628,N_14970,N_14832);
and UO_1629 (O_1629,N_14988,N_14855);
xnor UO_1630 (O_1630,N_14921,N_14896);
nor UO_1631 (O_1631,N_14869,N_14990);
and UO_1632 (O_1632,N_14936,N_14813);
or UO_1633 (O_1633,N_14828,N_14917);
or UO_1634 (O_1634,N_14900,N_14937);
nand UO_1635 (O_1635,N_14880,N_14814);
nand UO_1636 (O_1636,N_14960,N_14871);
or UO_1637 (O_1637,N_14907,N_14917);
nor UO_1638 (O_1638,N_14966,N_14916);
nand UO_1639 (O_1639,N_14857,N_14814);
xor UO_1640 (O_1640,N_14829,N_14979);
or UO_1641 (O_1641,N_14924,N_14928);
nor UO_1642 (O_1642,N_14908,N_14983);
nor UO_1643 (O_1643,N_14877,N_14807);
xor UO_1644 (O_1644,N_14898,N_14801);
and UO_1645 (O_1645,N_14986,N_14970);
and UO_1646 (O_1646,N_14961,N_14957);
nor UO_1647 (O_1647,N_14976,N_14993);
nand UO_1648 (O_1648,N_14857,N_14827);
xor UO_1649 (O_1649,N_14939,N_14992);
or UO_1650 (O_1650,N_14856,N_14982);
nand UO_1651 (O_1651,N_14988,N_14897);
or UO_1652 (O_1652,N_14892,N_14804);
xor UO_1653 (O_1653,N_14998,N_14911);
or UO_1654 (O_1654,N_14823,N_14978);
xnor UO_1655 (O_1655,N_14829,N_14924);
nor UO_1656 (O_1656,N_14962,N_14970);
nor UO_1657 (O_1657,N_14897,N_14946);
nand UO_1658 (O_1658,N_14997,N_14939);
nand UO_1659 (O_1659,N_14827,N_14938);
nor UO_1660 (O_1660,N_14854,N_14930);
nor UO_1661 (O_1661,N_14845,N_14908);
nor UO_1662 (O_1662,N_14834,N_14929);
nand UO_1663 (O_1663,N_14906,N_14940);
and UO_1664 (O_1664,N_14904,N_14984);
nand UO_1665 (O_1665,N_14928,N_14875);
nand UO_1666 (O_1666,N_14999,N_14896);
or UO_1667 (O_1667,N_14967,N_14962);
xnor UO_1668 (O_1668,N_14943,N_14870);
nor UO_1669 (O_1669,N_14934,N_14832);
and UO_1670 (O_1670,N_14971,N_14834);
nand UO_1671 (O_1671,N_14827,N_14989);
or UO_1672 (O_1672,N_14915,N_14890);
and UO_1673 (O_1673,N_14924,N_14989);
and UO_1674 (O_1674,N_14940,N_14999);
and UO_1675 (O_1675,N_14806,N_14888);
or UO_1676 (O_1676,N_14938,N_14989);
or UO_1677 (O_1677,N_14854,N_14931);
xnor UO_1678 (O_1678,N_14853,N_14929);
or UO_1679 (O_1679,N_14954,N_14902);
or UO_1680 (O_1680,N_14803,N_14966);
nand UO_1681 (O_1681,N_14998,N_14934);
nor UO_1682 (O_1682,N_14866,N_14938);
and UO_1683 (O_1683,N_14925,N_14963);
xor UO_1684 (O_1684,N_14837,N_14967);
nor UO_1685 (O_1685,N_14925,N_14823);
and UO_1686 (O_1686,N_14940,N_14805);
or UO_1687 (O_1687,N_14808,N_14815);
nand UO_1688 (O_1688,N_14801,N_14883);
or UO_1689 (O_1689,N_14852,N_14941);
xnor UO_1690 (O_1690,N_14946,N_14880);
or UO_1691 (O_1691,N_14847,N_14968);
nor UO_1692 (O_1692,N_14991,N_14890);
nand UO_1693 (O_1693,N_14938,N_14972);
nand UO_1694 (O_1694,N_14936,N_14888);
nor UO_1695 (O_1695,N_14847,N_14926);
or UO_1696 (O_1696,N_14926,N_14935);
or UO_1697 (O_1697,N_14975,N_14819);
xor UO_1698 (O_1698,N_14817,N_14847);
nand UO_1699 (O_1699,N_14953,N_14833);
and UO_1700 (O_1700,N_14874,N_14977);
nand UO_1701 (O_1701,N_14978,N_14879);
nor UO_1702 (O_1702,N_14994,N_14897);
nor UO_1703 (O_1703,N_14955,N_14975);
nor UO_1704 (O_1704,N_14852,N_14886);
xnor UO_1705 (O_1705,N_14848,N_14931);
nand UO_1706 (O_1706,N_14968,N_14954);
and UO_1707 (O_1707,N_14893,N_14846);
xor UO_1708 (O_1708,N_14949,N_14952);
and UO_1709 (O_1709,N_14974,N_14994);
and UO_1710 (O_1710,N_14951,N_14861);
xnor UO_1711 (O_1711,N_14969,N_14947);
nand UO_1712 (O_1712,N_14949,N_14984);
nand UO_1713 (O_1713,N_14903,N_14886);
and UO_1714 (O_1714,N_14815,N_14991);
xnor UO_1715 (O_1715,N_14973,N_14815);
xor UO_1716 (O_1716,N_14807,N_14876);
or UO_1717 (O_1717,N_14951,N_14879);
or UO_1718 (O_1718,N_14951,N_14935);
nor UO_1719 (O_1719,N_14944,N_14898);
nor UO_1720 (O_1720,N_14813,N_14853);
xor UO_1721 (O_1721,N_14844,N_14922);
xor UO_1722 (O_1722,N_14904,N_14918);
and UO_1723 (O_1723,N_14939,N_14816);
nor UO_1724 (O_1724,N_14835,N_14802);
nor UO_1725 (O_1725,N_14803,N_14991);
and UO_1726 (O_1726,N_14846,N_14843);
and UO_1727 (O_1727,N_14879,N_14853);
nor UO_1728 (O_1728,N_14907,N_14977);
xor UO_1729 (O_1729,N_14872,N_14993);
or UO_1730 (O_1730,N_14978,N_14862);
nand UO_1731 (O_1731,N_14970,N_14860);
and UO_1732 (O_1732,N_14863,N_14976);
nor UO_1733 (O_1733,N_14987,N_14946);
nand UO_1734 (O_1734,N_14975,N_14850);
nand UO_1735 (O_1735,N_14952,N_14871);
nand UO_1736 (O_1736,N_14819,N_14857);
nor UO_1737 (O_1737,N_14812,N_14966);
nor UO_1738 (O_1738,N_14912,N_14881);
and UO_1739 (O_1739,N_14965,N_14903);
nor UO_1740 (O_1740,N_14876,N_14986);
and UO_1741 (O_1741,N_14878,N_14895);
or UO_1742 (O_1742,N_14862,N_14827);
xor UO_1743 (O_1743,N_14831,N_14859);
nand UO_1744 (O_1744,N_14935,N_14965);
xnor UO_1745 (O_1745,N_14842,N_14993);
xor UO_1746 (O_1746,N_14918,N_14815);
xor UO_1747 (O_1747,N_14816,N_14835);
and UO_1748 (O_1748,N_14837,N_14812);
xor UO_1749 (O_1749,N_14900,N_14860);
xnor UO_1750 (O_1750,N_14918,N_14971);
or UO_1751 (O_1751,N_14882,N_14895);
nor UO_1752 (O_1752,N_14888,N_14981);
nand UO_1753 (O_1753,N_14994,N_14997);
xor UO_1754 (O_1754,N_14935,N_14918);
nor UO_1755 (O_1755,N_14853,N_14901);
and UO_1756 (O_1756,N_14890,N_14907);
or UO_1757 (O_1757,N_14826,N_14885);
or UO_1758 (O_1758,N_14871,N_14912);
nor UO_1759 (O_1759,N_14890,N_14950);
or UO_1760 (O_1760,N_14822,N_14863);
or UO_1761 (O_1761,N_14819,N_14856);
nand UO_1762 (O_1762,N_14825,N_14805);
and UO_1763 (O_1763,N_14990,N_14964);
or UO_1764 (O_1764,N_14885,N_14957);
or UO_1765 (O_1765,N_14870,N_14933);
or UO_1766 (O_1766,N_14896,N_14857);
nand UO_1767 (O_1767,N_14856,N_14942);
and UO_1768 (O_1768,N_14887,N_14973);
xnor UO_1769 (O_1769,N_14859,N_14934);
xnor UO_1770 (O_1770,N_14929,N_14922);
nor UO_1771 (O_1771,N_14893,N_14976);
and UO_1772 (O_1772,N_14908,N_14984);
and UO_1773 (O_1773,N_14817,N_14841);
or UO_1774 (O_1774,N_14999,N_14973);
nand UO_1775 (O_1775,N_14964,N_14993);
xor UO_1776 (O_1776,N_14831,N_14800);
nand UO_1777 (O_1777,N_14953,N_14897);
and UO_1778 (O_1778,N_14891,N_14818);
nor UO_1779 (O_1779,N_14948,N_14967);
or UO_1780 (O_1780,N_14933,N_14962);
nor UO_1781 (O_1781,N_14933,N_14810);
and UO_1782 (O_1782,N_14972,N_14948);
nor UO_1783 (O_1783,N_14904,N_14896);
or UO_1784 (O_1784,N_14957,N_14869);
xor UO_1785 (O_1785,N_14901,N_14850);
and UO_1786 (O_1786,N_14846,N_14964);
and UO_1787 (O_1787,N_14983,N_14950);
and UO_1788 (O_1788,N_14960,N_14984);
or UO_1789 (O_1789,N_14889,N_14831);
or UO_1790 (O_1790,N_14884,N_14845);
and UO_1791 (O_1791,N_14885,N_14897);
and UO_1792 (O_1792,N_14813,N_14982);
nand UO_1793 (O_1793,N_14843,N_14920);
nand UO_1794 (O_1794,N_14982,N_14873);
nor UO_1795 (O_1795,N_14891,N_14961);
or UO_1796 (O_1796,N_14917,N_14830);
nand UO_1797 (O_1797,N_14983,N_14915);
nor UO_1798 (O_1798,N_14906,N_14997);
xor UO_1799 (O_1799,N_14987,N_14870);
xor UO_1800 (O_1800,N_14906,N_14970);
nor UO_1801 (O_1801,N_14879,N_14816);
xor UO_1802 (O_1802,N_14916,N_14986);
nor UO_1803 (O_1803,N_14929,N_14842);
and UO_1804 (O_1804,N_14919,N_14902);
xnor UO_1805 (O_1805,N_14804,N_14953);
nor UO_1806 (O_1806,N_14803,N_14909);
or UO_1807 (O_1807,N_14894,N_14825);
nand UO_1808 (O_1808,N_14998,N_14842);
nand UO_1809 (O_1809,N_14953,N_14895);
xnor UO_1810 (O_1810,N_14806,N_14819);
nand UO_1811 (O_1811,N_14890,N_14921);
nor UO_1812 (O_1812,N_14820,N_14863);
and UO_1813 (O_1813,N_14978,N_14842);
or UO_1814 (O_1814,N_14849,N_14949);
and UO_1815 (O_1815,N_14860,N_14890);
and UO_1816 (O_1816,N_14970,N_14950);
nor UO_1817 (O_1817,N_14979,N_14856);
xor UO_1818 (O_1818,N_14918,N_14827);
nor UO_1819 (O_1819,N_14997,N_14920);
or UO_1820 (O_1820,N_14877,N_14817);
nand UO_1821 (O_1821,N_14972,N_14995);
nand UO_1822 (O_1822,N_14869,N_14902);
or UO_1823 (O_1823,N_14859,N_14806);
nor UO_1824 (O_1824,N_14937,N_14874);
or UO_1825 (O_1825,N_14885,N_14841);
nand UO_1826 (O_1826,N_14842,N_14811);
nand UO_1827 (O_1827,N_14979,N_14996);
and UO_1828 (O_1828,N_14974,N_14962);
nand UO_1829 (O_1829,N_14965,N_14806);
or UO_1830 (O_1830,N_14988,N_14862);
xnor UO_1831 (O_1831,N_14886,N_14890);
or UO_1832 (O_1832,N_14920,N_14995);
nor UO_1833 (O_1833,N_14939,N_14911);
or UO_1834 (O_1834,N_14928,N_14914);
or UO_1835 (O_1835,N_14914,N_14916);
nand UO_1836 (O_1836,N_14930,N_14979);
and UO_1837 (O_1837,N_14902,N_14938);
or UO_1838 (O_1838,N_14920,N_14852);
or UO_1839 (O_1839,N_14837,N_14897);
and UO_1840 (O_1840,N_14972,N_14906);
nand UO_1841 (O_1841,N_14972,N_14921);
nor UO_1842 (O_1842,N_14859,N_14882);
nor UO_1843 (O_1843,N_14929,N_14811);
or UO_1844 (O_1844,N_14908,N_14927);
or UO_1845 (O_1845,N_14819,N_14902);
or UO_1846 (O_1846,N_14888,N_14959);
or UO_1847 (O_1847,N_14817,N_14829);
xnor UO_1848 (O_1848,N_14827,N_14836);
and UO_1849 (O_1849,N_14811,N_14812);
xnor UO_1850 (O_1850,N_14960,N_14892);
xnor UO_1851 (O_1851,N_14851,N_14823);
or UO_1852 (O_1852,N_14865,N_14827);
nand UO_1853 (O_1853,N_14997,N_14818);
or UO_1854 (O_1854,N_14878,N_14918);
and UO_1855 (O_1855,N_14812,N_14866);
and UO_1856 (O_1856,N_14860,N_14968);
or UO_1857 (O_1857,N_14980,N_14821);
nor UO_1858 (O_1858,N_14887,N_14981);
or UO_1859 (O_1859,N_14915,N_14842);
xor UO_1860 (O_1860,N_14820,N_14869);
nand UO_1861 (O_1861,N_14874,N_14966);
or UO_1862 (O_1862,N_14927,N_14948);
or UO_1863 (O_1863,N_14851,N_14828);
and UO_1864 (O_1864,N_14973,N_14982);
nand UO_1865 (O_1865,N_14921,N_14855);
and UO_1866 (O_1866,N_14917,N_14972);
nor UO_1867 (O_1867,N_14907,N_14952);
or UO_1868 (O_1868,N_14813,N_14909);
and UO_1869 (O_1869,N_14896,N_14828);
and UO_1870 (O_1870,N_14859,N_14974);
and UO_1871 (O_1871,N_14967,N_14807);
xor UO_1872 (O_1872,N_14808,N_14830);
and UO_1873 (O_1873,N_14992,N_14832);
or UO_1874 (O_1874,N_14962,N_14883);
or UO_1875 (O_1875,N_14881,N_14854);
or UO_1876 (O_1876,N_14835,N_14973);
xor UO_1877 (O_1877,N_14966,N_14813);
xor UO_1878 (O_1878,N_14979,N_14850);
nor UO_1879 (O_1879,N_14908,N_14805);
xor UO_1880 (O_1880,N_14884,N_14963);
nand UO_1881 (O_1881,N_14865,N_14905);
nor UO_1882 (O_1882,N_14875,N_14906);
and UO_1883 (O_1883,N_14990,N_14950);
nor UO_1884 (O_1884,N_14913,N_14936);
or UO_1885 (O_1885,N_14950,N_14869);
nand UO_1886 (O_1886,N_14954,N_14959);
or UO_1887 (O_1887,N_14836,N_14912);
nand UO_1888 (O_1888,N_14830,N_14936);
nand UO_1889 (O_1889,N_14840,N_14953);
nand UO_1890 (O_1890,N_14813,N_14933);
nor UO_1891 (O_1891,N_14950,N_14994);
nor UO_1892 (O_1892,N_14816,N_14936);
xor UO_1893 (O_1893,N_14971,N_14852);
nor UO_1894 (O_1894,N_14936,N_14832);
or UO_1895 (O_1895,N_14953,N_14810);
nand UO_1896 (O_1896,N_14994,N_14976);
nand UO_1897 (O_1897,N_14873,N_14836);
or UO_1898 (O_1898,N_14814,N_14850);
xor UO_1899 (O_1899,N_14956,N_14815);
and UO_1900 (O_1900,N_14914,N_14818);
xnor UO_1901 (O_1901,N_14922,N_14805);
and UO_1902 (O_1902,N_14998,N_14864);
nand UO_1903 (O_1903,N_14967,N_14989);
and UO_1904 (O_1904,N_14877,N_14880);
or UO_1905 (O_1905,N_14940,N_14838);
or UO_1906 (O_1906,N_14945,N_14942);
and UO_1907 (O_1907,N_14870,N_14891);
nand UO_1908 (O_1908,N_14960,N_14983);
and UO_1909 (O_1909,N_14835,N_14996);
and UO_1910 (O_1910,N_14805,N_14974);
nand UO_1911 (O_1911,N_14817,N_14894);
nand UO_1912 (O_1912,N_14803,N_14834);
nand UO_1913 (O_1913,N_14973,N_14940);
or UO_1914 (O_1914,N_14964,N_14963);
nor UO_1915 (O_1915,N_14938,N_14941);
nand UO_1916 (O_1916,N_14959,N_14989);
nand UO_1917 (O_1917,N_14894,N_14985);
and UO_1918 (O_1918,N_14844,N_14925);
or UO_1919 (O_1919,N_14835,N_14959);
and UO_1920 (O_1920,N_14904,N_14859);
xnor UO_1921 (O_1921,N_14906,N_14822);
or UO_1922 (O_1922,N_14966,N_14902);
nor UO_1923 (O_1923,N_14965,N_14923);
xnor UO_1924 (O_1924,N_14954,N_14983);
or UO_1925 (O_1925,N_14881,N_14943);
nand UO_1926 (O_1926,N_14823,N_14876);
and UO_1927 (O_1927,N_14846,N_14925);
and UO_1928 (O_1928,N_14979,N_14990);
nor UO_1929 (O_1929,N_14984,N_14848);
nor UO_1930 (O_1930,N_14960,N_14953);
nor UO_1931 (O_1931,N_14928,N_14811);
or UO_1932 (O_1932,N_14931,N_14942);
and UO_1933 (O_1933,N_14879,N_14856);
nor UO_1934 (O_1934,N_14916,N_14808);
and UO_1935 (O_1935,N_14951,N_14983);
or UO_1936 (O_1936,N_14882,N_14807);
and UO_1937 (O_1937,N_14946,N_14948);
xnor UO_1938 (O_1938,N_14916,N_14883);
xnor UO_1939 (O_1939,N_14958,N_14932);
nor UO_1940 (O_1940,N_14905,N_14880);
nand UO_1941 (O_1941,N_14971,N_14833);
or UO_1942 (O_1942,N_14841,N_14954);
or UO_1943 (O_1943,N_14895,N_14885);
nand UO_1944 (O_1944,N_14871,N_14881);
nor UO_1945 (O_1945,N_14959,N_14859);
or UO_1946 (O_1946,N_14835,N_14839);
or UO_1947 (O_1947,N_14970,N_14817);
xnor UO_1948 (O_1948,N_14917,N_14859);
and UO_1949 (O_1949,N_14982,N_14961);
nand UO_1950 (O_1950,N_14963,N_14942);
or UO_1951 (O_1951,N_14929,N_14900);
or UO_1952 (O_1952,N_14898,N_14911);
or UO_1953 (O_1953,N_14997,N_14947);
and UO_1954 (O_1954,N_14983,N_14977);
nand UO_1955 (O_1955,N_14879,N_14850);
xor UO_1956 (O_1956,N_14954,N_14886);
and UO_1957 (O_1957,N_14978,N_14917);
or UO_1958 (O_1958,N_14848,N_14805);
nand UO_1959 (O_1959,N_14867,N_14970);
nand UO_1960 (O_1960,N_14947,N_14800);
nand UO_1961 (O_1961,N_14938,N_14872);
nor UO_1962 (O_1962,N_14992,N_14969);
xnor UO_1963 (O_1963,N_14985,N_14963);
or UO_1964 (O_1964,N_14835,N_14991);
and UO_1965 (O_1965,N_14978,N_14910);
and UO_1966 (O_1966,N_14901,N_14893);
nor UO_1967 (O_1967,N_14873,N_14994);
nand UO_1968 (O_1968,N_14806,N_14983);
and UO_1969 (O_1969,N_14843,N_14966);
or UO_1970 (O_1970,N_14882,N_14867);
and UO_1971 (O_1971,N_14807,N_14981);
xnor UO_1972 (O_1972,N_14929,N_14926);
and UO_1973 (O_1973,N_14971,N_14839);
and UO_1974 (O_1974,N_14861,N_14909);
and UO_1975 (O_1975,N_14916,N_14832);
and UO_1976 (O_1976,N_14886,N_14892);
nor UO_1977 (O_1977,N_14930,N_14829);
or UO_1978 (O_1978,N_14961,N_14838);
nand UO_1979 (O_1979,N_14853,N_14943);
xor UO_1980 (O_1980,N_14890,N_14964);
nor UO_1981 (O_1981,N_14996,N_14813);
and UO_1982 (O_1982,N_14963,N_14903);
xor UO_1983 (O_1983,N_14935,N_14928);
xor UO_1984 (O_1984,N_14945,N_14991);
nand UO_1985 (O_1985,N_14921,N_14800);
or UO_1986 (O_1986,N_14995,N_14882);
nor UO_1987 (O_1987,N_14814,N_14940);
nor UO_1988 (O_1988,N_14820,N_14946);
and UO_1989 (O_1989,N_14901,N_14846);
and UO_1990 (O_1990,N_14925,N_14812);
nor UO_1991 (O_1991,N_14960,N_14938);
xnor UO_1992 (O_1992,N_14932,N_14915);
nor UO_1993 (O_1993,N_14930,N_14939);
xnor UO_1994 (O_1994,N_14891,N_14871);
nor UO_1995 (O_1995,N_14916,N_14928);
or UO_1996 (O_1996,N_14843,N_14925);
xnor UO_1997 (O_1997,N_14825,N_14973);
or UO_1998 (O_1998,N_14976,N_14921);
and UO_1999 (O_1999,N_14894,N_14972);
endmodule