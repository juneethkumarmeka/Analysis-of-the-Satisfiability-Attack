module basic_750_5000_1000_5_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_85,In_555);
xnor U1 (N_1,In_118,In_523);
nor U2 (N_2,In_485,In_537);
nand U3 (N_3,In_551,In_27);
and U4 (N_4,In_449,In_512);
nand U5 (N_5,In_684,In_53);
nand U6 (N_6,In_114,In_8);
nor U7 (N_7,In_634,In_138);
nand U8 (N_8,In_58,In_683);
nand U9 (N_9,In_521,In_188);
or U10 (N_10,In_124,In_627);
xnor U11 (N_11,In_242,In_176);
and U12 (N_12,In_322,In_134);
nand U13 (N_13,In_214,In_606);
and U14 (N_14,In_246,In_365);
nand U15 (N_15,In_509,In_145);
nand U16 (N_16,In_552,In_12);
nor U17 (N_17,In_574,In_742);
nand U18 (N_18,In_143,In_724);
or U19 (N_19,In_387,In_557);
nor U20 (N_20,In_238,In_352);
xnor U21 (N_21,In_350,In_360);
or U22 (N_22,In_540,In_182);
and U23 (N_23,In_728,In_402);
and U24 (N_24,In_638,In_291);
and U25 (N_25,In_311,In_23);
and U26 (N_26,In_337,In_443);
nor U27 (N_27,In_177,In_63);
or U28 (N_28,In_279,In_416);
and U29 (N_29,In_426,In_155);
and U30 (N_30,In_692,In_91);
and U31 (N_31,In_423,In_111);
and U32 (N_32,In_212,In_483);
xor U33 (N_33,In_7,In_656);
and U34 (N_34,In_536,In_258);
or U35 (N_35,In_170,In_657);
or U36 (N_36,In_583,In_301);
nand U37 (N_37,In_206,In_378);
nand U38 (N_38,In_727,In_167);
xnor U39 (N_39,In_418,In_256);
and U40 (N_40,In_348,In_239);
and U41 (N_41,In_204,In_95);
nor U42 (N_42,In_486,In_590);
xnor U43 (N_43,In_132,In_399);
nor U44 (N_44,In_385,In_180);
nor U45 (N_45,In_667,In_500);
nand U46 (N_46,In_333,In_725);
or U47 (N_47,In_297,In_610);
nor U48 (N_48,In_151,In_202);
nand U49 (N_49,In_524,In_741);
or U50 (N_50,In_473,In_567);
nand U51 (N_51,In_603,In_144);
nor U52 (N_52,In_159,In_543);
nor U53 (N_53,In_332,In_288);
or U54 (N_54,In_459,In_183);
or U55 (N_55,In_193,In_45);
nand U56 (N_56,In_700,In_284);
or U57 (N_57,In_26,In_363);
and U58 (N_58,In_120,In_674);
or U59 (N_59,In_670,In_127);
and U60 (N_60,In_732,In_390);
and U61 (N_61,In_695,In_351);
or U62 (N_62,In_355,In_5);
xnor U63 (N_63,In_201,In_428);
nand U64 (N_64,In_326,In_442);
or U65 (N_65,In_141,In_130);
xnor U66 (N_66,In_382,In_222);
xor U67 (N_67,In_391,In_632);
nand U68 (N_68,In_717,In_266);
nand U69 (N_69,In_644,In_585);
or U70 (N_70,In_318,In_314);
nand U71 (N_71,In_469,In_296);
xnor U72 (N_72,In_715,In_317);
and U73 (N_73,In_3,In_298);
nor U74 (N_74,In_356,In_589);
nand U75 (N_75,In_331,In_735);
nand U76 (N_76,In_37,In_694);
xor U77 (N_77,In_146,In_662);
nand U78 (N_78,In_522,In_538);
nor U79 (N_79,In_56,In_542);
xor U80 (N_80,In_345,In_554);
nand U81 (N_81,In_6,In_75);
or U82 (N_82,In_18,In_397);
xnor U83 (N_83,In_566,In_497);
nand U84 (N_84,In_438,In_197);
xor U85 (N_85,In_461,In_172);
nand U86 (N_86,In_383,In_743);
or U87 (N_87,In_531,In_679);
nand U88 (N_88,In_471,In_584);
xnor U89 (N_89,In_731,In_546);
nor U90 (N_90,In_477,In_175);
or U91 (N_91,In_292,In_283);
or U92 (N_92,In_126,In_342);
nand U93 (N_93,In_109,In_139);
nand U94 (N_94,In_308,In_294);
or U95 (N_95,In_580,In_676);
or U96 (N_96,In_649,In_362);
nor U97 (N_97,In_441,In_166);
and U98 (N_98,In_709,In_270);
nor U99 (N_99,In_468,In_484);
nand U100 (N_100,In_336,In_346);
and U101 (N_101,In_65,In_226);
and U102 (N_102,In_429,In_516);
or U103 (N_103,In_2,In_456);
or U104 (N_104,In_431,In_185);
nor U105 (N_105,In_98,In_44);
or U106 (N_106,In_587,In_626);
nand U107 (N_107,In_687,In_257);
nor U108 (N_108,In_205,In_49);
nand U109 (N_109,In_324,In_406);
and U110 (N_110,In_330,In_450);
nand U111 (N_111,In_199,In_421);
or U112 (N_112,In_366,In_218);
xor U113 (N_113,In_614,In_154);
xnor U114 (N_114,In_248,In_510);
and U115 (N_115,In_492,In_217);
or U116 (N_116,In_152,In_161);
xor U117 (N_117,In_673,In_663);
and U118 (N_118,In_493,In_401);
and U119 (N_119,In_83,In_511);
nor U120 (N_120,In_94,In_179);
nor U121 (N_121,In_577,In_310);
or U122 (N_122,In_235,In_252);
and U123 (N_123,In_344,In_19);
nand U124 (N_124,In_737,In_300);
nand U125 (N_125,In_739,In_255);
or U126 (N_126,In_268,In_71);
or U127 (N_127,In_274,In_160);
nor U128 (N_128,In_282,In_530);
or U129 (N_129,In_495,In_488);
nor U130 (N_130,In_104,In_89);
or U131 (N_131,In_653,In_110);
and U132 (N_132,In_572,In_13);
or U133 (N_133,In_384,In_379);
or U134 (N_134,In_678,In_746);
nand U135 (N_135,In_55,In_377);
and U136 (N_136,In_93,In_73);
and U137 (N_137,In_631,In_341);
nor U138 (N_138,In_20,In_620);
nand U139 (N_139,In_101,In_404);
and U140 (N_140,In_487,In_68);
nor U141 (N_141,In_278,In_494);
and U142 (N_142,In_221,In_602);
nor U143 (N_143,In_745,In_502);
or U144 (N_144,In_565,In_398);
nor U145 (N_145,In_164,In_86);
and U146 (N_146,In_328,In_321);
and U147 (N_147,In_628,In_564);
nor U148 (N_148,In_329,In_665);
xnor U149 (N_149,In_437,In_581);
or U150 (N_150,In_479,In_714);
nor U151 (N_151,In_439,In_419);
nand U152 (N_152,In_169,In_153);
and U153 (N_153,In_570,In_573);
and U154 (N_154,In_107,In_425);
and U155 (N_155,In_61,In_386);
nor U156 (N_156,In_190,In_150);
and U157 (N_157,In_79,In_525);
or U158 (N_158,In_604,In_251);
nand U159 (N_159,In_70,In_67);
nor U160 (N_160,In_43,In_633);
nor U161 (N_161,In_254,In_607);
nor U162 (N_162,In_738,In_220);
and U163 (N_163,In_413,In_643);
nand U164 (N_164,In_417,In_508);
nand U165 (N_165,In_749,In_121);
nand U166 (N_166,In_722,In_102);
xnor U167 (N_167,In_637,In_88);
and U168 (N_168,In_527,In_22);
nor U169 (N_169,In_498,In_302);
nor U170 (N_170,In_376,In_553);
nor U171 (N_171,In_624,In_596);
and U172 (N_172,In_207,In_669);
or U173 (N_173,In_307,In_135);
xor U174 (N_174,In_285,In_327);
or U175 (N_175,In_748,In_690);
or U176 (N_176,In_476,In_373);
or U177 (N_177,In_9,In_358);
and U178 (N_178,In_629,In_81);
nand U179 (N_179,In_299,In_131);
xor U180 (N_180,In_592,In_460);
nand U181 (N_181,In_635,In_48);
nor U182 (N_182,In_113,In_710);
nor U183 (N_183,In_287,In_211);
or U184 (N_184,In_505,In_375);
or U185 (N_185,In_103,In_82);
or U186 (N_186,In_519,In_74);
nor U187 (N_187,In_489,In_414);
nand U188 (N_188,In_575,In_616);
and U189 (N_189,In_10,In_173);
nor U190 (N_190,In_474,In_200);
nor U191 (N_191,In_77,In_457);
or U192 (N_192,In_579,In_517);
nand U193 (N_193,In_29,In_306);
or U194 (N_194,In_196,In_452);
nor U195 (N_195,In_440,In_165);
nand U196 (N_196,In_210,In_528);
nand U197 (N_197,In_148,In_122);
and U198 (N_198,In_681,In_475);
nand U199 (N_199,In_303,In_253);
and U200 (N_200,In_707,In_586);
xor U201 (N_201,In_666,In_506);
and U202 (N_202,In_137,In_289);
and U203 (N_203,In_16,In_427);
nor U204 (N_204,In_280,In_216);
and U205 (N_205,In_593,In_393);
or U206 (N_206,In_482,In_123);
nand U207 (N_207,In_591,In_41);
nor U208 (N_208,In_69,In_194);
or U209 (N_209,In_462,In_617);
and U210 (N_210,In_233,In_231);
and U211 (N_211,In_520,In_719);
nand U212 (N_212,In_576,In_466);
and U213 (N_213,In_50,In_272);
and U214 (N_214,In_338,In_650);
and U215 (N_215,In_1,In_711);
or U216 (N_216,In_99,In_335);
and U217 (N_217,In_403,In_689);
nor U218 (N_218,In_90,In_685);
nor U219 (N_219,In_38,In_225);
nand U220 (N_220,In_415,In_693);
and U221 (N_221,In_312,In_87);
and U222 (N_222,In_313,In_168);
or U223 (N_223,In_436,In_136);
xor U224 (N_224,In_25,In_184);
and U225 (N_225,In_533,In_4);
nand U226 (N_226,In_556,In_304);
and U227 (N_227,In_504,In_192);
nor U228 (N_228,In_605,In_247);
nor U229 (N_229,In_513,In_52);
xnor U230 (N_230,In_716,In_733);
nand U231 (N_231,In_47,In_582);
xnor U232 (N_232,In_680,In_388);
or U233 (N_233,In_286,In_405);
nand U234 (N_234,In_187,In_347);
nor U235 (N_235,In_259,In_66);
nor U236 (N_236,In_648,In_721);
xor U237 (N_237,In_92,In_219);
and U238 (N_238,In_59,In_671);
xor U239 (N_239,In_0,In_613);
nand U240 (N_240,In_729,In_407);
and U241 (N_241,In_290,In_677);
xnor U242 (N_242,In_726,In_490);
and U243 (N_243,In_558,In_432);
and U244 (N_244,In_245,In_547);
and U245 (N_245,In_229,In_57);
nand U246 (N_246,In_367,In_659);
and U247 (N_247,In_125,In_641);
xnor U248 (N_248,In_411,In_424);
or U249 (N_249,In_171,In_622);
and U250 (N_250,In_642,In_534);
nand U251 (N_251,In_276,In_128);
xor U252 (N_252,In_147,In_51);
xor U253 (N_253,In_400,In_357);
or U254 (N_254,In_435,In_34);
xnor U255 (N_255,In_361,In_129);
nor U256 (N_256,In_112,In_30);
and U257 (N_257,In_682,In_526);
nor U258 (N_258,In_549,In_234);
and U259 (N_259,In_309,In_105);
nor U260 (N_260,In_699,In_181);
and U261 (N_261,In_712,In_244);
xnor U262 (N_262,In_600,In_623);
nand U263 (N_263,In_80,In_621);
nor U264 (N_264,In_544,In_609);
nand U265 (N_265,In_277,In_364);
and U266 (N_266,In_36,In_713);
nor U267 (N_267,In_394,In_17);
nor U268 (N_268,In_472,In_84);
nor U269 (N_269,In_97,In_507);
nor U270 (N_270,In_157,In_736);
nor U271 (N_271,In_453,In_619);
and U272 (N_272,In_655,In_11);
and U273 (N_273,In_744,In_24);
and U274 (N_274,In_28,In_40);
nand U275 (N_275,In_230,In_420);
and U276 (N_276,In_706,In_529);
and U277 (N_277,In_269,In_372);
nand U278 (N_278,In_227,In_325);
nor U279 (N_279,In_467,In_696);
or U280 (N_280,In_625,In_598);
or U281 (N_281,In_273,In_688);
or U282 (N_282,In_178,In_241);
or U283 (N_283,In_578,In_96);
nor U284 (N_284,In_371,In_651);
nand U285 (N_285,In_142,In_261);
or U286 (N_286,In_545,In_237);
or U287 (N_287,In_174,In_647);
and U288 (N_288,In_15,In_264);
nand U289 (N_289,In_535,In_448);
nor U290 (N_290,In_640,In_203);
nor U291 (N_291,In_133,In_664);
or U292 (N_292,In_447,In_189);
nor U293 (N_293,In_646,In_636);
and U294 (N_294,In_271,In_675);
xnor U295 (N_295,In_323,In_54);
nor U296 (N_296,In_156,In_100);
nor U297 (N_297,In_569,In_618);
or U298 (N_298,In_265,In_559);
nand U299 (N_299,In_454,In_597);
nand U300 (N_300,In_701,In_652);
nand U301 (N_301,In_78,In_560);
nand U302 (N_302,In_334,In_14);
or U303 (N_303,In_718,In_481);
nor U304 (N_304,In_704,In_223);
and U305 (N_305,In_686,In_645);
and U306 (N_306,In_720,In_563);
nand U307 (N_307,In_72,In_562);
nor U308 (N_308,In_354,In_550);
or U309 (N_309,In_599,In_470);
and U310 (N_310,In_21,In_353);
or U311 (N_311,In_380,In_639);
and U312 (N_312,In_615,In_162);
xor U313 (N_313,In_389,In_295);
nand U314 (N_314,In_262,In_374);
and U315 (N_315,In_658,In_455);
or U316 (N_316,In_412,In_433);
or U317 (N_317,In_316,In_518);
and U318 (N_318,In_465,In_561);
xnor U319 (N_319,In_568,In_548);
and U320 (N_320,In_740,In_35);
or U321 (N_321,In_611,In_734);
nor U322 (N_322,In_434,In_668);
nor U323 (N_323,In_260,In_195);
and U324 (N_324,In_571,In_46);
nor U325 (N_325,In_445,In_630);
nand U326 (N_326,In_339,In_464);
nor U327 (N_327,In_430,In_496);
nor U328 (N_328,In_240,In_119);
nor U329 (N_329,In_343,In_595);
nand U330 (N_330,In_250,In_395);
or U331 (N_331,In_446,In_39);
nand U332 (N_332,In_191,In_319);
nor U333 (N_333,In_236,In_503);
nand U334 (N_334,In_691,In_480);
xnor U335 (N_335,In_243,In_158);
nand U336 (N_336,In_463,In_116);
and U337 (N_337,In_198,In_410);
or U338 (N_338,In_349,In_305);
and U339 (N_339,In_532,In_730);
and U340 (N_340,In_232,In_224);
nand U341 (N_341,In_422,In_444);
and U342 (N_342,In_594,In_163);
or U343 (N_343,In_368,In_186);
nor U344 (N_344,In_588,In_705);
and U345 (N_345,In_315,In_381);
nor U346 (N_346,In_392,In_539);
nor U347 (N_347,In_654,In_149);
and U348 (N_348,In_31,In_267);
or U349 (N_349,In_370,In_320);
nand U350 (N_350,In_215,In_275);
and U351 (N_351,In_515,In_42);
or U352 (N_352,In_396,In_660);
nor U353 (N_353,In_458,In_293);
or U354 (N_354,In_747,In_359);
and U355 (N_355,In_499,In_76);
nor U356 (N_356,In_213,In_340);
nor U357 (N_357,In_117,In_478);
nand U358 (N_358,In_702,In_514);
or U359 (N_359,In_703,In_281);
nand U360 (N_360,In_115,In_698);
nand U361 (N_361,In_64,In_612);
nand U362 (N_362,In_541,In_672);
and U363 (N_363,In_661,In_106);
nor U364 (N_364,In_708,In_140);
or U365 (N_365,In_408,In_108);
and U366 (N_366,In_249,In_723);
nand U367 (N_367,In_60,In_501);
or U368 (N_368,In_209,In_369);
nor U369 (N_369,In_409,In_608);
nor U370 (N_370,In_228,In_33);
or U371 (N_371,In_32,In_451);
and U372 (N_372,In_263,In_697);
xnor U373 (N_373,In_208,In_601);
and U374 (N_374,In_491,In_62);
and U375 (N_375,In_69,In_591);
nor U376 (N_376,In_386,In_474);
and U377 (N_377,In_386,In_138);
nand U378 (N_378,In_442,In_160);
nand U379 (N_379,In_296,In_393);
nor U380 (N_380,In_140,In_152);
nor U381 (N_381,In_359,In_146);
nor U382 (N_382,In_522,In_32);
nand U383 (N_383,In_140,In_683);
nor U384 (N_384,In_108,In_257);
or U385 (N_385,In_658,In_145);
nor U386 (N_386,In_66,In_420);
xnor U387 (N_387,In_222,In_13);
nor U388 (N_388,In_386,In_589);
nand U389 (N_389,In_562,In_528);
and U390 (N_390,In_385,In_405);
or U391 (N_391,In_254,In_568);
or U392 (N_392,In_482,In_518);
nand U393 (N_393,In_687,In_740);
xnor U394 (N_394,In_722,In_314);
xor U395 (N_395,In_91,In_741);
xnor U396 (N_396,In_699,In_495);
nand U397 (N_397,In_522,In_506);
or U398 (N_398,In_656,In_505);
and U399 (N_399,In_561,In_370);
nand U400 (N_400,In_359,In_209);
xnor U401 (N_401,In_331,In_471);
and U402 (N_402,In_665,In_676);
nand U403 (N_403,In_722,In_525);
and U404 (N_404,In_90,In_360);
nor U405 (N_405,In_185,In_44);
nor U406 (N_406,In_197,In_539);
nor U407 (N_407,In_185,In_96);
and U408 (N_408,In_37,In_733);
nor U409 (N_409,In_517,In_418);
and U410 (N_410,In_556,In_521);
and U411 (N_411,In_620,In_77);
and U412 (N_412,In_36,In_35);
and U413 (N_413,In_412,In_409);
or U414 (N_414,In_358,In_681);
or U415 (N_415,In_323,In_560);
nand U416 (N_416,In_674,In_421);
or U417 (N_417,In_90,In_433);
nor U418 (N_418,In_677,In_253);
nor U419 (N_419,In_604,In_146);
or U420 (N_420,In_59,In_732);
nand U421 (N_421,In_288,In_465);
nor U422 (N_422,In_171,In_7);
xor U423 (N_423,In_708,In_233);
nor U424 (N_424,In_87,In_721);
and U425 (N_425,In_510,In_492);
nor U426 (N_426,In_264,In_590);
nor U427 (N_427,In_424,In_267);
and U428 (N_428,In_643,In_445);
or U429 (N_429,In_42,In_527);
or U430 (N_430,In_480,In_581);
and U431 (N_431,In_674,In_27);
and U432 (N_432,In_245,In_660);
nor U433 (N_433,In_631,In_453);
nand U434 (N_434,In_394,In_701);
nor U435 (N_435,In_480,In_39);
or U436 (N_436,In_462,In_360);
or U437 (N_437,In_431,In_500);
nor U438 (N_438,In_452,In_666);
nor U439 (N_439,In_467,In_580);
or U440 (N_440,In_677,In_57);
or U441 (N_441,In_745,In_298);
nor U442 (N_442,In_382,In_744);
nor U443 (N_443,In_447,In_313);
nor U444 (N_444,In_450,In_446);
and U445 (N_445,In_157,In_554);
and U446 (N_446,In_545,In_319);
nand U447 (N_447,In_4,In_539);
and U448 (N_448,In_171,In_320);
nand U449 (N_449,In_5,In_188);
or U450 (N_450,In_228,In_680);
xor U451 (N_451,In_9,In_672);
xor U452 (N_452,In_546,In_483);
nor U453 (N_453,In_294,In_142);
nor U454 (N_454,In_524,In_182);
or U455 (N_455,In_466,In_614);
nor U456 (N_456,In_88,In_292);
or U457 (N_457,In_253,In_441);
or U458 (N_458,In_621,In_232);
nand U459 (N_459,In_194,In_749);
and U460 (N_460,In_404,In_285);
or U461 (N_461,In_412,In_527);
xor U462 (N_462,In_184,In_45);
nor U463 (N_463,In_106,In_172);
or U464 (N_464,In_452,In_515);
and U465 (N_465,In_179,In_62);
and U466 (N_466,In_69,In_419);
nor U467 (N_467,In_178,In_490);
and U468 (N_468,In_161,In_164);
and U469 (N_469,In_478,In_30);
and U470 (N_470,In_194,In_548);
xnor U471 (N_471,In_218,In_727);
nor U472 (N_472,In_222,In_127);
nand U473 (N_473,In_236,In_178);
nand U474 (N_474,In_483,In_570);
xor U475 (N_475,In_378,In_53);
or U476 (N_476,In_529,In_452);
nor U477 (N_477,In_574,In_277);
xnor U478 (N_478,In_648,In_598);
xor U479 (N_479,In_113,In_8);
nor U480 (N_480,In_143,In_366);
xor U481 (N_481,In_566,In_608);
or U482 (N_482,In_703,In_579);
nand U483 (N_483,In_86,In_477);
nor U484 (N_484,In_297,In_284);
or U485 (N_485,In_156,In_18);
and U486 (N_486,In_281,In_74);
or U487 (N_487,In_390,In_615);
nand U488 (N_488,In_67,In_212);
and U489 (N_489,In_550,In_423);
nor U490 (N_490,In_294,In_540);
nand U491 (N_491,In_733,In_585);
nor U492 (N_492,In_256,In_242);
or U493 (N_493,In_496,In_587);
and U494 (N_494,In_357,In_526);
nand U495 (N_495,In_687,In_211);
nor U496 (N_496,In_515,In_100);
xnor U497 (N_497,In_631,In_368);
and U498 (N_498,In_633,In_406);
nor U499 (N_499,In_482,In_651);
or U500 (N_500,In_569,In_486);
xnor U501 (N_501,In_733,In_576);
and U502 (N_502,In_508,In_22);
and U503 (N_503,In_114,In_399);
and U504 (N_504,In_134,In_496);
and U505 (N_505,In_637,In_66);
xor U506 (N_506,In_449,In_676);
and U507 (N_507,In_305,In_442);
nor U508 (N_508,In_448,In_205);
or U509 (N_509,In_683,In_20);
nand U510 (N_510,In_6,In_361);
nand U511 (N_511,In_61,In_132);
nand U512 (N_512,In_193,In_112);
nand U513 (N_513,In_76,In_376);
nand U514 (N_514,In_588,In_204);
or U515 (N_515,In_672,In_693);
nand U516 (N_516,In_29,In_398);
and U517 (N_517,In_718,In_246);
and U518 (N_518,In_526,In_37);
nand U519 (N_519,In_400,In_610);
nor U520 (N_520,In_106,In_144);
and U521 (N_521,In_713,In_687);
nand U522 (N_522,In_272,In_47);
nor U523 (N_523,In_373,In_488);
nand U524 (N_524,In_28,In_566);
or U525 (N_525,In_718,In_85);
nor U526 (N_526,In_39,In_415);
nor U527 (N_527,In_16,In_596);
nand U528 (N_528,In_489,In_487);
xor U529 (N_529,In_59,In_255);
nor U530 (N_530,In_291,In_297);
nand U531 (N_531,In_200,In_710);
or U532 (N_532,In_491,In_540);
nor U533 (N_533,In_197,In_691);
and U534 (N_534,In_500,In_252);
and U535 (N_535,In_487,In_294);
or U536 (N_536,In_341,In_185);
and U537 (N_537,In_6,In_166);
and U538 (N_538,In_36,In_125);
or U539 (N_539,In_488,In_443);
nor U540 (N_540,In_371,In_6);
and U541 (N_541,In_565,In_596);
nor U542 (N_542,In_648,In_102);
and U543 (N_543,In_696,In_607);
xnor U544 (N_544,In_209,In_403);
nor U545 (N_545,In_226,In_704);
or U546 (N_546,In_418,In_471);
nand U547 (N_547,In_743,In_744);
and U548 (N_548,In_527,In_152);
nand U549 (N_549,In_571,In_197);
and U550 (N_550,In_440,In_628);
nand U551 (N_551,In_335,In_663);
or U552 (N_552,In_128,In_207);
and U553 (N_553,In_399,In_635);
nor U554 (N_554,In_552,In_654);
or U555 (N_555,In_213,In_579);
and U556 (N_556,In_73,In_162);
and U557 (N_557,In_317,In_41);
or U558 (N_558,In_638,In_473);
or U559 (N_559,In_703,In_612);
xnor U560 (N_560,In_445,In_13);
and U561 (N_561,In_338,In_678);
nand U562 (N_562,In_92,In_588);
nor U563 (N_563,In_656,In_571);
nor U564 (N_564,In_54,In_307);
nand U565 (N_565,In_484,In_334);
or U566 (N_566,In_326,In_508);
nand U567 (N_567,In_10,In_362);
or U568 (N_568,In_371,In_339);
nor U569 (N_569,In_425,In_506);
xnor U570 (N_570,In_252,In_308);
nor U571 (N_571,In_66,In_496);
or U572 (N_572,In_667,In_732);
nor U573 (N_573,In_609,In_470);
xnor U574 (N_574,In_429,In_411);
nand U575 (N_575,In_2,In_89);
or U576 (N_576,In_53,In_553);
nand U577 (N_577,In_246,In_579);
nand U578 (N_578,In_391,In_138);
nand U579 (N_579,In_348,In_620);
or U580 (N_580,In_430,In_662);
nand U581 (N_581,In_113,In_349);
and U582 (N_582,In_642,In_560);
nand U583 (N_583,In_674,In_70);
nand U584 (N_584,In_20,In_647);
nor U585 (N_585,In_271,In_383);
or U586 (N_586,In_302,In_502);
nand U587 (N_587,In_46,In_326);
nand U588 (N_588,In_567,In_623);
or U589 (N_589,In_535,In_572);
nor U590 (N_590,In_677,In_191);
nand U591 (N_591,In_309,In_496);
and U592 (N_592,In_69,In_731);
and U593 (N_593,In_434,In_193);
or U594 (N_594,In_254,In_38);
and U595 (N_595,In_748,In_62);
xnor U596 (N_596,In_748,In_238);
or U597 (N_597,In_523,In_543);
nand U598 (N_598,In_107,In_376);
nand U599 (N_599,In_437,In_612);
xnor U600 (N_600,In_503,In_669);
nor U601 (N_601,In_746,In_365);
nand U602 (N_602,In_110,In_339);
nand U603 (N_603,In_554,In_438);
or U604 (N_604,In_460,In_231);
or U605 (N_605,In_164,In_529);
and U606 (N_606,In_443,In_284);
or U607 (N_607,In_313,In_106);
nand U608 (N_608,In_478,In_641);
or U609 (N_609,In_214,In_211);
and U610 (N_610,In_570,In_50);
and U611 (N_611,In_463,In_615);
nand U612 (N_612,In_432,In_686);
nand U613 (N_613,In_509,In_117);
nor U614 (N_614,In_254,In_424);
nand U615 (N_615,In_192,In_142);
and U616 (N_616,In_262,In_127);
or U617 (N_617,In_432,In_723);
nor U618 (N_618,In_410,In_129);
and U619 (N_619,In_12,In_607);
nor U620 (N_620,In_192,In_598);
nor U621 (N_621,In_504,In_721);
and U622 (N_622,In_250,In_592);
nand U623 (N_623,In_181,In_713);
nand U624 (N_624,In_270,In_373);
and U625 (N_625,In_144,In_32);
or U626 (N_626,In_634,In_308);
and U627 (N_627,In_110,In_258);
nor U628 (N_628,In_280,In_645);
nand U629 (N_629,In_87,In_551);
or U630 (N_630,In_352,In_701);
nor U631 (N_631,In_278,In_618);
or U632 (N_632,In_483,In_73);
nand U633 (N_633,In_526,In_294);
and U634 (N_634,In_460,In_603);
nand U635 (N_635,In_402,In_514);
or U636 (N_636,In_710,In_527);
nand U637 (N_637,In_120,In_725);
nand U638 (N_638,In_539,In_57);
or U639 (N_639,In_107,In_665);
nand U640 (N_640,In_463,In_312);
xor U641 (N_641,In_683,In_658);
nand U642 (N_642,In_606,In_504);
or U643 (N_643,In_288,In_201);
or U644 (N_644,In_144,In_561);
and U645 (N_645,In_255,In_152);
nand U646 (N_646,In_634,In_625);
or U647 (N_647,In_335,In_372);
nand U648 (N_648,In_242,In_414);
or U649 (N_649,In_425,In_467);
nor U650 (N_650,In_332,In_569);
xor U651 (N_651,In_636,In_323);
xnor U652 (N_652,In_186,In_543);
or U653 (N_653,In_202,In_50);
nor U654 (N_654,In_428,In_10);
or U655 (N_655,In_175,In_561);
or U656 (N_656,In_74,In_482);
xor U657 (N_657,In_691,In_104);
nand U658 (N_658,In_724,In_285);
nor U659 (N_659,In_296,In_317);
and U660 (N_660,In_88,In_710);
and U661 (N_661,In_636,In_127);
or U662 (N_662,In_640,In_558);
xor U663 (N_663,In_72,In_740);
or U664 (N_664,In_621,In_54);
nor U665 (N_665,In_344,In_327);
or U666 (N_666,In_87,In_667);
and U667 (N_667,In_173,In_85);
nand U668 (N_668,In_681,In_323);
nand U669 (N_669,In_404,In_175);
nor U670 (N_670,In_339,In_554);
and U671 (N_671,In_515,In_6);
and U672 (N_672,In_472,In_520);
nor U673 (N_673,In_679,In_664);
or U674 (N_674,In_486,In_139);
nand U675 (N_675,In_346,In_223);
nor U676 (N_676,In_599,In_123);
xor U677 (N_677,In_44,In_267);
and U678 (N_678,In_274,In_560);
nand U679 (N_679,In_611,In_23);
xnor U680 (N_680,In_393,In_396);
nand U681 (N_681,In_655,In_41);
nor U682 (N_682,In_557,In_741);
nand U683 (N_683,In_220,In_66);
or U684 (N_684,In_371,In_322);
xor U685 (N_685,In_87,In_47);
nand U686 (N_686,In_376,In_535);
nor U687 (N_687,In_495,In_5);
or U688 (N_688,In_361,In_704);
and U689 (N_689,In_352,In_537);
and U690 (N_690,In_324,In_101);
nand U691 (N_691,In_406,In_452);
or U692 (N_692,In_116,In_400);
nor U693 (N_693,In_96,In_19);
nand U694 (N_694,In_646,In_663);
or U695 (N_695,In_437,In_191);
nand U696 (N_696,In_110,In_156);
nand U697 (N_697,In_383,In_695);
nor U698 (N_698,In_532,In_745);
and U699 (N_699,In_200,In_150);
nor U700 (N_700,In_153,In_712);
nor U701 (N_701,In_563,In_730);
or U702 (N_702,In_322,In_1);
or U703 (N_703,In_743,In_275);
xor U704 (N_704,In_594,In_94);
nor U705 (N_705,In_315,In_481);
and U706 (N_706,In_424,In_613);
nand U707 (N_707,In_637,In_485);
or U708 (N_708,In_114,In_270);
nand U709 (N_709,In_677,In_298);
nand U710 (N_710,In_139,In_479);
nand U711 (N_711,In_465,In_192);
nand U712 (N_712,In_407,In_553);
or U713 (N_713,In_30,In_699);
nand U714 (N_714,In_375,In_45);
nor U715 (N_715,In_177,In_625);
nor U716 (N_716,In_194,In_420);
nand U717 (N_717,In_648,In_351);
xnor U718 (N_718,In_285,In_628);
xnor U719 (N_719,In_477,In_724);
xor U720 (N_720,In_115,In_430);
and U721 (N_721,In_167,In_156);
or U722 (N_722,In_507,In_635);
and U723 (N_723,In_39,In_538);
or U724 (N_724,In_676,In_610);
or U725 (N_725,In_671,In_617);
and U726 (N_726,In_128,In_371);
xnor U727 (N_727,In_435,In_243);
and U728 (N_728,In_474,In_105);
xor U729 (N_729,In_647,In_496);
or U730 (N_730,In_369,In_646);
xnor U731 (N_731,In_680,In_299);
xnor U732 (N_732,In_104,In_80);
and U733 (N_733,In_194,In_472);
and U734 (N_734,In_189,In_740);
nand U735 (N_735,In_255,In_747);
nor U736 (N_736,In_26,In_697);
nor U737 (N_737,In_685,In_589);
xnor U738 (N_738,In_354,In_714);
nand U739 (N_739,In_244,In_339);
or U740 (N_740,In_692,In_344);
nor U741 (N_741,In_146,In_342);
nor U742 (N_742,In_580,In_473);
or U743 (N_743,In_234,In_615);
and U744 (N_744,In_254,In_269);
or U745 (N_745,In_345,In_226);
nor U746 (N_746,In_538,In_152);
or U747 (N_747,In_415,In_172);
or U748 (N_748,In_658,In_160);
and U749 (N_749,In_282,In_72);
nor U750 (N_750,In_454,In_217);
or U751 (N_751,In_378,In_471);
nand U752 (N_752,In_100,In_332);
xnor U753 (N_753,In_137,In_705);
nand U754 (N_754,In_678,In_662);
nand U755 (N_755,In_226,In_68);
nand U756 (N_756,In_198,In_637);
nand U757 (N_757,In_429,In_148);
or U758 (N_758,In_615,In_387);
nand U759 (N_759,In_474,In_568);
and U760 (N_760,In_47,In_295);
nand U761 (N_761,In_313,In_419);
and U762 (N_762,In_399,In_674);
or U763 (N_763,In_457,In_448);
nor U764 (N_764,In_458,In_313);
nor U765 (N_765,In_384,In_155);
nor U766 (N_766,In_317,In_607);
and U767 (N_767,In_392,In_17);
or U768 (N_768,In_602,In_247);
and U769 (N_769,In_127,In_239);
nor U770 (N_770,In_392,In_303);
or U771 (N_771,In_437,In_572);
and U772 (N_772,In_518,In_700);
nor U773 (N_773,In_249,In_46);
nand U774 (N_774,In_53,In_447);
and U775 (N_775,In_109,In_187);
or U776 (N_776,In_161,In_432);
nand U777 (N_777,In_364,In_341);
or U778 (N_778,In_371,In_530);
and U779 (N_779,In_379,In_366);
xor U780 (N_780,In_514,In_655);
and U781 (N_781,In_134,In_741);
and U782 (N_782,In_265,In_348);
or U783 (N_783,In_449,In_252);
xor U784 (N_784,In_430,In_631);
xor U785 (N_785,In_308,In_350);
nor U786 (N_786,In_9,In_443);
nor U787 (N_787,In_150,In_114);
and U788 (N_788,In_651,In_112);
nand U789 (N_789,In_402,In_238);
nand U790 (N_790,In_132,In_634);
nand U791 (N_791,In_736,In_230);
and U792 (N_792,In_661,In_116);
or U793 (N_793,In_55,In_22);
and U794 (N_794,In_283,In_421);
xor U795 (N_795,In_567,In_44);
and U796 (N_796,In_111,In_667);
or U797 (N_797,In_146,In_383);
nor U798 (N_798,In_396,In_492);
or U799 (N_799,In_109,In_466);
nand U800 (N_800,In_74,In_551);
xnor U801 (N_801,In_137,In_311);
nor U802 (N_802,In_477,In_648);
nand U803 (N_803,In_494,In_140);
nor U804 (N_804,In_332,In_647);
xnor U805 (N_805,In_592,In_111);
nand U806 (N_806,In_241,In_33);
nor U807 (N_807,In_737,In_534);
nor U808 (N_808,In_118,In_596);
xor U809 (N_809,In_348,In_354);
nand U810 (N_810,In_235,In_452);
and U811 (N_811,In_745,In_308);
and U812 (N_812,In_439,In_565);
nor U813 (N_813,In_732,In_408);
nor U814 (N_814,In_505,In_39);
nand U815 (N_815,In_555,In_184);
or U816 (N_816,In_482,In_732);
or U817 (N_817,In_634,In_233);
or U818 (N_818,In_47,In_704);
or U819 (N_819,In_646,In_69);
nand U820 (N_820,In_301,In_466);
or U821 (N_821,In_410,In_744);
and U822 (N_822,In_406,In_536);
and U823 (N_823,In_220,In_714);
and U824 (N_824,In_720,In_600);
xnor U825 (N_825,In_163,In_700);
or U826 (N_826,In_437,In_461);
or U827 (N_827,In_42,In_725);
nor U828 (N_828,In_516,In_328);
nand U829 (N_829,In_390,In_245);
nand U830 (N_830,In_81,In_361);
nand U831 (N_831,In_649,In_27);
nor U832 (N_832,In_451,In_250);
nand U833 (N_833,In_443,In_413);
nand U834 (N_834,In_674,In_469);
and U835 (N_835,In_417,In_722);
and U836 (N_836,In_294,In_530);
nor U837 (N_837,In_338,In_312);
and U838 (N_838,In_560,In_477);
nand U839 (N_839,In_223,In_82);
or U840 (N_840,In_181,In_100);
or U841 (N_841,In_278,In_353);
or U842 (N_842,In_130,In_30);
and U843 (N_843,In_486,In_538);
nand U844 (N_844,In_503,In_220);
and U845 (N_845,In_239,In_80);
nor U846 (N_846,In_452,In_728);
nand U847 (N_847,In_736,In_420);
and U848 (N_848,In_202,In_727);
nor U849 (N_849,In_138,In_137);
xor U850 (N_850,In_657,In_558);
and U851 (N_851,In_464,In_353);
and U852 (N_852,In_438,In_635);
nand U853 (N_853,In_65,In_500);
xor U854 (N_854,In_55,In_160);
nand U855 (N_855,In_206,In_464);
or U856 (N_856,In_523,In_129);
and U857 (N_857,In_365,In_472);
xnor U858 (N_858,In_292,In_705);
and U859 (N_859,In_160,In_550);
and U860 (N_860,In_169,In_193);
nand U861 (N_861,In_329,In_396);
nor U862 (N_862,In_731,In_123);
xor U863 (N_863,In_150,In_119);
xor U864 (N_864,In_746,In_210);
xnor U865 (N_865,In_148,In_363);
nand U866 (N_866,In_6,In_112);
or U867 (N_867,In_405,In_601);
and U868 (N_868,In_159,In_140);
and U869 (N_869,In_489,In_226);
or U870 (N_870,In_119,In_232);
nand U871 (N_871,In_459,In_178);
and U872 (N_872,In_515,In_288);
or U873 (N_873,In_420,In_577);
or U874 (N_874,In_123,In_144);
nand U875 (N_875,In_48,In_164);
and U876 (N_876,In_164,In_15);
xor U877 (N_877,In_409,In_484);
nand U878 (N_878,In_142,In_326);
nor U879 (N_879,In_407,In_19);
nand U880 (N_880,In_712,In_305);
or U881 (N_881,In_286,In_684);
nand U882 (N_882,In_587,In_633);
and U883 (N_883,In_362,In_372);
or U884 (N_884,In_89,In_164);
nand U885 (N_885,In_328,In_132);
and U886 (N_886,In_277,In_192);
nand U887 (N_887,In_718,In_576);
or U888 (N_888,In_454,In_474);
nand U889 (N_889,In_28,In_271);
or U890 (N_890,In_185,In_597);
and U891 (N_891,In_744,In_288);
nand U892 (N_892,In_637,In_501);
xor U893 (N_893,In_363,In_697);
nand U894 (N_894,In_378,In_680);
or U895 (N_895,In_657,In_689);
nor U896 (N_896,In_535,In_398);
nor U897 (N_897,In_521,In_531);
nor U898 (N_898,In_66,In_410);
xnor U899 (N_899,In_90,In_17);
nor U900 (N_900,In_383,In_610);
and U901 (N_901,In_490,In_350);
or U902 (N_902,In_218,In_550);
or U903 (N_903,In_189,In_104);
or U904 (N_904,In_471,In_506);
nor U905 (N_905,In_215,In_357);
xor U906 (N_906,In_475,In_217);
nand U907 (N_907,In_60,In_80);
nand U908 (N_908,In_639,In_58);
or U909 (N_909,In_17,In_229);
or U910 (N_910,In_352,In_636);
or U911 (N_911,In_92,In_256);
nor U912 (N_912,In_394,In_338);
and U913 (N_913,In_462,In_365);
xor U914 (N_914,In_620,In_284);
and U915 (N_915,In_601,In_522);
or U916 (N_916,In_354,In_385);
and U917 (N_917,In_389,In_120);
or U918 (N_918,In_275,In_385);
nor U919 (N_919,In_59,In_502);
and U920 (N_920,In_494,In_366);
xnor U921 (N_921,In_730,In_693);
xnor U922 (N_922,In_539,In_617);
and U923 (N_923,In_352,In_192);
and U924 (N_924,In_678,In_631);
nand U925 (N_925,In_642,In_556);
nor U926 (N_926,In_640,In_143);
nand U927 (N_927,In_27,In_249);
or U928 (N_928,In_687,In_564);
or U929 (N_929,In_8,In_530);
nor U930 (N_930,In_24,In_634);
or U931 (N_931,In_669,In_44);
or U932 (N_932,In_287,In_581);
nand U933 (N_933,In_717,In_441);
or U934 (N_934,In_661,In_133);
xnor U935 (N_935,In_167,In_201);
nor U936 (N_936,In_160,In_302);
nor U937 (N_937,In_257,In_360);
nor U938 (N_938,In_491,In_531);
nand U939 (N_939,In_214,In_534);
nor U940 (N_940,In_406,In_10);
or U941 (N_941,In_501,In_323);
and U942 (N_942,In_601,In_179);
nor U943 (N_943,In_148,In_312);
nand U944 (N_944,In_476,In_624);
nand U945 (N_945,In_369,In_73);
and U946 (N_946,In_204,In_198);
nor U947 (N_947,In_368,In_438);
xnor U948 (N_948,In_176,In_402);
nand U949 (N_949,In_656,In_590);
or U950 (N_950,In_193,In_521);
nor U951 (N_951,In_656,In_10);
nor U952 (N_952,In_550,In_363);
nand U953 (N_953,In_42,In_433);
xor U954 (N_954,In_330,In_346);
or U955 (N_955,In_458,In_596);
and U956 (N_956,In_414,In_617);
nand U957 (N_957,In_624,In_433);
nor U958 (N_958,In_621,In_78);
or U959 (N_959,In_86,In_106);
xnor U960 (N_960,In_84,In_76);
nand U961 (N_961,In_438,In_748);
or U962 (N_962,In_79,In_316);
nor U963 (N_963,In_117,In_276);
xor U964 (N_964,In_114,In_110);
or U965 (N_965,In_643,In_515);
nor U966 (N_966,In_463,In_336);
nor U967 (N_967,In_664,In_582);
or U968 (N_968,In_124,In_553);
xnor U969 (N_969,In_194,In_673);
nand U970 (N_970,In_314,In_484);
nand U971 (N_971,In_578,In_509);
xor U972 (N_972,In_574,In_350);
and U973 (N_973,In_271,In_690);
or U974 (N_974,In_442,In_439);
nor U975 (N_975,In_213,In_165);
nand U976 (N_976,In_683,In_368);
and U977 (N_977,In_440,In_226);
xor U978 (N_978,In_538,In_58);
nor U979 (N_979,In_367,In_201);
or U980 (N_980,In_27,In_168);
or U981 (N_981,In_424,In_433);
nor U982 (N_982,In_433,In_422);
or U983 (N_983,In_469,In_67);
nor U984 (N_984,In_161,In_66);
or U985 (N_985,In_583,In_61);
or U986 (N_986,In_275,In_718);
nand U987 (N_987,In_605,In_406);
and U988 (N_988,In_535,In_746);
and U989 (N_989,In_740,In_92);
or U990 (N_990,In_470,In_560);
or U991 (N_991,In_335,In_282);
nand U992 (N_992,In_365,In_624);
nor U993 (N_993,In_231,In_473);
nand U994 (N_994,In_46,In_393);
or U995 (N_995,In_654,In_638);
nand U996 (N_996,In_208,In_288);
xor U997 (N_997,In_518,In_565);
nor U998 (N_998,In_711,In_117);
and U999 (N_999,In_664,In_251);
nor U1000 (N_1000,N_412,N_210);
or U1001 (N_1001,N_946,N_987);
or U1002 (N_1002,N_608,N_2);
or U1003 (N_1003,N_22,N_661);
nor U1004 (N_1004,N_71,N_62);
nand U1005 (N_1005,N_984,N_129);
or U1006 (N_1006,N_406,N_739);
nand U1007 (N_1007,N_386,N_950);
nand U1008 (N_1008,N_11,N_324);
and U1009 (N_1009,N_228,N_758);
xor U1010 (N_1010,N_768,N_419);
or U1011 (N_1011,N_938,N_84);
and U1012 (N_1012,N_493,N_68);
nor U1013 (N_1013,N_301,N_403);
or U1014 (N_1014,N_839,N_340);
and U1015 (N_1015,N_439,N_919);
and U1016 (N_1016,N_445,N_172);
nor U1017 (N_1017,N_920,N_229);
or U1018 (N_1018,N_422,N_627);
and U1019 (N_1019,N_204,N_654);
nand U1020 (N_1020,N_619,N_113);
nor U1021 (N_1021,N_348,N_77);
or U1022 (N_1022,N_782,N_736);
and U1023 (N_1023,N_971,N_256);
nor U1024 (N_1024,N_826,N_365);
nor U1025 (N_1025,N_359,N_441);
nor U1026 (N_1026,N_752,N_440);
nor U1027 (N_1027,N_0,N_297);
or U1028 (N_1028,N_733,N_681);
and U1029 (N_1029,N_259,N_6);
xor U1030 (N_1030,N_590,N_100);
nand U1031 (N_1031,N_261,N_392);
or U1032 (N_1032,N_218,N_285);
xnor U1033 (N_1033,N_814,N_23);
and U1034 (N_1034,N_810,N_180);
nor U1035 (N_1035,N_21,N_416);
nand U1036 (N_1036,N_250,N_596);
nor U1037 (N_1037,N_99,N_454);
nand U1038 (N_1038,N_719,N_789);
nand U1039 (N_1039,N_330,N_630);
and U1040 (N_1040,N_5,N_927);
nand U1041 (N_1041,N_443,N_888);
nand U1042 (N_1042,N_294,N_199);
or U1043 (N_1043,N_354,N_90);
nor U1044 (N_1044,N_565,N_232);
nand U1045 (N_1045,N_50,N_308);
nand U1046 (N_1046,N_853,N_76);
nand U1047 (N_1047,N_155,N_185);
or U1048 (N_1048,N_512,N_379);
or U1049 (N_1049,N_552,N_871);
or U1050 (N_1050,N_929,N_751);
or U1051 (N_1051,N_299,N_508);
nor U1052 (N_1052,N_833,N_221);
nor U1053 (N_1053,N_290,N_216);
xor U1054 (N_1054,N_524,N_28);
and U1055 (N_1055,N_741,N_277);
or U1056 (N_1056,N_343,N_905);
and U1057 (N_1057,N_885,N_603);
nor U1058 (N_1058,N_790,N_135);
nor U1059 (N_1059,N_179,N_132);
xnor U1060 (N_1060,N_588,N_479);
nand U1061 (N_1061,N_579,N_561);
nor U1062 (N_1062,N_930,N_160);
nor U1063 (N_1063,N_27,N_628);
nor U1064 (N_1064,N_591,N_263);
and U1065 (N_1065,N_63,N_693);
or U1066 (N_1066,N_904,N_847);
nor U1067 (N_1067,N_15,N_917);
nand U1068 (N_1068,N_677,N_426);
and U1069 (N_1069,N_257,N_241);
xor U1070 (N_1070,N_535,N_842);
and U1071 (N_1071,N_240,N_815);
xnor U1072 (N_1072,N_388,N_742);
and U1073 (N_1073,N_183,N_762);
or U1074 (N_1074,N_883,N_560);
and U1075 (N_1075,N_691,N_641);
and U1076 (N_1076,N_338,N_491);
nor U1077 (N_1077,N_666,N_586);
xor U1078 (N_1078,N_320,N_60);
nand U1079 (N_1079,N_29,N_387);
nand U1080 (N_1080,N_634,N_427);
nor U1081 (N_1081,N_662,N_602);
and U1082 (N_1082,N_319,N_632);
nor U1083 (N_1083,N_333,N_342);
xor U1084 (N_1084,N_611,N_543);
nor U1085 (N_1085,N_248,N_209);
and U1086 (N_1086,N_214,N_570);
and U1087 (N_1087,N_796,N_188);
or U1088 (N_1088,N_501,N_797);
and U1089 (N_1089,N_408,N_486);
or U1090 (N_1090,N_435,N_989);
and U1091 (N_1091,N_442,N_222);
and U1092 (N_1092,N_192,N_521);
nor U1093 (N_1093,N_56,N_544);
and U1094 (N_1094,N_207,N_614);
xor U1095 (N_1095,N_566,N_609);
nand U1096 (N_1096,N_559,N_582);
xnor U1097 (N_1097,N_974,N_161);
or U1098 (N_1098,N_117,N_162);
and U1099 (N_1099,N_891,N_896);
nor U1100 (N_1100,N_546,N_410);
and U1101 (N_1101,N_889,N_146);
xnor U1102 (N_1102,N_487,N_404);
xor U1103 (N_1103,N_61,N_33);
nor U1104 (N_1104,N_370,N_541);
nor U1105 (N_1105,N_278,N_417);
nand U1106 (N_1106,N_265,N_383);
or U1107 (N_1107,N_728,N_139);
or U1108 (N_1108,N_35,N_38);
nor U1109 (N_1109,N_822,N_511);
or U1110 (N_1110,N_334,N_562);
nand U1111 (N_1111,N_931,N_345);
and U1112 (N_1112,N_481,N_536);
and U1113 (N_1113,N_202,N_203);
nor U1114 (N_1114,N_271,N_397);
and U1115 (N_1115,N_374,N_961);
nor U1116 (N_1116,N_494,N_563);
or U1117 (N_1117,N_322,N_775);
xor U1118 (N_1118,N_821,N_567);
and U1119 (N_1119,N_269,N_678);
or U1120 (N_1120,N_242,N_640);
nor U1121 (N_1121,N_391,N_451);
and U1122 (N_1122,N_252,N_761);
or U1123 (N_1123,N_41,N_85);
xor U1124 (N_1124,N_74,N_868);
or U1125 (N_1125,N_684,N_687);
or U1126 (N_1126,N_607,N_759);
nor U1127 (N_1127,N_16,N_114);
or U1128 (N_1128,N_154,N_850);
xor U1129 (N_1129,N_599,N_468);
and U1130 (N_1130,N_648,N_55);
or U1131 (N_1131,N_637,N_997);
or U1132 (N_1132,N_998,N_111);
or U1133 (N_1133,N_98,N_239);
nand U1134 (N_1134,N_288,N_353);
and U1135 (N_1135,N_610,N_975);
nand U1136 (N_1136,N_430,N_933);
nand U1137 (N_1137,N_206,N_131);
xor U1138 (N_1138,N_167,N_757);
or U1139 (N_1139,N_865,N_137);
or U1140 (N_1140,N_163,N_940);
and U1141 (N_1141,N_46,N_438);
and U1142 (N_1142,N_462,N_912);
or U1143 (N_1143,N_986,N_170);
nor U1144 (N_1144,N_247,N_522);
or U1145 (N_1145,N_300,N_86);
nand U1146 (N_1146,N_953,N_923);
and U1147 (N_1147,N_746,N_346);
nand U1148 (N_1148,N_787,N_159);
or U1149 (N_1149,N_688,N_621);
and U1150 (N_1150,N_956,N_53);
or U1151 (N_1151,N_502,N_166);
nor U1152 (N_1152,N_695,N_470);
nor U1153 (N_1153,N_367,N_431);
nor U1154 (N_1154,N_903,N_293);
nor U1155 (N_1155,N_42,N_776);
nor U1156 (N_1156,N_625,N_969);
nor U1157 (N_1157,N_716,N_496);
nor U1158 (N_1158,N_72,N_489);
nor U1159 (N_1159,N_58,N_574);
nor U1160 (N_1160,N_876,N_553);
nor U1161 (N_1161,N_44,N_725);
nand U1162 (N_1162,N_456,N_937);
and U1163 (N_1163,N_964,N_107);
and U1164 (N_1164,N_198,N_594);
and U1165 (N_1165,N_877,N_184);
or U1166 (N_1166,N_995,N_234);
and U1167 (N_1167,N_52,N_51);
nor U1168 (N_1168,N_676,N_492);
nand U1169 (N_1169,N_140,N_783);
or U1170 (N_1170,N_366,N_361);
nand U1171 (N_1171,N_701,N_474);
nand U1172 (N_1172,N_321,N_862);
or U1173 (N_1173,N_106,N_753);
or U1174 (N_1174,N_65,N_313);
nand U1175 (N_1175,N_395,N_193);
or U1176 (N_1176,N_517,N_380);
nand U1177 (N_1177,N_807,N_825);
and U1178 (N_1178,N_219,N_335);
or U1179 (N_1179,N_103,N_187);
or U1180 (N_1180,N_900,N_150);
or U1181 (N_1181,N_420,N_679);
or U1182 (N_1182,N_325,N_506);
and U1183 (N_1183,N_717,N_195);
nor U1184 (N_1184,N_573,N_755);
nand U1185 (N_1185,N_245,N_476);
and U1186 (N_1186,N_472,N_332);
nand U1187 (N_1187,N_875,N_663);
and U1188 (N_1188,N_978,N_429);
and U1189 (N_1189,N_399,N_151);
or U1190 (N_1190,N_837,N_972);
nand U1191 (N_1191,N_358,N_153);
and U1192 (N_1192,N_480,N_92);
nand U1193 (N_1193,N_942,N_624);
or U1194 (N_1194,N_460,N_623);
and U1195 (N_1195,N_326,N_727);
nand U1196 (N_1196,N_18,N_873);
nor U1197 (N_1197,N_707,N_384);
nand U1198 (N_1198,N_520,N_943);
and U1199 (N_1199,N_309,N_992);
or U1200 (N_1200,N_59,N_735);
xnor U1201 (N_1201,N_955,N_194);
and U1202 (N_1202,N_577,N_505);
xor U1203 (N_1203,N_670,N_977);
or U1204 (N_1204,N_482,N_771);
nand U1205 (N_1205,N_999,N_866);
and U1206 (N_1206,N_270,N_449);
and U1207 (N_1207,N_197,N_122);
nor U1208 (N_1208,N_740,N_777);
nor U1209 (N_1209,N_756,N_882);
or U1210 (N_1210,N_363,N_829);
and U1211 (N_1211,N_262,N_67);
nor U1212 (N_1212,N_519,N_144);
nand U1213 (N_1213,N_447,N_750);
and U1214 (N_1214,N_94,N_223);
or U1215 (N_1215,N_20,N_852);
or U1216 (N_1216,N_200,N_813);
nor U1217 (N_1217,N_601,N_948);
or U1218 (N_1218,N_105,N_69);
nor U1219 (N_1219,N_264,N_503);
or U1220 (N_1220,N_804,N_649);
nor U1221 (N_1221,N_455,N_980);
nor U1222 (N_1222,N_589,N_268);
or U1223 (N_1223,N_702,N_606);
or U1224 (N_1224,N_550,N_173);
nand U1225 (N_1225,N_851,N_409);
or U1226 (N_1226,N_729,N_638);
and U1227 (N_1227,N_500,N_737);
nor U1228 (N_1228,N_498,N_890);
nor U1229 (N_1229,N_220,N_652);
and U1230 (N_1230,N_918,N_414);
and U1231 (N_1231,N_238,N_721);
nor U1232 (N_1232,N_816,N_283);
xnor U1233 (N_1233,N_157,N_26);
nor U1234 (N_1234,N_504,N_659);
xor U1235 (N_1235,N_952,N_336);
or U1236 (N_1236,N_915,N_190);
xnor U1237 (N_1237,N_483,N_147);
or U1238 (N_1238,N_925,N_249);
nand U1239 (N_1239,N_723,N_916);
and U1240 (N_1240,N_463,N_660);
and U1241 (N_1241,N_9,N_898);
and U1242 (N_1242,N_525,N_317);
xor U1243 (N_1243,N_774,N_772);
nand U1244 (N_1244,N_243,N_713);
nor U1245 (N_1245,N_647,N_347);
nand U1246 (N_1246,N_32,N_703);
nand U1247 (N_1247,N_801,N_620);
or U1248 (N_1248,N_968,N_722);
nand U1249 (N_1249,N_415,N_78);
and U1250 (N_1250,N_475,N_726);
nand U1251 (N_1251,N_402,N_303);
nor U1252 (N_1252,N_724,N_863);
and U1253 (N_1253,N_31,N_845);
nand U1254 (N_1254,N_656,N_585);
and U1255 (N_1255,N_255,N_314);
nor U1256 (N_1256,N_108,N_189);
nand U1257 (N_1257,N_694,N_680);
or U1258 (N_1258,N_867,N_376);
nand U1259 (N_1259,N_328,N_683);
nor U1260 (N_1260,N_37,N_158);
or U1261 (N_1261,N_639,N_699);
and U1262 (N_1262,N_811,N_569);
and U1263 (N_1263,N_407,N_339);
nor U1264 (N_1264,N_149,N_584);
and U1265 (N_1265,N_175,N_548);
and U1266 (N_1266,N_692,N_509);
and U1267 (N_1267,N_64,N_284);
and U1268 (N_1268,N_327,N_864);
nor U1269 (N_1269,N_282,N_258);
nor U1270 (N_1270,N_650,N_371);
or U1271 (N_1271,N_949,N_24);
nand U1272 (N_1272,N_834,N_196);
and U1273 (N_1273,N_233,N_766);
and U1274 (N_1274,N_748,N_745);
nand U1275 (N_1275,N_617,N_141);
nand U1276 (N_1276,N_644,N_75);
xor U1277 (N_1277,N_469,N_484);
nand U1278 (N_1278,N_375,N_921);
and U1279 (N_1279,N_894,N_686);
or U1280 (N_1280,N_936,N_540);
xnor U1281 (N_1281,N_554,N_526);
and U1282 (N_1282,N_381,N_235);
or U1283 (N_1283,N_636,N_10);
nor U1284 (N_1284,N_965,N_398);
and U1285 (N_1285,N_527,N_629);
nor U1286 (N_1286,N_958,N_780);
and U1287 (N_1287,N_857,N_80);
or U1288 (N_1288,N_848,N_533);
nor U1289 (N_1289,N_884,N_858);
xnor U1290 (N_1290,N_685,N_682);
nand U1291 (N_1291,N_171,N_794);
nand U1292 (N_1292,N_444,N_529);
xnor U1293 (N_1293,N_134,N_537);
xor U1294 (N_1294,N_996,N_211);
xnor U1295 (N_1295,N_836,N_909);
and U1296 (N_1296,N_534,N_292);
nor U1297 (N_1297,N_458,N_928);
nand U1298 (N_1298,N_558,N_870);
xnor U1299 (N_1299,N_705,N_764);
and U1300 (N_1300,N_471,N_1);
nand U1301 (N_1301,N_859,N_423);
or U1302 (N_1302,N_612,N_156);
and U1303 (N_1303,N_645,N_785);
nand U1304 (N_1304,N_17,N_712);
and U1305 (N_1305,N_973,N_400);
or U1306 (N_1306,N_205,N_499);
nor U1307 (N_1307,N_838,N_213);
and U1308 (N_1308,N_227,N_30);
and U1309 (N_1309,N_176,N_805);
xor U1310 (N_1310,N_286,N_329);
or U1311 (N_1311,N_389,N_112);
and U1312 (N_1312,N_959,N_236);
nor U1313 (N_1313,N_275,N_369);
or U1314 (N_1314,N_854,N_13);
xor U1315 (N_1315,N_580,N_664);
nand U1316 (N_1316,N_267,N_164);
or U1317 (N_1317,N_800,N_911);
and U1318 (N_1318,N_360,N_101);
nor U1319 (N_1319,N_390,N_665);
and U1320 (N_1320,N_237,N_49);
xnor U1321 (N_1321,N_306,N_316);
nand U1322 (N_1322,N_467,N_799);
nand U1323 (N_1323,N_781,N_93);
and U1324 (N_1324,N_622,N_887);
or U1325 (N_1325,N_583,N_43);
or U1326 (N_1326,N_510,N_528);
and U1327 (N_1327,N_747,N_595);
nor U1328 (N_1328,N_643,N_605);
and U1329 (N_1329,N_177,N_516);
or U1330 (N_1330,N_564,N_507);
nand U1331 (N_1331,N_798,N_840);
nand U1332 (N_1332,N_899,N_715);
or U1333 (N_1333,N_73,N_254);
or U1334 (N_1334,N_276,N_675);
nor U1335 (N_1335,N_373,N_125);
and U1336 (N_1336,N_437,N_598);
xor U1337 (N_1337,N_217,N_362);
nor U1338 (N_1338,N_830,N_66);
or U1339 (N_1339,N_142,N_490);
nor U1340 (N_1340,N_658,N_831);
nand U1341 (N_1341,N_697,N_152);
xor U1342 (N_1342,N_424,N_224);
or U1343 (N_1343,N_130,N_418);
and U1344 (N_1344,N_597,N_372);
and U1345 (N_1345,N_604,N_689);
and U1346 (N_1346,N_947,N_96);
or U1347 (N_1347,N_411,N_954);
xor U1348 (N_1348,N_600,N_461);
and U1349 (N_1349,N_696,N_879);
nor U1350 (N_1350,N_57,N_350);
nor U1351 (N_1351,N_708,N_906);
and U1352 (N_1352,N_368,N_91);
and U1353 (N_1353,N_349,N_902);
nand U1354 (N_1354,N_874,N_260);
and U1355 (N_1355,N_48,N_143);
or U1356 (N_1356,N_802,N_817);
or U1357 (N_1357,N_531,N_298);
or U1358 (N_1358,N_136,N_668);
and U1359 (N_1359,N_749,N_364);
or U1360 (N_1360,N_532,N_642);
or U1361 (N_1361,N_618,N_655);
or U1362 (N_1362,N_450,N_846);
xnor U1363 (N_1363,N_849,N_844);
or U1364 (N_1364,N_121,N_653);
or U1365 (N_1365,N_119,N_148);
nor U1366 (N_1366,N_401,N_118);
or U1367 (N_1367,N_939,N_477);
nor U1368 (N_1368,N_806,N_786);
nand U1369 (N_1369,N_351,N_47);
nand U1370 (N_1370,N_88,N_993);
or U1371 (N_1371,N_672,N_710);
and U1372 (N_1372,N_792,N_626);
nand U1373 (N_1373,N_413,N_432);
nand U1374 (N_1374,N_273,N_542);
and U1375 (N_1375,N_901,N_215);
xor U1376 (N_1376,N_698,N_81);
nand U1377 (N_1377,N_377,N_545);
nor U1378 (N_1378,N_355,N_773);
nand U1379 (N_1379,N_913,N_289);
nand U1380 (N_1380,N_832,N_788);
and U1381 (N_1381,N_7,N_812);
or U1382 (N_1382,N_907,N_34);
or U1383 (N_1383,N_126,N_922);
nor U1384 (N_1384,N_89,N_79);
xnor U1385 (N_1385,N_881,N_895);
nor U1386 (N_1386,N_994,N_530);
and U1387 (N_1387,N_908,N_819);
xor U1388 (N_1388,N_791,N_557);
or U1389 (N_1389,N_356,N_754);
nor U1390 (N_1390,N_576,N_178);
or U1391 (N_1391,N_274,N_428);
or U1392 (N_1392,N_673,N_457);
nor U1393 (N_1393,N_760,N_572);
xor U1394 (N_1394,N_310,N_434);
nand U1395 (N_1395,N_495,N_935);
and U1396 (N_1396,N_244,N_83);
and U1397 (N_1397,N_425,N_892);
xor U1398 (N_1398,N_287,N_253);
or U1399 (N_1399,N_860,N_878);
and U1400 (N_1400,N_341,N_731);
nand U1401 (N_1401,N_344,N_87);
nor U1402 (N_1402,N_305,N_763);
xor U1403 (N_1403,N_824,N_593);
nand U1404 (N_1404,N_488,N_967);
nor U1405 (N_1405,N_835,N_128);
or U1406 (N_1406,N_657,N_872);
or U1407 (N_1407,N_133,N_843);
nand U1408 (N_1408,N_970,N_651);
xnor U1409 (N_1409,N_225,N_421);
or U1410 (N_1410,N_138,N_304);
xnor U1411 (N_1411,N_231,N_464);
or U1412 (N_1412,N_575,N_230);
and U1413 (N_1413,N_302,N_568);
or U1414 (N_1414,N_436,N_616);
nand U1415 (N_1415,N_944,N_646);
nor U1416 (N_1416,N_809,N_181);
nand U1417 (N_1417,N_631,N_587);
xnor U1418 (N_1418,N_97,N_39);
or U1419 (N_1419,N_704,N_497);
and U1420 (N_1420,N_910,N_478);
nor U1421 (N_1421,N_251,N_795);
xor U1422 (N_1422,N_4,N_592);
nor U1423 (N_1423,N_466,N_669);
and U1424 (N_1424,N_120,N_266);
or U1425 (N_1425,N_281,N_174);
or U1426 (N_1426,N_168,N_709);
and U1427 (N_1427,N_667,N_880);
xor U1428 (N_1428,N_485,N_893);
nor U1429 (N_1429,N_743,N_8);
xor U1430 (N_1430,N_979,N_945);
and U1431 (N_1431,N_808,N_615);
nor U1432 (N_1432,N_765,N_102);
or U1433 (N_1433,N_12,N_991);
nand U1434 (N_1434,N_394,N_538);
nand U1435 (N_1435,N_127,N_14);
nand U1436 (N_1436,N_291,N_784);
and U1437 (N_1437,N_433,N_337);
or U1438 (N_1438,N_555,N_3);
nand U1439 (N_1439,N_976,N_272);
and U1440 (N_1440,N_396,N_109);
nor U1441 (N_1441,N_123,N_983);
nand U1442 (N_1442,N_690,N_934);
nand U1443 (N_1443,N_70,N_962);
xor U1444 (N_1444,N_378,N_738);
nand U1445 (N_1445,N_452,N_246);
nor U1446 (N_1446,N_465,N_720);
nand U1447 (N_1447,N_770,N_95);
or U1448 (N_1448,N_331,N_393);
or U1449 (N_1449,N_473,N_182);
and U1450 (N_1450,N_523,N_966);
nand U1451 (N_1451,N_778,N_315);
and U1452 (N_1452,N_613,N_40);
and U1453 (N_1453,N_963,N_208);
or U1454 (N_1454,N_539,N_941);
nor U1455 (N_1455,N_820,N_960);
or U1456 (N_1456,N_191,N_116);
and U1457 (N_1457,N_54,N_855);
nor U1458 (N_1458,N_515,N_82);
and U1459 (N_1459,N_318,N_818);
or U1460 (N_1460,N_732,N_513);
nor U1461 (N_1461,N_212,N_803);
nand U1462 (N_1462,N_767,N_897);
nor U1463 (N_1463,N_549,N_985);
nor U1464 (N_1464,N_926,N_514);
nor U1465 (N_1465,N_571,N_700);
nor U1466 (N_1466,N_734,N_45);
or U1467 (N_1467,N_279,N_124);
or U1468 (N_1468,N_226,N_982);
or U1469 (N_1469,N_827,N_932);
and U1470 (N_1470,N_357,N_841);
or U1471 (N_1471,N_861,N_990);
nor U1472 (N_1472,N_110,N_793);
nor U1473 (N_1473,N_518,N_19);
or U1474 (N_1474,N_385,N_169);
and U1475 (N_1475,N_886,N_115);
xnor U1476 (N_1476,N_311,N_448);
or U1477 (N_1477,N_459,N_578);
nand U1478 (N_1478,N_914,N_671);
or U1479 (N_1479,N_453,N_405);
nand U1480 (N_1480,N_988,N_744);
xor U1481 (N_1481,N_280,N_924);
nor U1482 (N_1482,N_382,N_145);
and U1483 (N_1483,N_556,N_633);
and U1484 (N_1484,N_674,N_730);
nand U1485 (N_1485,N_165,N_856);
or U1486 (N_1486,N_323,N_714);
or U1487 (N_1487,N_312,N_828);
nand U1488 (N_1488,N_957,N_547);
nor U1489 (N_1489,N_201,N_951);
nor U1490 (N_1490,N_581,N_352);
nor U1491 (N_1491,N_981,N_307);
xor U1492 (N_1492,N_186,N_718);
nand U1493 (N_1493,N_25,N_769);
or U1494 (N_1494,N_869,N_551);
and U1495 (N_1495,N_823,N_706);
nor U1496 (N_1496,N_635,N_296);
or U1497 (N_1497,N_104,N_295);
nand U1498 (N_1498,N_36,N_446);
nand U1499 (N_1499,N_779,N_711);
or U1500 (N_1500,N_498,N_987);
and U1501 (N_1501,N_467,N_636);
nor U1502 (N_1502,N_995,N_10);
or U1503 (N_1503,N_83,N_111);
nor U1504 (N_1504,N_224,N_255);
or U1505 (N_1505,N_148,N_734);
nor U1506 (N_1506,N_305,N_289);
nor U1507 (N_1507,N_292,N_577);
or U1508 (N_1508,N_381,N_718);
nor U1509 (N_1509,N_921,N_292);
nand U1510 (N_1510,N_389,N_682);
nor U1511 (N_1511,N_678,N_102);
nand U1512 (N_1512,N_998,N_59);
nand U1513 (N_1513,N_49,N_171);
nand U1514 (N_1514,N_126,N_479);
and U1515 (N_1515,N_768,N_642);
nor U1516 (N_1516,N_953,N_190);
and U1517 (N_1517,N_295,N_729);
nand U1518 (N_1518,N_863,N_125);
nand U1519 (N_1519,N_605,N_214);
nand U1520 (N_1520,N_505,N_835);
nor U1521 (N_1521,N_83,N_956);
and U1522 (N_1522,N_853,N_825);
and U1523 (N_1523,N_807,N_900);
and U1524 (N_1524,N_214,N_569);
xnor U1525 (N_1525,N_149,N_314);
or U1526 (N_1526,N_125,N_404);
nor U1527 (N_1527,N_3,N_549);
or U1528 (N_1528,N_814,N_492);
and U1529 (N_1529,N_334,N_769);
and U1530 (N_1530,N_596,N_582);
nand U1531 (N_1531,N_169,N_724);
nor U1532 (N_1532,N_805,N_918);
or U1533 (N_1533,N_776,N_641);
nor U1534 (N_1534,N_878,N_898);
and U1535 (N_1535,N_686,N_709);
xnor U1536 (N_1536,N_493,N_381);
or U1537 (N_1537,N_105,N_429);
nand U1538 (N_1538,N_562,N_565);
and U1539 (N_1539,N_120,N_282);
nor U1540 (N_1540,N_861,N_862);
and U1541 (N_1541,N_345,N_114);
or U1542 (N_1542,N_676,N_707);
nor U1543 (N_1543,N_612,N_991);
or U1544 (N_1544,N_911,N_510);
nor U1545 (N_1545,N_558,N_728);
xor U1546 (N_1546,N_334,N_645);
and U1547 (N_1547,N_581,N_158);
and U1548 (N_1548,N_626,N_615);
xor U1549 (N_1549,N_605,N_218);
nand U1550 (N_1550,N_917,N_818);
or U1551 (N_1551,N_862,N_772);
nand U1552 (N_1552,N_431,N_723);
nand U1553 (N_1553,N_962,N_302);
or U1554 (N_1554,N_983,N_566);
and U1555 (N_1555,N_163,N_282);
and U1556 (N_1556,N_126,N_710);
xor U1557 (N_1557,N_376,N_428);
or U1558 (N_1558,N_560,N_948);
or U1559 (N_1559,N_619,N_36);
nor U1560 (N_1560,N_379,N_283);
nor U1561 (N_1561,N_552,N_415);
or U1562 (N_1562,N_637,N_15);
nand U1563 (N_1563,N_69,N_489);
xor U1564 (N_1564,N_875,N_467);
or U1565 (N_1565,N_939,N_510);
nand U1566 (N_1566,N_159,N_87);
and U1567 (N_1567,N_319,N_3);
or U1568 (N_1568,N_963,N_955);
nor U1569 (N_1569,N_581,N_323);
nor U1570 (N_1570,N_927,N_280);
or U1571 (N_1571,N_29,N_7);
nand U1572 (N_1572,N_239,N_517);
or U1573 (N_1573,N_233,N_280);
nor U1574 (N_1574,N_926,N_404);
or U1575 (N_1575,N_63,N_808);
nand U1576 (N_1576,N_729,N_499);
nor U1577 (N_1577,N_899,N_582);
nor U1578 (N_1578,N_942,N_846);
and U1579 (N_1579,N_255,N_94);
nor U1580 (N_1580,N_846,N_399);
nand U1581 (N_1581,N_349,N_289);
xnor U1582 (N_1582,N_787,N_273);
nand U1583 (N_1583,N_437,N_40);
nor U1584 (N_1584,N_429,N_418);
or U1585 (N_1585,N_554,N_828);
nor U1586 (N_1586,N_337,N_575);
nand U1587 (N_1587,N_689,N_670);
nor U1588 (N_1588,N_603,N_479);
and U1589 (N_1589,N_581,N_47);
nor U1590 (N_1590,N_221,N_748);
nand U1591 (N_1591,N_846,N_55);
and U1592 (N_1592,N_56,N_282);
and U1593 (N_1593,N_805,N_607);
xnor U1594 (N_1594,N_256,N_884);
and U1595 (N_1595,N_522,N_481);
nand U1596 (N_1596,N_524,N_945);
xnor U1597 (N_1597,N_235,N_621);
and U1598 (N_1598,N_313,N_891);
nor U1599 (N_1599,N_790,N_826);
nand U1600 (N_1600,N_589,N_58);
or U1601 (N_1601,N_851,N_616);
nor U1602 (N_1602,N_208,N_634);
nor U1603 (N_1603,N_250,N_65);
nand U1604 (N_1604,N_575,N_277);
nand U1605 (N_1605,N_637,N_460);
and U1606 (N_1606,N_235,N_182);
or U1607 (N_1607,N_896,N_574);
or U1608 (N_1608,N_25,N_989);
or U1609 (N_1609,N_585,N_677);
and U1610 (N_1610,N_894,N_992);
nand U1611 (N_1611,N_964,N_490);
or U1612 (N_1612,N_47,N_168);
or U1613 (N_1613,N_996,N_901);
nand U1614 (N_1614,N_332,N_670);
or U1615 (N_1615,N_538,N_94);
and U1616 (N_1616,N_259,N_770);
nor U1617 (N_1617,N_194,N_322);
nand U1618 (N_1618,N_937,N_370);
nand U1619 (N_1619,N_872,N_44);
nor U1620 (N_1620,N_92,N_303);
nand U1621 (N_1621,N_946,N_574);
or U1622 (N_1622,N_988,N_236);
nor U1623 (N_1623,N_490,N_924);
nand U1624 (N_1624,N_151,N_91);
or U1625 (N_1625,N_868,N_234);
nand U1626 (N_1626,N_714,N_134);
nand U1627 (N_1627,N_65,N_994);
xnor U1628 (N_1628,N_527,N_884);
nor U1629 (N_1629,N_912,N_345);
and U1630 (N_1630,N_81,N_270);
nand U1631 (N_1631,N_899,N_309);
nor U1632 (N_1632,N_270,N_76);
or U1633 (N_1633,N_746,N_568);
and U1634 (N_1634,N_767,N_305);
or U1635 (N_1635,N_78,N_463);
nor U1636 (N_1636,N_447,N_711);
or U1637 (N_1637,N_308,N_231);
or U1638 (N_1638,N_545,N_771);
xor U1639 (N_1639,N_514,N_643);
nor U1640 (N_1640,N_22,N_187);
and U1641 (N_1641,N_631,N_505);
nor U1642 (N_1642,N_698,N_349);
or U1643 (N_1643,N_176,N_168);
nand U1644 (N_1644,N_765,N_641);
nor U1645 (N_1645,N_699,N_636);
and U1646 (N_1646,N_31,N_315);
and U1647 (N_1647,N_830,N_718);
nand U1648 (N_1648,N_455,N_160);
nand U1649 (N_1649,N_152,N_189);
and U1650 (N_1650,N_747,N_535);
nand U1651 (N_1651,N_192,N_959);
xor U1652 (N_1652,N_781,N_633);
or U1653 (N_1653,N_18,N_225);
nand U1654 (N_1654,N_570,N_573);
xor U1655 (N_1655,N_175,N_700);
xor U1656 (N_1656,N_941,N_237);
nor U1657 (N_1657,N_816,N_942);
nor U1658 (N_1658,N_724,N_823);
nand U1659 (N_1659,N_390,N_604);
or U1660 (N_1660,N_188,N_343);
nand U1661 (N_1661,N_969,N_189);
nor U1662 (N_1662,N_439,N_202);
and U1663 (N_1663,N_196,N_607);
nor U1664 (N_1664,N_221,N_826);
and U1665 (N_1665,N_40,N_87);
nand U1666 (N_1666,N_120,N_225);
nor U1667 (N_1667,N_488,N_477);
or U1668 (N_1668,N_357,N_713);
and U1669 (N_1669,N_106,N_423);
and U1670 (N_1670,N_856,N_120);
or U1671 (N_1671,N_279,N_959);
or U1672 (N_1672,N_307,N_967);
nor U1673 (N_1673,N_588,N_1);
or U1674 (N_1674,N_95,N_277);
nand U1675 (N_1675,N_596,N_486);
and U1676 (N_1676,N_585,N_244);
and U1677 (N_1677,N_123,N_207);
xnor U1678 (N_1678,N_647,N_115);
and U1679 (N_1679,N_608,N_860);
nor U1680 (N_1680,N_640,N_154);
xnor U1681 (N_1681,N_764,N_976);
nor U1682 (N_1682,N_721,N_447);
nor U1683 (N_1683,N_639,N_161);
xor U1684 (N_1684,N_814,N_329);
or U1685 (N_1685,N_724,N_519);
or U1686 (N_1686,N_712,N_26);
or U1687 (N_1687,N_24,N_687);
nand U1688 (N_1688,N_954,N_893);
nor U1689 (N_1689,N_81,N_206);
or U1690 (N_1690,N_486,N_2);
or U1691 (N_1691,N_612,N_85);
or U1692 (N_1692,N_492,N_713);
nor U1693 (N_1693,N_321,N_228);
and U1694 (N_1694,N_356,N_92);
nand U1695 (N_1695,N_682,N_460);
nand U1696 (N_1696,N_540,N_506);
xor U1697 (N_1697,N_437,N_310);
nor U1698 (N_1698,N_486,N_956);
xnor U1699 (N_1699,N_591,N_12);
and U1700 (N_1700,N_297,N_482);
nor U1701 (N_1701,N_768,N_431);
nor U1702 (N_1702,N_763,N_20);
xnor U1703 (N_1703,N_309,N_70);
and U1704 (N_1704,N_881,N_884);
and U1705 (N_1705,N_628,N_91);
or U1706 (N_1706,N_314,N_741);
and U1707 (N_1707,N_708,N_589);
and U1708 (N_1708,N_91,N_950);
or U1709 (N_1709,N_360,N_672);
and U1710 (N_1710,N_254,N_573);
nor U1711 (N_1711,N_279,N_29);
nor U1712 (N_1712,N_914,N_82);
nand U1713 (N_1713,N_432,N_277);
or U1714 (N_1714,N_866,N_540);
xnor U1715 (N_1715,N_11,N_403);
nor U1716 (N_1716,N_558,N_813);
nand U1717 (N_1717,N_152,N_253);
nor U1718 (N_1718,N_143,N_255);
and U1719 (N_1719,N_459,N_871);
nand U1720 (N_1720,N_371,N_363);
or U1721 (N_1721,N_461,N_825);
nand U1722 (N_1722,N_978,N_838);
and U1723 (N_1723,N_145,N_142);
and U1724 (N_1724,N_531,N_902);
nor U1725 (N_1725,N_104,N_391);
xnor U1726 (N_1726,N_662,N_109);
nor U1727 (N_1727,N_881,N_458);
nor U1728 (N_1728,N_229,N_7);
nand U1729 (N_1729,N_291,N_803);
nor U1730 (N_1730,N_320,N_105);
nand U1731 (N_1731,N_223,N_289);
or U1732 (N_1732,N_594,N_595);
nor U1733 (N_1733,N_384,N_295);
nor U1734 (N_1734,N_693,N_158);
xor U1735 (N_1735,N_118,N_577);
and U1736 (N_1736,N_980,N_223);
and U1737 (N_1737,N_295,N_917);
and U1738 (N_1738,N_620,N_466);
nand U1739 (N_1739,N_703,N_188);
nand U1740 (N_1740,N_34,N_141);
nor U1741 (N_1741,N_757,N_766);
and U1742 (N_1742,N_270,N_350);
nor U1743 (N_1743,N_925,N_210);
and U1744 (N_1744,N_987,N_260);
or U1745 (N_1745,N_348,N_952);
nor U1746 (N_1746,N_869,N_649);
and U1747 (N_1747,N_144,N_830);
or U1748 (N_1748,N_658,N_746);
nor U1749 (N_1749,N_764,N_54);
nand U1750 (N_1750,N_24,N_96);
nand U1751 (N_1751,N_188,N_546);
nand U1752 (N_1752,N_816,N_365);
nor U1753 (N_1753,N_433,N_82);
or U1754 (N_1754,N_639,N_764);
or U1755 (N_1755,N_916,N_909);
and U1756 (N_1756,N_487,N_721);
xnor U1757 (N_1757,N_248,N_451);
and U1758 (N_1758,N_408,N_37);
xor U1759 (N_1759,N_368,N_403);
and U1760 (N_1760,N_268,N_721);
and U1761 (N_1761,N_569,N_490);
and U1762 (N_1762,N_32,N_165);
or U1763 (N_1763,N_796,N_219);
and U1764 (N_1764,N_596,N_584);
xor U1765 (N_1765,N_216,N_125);
and U1766 (N_1766,N_472,N_682);
nand U1767 (N_1767,N_483,N_355);
and U1768 (N_1768,N_555,N_594);
or U1769 (N_1769,N_499,N_560);
nor U1770 (N_1770,N_319,N_671);
or U1771 (N_1771,N_588,N_928);
and U1772 (N_1772,N_687,N_267);
or U1773 (N_1773,N_425,N_454);
nand U1774 (N_1774,N_969,N_39);
or U1775 (N_1775,N_839,N_564);
and U1776 (N_1776,N_570,N_484);
nor U1777 (N_1777,N_889,N_489);
xor U1778 (N_1778,N_487,N_795);
and U1779 (N_1779,N_569,N_188);
or U1780 (N_1780,N_269,N_938);
nand U1781 (N_1781,N_458,N_457);
nor U1782 (N_1782,N_827,N_746);
and U1783 (N_1783,N_230,N_246);
or U1784 (N_1784,N_48,N_598);
and U1785 (N_1785,N_532,N_285);
nor U1786 (N_1786,N_672,N_643);
xnor U1787 (N_1787,N_371,N_214);
nand U1788 (N_1788,N_974,N_102);
nor U1789 (N_1789,N_302,N_475);
xnor U1790 (N_1790,N_759,N_736);
and U1791 (N_1791,N_402,N_224);
nand U1792 (N_1792,N_225,N_561);
and U1793 (N_1793,N_652,N_186);
nor U1794 (N_1794,N_844,N_268);
or U1795 (N_1795,N_859,N_251);
or U1796 (N_1796,N_526,N_946);
and U1797 (N_1797,N_815,N_490);
nor U1798 (N_1798,N_107,N_679);
nand U1799 (N_1799,N_644,N_834);
nor U1800 (N_1800,N_995,N_670);
nor U1801 (N_1801,N_856,N_942);
and U1802 (N_1802,N_967,N_749);
nor U1803 (N_1803,N_4,N_76);
nand U1804 (N_1804,N_301,N_633);
xnor U1805 (N_1805,N_890,N_617);
and U1806 (N_1806,N_38,N_74);
or U1807 (N_1807,N_190,N_342);
or U1808 (N_1808,N_397,N_687);
nand U1809 (N_1809,N_800,N_275);
nand U1810 (N_1810,N_46,N_399);
nor U1811 (N_1811,N_399,N_733);
nand U1812 (N_1812,N_904,N_82);
nand U1813 (N_1813,N_992,N_614);
or U1814 (N_1814,N_10,N_562);
xnor U1815 (N_1815,N_770,N_192);
nor U1816 (N_1816,N_197,N_866);
and U1817 (N_1817,N_113,N_355);
nor U1818 (N_1818,N_552,N_812);
nor U1819 (N_1819,N_989,N_447);
or U1820 (N_1820,N_606,N_423);
nand U1821 (N_1821,N_333,N_574);
and U1822 (N_1822,N_139,N_612);
and U1823 (N_1823,N_681,N_563);
xor U1824 (N_1824,N_223,N_455);
nand U1825 (N_1825,N_406,N_760);
or U1826 (N_1826,N_812,N_768);
nor U1827 (N_1827,N_679,N_986);
or U1828 (N_1828,N_796,N_137);
xnor U1829 (N_1829,N_569,N_680);
nand U1830 (N_1830,N_966,N_472);
xnor U1831 (N_1831,N_951,N_599);
nor U1832 (N_1832,N_472,N_524);
nor U1833 (N_1833,N_566,N_689);
or U1834 (N_1834,N_734,N_503);
or U1835 (N_1835,N_663,N_802);
nand U1836 (N_1836,N_111,N_671);
and U1837 (N_1837,N_852,N_652);
or U1838 (N_1838,N_41,N_103);
nand U1839 (N_1839,N_454,N_885);
nor U1840 (N_1840,N_886,N_543);
or U1841 (N_1841,N_684,N_894);
or U1842 (N_1842,N_139,N_504);
nor U1843 (N_1843,N_260,N_565);
and U1844 (N_1844,N_150,N_67);
and U1845 (N_1845,N_736,N_581);
and U1846 (N_1846,N_26,N_629);
nand U1847 (N_1847,N_781,N_326);
nor U1848 (N_1848,N_348,N_663);
nor U1849 (N_1849,N_898,N_452);
or U1850 (N_1850,N_747,N_614);
and U1851 (N_1851,N_115,N_968);
or U1852 (N_1852,N_617,N_502);
nand U1853 (N_1853,N_22,N_441);
and U1854 (N_1854,N_495,N_171);
nor U1855 (N_1855,N_7,N_371);
or U1856 (N_1856,N_340,N_70);
nor U1857 (N_1857,N_906,N_777);
nor U1858 (N_1858,N_536,N_893);
nand U1859 (N_1859,N_891,N_667);
nand U1860 (N_1860,N_886,N_964);
nor U1861 (N_1861,N_586,N_241);
nor U1862 (N_1862,N_778,N_777);
nand U1863 (N_1863,N_708,N_369);
nor U1864 (N_1864,N_218,N_855);
nand U1865 (N_1865,N_18,N_270);
nor U1866 (N_1866,N_766,N_13);
nor U1867 (N_1867,N_475,N_71);
and U1868 (N_1868,N_925,N_752);
and U1869 (N_1869,N_869,N_264);
or U1870 (N_1870,N_957,N_897);
nand U1871 (N_1871,N_697,N_489);
or U1872 (N_1872,N_433,N_202);
or U1873 (N_1873,N_536,N_187);
or U1874 (N_1874,N_437,N_268);
nand U1875 (N_1875,N_53,N_713);
or U1876 (N_1876,N_145,N_529);
nor U1877 (N_1877,N_543,N_112);
nand U1878 (N_1878,N_308,N_295);
nor U1879 (N_1879,N_896,N_373);
xor U1880 (N_1880,N_365,N_703);
nand U1881 (N_1881,N_155,N_539);
or U1882 (N_1882,N_457,N_378);
nand U1883 (N_1883,N_509,N_695);
nand U1884 (N_1884,N_653,N_673);
nor U1885 (N_1885,N_884,N_80);
nor U1886 (N_1886,N_813,N_615);
nor U1887 (N_1887,N_746,N_761);
and U1888 (N_1888,N_19,N_665);
nor U1889 (N_1889,N_167,N_893);
nand U1890 (N_1890,N_840,N_325);
and U1891 (N_1891,N_933,N_563);
and U1892 (N_1892,N_21,N_270);
nand U1893 (N_1893,N_711,N_451);
or U1894 (N_1894,N_191,N_403);
xor U1895 (N_1895,N_670,N_768);
nand U1896 (N_1896,N_986,N_891);
and U1897 (N_1897,N_14,N_952);
nand U1898 (N_1898,N_185,N_828);
nor U1899 (N_1899,N_225,N_360);
or U1900 (N_1900,N_757,N_454);
xor U1901 (N_1901,N_264,N_899);
xor U1902 (N_1902,N_924,N_600);
nor U1903 (N_1903,N_357,N_983);
and U1904 (N_1904,N_962,N_385);
and U1905 (N_1905,N_660,N_665);
nand U1906 (N_1906,N_650,N_11);
or U1907 (N_1907,N_585,N_218);
nand U1908 (N_1908,N_12,N_914);
nand U1909 (N_1909,N_845,N_620);
and U1910 (N_1910,N_141,N_661);
nor U1911 (N_1911,N_417,N_507);
nand U1912 (N_1912,N_687,N_518);
nand U1913 (N_1913,N_734,N_660);
and U1914 (N_1914,N_254,N_983);
nand U1915 (N_1915,N_623,N_14);
nand U1916 (N_1916,N_174,N_58);
or U1917 (N_1917,N_254,N_616);
or U1918 (N_1918,N_290,N_355);
nor U1919 (N_1919,N_464,N_800);
and U1920 (N_1920,N_220,N_602);
or U1921 (N_1921,N_453,N_649);
nand U1922 (N_1922,N_298,N_111);
and U1923 (N_1923,N_682,N_401);
nand U1924 (N_1924,N_13,N_759);
nor U1925 (N_1925,N_481,N_65);
nor U1926 (N_1926,N_203,N_780);
or U1927 (N_1927,N_723,N_945);
and U1928 (N_1928,N_242,N_139);
or U1929 (N_1929,N_817,N_657);
xor U1930 (N_1930,N_726,N_457);
and U1931 (N_1931,N_204,N_286);
or U1932 (N_1932,N_14,N_739);
xnor U1933 (N_1933,N_808,N_117);
nor U1934 (N_1934,N_128,N_667);
or U1935 (N_1935,N_358,N_660);
nand U1936 (N_1936,N_87,N_766);
or U1937 (N_1937,N_713,N_774);
nand U1938 (N_1938,N_919,N_871);
xor U1939 (N_1939,N_542,N_787);
nand U1940 (N_1940,N_236,N_456);
xnor U1941 (N_1941,N_960,N_298);
and U1942 (N_1942,N_634,N_437);
and U1943 (N_1943,N_76,N_261);
or U1944 (N_1944,N_201,N_190);
nor U1945 (N_1945,N_942,N_397);
nand U1946 (N_1946,N_741,N_368);
xnor U1947 (N_1947,N_532,N_372);
nand U1948 (N_1948,N_726,N_809);
and U1949 (N_1949,N_214,N_194);
nor U1950 (N_1950,N_302,N_395);
nand U1951 (N_1951,N_509,N_144);
or U1952 (N_1952,N_159,N_103);
nand U1953 (N_1953,N_260,N_501);
or U1954 (N_1954,N_860,N_913);
nand U1955 (N_1955,N_95,N_107);
xnor U1956 (N_1956,N_974,N_259);
and U1957 (N_1957,N_694,N_641);
nand U1958 (N_1958,N_829,N_214);
nor U1959 (N_1959,N_613,N_624);
and U1960 (N_1960,N_341,N_653);
nand U1961 (N_1961,N_357,N_489);
nor U1962 (N_1962,N_239,N_846);
and U1963 (N_1963,N_721,N_818);
nand U1964 (N_1964,N_225,N_41);
nor U1965 (N_1965,N_447,N_962);
and U1966 (N_1966,N_780,N_595);
nor U1967 (N_1967,N_396,N_695);
and U1968 (N_1968,N_741,N_846);
nand U1969 (N_1969,N_415,N_500);
or U1970 (N_1970,N_417,N_720);
or U1971 (N_1971,N_750,N_556);
and U1972 (N_1972,N_854,N_116);
nand U1973 (N_1973,N_2,N_363);
or U1974 (N_1974,N_762,N_839);
nand U1975 (N_1975,N_932,N_883);
or U1976 (N_1976,N_149,N_980);
nand U1977 (N_1977,N_207,N_96);
nand U1978 (N_1978,N_124,N_309);
or U1979 (N_1979,N_381,N_127);
nand U1980 (N_1980,N_58,N_944);
and U1981 (N_1981,N_909,N_204);
nor U1982 (N_1982,N_279,N_465);
xnor U1983 (N_1983,N_649,N_486);
and U1984 (N_1984,N_934,N_641);
and U1985 (N_1985,N_620,N_560);
nor U1986 (N_1986,N_657,N_810);
or U1987 (N_1987,N_641,N_881);
nand U1988 (N_1988,N_585,N_833);
nand U1989 (N_1989,N_168,N_579);
or U1990 (N_1990,N_805,N_19);
nor U1991 (N_1991,N_400,N_895);
or U1992 (N_1992,N_990,N_544);
or U1993 (N_1993,N_595,N_149);
nand U1994 (N_1994,N_993,N_417);
nand U1995 (N_1995,N_19,N_615);
nor U1996 (N_1996,N_507,N_176);
or U1997 (N_1997,N_284,N_990);
nor U1998 (N_1998,N_174,N_214);
nand U1999 (N_1999,N_695,N_263);
and U2000 (N_2000,N_1835,N_1008);
nand U2001 (N_2001,N_1958,N_1720);
or U2002 (N_2002,N_1453,N_1095);
and U2003 (N_2003,N_1175,N_1595);
nor U2004 (N_2004,N_1754,N_1474);
or U2005 (N_2005,N_1235,N_1361);
nor U2006 (N_2006,N_1023,N_1108);
nor U2007 (N_2007,N_1421,N_1811);
nor U2008 (N_2008,N_1910,N_1204);
xor U2009 (N_2009,N_1368,N_1469);
and U2010 (N_2010,N_1858,N_1410);
nand U2011 (N_2011,N_1669,N_1889);
xnor U2012 (N_2012,N_1647,N_1945);
nand U2013 (N_2013,N_1930,N_1164);
and U2014 (N_2014,N_1168,N_1545);
and U2015 (N_2015,N_1067,N_1020);
nor U2016 (N_2016,N_1553,N_1846);
nand U2017 (N_2017,N_1541,N_1145);
nor U2018 (N_2018,N_1329,N_1941);
and U2019 (N_2019,N_1154,N_1908);
nand U2020 (N_2020,N_1507,N_1265);
nand U2021 (N_2021,N_1977,N_1755);
or U2022 (N_2022,N_1136,N_1639);
nor U2023 (N_2023,N_1686,N_1261);
xnor U2024 (N_2024,N_1853,N_1981);
or U2025 (N_2025,N_1491,N_1335);
or U2026 (N_2026,N_1216,N_1707);
or U2027 (N_2027,N_1670,N_1221);
nand U2028 (N_2028,N_1691,N_1439);
nand U2029 (N_2029,N_1867,N_1949);
xor U2030 (N_2030,N_1354,N_1071);
nand U2031 (N_2031,N_1940,N_1304);
or U2032 (N_2032,N_1400,N_1752);
and U2033 (N_2033,N_1231,N_1386);
nand U2034 (N_2034,N_1543,N_1785);
and U2035 (N_2035,N_1339,N_1897);
xnor U2036 (N_2036,N_1583,N_1925);
nor U2037 (N_2037,N_1655,N_1570);
and U2038 (N_2038,N_1320,N_1159);
nand U2039 (N_2039,N_1688,N_1578);
and U2040 (N_2040,N_1392,N_1419);
and U2041 (N_2041,N_1523,N_1267);
nor U2042 (N_2042,N_1012,N_1475);
or U2043 (N_2043,N_1600,N_1073);
or U2044 (N_2044,N_1103,N_1764);
nand U2045 (N_2045,N_1555,N_1114);
or U2046 (N_2046,N_1081,N_1378);
xor U2047 (N_2047,N_1139,N_1602);
nor U2048 (N_2048,N_1040,N_1127);
nor U2049 (N_2049,N_1591,N_1466);
nand U2050 (N_2050,N_1129,N_1879);
xor U2051 (N_2051,N_1025,N_1328);
and U2052 (N_2052,N_1573,N_1263);
nor U2053 (N_2053,N_1758,N_1124);
nand U2054 (N_2054,N_1151,N_1483);
nor U2055 (N_2055,N_1805,N_1515);
nand U2056 (N_2056,N_1778,N_1671);
or U2057 (N_2057,N_1633,N_1131);
nand U2058 (N_2058,N_1285,N_1387);
nor U2059 (N_2059,N_1196,N_1169);
and U2060 (N_2060,N_1975,N_1849);
nand U2061 (N_2061,N_1119,N_1253);
xor U2062 (N_2062,N_1607,N_1412);
or U2063 (N_2063,N_1834,N_1195);
nand U2064 (N_2064,N_1123,N_1465);
xnor U2065 (N_2065,N_1097,N_1799);
nand U2066 (N_2066,N_1251,N_1870);
xnor U2067 (N_2067,N_1919,N_1110);
and U2068 (N_2068,N_1309,N_1894);
nand U2069 (N_2069,N_1384,N_1260);
and U2070 (N_2070,N_1035,N_1153);
nand U2071 (N_2071,N_1830,N_1488);
nand U2072 (N_2072,N_1257,N_1068);
or U2073 (N_2073,N_1186,N_1030);
and U2074 (N_2074,N_1855,N_1616);
nor U2075 (N_2075,N_1118,N_1715);
nand U2076 (N_2076,N_1113,N_1874);
xor U2077 (N_2077,N_1604,N_1721);
nor U2078 (N_2078,N_1943,N_1682);
nor U2079 (N_2079,N_1821,N_1926);
nand U2080 (N_2080,N_1418,N_1240);
or U2081 (N_2081,N_1818,N_1214);
xnor U2082 (N_2082,N_1497,N_1057);
and U2083 (N_2083,N_1819,N_1988);
or U2084 (N_2084,N_1652,N_1447);
or U2085 (N_2085,N_1225,N_1202);
or U2086 (N_2086,N_1581,N_1401);
and U2087 (N_2087,N_1531,N_1058);
or U2088 (N_2088,N_1489,N_1224);
or U2089 (N_2089,N_1615,N_1403);
nor U2090 (N_2090,N_1314,N_1163);
xor U2091 (N_2091,N_1559,N_1112);
or U2092 (N_2092,N_1801,N_1086);
nor U2093 (N_2093,N_1413,N_1406);
nand U2094 (N_2094,N_1603,N_1551);
and U2095 (N_2095,N_1579,N_1964);
and U2096 (N_2096,N_1959,N_1997);
or U2097 (N_2097,N_1606,N_1311);
nor U2098 (N_2098,N_1457,N_1428);
xor U2099 (N_2099,N_1229,N_1994);
nand U2100 (N_2100,N_1634,N_1310);
or U2101 (N_2101,N_1006,N_1954);
and U2102 (N_2102,N_1967,N_1768);
and U2103 (N_2103,N_1415,N_1293);
xor U2104 (N_2104,N_1459,N_1336);
and U2105 (N_2105,N_1382,N_1659);
or U2106 (N_2106,N_1034,N_1101);
or U2107 (N_2107,N_1674,N_1672);
nor U2108 (N_2108,N_1243,N_1269);
nand U2109 (N_2109,N_1582,N_1249);
or U2110 (N_2110,N_1019,N_1083);
nor U2111 (N_2111,N_1362,N_1769);
nor U2112 (N_2112,N_1286,N_1150);
and U2113 (N_2113,N_1003,N_1741);
or U2114 (N_2114,N_1653,N_1301);
nor U2115 (N_2115,N_1203,N_1612);
nand U2116 (N_2116,N_1143,N_1632);
nand U2117 (N_2117,N_1275,N_1585);
or U2118 (N_2118,N_1179,N_1623);
nand U2119 (N_2119,N_1167,N_1201);
nor U2120 (N_2120,N_1004,N_1147);
nor U2121 (N_2121,N_1353,N_1845);
nor U2122 (N_2122,N_1347,N_1077);
or U2123 (N_2123,N_1341,N_1728);
and U2124 (N_2124,N_1844,N_1296);
nor U2125 (N_2125,N_1274,N_1241);
xnor U2126 (N_2126,N_1084,N_1098);
or U2127 (N_2127,N_1505,N_1213);
xnor U2128 (N_2128,N_1132,N_1529);
nand U2129 (N_2129,N_1970,N_1363);
or U2130 (N_2130,N_1899,N_1405);
xor U2131 (N_2131,N_1770,N_1714);
and U2132 (N_2132,N_1370,N_1727);
or U2133 (N_2133,N_1436,N_1513);
nand U2134 (N_2134,N_1776,N_1443);
nor U2135 (N_2135,N_1588,N_1010);
or U2136 (N_2136,N_1978,N_1598);
nor U2137 (N_2137,N_1495,N_1510);
nor U2138 (N_2138,N_1944,N_1539);
nand U2139 (N_2139,N_1451,N_1237);
and U2140 (N_2140,N_1712,N_1115);
nor U2141 (N_2141,N_1589,N_1059);
nand U2142 (N_2142,N_1854,N_1654);
nor U2143 (N_2143,N_1885,N_1478);
nand U2144 (N_2144,N_1393,N_1868);
nand U2145 (N_2145,N_1924,N_1972);
nor U2146 (N_2146,N_1360,N_1255);
nand U2147 (N_2147,N_1839,N_1399);
nand U2148 (N_2148,N_1548,N_1259);
or U2149 (N_2149,N_1638,N_1450);
nand U2150 (N_2150,N_1961,N_1575);
or U2151 (N_2151,N_1998,N_1174);
nor U2152 (N_2152,N_1248,N_1048);
nor U2153 (N_2153,N_1376,N_1391);
and U2154 (N_2154,N_1773,N_1002);
nor U2155 (N_2155,N_1487,N_1508);
nand U2156 (N_2156,N_1909,N_1383);
xor U2157 (N_2157,N_1367,N_1802);
or U2158 (N_2158,N_1976,N_1394);
nor U2159 (N_2159,N_1512,N_1927);
and U2160 (N_2160,N_1463,N_1054);
or U2161 (N_2161,N_1321,N_1324);
xor U2162 (N_2162,N_1922,N_1611);
xnor U2163 (N_2163,N_1697,N_1571);
or U2164 (N_2164,N_1526,N_1883);
and U2165 (N_2165,N_1683,N_1540);
nor U2166 (N_2166,N_1562,N_1481);
and U2167 (N_2167,N_1678,N_1303);
nor U2168 (N_2168,N_1847,N_1856);
nor U2169 (N_2169,N_1080,N_1056);
nand U2170 (N_2170,N_1902,N_1871);
nand U2171 (N_2171,N_1733,N_1695);
nand U2172 (N_2172,N_1706,N_1280);
nand U2173 (N_2173,N_1781,N_1432);
or U2174 (N_2174,N_1624,N_1290);
or U2175 (N_2175,N_1843,N_1992);
xnor U2176 (N_2176,N_1137,N_1864);
nor U2177 (N_2177,N_1026,N_1504);
nand U2178 (N_2178,N_1534,N_1128);
nor U2179 (N_2179,N_1130,N_1857);
nand U2180 (N_2180,N_1957,N_1337);
nor U2181 (N_2181,N_1527,N_1979);
or U2182 (N_2182,N_1066,N_1190);
nand U2183 (N_2183,N_1182,N_1788);
or U2184 (N_2184,N_1605,N_1178);
nor U2185 (N_2185,N_1055,N_1111);
and U2186 (N_2186,N_1028,N_1456);
nor U2187 (N_2187,N_1094,N_1484);
nand U2188 (N_2188,N_1158,N_1537);
and U2189 (N_2189,N_1172,N_1519);
xor U2190 (N_2190,N_1312,N_1787);
and U2191 (N_2191,N_1593,N_1913);
and U2192 (N_2192,N_1656,N_1013);
or U2193 (N_2193,N_1380,N_1905);
or U2194 (N_2194,N_1062,N_1138);
and U2195 (N_2195,N_1051,N_1171);
and U2196 (N_2196,N_1866,N_1516);
nand U2197 (N_2197,N_1011,N_1955);
nor U2198 (N_2198,N_1668,N_1236);
and U2199 (N_2199,N_1891,N_1798);
or U2200 (N_2200,N_1993,N_1677);
nor U2201 (N_2201,N_1794,N_1226);
xnor U2202 (N_2202,N_1087,N_1359);
xor U2203 (N_2203,N_1365,N_1522);
nand U2204 (N_2204,N_1528,N_1152);
nand U2205 (N_2205,N_1468,N_1185);
nand U2206 (N_2206,N_1631,N_1476);
xnor U2207 (N_2207,N_1968,N_1765);
nor U2208 (N_2208,N_1509,N_1822);
and U2209 (N_2209,N_1831,N_1708);
or U2210 (N_2210,N_1161,N_1414);
nand U2211 (N_2211,N_1936,N_1282);
nor U2212 (N_2212,N_1660,N_1210);
nor U2213 (N_2213,N_1829,N_1751);
or U2214 (N_2214,N_1090,N_1971);
and U2215 (N_2215,N_1338,N_1791);
and U2216 (N_2216,N_1731,N_1999);
and U2217 (N_2217,N_1180,N_1800);
xnor U2218 (N_2218,N_1460,N_1824);
nor U2219 (N_2219,N_1326,N_1219);
or U2220 (N_2220,N_1379,N_1861);
and U2221 (N_2221,N_1395,N_1350);
or U2222 (N_2222,N_1449,N_1875);
nand U2223 (N_2223,N_1334,N_1141);
and U2224 (N_2224,N_1547,N_1100);
nand U2225 (N_2225,N_1735,N_1356);
nand U2226 (N_2226,N_1932,N_1506);
or U2227 (N_2227,N_1223,N_1895);
or U2228 (N_2228,N_1825,N_1782);
nor U2229 (N_2229,N_1815,N_1315);
nor U2230 (N_2230,N_1601,N_1796);
xor U2231 (N_2231,N_1502,N_1610);
nor U2232 (N_2232,N_1766,N_1763);
xnor U2233 (N_2233,N_1740,N_1292);
nor U2234 (N_2234,N_1031,N_1279);
or U2235 (N_2235,N_1121,N_1166);
nor U2236 (N_2236,N_1746,N_1646);
or U2237 (N_2237,N_1809,N_1572);
or U2238 (N_2238,N_1725,N_1703);
nand U2239 (N_2239,N_1916,N_1117);
nor U2240 (N_2240,N_1577,N_1629);
or U2241 (N_2241,N_1014,N_1467);
nor U2242 (N_2242,N_1783,N_1276);
or U2243 (N_2243,N_1357,N_1064);
nor U2244 (N_2244,N_1142,N_1107);
nor U2245 (N_2245,N_1650,N_1409);
xnor U2246 (N_2246,N_1156,N_1348);
nand U2247 (N_2247,N_1774,N_1877);
nor U2248 (N_2248,N_1973,N_1744);
and U2249 (N_2249,N_1907,N_1584);
nor U2250 (N_2250,N_1761,N_1881);
or U2251 (N_2251,N_1896,N_1912);
nor U2252 (N_2252,N_1024,N_1254);
nor U2253 (N_2253,N_1300,N_1184);
nor U2254 (N_2254,N_1250,N_1162);
xnor U2255 (N_2255,N_1425,N_1188);
nor U2256 (N_2256,N_1649,N_1745);
nand U2257 (N_2257,N_1288,N_1037);
nor U2258 (N_2258,N_1832,N_1814);
nor U2259 (N_2259,N_1893,N_1092);
and U2260 (N_2260,N_1284,N_1810);
and U2261 (N_2261,N_1189,N_1287);
nand U2262 (N_2262,N_1327,N_1762);
nor U2263 (N_2263,N_1619,N_1760);
and U2264 (N_2264,N_1576,N_1352);
nor U2265 (N_2265,N_1542,N_1369);
or U2266 (N_2266,N_1699,N_1613);
xnor U2267 (N_2267,N_1625,N_1749);
nand U2268 (N_2268,N_1797,N_1828);
nand U2269 (N_2269,N_1396,N_1313);
nor U2270 (N_2270,N_1717,N_1305);
or U2271 (N_2271,N_1433,N_1272);
and U2272 (N_2272,N_1739,N_1549);
or U2273 (N_2273,N_1344,N_1206);
nor U2274 (N_2274,N_1455,N_1429);
nor U2275 (N_2275,N_1345,N_1618);
and U2276 (N_2276,N_1452,N_1804);
and U2277 (N_2277,N_1586,N_1397);
and U2278 (N_2278,N_1085,N_1298);
or U2279 (N_2279,N_1351,N_1730);
nand U2280 (N_2280,N_1742,N_1530);
nand U2281 (N_2281,N_1914,N_1738);
xnor U2282 (N_2282,N_1535,N_1050);
nand U2283 (N_2283,N_1795,N_1297);
nor U2284 (N_2284,N_1060,N_1388);
nor U2285 (N_2285,N_1042,N_1679);
nor U2286 (N_2286,N_1713,N_1826);
or U2287 (N_2287,N_1722,N_1183);
or U2288 (N_2288,N_1375,N_1473);
nor U2289 (N_2289,N_1817,N_1173);
nand U2290 (N_2290,N_1317,N_1374);
or U2291 (N_2291,N_1022,N_1330);
nand U2292 (N_2292,N_1748,N_1533);
or U2293 (N_2293,N_1590,N_1675);
nor U2294 (N_2294,N_1962,N_1233);
nand U2295 (N_2295,N_1033,N_1892);
or U2296 (N_2296,N_1245,N_1833);
and U2297 (N_2297,N_1876,N_1685);
nand U2298 (N_2298,N_1482,N_1995);
or U2299 (N_2299,N_1934,N_1015);
nor U2300 (N_2300,N_1270,N_1718);
nand U2301 (N_2301,N_1385,N_1041);
nor U2302 (N_2302,N_1753,N_1120);
nor U2303 (N_2303,N_1990,N_1258);
nand U2304 (N_2304,N_1942,N_1209);
nand U2305 (N_2305,N_1594,N_1125);
and U2306 (N_2306,N_1364,N_1283);
nand U2307 (N_2307,N_1492,N_1480);
xnor U2308 (N_2308,N_1786,N_1991);
nor U2309 (N_2309,N_1644,N_1775);
nor U2310 (N_2310,N_1793,N_1426);
nor U2311 (N_2311,N_1464,N_1701);
xor U2312 (N_2312,N_1372,N_1458);
and U2313 (N_2313,N_1651,N_1256);
nor U2314 (N_2314,N_1935,N_1729);
or U2315 (N_2315,N_1886,N_1016);
nand U2316 (N_2316,N_1777,N_1772);
nand U2317 (N_2317,N_1416,N_1716);
and U2318 (N_2318,N_1155,N_1641);
nand U2319 (N_2319,N_1756,N_1663);
nor U2320 (N_2320,N_1937,N_1734);
nand U2321 (N_2321,N_1218,N_1622);
or U2322 (N_2322,N_1342,N_1343);
and U2323 (N_2323,N_1931,N_1518);
and U2324 (N_2324,N_1238,N_1851);
or U2325 (N_2325,N_1318,N_1242);
and U2326 (N_2326,N_1692,N_1036);
nor U2327 (N_2327,N_1278,N_1838);
and U2328 (N_2328,N_1027,N_1207);
or U2329 (N_2329,N_1194,N_1974);
nor U2330 (N_2330,N_1007,N_1234);
and U2331 (N_2331,N_1784,N_1331);
nor U2332 (N_2332,N_1454,N_1091);
or U2333 (N_2333,N_1322,N_1122);
xnor U2334 (N_2334,N_1517,N_1918);
nand U2335 (N_2335,N_1938,N_1863);
nor U2336 (N_2336,N_1486,N_1479);
nor U2337 (N_2337,N_1192,N_1966);
or U2338 (N_2338,N_1608,N_1099);
nor U2339 (N_2339,N_1599,N_1850);
or U2340 (N_2340,N_1664,N_1047);
nor U2341 (N_2341,N_1319,N_1211);
nand U2342 (N_2342,N_1956,N_1227);
and U2343 (N_2343,N_1948,N_1205);
nor U2344 (N_2344,N_1790,N_1951);
nor U2345 (N_2345,N_1157,N_1140);
nor U2346 (N_2346,N_1690,N_1438);
nor U2347 (N_2347,N_1381,N_1032);
or U2348 (N_2348,N_1884,N_1061);
nand U2349 (N_2349,N_1435,N_1643);
and U2350 (N_2350,N_1557,N_1422);
or U2351 (N_2351,N_1440,N_1308);
or U2352 (N_2352,N_1521,N_1018);
xnor U2353 (N_2353,N_1779,N_1597);
nand U2354 (N_2354,N_1009,N_1333);
nand U2355 (N_2355,N_1088,N_1880);
nor U2356 (N_2356,N_1666,N_1001);
nand U2357 (N_2357,N_1273,N_1493);
and U2358 (N_2358,N_1984,N_1355);
nand U2359 (N_2359,N_1038,N_1848);
nand U2360 (N_2360,N_1823,N_1911);
or U2361 (N_2361,N_1808,N_1552);
and U2362 (N_2362,N_1732,N_1053);
nor U2363 (N_2363,N_1719,N_1840);
and U2364 (N_2364,N_1681,N_1498);
or U2365 (N_2365,N_1029,N_1039);
nand U2366 (N_2366,N_1230,N_1000);
nand U2367 (N_2367,N_1462,N_1789);
nand U2368 (N_2368,N_1191,N_1621);
nor U2369 (N_2369,N_1915,N_1694);
nor U2370 (N_2370,N_1228,N_1642);
and U2371 (N_2371,N_1747,N_1524);
and U2372 (N_2372,N_1820,N_1045);
or U2373 (N_2373,N_1427,N_1920);
and U2374 (N_2374,N_1665,N_1323);
or U2375 (N_2375,N_1561,N_1544);
or U2376 (N_2376,N_1176,N_1812);
or U2377 (N_2377,N_1349,N_1430);
and U2378 (N_2378,N_1563,N_1044);
and U2379 (N_2379,N_1700,N_1501);
and U2380 (N_2380,N_1461,N_1662);
and U2381 (N_2381,N_1135,N_1536);
nor U2382 (N_2382,N_1408,N_1837);
or U2383 (N_2383,N_1836,N_1511);
nor U2384 (N_2384,N_1217,N_1208);
xor U2385 (N_2385,N_1596,N_1093);
nand U2386 (N_2386,N_1564,N_1373);
and U2387 (N_2387,N_1133,N_1710);
or U2388 (N_2388,N_1969,N_1950);
and U2389 (N_2389,N_1687,N_1423);
and U2390 (N_2390,N_1841,N_1407);
nand U2391 (N_2391,N_1496,N_1878);
xor U2392 (N_2392,N_1723,N_1193);
or U2393 (N_2393,N_1134,N_1398);
nand U2394 (N_2394,N_1069,N_1445);
nor U2395 (N_2395,N_1661,N_1565);
and U2396 (N_2396,N_1444,N_1271);
nor U2397 (N_2397,N_1554,N_1630);
nand U2398 (N_2398,N_1702,N_1989);
and U2399 (N_2399,N_1500,N_1485);
nand U2400 (N_2400,N_1737,N_1628);
xnor U2401 (N_2401,N_1448,N_1377);
nor U2402 (N_2402,N_1635,N_1126);
and U2403 (N_2403,N_1181,N_1177);
xnor U2404 (N_2404,N_1525,N_1197);
and U2405 (N_2405,N_1558,N_1471);
xnor U2406 (N_2406,N_1640,N_1767);
nor U2407 (N_2407,N_1294,N_1903);
nand U2408 (N_2408,N_1149,N_1983);
nand U2409 (N_2409,N_1566,N_1222);
or U2410 (N_2410,N_1340,N_1215);
and U2411 (N_2411,N_1089,N_1645);
xor U2412 (N_2412,N_1921,N_1901);
nand U2413 (N_2413,N_1890,N_1757);
nor U2414 (N_2414,N_1281,N_1244);
and U2415 (N_2415,N_1986,N_1648);
or U2416 (N_2416,N_1860,N_1490);
and U2417 (N_2417,N_1499,N_1614);
and U2418 (N_2418,N_1316,N_1146);
and U2419 (N_2419,N_1232,N_1803);
and U2420 (N_2420,N_1568,N_1743);
and U2421 (N_2421,N_1947,N_1705);
nand U2422 (N_2422,N_1404,N_1587);
or U2423 (N_2423,N_1813,N_1900);
or U2424 (N_2424,N_1105,N_1239);
and U2425 (N_2425,N_1431,N_1567);
or U2426 (N_2426,N_1704,N_1072);
or U2427 (N_2427,N_1358,N_1680);
or U2428 (N_2428,N_1109,N_1987);
nand U2429 (N_2429,N_1477,N_1676);
and U2430 (N_2430,N_1520,N_1199);
or U2431 (N_2431,N_1882,N_1417);
or U2432 (N_2432,N_1332,N_1698);
or U2433 (N_2433,N_1366,N_1532);
nor U2434 (N_2434,N_1574,N_1887);
and U2435 (N_2435,N_1268,N_1005);
nand U2436 (N_2436,N_1620,N_1696);
and U2437 (N_2437,N_1569,N_1626);
and U2438 (N_2438,N_1933,N_1965);
or U2439 (N_2439,N_1859,N_1220);
nor U2440 (N_2440,N_1021,N_1673);
and U2441 (N_2441,N_1869,N_1580);
or U2442 (N_2442,N_1917,N_1538);
nor U2443 (N_2443,N_1667,N_1411);
xnor U2444 (N_2444,N_1560,N_1658);
nand U2445 (N_2445,N_1277,N_1724);
and U2446 (N_2446,N_1390,N_1771);
or U2447 (N_2447,N_1939,N_1470);
and U2448 (N_2448,N_1043,N_1982);
and U2449 (N_2449,N_1104,N_1636);
xnor U2450 (N_2450,N_1371,N_1075);
nand U2451 (N_2451,N_1434,N_1514);
or U2452 (N_2452,N_1252,N_1295);
nand U2453 (N_2453,N_1441,N_1693);
nor U2454 (N_2454,N_1306,N_1550);
nor U2455 (N_2455,N_1472,N_1446);
nand U2456 (N_2456,N_1709,N_1494);
and U2457 (N_2457,N_1852,N_1160);
nor U2458 (N_2458,N_1074,N_1637);
and U2459 (N_2459,N_1960,N_1928);
nor U2460 (N_2460,N_1264,N_1052);
nor U2461 (N_2461,N_1906,N_1106);
or U2462 (N_2462,N_1816,N_1556);
or U2463 (N_2463,N_1617,N_1302);
or U2464 (N_2464,N_1246,N_1546);
and U2465 (N_2465,N_1923,N_1503);
nor U2466 (N_2466,N_1888,N_1420);
nor U2467 (N_2467,N_1198,N_1424);
or U2468 (N_2468,N_1929,N_1726);
or U2469 (N_2469,N_1187,N_1079);
nand U2470 (N_2470,N_1684,N_1402);
or U2471 (N_2471,N_1325,N_1289);
and U2472 (N_2472,N_1082,N_1953);
nand U2473 (N_2473,N_1266,N_1898);
nand U2474 (N_2474,N_1996,N_1307);
nor U2475 (N_2475,N_1049,N_1389);
and U2476 (N_2476,N_1065,N_1980);
nor U2477 (N_2477,N_1102,N_1862);
nand U2478 (N_2478,N_1657,N_1346);
or U2479 (N_2479,N_1807,N_1827);
and U2480 (N_2480,N_1096,N_1792);
nand U2481 (N_2481,N_1946,N_1165);
or U2482 (N_2482,N_1070,N_1291);
or U2483 (N_2483,N_1780,N_1170);
nor U2484 (N_2484,N_1437,N_1865);
nor U2485 (N_2485,N_1017,N_1711);
nor U2486 (N_2486,N_1736,N_1442);
nand U2487 (N_2487,N_1212,N_1063);
and U2488 (N_2488,N_1046,N_1904);
nor U2489 (N_2489,N_1609,N_1076);
xor U2490 (N_2490,N_1689,N_1952);
or U2491 (N_2491,N_1078,N_1963);
or U2492 (N_2492,N_1806,N_1985);
nand U2493 (N_2493,N_1759,N_1842);
nor U2494 (N_2494,N_1247,N_1116);
nor U2495 (N_2495,N_1144,N_1592);
nand U2496 (N_2496,N_1627,N_1299);
nor U2497 (N_2497,N_1873,N_1148);
xor U2498 (N_2498,N_1872,N_1262);
or U2499 (N_2499,N_1750,N_1200);
nand U2500 (N_2500,N_1547,N_1999);
nor U2501 (N_2501,N_1963,N_1052);
nor U2502 (N_2502,N_1278,N_1753);
and U2503 (N_2503,N_1235,N_1204);
nand U2504 (N_2504,N_1587,N_1528);
xor U2505 (N_2505,N_1611,N_1484);
and U2506 (N_2506,N_1725,N_1474);
or U2507 (N_2507,N_1152,N_1668);
and U2508 (N_2508,N_1308,N_1829);
or U2509 (N_2509,N_1864,N_1332);
and U2510 (N_2510,N_1081,N_1909);
and U2511 (N_2511,N_1041,N_1959);
and U2512 (N_2512,N_1365,N_1763);
nor U2513 (N_2513,N_1682,N_1808);
or U2514 (N_2514,N_1780,N_1696);
nand U2515 (N_2515,N_1779,N_1550);
xnor U2516 (N_2516,N_1047,N_1363);
nor U2517 (N_2517,N_1001,N_1050);
nand U2518 (N_2518,N_1480,N_1047);
nor U2519 (N_2519,N_1621,N_1896);
nor U2520 (N_2520,N_1701,N_1219);
nor U2521 (N_2521,N_1060,N_1700);
and U2522 (N_2522,N_1999,N_1949);
xnor U2523 (N_2523,N_1122,N_1062);
or U2524 (N_2524,N_1694,N_1863);
and U2525 (N_2525,N_1204,N_1255);
and U2526 (N_2526,N_1304,N_1114);
xnor U2527 (N_2527,N_1106,N_1736);
nand U2528 (N_2528,N_1052,N_1406);
and U2529 (N_2529,N_1006,N_1649);
nor U2530 (N_2530,N_1530,N_1591);
or U2531 (N_2531,N_1561,N_1868);
or U2532 (N_2532,N_1385,N_1657);
nand U2533 (N_2533,N_1692,N_1572);
nor U2534 (N_2534,N_1139,N_1269);
and U2535 (N_2535,N_1277,N_1284);
nand U2536 (N_2536,N_1798,N_1113);
and U2537 (N_2537,N_1333,N_1848);
xnor U2538 (N_2538,N_1241,N_1040);
and U2539 (N_2539,N_1049,N_1028);
or U2540 (N_2540,N_1000,N_1227);
or U2541 (N_2541,N_1954,N_1735);
nor U2542 (N_2542,N_1370,N_1709);
nor U2543 (N_2543,N_1504,N_1623);
or U2544 (N_2544,N_1115,N_1434);
or U2545 (N_2545,N_1225,N_1014);
nand U2546 (N_2546,N_1425,N_1354);
nand U2547 (N_2547,N_1261,N_1642);
and U2548 (N_2548,N_1302,N_1391);
xnor U2549 (N_2549,N_1075,N_1725);
or U2550 (N_2550,N_1136,N_1364);
nor U2551 (N_2551,N_1088,N_1789);
and U2552 (N_2552,N_1740,N_1871);
nor U2553 (N_2553,N_1919,N_1817);
or U2554 (N_2554,N_1150,N_1910);
or U2555 (N_2555,N_1209,N_1625);
or U2556 (N_2556,N_1247,N_1400);
and U2557 (N_2557,N_1622,N_1536);
xor U2558 (N_2558,N_1701,N_1045);
and U2559 (N_2559,N_1166,N_1619);
xor U2560 (N_2560,N_1518,N_1485);
or U2561 (N_2561,N_1331,N_1316);
nor U2562 (N_2562,N_1842,N_1112);
nor U2563 (N_2563,N_1068,N_1662);
and U2564 (N_2564,N_1424,N_1518);
and U2565 (N_2565,N_1633,N_1538);
nor U2566 (N_2566,N_1694,N_1157);
xor U2567 (N_2567,N_1980,N_1650);
nand U2568 (N_2568,N_1767,N_1254);
nand U2569 (N_2569,N_1972,N_1631);
or U2570 (N_2570,N_1799,N_1407);
or U2571 (N_2571,N_1519,N_1526);
xor U2572 (N_2572,N_1531,N_1829);
nand U2573 (N_2573,N_1358,N_1836);
and U2574 (N_2574,N_1255,N_1465);
xnor U2575 (N_2575,N_1207,N_1921);
nor U2576 (N_2576,N_1558,N_1993);
nand U2577 (N_2577,N_1516,N_1739);
xnor U2578 (N_2578,N_1580,N_1434);
or U2579 (N_2579,N_1090,N_1115);
nand U2580 (N_2580,N_1552,N_1361);
nand U2581 (N_2581,N_1645,N_1863);
or U2582 (N_2582,N_1091,N_1833);
and U2583 (N_2583,N_1912,N_1602);
nand U2584 (N_2584,N_1656,N_1735);
and U2585 (N_2585,N_1946,N_1832);
nor U2586 (N_2586,N_1443,N_1481);
nor U2587 (N_2587,N_1332,N_1397);
nor U2588 (N_2588,N_1639,N_1531);
nor U2589 (N_2589,N_1310,N_1921);
nor U2590 (N_2590,N_1541,N_1308);
nor U2591 (N_2591,N_1945,N_1778);
nor U2592 (N_2592,N_1084,N_1251);
xnor U2593 (N_2593,N_1931,N_1730);
and U2594 (N_2594,N_1473,N_1760);
nand U2595 (N_2595,N_1253,N_1423);
nand U2596 (N_2596,N_1492,N_1867);
nor U2597 (N_2597,N_1187,N_1570);
and U2598 (N_2598,N_1838,N_1422);
and U2599 (N_2599,N_1673,N_1598);
and U2600 (N_2600,N_1603,N_1396);
xnor U2601 (N_2601,N_1436,N_1509);
or U2602 (N_2602,N_1951,N_1113);
nand U2603 (N_2603,N_1139,N_1875);
nor U2604 (N_2604,N_1690,N_1054);
nor U2605 (N_2605,N_1403,N_1995);
nand U2606 (N_2606,N_1475,N_1745);
xnor U2607 (N_2607,N_1508,N_1522);
nor U2608 (N_2608,N_1118,N_1940);
nor U2609 (N_2609,N_1191,N_1695);
or U2610 (N_2610,N_1342,N_1077);
and U2611 (N_2611,N_1178,N_1149);
or U2612 (N_2612,N_1041,N_1999);
nand U2613 (N_2613,N_1959,N_1902);
nor U2614 (N_2614,N_1289,N_1368);
or U2615 (N_2615,N_1983,N_1905);
or U2616 (N_2616,N_1914,N_1354);
or U2617 (N_2617,N_1328,N_1647);
xor U2618 (N_2618,N_1364,N_1264);
nor U2619 (N_2619,N_1318,N_1623);
and U2620 (N_2620,N_1413,N_1489);
or U2621 (N_2621,N_1952,N_1839);
nor U2622 (N_2622,N_1844,N_1478);
or U2623 (N_2623,N_1609,N_1410);
or U2624 (N_2624,N_1552,N_1313);
and U2625 (N_2625,N_1004,N_1008);
and U2626 (N_2626,N_1464,N_1077);
nor U2627 (N_2627,N_1345,N_1212);
and U2628 (N_2628,N_1007,N_1973);
or U2629 (N_2629,N_1729,N_1842);
and U2630 (N_2630,N_1771,N_1343);
nor U2631 (N_2631,N_1082,N_1779);
and U2632 (N_2632,N_1939,N_1573);
nor U2633 (N_2633,N_1017,N_1557);
nand U2634 (N_2634,N_1144,N_1517);
xor U2635 (N_2635,N_1187,N_1167);
xnor U2636 (N_2636,N_1578,N_1331);
nand U2637 (N_2637,N_1238,N_1641);
xor U2638 (N_2638,N_1797,N_1316);
nor U2639 (N_2639,N_1226,N_1598);
nor U2640 (N_2640,N_1464,N_1327);
nand U2641 (N_2641,N_1245,N_1993);
nor U2642 (N_2642,N_1786,N_1735);
nor U2643 (N_2643,N_1880,N_1403);
nand U2644 (N_2644,N_1844,N_1082);
and U2645 (N_2645,N_1172,N_1207);
nand U2646 (N_2646,N_1903,N_1819);
and U2647 (N_2647,N_1978,N_1150);
and U2648 (N_2648,N_1341,N_1748);
nor U2649 (N_2649,N_1882,N_1791);
or U2650 (N_2650,N_1550,N_1964);
xor U2651 (N_2651,N_1893,N_1753);
or U2652 (N_2652,N_1981,N_1628);
xnor U2653 (N_2653,N_1224,N_1273);
nand U2654 (N_2654,N_1558,N_1303);
and U2655 (N_2655,N_1368,N_1058);
or U2656 (N_2656,N_1943,N_1206);
nor U2657 (N_2657,N_1640,N_1129);
or U2658 (N_2658,N_1024,N_1229);
nor U2659 (N_2659,N_1530,N_1706);
nand U2660 (N_2660,N_1707,N_1267);
or U2661 (N_2661,N_1524,N_1789);
or U2662 (N_2662,N_1300,N_1727);
nand U2663 (N_2663,N_1493,N_1539);
nor U2664 (N_2664,N_1298,N_1843);
xor U2665 (N_2665,N_1406,N_1945);
nand U2666 (N_2666,N_1742,N_1502);
nor U2667 (N_2667,N_1188,N_1549);
and U2668 (N_2668,N_1776,N_1142);
xor U2669 (N_2669,N_1247,N_1258);
xor U2670 (N_2670,N_1041,N_1207);
or U2671 (N_2671,N_1783,N_1250);
nor U2672 (N_2672,N_1489,N_1924);
and U2673 (N_2673,N_1832,N_1972);
or U2674 (N_2674,N_1755,N_1442);
nand U2675 (N_2675,N_1175,N_1304);
and U2676 (N_2676,N_1094,N_1441);
or U2677 (N_2677,N_1066,N_1937);
nor U2678 (N_2678,N_1499,N_1803);
and U2679 (N_2679,N_1280,N_1134);
nand U2680 (N_2680,N_1041,N_1973);
nand U2681 (N_2681,N_1094,N_1522);
nand U2682 (N_2682,N_1668,N_1008);
xnor U2683 (N_2683,N_1265,N_1662);
nor U2684 (N_2684,N_1512,N_1382);
nand U2685 (N_2685,N_1336,N_1911);
nand U2686 (N_2686,N_1703,N_1868);
xnor U2687 (N_2687,N_1846,N_1313);
nand U2688 (N_2688,N_1179,N_1033);
and U2689 (N_2689,N_1353,N_1068);
or U2690 (N_2690,N_1082,N_1509);
nor U2691 (N_2691,N_1140,N_1457);
or U2692 (N_2692,N_1868,N_1438);
or U2693 (N_2693,N_1809,N_1605);
and U2694 (N_2694,N_1651,N_1523);
and U2695 (N_2695,N_1554,N_1034);
nand U2696 (N_2696,N_1355,N_1533);
or U2697 (N_2697,N_1860,N_1045);
nor U2698 (N_2698,N_1275,N_1741);
nor U2699 (N_2699,N_1628,N_1153);
nor U2700 (N_2700,N_1050,N_1394);
and U2701 (N_2701,N_1797,N_1481);
and U2702 (N_2702,N_1620,N_1451);
and U2703 (N_2703,N_1803,N_1278);
nor U2704 (N_2704,N_1152,N_1808);
or U2705 (N_2705,N_1968,N_1321);
or U2706 (N_2706,N_1243,N_1029);
or U2707 (N_2707,N_1110,N_1661);
nor U2708 (N_2708,N_1847,N_1052);
nand U2709 (N_2709,N_1041,N_1644);
or U2710 (N_2710,N_1215,N_1834);
xnor U2711 (N_2711,N_1851,N_1877);
or U2712 (N_2712,N_1858,N_1503);
or U2713 (N_2713,N_1338,N_1469);
or U2714 (N_2714,N_1765,N_1032);
or U2715 (N_2715,N_1034,N_1057);
and U2716 (N_2716,N_1782,N_1427);
or U2717 (N_2717,N_1256,N_1216);
nand U2718 (N_2718,N_1759,N_1369);
or U2719 (N_2719,N_1597,N_1793);
nor U2720 (N_2720,N_1520,N_1556);
nand U2721 (N_2721,N_1654,N_1326);
and U2722 (N_2722,N_1823,N_1646);
or U2723 (N_2723,N_1949,N_1345);
or U2724 (N_2724,N_1597,N_1667);
nor U2725 (N_2725,N_1349,N_1964);
nand U2726 (N_2726,N_1320,N_1992);
nor U2727 (N_2727,N_1968,N_1905);
and U2728 (N_2728,N_1922,N_1630);
nand U2729 (N_2729,N_1205,N_1749);
or U2730 (N_2730,N_1582,N_1387);
xnor U2731 (N_2731,N_1352,N_1766);
nor U2732 (N_2732,N_1139,N_1594);
nor U2733 (N_2733,N_1495,N_1103);
xor U2734 (N_2734,N_1033,N_1552);
nor U2735 (N_2735,N_1749,N_1553);
and U2736 (N_2736,N_1577,N_1646);
and U2737 (N_2737,N_1068,N_1650);
and U2738 (N_2738,N_1242,N_1806);
nand U2739 (N_2739,N_1887,N_1236);
and U2740 (N_2740,N_1840,N_1344);
nor U2741 (N_2741,N_1137,N_1083);
nor U2742 (N_2742,N_1434,N_1645);
nor U2743 (N_2743,N_1225,N_1999);
nand U2744 (N_2744,N_1288,N_1567);
nand U2745 (N_2745,N_1514,N_1734);
nor U2746 (N_2746,N_1185,N_1765);
and U2747 (N_2747,N_1318,N_1554);
xnor U2748 (N_2748,N_1499,N_1063);
xor U2749 (N_2749,N_1008,N_1788);
nand U2750 (N_2750,N_1428,N_1171);
nor U2751 (N_2751,N_1804,N_1670);
and U2752 (N_2752,N_1199,N_1976);
nand U2753 (N_2753,N_1158,N_1327);
and U2754 (N_2754,N_1528,N_1918);
nand U2755 (N_2755,N_1972,N_1375);
nand U2756 (N_2756,N_1294,N_1803);
or U2757 (N_2757,N_1429,N_1661);
or U2758 (N_2758,N_1474,N_1604);
or U2759 (N_2759,N_1118,N_1883);
or U2760 (N_2760,N_1423,N_1745);
nand U2761 (N_2761,N_1494,N_1037);
nor U2762 (N_2762,N_1600,N_1657);
or U2763 (N_2763,N_1932,N_1994);
and U2764 (N_2764,N_1365,N_1157);
and U2765 (N_2765,N_1999,N_1257);
xnor U2766 (N_2766,N_1684,N_1126);
nand U2767 (N_2767,N_1080,N_1464);
and U2768 (N_2768,N_1689,N_1337);
nor U2769 (N_2769,N_1969,N_1851);
or U2770 (N_2770,N_1859,N_1262);
or U2771 (N_2771,N_1624,N_1729);
nand U2772 (N_2772,N_1499,N_1494);
nand U2773 (N_2773,N_1385,N_1529);
and U2774 (N_2774,N_1166,N_1724);
and U2775 (N_2775,N_1041,N_1324);
xnor U2776 (N_2776,N_1148,N_1264);
xnor U2777 (N_2777,N_1871,N_1128);
or U2778 (N_2778,N_1939,N_1338);
or U2779 (N_2779,N_1366,N_1027);
nand U2780 (N_2780,N_1784,N_1513);
or U2781 (N_2781,N_1430,N_1843);
xnor U2782 (N_2782,N_1889,N_1769);
or U2783 (N_2783,N_1720,N_1481);
nor U2784 (N_2784,N_1906,N_1732);
and U2785 (N_2785,N_1542,N_1116);
nor U2786 (N_2786,N_1279,N_1774);
nor U2787 (N_2787,N_1840,N_1515);
nand U2788 (N_2788,N_1687,N_1249);
xor U2789 (N_2789,N_1549,N_1399);
nand U2790 (N_2790,N_1968,N_1315);
or U2791 (N_2791,N_1207,N_1686);
or U2792 (N_2792,N_1311,N_1613);
xor U2793 (N_2793,N_1191,N_1107);
nor U2794 (N_2794,N_1658,N_1885);
nand U2795 (N_2795,N_1363,N_1659);
xnor U2796 (N_2796,N_1126,N_1245);
xor U2797 (N_2797,N_1739,N_1579);
or U2798 (N_2798,N_1225,N_1872);
and U2799 (N_2799,N_1613,N_1060);
nand U2800 (N_2800,N_1357,N_1412);
and U2801 (N_2801,N_1063,N_1637);
or U2802 (N_2802,N_1877,N_1379);
nand U2803 (N_2803,N_1934,N_1725);
or U2804 (N_2804,N_1339,N_1923);
and U2805 (N_2805,N_1806,N_1758);
or U2806 (N_2806,N_1520,N_1300);
or U2807 (N_2807,N_1865,N_1004);
nor U2808 (N_2808,N_1615,N_1355);
nand U2809 (N_2809,N_1931,N_1821);
or U2810 (N_2810,N_1014,N_1988);
and U2811 (N_2811,N_1652,N_1311);
or U2812 (N_2812,N_1075,N_1442);
or U2813 (N_2813,N_1939,N_1315);
or U2814 (N_2814,N_1265,N_1737);
nor U2815 (N_2815,N_1657,N_1539);
and U2816 (N_2816,N_1708,N_1477);
or U2817 (N_2817,N_1298,N_1942);
and U2818 (N_2818,N_1409,N_1827);
nand U2819 (N_2819,N_1137,N_1127);
or U2820 (N_2820,N_1318,N_1638);
nand U2821 (N_2821,N_1556,N_1974);
and U2822 (N_2822,N_1984,N_1597);
nand U2823 (N_2823,N_1908,N_1423);
nand U2824 (N_2824,N_1753,N_1315);
or U2825 (N_2825,N_1445,N_1041);
nor U2826 (N_2826,N_1864,N_1494);
nand U2827 (N_2827,N_1937,N_1634);
nor U2828 (N_2828,N_1943,N_1074);
or U2829 (N_2829,N_1109,N_1874);
nor U2830 (N_2830,N_1636,N_1281);
or U2831 (N_2831,N_1903,N_1849);
and U2832 (N_2832,N_1921,N_1012);
nor U2833 (N_2833,N_1815,N_1027);
nor U2834 (N_2834,N_1103,N_1606);
or U2835 (N_2835,N_1276,N_1392);
or U2836 (N_2836,N_1246,N_1472);
nor U2837 (N_2837,N_1124,N_1289);
nor U2838 (N_2838,N_1638,N_1030);
and U2839 (N_2839,N_1118,N_1853);
and U2840 (N_2840,N_1158,N_1789);
xnor U2841 (N_2841,N_1158,N_1783);
and U2842 (N_2842,N_1338,N_1370);
nand U2843 (N_2843,N_1863,N_1767);
nand U2844 (N_2844,N_1362,N_1713);
and U2845 (N_2845,N_1813,N_1234);
nor U2846 (N_2846,N_1208,N_1181);
or U2847 (N_2847,N_1497,N_1478);
nor U2848 (N_2848,N_1330,N_1242);
nor U2849 (N_2849,N_1101,N_1239);
nand U2850 (N_2850,N_1780,N_1820);
nor U2851 (N_2851,N_1308,N_1368);
or U2852 (N_2852,N_1396,N_1617);
nand U2853 (N_2853,N_1033,N_1275);
or U2854 (N_2854,N_1828,N_1706);
or U2855 (N_2855,N_1395,N_1232);
xnor U2856 (N_2856,N_1466,N_1521);
xor U2857 (N_2857,N_1326,N_1225);
nor U2858 (N_2858,N_1207,N_1581);
xor U2859 (N_2859,N_1180,N_1417);
or U2860 (N_2860,N_1577,N_1243);
xnor U2861 (N_2861,N_1185,N_1107);
nor U2862 (N_2862,N_1568,N_1155);
nand U2863 (N_2863,N_1374,N_1668);
nand U2864 (N_2864,N_1211,N_1085);
or U2865 (N_2865,N_1810,N_1692);
xor U2866 (N_2866,N_1167,N_1880);
or U2867 (N_2867,N_1159,N_1194);
nand U2868 (N_2868,N_1333,N_1409);
or U2869 (N_2869,N_1821,N_1295);
or U2870 (N_2870,N_1837,N_1838);
or U2871 (N_2871,N_1593,N_1371);
or U2872 (N_2872,N_1498,N_1544);
and U2873 (N_2873,N_1674,N_1208);
nor U2874 (N_2874,N_1987,N_1733);
nor U2875 (N_2875,N_1295,N_1782);
nand U2876 (N_2876,N_1679,N_1170);
or U2877 (N_2877,N_1015,N_1546);
and U2878 (N_2878,N_1483,N_1378);
or U2879 (N_2879,N_1208,N_1442);
nor U2880 (N_2880,N_1686,N_1900);
and U2881 (N_2881,N_1623,N_1825);
nand U2882 (N_2882,N_1519,N_1265);
nor U2883 (N_2883,N_1336,N_1381);
xor U2884 (N_2884,N_1849,N_1696);
nor U2885 (N_2885,N_1430,N_1013);
and U2886 (N_2886,N_1156,N_1683);
nand U2887 (N_2887,N_1065,N_1949);
xnor U2888 (N_2888,N_1485,N_1211);
or U2889 (N_2889,N_1000,N_1918);
and U2890 (N_2890,N_1074,N_1379);
and U2891 (N_2891,N_1908,N_1984);
and U2892 (N_2892,N_1205,N_1747);
or U2893 (N_2893,N_1949,N_1813);
nor U2894 (N_2894,N_1516,N_1533);
nor U2895 (N_2895,N_1831,N_1401);
and U2896 (N_2896,N_1346,N_1985);
xnor U2897 (N_2897,N_1489,N_1775);
or U2898 (N_2898,N_1050,N_1042);
nand U2899 (N_2899,N_1839,N_1892);
and U2900 (N_2900,N_1461,N_1027);
and U2901 (N_2901,N_1782,N_1000);
nand U2902 (N_2902,N_1074,N_1155);
xnor U2903 (N_2903,N_1807,N_1509);
xnor U2904 (N_2904,N_1588,N_1753);
nand U2905 (N_2905,N_1352,N_1914);
xor U2906 (N_2906,N_1554,N_1224);
or U2907 (N_2907,N_1292,N_1291);
xnor U2908 (N_2908,N_1646,N_1091);
nand U2909 (N_2909,N_1958,N_1424);
nor U2910 (N_2910,N_1724,N_1843);
nand U2911 (N_2911,N_1032,N_1370);
xor U2912 (N_2912,N_1240,N_1363);
or U2913 (N_2913,N_1650,N_1325);
nor U2914 (N_2914,N_1451,N_1691);
nor U2915 (N_2915,N_1597,N_1290);
and U2916 (N_2916,N_1658,N_1059);
or U2917 (N_2917,N_1226,N_1606);
nand U2918 (N_2918,N_1002,N_1232);
nand U2919 (N_2919,N_1020,N_1361);
and U2920 (N_2920,N_1203,N_1464);
and U2921 (N_2921,N_1422,N_1578);
and U2922 (N_2922,N_1309,N_1608);
and U2923 (N_2923,N_1108,N_1227);
and U2924 (N_2924,N_1320,N_1155);
and U2925 (N_2925,N_1758,N_1817);
nand U2926 (N_2926,N_1359,N_1545);
or U2927 (N_2927,N_1507,N_1269);
xor U2928 (N_2928,N_1239,N_1854);
or U2929 (N_2929,N_1167,N_1430);
nor U2930 (N_2930,N_1737,N_1882);
nor U2931 (N_2931,N_1417,N_1748);
nor U2932 (N_2932,N_1480,N_1906);
nor U2933 (N_2933,N_1823,N_1987);
nand U2934 (N_2934,N_1392,N_1063);
nor U2935 (N_2935,N_1333,N_1161);
or U2936 (N_2936,N_1544,N_1720);
nand U2937 (N_2937,N_1290,N_1273);
and U2938 (N_2938,N_1327,N_1162);
nand U2939 (N_2939,N_1392,N_1381);
and U2940 (N_2940,N_1840,N_1819);
and U2941 (N_2941,N_1356,N_1120);
or U2942 (N_2942,N_1130,N_1609);
nand U2943 (N_2943,N_1622,N_1750);
and U2944 (N_2944,N_1858,N_1417);
or U2945 (N_2945,N_1726,N_1947);
xor U2946 (N_2946,N_1669,N_1396);
and U2947 (N_2947,N_1346,N_1673);
nor U2948 (N_2948,N_1468,N_1879);
xnor U2949 (N_2949,N_1863,N_1510);
nand U2950 (N_2950,N_1950,N_1307);
xnor U2951 (N_2951,N_1717,N_1389);
and U2952 (N_2952,N_1846,N_1378);
xor U2953 (N_2953,N_1304,N_1186);
nand U2954 (N_2954,N_1928,N_1498);
or U2955 (N_2955,N_1828,N_1133);
nor U2956 (N_2956,N_1602,N_1243);
or U2957 (N_2957,N_1522,N_1061);
and U2958 (N_2958,N_1554,N_1872);
and U2959 (N_2959,N_1003,N_1126);
nor U2960 (N_2960,N_1989,N_1021);
and U2961 (N_2961,N_1895,N_1642);
or U2962 (N_2962,N_1258,N_1789);
nand U2963 (N_2963,N_1467,N_1649);
nand U2964 (N_2964,N_1150,N_1678);
nor U2965 (N_2965,N_1551,N_1386);
or U2966 (N_2966,N_1333,N_1894);
nand U2967 (N_2967,N_1763,N_1914);
xor U2968 (N_2968,N_1323,N_1511);
or U2969 (N_2969,N_1033,N_1594);
nor U2970 (N_2970,N_1976,N_1759);
nor U2971 (N_2971,N_1212,N_1203);
and U2972 (N_2972,N_1728,N_1769);
or U2973 (N_2973,N_1468,N_1280);
xnor U2974 (N_2974,N_1517,N_1539);
nor U2975 (N_2975,N_1795,N_1352);
nor U2976 (N_2976,N_1565,N_1829);
or U2977 (N_2977,N_1471,N_1474);
or U2978 (N_2978,N_1342,N_1412);
or U2979 (N_2979,N_1281,N_1228);
or U2980 (N_2980,N_1216,N_1827);
nand U2981 (N_2981,N_1279,N_1786);
xor U2982 (N_2982,N_1096,N_1088);
or U2983 (N_2983,N_1053,N_1540);
and U2984 (N_2984,N_1553,N_1110);
nand U2985 (N_2985,N_1727,N_1111);
xnor U2986 (N_2986,N_1473,N_1253);
or U2987 (N_2987,N_1491,N_1410);
and U2988 (N_2988,N_1276,N_1767);
nand U2989 (N_2989,N_1437,N_1591);
nor U2990 (N_2990,N_1592,N_1377);
xnor U2991 (N_2991,N_1877,N_1170);
nor U2992 (N_2992,N_1291,N_1096);
or U2993 (N_2993,N_1790,N_1373);
xnor U2994 (N_2994,N_1902,N_1555);
or U2995 (N_2995,N_1253,N_1975);
nor U2996 (N_2996,N_1113,N_1174);
nand U2997 (N_2997,N_1408,N_1516);
xnor U2998 (N_2998,N_1300,N_1210);
and U2999 (N_2999,N_1066,N_1339);
nor U3000 (N_3000,N_2307,N_2985);
xnor U3001 (N_3001,N_2828,N_2272);
nor U3002 (N_3002,N_2552,N_2295);
or U3003 (N_3003,N_2490,N_2656);
nor U3004 (N_3004,N_2485,N_2319);
or U3005 (N_3005,N_2332,N_2971);
nand U3006 (N_3006,N_2080,N_2758);
nand U3007 (N_3007,N_2394,N_2683);
and U3008 (N_3008,N_2854,N_2056);
nor U3009 (N_3009,N_2499,N_2810);
nor U3010 (N_3010,N_2927,N_2739);
or U3011 (N_3011,N_2035,N_2231);
and U3012 (N_3012,N_2510,N_2716);
nor U3013 (N_3013,N_2778,N_2199);
or U3014 (N_3014,N_2823,N_2809);
or U3015 (N_3015,N_2302,N_2724);
or U3016 (N_3016,N_2795,N_2062);
and U3017 (N_3017,N_2557,N_2110);
and U3018 (N_3018,N_2010,N_2844);
xor U3019 (N_3019,N_2775,N_2234);
nand U3020 (N_3020,N_2802,N_2240);
nand U3021 (N_3021,N_2569,N_2322);
and U3022 (N_3022,N_2507,N_2696);
xnor U3023 (N_3023,N_2467,N_2296);
xnor U3024 (N_3024,N_2556,N_2201);
and U3025 (N_3025,N_2738,N_2550);
nand U3026 (N_3026,N_2612,N_2965);
nand U3027 (N_3027,N_2089,N_2131);
xnor U3028 (N_3028,N_2482,N_2388);
or U3029 (N_3029,N_2674,N_2229);
xor U3030 (N_3030,N_2937,N_2679);
nand U3031 (N_3031,N_2226,N_2179);
nand U3032 (N_3032,N_2324,N_2602);
nand U3033 (N_3033,N_2061,N_2200);
or U3034 (N_3034,N_2432,N_2911);
nor U3035 (N_3035,N_2017,N_2230);
nand U3036 (N_3036,N_2641,N_2814);
and U3037 (N_3037,N_2681,N_2456);
or U3038 (N_3038,N_2190,N_2816);
or U3039 (N_3039,N_2955,N_2022);
nand U3040 (N_3040,N_2609,N_2578);
nor U3041 (N_3041,N_2437,N_2594);
nor U3042 (N_3042,N_2559,N_2400);
or U3043 (N_3043,N_2922,N_2285);
and U3044 (N_3044,N_2355,N_2849);
and U3045 (N_3045,N_2077,N_2317);
or U3046 (N_3046,N_2289,N_2518);
xor U3047 (N_3047,N_2514,N_2275);
or U3048 (N_3048,N_2459,N_2779);
and U3049 (N_3049,N_2380,N_2172);
nor U3050 (N_3050,N_2105,N_2078);
or U3051 (N_3051,N_2255,N_2541);
nand U3052 (N_3052,N_2263,N_2382);
and U3053 (N_3053,N_2721,N_2577);
or U3054 (N_3054,N_2053,N_2977);
nand U3055 (N_3055,N_2712,N_2100);
xor U3056 (N_3056,N_2214,N_2174);
and U3057 (N_3057,N_2206,N_2236);
nor U3058 (N_3058,N_2149,N_2970);
nor U3059 (N_3059,N_2335,N_2422);
nand U3060 (N_3060,N_2649,N_2143);
or U3061 (N_3061,N_2710,N_2827);
xnor U3062 (N_3062,N_2479,N_2204);
and U3063 (N_3063,N_2919,N_2283);
nand U3064 (N_3064,N_2789,N_2469);
nor U3065 (N_3065,N_2227,N_2237);
or U3066 (N_3066,N_2278,N_2112);
nand U3067 (N_3067,N_2326,N_2808);
nand U3068 (N_3068,N_2320,N_2655);
nor U3069 (N_3069,N_2043,N_2342);
nand U3070 (N_3070,N_2014,N_2057);
xnor U3071 (N_3071,N_2622,N_2385);
nor U3072 (N_3072,N_2763,N_2718);
or U3073 (N_3073,N_2114,N_2512);
xnor U3074 (N_3074,N_2680,N_2973);
nand U3075 (N_3075,N_2566,N_2892);
and U3076 (N_3076,N_2187,N_2393);
or U3077 (N_3077,N_2901,N_2635);
nand U3078 (N_3078,N_2733,N_2740);
nor U3079 (N_3079,N_2625,N_2856);
nand U3080 (N_3080,N_2580,N_2815);
nor U3081 (N_3081,N_2637,N_2817);
and U3082 (N_3082,N_2346,N_2480);
nor U3083 (N_3083,N_2157,N_2395);
or U3084 (N_3084,N_2158,N_2208);
nand U3085 (N_3085,N_2491,N_2451);
and U3086 (N_3086,N_2787,N_2313);
or U3087 (N_3087,N_2867,N_2636);
or U3088 (N_3088,N_2345,N_2835);
or U3089 (N_3089,N_2101,N_2581);
and U3090 (N_3090,N_2306,N_2952);
and U3091 (N_3091,N_2308,N_2162);
nor U3092 (N_3092,N_2755,N_2483);
nand U3093 (N_3093,N_2545,N_2800);
nor U3094 (N_3094,N_2026,N_2711);
nor U3095 (N_3095,N_2608,N_2847);
nand U3096 (N_3096,N_2966,N_2735);
and U3097 (N_3097,N_2309,N_2979);
or U3098 (N_3098,N_2438,N_2826);
xnor U3099 (N_3099,N_2825,N_2205);
or U3100 (N_3100,N_2877,N_2381);
nand U3101 (N_3101,N_2799,N_2920);
or U3102 (N_3102,N_2671,N_2249);
nand U3103 (N_3103,N_2722,N_2829);
or U3104 (N_3104,N_2846,N_2848);
xnor U3105 (N_3105,N_2325,N_2423);
nand U3106 (N_3106,N_2543,N_2900);
nor U3107 (N_3107,N_2344,N_2639);
or U3108 (N_3108,N_2812,N_2503);
xor U3109 (N_3109,N_2832,N_2097);
nor U3110 (N_3110,N_2003,N_2780);
nand U3111 (N_3111,N_2551,N_2059);
nor U3112 (N_3112,N_2277,N_2408);
nand U3113 (N_3113,N_2173,N_2606);
xnor U3114 (N_3114,N_2638,N_2153);
or U3115 (N_3115,N_2669,N_2314);
nor U3116 (N_3116,N_2235,N_2884);
nand U3117 (N_3117,N_2837,N_2659);
nand U3118 (N_3118,N_2215,N_2796);
nand U3119 (N_3119,N_2387,N_2851);
nor U3120 (N_3120,N_2122,N_2331);
nand U3121 (N_3121,N_2372,N_2833);
and U3122 (N_3122,N_2488,N_2221);
nand U3123 (N_3123,N_2968,N_2634);
and U3124 (N_3124,N_2442,N_2535);
nor U3125 (N_3125,N_2055,N_2133);
or U3126 (N_3126,N_2468,N_2899);
and U3127 (N_3127,N_2769,N_2751);
or U3128 (N_3128,N_2560,N_2219);
and U3129 (N_3129,N_2086,N_2245);
nor U3130 (N_3130,N_2781,N_2111);
nand U3131 (N_3131,N_2487,N_2529);
nor U3132 (N_3132,N_2357,N_2925);
nand U3133 (N_3133,N_2371,N_2969);
nor U3134 (N_3134,N_2623,N_2861);
and U3135 (N_3135,N_2806,N_2183);
nand U3136 (N_3136,N_2521,N_2081);
or U3137 (N_3137,N_2840,N_2553);
or U3138 (N_3138,N_2707,N_2239);
and U3139 (N_3139,N_2185,N_2992);
and U3140 (N_3140,N_2786,N_2443);
nor U3141 (N_3141,N_2348,N_2269);
xnor U3142 (N_3142,N_2494,N_2378);
xor U3143 (N_3143,N_2138,N_2182);
nand U3144 (N_3144,N_2211,N_2058);
and U3145 (N_3145,N_2570,N_2708);
nor U3146 (N_3146,N_2504,N_2736);
nand U3147 (N_3147,N_2938,N_2359);
or U3148 (N_3148,N_2500,N_2567);
and U3149 (N_3149,N_2008,N_2429);
nand U3150 (N_3150,N_2954,N_2714);
and U3151 (N_3151,N_2343,N_2098);
nor U3152 (N_3152,N_2960,N_2990);
or U3153 (N_3153,N_2210,N_2607);
or U3154 (N_3154,N_2465,N_2785);
nand U3155 (N_3155,N_2374,N_2694);
and U3156 (N_3156,N_2804,N_2794);
and U3157 (N_3157,N_2753,N_2449);
nand U3158 (N_3158,N_2752,N_2166);
nor U3159 (N_3159,N_2905,N_2540);
and U3160 (N_3160,N_2011,N_2599);
or U3161 (N_3161,N_2771,N_2116);
and U3162 (N_3162,N_2093,N_2007);
or U3163 (N_3163,N_2522,N_2168);
nor U3164 (N_3164,N_2018,N_2742);
and U3165 (N_3165,N_2349,N_2247);
and U3166 (N_3166,N_2460,N_2617);
nor U3167 (N_3167,N_2863,N_2384);
or U3168 (N_3168,N_2147,N_2558);
xnor U3169 (N_3169,N_2536,N_2923);
or U3170 (N_3170,N_2417,N_2360);
nand U3171 (N_3171,N_2843,N_2462);
xor U3172 (N_3172,N_2083,N_2874);
or U3173 (N_3173,N_2358,N_2627);
and U3174 (N_3174,N_2931,N_2252);
nor U3175 (N_3175,N_2261,N_2537);
or U3176 (N_3176,N_2509,N_2389);
nor U3177 (N_3177,N_2879,N_2321);
nor U3178 (N_3178,N_2069,N_2644);
nand U3179 (N_3179,N_2405,N_2663);
or U3180 (N_3180,N_2130,N_2244);
or U3181 (N_3181,N_2421,N_2126);
xor U3182 (N_3182,N_2783,N_2547);
xor U3183 (N_3183,N_2333,N_2697);
and U3184 (N_3184,N_2180,N_2464);
nand U3185 (N_3185,N_2142,N_2109);
and U3186 (N_3186,N_2782,N_2565);
nor U3187 (N_3187,N_2652,N_2818);
and U3188 (N_3188,N_2555,N_2542);
nor U3189 (N_3189,N_2095,N_2998);
nor U3190 (N_3190,N_2232,N_2618);
and U3191 (N_3191,N_2759,N_2616);
or U3192 (N_3192,N_2648,N_2868);
nor U3193 (N_3193,N_2734,N_2534);
xnor U3194 (N_3194,N_2890,N_2129);
xnor U3195 (N_3195,N_2945,N_2439);
nand U3196 (N_3196,N_2259,N_2489);
or U3197 (N_3197,N_2222,N_2628);
or U3198 (N_3198,N_2171,N_2450);
xor U3199 (N_3199,N_2192,N_2476);
xor U3200 (N_3200,N_2574,N_2719);
xor U3201 (N_3201,N_2746,N_2016);
and U3202 (N_3202,N_2598,N_2473);
nor U3203 (N_3203,N_2506,N_2788);
and U3204 (N_3204,N_2398,N_2297);
or U3205 (N_3205,N_2959,N_2702);
nor U3206 (N_3206,N_2591,N_2562);
nor U3207 (N_3207,N_2997,N_2132);
nor U3208 (N_3208,N_2015,N_2871);
or U3209 (N_3209,N_2903,N_2466);
nand U3210 (N_3210,N_2023,N_2411);
nor U3211 (N_3211,N_2647,N_2596);
nor U3212 (N_3212,N_2528,N_2425);
nand U3213 (N_3213,N_2072,N_2403);
and U3214 (N_3214,N_2957,N_2691);
nand U3215 (N_3215,N_2312,N_2709);
nor U3216 (N_3216,N_2517,N_2548);
nor U3217 (N_3217,N_2113,N_2327);
nand U3218 (N_3218,N_2820,N_2094);
and U3219 (N_3219,N_2493,N_2878);
or U3220 (N_3220,N_2502,N_2791);
nand U3221 (N_3221,N_2049,N_2564);
xnor U3222 (N_3222,N_2981,N_2305);
nand U3223 (N_3223,N_2298,N_2141);
and U3224 (N_3224,N_2063,N_2207);
nand U3225 (N_3225,N_2995,N_2224);
xor U3226 (N_3226,N_2315,N_2178);
nor U3227 (N_3227,N_2964,N_2978);
or U3228 (N_3228,N_2603,N_2184);
nor U3229 (N_3229,N_2044,N_2583);
nand U3230 (N_3230,N_2601,N_2862);
nand U3231 (N_3231,N_2513,N_2128);
nand U3232 (N_3232,N_2203,N_2433);
or U3233 (N_3233,N_2629,N_2568);
nor U3234 (N_3234,N_2853,N_2765);
nand U3235 (N_3235,N_2376,N_2961);
and U3236 (N_3236,N_2164,N_2684);
nand U3237 (N_3237,N_2276,N_2197);
and U3238 (N_3238,N_2370,N_2073);
and U3239 (N_3239,N_2136,N_2692);
nand U3240 (N_3240,N_2757,N_2090);
and U3241 (N_3241,N_2323,N_2698);
or U3242 (N_3242,N_2084,N_2895);
nor U3243 (N_3243,N_2118,N_2060);
nand U3244 (N_3244,N_2962,N_2163);
nand U3245 (N_3245,N_2646,N_2658);
nand U3246 (N_3246,N_2108,N_2350);
and U3247 (N_3247,N_2621,N_2916);
and U3248 (N_3248,N_2434,N_2589);
nand U3249 (N_3249,N_2025,N_2071);
or U3250 (N_3250,N_2793,N_2196);
nand U3251 (N_3251,N_2531,N_2446);
nand U3252 (N_3252,N_2918,N_2909);
xor U3253 (N_3253,N_2883,N_2511);
and U3254 (N_3254,N_2988,N_2497);
nand U3255 (N_3255,N_2299,N_2989);
or U3256 (N_3256,N_2904,N_2134);
nor U3257 (N_3257,N_2140,N_2642);
nor U3258 (N_3258,N_2032,N_2139);
or U3259 (N_3259,N_2650,N_2125);
and U3260 (N_3260,N_2665,N_2361);
nor U3261 (N_3261,N_2260,N_2445);
and U3262 (N_3262,N_2731,N_2310);
nor U3263 (N_3263,N_2910,N_2986);
nor U3264 (N_3264,N_2248,N_2492);
or U3265 (N_3265,N_2756,N_2075);
xor U3266 (N_3266,N_2087,N_2413);
nor U3267 (N_3267,N_2773,N_2369);
and U3268 (N_3268,N_2582,N_2631);
and U3269 (N_3269,N_2519,N_2364);
nand U3270 (N_3270,N_2882,N_2889);
or U3271 (N_3271,N_2914,N_2803);
xnor U3272 (N_3272,N_2447,N_2524);
or U3273 (N_3273,N_2501,N_2191);
nand U3274 (N_3274,N_2311,N_2082);
xor U3275 (N_3275,N_2830,N_2407);
nor U3276 (N_3276,N_2597,N_2967);
nor U3277 (N_3277,N_2726,N_2304);
or U3278 (N_3278,N_2934,N_2186);
nor U3279 (N_3279,N_2744,N_2024);
and U3280 (N_3280,N_2091,N_2974);
nand U3281 (N_3281,N_2643,N_2028);
nor U3282 (N_3282,N_2424,N_2188);
xor U3283 (N_3283,N_2160,N_2949);
xnor U3284 (N_3284,N_2761,N_2031);
or U3285 (N_3285,N_2996,N_2675);
nor U3286 (N_3286,N_2404,N_2328);
or U3287 (N_3287,N_2748,N_2441);
xnor U3288 (N_3288,N_2613,N_2444);
or U3289 (N_3289,N_2645,N_2620);
and U3290 (N_3290,N_2956,N_2561);
xnor U3291 (N_3291,N_2271,N_2842);
nand U3292 (N_3292,N_2605,N_2181);
or U3293 (N_3293,N_2347,N_2019);
or U3294 (N_3294,N_2657,N_2088);
or U3295 (N_3295,N_2984,N_2339);
nand U3296 (N_3296,N_2584,N_2839);
and U3297 (N_3297,N_2390,N_2508);
and U3298 (N_3298,N_2653,N_2928);
xnor U3299 (N_3299,N_2399,N_2885);
and U3300 (N_3300,N_2866,N_2764);
nor U3301 (N_3301,N_2664,N_2801);
nand U3302 (N_3302,N_2983,N_2316);
nand U3303 (N_3303,N_2588,N_2530);
and U3304 (N_3304,N_2571,N_2693);
xnor U3305 (N_3305,N_2033,N_2994);
or U3306 (N_3306,N_2048,N_2189);
nand U3307 (N_3307,N_2170,N_2265);
or U3308 (N_3308,N_2064,N_2209);
nand U3309 (N_3309,N_2030,N_2458);
nand U3310 (N_3310,N_2610,N_2366);
nor U3311 (N_3311,N_2167,N_2704);
and U3312 (N_3312,N_2807,N_2337);
nand U3313 (N_3313,N_2103,N_2662);
nor U3314 (N_3314,N_2148,N_2120);
nor U3315 (N_3315,N_2478,N_2563);
and U3316 (N_3316,N_2668,N_2932);
nor U3317 (N_3317,N_2750,N_2611);
nand U3318 (N_3318,N_2216,N_2586);
or U3319 (N_3319,N_2150,N_2870);
nand U3320 (N_3320,N_2824,N_2225);
nor U3321 (N_3321,N_2749,N_2852);
nor U3322 (N_3322,N_2195,N_2772);
or U3323 (N_3323,N_2373,N_2029);
or U3324 (N_3324,N_2041,N_2367);
or U3325 (N_3325,N_2270,N_2452);
nor U3326 (N_3326,N_2595,N_2435);
nand U3327 (N_3327,N_2544,N_2415);
nor U3328 (N_3328,N_2947,N_2362);
or U3329 (N_3329,N_2732,N_2006);
or U3330 (N_3330,N_2165,N_2689);
nor U3331 (N_3331,N_2288,N_2220);
and U3332 (N_3332,N_2907,N_2291);
nor U3333 (N_3333,N_2104,N_2391);
nor U3334 (N_3334,N_2194,N_2695);
or U3335 (N_3335,N_2127,N_2729);
nor U3336 (N_3336,N_2869,N_2338);
nor U3337 (N_3337,N_2754,N_2677);
nor U3338 (N_3338,N_2632,N_2004);
or U3339 (N_3339,N_2070,N_2515);
or U3340 (N_3340,N_2119,N_2768);
or U3341 (N_3341,N_2250,N_2054);
nor U3342 (N_3342,N_2202,N_2575);
nand U3343 (N_3343,N_2144,N_2484);
xnor U3344 (N_3344,N_2893,N_2121);
or U3345 (N_3345,N_2290,N_2600);
nor U3346 (N_3346,N_2274,N_2766);
and U3347 (N_3347,N_2857,N_2212);
nand U3348 (N_3348,N_2046,N_2264);
nor U3349 (N_3349,N_2036,N_2177);
xnor U3350 (N_3350,N_2115,N_2409);
and U3351 (N_3351,N_2790,N_2747);
or U3352 (N_3352,N_2213,N_2615);
and U3353 (N_3353,N_2811,N_2300);
nor U3354 (N_3354,N_2065,N_2682);
nor U3355 (N_3355,N_2774,N_2092);
nand U3356 (N_3356,N_2539,N_2525);
and U3357 (N_3357,N_2477,N_2619);
nor U3358 (N_3358,N_2526,N_2397);
nand U3359 (N_3359,N_2864,N_2865);
nor U3360 (N_3360,N_2135,N_2876);
nand U3361 (N_3361,N_2418,N_2258);
or U3362 (N_3362,N_2000,N_2038);
nor U3363 (N_3363,N_2392,N_2218);
nand U3364 (N_3364,N_2944,N_2303);
nor U3365 (N_3365,N_2020,N_2156);
and U3366 (N_3366,N_2730,N_2262);
nor U3367 (N_3367,N_2760,N_2329);
nand U3368 (N_3368,N_2436,N_2334);
xor U3369 (N_3369,N_2942,N_2427);
or U3370 (N_3370,N_2688,N_2352);
and U3371 (N_3371,N_2654,N_2743);
nand U3372 (N_3372,N_2268,N_2318);
nand U3373 (N_3373,N_2386,N_2770);
nor U3374 (N_3374,N_2117,N_2254);
nor U3375 (N_3375,N_2193,N_2715);
or U3376 (N_3376,N_2472,N_2107);
and U3377 (N_3377,N_2838,N_2353);
or U3378 (N_3378,N_2440,N_2685);
nand U3379 (N_3379,N_2430,N_2396);
nor U3380 (N_3380,N_2898,N_2950);
and U3381 (N_3381,N_2894,N_2717);
and U3382 (N_3382,N_2940,N_2673);
or U3383 (N_3383,N_2845,N_2836);
nor U3384 (N_3384,N_2354,N_2912);
and U3385 (N_3385,N_2587,N_2953);
or U3386 (N_3386,N_2039,N_2917);
nor U3387 (N_3387,N_2414,N_2527);
or U3388 (N_3388,N_2076,N_2453);
nand U3389 (N_3389,N_2256,N_2474);
nand U3390 (N_3390,N_2151,N_2406);
nand U3391 (N_3391,N_2936,N_2496);
nand U3392 (N_3392,N_2850,N_2410);
and U3393 (N_3393,N_2266,N_2972);
nand U3394 (N_3394,N_2175,N_2047);
or U3395 (N_3395,N_2027,N_2891);
nand U3396 (N_3396,N_2713,N_2287);
or U3397 (N_3397,N_2154,N_2533);
nor U3398 (N_3398,N_2908,N_2251);
and U3399 (N_3399,N_2982,N_2448);
and U3400 (N_3400,N_2886,N_2822);
nand U3401 (N_3401,N_2340,N_2939);
or U3402 (N_3402,N_2687,N_2686);
nor U3403 (N_3403,N_2705,N_2915);
and U3404 (N_3404,N_2798,N_2002);
nor U3405 (N_3405,N_2246,N_2124);
or U3406 (N_3406,N_2935,N_2672);
and U3407 (N_3407,N_2626,N_2068);
nor U3408 (N_3408,N_2855,N_2051);
nor U3409 (N_3409,N_2975,N_2420);
xor U3410 (N_3410,N_2470,N_2253);
nand U3411 (N_3411,N_2538,N_2573);
nand U3412 (N_3412,N_2858,N_2926);
nor U3413 (N_3413,N_2426,N_2012);
and U3414 (N_3414,N_2859,N_2585);
nand U3415 (N_3415,N_2102,N_2099);
or U3416 (N_3416,N_2767,N_2416);
and U3417 (N_3417,N_2777,N_2630);
and U3418 (N_3418,N_2106,N_2282);
or U3419 (N_3419,N_2377,N_2419);
nand U3420 (N_3420,N_2896,N_2085);
or U3421 (N_3421,N_2660,N_2379);
nand U3422 (N_3422,N_2454,N_2703);
or U3423 (N_3423,N_2880,N_2273);
nor U3424 (N_3424,N_2152,N_2486);
or U3425 (N_3425,N_2176,N_2728);
nor U3426 (N_3426,N_2351,N_2554);
and U3427 (N_3427,N_2725,N_2881);
and U3428 (N_3428,N_2281,N_2873);
nand U3429 (N_3429,N_2243,N_2279);
nand U3430 (N_3430,N_2592,N_2897);
nand U3431 (N_3431,N_2549,N_2745);
nand U3432 (N_3432,N_2516,N_2079);
nor U3433 (N_3433,N_2267,N_2670);
or U3434 (N_3434,N_2875,N_2096);
xor U3435 (N_3435,N_2676,N_2284);
nand U3436 (N_3436,N_2951,N_2941);
nor U3437 (N_3437,N_2831,N_2902);
nor U3438 (N_3438,N_2330,N_2727);
xnor U3439 (N_3439,N_2021,N_2375);
nand U3440 (N_3440,N_2523,N_2706);
or U3441 (N_3441,N_2888,N_2633);
nand U3442 (N_3442,N_2495,N_2921);
nor U3443 (N_3443,N_2813,N_2286);
and U3444 (N_3444,N_2013,N_2701);
nor U3445 (N_3445,N_2457,N_2368);
nor U3446 (N_3446,N_2431,N_2841);
and U3447 (N_3447,N_2572,N_2009);
nor U3448 (N_3448,N_2471,N_2034);
and U3449 (N_3449,N_2301,N_2699);
xnor U3450 (N_3450,N_2906,N_2242);
and U3451 (N_3451,N_2257,N_2241);
nor U3452 (N_3452,N_2872,N_2741);
nand U3453 (N_3453,N_2402,N_2924);
or U3454 (N_3454,N_2481,N_2228);
nand U3455 (N_3455,N_2948,N_2280);
nor U3456 (N_3456,N_2356,N_2797);
nand U3457 (N_3457,N_2700,N_2963);
or U3458 (N_3458,N_2042,N_2834);
and U3459 (N_3459,N_2661,N_2475);
and U3460 (N_3460,N_2576,N_2604);
and U3461 (N_3461,N_2401,N_2943);
or U3462 (N_3462,N_2365,N_2145);
and U3463 (N_3463,N_2987,N_2037);
nand U3464 (N_3464,N_2532,N_2593);
nor U3465 (N_3465,N_2498,N_2428);
and U3466 (N_3466,N_2913,N_2930);
nor U3467 (N_3467,N_2720,N_2958);
nand U3468 (N_3468,N_2238,N_2293);
nand U3469 (N_3469,N_2045,N_2336);
and U3470 (N_3470,N_2678,N_2123);
and U3471 (N_3471,N_2074,N_2946);
and U3472 (N_3472,N_2976,N_2161);
nand U3473 (N_3473,N_2233,N_2223);
or U3474 (N_3474,N_2001,N_2784);
nor U3475 (N_3475,N_2723,N_2217);
nand U3476 (N_3476,N_2137,N_2933);
nor U3477 (N_3477,N_2651,N_2737);
nor U3478 (N_3478,N_2505,N_2412);
and U3479 (N_3479,N_2579,N_2292);
nand U3480 (N_3480,N_2155,N_2929);
or U3481 (N_3481,N_2993,N_2887);
nand U3482 (N_3482,N_2198,N_2821);
xor U3483 (N_3483,N_2363,N_2640);
and U3484 (N_3484,N_2383,N_2066);
nor U3485 (N_3485,N_2690,N_2666);
nor U3486 (N_3486,N_2546,N_2860);
nand U3487 (N_3487,N_2294,N_2169);
or U3488 (N_3488,N_2776,N_2762);
xnor U3489 (N_3489,N_2005,N_2067);
nor U3490 (N_3490,N_2052,N_2792);
or U3491 (N_3491,N_2146,N_2805);
nand U3492 (N_3492,N_2461,N_2050);
and U3493 (N_3493,N_2341,N_2624);
nor U3494 (N_3494,N_2819,N_2040);
nand U3495 (N_3495,N_2520,N_2667);
nor U3496 (N_3496,N_2980,N_2159);
xnor U3497 (N_3497,N_2463,N_2614);
xor U3498 (N_3498,N_2999,N_2590);
and U3499 (N_3499,N_2455,N_2991);
and U3500 (N_3500,N_2072,N_2174);
nor U3501 (N_3501,N_2075,N_2250);
nand U3502 (N_3502,N_2642,N_2275);
nand U3503 (N_3503,N_2458,N_2409);
nor U3504 (N_3504,N_2972,N_2821);
nand U3505 (N_3505,N_2081,N_2662);
or U3506 (N_3506,N_2361,N_2833);
or U3507 (N_3507,N_2703,N_2569);
and U3508 (N_3508,N_2688,N_2572);
or U3509 (N_3509,N_2087,N_2828);
or U3510 (N_3510,N_2207,N_2521);
or U3511 (N_3511,N_2977,N_2465);
or U3512 (N_3512,N_2180,N_2696);
or U3513 (N_3513,N_2834,N_2154);
and U3514 (N_3514,N_2016,N_2686);
nand U3515 (N_3515,N_2495,N_2084);
nor U3516 (N_3516,N_2778,N_2498);
nand U3517 (N_3517,N_2970,N_2143);
or U3518 (N_3518,N_2194,N_2869);
or U3519 (N_3519,N_2451,N_2060);
and U3520 (N_3520,N_2782,N_2129);
nand U3521 (N_3521,N_2269,N_2450);
and U3522 (N_3522,N_2777,N_2474);
and U3523 (N_3523,N_2425,N_2238);
or U3524 (N_3524,N_2388,N_2437);
xor U3525 (N_3525,N_2709,N_2023);
nor U3526 (N_3526,N_2819,N_2413);
xnor U3527 (N_3527,N_2832,N_2973);
and U3528 (N_3528,N_2783,N_2673);
or U3529 (N_3529,N_2092,N_2658);
and U3530 (N_3530,N_2010,N_2227);
nor U3531 (N_3531,N_2264,N_2375);
nor U3532 (N_3532,N_2127,N_2409);
nor U3533 (N_3533,N_2218,N_2787);
and U3534 (N_3534,N_2962,N_2469);
and U3535 (N_3535,N_2068,N_2516);
nand U3536 (N_3536,N_2015,N_2133);
and U3537 (N_3537,N_2000,N_2060);
xor U3538 (N_3538,N_2837,N_2719);
and U3539 (N_3539,N_2164,N_2339);
and U3540 (N_3540,N_2473,N_2887);
nand U3541 (N_3541,N_2243,N_2407);
nor U3542 (N_3542,N_2274,N_2738);
or U3543 (N_3543,N_2228,N_2363);
nor U3544 (N_3544,N_2571,N_2723);
nor U3545 (N_3545,N_2742,N_2267);
and U3546 (N_3546,N_2306,N_2372);
nor U3547 (N_3547,N_2931,N_2778);
xor U3548 (N_3548,N_2368,N_2473);
or U3549 (N_3549,N_2815,N_2498);
xnor U3550 (N_3550,N_2307,N_2940);
or U3551 (N_3551,N_2943,N_2054);
and U3552 (N_3552,N_2575,N_2686);
and U3553 (N_3553,N_2866,N_2571);
or U3554 (N_3554,N_2090,N_2846);
nor U3555 (N_3555,N_2392,N_2689);
or U3556 (N_3556,N_2322,N_2176);
xnor U3557 (N_3557,N_2213,N_2546);
nor U3558 (N_3558,N_2499,N_2169);
and U3559 (N_3559,N_2940,N_2081);
or U3560 (N_3560,N_2700,N_2144);
and U3561 (N_3561,N_2500,N_2188);
nor U3562 (N_3562,N_2959,N_2067);
and U3563 (N_3563,N_2508,N_2172);
or U3564 (N_3564,N_2236,N_2189);
nor U3565 (N_3565,N_2224,N_2361);
nand U3566 (N_3566,N_2597,N_2712);
nor U3567 (N_3567,N_2483,N_2488);
nand U3568 (N_3568,N_2355,N_2915);
nor U3569 (N_3569,N_2627,N_2452);
nor U3570 (N_3570,N_2312,N_2482);
nand U3571 (N_3571,N_2863,N_2737);
and U3572 (N_3572,N_2278,N_2846);
or U3573 (N_3573,N_2779,N_2972);
and U3574 (N_3574,N_2008,N_2233);
nand U3575 (N_3575,N_2527,N_2608);
nor U3576 (N_3576,N_2677,N_2243);
and U3577 (N_3577,N_2055,N_2082);
xnor U3578 (N_3578,N_2846,N_2794);
nor U3579 (N_3579,N_2477,N_2070);
or U3580 (N_3580,N_2900,N_2444);
nand U3581 (N_3581,N_2922,N_2889);
nor U3582 (N_3582,N_2173,N_2942);
and U3583 (N_3583,N_2347,N_2286);
or U3584 (N_3584,N_2215,N_2681);
and U3585 (N_3585,N_2898,N_2220);
and U3586 (N_3586,N_2446,N_2761);
and U3587 (N_3587,N_2583,N_2740);
or U3588 (N_3588,N_2791,N_2586);
nor U3589 (N_3589,N_2011,N_2387);
nand U3590 (N_3590,N_2430,N_2608);
nor U3591 (N_3591,N_2879,N_2239);
or U3592 (N_3592,N_2250,N_2522);
and U3593 (N_3593,N_2506,N_2599);
xnor U3594 (N_3594,N_2929,N_2150);
and U3595 (N_3595,N_2623,N_2939);
nand U3596 (N_3596,N_2945,N_2869);
and U3597 (N_3597,N_2080,N_2651);
nor U3598 (N_3598,N_2829,N_2370);
and U3599 (N_3599,N_2944,N_2787);
or U3600 (N_3600,N_2572,N_2313);
nand U3601 (N_3601,N_2208,N_2282);
and U3602 (N_3602,N_2362,N_2804);
or U3603 (N_3603,N_2697,N_2131);
nor U3604 (N_3604,N_2455,N_2148);
xnor U3605 (N_3605,N_2840,N_2130);
nor U3606 (N_3606,N_2815,N_2067);
xor U3607 (N_3607,N_2985,N_2531);
and U3608 (N_3608,N_2051,N_2113);
and U3609 (N_3609,N_2133,N_2895);
and U3610 (N_3610,N_2569,N_2557);
nor U3611 (N_3611,N_2843,N_2501);
nand U3612 (N_3612,N_2468,N_2731);
nor U3613 (N_3613,N_2124,N_2839);
nand U3614 (N_3614,N_2095,N_2061);
and U3615 (N_3615,N_2173,N_2807);
or U3616 (N_3616,N_2299,N_2542);
and U3617 (N_3617,N_2551,N_2462);
xnor U3618 (N_3618,N_2289,N_2306);
or U3619 (N_3619,N_2989,N_2704);
nor U3620 (N_3620,N_2657,N_2895);
xnor U3621 (N_3621,N_2141,N_2262);
and U3622 (N_3622,N_2147,N_2761);
or U3623 (N_3623,N_2124,N_2853);
nor U3624 (N_3624,N_2113,N_2771);
and U3625 (N_3625,N_2289,N_2749);
or U3626 (N_3626,N_2983,N_2881);
and U3627 (N_3627,N_2796,N_2949);
or U3628 (N_3628,N_2616,N_2131);
nor U3629 (N_3629,N_2581,N_2368);
and U3630 (N_3630,N_2808,N_2990);
and U3631 (N_3631,N_2421,N_2255);
or U3632 (N_3632,N_2109,N_2108);
and U3633 (N_3633,N_2401,N_2106);
nand U3634 (N_3634,N_2416,N_2215);
or U3635 (N_3635,N_2686,N_2132);
or U3636 (N_3636,N_2854,N_2448);
and U3637 (N_3637,N_2565,N_2669);
or U3638 (N_3638,N_2324,N_2119);
nand U3639 (N_3639,N_2624,N_2599);
nand U3640 (N_3640,N_2850,N_2503);
nor U3641 (N_3641,N_2185,N_2416);
nor U3642 (N_3642,N_2561,N_2882);
or U3643 (N_3643,N_2470,N_2432);
nand U3644 (N_3644,N_2342,N_2078);
nand U3645 (N_3645,N_2179,N_2354);
nand U3646 (N_3646,N_2206,N_2834);
nor U3647 (N_3647,N_2126,N_2125);
and U3648 (N_3648,N_2118,N_2055);
and U3649 (N_3649,N_2264,N_2316);
nor U3650 (N_3650,N_2674,N_2073);
and U3651 (N_3651,N_2327,N_2007);
and U3652 (N_3652,N_2494,N_2866);
or U3653 (N_3653,N_2491,N_2716);
and U3654 (N_3654,N_2827,N_2603);
nor U3655 (N_3655,N_2371,N_2956);
nor U3656 (N_3656,N_2285,N_2553);
and U3657 (N_3657,N_2322,N_2689);
and U3658 (N_3658,N_2211,N_2164);
nor U3659 (N_3659,N_2574,N_2538);
nor U3660 (N_3660,N_2637,N_2880);
nand U3661 (N_3661,N_2834,N_2359);
and U3662 (N_3662,N_2935,N_2212);
or U3663 (N_3663,N_2066,N_2288);
nor U3664 (N_3664,N_2694,N_2691);
or U3665 (N_3665,N_2608,N_2308);
or U3666 (N_3666,N_2269,N_2138);
and U3667 (N_3667,N_2910,N_2294);
nand U3668 (N_3668,N_2025,N_2605);
xnor U3669 (N_3669,N_2735,N_2534);
or U3670 (N_3670,N_2958,N_2324);
and U3671 (N_3671,N_2806,N_2887);
xnor U3672 (N_3672,N_2834,N_2484);
and U3673 (N_3673,N_2479,N_2394);
nor U3674 (N_3674,N_2126,N_2974);
or U3675 (N_3675,N_2561,N_2467);
nand U3676 (N_3676,N_2479,N_2015);
nor U3677 (N_3677,N_2653,N_2241);
and U3678 (N_3678,N_2830,N_2257);
nor U3679 (N_3679,N_2495,N_2309);
xor U3680 (N_3680,N_2901,N_2281);
and U3681 (N_3681,N_2511,N_2956);
and U3682 (N_3682,N_2824,N_2955);
xor U3683 (N_3683,N_2484,N_2524);
nor U3684 (N_3684,N_2981,N_2422);
nor U3685 (N_3685,N_2819,N_2848);
and U3686 (N_3686,N_2000,N_2664);
or U3687 (N_3687,N_2009,N_2771);
nor U3688 (N_3688,N_2373,N_2998);
nand U3689 (N_3689,N_2571,N_2243);
nand U3690 (N_3690,N_2241,N_2056);
nand U3691 (N_3691,N_2912,N_2994);
nand U3692 (N_3692,N_2463,N_2010);
nor U3693 (N_3693,N_2959,N_2145);
and U3694 (N_3694,N_2350,N_2646);
and U3695 (N_3695,N_2373,N_2495);
and U3696 (N_3696,N_2970,N_2843);
nand U3697 (N_3697,N_2751,N_2599);
or U3698 (N_3698,N_2975,N_2217);
nor U3699 (N_3699,N_2852,N_2752);
nor U3700 (N_3700,N_2352,N_2825);
and U3701 (N_3701,N_2379,N_2026);
nor U3702 (N_3702,N_2165,N_2946);
nand U3703 (N_3703,N_2498,N_2378);
and U3704 (N_3704,N_2856,N_2101);
xnor U3705 (N_3705,N_2912,N_2074);
or U3706 (N_3706,N_2353,N_2047);
nor U3707 (N_3707,N_2760,N_2484);
nor U3708 (N_3708,N_2638,N_2922);
or U3709 (N_3709,N_2644,N_2391);
or U3710 (N_3710,N_2122,N_2882);
nand U3711 (N_3711,N_2429,N_2482);
or U3712 (N_3712,N_2471,N_2624);
nand U3713 (N_3713,N_2219,N_2602);
or U3714 (N_3714,N_2165,N_2364);
nor U3715 (N_3715,N_2232,N_2488);
nand U3716 (N_3716,N_2792,N_2328);
and U3717 (N_3717,N_2503,N_2424);
nor U3718 (N_3718,N_2276,N_2329);
or U3719 (N_3719,N_2819,N_2037);
nand U3720 (N_3720,N_2600,N_2991);
nor U3721 (N_3721,N_2172,N_2209);
nand U3722 (N_3722,N_2293,N_2484);
or U3723 (N_3723,N_2374,N_2434);
xor U3724 (N_3724,N_2130,N_2974);
nor U3725 (N_3725,N_2490,N_2003);
xor U3726 (N_3726,N_2241,N_2457);
xor U3727 (N_3727,N_2199,N_2545);
nand U3728 (N_3728,N_2086,N_2120);
and U3729 (N_3729,N_2889,N_2811);
nor U3730 (N_3730,N_2051,N_2985);
xnor U3731 (N_3731,N_2319,N_2479);
or U3732 (N_3732,N_2732,N_2444);
nand U3733 (N_3733,N_2011,N_2893);
nand U3734 (N_3734,N_2070,N_2701);
xnor U3735 (N_3735,N_2977,N_2760);
nand U3736 (N_3736,N_2088,N_2615);
nand U3737 (N_3737,N_2512,N_2936);
nor U3738 (N_3738,N_2202,N_2857);
and U3739 (N_3739,N_2900,N_2001);
or U3740 (N_3740,N_2642,N_2875);
and U3741 (N_3741,N_2757,N_2099);
or U3742 (N_3742,N_2179,N_2426);
nor U3743 (N_3743,N_2212,N_2072);
xor U3744 (N_3744,N_2759,N_2134);
and U3745 (N_3745,N_2588,N_2986);
and U3746 (N_3746,N_2901,N_2194);
nand U3747 (N_3747,N_2543,N_2822);
and U3748 (N_3748,N_2275,N_2006);
xnor U3749 (N_3749,N_2062,N_2514);
xor U3750 (N_3750,N_2586,N_2808);
or U3751 (N_3751,N_2642,N_2526);
nor U3752 (N_3752,N_2265,N_2862);
or U3753 (N_3753,N_2197,N_2845);
nand U3754 (N_3754,N_2206,N_2020);
or U3755 (N_3755,N_2576,N_2742);
nand U3756 (N_3756,N_2350,N_2337);
nand U3757 (N_3757,N_2889,N_2880);
xor U3758 (N_3758,N_2788,N_2271);
nand U3759 (N_3759,N_2632,N_2158);
nor U3760 (N_3760,N_2129,N_2957);
and U3761 (N_3761,N_2582,N_2136);
nand U3762 (N_3762,N_2074,N_2156);
and U3763 (N_3763,N_2853,N_2421);
nand U3764 (N_3764,N_2282,N_2442);
or U3765 (N_3765,N_2321,N_2430);
nor U3766 (N_3766,N_2985,N_2113);
or U3767 (N_3767,N_2806,N_2034);
nor U3768 (N_3768,N_2963,N_2780);
and U3769 (N_3769,N_2936,N_2472);
nor U3770 (N_3770,N_2131,N_2198);
nor U3771 (N_3771,N_2494,N_2661);
nor U3772 (N_3772,N_2625,N_2994);
nor U3773 (N_3773,N_2660,N_2216);
nor U3774 (N_3774,N_2039,N_2147);
or U3775 (N_3775,N_2948,N_2082);
xnor U3776 (N_3776,N_2785,N_2588);
or U3777 (N_3777,N_2807,N_2461);
xnor U3778 (N_3778,N_2879,N_2990);
nand U3779 (N_3779,N_2300,N_2378);
and U3780 (N_3780,N_2869,N_2527);
and U3781 (N_3781,N_2132,N_2682);
nor U3782 (N_3782,N_2964,N_2807);
nor U3783 (N_3783,N_2626,N_2423);
or U3784 (N_3784,N_2692,N_2696);
nor U3785 (N_3785,N_2760,N_2763);
nor U3786 (N_3786,N_2765,N_2624);
or U3787 (N_3787,N_2118,N_2738);
nand U3788 (N_3788,N_2329,N_2789);
nand U3789 (N_3789,N_2653,N_2979);
nand U3790 (N_3790,N_2566,N_2296);
nand U3791 (N_3791,N_2393,N_2021);
nor U3792 (N_3792,N_2044,N_2779);
or U3793 (N_3793,N_2878,N_2140);
or U3794 (N_3794,N_2020,N_2818);
or U3795 (N_3795,N_2394,N_2424);
and U3796 (N_3796,N_2524,N_2055);
and U3797 (N_3797,N_2558,N_2836);
xnor U3798 (N_3798,N_2006,N_2987);
and U3799 (N_3799,N_2611,N_2211);
and U3800 (N_3800,N_2070,N_2810);
nand U3801 (N_3801,N_2317,N_2033);
xnor U3802 (N_3802,N_2150,N_2060);
or U3803 (N_3803,N_2903,N_2524);
and U3804 (N_3804,N_2287,N_2954);
nand U3805 (N_3805,N_2823,N_2839);
nor U3806 (N_3806,N_2082,N_2419);
nor U3807 (N_3807,N_2752,N_2879);
nor U3808 (N_3808,N_2880,N_2768);
nor U3809 (N_3809,N_2344,N_2208);
xor U3810 (N_3810,N_2765,N_2572);
and U3811 (N_3811,N_2914,N_2494);
and U3812 (N_3812,N_2974,N_2190);
nand U3813 (N_3813,N_2732,N_2384);
nand U3814 (N_3814,N_2886,N_2489);
and U3815 (N_3815,N_2871,N_2725);
and U3816 (N_3816,N_2905,N_2615);
or U3817 (N_3817,N_2931,N_2729);
nor U3818 (N_3818,N_2283,N_2129);
nand U3819 (N_3819,N_2836,N_2659);
nor U3820 (N_3820,N_2808,N_2026);
xor U3821 (N_3821,N_2632,N_2709);
or U3822 (N_3822,N_2609,N_2652);
or U3823 (N_3823,N_2578,N_2977);
or U3824 (N_3824,N_2432,N_2259);
and U3825 (N_3825,N_2232,N_2571);
or U3826 (N_3826,N_2502,N_2874);
xor U3827 (N_3827,N_2647,N_2053);
nand U3828 (N_3828,N_2578,N_2270);
xnor U3829 (N_3829,N_2202,N_2597);
xor U3830 (N_3830,N_2706,N_2575);
and U3831 (N_3831,N_2802,N_2482);
nand U3832 (N_3832,N_2979,N_2257);
xnor U3833 (N_3833,N_2373,N_2800);
nand U3834 (N_3834,N_2127,N_2577);
or U3835 (N_3835,N_2459,N_2544);
and U3836 (N_3836,N_2404,N_2417);
and U3837 (N_3837,N_2319,N_2852);
nor U3838 (N_3838,N_2422,N_2532);
nor U3839 (N_3839,N_2384,N_2561);
nand U3840 (N_3840,N_2357,N_2921);
nor U3841 (N_3841,N_2361,N_2773);
nand U3842 (N_3842,N_2730,N_2598);
and U3843 (N_3843,N_2252,N_2429);
nor U3844 (N_3844,N_2890,N_2198);
and U3845 (N_3845,N_2909,N_2111);
xor U3846 (N_3846,N_2528,N_2865);
nor U3847 (N_3847,N_2243,N_2304);
nand U3848 (N_3848,N_2742,N_2700);
and U3849 (N_3849,N_2149,N_2717);
and U3850 (N_3850,N_2721,N_2873);
or U3851 (N_3851,N_2260,N_2694);
nor U3852 (N_3852,N_2096,N_2016);
xnor U3853 (N_3853,N_2818,N_2568);
nand U3854 (N_3854,N_2190,N_2243);
nand U3855 (N_3855,N_2369,N_2546);
xnor U3856 (N_3856,N_2457,N_2708);
or U3857 (N_3857,N_2173,N_2352);
nand U3858 (N_3858,N_2806,N_2698);
and U3859 (N_3859,N_2513,N_2715);
nor U3860 (N_3860,N_2765,N_2058);
and U3861 (N_3861,N_2844,N_2801);
nand U3862 (N_3862,N_2641,N_2254);
or U3863 (N_3863,N_2172,N_2681);
nand U3864 (N_3864,N_2364,N_2973);
or U3865 (N_3865,N_2761,N_2059);
and U3866 (N_3866,N_2765,N_2079);
nand U3867 (N_3867,N_2673,N_2238);
or U3868 (N_3868,N_2274,N_2005);
or U3869 (N_3869,N_2659,N_2441);
nor U3870 (N_3870,N_2466,N_2113);
nand U3871 (N_3871,N_2294,N_2944);
and U3872 (N_3872,N_2479,N_2475);
and U3873 (N_3873,N_2234,N_2755);
xnor U3874 (N_3874,N_2727,N_2368);
nand U3875 (N_3875,N_2723,N_2279);
and U3876 (N_3876,N_2089,N_2782);
or U3877 (N_3877,N_2974,N_2169);
nor U3878 (N_3878,N_2836,N_2613);
and U3879 (N_3879,N_2681,N_2613);
or U3880 (N_3880,N_2329,N_2274);
nand U3881 (N_3881,N_2598,N_2674);
nand U3882 (N_3882,N_2283,N_2338);
nand U3883 (N_3883,N_2602,N_2381);
or U3884 (N_3884,N_2843,N_2741);
xnor U3885 (N_3885,N_2017,N_2180);
nand U3886 (N_3886,N_2066,N_2632);
nand U3887 (N_3887,N_2722,N_2872);
and U3888 (N_3888,N_2557,N_2330);
xnor U3889 (N_3889,N_2989,N_2092);
nor U3890 (N_3890,N_2708,N_2728);
and U3891 (N_3891,N_2368,N_2518);
or U3892 (N_3892,N_2116,N_2729);
nand U3893 (N_3893,N_2381,N_2348);
and U3894 (N_3894,N_2033,N_2694);
nor U3895 (N_3895,N_2478,N_2804);
nor U3896 (N_3896,N_2727,N_2532);
and U3897 (N_3897,N_2271,N_2681);
nand U3898 (N_3898,N_2770,N_2997);
and U3899 (N_3899,N_2406,N_2499);
or U3900 (N_3900,N_2912,N_2552);
and U3901 (N_3901,N_2949,N_2937);
or U3902 (N_3902,N_2193,N_2937);
and U3903 (N_3903,N_2097,N_2286);
nand U3904 (N_3904,N_2524,N_2968);
nand U3905 (N_3905,N_2671,N_2856);
nand U3906 (N_3906,N_2569,N_2419);
nor U3907 (N_3907,N_2164,N_2892);
and U3908 (N_3908,N_2951,N_2536);
and U3909 (N_3909,N_2449,N_2629);
xor U3910 (N_3910,N_2082,N_2133);
or U3911 (N_3911,N_2528,N_2395);
or U3912 (N_3912,N_2963,N_2232);
nand U3913 (N_3913,N_2989,N_2012);
or U3914 (N_3914,N_2297,N_2746);
xor U3915 (N_3915,N_2878,N_2382);
or U3916 (N_3916,N_2767,N_2372);
or U3917 (N_3917,N_2945,N_2834);
xnor U3918 (N_3918,N_2902,N_2263);
nand U3919 (N_3919,N_2800,N_2047);
and U3920 (N_3920,N_2269,N_2728);
or U3921 (N_3921,N_2412,N_2276);
and U3922 (N_3922,N_2291,N_2441);
and U3923 (N_3923,N_2719,N_2978);
or U3924 (N_3924,N_2083,N_2768);
nand U3925 (N_3925,N_2189,N_2368);
nor U3926 (N_3926,N_2693,N_2989);
and U3927 (N_3927,N_2631,N_2578);
nand U3928 (N_3928,N_2845,N_2173);
or U3929 (N_3929,N_2220,N_2268);
xor U3930 (N_3930,N_2049,N_2721);
and U3931 (N_3931,N_2605,N_2374);
or U3932 (N_3932,N_2321,N_2716);
or U3933 (N_3933,N_2976,N_2363);
and U3934 (N_3934,N_2784,N_2556);
nand U3935 (N_3935,N_2939,N_2840);
nand U3936 (N_3936,N_2820,N_2855);
or U3937 (N_3937,N_2682,N_2208);
nor U3938 (N_3938,N_2307,N_2058);
nor U3939 (N_3939,N_2093,N_2575);
nand U3940 (N_3940,N_2512,N_2842);
nor U3941 (N_3941,N_2551,N_2496);
nor U3942 (N_3942,N_2651,N_2137);
nand U3943 (N_3943,N_2854,N_2311);
and U3944 (N_3944,N_2566,N_2915);
or U3945 (N_3945,N_2715,N_2869);
nor U3946 (N_3946,N_2729,N_2688);
or U3947 (N_3947,N_2472,N_2874);
xnor U3948 (N_3948,N_2278,N_2131);
and U3949 (N_3949,N_2584,N_2028);
nor U3950 (N_3950,N_2807,N_2915);
nor U3951 (N_3951,N_2127,N_2709);
nand U3952 (N_3952,N_2522,N_2084);
and U3953 (N_3953,N_2321,N_2755);
and U3954 (N_3954,N_2060,N_2360);
nand U3955 (N_3955,N_2121,N_2509);
or U3956 (N_3956,N_2610,N_2716);
nand U3957 (N_3957,N_2088,N_2528);
nand U3958 (N_3958,N_2509,N_2322);
nand U3959 (N_3959,N_2751,N_2863);
nand U3960 (N_3960,N_2939,N_2956);
nor U3961 (N_3961,N_2451,N_2401);
nand U3962 (N_3962,N_2780,N_2620);
nor U3963 (N_3963,N_2851,N_2618);
or U3964 (N_3964,N_2464,N_2843);
and U3965 (N_3965,N_2795,N_2189);
or U3966 (N_3966,N_2611,N_2585);
nand U3967 (N_3967,N_2996,N_2052);
and U3968 (N_3968,N_2634,N_2309);
and U3969 (N_3969,N_2226,N_2269);
nand U3970 (N_3970,N_2159,N_2117);
or U3971 (N_3971,N_2733,N_2136);
nor U3972 (N_3972,N_2015,N_2497);
nor U3973 (N_3973,N_2655,N_2109);
nand U3974 (N_3974,N_2750,N_2263);
or U3975 (N_3975,N_2659,N_2815);
and U3976 (N_3976,N_2043,N_2557);
or U3977 (N_3977,N_2450,N_2966);
or U3978 (N_3978,N_2424,N_2389);
nor U3979 (N_3979,N_2822,N_2960);
and U3980 (N_3980,N_2525,N_2701);
or U3981 (N_3981,N_2615,N_2248);
or U3982 (N_3982,N_2876,N_2508);
and U3983 (N_3983,N_2691,N_2968);
or U3984 (N_3984,N_2377,N_2528);
nor U3985 (N_3985,N_2963,N_2695);
and U3986 (N_3986,N_2301,N_2364);
nand U3987 (N_3987,N_2157,N_2072);
or U3988 (N_3988,N_2412,N_2472);
nor U3989 (N_3989,N_2897,N_2356);
and U3990 (N_3990,N_2227,N_2692);
or U3991 (N_3991,N_2185,N_2658);
or U3992 (N_3992,N_2748,N_2206);
nor U3993 (N_3993,N_2710,N_2106);
nand U3994 (N_3994,N_2593,N_2825);
nor U3995 (N_3995,N_2383,N_2959);
xor U3996 (N_3996,N_2032,N_2869);
xor U3997 (N_3997,N_2517,N_2819);
nor U3998 (N_3998,N_2747,N_2350);
nor U3999 (N_3999,N_2020,N_2420);
nand U4000 (N_4000,N_3257,N_3287);
nor U4001 (N_4001,N_3928,N_3546);
nand U4002 (N_4002,N_3249,N_3620);
nand U4003 (N_4003,N_3172,N_3899);
and U4004 (N_4004,N_3554,N_3777);
nand U4005 (N_4005,N_3232,N_3355);
or U4006 (N_4006,N_3411,N_3216);
or U4007 (N_4007,N_3146,N_3823);
nand U4008 (N_4008,N_3154,N_3288);
nor U4009 (N_4009,N_3119,N_3342);
and U4010 (N_4010,N_3908,N_3965);
xor U4011 (N_4011,N_3260,N_3785);
nand U4012 (N_4012,N_3212,N_3250);
and U4013 (N_4013,N_3802,N_3158);
and U4014 (N_4014,N_3023,N_3134);
xnor U4015 (N_4015,N_3649,N_3731);
or U4016 (N_4016,N_3383,N_3251);
xnor U4017 (N_4017,N_3289,N_3660);
and U4018 (N_4018,N_3892,N_3078);
or U4019 (N_4019,N_3780,N_3829);
and U4020 (N_4020,N_3306,N_3711);
and U4021 (N_4021,N_3324,N_3339);
and U4022 (N_4022,N_3644,N_3227);
nor U4023 (N_4023,N_3922,N_3063);
nor U4024 (N_4024,N_3416,N_3656);
and U4025 (N_4025,N_3543,N_3203);
or U4026 (N_4026,N_3812,N_3431);
xnor U4027 (N_4027,N_3748,N_3944);
and U4028 (N_4028,N_3394,N_3261);
or U4029 (N_4029,N_3076,N_3448);
nor U4030 (N_4030,N_3304,N_3198);
xnor U4031 (N_4031,N_3327,N_3204);
nor U4032 (N_4032,N_3523,N_3853);
or U4033 (N_4033,N_3437,N_3915);
and U4034 (N_4034,N_3498,N_3841);
and U4035 (N_4035,N_3599,N_3640);
and U4036 (N_4036,N_3987,N_3643);
and U4037 (N_4037,N_3392,N_3461);
nor U4038 (N_4038,N_3292,N_3947);
and U4039 (N_4039,N_3894,N_3704);
and U4040 (N_4040,N_3440,N_3809);
nor U4041 (N_4041,N_3091,N_3627);
nor U4042 (N_4042,N_3034,N_3576);
and U4043 (N_4043,N_3485,N_3037);
nor U4044 (N_4044,N_3079,N_3560);
nor U4045 (N_4045,N_3558,N_3487);
or U4046 (N_4046,N_3848,N_3343);
xnor U4047 (N_4047,N_3021,N_3492);
or U4048 (N_4048,N_3329,N_3563);
and U4049 (N_4049,N_3345,N_3028);
nand U4050 (N_4050,N_3067,N_3265);
and U4051 (N_4051,N_3208,N_3629);
nor U4052 (N_4052,N_3992,N_3990);
and U4053 (N_4053,N_3321,N_3226);
xnor U4054 (N_4054,N_3835,N_3156);
nor U4055 (N_4055,N_3150,N_3976);
xnor U4056 (N_4056,N_3542,N_3065);
or U4057 (N_4057,N_3273,N_3458);
and U4058 (N_4058,N_3998,N_3513);
nor U4059 (N_4059,N_3775,N_3594);
xnor U4060 (N_4060,N_3387,N_3564);
nor U4061 (N_4061,N_3732,N_3259);
and U4062 (N_4062,N_3282,N_3057);
nor U4063 (N_4063,N_3141,N_3167);
nand U4064 (N_4064,N_3147,N_3330);
and U4065 (N_4065,N_3223,N_3791);
xor U4066 (N_4066,N_3420,N_3493);
nor U4067 (N_4067,N_3544,N_3967);
and U4068 (N_4068,N_3462,N_3618);
nor U4069 (N_4069,N_3230,N_3982);
and U4070 (N_4070,N_3932,N_3478);
or U4071 (N_4071,N_3938,N_3789);
nand U4072 (N_4072,N_3665,N_3765);
or U4073 (N_4073,N_3984,N_3929);
or U4074 (N_4074,N_3733,N_3476);
xnor U4075 (N_4075,N_3397,N_3913);
and U4076 (N_4076,N_3676,N_3041);
nand U4077 (N_4077,N_3298,N_3657);
nor U4078 (N_4078,N_3426,N_3309);
nand U4079 (N_4079,N_3299,N_3547);
or U4080 (N_4080,N_3975,N_3744);
nand U4081 (N_4081,N_3926,N_3541);
nand U4082 (N_4082,N_3334,N_3969);
nand U4083 (N_4083,N_3830,N_3441);
or U4084 (N_4084,N_3845,N_3794);
nor U4085 (N_4085,N_3677,N_3589);
xor U4086 (N_4086,N_3127,N_3055);
or U4087 (N_4087,N_3625,N_3857);
or U4088 (N_4088,N_3503,N_3593);
or U4089 (N_4089,N_3601,N_3362);
and U4090 (N_4090,N_3070,N_3693);
xnor U4091 (N_4091,N_3798,N_3453);
and U4092 (N_4092,N_3140,N_3116);
nor U4093 (N_4093,N_3105,N_3702);
or U4094 (N_4094,N_3528,N_3066);
and U4095 (N_4095,N_3222,N_3778);
nor U4096 (N_4096,N_3524,N_3169);
nor U4097 (N_4097,N_3717,N_3590);
and U4098 (N_4098,N_3782,N_3470);
and U4099 (N_4099,N_3201,N_3132);
nor U4100 (N_4100,N_3696,N_3698);
nor U4101 (N_4101,N_3253,N_3758);
xnor U4102 (N_4102,N_3876,N_3194);
nor U4103 (N_4103,N_3851,N_3786);
and U4104 (N_4104,N_3945,N_3122);
nand U4105 (N_4105,N_3935,N_3395);
or U4106 (N_4106,N_3166,N_3549);
nor U4107 (N_4107,N_3059,N_3805);
nor U4108 (N_4108,N_3400,N_3797);
nor U4109 (N_4109,N_3774,N_3190);
or U4110 (N_4110,N_3999,N_3189);
and U4111 (N_4111,N_3019,N_3866);
nor U4112 (N_4112,N_3772,N_3391);
and U4113 (N_4113,N_3377,N_3526);
or U4114 (N_4114,N_3511,N_3165);
xor U4115 (N_4115,N_3779,N_3701);
xor U4116 (N_4116,N_3887,N_3946);
nand U4117 (N_4117,N_3556,N_3636);
nor U4118 (N_4118,N_3096,N_3923);
nand U4119 (N_4119,N_3270,N_3068);
nand U4120 (N_4120,N_3597,N_3358);
or U4121 (N_4121,N_3489,N_3705);
and U4122 (N_4122,N_3691,N_3767);
or U4123 (N_4123,N_3860,N_3678);
xor U4124 (N_4124,N_3628,N_3981);
and U4125 (N_4125,N_3181,N_3592);
or U4126 (N_4126,N_3726,N_3171);
nand U4127 (N_4127,N_3410,N_3720);
xor U4128 (N_4128,N_3684,N_3750);
nand U4129 (N_4129,N_3415,N_3124);
nand U4130 (N_4130,N_3813,N_3266);
or U4131 (N_4131,N_3084,N_3173);
and U4132 (N_4132,N_3854,N_3514);
nand U4133 (N_4133,N_3714,N_3933);
or U4134 (N_4134,N_3648,N_3904);
nor U4135 (N_4135,N_3615,N_3865);
xor U4136 (N_4136,N_3793,N_3344);
or U4137 (N_4137,N_3583,N_3195);
nor U4138 (N_4138,N_3252,N_3905);
and U4139 (N_4139,N_3241,N_3637);
xor U4140 (N_4140,N_3533,N_3425);
xor U4141 (N_4141,N_3634,N_3930);
or U4142 (N_4142,N_3182,N_3090);
or U4143 (N_4143,N_3529,N_3495);
xor U4144 (N_4144,N_3099,N_3418);
and U4145 (N_4145,N_3092,N_3776);
xnor U4146 (N_4146,N_3010,N_3246);
and U4147 (N_4147,N_3510,N_3332);
or U4148 (N_4148,N_3402,N_3742);
or U4149 (N_4149,N_3484,N_3584);
or U4150 (N_4150,N_3110,N_3109);
or U4151 (N_4151,N_3995,N_3029);
nand U4152 (N_4152,N_3032,N_3550);
nand U4153 (N_4153,N_3294,N_3404);
nor U4154 (N_4154,N_3821,N_3569);
or U4155 (N_4155,N_3434,N_3356);
or U4156 (N_4156,N_3910,N_3471);
or U4157 (N_4157,N_3046,N_3061);
nor U4158 (N_4158,N_3459,N_3650);
nor U4159 (N_4159,N_3113,N_3423);
nor U4160 (N_4160,N_3697,N_3228);
or U4161 (N_4161,N_3752,N_3341);
nand U4162 (N_4162,N_3325,N_3145);
nand U4163 (N_4163,N_3371,N_3421);
and U4164 (N_4164,N_3308,N_3472);
and U4165 (N_4165,N_3011,N_3924);
nor U4166 (N_4166,N_3429,N_3960);
nand U4167 (N_4167,N_3517,N_3388);
or U4168 (N_4168,N_3316,N_3357);
nor U4169 (N_4169,N_3667,N_3483);
or U4170 (N_4170,N_3931,N_3218);
xnor U4171 (N_4171,N_3559,N_3381);
or U4172 (N_4172,N_3346,N_3837);
nor U4173 (N_4173,N_3438,N_3571);
and U4174 (N_4174,N_3219,N_3762);
and U4175 (N_4175,N_3211,N_3681);
nand U4176 (N_4176,N_3846,N_3401);
nand U4177 (N_4177,N_3598,N_3300);
nand U4178 (N_4178,N_3670,N_3467);
or U4179 (N_4179,N_3235,N_3700);
and U4180 (N_4180,N_3602,N_3985);
and U4181 (N_4181,N_3269,N_3446);
or U4182 (N_4182,N_3000,N_3902);
nand U4183 (N_4183,N_3885,N_3532);
or U4184 (N_4184,N_3530,N_3534);
and U4185 (N_4185,N_3445,N_3961);
or U4186 (N_4186,N_3281,N_3687);
xnor U4187 (N_4187,N_3311,N_3539);
or U4188 (N_4188,N_3314,N_3364);
and U4189 (N_4189,N_3663,N_3280);
and U4190 (N_4190,N_3002,N_3808);
nand U4191 (N_4191,N_3035,N_3608);
nor U4192 (N_4192,N_3380,N_3536);
nor U4193 (N_4193,N_3595,N_3499);
or U4194 (N_4194,N_3365,N_3614);
and U4195 (N_4195,N_3831,N_3879);
nand U4196 (N_4196,N_3340,N_3062);
or U4197 (N_4197,N_3896,N_3137);
xnor U4198 (N_4198,N_3112,N_3015);
nor U4199 (N_4199,N_3163,N_3582);
nand U4200 (N_4200,N_3213,N_3801);
nand U4201 (N_4201,N_3966,N_3638);
nor U4202 (N_4202,N_3540,N_3473);
nand U4203 (N_4203,N_3087,N_3690);
and U4204 (N_4204,N_3297,N_3979);
or U4205 (N_4205,N_3822,N_3954);
nand U4206 (N_4206,N_3565,N_3085);
and U4207 (N_4207,N_3326,N_3399);
and U4208 (N_4208,N_3175,N_3725);
nor U4209 (N_4209,N_3054,N_3243);
and U4210 (N_4210,N_3825,N_3939);
nor U4211 (N_4211,N_3086,N_3052);
nand U4212 (N_4212,N_3474,N_3274);
or U4213 (N_4213,N_3012,N_3502);
nand U4214 (N_4214,N_3941,N_3631);
or U4215 (N_4215,N_3898,N_3736);
nor U4216 (N_4216,N_3414,N_3180);
nand U4217 (N_4217,N_3844,N_3570);
nand U4218 (N_4218,N_3433,N_3895);
nand U4219 (N_4219,N_3828,N_3217);
and U4220 (N_4220,N_3196,N_3008);
and U4221 (N_4221,N_3031,N_3361);
or U4222 (N_4222,N_3973,N_3500);
nand U4223 (N_4223,N_3537,N_3375);
and U4224 (N_4224,N_3385,N_3347);
nand U4225 (N_4225,N_3111,N_3174);
and U4226 (N_4226,N_3221,N_3064);
nor U4227 (N_4227,N_3275,N_3911);
nand U4228 (N_4228,N_3318,N_3125);
nand U4229 (N_4229,N_3100,N_3220);
nor U4230 (N_4230,N_3465,N_3735);
and U4231 (N_4231,N_3396,N_3408);
or U4232 (N_4232,N_3293,N_3768);
nand U4233 (N_4233,N_3291,N_3655);
nor U4234 (N_4234,N_3186,N_3215);
nor U4235 (N_4235,N_3501,N_3873);
or U4236 (N_4236,N_3679,N_3382);
nand U4237 (N_4237,N_3143,N_3026);
nor U4238 (N_4238,N_3353,N_3089);
nor U4239 (N_4239,N_3464,N_3335);
and U4240 (N_4240,N_3551,N_3136);
xnor U4241 (N_4241,N_3024,N_3160);
nor U4242 (N_4242,N_3950,N_3814);
and U4243 (N_4243,N_3680,N_3925);
or U4244 (N_4244,N_3914,N_3977);
nor U4245 (N_4245,N_3454,N_3578);
or U4246 (N_4246,N_3295,N_3001);
and U4247 (N_4247,N_3242,N_3872);
or U4248 (N_4248,N_3386,N_3897);
and U4249 (N_4249,N_3117,N_3760);
or U4250 (N_4250,N_3622,N_3206);
or U4251 (N_4251,N_3949,N_3527);
nor U4252 (N_4252,N_3191,N_3393);
and U4253 (N_4253,N_3197,N_3888);
and U4254 (N_4254,N_3942,N_3372);
or U4255 (N_4255,N_3018,N_3943);
and U4256 (N_4256,N_3900,N_3322);
or U4257 (N_4257,N_3210,N_3451);
and U4258 (N_4258,N_3607,N_3972);
nor U4259 (N_4259,N_3713,N_3267);
and U4260 (N_4260,N_3020,N_3682);
or U4261 (N_4261,N_3447,N_3811);
xnor U4262 (N_4262,N_3766,N_3104);
and U4263 (N_4263,N_3738,N_3310);
xor U4264 (N_4264,N_3138,N_3955);
and U4265 (N_4265,N_3368,N_3818);
xnor U4266 (N_4266,N_3722,N_3795);
xnor U4267 (N_4267,N_3192,N_3097);
nor U4268 (N_4268,N_3820,N_3600);
nand U4269 (N_4269,N_3016,N_3148);
nor U4270 (N_4270,N_3286,N_3225);
nand U4271 (N_4271,N_3989,N_3053);
nor U4272 (N_4272,N_3773,N_3139);
or U4273 (N_4273,N_3787,N_3033);
or U4274 (N_4274,N_3477,N_3918);
xnor U4275 (N_4275,N_3877,N_3452);
and U4276 (N_4276,N_3179,N_3048);
or U4277 (N_4277,N_3479,N_3610);
or U4278 (N_4278,N_3200,N_3359);
nand U4279 (N_4279,N_3756,N_3834);
nand U4280 (N_4280,N_3840,N_3229);
or U4281 (N_4281,N_3460,N_3666);
or U4282 (N_4282,N_3991,N_3102);
nand U4283 (N_4283,N_3604,N_3727);
and U4284 (N_4284,N_3135,N_3639);
nor U4285 (N_4285,N_3443,N_3348);
or U4286 (N_4286,N_3870,N_3168);
or U4287 (N_4287,N_3716,N_3964);
and U4288 (N_4288,N_3207,N_3968);
nand U4289 (N_4289,N_3504,N_3729);
or U4290 (N_4290,N_3646,N_3161);
or U4291 (N_4291,N_3611,N_3074);
nor U4292 (N_4292,N_3237,N_3612);
or U4293 (N_4293,N_3370,N_3686);
nand U4294 (N_4294,N_3893,N_3036);
and U4295 (N_4295,N_3863,N_3264);
xnor U4296 (N_4296,N_3781,N_3296);
xor U4297 (N_4297,N_3996,N_3757);
or U4298 (N_4298,N_3997,N_3069);
xor U4299 (N_4299,N_3328,N_3839);
nand U4300 (N_4300,N_3959,N_3424);
or U4301 (N_4301,N_3800,N_3552);
nor U4302 (N_4302,N_3350,N_3632);
or U4303 (N_4303,N_3715,N_3689);
xnor U4304 (N_4304,N_3878,N_3337);
nor U4305 (N_4305,N_3613,N_3919);
and U4306 (N_4306,N_3248,N_3520);
or U4307 (N_4307,N_3567,N_3624);
and U4308 (N_4308,N_3307,N_3609);
and U4309 (N_4309,N_3022,N_3121);
or U4310 (N_4310,N_3419,N_3816);
nand U4311 (N_4311,N_3784,N_3792);
nor U4312 (N_4312,N_3412,N_3014);
nand U4313 (N_4313,N_3349,N_3149);
or U4314 (N_4314,N_3317,N_3566);
nand U4315 (N_4315,N_3754,N_3626);
nor U4316 (N_4316,N_3255,N_3710);
and U4317 (N_4317,N_3858,N_3668);
nand U4318 (N_4318,N_3155,N_3422);
or U4319 (N_4319,N_3098,N_3247);
nand U4320 (N_4320,N_3616,N_3561);
or U4321 (N_4321,N_3262,N_3788);
nand U4322 (N_4322,N_3747,N_3491);
nor U4323 (N_4323,N_3301,N_3662);
nand U4324 (N_4324,N_3940,N_3849);
nand U4325 (N_4325,N_3374,N_3586);
and U4326 (N_4326,N_3151,N_3882);
and U4327 (N_4327,N_3367,N_3993);
nor U4328 (N_4328,N_3581,N_3005);
or U4329 (N_4329,N_3506,N_3706);
nor U4330 (N_4330,N_3129,N_3231);
or U4331 (N_4331,N_3512,N_3468);
nor U4332 (N_4332,N_3436,N_3469);
nor U4333 (N_4333,N_3994,N_3585);
nand U4334 (N_4334,N_3623,N_3077);
or U4335 (N_4335,N_3130,N_3661);
nor U4336 (N_4336,N_3088,N_3373);
xnor U4337 (N_4337,N_3633,N_3009);
or U4338 (N_4338,N_3508,N_3859);
and U4339 (N_4339,N_3323,N_3674);
or U4340 (N_4340,N_3336,N_3951);
and U4341 (N_4341,N_3183,N_3177);
or U4342 (N_4342,N_3912,N_3695);
nand U4343 (N_4343,N_3804,N_3038);
xor U4344 (N_4344,N_3741,N_3745);
or U4345 (N_4345,N_3376,N_3770);
xor U4346 (N_4346,N_3783,N_3043);
or U4347 (N_4347,N_3664,N_3619);
or U4348 (N_4348,N_3574,N_3120);
xor U4349 (N_4349,N_3963,N_3379);
or U4350 (N_4350,N_3060,N_3115);
nand U4351 (N_4351,N_3279,N_3004);
or U4352 (N_4352,N_3980,N_3101);
and U4353 (N_4353,N_3003,N_3621);
or U4354 (N_4354,N_3759,N_3852);
xor U4355 (N_4355,N_3806,N_3118);
nand U4356 (N_4356,N_3916,N_3427);
or U4357 (N_4357,N_3958,N_3013);
and U4358 (N_4358,N_3413,N_3490);
and U4359 (N_4359,N_3952,N_3833);
or U4360 (N_4360,N_3647,N_3901);
xnor U4361 (N_4361,N_3093,N_3824);
nand U4362 (N_4362,N_3268,N_3538);
and U4363 (N_4363,N_3974,N_3187);
and U4364 (N_4364,N_3836,N_3214);
nand U4365 (N_4365,N_3724,N_3103);
or U4366 (N_4366,N_3861,N_3058);
nand U4367 (N_4367,N_3548,N_3428);
and U4368 (N_4368,N_3692,N_3719);
nand U4369 (N_4369,N_3290,N_3790);
nor U4370 (N_4370,N_3703,N_3236);
xor U4371 (N_4371,N_3707,N_3338);
and U4372 (N_4372,N_3557,N_3525);
or U4373 (N_4373,N_3838,N_3988);
nor U4374 (N_4374,N_3606,N_3176);
nor U4375 (N_4375,N_3193,N_3114);
nor U4376 (N_4376,N_3740,N_3108);
nor U4377 (N_4377,N_3083,N_3708);
nor U4378 (N_4378,N_3039,N_3807);
nand U4379 (N_4379,N_3868,N_3164);
nand U4380 (N_4380,N_3044,N_3856);
and U4381 (N_4381,N_3763,N_3234);
nor U4382 (N_4382,N_3568,N_3843);
nand U4383 (N_4383,N_3683,N_3170);
and U4384 (N_4384,N_3285,N_3771);
or U4385 (N_4385,N_3407,N_3723);
and U4386 (N_4386,N_3751,N_3050);
and U4387 (N_4387,N_3755,N_3588);
nand U4388 (N_4388,N_3354,N_3934);
nor U4389 (N_4389,N_3986,N_3435);
nand U4390 (N_4390,N_3577,N_3743);
nor U4391 (N_4391,N_3535,N_3030);
and U4392 (N_4392,N_3737,N_3749);
and U4393 (N_4393,N_3669,N_3482);
nor U4394 (N_4394,N_3953,N_3718);
nor U4395 (N_4395,N_3475,N_3254);
nand U4396 (N_4396,N_3486,N_3764);
and U4397 (N_4397,N_3047,N_3403);
or U4398 (N_4398,N_3185,N_3730);
nand U4399 (N_4399,N_3072,N_3305);
nand U4400 (N_4400,N_3283,N_3398);
or U4401 (N_4401,N_3983,N_3591);
and U4402 (N_4402,N_3017,N_3258);
and U4403 (N_4403,N_3157,N_3244);
or U4404 (N_4404,N_3886,N_3796);
nor U4405 (N_4405,N_3095,N_3871);
or U4406 (N_4406,N_3494,N_3579);
nand U4407 (N_4407,N_3936,N_3430);
and U4408 (N_4408,N_3874,N_3761);
xnor U4409 (N_4409,N_3366,N_3128);
or U4410 (N_4410,N_3442,N_3880);
nor U4411 (N_4411,N_3082,N_3466);
nand U4412 (N_4412,N_3653,N_3094);
and U4413 (N_4413,N_3144,N_3921);
or U4414 (N_4414,N_3555,N_3685);
nand U4415 (N_4415,N_3042,N_3051);
or U4416 (N_4416,N_3562,N_3378);
and U4417 (N_4417,N_3071,N_3675);
nor U4418 (N_4418,N_3842,N_3572);
and U4419 (N_4419,N_3688,N_3862);
nor U4420 (N_4420,N_3654,N_3850);
and U4421 (N_4421,N_3753,N_3746);
nor U4422 (N_4422,N_3521,N_3927);
nor U4423 (N_4423,N_3488,N_3153);
and U4424 (N_4424,N_3457,N_3651);
nand U4425 (N_4425,N_3224,N_3439);
xnor U4426 (N_4426,N_3652,N_3505);
nor U4427 (N_4427,N_3815,N_3970);
nand U4428 (N_4428,N_3962,N_3271);
or U4429 (N_4429,N_3417,N_3178);
nor U4430 (N_4430,N_3580,N_3699);
nor U4431 (N_4431,N_3320,N_3075);
nor U4432 (N_4432,N_3481,N_3956);
nand U4433 (N_4433,N_3277,N_3238);
and U4434 (N_4434,N_3480,N_3497);
nand U4435 (N_4435,N_3957,N_3883);
nor U4436 (N_4436,N_3199,N_3162);
and U4437 (N_4437,N_3363,N_3889);
nor U4438 (N_4438,N_3603,N_3073);
and U4439 (N_4439,N_3331,N_3025);
and U4440 (N_4440,N_3769,N_3721);
or U4441 (N_4441,N_3081,N_3906);
or U4442 (N_4442,N_3106,N_3312);
nand U4443 (N_4443,N_3673,N_3630);
nor U4444 (N_4444,N_3126,N_3658);
xnor U4445 (N_4445,N_3184,N_3390);
or U4446 (N_4446,N_3496,N_3909);
nor U4447 (N_4447,N_3333,N_3855);
or U4448 (N_4448,N_3006,N_3867);
xnor U4449 (N_4449,N_3573,N_3739);
nand U4450 (N_4450,N_3864,N_3937);
and U4451 (N_4451,N_3827,N_3152);
or U4452 (N_4452,N_3881,N_3007);
xor U4453 (N_4453,N_3409,N_3803);
and U4454 (N_4454,N_3728,N_3659);
or U4455 (N_4455,N_3245,N_3617);
and U4456 (N_4456,N_3384,N_3891);
or U4457 (N_4457,N_3389,N_3056);
nor U4458 (N_4458,N_3522,N_3832);
nand U4459 (N_4459,N_3531,N_3272);
and U4460 (N_4460,N_3971,N_3712);
nor U4461 (N_4461,N_3635,N_3515);
nand U4462 (N_4462,N_3507,N_3645);
nor U4463 (N_4463,N_3303,N_3455);
nand U4464 (N_4464,N_3826,N_3575);
and U4465 (N_4465,N_3672,N_3907);
nor U4466 (N_4466,N_3641,N_3819);
or U4467 (N_4467,N_3123,N_3205);
nand U4468 (N_4468,N_3319,N_3456);
and U4469 (N_4469,N_3159,N_3587);
xnor U4470 (N_4470,N_3516,N_3920);
nor U4471 (N_4471,N_3545,N_3045);
or U4472 (N_4472,N_3049,N_3903);
xnor U4473 (N_4473,N_3133,N_3278);
or U4474 (N_4474,N_3360,N_3817);
and U4475 (N_4475,N_3694,N_3405);
and U4476 (N_4476,N_3596,N_3369);
nor U4477 (N_4477,N_3709,N_3142);
and U4478 (N_4478,N_3948,N_3463);
nand U4479 (N_4479,N_3209,N_3799);
xnor U4480 (N_4480,N_3509,N_3642);
or U4481 (N_4481,N_3884,N_3734);
and U4482 (N_4482,N_3263,N_3352);
and U4483 (N_4483,N_3406,N_3313);
xor U4484 (N_4484,N_3027,N_3875);
or U4485 (N_4485,N_3450,N_3302);
or U4486 (N_4486,N_3890,N_3671);
or U4487 (N_4487,N_3276,N_3810);
nand U4488 (N_4488,N_3080,N_3847);
nor U4489 (N_4489,N_3107,N_3188);
or U4490 (N_4490,N_3444,N_3553);
and U4491 (N_4491,N_3869,N_3519);
nand U4492 (N_4492,N_3233,N_3978);
and U4493 (N_4493,N_3351,N_3240);
xnor U4494 (N_4494,N_3131,N_3284);
nor U4495 (N_4495,N_3449,N_3315);
nor U4496 (N_4496,N_3605,N_3040);
or U4497 (N_4497,N_3432,N_3256);
xor U4498 (N_4498,N_3917,N_3202);
nor U4499 (N_4499,N_3518,N_3239);
or U4500 (N_4500,N_3547,N_3770);
or U4501 (N_4501,N_3503,N_3355);
xnor U4502 (N_4502,N_3196,N_3264);
and U4503 (N_4503,N_3239,N_3022);
or U4504 (N_4504,N_3450,N_3103);
nor U4505 (N_4505,N_3384,N_3813);
nor U4506 (N_4506,N_3331,N_3918);
nand U4507 (N_4507,N_3767,N_3261);
and U4508 (N_4508,N_3013,N_3642);
or U4509 (N_4509,N_3197,N_3489);
nand U4510 (N_4510,N_3634,N_3050);
nand U4511 (N_4511,N_3872,N_3141);
nor U4512 (N_4512,N_3357,N_3374);
and U4513 (N_4513,N_3591,N_3690);
xnor U4514 (N_4514,N_3793,N_3846);
nand U4515 (N_4515,N_3442,N_3561);
and U4516 (N_4516,N_3396,N_3221);
or U4517 (N_4517,N_3677,N_3114);
or U4518 (N_4518,N_3920,N_3963);
nand U4519 (N_4519,N_3894,N_3314);
nand U4520 (N_4520,N_3954,N_3690);
or U4521 (N_4521,N_3515,N_3734);
and U4522 (N_4522,N_3141,N_3274);
or U4523 (N_4523,N_3520,N_3636);
and U4524 (N_4524,N_3364,N_3670);
or U4525 (N_4525,N_3523,N_3869);
nand U4526 (N_4526,N_3823,N_3203);
and U4527 (N_4527,N_3885,N_3905);
nor U4528 (N_4528,N_3161,N_3337);
xor U4529 (N_4529,N_3667,N_3115);
and U4530 (N_4530,N_3391,N_3612);
nor U4531 (N_4531,N_3549,N_3692);
nor U4532 (N_4532,N_3738,N_3776);
and U4533 (N_4533,N_3779,N_3284);
and U4534 (N_4534,N_3955,N_3153);
nor U4535 (N_4535,N_3064,N_3202);
nor U4536 (N_4536,N_3147,N_3180);
or U4537 (N_4537,N_3170,N_3530);
or U4538 (N_4538,N_3562,N_3115);
nor U4539 (N_4539,N_3630,N_3396);
nor U4540 (N_4540,N_3559,N_3607);
nand U4541 (N_4541,N_3047,N_3056);
nor U4542 (N_4542,N_3891,N_3912);
nor U4543 (N_4543,N_3373,N_3300);
nor U4544 (N_4544,N_3420,N_3174);
nor U4545 (N_4545,N_3286,N_3317);
or U4546 (N_4546,N_3668,N_3295);
and U4547 (N_4547,N_3638,N_3849);
nor U4548 (N_4548,N_3031,N_3553);
and U4549 (N_4549,N_3137,N_3975);
nand U4550 (N_4550,N_3424,N_3040);
and U4551 (N_4551,N_3367,N_3067);
nand U4552 (N_4552,N_3001,N_3972);
nor U4553 (N_4553,N_3542,N_3483);
and U4554 (N_4554,N_3781,N_3912);
nand U4555 (N_4555,N_3549,N_3982);
xor U4556 (N_4556,N_3770,N_3301);
and U4557 (N_4557,N_3881,N_3106);
xor U4558 (N_4558,N_3498,N_3605);
nand U4559 (N_4559,N_3392,N_3237);
and U4560 (N_4560,N_3863,N_3786);
and U4561 (N_4561,N_3447,N_3908);
or U4562 (N_4562,N_3432,N_3508);
or U4563 (N_4563,N_3033,N_3140);
and U4564 (N_4564,N_3122,N_3148);
nand U4565 (N_4565,N_3337,N_3873);
nand U4566 (N_4566,N_3807,N_3419);
xor U4567 (N_4567,N_3620,N_3217);
and U4568 (N_4568,N_3806,N_3151);
nor U4569 (N_4569,N_3221,N_3003);
and U4570 (N_4570,N_3355,N_3476);
nand U4571 (N_4571,N_3757,N_3768);
nand U4572 (N_4572,N_3959,N_3373);
nand U4573 (N_4573,N_3214,N_3410);
xnor U4574 (N_4574,N_3711,N_3331);
nor U4575 (N_4575,N_3991,N_3278);
nor U4576 (N_4576,N_3204,N_3218);
or U4577 (N_4577,N_3834,N_3918);
or U4578 (N_4578,N_3222,N_3858);
nand U4579 (N_4579,N_3723,N_3539);
and U4580 (N_4580,N_3162,N_3298);
and U4581 (N_4581,N_3111,N_3703);
and U4582 (N_4582,N_3324,N_3249);
or U4583 (N_4583,N_3547,N_3690);
nand U4584 (N_4584,N_3312,N_3381);
and U4585 (N_4585,N_3409,N_3265);
xnor U4586 (N_4586,N_3527,N_3642);
and U4587 (N_4587,N_3514,N_3960);
nand U4588 (N_4588,N_3685,N_3285);
and U4589 (N_4589,N_3107,N_3063);
and U4590 (N_4590,N_3622,N_3194);
xor U4591 (N_4591,N_3545,N_3288);
xnor U4592 (N_4592,N_3594,N_3685);
and U4593 (N_4593,N_3589,N_3635);
or U4594 (N_4594,N_3664,N_3950);
and U4595 (N_4595,N_3124,N_3780);
nor U4596 (N_4596,N_3796,N_3089);
or U4597 (N_4597,N_3336,N_3720);
or U4598 (N_4598,N_3663,N_3764);
or U4599 (N_4599,N_3477,N_3215);
and U4600 (N_4600,N_3966,N_3237);
or U4601 (N_4601,N_3549,N_3187);
and U4602 (N_4602,N_3636,N_3543);
or U4603 (N_4603,N_3605,N_3900);
nand U4604 (N_4604,N_3193,N_3946);
or U4605 (N_4605,N_3734,N_3398);
nor U4606 (N_4606,N_3159,N_3329);
xor U4607 (N_4607,N_3680,N_3587);
nand U4608 (N_4608,N_3026,N_3204);
xnor U4609 (N_4609,N_3628,N_3209);
or U4610 (N_4610,N_3987,N_3523);
nor U4611 (N_4611,N_3258,N_3398);
or U4612 (N_4612,N_3201,N_3750);
or U4613 (N_4613,N_3462,N_3405);
nor U4614 (N_4614,N_3056,N_3388);
or U4615 (N_4615,N_3802,N_3033);
and U4616 (N_4616,N_3483,N_3789);
nand U4617 (N_4617,N_3945,N_3975);
and U4618 (N_4618,N_3014,N_3101);
nand U4619 (N_4619,N_3550,N_3717);
nor U4620 (N_4620,N_3574,N_3612);
or U4621 (N_4621,N_3110,N_3031);
or U4622 (N_4622,N_3267,N_3845);
or U4623 (N_4623,N_3224,N_3780);
nand U4624 (N_4624,N_3143,N_3575);
nand U4625 (N_4625,N_3926,N_3047);
xnor U4626 (N_4626,N_3837,N_3174);
nand U4627 (N_4627,N_3359,N_3546);
or U4628 (N_4628,N_3524,N_3857);
nand U4629 (N_4629,N_3925,N_3440);
or U4630 (N_4630,N_3834,N_3155);
or U4631 (N_4631,N_3654,N_3135);
and U4632 (N_4632,N_3118,N_3169);
or U4633 (N_4633,N_3804,N_3178);
or U4634 (N_4634,N_3820,N_3845);
or U4635 (N_4635,N_3210,N_3241);
nor U4636 (N_4636,N_3829,N_3303);
nand U4637 (N_4637,N_3046,N_3016);
or U4638 (N_4638,N_3511,N_3908);
or U4639 (N_4639,N_3599,N_3027);
nand U4640 (N_4640,N_3412,N_3947);
nand U4641 (N_4641,N_3301,N_3165);
nor U4642 (N_4642,N_3969,N_3727);
nor U4643 (N_4643,N_3240,N_3859);
or U4644 (N_4644,N_3582,N_3075);
and U4645 (N_4645,N_3643,N_3230);
or U4646 (N_4646,N_3626,N_3161);
nand U4647 (N_4647,N_3821,N_3321);
or U4648 (N_4648,N_3760,N_3636);
and U4649 (N_4649,N_3013,N_3508);
or U4650 (N_4650,N_3068,N_3011);
nor U4651 (N_4651,N_3065,N_3326);
nand U4652 (N_4652,N_3650,N_3627);
nand U4653 (N_4653,N_3865,N_3769);
nand U4654 (N_4654,N_3595,N_3365);
nor U4655 (N_4655,N_3613,N_3774);
nand U4656 (N_4656,N_3839,N_3002);
xor U4657 (N_4657,N_3639,N_3419);
and U4658 (N_4658,N_3324,N_3042);
or U4659 (N_4659,N_3224,N_3500);
nor U4660 (N_4660,N_3395,N_3982);
or U4661 (N_4661,N_3047,N_3691);
nand U4662 (N_4662,N_3104,N_3380);
nor U4663 (N_4663,N_3123,N_3677);
nor U4664 (N_4664,N_3298,N_3044);
nor U4665 (N_4665,N_3995,N_3208);
xnor U4666 (N_4666,N_3447,N_3964);
nor U4667 (N_4667,N_3022,N_3930);
or U4668 (N_4668,N_3079,N_3596);
nand U4669 (N_4669,N_3749,N_3209);
or U4670 (N_4670,N_3380,N_3926);
and U4671 (N_4671,N_3811,N_3075);
and U4672 (N_4672,N_3601,N_3914);
nor U4673 (N_4673,N_3497,N_3810);
or U4674 (N_4674,N_3597,N_3300);
nor U4675 (N_4675,N_3102,N_3756);
nand U4676 (N_4676,N_3080,N_3519);
nor U4677 (N_4677,N_3240,N_3539);
and U4678 (N_4678,N_3922,N_3117);
and U4679 (N_4679,N_3596,N_3223);
nor U4680 (N_4680,N_3672,N_3826);
or U4681 (N_4681,N_3471,N_3682);
nor U4682 (N_4682,N_3015,N_3605);
nor U4683 (N_4683,N_3287,N_3655);
nor U4684 (N_4684,N_3162,N_3270);
xor U4685 (N_4685,N_3521,N_3995);
or U4686 (N_4686,N_3402,N_3048);
and U4687 (N_4687,N_3353,N_3416);
and U4688 (N_4688,N_3890,N_3479);
and U4689 (N_4689,N_3605,N_3725);
nand U4690 (N_4690,N_3670,N_3915);
nor U4691 (N_4691,N_3590,N_3785);
or U4692 (N_4692,N_3451,N_3638);
xor U4693 (N_4693,N_3843,N_3932);
nor U4694 (N_4694,N_3745,N_3274);
or U4695 (N_4695,N_3376,N_3019);
nor U4696 (N_4696,N_3871,N_3057);
nand U4697 (N_4697,N_3444,N_3891);
xor U4698 (N_4698,N_3065,N_3131);
xnor U4699 (N_4699,N_3050,N_3208);
and U4700 (N_4700,N_3932,N_3404);
or U4701 (N_4701,N_3526,N_3727);
and U4702 (N_4702,N_3685,N_3096);
nand U4703 (N_4703,N_3036,N_3195);
nand U4704 (N_4704,N_3261,N_3864);
nor U4705 (N_4705,N_3354,N_3186);
nand U4706 (N_4706,N_3116,N_3229);
and U4707 (N_4707,N_3880,N_3488);
nand U4708 (N_4708,N_3434,N_3695);
nor U4709 (N_4709,N_3715,N_3147);
nand U4710 (N_4710,N_3523,N_3484);
and U4711 (N_4711,N_3614,N_3872);
or U4712 (N_4712,N_3677,N_3027);
or U4713 (N_4713,N_3630,N_3749);
or U4714 (N_4714,N_3201,N_3999);
or U4715 (N_4715,N_3513,N_3532);
and U4716 (N_4716,N_3092,N_3553);
nand U4717 (N_4717,N_3218,N_3112);
xor U4718 (N_4718,N_3102,N_3526);
or U4719 (N_4719,N_3735,N_3701);
nor U4720 (N_4720,N_3105,N_3226);
or U4721 (N_4721,N_3247,N_3402);
nand U4722 (N_4722,N_3515,N_3646);
and U4723 (N_4723,N_3367,N_3360);
nor U4724 (N_4724,N_3413,N_3780);
nand U4725 (N_4725,N_3907,N_3314);
and U4726 (N_4726,N_3104,N_3000);
or U4727 (N_4727,N_3579,N_3408);
nor U4728 (N_4728,N_3039,N_3763);
and U4729 (N_4729,N_3468,N_3618);
nand U4730 (N_4730,N_3314,N_3604);
and U4731 (N_4731,N_3188,N_3246);
xnor U4732 (N_4732,N_3460,N_3227);
and U4733 (N_4733,N_3354,N_3589);
and U4734 (N_4734,N_3845,N_3806);
and U4735 (N_4735,N_3776,N_3537);
and U4736 (N_4736,N_3302,N_3416);
and U4737 (N_4737,N_3819,N_3445);
nand U4738 (N_4738,N_3033,N_3766);
and U4739 (N_4739,N_3797,N_3123);
nand U4740 (N_4740,N_3733,N_3124);
and U4741 (N_4741,N_3826,N_3301);
nand U4742 (N_4742,N_3982,N_3698);
or U4743 (N_4743,N_3590,N_3583);
or U4744 (N_4744,N_3475,N_3123);
nor U4745 (N_4745,N_3435,N_3922);
or U4746 (N_4746,N_3082,N_3515);
nand U4747 (N_4747,N_3151,N_3914);
nand U4748 (N_4748,N_3072,N_3744);
nand U4749 (N_4749,N_3106,N_3461);
or U4750 (N_4750,N_3007,N_3128);
and U4751 (N_4751,N_3179,N_3176);
nor U4752 (N_4752,N_3812,N_3863);
xnor U4753 (N_4753,N_3858,N_3382);
nor U4754 (N_4754,N_3671,N_3910);
and U4755 (N_4755,N_3763,N_3845);
nand U4756 (N_4756,N_3837,N_3520);
or U4757 (N_4757,N_3161,N_3587);
nor U4758 (N_4758,N_3393,N_3660);
nand U4759 (N_4759,N_3073,N_3007);
or U4760 (N_4760,N_3170,N_3520);
nand U4761 (N_4761,N_3804,N_3106);
nand U4762 (N_4762,N_3490,N_3520);
nor U4763 (N_4763,N_3097,N_3844);
nor U4764 (N_4764,N_3592,N_3947);
nor U4765 (N_4765,N_3729,N_3210);
and U4766 (N_4766,N_3402,N_3033);
and U4767 (N_4767,N_3812,N_3707);
or U4768 (N_4768,N_3822,N_3743);
or U4769 (N_4769,N_3209,N_3379);
xor U4770 (N_4770,N_3067,N_3766);
xnor U4771 (N_4771,N_3593,N_3786);
and U4772 (N_4772,N_3089,N_3186);
xor U4773 (N_4773,N_3033,N_3229);
and U4774 (N_4774,N_3483,N_3646);
or U4775 (N_4775,N_3920,N_3165);
and U4776 (N_4776,N_3541,N_3290);
xnor U4777 (N_4777,N_3647,N_3038);
nand U4778 (N_4778,N_3995,N_3285);
and U4779 (N_4779,N_3672,N_3490);
or U4780 (N_4780,N_3253,N_3166);
nor U4781 (N_4781,N_3632,N_3899);
xor U4782 (N_4782,N_3173,N_3082);
nand U4783 (N_4783,N_3238,N_3831);
or U4784 (N_4784,N_3700,N_3259);
or U4785 (N_4785,N_3965,N_3508);
nor U4786 (N_4786,N_3700,N_3097);
nand U4787 (N_4787,N_3174,N_3446);
and U4788 (N_4788,N_3655,N_3181);
or U4789 (N_4789,N_3537,N_3035);
and U4790 (N_4790,N_3910,N_3655);
and U4791 (N_4791,N_3080,N_3702);
and U4792 (N_4792,N_3551,N_3834);
nand U4793 (N_4793,N_3001,N_3170);
nand U4794 (N_4794,N_3857,N_3757);
or U4795 (N_4795,N_3398,N_3131);
or U4796 (N_4796,N_3219,N_3640);
nand U4797 (N_4797,N_3602,N_3056);
nor U4798 (N_4798,N_3288,N_3085);
nor U4799 (N_4799,N_3372,N_3969);
nor U4800 (N_4800,N_3729,N_3129);
xnor U4801 (N_4801,N_3169,N_3491);
nor U4802 (N_4802,N_3710,N_3377);
and U4803 (N_4803,N_3229,N_3925);
nand U4804 (N_4804,N_3139,N_3127);
nor U4805 (N_4805,N_3002,N_3419);
or U4806 (N_4806,N_3264,N_3596);
nand U4807 (N_4807,N_3123,N_3353);
and U4808 (N_4808,N_3617,N_3635);
xor U4809 (N_4809,N_3466,N_3338);
nor U4810 (N_4810,N_3116,N_3106);
nand U4811 (N_4811,N_3963,N_3671);
or U4812 (N_4812,N_3798,N_3116);
xor U4813 (N_4813,N_3430,N_3047);
xnor U4814 (N_4814,N_3679,N_3839);
nor U4815 (N_4815,N_3242,N_3399);
nor U4816 (N_4816,N_3735,N_3475);
and U4817 (N_4817,N_3551,N_3129);
and U4818 (N_4818,N_3849,N_3319);
nor U4819 (N_4819,N_3560,N_3867);
xnor U4820 (N_4820,N_3682,N_3440);
nand U4821 (N_4821,N_3074,N_3372);
nand U4822 (N_4822,N_3752,N_3365);
xor U4823 (N_4823,N_3593,N_3173);
nor U4824 (N_4824,N_3845,N_3839);
or U4825 (N_4825,N_3281,N_3402);
nand U4826 (N_4826,N_3117,N_3369);
nor U4827 (N_4827,N_3518,N_3641);
nand U4828 (N_4828,N_3251,N_3439);
xor U4829 (N_4829,N_3910,N_3337);
or U4830 (N_4830,N_3805,N_3581);
nor U4831 (N_4831,N_3778,N_3807);
and U4832 (N_4832,N_3187,N_3056);
nand U4833 (N_4833,N_3461,N_3112);
nor U4834 (N_4834,N_3785,N_3491);
nor U4835 (N_4835,N_3913,N_3309);
or U4836 (N_4836,N_3822,N_3741);
xor U4837 (N_4837,N_3951,N_3673);
and U4838 (N_4838,N_3708,N_3951);
nand U4839 (N_4839,N_3493,N_3147);
or U4840 (N_4840,N_3461,N_3712);
nand U4841 (N_4841,N_3129,N_3899);
or U4842 (N_4842,N_3439,N_3941);
xor U4843 (N_4843,N_3917,N_3495);
nor U4844 (N_4844,N_3978,N_3278);
nor U4845 (N_4845,N_3612,N_3461);
or U4846 (N_4846,N_3686,N_3297);
nor U4847 (N_4847,N_3695,N_3711);
or U4848 (N_4848,N_3205,N_3609);
nand U4849 (N_4849,N_3936,N_3843);
and U4850 (N_4850,N_3475,N_3085);
and U4851 (N_4851,N_3991,N_3694);
or U4852 (N_4852,N_3754,N_3098);
and U4853 (N_4853,N_3110,N_3483);
nand U4854 (N_4854,N_3065,N_3961);
and U4855 (N_4855,N_3887,N_3414);
and U4856 (N_4856,N_3450,N_3601);
nand U4857 (N_4857,N_3919,N_3554);
nand U4858 (N_4858,N_3413,N_3451);
xnor U4859 (N_4859,N_3838,N_3598);
nand U4860 (N_4860,N_3832,N_3525);
nor U4861 (N_4861,N_3633,N_3137);
and U4862 (N_4862,N_3214,N_3136);
xnor U4863 (N_4863,N_3162,N_3862);
and U4864 (N_4864,N_3604,N_3117);
nand U4865 (N_4865,N_3248,N_3450);
and U4866 (N_4866,N_3116,N_3385);
xor U4867 (N_4867,N_3091,N_3824);
or U4868 (N_4868,N_3097,N_3959);
nor U4869 (N_4869,N_3800,N_3458);
nor U4870 (N_4870,N_3231,N_3793);
nand U4871 (N_4871,N_3379,N_3520);
nand U4872 (N_4872,N_3958,N_3844);
nor U4873 (N_4873,N_3261,N_3047);
nand U4874 (N_4874,N_3183,N_3204);
nor U4875 (N_4875,N_3655,N_3789);
nor U4876 (N_4876,N_3214,N_3668);
or U4877 (N_4877,N_3399,N_3213);
or U4878 (N_4878,N_3359,N_3788);
nor U4879 (N_4879,N_3632,N_3607);
or U4880 (N_4880,N_3183,N_3446);
or U4881 (N_4881,N_3693,N_3458);
or U4882 (N_4882,N_3799,N_3338);
and U4883 (N_4883,N_3193,N_3662);
or U4884 (N_4884,N_3616,N_3488);
or U4885 (N_4885,N_3445,N_3531);
nand U4886 (N_4886,N_3913,N_3458);
nand U4887 (N_4887,N_3572,N_3072);
or U4888 (N_4888,N_3553,N_3540);
or U4889 (N_4889,N_3777,N_3113);
or U4890 (N_4890,N_3335,N_3312);
and U4891 (N_4891,N_3447,N_3909);
and U4892 (N_4892,N_3500,N_3355);
nand U4893 (N_4893,N_3714,N_3389);
and U4894 (N_4894,N_3384,N_3694);
or U4895 (N_4895,N_3320,N_3555);
nand U4896 (N_4896,N_3119,N_3418);
nand U4897 (N_4897,N_3522,N_3512);
or U4898 (N_4898,N_3267,N_3115);
xor U4899 (N_4899,N_3573,N_3427);
nand U4900 (N_4900,N_3436,N_3050);
nor U4901 (N_4901,N_3065,N_3072);
nand U4902 (N_4902,N_3513,N_3767);
or U4903 (N_4903,N_3359,N_3362);
nor U4904 (N_4904,N_3676,N_3540);
xnor U4905 (N_4905,N_3709,N_3887);
nor U4906 (N_4906,N_3228,N_3629);
nand U4907 (N_4907,N_3967,N_3150);
nand U4908 (N_4908,N_3807,N_3122);
nand U4909 (N_4909,N_3140,N_3794);
xnor U4910 (N_4910,N_3467,N_3672);
nand U4911 (N_4911,N_3086,N_3205);
and U4912 (N_4912,N_3549,N_3811);
or U4913 (N_4913,N_3165,N_3222);
and U4914 (N_4914,N_3929,N_3687);
xor U4915 (N_4915,N_3710,N_3663);
nor U4916 (N_4916,N_3067,N_3607);
nor U4917 (N_4917,N_3962,N_3339);
and U4918 (N_4918,N_3930,N_3021);
nor U4919 (N_4919,N_3742,N_3210);
xnor U4920 (N_4920,N_3946,N_3422);
nor U4921 (N_4921,N_3663,N_3960);
nand U4922 (N_4922,N_3259,N_3268);
or U4923 (N_4923,N_3068,N_3570);
nand U4924 (N_4924,N_3806,N_3173);
or U4925 (N_4925,N_3075,N_3057);
nor U4926 (N_4926,N_3569,N_3730);
and U4927 (N_4927,N_3031,N_3047);
xor U4928 (N_4928,N_3527,N_3894);
nand U4929 (N_4929,N_3856,N_3729);
nor U4930 (N_4930,N_3118,N_3874);
nor U4931 (N_4931,N_3689,N_3198);
and U4932 (N_4932,N_3923,N_3822);
nor U4933 (N_4933,N_3093,N_3612);
xnor U4934 (N_4934,N_3929,N_3952);
nor U4935 (N_4935,N_3233,N_3468);
or U4936 (N_4936,N_3407,N_3515);
or U4937 (N_4937,N_3391,N_3968);
and U4938 (N_4938,N_3240,N_3256);
and U4939 (N_4939,N_3231,N_3908);
nor U4940 (N_4940,N_3349,N_3737);
and U4941 (N_4941,N_3580,N_3963);
nand U4942 (N_4942,N_3274,N_3614);
or U4943 (N_4943,N_3475,N_3322);
and U4944 (N_4944,N_3880,N_3866);
or U4945 (N_4945,N_3888,N_3196);
nand U4946 (N_4946,N_3678,N_3361);
nor U4947 (N_4947,N_3117,N_3508);
xor U4948 (N_4948,N_3020,N_3968);
and U4949 (N_4949,N_3835,N_3703);
and U4950 (N_4950,N_3037,N_3863);
nand U4951 (N_4951,N_3766,N_3745);
and U4952 (N_4952,N_3747,N_3825);
and U4953 (N_4953,N_3856,N_3076);
and U4954 (N_4954,N_3632,N_3557);
nand U4955 (N_4955,N_3463,N_3484);
or U4956 (N_4956,N_3871,N_3324);
and U4957 (N_4957,N_3618,N_3404);
nand U4958 (N_4958,N_3105,N_3843);
nor U4959 (N_4959,N_3697,N_3252);
nor U4960 (N_4960,N_3528,N_3141);
and U4961 (N_4961,N_3855,N_3400);
xor U4962 (N_4962,N_3712,N_3725);
and U4963 (N_4963,N_3670,N_3891);
nand U4964 (N_4964,N_3846,N_3597);
xor U4965 (N_4965,N_3921,N_3709);
and U4966 (N_4966,N_3782,N_3187);
nand U4967 (N_4967,N_3505,N_3624);
nand U4968 (N_4968,N_3625,N_3191);
or U4969 (N_4969,N_3019,N_3073);
and U4970 (N_4970,N_3223,N_3710);
nor U4971 (N_4971,N_3576,N_3134);
and U4972 (N_4972,N_3702,N_3650);
nor U4973 (N_4973,N_3458,N_3784);
nor U4974 (N_4974,N_3702,N_3934);
nor U4975 (N_4975,N_3766,N_3076);
or U4976 (N_4976,N_3275,N_3665);
and U4977 (N_4977,N_3729,N_3205);
nor U4978 (N_4978,N_3953,N_3440);
nor U4979 (N_4979,N_3588,N_3999);
nand U4980 (N_4980,N_3758,N_3733);
xor U4981 (N_4981,N_3582,N_3156);
xnor U4982 (N_4982,N_3847,N_3449);
or U4983 (N_4983,N_3864,N_3450);
nand U4984 (N_4984,N_3864,N_3218);
nand U4985 (N_4985,N_3274,N_3372);
nand U4986 (N_4986,N_3356,N_3015);
or U4987 (N_4987,N_3633,N_3357);
xor U4988 (N_4988,N_3950,N_3252);
and U4989 (N_4989,N_3783,N_3577);
nand U4990 (N_4990,N_3583,N_3268);
and U4991 (N_4991,N_3834,N_3352);
or U4992 (N_4992,N_3200,N_3368);
xor U4993 (N_4993,N_3796,N_3665);
and U4994 (N_4994,N_3127,N_3003);
nor U4995 (N_4995,N_3147,N_3433);
nor U4996 (N_4996,N_3024,N_3323);
nand U4997 (N_4997,N_3614,N_3151);
nor U4998 (N_4998,N_3421,N_3090);
nor U4999 (N_4999,N_3689,N_3497);
nor UO_0 (O_0,N_4535,N_4837);
and UO_1 (O_1,N_4435,N_4739);
nor UO_2 (O_2,N_4668,N_4222);
and UO_3 (O_3,N_4450,N_4298);
nor UO_4 (O_4,N_4604,N_4143);
nand UO_5 (O_5,N_4832,N_4314);
and UO_6 (O_6,N_4133,N_4592);
nor UO_7 (O_7,N_4156,N_4264);
nor UO_8 (O_8,N_4577,N_4751);
nand UO_9 (O_9,N_4157,N_4415);
or UO_10 (O_10,N_4140,N_4362);
and UO_11 (O_11,N_4642,N_4371);
xor UO_12 (O_12,N_4386,N_4276);
nor UO_13 (O_13,N_4902,N_4165);
or UO_14 (O_14,N_4137,N_4227);
xor UO_15 (O_15,N_4570,N_4601);
and UO_16 (O_16,N_4652,N_4387);
and UO_17 (O_17,N_4017,N_4062);
nor UO_18 (O_18,N_4922,N_4281);
nor UO_19 (O_19,N_4052,N_4731);
nand UO_20 (O_20,N_4448,N_4468);
and UO_21 (O_21,N_4269,N_4506);
or UO_22 (O_22,N_4743,N_4584);
nand UO_23 (O_23,N_4383,N_4812);
and UO_24 (O_24,N_4877,N_4033);
or UO_25 (O_25,N_4149,N_4633);
xor UO_26 (O_26,N_4925,N_4817);
and UO_27 (O_27,N_4037,N_4354);
or UO_28 (O_28,N_4238,N_4193);
xnor UO_29 (O_29,N_4809,N_4689);
xor UO_30 (O_30,N_4217,N_4792);
or UO_31 (O_31,N_4000,N_4836);
nor UO_32 (O_32,N_4928,N_4657);
nand UO_33 (O_33,N_4016,N_4352);
nand UO_34 (O_34,N_4816,N_4935);
or UO_35 (O_35,N_4180,N_4789);
and UO_36 (O_36,N_4848,N_4983);
or UO_37 (O_37,N_4503,N_4628);
or UO_38 (O_38,N_4097,N_4481);
nand UO_39 (O_39,N_4700,N_4552);
and UO_40 (O_40,N_4838,N_4365);
and UO_41 (O_41,N_4230,N_4718);
nor UO_42 (O_42,N_4463,N_4617);
and UO_43 (O_43,N_4954,N_4969);
nor UO_44 (O_44,N_4754,N_4393);
nand UO_45 (O_45,N_4830,N_4405);
nand UO_46 (O_46,N_4914,N_4522);
or UO_47 (O_47,N_4758,N_4762);
and UO_48 (O_48,N_4317,N_4429);
nand UO_49 (O_49,N_4963,N_4727);
and UO_50 (O_50,N_4786,N_4400);
or UO_51 (O_51,N_4790,N_4443);
nand UO_52 (O_52,N_4857,N_4005);
nand UO_53 (O_53,N_4986,N_4413);
nor UO_54 (O_54,N_4434,N_4795);
nor UO_55 (O_55,N_4760,N_4350);
or UO_56 (O_56,N_4373,N_4224);
nand UO_57 (O_57,N_4253,N_4273);
and UO_58 (O_58,N_4102,N_4814);
nand UO_59 (O_59,N_4810,N_4012);
nand UO_60 (O_60,N_4977,N_4794);
and UO_61 (O_61,N_4082,N_4894);
or UO_62 (O_62,N_4081,N_4305);
xnor UO_63 (O_63,N_4858,N_4882);
nor UO_64 (O_64,N_4579,N_4591);
and UO_65 (O_65,N_4239,N_4993);
nor UO_66 (O_66,N_4099,N_4865);
and UO_67 (O_67,N_4994,N_4874);
and UO_68 (O_68,N_4337,N_4476);
or UO_69 (O_69,N_4009,N_4211);
nor UO_70 (O_70,N_4161,N_4875);
xnor UO_71 (O_71,N_4145,N_4901);
nand UO_72 (O_72,N_4975,N_4849);
or UO_73 (O_73,N_4195,N_4670);
nor UO_74 (O_74,N_4712,N_4755);
and UO_75 (O_75,N_4656,N_4338);
or UO_76 (O_76,N_4333,N_4171);
nor UO_77 (O_77,N_4547,N_4439);
nor UO_78 (O_78,N_4205,N_4997);
nand UO_79 (O_79,N_4961,N_4254);
and UO_80 (O_80,N_4376,N_4461);
or UO_81 (O_81,N_4626,N_4212);
nand UO_82 (O_82,N_4436,N_4864);
and UO_83 (O_83,N_4471,N_4131);
and UO_84 (O_84,N_4866,N_4699);
nor UO_85 (O_85,N_4638,N_4366);
xor UO_86 (O_86,N_4920,N_4950);
nor UO_87 (O_87,N_4136,N_4730);
xnor UO_88 (O_88,N_4843,N_4500);
nor UO_89 (O_89,N_4528,N_4339);
and UO_90 (O_90,N_4181,N_4342);
and UO_91 (O_91,N_4134,N_4976);
nor UO_92 (O_92,N_4530,N_4597);
nand UO_93 (O_93,N_4655,N_4927);
and UO_94 (O_94,N_4207,N_4290);
nand UO_95 (O_95,N_4879,N_4960);
and UO_96 (O_96,N_4662,N_4771);
and UO_97 (O_97,N_4844,N_4475);
or UO_98 (O_98,N_4806,N_4382);
and UO_99 (O_99,N_4752,N_4368);
nand UO_100 (O_100,N_4142,N_4074);
nor UO_101 (O_101,N_4833,N_4458);
nor UO_102 (O_102,N_4018,N_4659);
and UO_103 (O_103,N_4644,N_4129);
or UO_104 (O_104,N_4462,N_4722);
and UO_105 (O_105,N_4115,N_4572);
or UO_106 (O_106,N_4952,N_4198);
or UO_107 (O_107,N_4460,N_4828);
xor UO_108 (O_108,N_4892,N_4681);
nand UO_109 (O_109,N_4456,N_4199);
or UO_110 (O_110,N_4085,N_4958);
nor UO_111 (O_111,N_4507,N_4703);
xor UO_112 (O_112,N_4084,N_4259);
and UO_113 (O_113,N_4293,N_4770);
nand UO_114 (O_114,N_4164,N_4682);
xor UO_115 (O_115,N_4100,N_4043);
nor UO_116 (O_116,N_4155,N_4791);
nand UO_117 (O_117,N_4728,N_4067);
and UO_118 (O_118,N_4302,N_4380);
nor UO_119 (O_119,N_4929,N_4417);
or UO_120 (O_120,N_4072,N_4614);
xnor UO_121 (O_121,N_4459,N_4797);
nand UO_122 (O_122,N_4824,N_4745);
nand UO_123 (O_123,N_4683,N_4721);
and UO_124 (O_124,N_4690,N_4058);
and UO_125 (O_125,N_4003,N_4498);
or UO_126 (O_126,N_4867,N_4559);
or UO_127 (O_127,N_4412,N_4765);
nand UO_128 (O_128,N_4854,N_4815);
and UO_129 (O_129,N_4374,N_4303);
or UO_130 (O_130,N_4004,N_4457);
nor UO_131 (O_131,N_4422,N_4182);
nor UO_132 (O_132,N_4737,N_4971);
and UO_133 (O_133,N_4263,N_4669);
nor UO_134 (O_134,N_4593,N_4916);
nand UO_135 (O_135,N_4206,N_4545);
or UO_136 (O_136,N_4150,N_4379);
or UO_137 (O_137,N_4146,N_4713);
nand UO_138 (O_138,N_4138,N_4911);
and UO_139 (O_139,N_4203,N_4846);
nor UO_140 (O_140,N_4079,N_4649);
nand UO_141 (O_141,N_4361,N_4953);
xor UO_142 (O_142,N_4951,N_4433);
nand UO_143 (O_143,N_4031,N_4035);
nor UO_144 (O_144,N_4757,N_4391);
or UO_145 (O_145,N_4736,N_4675);
or UO_146 (O_146,N_4325,N_4359);
nor UO_147 (O_147,N_4635,N_4860);
and UO_148 (O_148,N_4621,N_4111);
nor UO_149 (O_149,N_4453,N_4201);
and UO_150 (O_150,N_4266,N_4309);
nor UO_151 (O_151,N_4640,N_4539);
or UO_152 (O_152,N_4784,N_4119);
nand UO_153 (O_153,N_4349,N_4389);
nand UO_154 (O_154,N_4820,N_4039);
nand UO_155 (O_155,N_4533,N_4015);
xnor UO_156 (O_156,N_4934,N_4607);
nor UO_157 (O_157,N_4265,N_4568);
and UO_158 (O_158,N_4447,N_4327);
and UO_159 (O_159,N_4974,N_4377);
and UO_160 (O_160,N_4945,N_4851);
or UO_161 (O_161,N_4488,N_4036);
nand UO_162 (O_162,N_4020,N_4711);
and UO_163 (O_163,N_4873,N_4247);
nor UO_164 (O_164,N_4536,N_4442);
and UO_165 (O_165,N_4550,N_4701);
xor UO_166 (O_166,N_4622,N_4554);
nand UO_167 (O_167,N_4397,N_4586);
nand UO_168 (O_168,N_4895,N_4250);
and UO_169 (O_169,N_4204,N_4286);
xnor UO_170 (O_170,N_4884,N_4924);
nand UO_171 (O_171,N_4335,N_4808);
xor UO_172 (O_172,N_4772,N_4834);
and UO_173 (O_173,N_4048,N_4496);
xnor UO_174 (O_174,N_4982,N_4685);
nor UO_175 (O_175,N_4517,N_4667);
nand UO_176 (O_176,N_4556,N_4278);
nor UO_177 (O_177,N_4847,N_4919);
nor UO_178 (O_178,N_4546,N_4418);
nor UO_179 (O_179,N_4540,N_4190);
and UO_180 (O_180,N_4819,N_4676);
or UO_181 (O_181,N_4571,N_4872);
or UO_182 (O_182,N_4542,N_4581);
nor UO_183 (O_183,N_4600,N_4179);
or UO_184 (O_184,N_4272,N_4406);
nand UO_185 (O_185,N_4779,N_4232);
or UO_186 (O_186,N_4103,N_4316);
and UO_187 (O_187,N_4811,N_4262);
and UO_188 (O_188,N_4355,N_4705);
nand UO_189 (O_189,N_4852,N_4825);
xnor UO_190 (O_190,N_4501,N_4147);
nor UO_191 (O_191,N_4735,N_4534);
and UO_192 (O_192,N_4774,N_4257);
nand UO_193 (O_193,N_4274,N_4077);
or UO_194 (O_194,N_4941,N_4886);
xor UO_195 (O_195,N_4891,N_4491);
nand UO_196 (O_196,N_4162,N_4023);
nand UO_197 (O_197,N_4548,N_4256);
xnor UO_198 (O_198,N_4831,N_4300);
and UO_199 (O_199,N_4484,N_4242);
or UO_200 (O_200,N_4856,N_4385);
nor UO_201 (O_201,N_4279,N_4594);
and UO_202 (O_202,N_4378,N_4096);
or UO_203 (O_203,N_4510,N_4673);
nand UO_204 (O_204,N_4589,N_4940);
or UO_205 (O_205,N_4798,N_4564);
xnor UO_206 (O_206,N_4707,N_4987);
xnor UO_207 (O_207,N_4562,N_4513);
nor UO_208 (O_208,N_4060,N_4189);
nand UO_209 (O_209,N_4040,N_4126);
nand UO_210 (O_210,N_4208,N_4170);
nor UO_211 (O_211,N_4154,N_4942);
nor UO_212 (O_212,N_4807,N_4729);
or UO_213 (O_213,N_4610,N_4973);
or UO_214 (O_214,N_4527,N_4066);
or UO_215 (O_215,N_4346,N_4076);
nor UO_216 (O_216,N_4748,N_4110);
and UO_217 (O_217,N_4215,N_4645);
nand UO_218 (O_218,N_4679,N_4416);
xor UO_219 (O_219,N_4905,N_4663);
nand UO_220 (O_220,N_4078,N_4859);
and UO_221 (O_221,N_4850,N_4432);
nor UO_222 (O_222,N_4933,N_4135);
nor UO_223 (O_223,N_4245,N_4310);
nand UO_224 (O_224,N_4744,N_4411);
and UO_225 (O_225,N_4213,N_4915);
nor UO_226 (O_226,N_4069,N_4647);
nor UO_227 (O_227,N_4661,N_4778);
xnor UO_228 (O_228,N_4616,N_4014);
nor UO_229 (O_229,N_4602,N_4151);
and UO_230 (O_230,N_4909,N_4306);
or UO_231 (O_231,N_4061,N_4561);
xor UO_232 (O_232,N_4184,N_4297);
or UO_233 (O_233,N_4390,N_4392);
nand UO_234 (O_234,N_4674,N_4172);
nor UO_235 (O_235,N_4629,N_4876);
nor UO_236 (O_236,N_4719,N_4341);
or UO_237 (O_237,N_4292,N_4419);
nor UO_238 (O_238,N_4426,N_4637);
nor UO_239 (O_239,N_4324,N_4803);
nor UO_240 (O_240,N_4261,N_4258);
nor UO_241 (O_241,N_4399,N_4908);
and UO_242 (O_242,N_4381,N_4989);
nand UO_243 (O_243,N_4630,N_4428);
and UO_244 (O_244,N_4050,N_4835);
nand UO_245 (O_245,N_4479,N_4243);
or UO_246 (O_246,N_4367,N_4560);
and UO_247 (O_247,N_4868,N_4421);
and UO_248 (O_248,N_4880,N_4401);
and UO_249 (O_249,N_4687,N_4704);
xor UO_250 (O_250,N_4631,N_4906);
xnor UO_251 (O_251,N_4431,N_4214);
nand UO_252 (O_252,N_4191,N_4108);
nor UO_253 (O_253,N_4148,N_4294);
and UO_254 (O_254,N_4492,N_4351);
nand UO_255 (O_255,N_4715,N_4627);
or UO_256 (O_256,N_4862,N_4032);
xor UO_257 (O_257,N_4968,N_4101);
nand UO_258 (O_258,N_4904,N_4684);
or UO_259 (O_259,N_4839,N_4277);
nor UO_260 (O_260,N_4080,N_4139);
and UO_261 (O_261,N_4364,N_4311);
and UO_262 (O_262,N_4781,N_4956);
and UO_263 (O_263,N_4223,N_4802);
nor UO_264 (O_264,N_4537,N_4175);
or UO_265 (O_265,N_4580,N_4287);
and UO_266 (O_266,N_4123,N_4329);
nand UO_267 (O_267,N_4252,N_4246);
nand UO_268 (O_268,N_4529,N_4965);
and UO_269 (O_269,N_4955,N_4499);
nor UO_270 (O_270,N_4469,N_4502);
or UO_271 (O_271,N_4709,N_4551);
nand UO_272 (O_272,N_4793,N_4444);
and UO_273 (O_273,N_4888,N_4130);
or UO_274 (O_274,N_4724,N_4677);
and UO_275 (O_275,N_4008,N_4696);
nor UO_276 (O_276,N_4410,N_4787);
nor UO_277 (O_277,N_4296,N_4932);
and UO_278 (O_278,N_4898,N_4420);
nand UO_279 (O_279,N_4026,N_4720);
and UO_280 (O_280,N_4717,N_4508);
nor UO_281 (O_281,N_4240,N_4966);
or UO_282 (O_282,N_4512,N_4714);
xnor UO_283 (O_283,N_4768,N_4219);
and UO_284 (O_284,N_4588,N_4896);
nor UO_285 (O_285,N_4693,N_4192);
nand UO_286 (O_286,N_4596,N_4235);
or UO_287 (O_287,N_4912,N_4907);
and UO_288 (O_288,N_4007,N_4144);
nor UO_289 (O_289,N_4978,N_4634);
nand UO_290 (O_290,N_4054,N_4396);
or UO_291 (O_291,N_4599,N_4363);
nand UO_292 (O_292,N_4315,N_4438);
nand UO_293 (O_293,N_4334,N_4318);
or UO_294 (O_294,N_4782,N_4002);
nand UO_295 (O_295,N_4231,N_4805);
nand UO_296 (O_296,N_4641,N_4489);
nand UO_297 (O_297,N_4511,N_4086);
nand UO_298 (O_298,N_4326,N_4585);
nor UO_299 (O_299,N_4943,N_4913);
nor UO_300 (O_300,N_4590,N_4611);
nand UO_301 (O_301,N_4283,N_4509);
and UO_302 (O_302,N_4959,N_4988);
or UO_303 (O_303,N_4163,N_4057);
nand UO_304 (O_304,N_4910,N_4578);
nor UO_305 (O_305,N_4490,N_4995);
nor UO_306 (O_306,N_4716,N_4042);
or UO_307 (O_307,N_4372,N_4021);
nand UO_308 (O_308,N_4220,N_4090);
nor UO_309 (O_309,N_4408,N_4524);
and UO_310 (O_310,N_4046,N_4347);
or UO_311 (O_311,N_4775,N_4783);
nor UO_312 (O_312,N_4799,N_4188);
or UO_313 (O_313,N_4092,N_4024);
nand UO_314 (O_314,N_4288,N_4889);
or UO_315 (O_315,N_4939,N_4019);
or UO_316 (O_316,N_4075,N_4531);
nor UO_317 (O_317,N_4885,N_4826);
nand UO_318 (O_318,N_4555,N_4653);
or UO_319 (O_319,N_4344,N_4345);
and UO_320 (O_320,N_4395,N_4726);
or UO_321 (O_321,N_4255,N_4981);
nand UO_322 (O_322,N_4313,N_4064);
nand UO_323 (O_323,N_4407,N_4625);
nor UO_324 (O_324,N_4823,N_4112);
nand UO_325 (O_325,N_4451,N_4068);
or UO_326 (O_326,N_4998,N_4900);
or UO_327 (O_327,N_4893,N_4121);
or UO_328 (O_328,N_4738,N_4369);
nand UO_329 (O_329,N_4249,N_4595);
and UO_330 (O_330,N_4917,N_4473);
nand UO_331 (O_331,N_4105,N_4178);
or UO_332 (O_332,N_4109,N_4404);
or UO_333 (O_333,N_4241,N_4741);
xor UO_334 (O_334,N_4152,N_4120);
and UO_335 (O_335,N_4887,N_4788);
nor UO_336 (O_336,N_4226,N_4780);
and UO_337 (O_337,N_4284,N_4514);
xor UO_338 (O_338,N_4660,N_4526);
or UO_339 (O_339,N_4495,N_4937);
nand UO_340 (O_340,N_4938,N_4763);
nand UO_341 (O_341,N_4665,N_4518);
and UO_342 (O_342,N_4127,N_4466);
nand UO_343 (O_343,N_4425,N_4169);
nor UO_344 (O_344,N_4010,N_4210);
or UO_345 (O_345,N_4800,N_4025);
nor UO_346 (O_346,N_4636,N_4285);
and UO_347 (O_347,N_4767,N_4801);
nor UO_348 (O_348,N_4878,N_4861);
or UO_349 (O_349,N_4776,N_4761);
nor UO_350 (O_350,N_4478,N_4984);
xor UO_351 (O_351,N_4044,N_4691);
nand UO_352 (O_352,N_4903,N_4117);
nor UO_353 (O_353,N_4944,N_4173);
and UO_354 (O_354,N_4863,N_4702);
nor UO_355 (O_355,N_4615,N_4268);
nor UO_356 (O_356,N_4710,N_4124);
nand UO_357 (O_357,N_4946,N_4999);
nand UO_358 (O_358,N_4356,N_4557);
nand UO_359 (O_359,N_4624,N_4218);
and UO_360 (O_360,N_4605,N_4482);
xnor UO_361 (O_361,N_4360,N_4308);
nand UO_362 (O_362,N_4609,N_4962);
nand UO_363 (O_363,N_4125,N_4582);
or UO_364 (O_364,N_4107,N_4918);
nor UO_365 (O_365,N_4104,N_4516);
nand UO_366 (O_366,N_4643,N_4197);
or UO_367 (O_367,N_4304,N_4094);
nor UO_368 (O_368,N_4985,N_4957);
nor UO_369 (O_369,N_4132,N_4445);
and UO_370 (O_370,N_4764,N_4299);
nand UO_371 (O_371,N_4260,N_4098);
and UO_372 (O_372,N_4370,N_4295);
nor UO_373 (O_373,N_4723,N_4688);
nor UO_374 (O_374,N_4055,N_4027);
nor UO_375 (O_375,N_4821,N_4883);
nand UO_376 (O_376,N_4307,N_4523);
or UO_377 (O_377,N_4237,N_4011);
and UO_378 (O_378,N_4549,N_4678);
nor UO_379 (O_379,N_4174,N_4612);
xnor UO_380 (O_380,N_4095,N_4398);
nand UO_381 (O_381,N_4493,N_4613);
or UO_382 (O_382,N_4343,N_4071);
or UO_383 (O_383,N_4452,N_4186);
nand UO_384 (O_384,N_4931,N_4056);
nand UO_385 (O_385,N_4271,N_4244);
and UO_386 (O_386,N_4477,N_4646);
nor UO_387 (O_387,N_4006,N_4598);
and UO_388 (O_388,N_4870,N_4454);
nor UO_389 (O_389,N_4167,N_4070);
nand UO_390 (O_390,N_4725,N_4756);
nor UO_391 (O_391,N_4441,N_4202);
and UO_392 (O_392,N_4521,N_4996);
or UO_393 (O_393,N_4708,N_4472);
nor UO_394 (O_394,N_4449,N_4541);
or UO_395 (O_395,N_4323,N_4575);
and UO_396 (O_396,N_4566,N_4427);
nand UO_397 (O_397,N_4990,N_4567);
xnor UO_398 (O_398,N_4773,N_4948);
xnor UO_399 (O_399,N_4038,N_4234);
and UO_400 (O_400,N_4087,N_4291);
xor UO_401 (O_401,N_4553,N_4648);
or UO_402 (O_402,N_4280,N_4194);
nand UO_403 (O_403,N_4289,N_4047);
xor UO_404 (O_404,N_4979,N_4248);
nand UO_405 (O_405,N_4651,N_4409);
and UO_406 (O_406,N_4028,N_4930);
and UO_407 (O_407,N_4113,N_4620);
nand UO_408 (O_408,N_4251,N_4606);
or UO_409 (O_409,N_4632,N_4936);
nand UO_410 (O_410,N_4753,N_4497);
nor UO_411 (O_411,N_4991,N_4470);
and UO_412 (O_412,N_4947,N_4766);
nor UO_413 (O_413,N_4001,N_4200);
or UO_414 (O_414,N_4970,N_4746);
or UO_415 (O_415,N_4437,N_4742);
xnor UO_416 (O_416,N_4225,N_4650);
or UO_417 (O_417,N_4827,N_4654);
nand UO_418 (O_418,N_4336,N_4855);
or UO_419 (O_419,N_4576,N_4890);
and UO_420 (O_420,N_4623,N_4465);
nor UO_421 (O_421,N_4394,N_4270);
nand UO_422 (O_422,N_4357,N_4899);
nor UO_423 (O_423,N_4680,N_4992);
xnor UO_424 (O_424,N_4525,N_4089);
and UO_425 (O_425,N_4051,N_4664);
nor UO_426 (O_426,N_4740,N_4221);
nand UO_427 (O_427,N_4332,N_4563);
xnor UO_428 (O_428,N_4515,N_4053);
or UO_429 (O_429,N_4686,N_4176);
nand UO_430 (O_430,N_4538,N_4750);
nor UO_431 (O_431,N_4840,N_4759);
or UO_432 (O_432,N_4639,N_4695);
and UO_433 (O_433,N_4116,N_4822);
nor UO_434 (O_434,N_4073,N_4574);
nand UO_435 (O_435,N_4348,N_4697);
and UO_436 (O_436,N_4059,N_4177);
and UO_437 (O_437,N_4088,N_4532);
nand UO_438 (O_438,N_4328,N_4233);
or UO_439 (O_439,N_4504,N_4565);
and UO_440 (O_440,N_4423,N_4330);
nand UO_441 (O_441,N_4187,N_4569);
xnor UO_442 (O_442,N_4083,N_4467);
and UO_443 (O_443,N_4505,N_4480);
or UO_444 (O_444,N_4049,N_4732);
or UO_445 (O_445,N_4464,N_4777);
or UO_446 (O_446,N_4749,N_4353);
or UO_447 (O_447,N_4029,N_4694);
nor UO_448 (O_448,N_4446,N_4603);
xor UO_449 (O_449,N_4159,N_4091);
nand UO_450 (O_450,N_4440,N_4331);
or UO_451 (O_451,N_4402,N_4388);
or UO_452 (O_452,N_4671,N_4964);
nand UO_453 (O_453,N_4698,N_4034);
xnor UO_454 (O_454,N_4319,N_4871);
xnor UO_455 (O_455,N_4706,N_4375);
xor UO_456 (O_456,N_4168,N_4485);
and UO_457 (O_457,N_4487,N_4845);
nor UO_458 (O_458,N_4796,N_4322);
xor UO_459 (O_459,N_4185,N_4747);
or UO_460 (O_460,N_4128,N_4692);
xor UO_461 (O_461,N_4818,N_4430);
or UO_462 (O_462,N_4923,N_4065);
nand UO_463 (O_463,N_4573,N_4587);
and UO_464 (O_464,N_4926,N_4804);
xor UO_465 (O_465,N_4813,N_4734);
or UO_466 (O_466,N_4869,N_4106);
nand UO_467 (O_467,N_4114,N_4340);
and UO_468 (O_468,N_4520,N_4897);
nand UO_469 (O_469,N_4196,N_4483);
nor UO_470 (O_470,N_4045,N_4141);
and UO_471 (O_471,N_4785,N_4041);
and UO_472 (O_472,N_4320,N_4030);
and UO_473 (O_473,N_4312,N_4013);
or UO_474 (O_474,N_4158,N_4209);
nand UO_475 (O_475,N_4921,N_4967);
nor UO_476 (O_476,N_4829,N_4881);
nand UO_477 (O_477,N_4558,N_4486);
nand UO_478 (O_478,N_4544,N_4658);
nor UO_479 (O_479,N_4267,N_4769);
and UO_480 (O_480,N_4583,N_4853);
nor UO_481 (O_481,N_4321,N_4842);
and UO_482 (O_482,N_4733,N_4122);
nand UO_483 (O_483,N_4160,N_4358);
xnor UO_484 (O_484,N_4474,N_4424);
nor UO_485 (O_485,N_4414,N_4153);
xor UO_486 (O_486,N_4841,N_4980);
nor UO_487 (O_487,N_4949,N_4455);
nor UO_488 (O_488,N_4229,N_4618);
nand UO_489 (O_489,N_4543,N_4403);
and UO_490 (O_490,N_4118,N_4519);
nand UO_491 (O_491,N_4236,N_4166);
nor UO_492 (O_492,N_4022,N_4619);
nor UO_493 (O_493,N_4228,N_4282);
and UO_494 (O_494,N_4216,N_4384);
or UO_495 (O_495,N_4275,N_4666);
and UO_496 (O_496,N_4093,N_4301);
nor UO_497 (O_497,N_4672,N_4608);
nor UO_498 (O_498,N_4494,N_4972);
nand UO_499 (O_499,N_4183,N_4063);
and UO_500 (O_500,N_4763,N_4382);
xor UO_501 (O_501,N_4023,N_4628);
nor UO_502 (O_502,N_4798,N_4072);
and UO_503 (O_503,N_4795,N_4447);
or UO_504 (O_504,N_4878,N_4124);
nand UO_505 (O_505,N_4347,N_4894);
nand UO_506 (O_506,N_4195,N_4201);
and UO_507 (O_507,N_4542,N_4349);
and UO_508 (O_508,N_4428,N_4444);
nor UO_509 (O_509,N_4374,N_4751);
nand UO_510 (O_510,N_4590,N_4303);
or UO_511 (O_511,N_4645,N_4667);
and UO_512 (O_512,N_4424,N_4127);
or UO_513 (O_513,N_4708,N_4638);
and UO_514 (O_514,N_4792,N_4074);
xnor UO_515 (O_515,N_4332,N_4810);
and UO_516 (O_516,N_4695,N_4552);
nor UO_517 (O_517,N_4818,N_4857);
nand UO_518 (O_518,N_4149,N_4860);
and UO_519 (O_519,N_4413,N_4115);
nand UO_520 (O_520,N_4387,N_4982);
or UO_521 (O_521,N_4466,N_4776);
or UO_522 (O_522,N_4900,N_4099);
and UO_523 (O_523,N_4889,N_4366);
nand UO_524 (O_524,N_4398,N_4330);
or UO_525 (O_525,N_4107,N_4616);
and UO_526 (O_526,N_4965,N_4302);
or UO_527 (O_527,N_4913,N_4290);
or UO_528 (O_528,N_4224,N_4394);
nand UO_529 (O_529,N_4706,N_4494);
nand UO_530 (O_530,N_4271,N_4055);
xnor UO_531 (O_531,N_4372,N_4863);
nand UO_532 (O_532,N_4376,N_4507);
or UO_533 (O_533,N_4578,N_4418);
and UO_534 (O_534,N_4159,N_4213);
and UO_535 (O_535,N_4993,N_4588);
and UO_536 (O_536,N_4950,N_4902);
nor UO_537 (O_537,N_4935,N_4308);
or UO_538 (O_538,N_4362,N_4480);
xor UO_539 (O_539,N_4960,N_4961);
and UO_540 (O_540,N_4090,N_4558);
xor UO_541 (O_541,N_4778,N_4928);
or UO_542 (O_542,N_4776,N_4889);
nand UO_543 (O_543,N_4220,N_4538);
nand UO_544 (O_544,N_4785,N_4331);
nand UO_545 (O_545,N_4869,N_4804);
xor UO_546 (O_546,N_4428,N_4237);
nand UO_547 (O_547,N_4013,N_4188);
and UO_548 (O_548,N_4837,N_4257);
nand UO_549 (O_549,N_4372,N_4549);
nor UO_550 (O_550,N_4986,N_4889);
nand UO_551 (O_551,N_4030,N_4137);
or UO_552 (O_552,N_4366,N_4729);
nand UO_553 (O_553,N_4426,N_4503);
or UO_554 (O_554,N_4907,N_4751);
and UO_555 (O_555,N_4885,N_4511);
or UO_556 (O_556,N_4750,N_4272);
or UO_557 (O_557,N_4997,N_4481);
or UO_558 (O_558,N_4843,N_4817);
or UO_559 (O_559,N_4672,N_4118);
and UO_560 (O_560,N_4455,N_4467);
and UO_561 (O_561,N_4637,N_4173);
and UO_562 (O_562,N_4576,N_4959);
nor UO_563 (O_563,N_4098,N_4208);
xor UO_564 (O_564,N_4125,N_4602);
nand UO_565 (O_565,N_4372,N_4952);
and UO_566 (O_566,N_4987,N_4547);
nor UO_567 (O_567,N_4763,N_4080);
nand UO_568 (O_568,N_4873,N_4817);
nor UO_569 (O_569,N_4912,N_4401);
or UO_570 (O_570,N_4729,N_4099);
nand UO_571 (O_571,N_4760,N_4953);
and UO_572 (O_572,N_4330,N_4345);
nand UO_573 (O_573,N_4579,N_4055);
and UO_574 (O_574,N_4707,N_4435);
and UO_575 (O_575,N_4365,N_4720);
or UO_576 (O_576,N_4189,N_4917);
nor UO_577 (O_577,N_4724,N_4818);
nand UO_578 (O_578,N_4226,N_4867);
xnor UO_579 (O_579,N_4220,N_4016);
nor UO_580 (O_580,N_4724,N_4419);
or UO_581 (O_581,N_4982,N_4313);
nor UO_582 (O_582,N_4424,N_4282);
and UO_583 (O_583,N_4357,N_4666);
or UO_584 (O_584,N_4863,N_4586);
and UO_585 (O_585,N_4316,N_4256);
or UO_586 (O_586,N_4760,N_4473);
or UO_587 (O_587,N_4482,N_4151);
nor UO_588 (O_588,N_4815,N_4951);
xor UO_589 (O_589,N_4460,N_4711);
nand UO_590 (O_590,N_4029,N_4119);
nor UO_591 (O_591,N_4191,N_4681);
nor UO_592 (O_592,N_4061,N_4281);
or UO_593 (O_593,N_4728,N_4089);
nor UO_594 (O_594,N_4182,N_4662);
and UO_595 (O_595,N_4789,N_4772);
nand UO_596 (O_596,N_4261,N_4167);
nor UO_597 (O_597,N_4070,N_4571);
and UO_598 (O_598,N_4181,N_4842);
xnor UO_599 (O_599,N_4435,N_4928);
and UO_600 (O_600,N_4474,N_4653);
and UO_601 (O_601,N_4322,N_4389);
and UO_602 (O_602,N_4685,N_4431);
nor UO_603 (O_603,N_4651,N_4082);
nor UO_604 (O_604,N_4123,N_4110);
or UO_605 (O_605,N_4195,N_4514);
nand UO_606 (O_606,N_4887,N_4496);
or UO_607 (O_607,N_4865,N_4498);
nand UO_608 (O_608,N_4499,N_4131);
nor UO_609 (O_609,N_4584,N_4583);
nor UO_610 (O_610,N_4122,N_4842);
nor UO_611 (O_611,N_4742,N_4258);
and UO_612 (O_612,N_4982,N_4281);
or UO_613 (O_613,N_4195,N_4556);
xor UO_614 (O_614,N_4440,N_4475);
and UO_615 (O_615,N_4956,N_4851);
nor UO_616 (O_616,N_4212,N_4902);
nor UO_617 (O_617,N_4974,N_4492);
or UO_618 (O_618,N_4679,N_4382);
nor UO_619 (O_619,N_4429,N_4790);
and UO_620 (O_620,N_4703,N_4353);
xnor UO_621 (O_621,N_4493,N_4523);
and UO_622 (O_622,N_4188,N_4479);
nor UO_623 (O_623,N_4030,N_4144);
nor UO_624 (O_624,N_4822,N_4189);
nand UO_625 (O_625,N_4263,N_4872);
nand UO_626 (O_626,N_4432,N_4001);
nor UO_627 (O_627,N_4614,N_4659);
or UO_628 (O_628,N_4607,N_4701);
and UO_629 (O_629,N_4590,N_4197);
or UO_630 (O_630,N_4250,N_4840);
or UO_631 (O_631,N_4515,N_4662);
and UO_632 (O_632,N_4610,N_4734);
nor UO_633 (O_633,N_4042,N_4639);
and UO_634 (O_634,N_4848,N_4642);
nor UO_635 (O_635,N_4001,N_4540);
or UO_636 (O_636,N_4617,N_4014);
and UO_637 (O_637,N_4171,N_4115);
nand UO_638 (O_638,N_4377,N_4887);
and UO_639 (O_639,N_4070,N_4099);
and UO_640 (O_640,N_4957,N_4851);
or UO_641 (O_641,N_4302,N_4768);
nand UO_642 (O_642,N_4887,N_4078);
and UO_643 (O_643,N_4060,N_4590);
nor UO_644 (O_644,N_4227,N_4952);
and UO_645 (O_645,N_4061,N_4830);
or UO_646 (O_646,N_4517,N_4189);
nor UO_647 (O_647,N_4631,N_4048);
or UO_648 (O_648,N_4936,N_4907);
or UO_649 (O_649,N_4507,N_4326);
xnor UO_650 (O_650,N_4823,N_4029);
and UO_651 (O_651,N_4855,N_4806);
xnor UO_652 (O_652,N_4064,N_4540);
and UO_653 (O_653,N_4501,N_4567);
and UO_654 (O_654,N_4206,N_4833);
nor UO_655 (O_655,N_4472,N_4895);
and UO_656 (O_656,N_4373,N_4082);
and UO_657 (O_657,N_4365,N_4579);
or UO_658 (O_658,N_4076,N_4503);
nor UO_659 (O_659,N_4905,N_4287);
or UO_660 (O_660,N_4201,N_4006);
and UO_661 (O_661,N_4103,N_4783);
nand UO_662 (O_662,N_4408,N_4261);
xor UO_663 (O_663,N_4571,N_4238);
and UO_664 (O_664,N_4124,N_4572);
and UO_665 (O_665,N_4006,N_4541);
nor UO_666 (O_666,N_4621,N_4568);
and UO_667 (O_667,N_4411,N_4200);
and UO_668 (O_668,N_4977,N_4391);
or UO_669 (O_669,N_4853,N_4719);
xor UO_670 (O_670,N_4830,N_4614);
nor UO_671 (O_671,N_4930,N_4669);
and UO_672 (O_672,N_4928,N_4023);
xor UO_673 (O_673,N_4231,N_4485);
nor UO_674 (O_674,N_4886,N_4351);
or UO_675 (O_675,N_4476,N_4900);
xor UO_676 (O_676,N_4835,N_4193);
nor UO_677 (O_677,N_4722,N_4908);
nand UO_678 (O_678,N_4320,N_4746);
nor UO_679 (O_679,N_4148,N_4223);
and UO_680 (O_680,N_4111,N_4728);
nand UO_681 (O_681,N_4920,N_4012);
and UO_682 (O_682,N_4746,N_4070);
nand UO_683 (O_683,N_4372,N_4743);
and UO_684 (O_684,N_4534,N_4459);
nand UO_685 (O_685,N_4234,N_4855);
or UO_686 (O_686,N_4781,N_4817);
or UO_687 (O_687,N_4078,N_4446);
xor UO_688 (O_688,N_4879,N_4340);
nor UO_689 (O_689,N_4204,N_4445);
and UO_690 (O_690,N_4649,N_4298);
nor UO_691 (O_691,N_4699,N_4638);
and UO_692 (O_692,N_4497,N_4032);
and UO_693 (O_693,N_4231,N_4342);
nor UO_694 (O_694,N_4340,N_4145);
or UO_695 (O_695,N_4209,N_4422);
nand UO_696 (O_696,N_4239,N_4084);
and UO_697 (O_697,N_4905,N_4102);
and UO_698 (O_698,N_4980,N_4995);
or UO_699 (O_699,N_4043,N_4264);
nor UO_700 (O_700,N_4026,N_4574);
or UO_701 (O_701,N_4229,N_4377);
xnor UO_702 (O_702,N_4051,N_4009);
nor UO_703 (O_703,N_4020,N_4905);
or UO_704 (O_704,N_4208,N_4152);
and UO_705 (O_705,N_4530,N_4242);
or UO_706 (O_706,N_4275,N_4929);
nand UO_707 (O_707,N_4080,N_4688);
nand UO_708 (O_708,N_4902,N_4725);
nor UO_709 (O_709,N_4102,N_4460);
or UO_710 (O_710,N_4839,N_4128);
nor UO_711 (O_711,N_4386,N_4086);
nand UO_712 (O_712,N_4175,N_4187);
nand UO_713 (O_713,N_4952,N_4569);
xnor UO_714 (O_714,N_4988,N_4806);
or UO_715 (O_715,N_4873,N_4851);
and UO_716 (O_716,N_4200,N_4906);
nand UO_717 (O_717,N_4195,N_4555);
and UO_718 (O_718,N_4000,N_4182);
nand UO_719 (O_719,N_4861,N_4276);
xnor UO_720 (O_720,N_4684,N_4536);
nor UO_721 (O_721,N_4751,N_4334);
or UO_722 (O_722,N_4063,N_4004);
nand UO_723 (O_723,N_4941,N_4502);
nor UO_724 (O_724,N_4195,N_4681);
nor UO_725 (O_725,N_4947,N_4399);
nor UO_726 (O_726,N_4674,N_4454);
or UO_727 (O_727,N_4895,N_4727);
and UO_728 (O_728,N_4204,N_4627);
nand UO_729 (O_729,N_4862,N_4904);
nor UO_730 (O_730,N_4530,N_4598);
nor UO_731 (O_731,N_4794,N_4168);
nand UO_732 (O_732,N_4490,N_4541);
nor UO_733 (O_733,N_4217,N_4710);
or UO_734 (O_734,N_4431,N_4312);
nor UO_735 (O_735,N_4721,N_4566);
or UO_736 (O_736,N_4796,N_4286);
nand UO_737 (O_737,N_4031,N_4474);
nand UO_738 (O_738,N_4594,N_4040);
or UO_739 (O_739,N_4388,N_4103);
xor UO_740 (O_740,N_4611,N_4356);
xnor UO_741 (O_741,N_4105,N_4638);
nor UO_742 (O_742,N_4026,N_4603);
nor UO_743 (O_743,N_4206,N_4356);
or UO_744 (O_744,N_4089,N_4397);
nor UO_745 (O_745,N_4377,N_4531);
or UO_746 (O_746,N_4967,N_4140);
nor UO_747 (O_747,N_4053,N_4163);
nor UO_748 (O_748,N_4656,N_4973);
nand UO_749 (O_749,N_4327,N_4948);
and UO_750 (O_750,N_4998,N_4626);
nor UO_751 (O_751,N_4716,N_4199);
nand UO_752 (O_752,N_4539,N_4962);
nand UO_753 (O_753,N_4107,N_4931);
nand UO_754 (O_754,N_4888,N_4283);
and UO_755 (O_755,N_4523,N_4023);
nand UO_756 (O_756,N_4009,N_4586);
nand UO_757 (O_757,N_4753,N_4849);
nand UO_758 (O_758,N_4848,N_4784);
nor UO_759 (O_759,N_4558,N_4948);
or UO_760 (O_760,N_4595,N_4615);
or UO_761 (O_761,N_4322,N_4449);
nand UO_762 (O_762,N_4775,N_4406);
or UO_763 (O_763,N_4262,N_4638);
nor UO_764 (O_764,N_4349,N_4321);
nand UO_765 (O_765,N_4102,N_4477);
and UO_766 (O_766,N_4331,N_4563);
or UO_767 (O_767,N_4046,N_4374);
and UO_768 (O_768,N_4179,N_4056);
or UO_769 (O_769,N_4826,N_4271);
nor UO_770 (O_770,N_4872,N_4568);
nor UO_771 (O_771,N_4390,N_4818);
and UO_772 (O_772,N_4746,N_4774);
or UO_773 (O_773,N_4160,N_4708);
nand UO_774 (O_774,N_4993,N_4972);
xnor UO_775 (O_775,N_4450,N_4946);
nand UO_776 (O_776,N_4432,N_4887);
nand UO_777 (O_777,N_4112,N_4787);
or UO_778 (O_778,N_4485,N_4584);
nor UO_779 (O_779,N_4833,N_4992);
nor UO_780 (O_780,N_4636,N_4161);
nand UO_781 (O_781,N_4617,N_4942);
nand UO_782 (O_782,N_4804,N_4148);
or UO_783 (O_783,N_4485,N_4011);
nor UO_784 (O_784,N_4105,N_4108);
or UO_785 (O_785,N_4505,N_4174);
nor UO_786 (O_786,N_4301,N_4903);
and UO_787 (O_787,N_4307,N_4304);
or UO_788 (O_788,N_4956,N_4223);
nand UO_789 (O_789,N_4884,N_4210);
xor UO_790 (O_790,N_4140,N_4207);
and UO_791 (O_791,N_4358,N_4038);
nor UO_792 (O_792,N_4715,N_4685);
xnor UO_793 (O_793,N_4935,N_4771);
or UO_794 (O_794,N_4387,N_4226);
nand UO_795 (O_795,N_4079,N_4351);
or UO_796 (O_796,N_4334,N_4416);
nand UO_797 (O_797,N_4478,N_4329);
or UO_798 (O_798,N_4276,N_4555);
or UO_799 (O_799,N_4550,N_4624);
or UO_800 (O_800,N_4271,N_4779);
nand UO_801 (O_801,N_4534,N_4288);
xnor UO_802 (O_802,N_4631,N_4061);
nand UO_803 (O_803,N_4108,N_4783);
nor UO_804 (O_804,N_4680,N_4049);
nor UO_805 (O_805,N_4069,N_4036);
xor UO_806 (O_806,N_4706,N_4893);
nor UO_807 (O_807,N_4887,N_4216);
and UO_808 (O_808,N_4992,N_4884);
nand UO_809 (O_809,N_4975,N_4363);
xor UO_810 (O_810,N_4241,N_4583);
or UO_811 (O_811,N_4215,N_4197);
and UO_812 (O_812,N_4282,N_4895);
nand UO_813 (O_813,N_4738,N_4043);
nand UO_814 (O_814,N_4796,N_4478);
nor UO_815 (O_815,N_4973,N_4861);
nand UO_816 (O_816,N_4196,N_4110);
or UO_817 (O_817,N_4708,N_4930);
xor UO_818 (O_818,N_4350,N_4542);
or UO_819 (O_819,N_4061,N_4958);
or UO_820 (O_820,N_4898,N_4201);
xnor UO_821 (O_821,N_4516,N_4695);
or UO_822 (O_822,N_4948,N_4374);
nand UO_823 (O_823,N_4066,N_4458);
or UO_824 (O_824,N_4997,N_4306);
nor UO_825 (O_825,N_4547,N_4252);
or UO_826 (O_826,N_4086,N_4969);
and UO_827 (O_827,N_4479,N_4780);
nand UO_828 (O_828,N_4359,N_4703);
nor UO_829 (O_829,N_4507,N_4355);
or UO_830 (O_830,N_4214,N_4511);
nor UO_831 (O_831,N_4053,N_4613);
nor UO_832 (O_832,N_4397,N_4504);
nor UO_833 (O_833,N_4226,N_4613);
or UO_834 (O_834,N_4249,N_4641);
and UO_835 (O_835,N_4272,N_4734);
and UO_836 (O_836,N_4369,N_4291);
nand UO_837 (O_837,N_4458,N_4632);
nor UO_838 (O_838,N_4115,N_4103);
or UO_839 (O_839,N_4036,N_4110);
nand UO_840 (O_840,N_4813,N_4134);
nor UO_841 (O_841,N_4415,N_4120);
nand UO_842 (O_842,N_4510,N_4154);
and UO_843 (O_843,N_4761,N_4136);
or UO_844 (O_844,N_4880,N_4652);
nand UO_845 (O_845,N_4164,N_4034);
and UO_846 (O_846,N_4708,N_4647);
and UO_847 (O_847,N_4200,N_4431);
and UO_848 (O_848,N_4662,N_4464);
nand UO_849 (O_849,N_4587,N_4266);
nor UO_850 (O_850,N_4356,N_4208);
nor UO_851 (O_851,N_4311,N_4368);
xor UO_852 (O_852,N_4987,N_4316);
or UO_853 (O_853,N_4606,N_4905);
nand UO_854 (O_854,N_4274,N_4170);
xnor UO_855 (O_855,N_4654,N_4971);
and UO_856 (O_856,N_4156,N_4714);
nor UO_857 (O_857,N_4433,N_4561);
nand UO_858 (O_858,N_4508,N_4654);
and UO_859 (O_859,N_4582,N_4045);
nand UO_860 (O_860,N_4822,N_4368);
and UO_861 (O_861,N_4848,N_4063);
or UO_862 (O_862,N_4046,N_4898);
or UO_863 (O_863,N_4903,N_4767);
and UO_864 (O_864,N_4958,N_4516);
and UO_865 (O_865,N_4774,N_4023);
and UO_866 (O_866,N_4166,N_4249);
nand UO_867 (O_867,N_4124,N_4371);
xnor UO_868 (O_868,N_4481,N_4131);
nor UO_869 (O_869,N_4934,N_4688);
nand UO_870 (O_870,N_4451,N_4565);
or UO_871 (O_871,N_4372,N_4165);
and UO_872 (O_872,N_4311,N_4825);
and UO_873 (O_873,N_4987,N_4552);
nand UO_874 (O_874,N_4908,N_4755);
and UO_875 (O_875,N_4710,N_4521);
and UO_876 (O_876,N_4973,N_4277);
and UO_877 (O_877,N_4158,N_4983);
xnor UO_878 (O_878,N_4719,N_4582);
nor UO_879 (O_879,N_4338,N_4296);
or UO_880 (O_880,N_4418,N_4018);
nand UO_881 (O_881,N_4105,N_4771);
xor UO_882 (O_882,N_4972,N_4943);
nor UO_883 (O_883,N_4414,N_4042);
nor UO_884 (O_884,N_4197,N_4688);
nor UO_885 (O_885,N_4346,N_4936);
xor UO_886 (O_886,N_4248,N_4582);
nor UO_887 (O_887,N_4201,N_4582);
or UO_888 (O_888,N_4348,N_4973);
or UO_889 (O_889,N_4596,N_4716);
and UO_890 (O_890,N_4886,N_4464);
nand UO_891 (O_891,N_4071,N_4187);
nor UO_892 (O_892,N_4156,N_4786);
xor UO_893 (O_893,N_4448,N_4556);
xor UO_894 (O_894,N_4583,N_4312);
or UO_895 (O_895,N_4031,N_4667);
nor UO_896 (O_896,N_4886,N_4219);
xor UO_897 (O_897,N_4862,N_4445);
or UO_898 (O_898,N_4584,N_4852);
nor UO_899 (O_899,N_4674,N_4893);
nor UO_900 (O_900,N_4660,N_4518);
nand UO_901 (O_901,N_4587,N_4690);
and UO_902 (O_902,N_4075,N_4295);
nand UO_903 (O_903,N_4026,N_4964);
or UO_904 (O_904,N_4964,N_4177);
xor UO_905 (O_905,N_4716,N_4715);
nand UO_906 (O_906,N_4088,N_4869);
and UO_907 (O_907,N_4066,N_4983);
or UO_908 (O_908,N_4778,N_4386);
nand UO_909 (O_909,N_4342,N_4053);
and UO_910 (O_910,N_4237,N_4564);
xnor UO_911 (O_911,N_4418,N_4159);
nand UO_912 (O_912,N_4256,N_4822);
or UO_913 (O_913,N_4170,N_4118);
xor UO_914 (O_914,N_4615,N_4105);
and UO_915 (O_915,N_4609,N_4700);
nor UO_916 (O_916,N_4114,N_4153);
nor UO_917 (O_917,N_4366,N_4416);
and UO_918 (O_918,N_4787,N_4327);
nand UO_919 (O_919,N_4191,N_4464);
nand UO_920 (O_920,N_4582,N_4615);
or UO_921 (O_921,N_4839,N_4391);
nand UO_922 (O_922,N_4562,N_4738);
nor UO_923 (O_923,N_4233,N_4589);
and UO_924 (O_924,N_4831,N_4426);
nand UO_925 (O_925,N_4111,N_4818);
and UO_926 (O_926,N_4957,N_4767);
nand UO_927 (O_927,N_4465,N_4337);
or UO_928 (O_928,N_4908,N_4329);
or UO_929 (O_929,N_4605,N_4538);
nand UO_930 (O_930,N_4121,N_4804);
or UO_931 (O_931,N_4157,N_4706);
nand UO_932 (O_932,N_4750,N_4869);
nand UO_933 (O_933,N_4757,N_4286);
nand UO_934 (O_934,N_4614,N_4068);
nand UO_935 (O_935,N_4437,N_4099);
and UO_936 (O_936,N_4235,N_4940);
and UO_937 (O_937,N_4737,N_4791);
and UO_938 (O_938,N_4242,N_4832);
or UO_939 (O_939,N_4604,N_4566);
nand UO_940 (O_940,N_4818,N_4886);
xnor UO_941 (O_941,N_4595,N_4063);
and UO_942 (O_942,N_4560,N_4549);
and UO_943 (O_943,N_4338,N_4351);
nor UO_944 (O_944,N_4859,N_4545);
or UO_945 (O_945,N_4124,N_4046);
or UO_946 (O_946,N_4287,N_4982);
nor UO_947 (O_947,N_4604,N_4193);
or UO_948 (O_948,N_4369,N_4284);
nor UO_949 (O_949,N_4143,N_4102);
or UO_950 (O_950,N_4850,N_4098);
nor UO_951 (O_951,N_4953,N_4541);
and UO_952 (O_952,N_4132,N_4591);
xnor UO_953 (O_953,N_4015,N_4381);
xnor UO_954 (O_954,N_4118,N_4504);
or UO_955 (O_955,N_4712,N_4699);
or UO_956 (O_956,N_4891,N_4751);
or UO_957 (O_957,N_4709,N_4688);
or UO_958 (O_958,N_4237,N_4665);
nand UO_959 (O_959,N_4895,N_4949);
or UO_960 (O_960,N_4989,N_4574);
nand UO_961 (O_961,N_4239,N_4162);
or UO_962 (O_962,N_4727,N_4571);
nor UO_963 (O_963,N_4874,N_4989);
nand UO_964 (O_964,N_4105,N_4534);
nand UO_965 (O_965,N_4757,N_4773);
or UO_966 (O_966,N_4195,N_4718);
nand UO_967 (O_967,N_4656,N_4876);
xor UO_968 (O_968,N_4541,N_4472);
or UO_969 (O_969,N_4043,N_4581);
and UO_970 (O_970,N_4898,N_4308);
or UO_971 (O_971,N_4043,N_4106);
or UO_972 (O_972,N_4903,N_4680);
and UO_973 (O_973,N_4239,N_4096);
and UO_974 (O_974,N_4914,N_4148);
nand UO_975 (O_975,N_4185,N_4555);
and UO_976 (O_976,N_4726,N_4468);
nand UO_977 (O_977,N_4718,N_4781);
or UO_978 (O_978,N_4992,N_4539);
nor UO_979 (O_979,N_4537,N_4723);
or UO_980 (O_980,N_4282,N_4301);
and UO_981 (O_981,N_4873,N_4156);
xor UO_982 (O_982,N_4759,N_4825);
nand UO_983 (O_983,N_4168,N_4891);
nor UO_984 (O_984,N_4894,N_4258);
and UO_985 (O_985,N_4536,N_4941);
or UO_986 (O_986,N_4012,N_4891);
or UO_987 (O_987,N_4600,N_4623);
nand UO_988 (O_988,N_4607,N_4150);
nand UO_989 (O_989,N_4643,N_4494);
and UO_990 (O_990,N_4990,N_4295);
and UO_991 (O_991,N_4806,N_4542);
and UO_992 (O_992,N_4427,N_4313);
nor UO_993 (O_993,N_4581,N_4558);
or UO_994 (O_994,N_4034,N_4358);
and UO_995 (O_995,N_4183,N_4454);
and UO_996 (O_996,N_4728,N_4413);
or UO_997 (O_997,N_4130,N_4590);
and UO_998 (O_998,N_4093,N_4653);
or UO_999 (O_999,N_4230,N_4484);
endmodule