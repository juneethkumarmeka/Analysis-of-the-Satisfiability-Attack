module basic_750_5000_1000_10_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_166,In_424);
or U1 (N_1,In_388,In_581);
and U2 (N_2,In_216,In_685);
nor U3 (N_3,In_105,In_680);
nor U4 (N_4,In_236,In_360);
nand U5 (N_5,In_645,In_138);
nand U6 (N_6,In_295,In_268);
nor U7 (N_7,In_541,In_239);
xor U8 (N_8,In_475,In_395);
or U9 (N_9,In_525,In_662);
xnor U10 (N_10,In_492,In_255);
or U11 (N_11,In_269,In_337);
or U12 (N_12,In_693,In_387);
nor U13 (N_13,In_65,In_543);
or U14 (N_14,In_554,In_526);
or U15 (N_15,In_565,In_77);
xnor U16 (N_16,In_35,In_466);
nand U17 (N_17,In_98,In_636);
nor U18 (N_18,In_155,In_21);
or U19 (N_19,In_352,In_444);
nand U20 (N_20,In_384,In_39);
or U21 (N_21,In_451,In_81);
or U22 (N_22,In_745,In_373);
nand U23 (N_23,In_506,In_717);
nor U24 (N_24,In_383,In_176);
and U25 (N_25,In_464,In_487);
nor U26 (N_26,In_127,In_143);
nor U27 (N_27,In_686,In_282);
xor U28 (N_28,In_440,In_202);
nor U29 (N_29,In_528,In_746);
nor U30 (N_30,In_0,In_28);
and U31 (N_31,In_262,In_347);
nor U32 (N_32,In_296,In_692);
or U33 (N_33,In_483,In_720);
and U34 (N_34,In_86,In_722);
or U35 (N_35,In_307,In_469);
nand U36 (N_36,In_731,In_635);
nor U37 (N_37,In_69,In_736);
nand U38 (N_38,In_364,In_376);
and U39 (N_39,In_343,In_418);
or U40 (N_40,In_442,In_749);
nand U41 (N_41,In_718,In_672);
nor U42 (N_42,In_460,In_571);
and U43 (N_43,In_50,In_289);
nor U44 (N_44,In_169,In_73);
or U45 (N_45,In_597,In_198);
nand U46 (N_46,In_321,In_305);
nand U47 (N_47,In_192,In_697);
and U48 (N_48,In_682,In_485);
or U49 (N_49,In_38,In_304);
nor U50 (N_50,In_429,In_389);
nor U51 (N_51,In_471,In_664);
and U52 (N_52,In_29,In_181);
and U53 (N_53,In_103,In_154);
or U54 (N_54,In_27,In_342);
nand U55 (N_55,In_194,In_445);
nand U56 (N_56,In_625,In_533);
nand U57 (N_57,In_443,In_125);
or U58 (N_58,In_520,In_41);
and U59 (N_59,In_354,In_548);
and U60 (N_60,In_341,In_264);
xor U61 (N_61,In_71,In_546);
nand U62 (N_62,In_441,In_674);
or U63 (N_63,In_57,In_617);
and U64 (N_64,In_695,In_159);
xnor U65 (N_65,In_472,In_94);
and U66 (N_66,In_286,In_719);
or U67 (N_67,In_509,In_284);
or U68 (N_68,In_299,In_660);
nor U69 (N_69,In_704,In_164);
nor U70 (N_70,In_335,In_333);
or U71 (N_71,In_739,In_233);
xnor U72 (N_72,In_40,In_80);
and U73 (N_73,In_409,In_477);
and U74 (N_74,In_728,In_14);
or U75 (N_75,In_663,In_539);
and U76 (N_76,In_671,In_238);
xnor U77 (N_77,In_129,In_147);
xor U78 (N_78,In_721,In_36);
nand U79 (N_79,In_223,In_687);
nor U80 (N_80,In_288,In_427);
and U81 (N_81,In_495,In_186);
or U82 (N_82,In_455,In_742);
xnor U83 (N_83,In_173,In_730);
nand U84 (N_84,In_535,In_684);
nor U85 (N_85,In_627,In_47);
and U86 (N_86,In_414,In_690);
or U87 (N_87,In_560,In_74);
and U88 (N_88,In_263,In_331);
and U89 (N_89,In_568,In_380);
nor U90 (N_90,In_408,In_608);
xnor U91 (N_91,In_346,In_698);
nor U92 (N_92,In_142,In_538);
and U93 (N_93,In_213,In_24);
and U94 (N_94,In_274,In_378);
nor U95 (N_95,In_273,In_97);
xnor U96 (N_96,In_6,In_430);
or U97 (N_97,In_700,In_590);
xor U98 (N_98,In_523,In_167);
nand U99 (N_99,In_531,In_639);
nand U100 (N_100,In_334,In_200);
or U101 (N_101,In_20,In_115);
or U102 (N_102,In_740,In_620);
xor U103 (N_103,In_610,In_163);
and U104 (N_104,In_175,In_92);
nor U105 (N_105,In_479,In_615);
and U106 (N_106,In_577,In_641);
nand U107 (N_107,In_706,In_275);
nor U108 (N_108,In_206,In_209);
xor U109 (N_109,In_715,In_658);
or U110 (N_110,In_398,In_667);
nor U111 (N_111,In_432,In_569);
nor U112 (N_112,In_132,In_505);
and U113 (N_113,In_504,In_499);
xnor U114 (N_114,In_43,In_478);
nand U115 (N_115,In_95,In_183);
and U116 (N_116,In_621,In_292);
xnor U117 (N_117,In_688,In_19);
and U118 (N_118,In_324,In_253);
nand U119 (N_119,In_247,In_707);
xnor U120 (N_120,In_351,In_270);
or U121 (N_121,In_184,In_600);
and U122 (N_122,In_592,In_566);
or U123 (N_123,In_649,In_177);
and U124 (N_124,In_725,In_422);
and U125 (N_125,In_659,In_574);
or U126 (N_126,In_521,In_594);
nand U127 (N_127,In_653,In_117);
xnor U128 (N_128,In_677,In_748);
or U129 (N_129,In_189,In_630);
xnor U130 (N_130,In_399,In_67);
nor U131 (N_131,In_205,In_503);
or U132 (N_132,In_542,In_433);
and U133 (N_133,In_151,In_15);
or U134 (N_134,In_493,In_290);
and U135 (N_135,In_723,In_26);
nand U136 (N_136,In_355,In_496);
nand U137 (N_137,In_573,In_410);
xor U138 (N_138,In_515,In_371);
nor U139 (N_139,In_579,In_328);
xnor U140 (N_140,In_283,In_586);
xor U141 (N_141,In_702,In_243);
and U142 (N_142,In_224,In_204);
and U143 (N_143,In_137,In_570);
or U144 (N_144,In_744,In_327);
nor U145 (N_145,In_381,In_517);
xnor U146 (N_146,In_114,In_456);
or U147 (N_147,In_439,In_589);
xnor U148 (N_148,In_168,In_416);
and U149 (N_149,In_710,In_102);
xnor U150 (N_150,In_195,In_88);
xnor U151 (N_151,In_591,In_231);
and U152 (N_152,In_593,In_368);
nor U153 (N_153,In_193,In_647);
nand U154 (N_154,In_618,In_544);
and U155 (N_155,In_747,In_447);
nand U156 (N_156,In_488,In_406);
xor U157 (N_157,In_90,In_258);
nand U158 (N_158,In_512,In_446);
nor U159 (N_159,In_507,In_82);
nand U160 (N_160,In_85,In_55);
nor U161 (N_161,In_259,In_345);
nand U162 (N_162,In_582,In_500);
or U163 (N_163,In_732,In_153);
and U164 (N_164,In_735,In_482);
xor U165 (N_165,In_614,In_470);
nor U166 (N_166,In_476,In_452);
and U167 (N_167,In_121,In_363);
xor U168 (N_168,In_453,In_673);
nand U169 (N_169,In_87,In_437);
and U170 (N_170,In_126,In_108);
or U171 (N_171,In_413,In_415);
xor U172 (N_172,In_237,In_724);
xor U173 (N_173,In_37,In_370);
nor U174 (N_174,In_514,In_448);
xor U175 (N_175,In_598,In_584);
nor U176 (N_176,In_489,In_332);
and U177 (N_177,In_457,In_72);
nor U178 (N_178,In_361,In_134);
and U179 (N_179,In_522,In_42);
and U180 (N_180,In_675,In_314);
nand U181 (N_181,In_423,In_652);
and U182 (N_182,In_218,In_481);
or U183 (N_183,In_711,In_320);
xnor U184 (N_184,In_254,In_315);
nand U185 (N_185,In_642,In_267);
nand U186 (N_186,In_135,In_330);
or U187 (N_187,In_136,In_665);
nor U188 (N_188,In_465,In_683);
nor U189 (N_189,In_729,In_609);
and U190 (N_190,In_63,In_16);
nand U191 (N_191,In_449,In_587);
nor U192 (N_192,In_54,In_172);
and U193 (N_193,In_245,In_34);
nand U194 (N_194,In_30,In_377);
or U195 (N_195,In_393,In_511);
nor U196 (N_196,In_553,In_124);
or U197 (N_197,In_285,In_123);
and U198 (N_198,In_300,In_712);
nor U199 (N_199,In_188,In_336);
or U200 (N_200,In_668,In_165);
nor U201 (N_201,In_228,In_644);
and U202 (N_202,In_353,In_508);
nand U203 (N_203,In_180,In_524);
and U204 (N_204,In_329,In_657);
or U205 (N_205,In_310,In_709);
and U206 (N_206,In_556,In_149);
and U207 (N_207,In_66,In_601);
xnor U208 (N_208,In_100,In_128);
and U209 (N_209,In_434,In_234);
or U210 (N_210,In_89,In_348);
xnor U211 (N_211,In_250,In_713);
nand U212 (N_212,In_616,In_294);
or U213 (N_213,In_25,In_741);
nor U214 (N_214,In_530,In_191);
or U215 (N_215,In_669,In_411);
or U216 (N_216,In_559,In_139);
nand U217 (N_217,In_44,In_372);
xnor U218 (N_218,In_144,In_461);
nor U219 (N_219,In_575,In_557);
xnor U220 (N_220,In_612,In_394);
xnor U221 (N_221,In_678,In_58);
or U222 (N_222,In_547,In_705);
xor U223 (N_223,In_431,In_280);
nor U224 (N_224,In_648,In_112);
and U225 (N_225,In_157,In_580);
and U226 (N_226,In_109,In_497);
or U227 (N_227,In_146,In_291);
and U228 (N_228,In_359,In_46);
and U229 (N_229,In_111,In_96);
and U230 (N_230,In_11,In_532);
xnor U231 (N_231,In_306,In_595);
or U232 (N_232,In_484,In_362);
or U233 (N_233,In_252,In_634);
nand U234 (N_234,In_651,In_61);
nand U235 (N_235,In_1,In_502);
nor U236 (N_236,In_474,In_459);
xor U237 (N_237,In_170,In_156);
and U238 (N_238,In_32,In_537);
nand U239 (N_239,In_162,In_199);
and U240 (N_240,In_344,In_501);
xor U241 (N_241,In_585,In_679);
nand U242 (N_242,In_249,In_179);
xor U243 (N_243,In_490,In_605);
and U244 (N_244,In_450,In_402);
nor U245 (N_245,In_628,In_726);
nand U246 (N_246,In_576,In_552);
nand U247 (N_247,In_436,In_208);
or U248 (N_248,In_369,In_318);
nor U249 (N_249,In_303,In_257);
nor U250 (N_250,In_604,In_83);
and U251 (N_251,In_221,In_248);
nor U252 (N_252,In_438,In_242);
xnor U253 (N_253,In_53,In_646);
nor U254 (N_254,In_222,In_558);
nand U255 (N_255,In_549,In_311);
or U256 (N_256,In_737,In_386);
xor U257 (N_257,In_681,In_9);
xor U258 (N_258,In_670,In_76);
xor U259 (N_259,In_240,In_494);
nand U260 (N_260,In_174,In_317);
and U261 (N_261,In_666,In_110);
and U262 (N_262,In_64,In_229);
and U263 (N_263,In_420,In_407);
nand U264 (N_264,In_227,In_419);
nand U265 (N_265,In_272,In_271);
nor U266 (N_266,In_349,In_301);
nand U267 (N_267,In_458,In_550);
nand U268 (N_268,In_251,In_101);
nor U269 (N_269,In_405,In_603);
nor U270 (N_270,In_160,In_417);
or U271 (N_271,In_7,In_703);
nand U272 (N_272,In_210,In_122);
and U273 (N_273,In_365,In_308);
xnor U274 (N_274,In_59,In_93);
nand U275 (N_275,In_326,In_340);
xnor U276 (N_276,In_319,In_623);
xor U277 (N_277,In_276,In_150);
xor U278 (N_278,In_435,In_701);
or U279 (N_279,In_567,In_397);
xor U280 (N_280,In_131,In_226);
nor U281 (N_281,In_211,In_12);
and U282 (N_282,In_691,In_8);
or U283 (N_283,In_31,In_588);
xnor U284 (N_284,In_385,In_694);
nand U285 (N_285,In_3,In_350);
and U286 (N_286,In_187,In_197);
nor U287 (N_287,In_622,In_426);
nor U288 (N_288,In_5,In_611);
nor U289 (N_289,In_13,In_467);
or U290 (N_290,In_178,In_281);
and U291 (N_291,In_79,In_104);
and U292 (N_292,In_637,In_734);
or U293 (N_293,In_358,In_33);
and U294 (N_294,In_141,In_486);
or U295 (N_295,In_562,In_75);
xor U296 (N_296,In_638,In_322);
xnor U297 (N_297,In_716,In_140);
nand U298 (N_298,In_390,In_106);
nand U299 (N_299,In_599,In_545);
nor U300 (N_300,In_52,In_357);
xor U301 (N_301,In_17,In_561);
or U302 (N_302,In_220,In_325);
and U303 (N_303,In_309,In_374);
nor U304 (N_304,In_624,In_632);
nand U305 (N_305,In_412,In_727);
and U306 (N_306,In_171,In_696);
nor U307 (N_307,In_219,In_404);
xor U308 (N_308,In_714,In_656);
xor U309 (N_309,In_743,In_244);
nor U310 (N_310,In_116,In_68);
xnor U311 (N_311,In_607,In_2);
nand U312 (N_312,In_99,In_463);
nor U313 (N_313,In_62,In_392);
xnor U314 (N_314,In_48,In_733);
nor U315 (N_315,In_602,In_51);
nor U316 (N_316,In_230,In_78);
xor U317 (N_317,In_454,In_215);
xor U318 (N_318,In_260,In_400);
xnor U319 (N_319,In_339,In_689);
and U320 (N_320,In_107,In_613);
nor U321 (N_321,In_473,In_148);
xnor U322 (N_322,In_516,In_241);
or U323 (N_323,In_676,In_498);
or U324 (N_324,In_375,In_428);
nand U325 (N_325,In_396,In_382);
or U326 (N_326,In_91,In_118);
and U327 (N_327,In_572,In_555);
nor U328 (N_328,In_661,In_391);
and U329 (N_329,In_643,In_619);
and U330 (N_330,In_297,In_261);
xor U331 (N_331,In_133,In_425);
nand U332 (N_332,In_212,In_232);
or U333 (N_333,In_185,In_738);
nand U334 (N_334,In_563,In_640);
xnor U335 (N_335,In_654,In_519);
nor U336 (N_336,In_246,In_190);
xor U337 (N_337,In_84,In_534);
nor U338 (N_338,In_564,In_338);
xor U339 (N_339,In_23,In_145);
or U340 (N_340,In_480,In_699);
nand U341 (N_341,In_462,In_596);
xnor U342 (N_342,In_278,In_203);
nor U343 (N_343,In_529,In_302);
nor U344 (N_344,In_22,In_152);
or U345 (N_345,In_421,In_120);
or U346 (N_346,In_45,In_225);
nand U347 (N_347,In_277,In_161);
xnor U348 (N_348,In_287,In_626);
nor U349 (N_349,In_629,In_323);
nor U350 (N_350,In_56,In_113);
nand U351 (N_351,In_119,In_214);
nor U352 (N_352,In_583,In_366);
and U353 (N_353,In_403,In_293);
nand U354 (N_354,In_708,In_578);
nor U355 (N_355,In_49,In_631);
or U356 (N_356,In_158,In_316);
or U357 (N_357,In_207,In_367);
or U358 (N_358,In_379,In_401);
or U359 (N_359,In_4,In_655);
and U360 (N_360,In_551,In_201);
or U361 (N_361,In_60,In_18);
xnor U362 (N_362,In_513,In_256);
nand U363 (N_363,In_536,In_312);
nand U364 (N_364,In_265,In_313);
nand U365 (N_365,In_633,In_10);
and U366 (N_366,In_182,In_650);
or U367 (N_367,In_217,In_356);
or U368 (N_368,In_266,In_491);
or U369 (N_369,In_540,In_468);
or U370 (N_370,In_70,In_196);
or U371 (N_371,In_279,In_527);
xnor U372 (N_372,In_518,In_298);
or U373 (N_373,In_130,In_606);
and U374 (N_374,In_235,In_510);
nor U375 (N_375,In_507,In_678);
and U376 (N_376,In_375,In_40);
nor U377 (N_377,In_594,In_600);
nor U378 (N_378,In_177,In_630);
nand U379 (N_379,In_175,In_394);
and U380 (N_380,In_446,In_270);
nand U381 (N_381,In_439,In_67);
or U382 (N_382,In_372,In_391);
and U383 (N_383,In_243,In_413);
nor U384 (N_384,In_367,In_555);
nor U385 (N_385,In_644,In_219);
xnor U386 (N_386,In_193,In_649);
nand U387 (N_387,In_242,In_268);
nor U388 (N_388,In_541,In_248);
nand U389 (N_389,In_200,In_10);
and U390 (N_390,In_220,In_138);
nand U391 (N_391,In_723,In_193);
xnor U392 (N_392,In_525,In_533);
nor U393 (N_393,In_419,In_718);
xor U394 (N_394,In_400,In_250);
and U395 (N_395,In_486,In_389);
or U396 (N_396,In_48,In_642);
nand U397 (N_397,In_614,In_704);
xor U398 (N_398,In_420,In_455);
nor U399 (N_399,In_512,In_341);
xnor U400 (N_400,In_259,In_539);
nor U401 (N_401,In_434,In_402);
nor U402 (N_402,In_321,In_181);
xnor U403 (N_403,In_512,In_483);
and U404 (N_404,In_283,In_417);
and U405 (N_405,In_678,In_607);
and U406 (N_406,In_307,In_654);
nor U407 (N_407,In_194,In_665);
nor U408 (N_408,In_495,In_360);
and U409 (N_409,In_726,In_511);
xnor U410 (N_410,In_228,In_264);
xor U411 (N_411,In_513,In_509);
and U412 (N_412,In_249,In_98);
xor U413 (N_413,In_143,In_595);
or U414 (N_414,In_4,In_381);
and U415 (N_415,In_139,In_436);
xor U416 (N_416,In_467,In_217);
and U417 (N_417,In_56,In_202);
xor U418 (N_418,In_545,In_353);
nand U419 (N_419,In_500,In_261);
or U420 (N_420,In_724,In_625);
or U421 (N_421,In_47,In_243);
xor U422 (N_422,In_244,In_193);
or U423 (N_423,In_566,In_672);
or U424 (N_424,In_525,In_260);
nor U425 (N_425,In_745,In_296);
and U426 (N_426,In_73,In_40);
nor U427 (N_427,In_20,In_178);
nand U428 (N_428,In_265,In_7);
or U429 (N_429,In_54,In_100);
and U430 (N_430,In_544,In_26);
nor U431 (N_431,In_91,In_322);
and U432 (N_432,In_309,In_23);
or U433 (N_433,In_653,In_132);
xor U434 (N_434,In_637,In_274);
and U435 (N_435,In_201,In_507);
xor U436 (N_436,In_288,In_421);
or U437 (N_437,In_500,In_43);
nor U438 (N_438,In_200,In_719);
nand U439 (N_439,In_443,In_676);
xnor U440 (N_440,In_96,In_533);
or U441 (N_441,In_558,In_478);
xor U442 (N_442,In_372,In_739);
or U443 (N_443,In_97,In_10);
nand U444 (N_444,In_13,In_142);
and U445 (N_445,In_51,In_202);
xor U446 (N_446,In_129,In_438);
or U447 (N_447,In_74,In_214);
nand U448 (N_448,In_748,In_7);
xnor U449 (N_449,In_27,In_537);
and U450 (N_450,In_249,In_554);
nor U451 (N_451,In_342,In_473);
and U452 (N_452,In_83,In_166);
or U453 (N_453,In_142,In_629);
nor U454 (N_454,In_107,In_685);
nand U455 (N_455,In_367,In_480);
nand U456 (N_456,In_11,In_629);
xor U457 (N_457,In_206,In_20);
xor U458 (N_458,In_554,In_577);
nand U459 (N_459,In_551,In_96);
and U460 (N_460,In_306,In_123);
or U461 (N_461,In_609,In_306);
and U462 (N_462,In_42,In_464);
nor U463 (N_463,In_27,In_4);
nor U464 (N_464,In_277,In_335);
and U465 (N_465,In_410,In_143);
nand U466 (N_466,In_49,In_471);
or U467 (N_467,In_352,In_540);
or U468 (N_468,In_470,In_248);
xnor U469 (N_469,In_153,In_606);
nor U470 (N_470,In_605,In_179);
nor U471 (N_471,In_647,In_29);
nor U472 (N_472,In_155,In_120);
nand U473 (N_473,In_213,In_216);
xor U474 (N_474,In_632,In_542);
xor U475 (N_475,In_344,In_361);
nor U476 (N_476,In_688,In_599);
and U477 (N_477,In_282,In_267);
nand U478 (N_478,In_733,In_116);
nand U479 (N_479,In_532,In_407);
nand U480 (N_480,In_21,In_138);
nand U481 (N_481,In_415,In_500);
or U482 (N_482,In_725,In_714);
and U483 (N_483,In_502,In_492);
xor U484 (N_484,In_730,In_297);
nor U485 (N_485,In_577,In_546);
xor U486 (N_486,In_569,In_15);
nand U487 (N_487,In_577,In_306);
nor U488 (N_488,In_373,In_232);
and U489 (N_489,In_421,In_301);
and U490 (N_490,In_541,In_110);
nor U491 (N_491,In_448,In_22);
xnor U492 (N_492,In_601,In_69);
nor U493 (N_493,In_250,In_130);
nand U494 (N_494,In_133,In_175);
nor U495 (N_495,In_740,In_738);
and U496 (N_496,In_409,In_111);
and U497 (N_497,In_97,In_729);
and U498 (N_498,In_402,In_629);
xnor U499 (N_499,In_37,In_741);
xor U500 (N_500,N_54,N_194);
or U501 (N_501,N_19,N_239);
nand U502 (N_502,N_353,N_136);
nor U503 (N_503,N_79,N_477);
nor U504 (N_504,N_163,N_62);
nor U505 (N_505,N_7,N_80);
or U506 (N_506,N_170,N_96);
xor U507 (N_507,N_15,N_2);
xor U508 (N_508,N_494,N_81);
xnor U509 (N_509,N_470,N_16);
xnor U510 (N_510,N_243,N_41);
xor U511 (N_511,N_162,N_236);
nor U512 (N_512,N_297,N_75);
nor U513 (N_513,N_175,N_283);
xnor U514 (N_514,N_418,N_231);
or U515 (N_515,N_390,N_253);
xnor U516 (N_516,N_171,N_109);
nand U517 (N_517,N_399,N_356);
nor U518 (N_518,N_174,N_310);
xnor U519 (N_519,N_13,N_201);
xnor U520 (N_520,N_261,N_139);
nand U521 (N_521,N_141,N_255);
nand U522 (N_522,N_188,N_360);
xor U523 (N_523,N_370,N_159);
and U524 (N_524,N_213,N_73);
nand U525 (N_525,N_298,N_212);
xor U526 (N_526,N_44,N_345);
and U527 (N_527,N_413,N_180);
or U528 (N_528,N_135,N_259);
or U529 (N_529,N_492,N_299);
or U530 (N_530,N_242,N_55);
and U531 (N_531,N_332,N_473);
nand U532 (N_532,N_300,N_435);
and U533 (N_533,N_486,N_344);
nand U534 (N_534,N_158,N_87);
nand U535 (N_535,N_206,N_482);
nor U536 (N_536,N_260,N_407);
nand U537 (N_537,N_191,N_184);
or U538 (N_538,N_207,N_113);
or U539 (N_539,N_308,N_319);
xnor U540 (N_540,N_257,N_46);
or U541 (N_541,N_409,N_265);
nor U542 (N_542,N_357,N_363);
xor U543 (N_543,N_183,N_304);
xor U544 (N_544,N_121,N_104);
and U545 (N_545,N_458,N_342);
xnor U546 (N_546,N_369,N_440);
or U547 (N_547,N_307,N_3);
and U548 (N_548,N_18,N_114);
nor U549 (N_549,N_416,N_425);
nor U550 (N_550,N_149,N_223);
nor U551 (N_551,N_336,N_66);
and U552 (N_552,N_388,N_221);
or U553 (N_553,N_35,N_431);
nand U554 (N_554,N_364,N_281);
nor U555 (N_555,N_325,N_177);
nor U556 (N_556,N_396,N_219);
nand U557 (N_557,N_198,N_67);
nand U558 (N_558,N_144,N_301);
and U559 (N_559,N_199,N_309);
nor U560 (N_560,N_89,N_200);
xor U561 (N_561,N_93,N_468);
or U562 (N_562,N_465,N_1);
and U563 (N_563,N_272,N_28);
xnor U564 (N_564,N_439,N_154);
or U565 (N_565,N_164,N_57);
and U566 (N_566,N_346,N_220);
or U567 (N_567,N_436,N_316);
nand U568 (N_568,N_197,N_419);
and U569 (N_569,N_248,N_90);
or U570 (N_570,N_64,N_25);
and U571 (N_571,N_214,N_444);
nand U572 (N_572,N_426,N_182);
xor U573 (N_573,N_112,N_71);
nand U574 (N_574,N_340,N_403);
or U575 (N_575,N_324,N_230);
and U576 (N_576,N_485,N_411);
xnor U577 (N_577,N_138,N_497);
nand U578 (N_578,N_251,N_445);
and U579 (N_579,N_499,N_6);
nor U580 (N_580,N_326,N_462);
or U581 (N_581,N_153,N_83);
nand U582 (N_582,N_186,N_247);
xnor U583 (N_583,N_480,N_21);
or U584 (N_584,N_467,N_389);
nand U585 (N_585,N_61,N_487);
nand U586 (N_586,N_250,N_289);
xor U587 (N_587,N_358,N_86);
xnor U588 (N_588,N_254,N_398);
xor U589 (N_589,N_117,N_167);
and U590 (N_590,N_120,N_422);
nand U591 (N_591,N_216,N_68);
nor U592 (N_592,N_447,N_394);
or U593 (N_593,N_208,N_305);
xnor U594 (N_594,N_382,N_488);
nand U595 (N_595,N_408,N_268);
or U596 (N_596,N_165,N_82);
and U597 (N_597,N_102,N_58);
and U598 (N_598,N_122,N_119);
xor U599 (N_599,N_267,N_116);
xnor U600 (N_600,N_65,N_293);
nand U601 (N_601,N_496,N_37);
nor U602 (N_602,N_303,N_217);
nand U603 (N_603,N_56,N_450);
nand U604 (N_604,N_78,N_161);
nor U605 (N_605,N_205,N_442);
xnor U606 (N_606,N_264,N_453);
or U607 (N_607,N_459,N_195);
or U608 (N_608,N_203,N_193);
nand U609 (N_609,N_52,N_328);
xor U610 (N_610,N_22,N_60);
or U611 (N_611,N_238,N_125);
or U612 (N_612,N_270,N_244);
nand U613 (N_613,N_352,N_155);
or U614 (N_614,N_263,N_245);
xor U615 (N_615,N_276,N_51);
xor U616 (N_616,N_140,N_282);
or U617 (N_617,N_339,N_373);
or U618 (N_618,N_126,N_329);
or U619 (N_619,N_348,N_24);
and U620 (N_620,N_38,N_279);
and U621 (N_621,N_386,N_266);
xnor U622 (N_622,N_45,N_375);
nand U623 (N_623,N_249,N_258);
and U624 (N_624,N_202,N_420);
xor U625 (N_625,N_189,N_311);
or U626 (N_626,N_72,N_150);
nor U627 (N_627,N_85,N_464);
nor U628 (N_628,N_179,N_443);
xor U629 (N_629,N_76,N_40);
xnor U630 (N_630,N_351,N_412);
or U631 (N_631,N_156,N_365);
xnor U632 (N_632,N_424,N_347);
nand U633 (N_633,N_317,N_63);
xnor U634 (N_634,N_315,N_457);
xor U635 (N_635,N_479,N_438);
and U636 (N_636,N_362,N_210);
nand U637 (N_637,N_70,N_49);
nor U638 (N_638,N_48,N_449);
or U639 (N_639,N_108,N_387);
nand U640 (N_640,N_277,N_490);
xnor U641 (N_641,N_423,N_133);
nand U642 (N_642,N_240,N_157);
nor U643 (N_643,N_50,N_484);
nor U644 (N_644,N_107,N_456);
or U645 (N_645,N_454,N_53);
nand U646 (N_646,N_404,N_94);
and U647 (N_647,N_4,N_137);
xor U648 (N_648,N_185,N_493);
and U649 (N_649,N_100,N_432);
nor U650 (N_650,N_291,N_290);
and U651 (N_651,N_256,N_475);
xnor U652 (N_652,N_30,N_483);
or U653 (N_653,N_173,N_478);
and U654 (N_654,N_190,N_84);
nor U655 (N_655,N_361,N_376);
xor U656 (N_656,N_43,N_211);
nand U657 (N_657,N_350,N_74);
and U658 (N_658,N_395,N_5);
and U659 (N_659,N_98,N_36);
nor U660 (N_660,N_323,N_381);
and U661 (N_661,N_318,N_481);
nor U662 (N_662,N_379,N_469);
nand U663 (N_663,N_143,N_437);
or U664 (N_664,N_218,N_131);
and U665 (N_665,N_17,N_451);
nor U666 (N_666,N_103,N_271);
xor U667 (N_667,N_26,N_47);
nor U668 (N_668,N_400,N_147);
xor U669 (N_669,N_384,N_430);
nor U670 (N_670,N_33,N_241);
nor U671 (N_671,N_142,N_472);
or U672 (N_672,N_225,N_287);
or U673 (N_673,N_355,N_8);
nor U674 (N_674,N_101,N_383);
or U675 (N_675,N_275,N_441);
and U676 (N_676,N_273,N_397);
or U677 (N_677,N_495,N_129);
nand U678 (N_678,N_229,N_295);
nor U679 (N_679,N_434,N_463);
nand U680 (N_680,N_343,N_335);
nand U681 (N_681,N_402,N_330);
and U682 (N_682,N_11,N_23);
nand U683 (N_683,N_14,N_172);
nand U684 (N_684,N_77,N_88);
nand U685 (N_685,N_127,N_392);
or U686 (N_686,N_187,N_476);
nand U687 (N_687,N_354,N_417);
nor U688 (N_688,N_331,N_237);
nand U689 (N_689,N_294,N_209);
or U690 (N_690,N_115,N_91);
nor U691 (N_691,N_489,N_192);
or U692 (N_692,N_372,N_92);
or U693 (N_693,N_146,N_320);
nand U694 (N_694,N_302,N_228);
or U695 (N_695,N_9,N_349);
xnor U696 (N_696,N_128,N_39);
and U697 (N_697,N_69,N_491);
nand U698 (N_698,N_366,N_429);
xnor U699 (N_699,N_160,N_274);
or U700 (N_700,N_460,N_176);
or U701 (N_701,N_59,N_284);
and U702 (N_702,N_168,N_410);
nor U703 (N_703,N_428,N_322);
and U704 (N_704,N_196,N_232);
or U705 (N_705,N_148,N_262);
and U706 (N_706,N_20,N_204);
and U707 (N_707,N_452,N_312);
nand U708 (N_708,N_433,N_393);
or U709 (N_709,N_246,N_29);
or U710 (N_710,N_466,N_314);
nand U711 (N_711,N_227,N_448);
xnor U712 (N_712,N_333,N_421);
xnor U713 (N_713,N_415,N_313);
or U714 (N_714,N_474,N_132);
and U715 (N_715,N_111,N_145);
nand U716 (N_716,N_105,N_374);
nor U717 (N_717,N_169,N_446);
or U718 (N_718,N_27,N_42);
nand U719 (N_719,N_178,N_461);
nor U720 (N_720,N_296,N_371);
or U721 (N_721,N_34,N_367);
nand U722 (N_722,N_124,N_368);
xor U723 (N_723,N_222,N_455);
nand U724 (N_724,N_130,N_405);
nor U725 (N_725,N_233,N_406);
xor U726 (N_726,N_414,N_134);
nand U727 (N_727,N_252,N_401);
xnor U728 (N_728,N_391,N_215);
and U729 (N_729,N_380,N_234);
and U730 (N_730,N_110,N_151);
and U731 (N_731,N_0,N_285);
or U732 (N_732,N_97,N_10);
xnor U733 (N_733,N_327,N_152);
or U734 (N_734,N_31,N_337);
or U735 (N_735,N_292,N_235);
nand U736 (N_736,N_338,N_359);
and U737 (N_737,N_32,N_226);
nand U738 (N_738,N_321,N_95);
or U739 (N_739,N_123,N_334);
nand U740 (N_740,N_377,N_269);
nand U741 (N_741,N_166,N_385);
or U742 (N_742,N_498,N_378);
nor U743 (N_743,N_306,N_286);
or U744 (N_744,N_341,N_288);
nand U745 (N_745,N_106,N_280);
or U746 (N_746,N_471,N_12);
xnor U747 (N_747,N_278,N_99);
and U748 (N_748,N_427,N_224);
and U749 (N_749,N_181,N_118);
nand U750 (N_750,N_112,N_89);
or U751 (N_751,N_178,N_239);
nor U752 (N_752,N_314,N_75);
nand U753 (N_753,N_257,N_218);
nor U754 (N_754,N_31,N_90);
nor U755 (N_755,N_148,N_440);
and U756 (N_756,N_324,N_326);
nand U757 (N_757,N_346,N_443);
nor U758 (N_758,N_423,N_238);
nor U759 (N_759,N_497,N_289);
xor U760 (N_760,N_319,N_171);
xor U761 (N_761,N_364,N_305);
nand U762 (N_762,N_323,N_27);
nand U763 (N_763,N_326,N_65);
or U764 (N_764,N_492,N_78);
nand U765 (N_765,N_52,N_467);
xor U766 (N_766,N_156,N_35);
and U767 (N_767,N_71,N_159);
and U768 (N_768,N_271,N_15);
and U769 (N_769,N_51,N_99);
nor U770 (N_770,N_355,N_26);
nand U771 (N_771,N_473,N_19);
nor U772 (N_772,N_444,N_29);
xnor U773 (N_773,N_351,N_461);
or U774 (N_774,N_30,N_222);
and U775 (N_775,N_175,N_465);
and U776 (N_776,N_476,N_354);
and U777 (N_777,N_445,N_439);
and U778 (N_778,N_364,N_491);
and U779 (N_779,N_61,N_101);
nand U780 (N_780,N_422,N_311);
xor U781 (N_781,N_458,N_405);
nor U782 (N_782,N_171,N_498);
nand U783 (N_783,N_269,N_271);
xor U784 (N_784,N_166,N_227);
nand U785 (N_785,N_250,N_370);
xor U786 (N_786,N_480,N_360);
or U787 (N_787,N_359,N_412);
and U788 (N_788,N_105,N_379);
nor U789 (N_789,N_117,N_168);
nor U790 (N_790,N_394,N_73);
and U791 (N_791,N_22,N_111);
or U792 (N_792,N_381,N_232);
nor U793 (N_793,N_241,N_114);
nand U794 (N_794,N_203,N_306);
nor U795 (N_795,N_17,N_480);
nand U796 (N_796,N_188,N_436);
or U797 (N_797,N_96,N_228);
nand U798 (N_798,N_36,N_413);
and U799 (N_799,N_4,N_315);
nor U800 (N_800,N_358,N_160);
nor U801 (N_801,N_104,N_311);
and U802 (N_802,N_425,N_451);
nand U803 (N_803,N_322,N_117);
and U804 (N_804,N_86,N_233);
nand U805 (N_805,N_158,N_78);
xor U806 (N_806,N_277,N_265);
nor U807 (N_807,N_29,N_102);
nor U808 (N_808,N_429,N_343);
or U809 (N_809,N_355,N_152);
xor U810 (N_810,N_305,N_430);
or U811 (N_811,N_206,N_192);
and U812 (N_812,N_316,N_166);
nor U813 (N_813,N_391,N_51);
or U814 (N_814,N_472,N_27);
or U815 (N_815,N_409,N_69);
nand U816 (N_816,N_133,N_353);
or U817 (N_817,N_44,N_363);
and U818 (N_818,N_385,N_437);
xor U819 (N_819,N_424,N_300);
nor U820 (N_820,N_358,N_435);
xor U821 (N_821,N_426,N_113);
or U822 (N_822,N_299,N_209);
nor U823 (N_823,N_53,N_174);
or U824 (N_824,N_48,N_204);
and U825 (N_825,N_335,N_292);
or U826 (N_826,N_329,N_209);
or U827 (N_827,N_330,N_371);
nand U828 (N_828,N_143,N_168);
nor U829 (N_829,N_282,N_217);
or U830 (N_830,N_289,N_304);
nor U831 (N_831,N_116,N_178);
nor U832 (N_832,N_155,N_83);
xnor U833 (N_833,N_140,N_453);
and U834 (N_834,N_226,N_61);
and U835 (N_835,N_275,N_94);
nand U836 (N_836,N_187,N_239);
xor U837 (N_837,N_353,N_486);
xnor U838 (N_838,N_193,N_459);
nor U839 (N_839,N_166,N_17);
and U840 (N_840,N_471,N_341);
xnor U841 (N_841,N_354,N_74);
or U842 (N_842,N_367,N_332);
or U843 (N_843,N_252,N_129);
xor U844 (N_844,N_64,N_266);
or U845 (N_845,N_191,N_168);
nor U846 (N_846,N_400,N_379);
nand U847 (N_847,N_259,N_106);
or U848 (N_848,N_94,N_39);
or U849 (N_849,N_492,N_384);
nor U850 (N_850,N_450,N_364);
and U851 (N_851,N_463,N_269);
xnor U852 (N_852,N_483,N_6);
and U853 (N_853,N_384,N_381);
nand U854 (N_854,N_26,N_406);
nor U855 (N_855,N_488,N_289);
and U856 (N_856,N_115,N_194);
or U857 (N_857,N_327,N_148);
or U858 (N_858,N_321,N_212);
nand U859 (N_859,N_481,N_483);
nand U860 (N_860,N_343,N_307);
or U861 (N_861,N_228,N_219);
nand U862 (N_862,N_7,N_193);
nor U863 (N_863,N_425,N_364);
xor U864 (N_864,N_415,N_271);
nand U865 (N_865,N_469,N_63);
or U866 (N_866,N_360,N_323);
xnor U867 (N_867,N_50,N_243);
xnor U868 (N_868,N_80,N_490);
xor U869 (N_869,N_16,N_379);
nor U870 (N_870,N_16,N_390);
nor U871 (N_871,N_177,N_15);
and U872 (N_872,N_66,N_43);
nand U873 (N_873,N_185,N_140);
and U874 (N_874,N_314,N_450);
xnor U875 (N_875,N_295,N_48);
nor U876 (N_876,N_279,N_345);
nor U877 (N_877,N_135,N_293);
and U878 (N_878,N_363,N_494);
and U879 (N_879,N_303,N_21);
nor U880 (N_880,N_419,N_392);
xnor U881 (N_881,N_82,N_383);
or U882 (N_882,N_339,N_233);
or U883 (N_883,N_362,N_293);
nand U884 (N_884,N_222,N_398);
or U885 (N_885,N_309,N_76);
nor U886 (N_886,N_182,N_354);
or U887 (N_887,N_0,N_401);
or U888 (N_888,N_188,N_77);
nor U889 (N_889,N_368,N_406);
or U890 (N_890,N_319,N_278);
or U891 (N_891,N_57,N_337);
or U892 (N_892,N_392,N_310);
or U893 (N_893,N_175,N_362);
xnor U894 (N_894,N_226,N_140);
and U895 (N_895,N_411,N_0);
nor U896 (N_896,N_443,N_25);
xnor U897 (N_897,N_480,N_54);
and U898 (N_898,N_484,N_372);
nor U899 (N_899,N_78,N_435);
and U900 (N_900,N_256,N_407);
xor U901 (N_901,N_292,N_461);
xnor U902 (N_902,N_161,N_269);
or U903 (N_903,N_401,N_178);
and U904 (N_904,N_0,N_361);
or U905 (N_905,N_332,N_386);
and U906 (N_906,N_438,N_0);
nor U907 (N_907,N_316,N_161);
nand U908 (N_908,N_246,N_71);
or U909 (N_909,N_93,N_216);
xor U910 (N_910,N_60,N_100);
nand U911 (N_911,N_381,N_237);
nand U912 (N_912,N_437,N_444);
nand U913 (N_913,N_8,N_290);
and U914 (N_914,N_469,N_38);
nor U915 (N_915,N_377,N_415);
nand U916 (N_916,N_449,N_269);
or U917 (N_917,N_113,N_95);
xor U918 (N_918,N_354,N_349);
nor U919 (N_919,N_13,N_153);
or U920 (N_920,N_231,N_406);
nand U921 (N_921,N_154,N_441);
xor U922 (N_922,N_242,N_376);
nor U923 (N_923,N_60,N_111);
nand U924 (N_924,N_209,N_347);
and U925 (N_925,N_13,N_241);
or U926 (N_926,N_80,N_240);
xnor U927 (N_927,N_307,N_108);
nand U928 (N_928,N_331,N_157);
nor U929 (N_929,N_480,N_16);
nor U930 (N_930,N_276,N_486);
or U931 (N_931,N_189,N_136);
and U932 (N_932,N_192,N_166);
nand U933 (N_933,N_226,N_87);
xor U934 (N_934,N_347,N_167);
and U935 (N_935,N_413,N_383);
xor U936 (N_936,N_7,N_229);
nor U937 (N_937,N_360,N_245);
xor U938 (N_938,N_115,N_150);
or U939 (N_939,N_350,N_292);
xnor U940 (N_940,N_30,N_421);
nor U941 (N_941,N_295,N_158);
and U942 (N_942,N_423,N_242);
and U943 (N_943,N_342,N_392);
nand U944 (N_944,N_452,N_310);
or U945 (N_945,N_26,N_290);
nor U946 (N_946,N_452,N_174);
or U947 (N_947,N_424,N_238);
or U948 (N_948,N_163,N_479);
nor U949 (N_949,N_428,N_215);
or U950 (N_950,N_453,N_392);
nand U951 (N_951,N_100,N_156);
or U952 (N_952,N_446,N_406);
nand U953 (N_953,N_37,N_96);
nand U954 (N_954,N_34,N_91);
and U955 (N_955,N_61,N_24);
nand U956 (N_956,N_160,N_89);
nand U957 (N_957,N_204,N_14);
and U958 (N_958,N_432,N_113);
nor U959 (N_959,N_437,N_264);
nand U960 (N_960,N_240,N_309);
and U961 (N_961,N_24,N_498);
nor U962 (N_962,N_146,N_83);
xnor U963 (N_963,N_193,N_426);
nor U964 (N_964,N_496,N_380);
xor U965 (N_965,N_24,N_18);
nor U966 (N_966,N_244,N_414);
and U967 (N_967,N_405,N_320);
nand U968 (N_968,N_104,N_370);
and U969 (N_969,N_367,N_144);
nor U970 (N_970,N_310,N_371);
or U971 (N_971,N_241,N_370);
and U972 (N_972,N_110,N_143);
xnor U973 (N_973,N_332,N_477);
nand U974 (N_974,N_221,N_137);
xnor U975 (N_975,N_377,N_111);
and U976 (N_976,N_383,N_370);
nand U977 (N_977,N_371,N_430);
nor U978 (N_978,N_290,N_99);
xor U979 (N_979,N_66,N_369);
and U980 (N_980,N_487,N_436);
and U981 (N_981,N_101,N_357);
or U982 (N_982,N_71,N_97);
and U983 (N_983,N_425,N_437);
or U984 (N_984,N_289,N_109);
nand U985 (N_985,N_442,N_3);
nor U986 (N_986,N_341,N_97);
or U987 (N_987,N_294,N_397);
and U988 (N_988,N_189,N_310);
nand U989 (N_989,N_366,N_352);
nor U990 (N_990,N_171,N_49);
nor U991 (N_991,N_481,N_407);
nor U992 (N_992,N_75,N_186);
nor U993 (N_993,N_481,N_221);
or U994 (N_994,N_382,N_277);
and U995 (N_995,N_325,N_74);
xnor U996 (N_996,N_495,N_444);
nand U997 (N_997,N_485,N_313);
nand U998 (N_998,N_108,N_278);
nor U999 (N_999,N_275,N_322);
xnor U1000 (N_1000,N_569,N_998);
or U1001 (N_1001,N_836,N_536);
or U1002 (N_1002,N_814,N_667);
xnor U1003 (N_1003,N_744,N_834);
nand U1004 (N_1004,N_660,N_523);
nor U1005 (N_1005,N_923,N_788);
nor U1006 (N_1006,N_764,N_867);
nor U1007 (N_1007,N_518,N_960);
or U1008 (N_1008,N_855,N_608);
nand U1009 (N_1009,N_880,N_731);
or U1010 (N_1010,N_500,N_884);
nand U1011 (N_1011,N_937,N_721);
nand U1012 (N_1012,N_758,N_784);
or U1013 (N_1013,N_771,N_975);
or U1014 (N_1014,N_920,N_850);
or U1015 (N_1015,N_635,N_773);
xnor U1016 (N_1016,N_992,N_597);
nor U1017 (N_1017,N_696,N_989);
nor U1018 (N_1018,N_822,N_887);
nor U1019 (N_1019,N_882,N_800);
nand U1020 (N_1020,N_554,N_953);
or U1021 (N_1021,N_748,N_645);
nand U1022 (N_1022,N_900,N_795);
nor U1023 (N_1023,N_540,N_665);
xnor U1024 (N_1024,N_873,N_976);
and U1025 (N_1025,N_985,N_827);
xnor U1026 (N_1026,N_664,N_505);
or U1027 (N_1027,N_737,N_778);
xor U1028 (N_1028,N_627,N_993);
nor U1029 (N_1029,N_863,N_915);
or U1030 (N_1030,N_934,N_720);
xor U1031 (N_1031,N_925,N_892);
and U1032 (N_1032,N_755,N_751);
nand U1033 (N_1033,N_969,N_567);
nand U1034 (N_1034,N_579,N_545);
xor U1035 (N_1035,N_534,N_668);
nor U1036 (N_1036,N_564,N_675);
nand U1037 (N_1037,N_861,N_826);
or U1038 (N_1038,N_657,N_946);
xnor U1039 (N_1039,N_609,N_595);
or U1040 (N_1040,N_772,N_648);
and U1041 (N_1041,N_869,N_835);
or U1042 (N_1042,N_629,N_914);
or U1043 (N_1043,N_824,N_565);
xnor U1044 (N_1044,N_828,N_733);
xor U1045 (N_1045,N_522,N_694);
nand U1046 (N_1046,N_739,N_762);
nor U1047 (N_1047,N_947,N_966);
nor U1048 (N_1048,N_705,N_576);
and U1049 (N_1049,N_654,N_699);
and U1050 (N_1050,N_890,N_805);
and U1051 (N_1051,N_622,N_789);
xor U1052 (N_1052,N_911,N_531);
xor U1053 (N_1053,N_831,N_996);
nand U1054 (N_1054,N_501,N_590);
or U1055 (N_1055,N_905,N_986);
nand U1056 (N_1056,N_601,N_700);
and U1057 (N_1057,N_684,N_899);
or U1058 (N_1058,N_987,N_752);
and U1059 (N_1059,N_922,N_671);
and U1060 (N_1060,N_803,N_901);
and U1061 (N_1061,N_709,N_820);
and U1062 (N_1062,N_678,N_723);
nand U1063 (N_1063,N_630,N_692);
nand U1064 (N_1064,N_906,N_853);
nor U1065 (N_1065,N_729,N_988);
nor U1066 (N_1066,N_690,N_766);
nand U1067 (N_1067,N_504,N_971);
nor U1068 (N_1068,N_647,N_615);
xor U1069 (N_1069,N_706,N_735);
nand U1070 (N_1070,N_812,N_963);
or U1071 (N_1071,N_682,N_715);
xor U1072 (N_1072,N_825,N_883);
nor U1073 (N_1073,N_859,N_991);
or U1074 (N_1074,N_543,N_559);
or U1075 (N_1075,N_525,N_613);
xor U1076 (N_1076,N_703,N_769);
nor U1077 (N_1077,N_984,N_681);
xnor U1078 (N_1078,N_982,N_624);
xnor U1079 (N_1079,N_929,N_978);
xor U1080 (N_1080,N_584,N_713);
nand U1081 (N_1081,N_550,N_908);
nand U1082 (N_1082,N_589,N_626);
and U1083 (N_1083,N_943,N_889);
and U1084 (N_1084,N_756,N_782);
and U1085 (N_1085,N_533,N_885);
nand U1086 (N_1086,N_964,N_509);
nand U1087 (N_1087,N_602,N_549);
nor U1088 (N_1088,N_585,N_542);
and U1089 (N_1089,N_651,N_895);
nand U1090 (N_1090,N_663,N_572);
or U1091 (N_1091,N_616,N_801);
xnor U1092 (N_1092,N_990,N_672);
xnor U1093 (N_1093,N_631,N_860);
nand U1094 (N_1094,N_965,N_979);
and U1095 (N_1095,N_575,N_952);
and U1096 (N_1096,N_718,N_605);
nor U1097 (N_1097,N_747,N_833);
or U1098 (N_1098,N_750,N_650);
xor U1099 (N_1099,N_661,N_693);
xor U1100 (N_1100,N_849,N_552);
xnor U1101 (N_1101,N_865,N_621);
xor U1102 (N_1102,N_872,N_603);
xnor U1103 (N_1103,N_819,N_902);
nand U1104 (N_1104,N_507,N_817);
nor U1105 (N_1105,N_674,N_972);
and U1106 (N_1106,N_583,N_913);
and U1107 (N_1107,N_931,N_529);
or U1108 (N_1108,N_767,N_754);
nand U1109 (N_1109,N_717,N_612);
xnor U1110 (N_1110,N_578,N_786);
or U1111 (N_1111,N_916,N_673);
and U1112 (N_1112,N_761,N_727);
nand U1113 (N_1113,N_864,N_832);
xnor U1114 (N_1114,N_676,N_888);
nor U1115 (N_1115,N_924,N_806);
and U1116 (N_1116,N_740,N_598);
nor U1117 (N_1117,N_607,N_876);
nor U1118 (N_1118,N_926,N_845);
nor U1119 (N_1119,N_556,N_874);
nand U1120 (N_1120,N_881,N_830);
nor U1121 (N_1121,N_539,N_623);
nor U1122 (N_1122,N_956,N_821);
nand U1123 (N_1123,N_907,N_637);
nand U1124 (N_1124,N_712,N_516);
and U1125 (N_1125,N_999,N_606);
and U1126 (N_1126,N_753,N_512);
nand U1127 (N_1127,N_967,N_646);
and U1128 (N_1128,N_639,N_701);
nor U1129 (N_1129,N_599,N_878);
or U1130 (N_1130,N_958,N_927);
xnor U1131 (N_1131,N_765,N_847);
xor U1132 (N_1132,N_634,N_877);
or U1133 (N_1133,N_759,N_656);
or U1134 (N_1134,N_810,N_617);
nand U1135 (N_1135,N_632,N_734);
nor U1136 (N_1136,N_823,N_796);
nand U1137 (N_1137,N_513,N_840);
nor U1138 (N_1138,N_535,N_560);
xnor U1139 (N_1139,N_918,N_868);
xnor U1140 (N_1140,N_571,N_891);
and U1141 (N_1141,N_614,N_945);
xnor U1142 (N_1142,N_852,N_866);
and U1143 (N_1143,N_798,N_679);
and U1144 (N_1144,N_577,N_879);
or U1145 (N_1145,N_746,N_936);
nor U1146 (N_1146,N_686,N_846);
nor U1147 (N_1147,N_994,N_652);
and U1148 (N_1148,N_837,N_582);
or U1149 (N_1149,N_511,N_625);
or U1150 (N_1150,N_611,N_618);
xnor U1151 (N_1151,N_983,N_558);
xor U1152 (N_1152,N_555,N_593);
xnor U1153 (N_1153,N_851,N_655);
and U1154 (N_1154,N_677,N_815);
and U1155 (N_1155,N_757,N_544);
and U1156 (N_1156,N_980,N_763);
and U1157 (N_1157,N_955,N_743);
and U1158 (N_1158,N_548,N_526);
xor U1159 (N_1159,N_521,N_697);
nor U1160 (N_1160,N_856,N_776);
xor U1161 (N_1161,N_875,N_503);
nor U1162 (N_1162,N_506,N_928);
or U1163 (N_1163,N_502,N_530);
nand U1164 (N_1164,N_508,N_592);
or U1165 (N_1165,N_981,N_843);
or U1166 (N_1166,N_790,N_581);
or U1167 (N_1167,N_719,N_642);
nand U1168 (N_1168,N_760,N_961);
nor U1169 (N_1169,N_939,N_780);
and U1170 (N_1170,N_546,N_933);
or U1171 (N_1171,N_551,N_722);
or U1172 (N_1172,N_842,N_775);
nor U1173 (N_1173,N_968,N_527);
xnor U1174 (N_1174,N_745,N_944);
and U1175 (N_1175,N_689,N_970);
nor U1176 (N_1176,N_553,N_770);
xor U1177 (N_1177,N_586,N_519);
xnor U1178 (N_1178,N_666,N_844);
xnor U1179 (N_1179,N_561,N_580);
nor U1180 (N_1180,N_841,N_711);
xnor U1181 (N_1181,N_541,N_949);
xnor U1182 (N_1182,N_816,N_641);
nand U1183 (N_1183,N_691,N_520);
xnor U1184 (N_1184,N_594,N_683);
nand U1185 (N_1185,N_610,N_685);
nor U1186 (N_1186,N_557,N_951);
xor U1187 (N_1187,N_793,N_716);
nand U1188 (N_1188,N_620,N_932);
nor U1189 (N_1189,N_724,N_959);
nand U1190 (N_1190,N_568,N_858);
nor U1191 (N_1191,N_813,N_871);
xnor U1192 (N_1192,N_818,N_510);
or U1193 (N_1193,N_538,N_909);
xnor U1194 (N_1194,N_997,N_741);
or U1195 (N_1195,N_562,N_854);
and U1196 (N_1196,N_528,N_862);
and U1197 (N_1197,N_948,N_728);
or U1198 (N_1198,N_942,N_628);
nor U1199 (N_1199,N_829,N_941);
xnor U1200 (N_1200,N_777,N_514);
nand U1201 (N_1201,N_768,N_649);
or U1202 (N_1202,N_710,N_794);
xor U1203 (N_1203,N_566,N_698);
nand U1204 (N_1204,N_687,N_604);
and U1205 (N_1205,N_524,N_848);
and U1206 (N_1206,N_930,N_898);
nand U1207 (N_1207,N_730,N_957);
xor U1208 (N_1208,N_659,N_783);
and U1209 (N_1209,N_532,N_894);
nor U1210 (N_1210,N_940,N_839);
xnor U1211 (N_1211,N_857,N_954);
nor U1212 (N_1212,N_702,N_738);
xnor U1213 (N_1213,N_732,N_726);
or U1214 (N_1214,N_785,N_973);
xnor U1215 (N_1215,N_636,N_977);
or U1216 (N_1216,N_791,N_633);
nor U1217 (N_1217,N_809,N_537);
nor U1218 (N_1218,N_570,N_781);
xnor U1219 (N_1219,N_870,N_670);
nor U1220 (N_1220,N_662,N_669);
and U1221 (N_1221,N_688,N_574);
xor U1222 (N_1222,N_680,N_787);
and U1223 (N_1223,N_725,N_910);
and U1224 (N_1224,N_792,N_695);
nor U1225 (N_1225,N_591,N_749);
nor U1226 (N_1226,N_802,N_950);
or U1227 (N_1227,N_904,N_807);
nand U1228 (N_1228,N_573,N_774);
or U1229 (N_1229,N_547,N_779);
nor U1230 (N_1230,N_896,N_515);
xnor U1231 (N_1231,N_919,N_797);
nor U1232 (N_1232,N_912,N_903);
and U1233 (N_1233,N_563,N_838);
or U1234 (N_1234,N_653,N_707);
nor U1235 (N_1235,N_704,N_893);
xor U1236 (N_1236,N_742,N_587);
xnor U1237 (N_1237,N_886,N_808);
nor U1238 (N_1238,N_658,N_995);
nand U1239 (N_1239,N_799,N_588);
nor U1240 (N_1240,N_600,N_935);
and U1241 (N_1241,N_714,N_974);
or U1242 (N_1242,N_811,N_644);
nand U1243 (N_1243,N_596,N_643);
nand U1244 (N_1244,N_921,N_638);
nor U1245 (N_1245,N_917,N_708);
nand U1246 (N_1246,N_938,N_804);
or U1247 (N_1247,N_736,N_640);
xnor U1248 (N_1248,N_897,N_962);
xor U1249 (N_1249,N_517,N_619);
and U1250 (N_1250,N_632,N_822);
nand U1251 (N_1251,N_641,N_558);
nor U1252 (N_1252,N_682,N_767);
nand U1253 (N_1253,N_749,N_729);
or U1254 (N_1254,N_684,N_523);
or U1255 (N_1255,N_873,N_798);
nand U1256 (N_1256,N_733,N_746);
or U1257 (N_1257,N_624,N_986);
or U1258 (N_1258,N_904,N_994);
nand U1259 (N_1259,N_863,N_855);
and U1260 (N_1260,N_977,N_862);
xnor U1261 (N_1261,N_538,N_963);
and U1262 (N_1262,N_601,N_811);
nand U1263 (N_1263,N_856,N_583);
nor U1264 (N_1264,N_646,N_891);
nand U1265 (N_1265,N_562,N_528);
nand U1266 (N_1266,N_673,N_925);
nand U1267 (N_1267,N_876,N_958);
nand U1268 (N_1268,N_608,N_739);
or U1269 (N_1269,N_807,N_731);
or U1270 (N_1270,N_891,N_789);
or U1271 (N_1271,N_789,N_661);
nand U1272 (N_1272,N_894,N_969);
nand U1273 (N_1273,N_539,N_603);
nor U1274 (N_1274,N_556,N_807);
xor U1275 (N_1275,N_813,N_951);
nor U1276 (N_1276,N_635,N_584);
or U1277 (N_1277,N_994,N_503);
or U1278 (N_1278,N_850,N_703);
and U1279 (N_1279,N_550,N_812);
and U1280 (N_1280,N_938,N_726);
xnor U1281 (N_1281,N_920,N_977);
xnor U1282 (N_1282,N_906,N_947);
nand U1283 (N_1283,N_834,N_641);
nor U1284 (N_1284,N_829,N_692);
nor U1285 (N_1285,N_844,N_660);
xnor U1286 (N_1286,N_871,N_884);
xnor U1287 (N_1287,N_985,N_568);
nor U1288 (N_1288,N_557,N_706);
nor U1289 (N_1289,N_997,N_515);
or U1290 (N_1290,N_672,N_749);
and U1291 (N_1291,N_851,N_782);
xnor U1292 (N_1292,N_671,N_604);
xnor U1293 (N_1293,N_716,N_837);
or U1294 (N_1294,N_606,N_621);
nand U1295 (N_1295,N_949,N_670);
and U1296 (N_1296,N_984,N_537);
or U1297 (N_1297,N_870,N_794);
xor U1298 (N_1298,N_693,N_634);
nor U1299 (N_1299,N_621,N_728);
and U1300 (N_1300,N_926,N_980);
xor U1301 (N_1301,N_904,N_688);
xnor U1302 (N_1302,N_544,N_712);
nand U1303 (N_1303,N_810,N_654);
or U1304 (N_1304,N_952,N_679);
and U1305 (N_1305,N_593,N_540);
nand U1306 (N_1306,N_966,N_682);
nand U1307 (N_1307,N_584,N_887);
or U1308 (N_1308,N_823,N_592);
nor U1309 (N_1309,N_525,N_758);
and U1310 (N_1310,N_642,N_966);
xnor U1311 (N_1311,N_931,N_803);
xor U1312 (N_1312,N_638,N_569);
xnor U1313 (N_1313,N_621,N_507);
nand U1314 (N_1314,N_720,N_794);
and U1315 (N_1315,N_646,N_634);
nand U1316 (N_1316,N_811,N_599);
nand U1317 (N_1317,N_618,N_796);
or U1318 (N_1318,N_854,N_834);
nor U1319 (N_1319,N_867,N_963);
nor U1320 (N_1320,N_808,N_836);
nor U1321 (N_1321,N_720,N_572);
xor U1322 (N_1322,N_616,N_659);
nor U1323 (N_1323,N_573,N_949);
nand U1324 (N_1324,N_620,N_763);
nor U1325 (N_1325,N_541,N_804);
nand U1326 (N_1326,N_990,N_896);
xnor U1327 (N_1327,N_839,N_659);
and U1328 (N_1328,N_544,N_950);
nand U1329 (N_1329,N_730,N_699);
or U1330 (N_1330,N_892,N_814);
and U1331 (N_1331,N_680,N_524);
and U1332 (N_1332,N_886,N_757);
xnor U1333 (N_1333,N_647,N_906);
nor U1334 (N_1334,N_873,N_672);
or U1335 (N_1335,N_717,N_607);
and U1336 (N_1336,N_600,N_877);
or U1337 (N_1337,N_819,N_559);
nand U1338 (N_1338,N_784,N_891);
and U1339 (N_1339,N_678,N_544);
xnor U1340 (N_1340,N_899,N_812);
xor U1341 (N_1341,N_898,N_792);
nand U1342 (N_1342,N_610,N_876);
nor U1343 (N_1343,N_620,N_660);
nand U1344 (N_1344,N_701,N_553);
and U1345 (N_1345,N_655,N_627);
and U1346 (N_1346,N_610,N_874);
and U1347 (N_1347,N_527,N_992);
nor U1348 (N_1348,N_955,N_854);
nand U1349 (N_1349,N_505,N_636);
nor U1350 (N_1350,N_558,N_708);
nand U1351 (N_1351,N_634,N_916);
and U1352 (N_1352,N_586,N_671);
and U1353 (N_1353,N_820,N_878);
and U1354 (N_1354,N_500,N_740);
or U1355 (N_1355,N_993,N_579);
and U1356 (N_1356,N_502,N_597);
xnor U1357 (N_1357,N_943,N_580);
and U1358 (N_1358,N_719,N_994);
or U1359 (N_1359,N_951,N_552);
nand U1360 (N_1360,N_817,N_502);
xnor U1361 (N_1361,N_810,N_695);
and U1362 (N_1362,N_793,N_995);
nand U1363 (N_1363,N_993,N_804);
nor U1364 (N_1364,N_571,N_986);
nand U1365 (N_1365,N_664,N_762);
and U1366 (N_1366,N_946,N_725);
and U1367 (N_1367,N_961,N_605);
nand U1368 (N_1368,N_591,N_805);
or U1369 (N_1369,N_912,N_919);
xor U1370 (N_1370,N_546,N_720);
or U1371 (N_1371,N_799,N_762);
and U1372 (N_1372,N_574,N_828);
or U1373 (N_1373,N_514,N_973);
nand U1374 (N_1374,N_605,N_936);
and U1375 (N_1375,N_598,N_803);
and U1376 (N_1376,N_713,N_662);
and U1377 (N_1377,N_588,N_955);
or U1378 (N_1378,N_748,N_807);
nand U1379 (N_1379,N_931,N_690);
nor U1380 (N_1380,N_993,N_714);
xnor U1381 (N_1381,N_919,N_994);
nand U1382 (N_1382,N_775,N_962);
nand U1383 (N_1383,N_978,N_859);
nand U1384 (N_1384,N_653,N_684);
nor U1385 (N_1385,N_900,N_853);
or U1386 (N_1386,N_703,N_809);
or U1387 (N_1387,N_779,N_832);
nand U1388 (N_1388,N_521,N_684);
nand U1389 (N_1389,N_957,N_530);
or U1390 (N_1390,N_628,N_649);
nor U1391 (N_1391,N_721,N_674);
xor U1392 (N_1392,N_666,N_965);
and U1393 (N_1393,N_507,N_658);
or U1394 (N_1394,N_728,N_603);
or U1395 (N_1395,N_545,N_617);
nand U1396 (N_1396,N_853,N_627);
or U1397 (N_1397,N_799,N_887);
or U1398 (N_1398,N_910,N_797);
nand U1399 (N_1399,N_832,N_532);
and U1400 (N_1400,N_644,N_604);
nand U1401 (N_1401,N_825,N_872);
nand U1402 (N_1402,N_886,N_799);
or U1403 (N_1403,N_990,N_879);
nor U1404 (N_1404,N_910,N_552);
or U1405 (N_1405,N_574,N_970);
nand U1406 (N_1406,N_788,N_603);
or U1407 (N_1407,N_735,N_894);
nor U1408 (N_1408,N_692,N_570);
xor U1409 (N_1409,N_641,N_801);
nor U1410 (N_1410,N_604,N_605);
or U1411 (N_1411,N_594,N_883);
and U1412 (N_1412,N_595,N_656);
nor U1413 (N_1413,N_600,N_691);
or U1414 (N_1414,N_723,N_807);
xnor U1415 (N_1415,N_908,N_500);
nor U1416 (N_1416,N_907,N_814);
nand U1417 (N_1417,N_570,N_816);
and U1418 (N_1418,N_905,N_845);
and U1419 (N_1419,N_879,N_819);
nor U1420 (N_1420,N_574,N_640);
or U1421 (N_1421,N_770,N_579);
nor U1422 (N_1422,N_657,N_567);
nand U1423 (N_1423,N_968,N_877);
and U1424 (N_1424,N_792,N_615);
or U1425 (N_1425,N_552,N_639);
nor U1426 (N_1426,N_519,N_555);
nor U1427 (N_1427,N_517,N_681);
xnor U1428 (N_1428,N_506,N_855);
nor U1429 (N_1429,N_561,N_963);
nor U1430 (N_1430,N_750,N_639);
nor U1431 (N_1431,N_800,N_623);
and U1432 (N_1432,N_619,N_597);
or U1433 (N_1433,N_572,N_745);
and U1434 (N_1434,N_846,N_687);
nand U1435 (N_1435,N_625,N_555);
xor U1436 (N_1436,N_816,N_624);
nor U1437 (N_1437,N_638,N_564);
or U1438 (N_1438,N_910,N_613);
or U1439 (N_1439,N_714,N_764);
and U1440 (N_1440,N_748,N_865);
or U1441 (N_1441,N_887,N_756);
nand U1442 (N_1442,N_648,N_562);
nand U1443 (N_1443,N_528,N_704);
and U1444 (N_1444,N_788,N_550);
nand U1445 (N_1445,N_606,N_746);
xnor U1446 (N_1446,N_898,N_660);
or U1447 (N_1447,N_695,N_540);
nand U1448 (N_1448,N_924,N_872);
and U1449 (N_1449,N_968,N_685);
and U1450 (N_1450,N_677,N_574);
or U1451 (N_1451,N_770,N_560);
xnor U1452 (N_1452,N_870,N_756);
or U1453 (N_1453,N_631,N_994);
nor U1454 (N_1454,N_916,N_748);
nor U1455 (N_1455,N_631,N_996);
nand U1456 (N_1456,N_874,N_550);
and U1457 (N_1457,N_678,N_809);
nor U1458 (N_1458,N_831,N_827);
or U1459 (N_1459,N_905,N_547);
or U1460 (N_1460,N_724,N_520);
or U1461 (N_1461,N_924,N_786);
xnor U1462 (N_1462,N_736,N_660);
xnor U1463 (N_1463,N_719,N_916);
or U1464 (N_1464,N_969,N_775);
or U1465 (N_1465,N_574,N_861);
nor U1466 (N_1466,N_520,N_631);
nor U1467 (N_1467,N_763,N_589);
nand U1468 (N_1468,N_500,N_705);
and U1469 (N_1469,N_576,N_939);
and U1470 (N_1470,N_581,N_793);
nor U1471 (N_1471,N_658,N_721);
or U1472 (N_1472,N_733,N_861);
nor U1473 (N_1473,N_685,N_603);
or U1474 (N_1474,N_767,N_716);
and U1475 (N_1475,N_720,N_765);
nand U1476 (N_1476,N_995,N_810);
and U1477 (N_1477,N_611,N_815);
or U1478 (N_1478,N_650,N_510);
xnor U1479 (N_1479,N_995,N_781);
nor U1480 (N_1480,N_923,N_744);
xnor U1481 (N_1481,N_648,N_766);
xor U1482 (N_1482,N_568,N_731);
and U1483 (N_1483,N_670,N_965);
nor U1484 (N_1484,N_953,N_862);
or U1485 (N_1485,N_903,N_849);
nor U1486 (N_1486,N_576,N_754);
and U1487 (N_1487,N_965,N_795);
and U1488 (N_1488,N_718,N_563);
xnor U1489 (N_1489,N_550,N_725);
xnor U1490 (N_1490,N_698,N_930);
or U1491 (N_1491,N_955,N_862);
xor U1492 (N_1492,N_693,N_620);
nand U1493 (N_1493,N_837,N_520);
nand U1494 (N_1494,N_621,N_820);
nand U1495 (N_1495,N_649,N_762);
nor U1496 (N_1496,N_982,N_888);
xnor U1497 (N_1497,N_764,N_579);
or U1498 (N_1498,N_921,N_720);
xor U1499 (N_1499,N_896,N_662);
xor U1500 (N_1500,N_1400,N_1037);
xor U1501 (N_1501,N_1484,N_1067);
nand U1502 (N_1502,N_1051,N_1423);
xnor U1503 (N_1503,N_1015,N_1011);
xor U1504 (N_1504,N_1379,N_1445);
and U1505 (N_1505,N_1338,N_1381);
nor U1506 (N_1506,N_1157,N_1256);
nor U1507 (N_1507,N_1479,N_1411);
or U1508 (N_1508,N_1207,N_1419);
or U1509 (N_1509,N_1402,N_1125);
and U1510 (N_1510,N_1388,N_1000);
or U1511 (N_1511,N_1174,N_1196);
nor U1512 (N_1512,N_1418,N_1105);
nand U1513 (N_1513,N_1062,N_1261);
nor U1514 (N_1514,N_1211,N_1118);
xor U1515 (N_1515,N_1336,N_1109);
xnor U1516 (N_1516,N_1122,N_1425);
xnor U1517 (N_1517,N_1112,N_1369);
or U1518 (N_1518,N_1343,N_1415);
or U1519 (N_1519,N_1202,N_1451);
xnor U1520 (N_1520,N_1367,N_1263);
nor U1521 (N_1521,N_1018,N_1088);
and U1522 (N_1522,N_1454,N_1021);
or U1523 (N_1523,N_1246,N_1030);
and U1524 (N_1524,N_1189,N_1465);
or U1525 (N_1525,N_1123,N_1007);
nor U1526 (N_1526,N_1472,N_1329);
or U1527 (N_1527,N_1072,N_1092);
nand U1528 (N_1528,N_1310,N_1097);
nor U1529 (N_1529,N_1131,N_1198);
or U1530 (N_1530,N_1101,N_1354);
nand U1531 (N_1531,N_1426,N_1351);
and U1532 (N_1532,N_1158,N_1442);
and U1533 (N_1533,N_1399,N_1382);
nand U1534 (N_1534,N_1358,N_1165);
or U1535 (N_1535,N_1141,N_1446);
xnor U1536 (N_1536,N_1373,N_1473);
nand U1537 (N_1537,N_1176,N_1318);
xnor U1538 (N_1538,N_1283,N_1124);
nand U1539 (N_1539,N_1155,N_1466);
xnor U1540 (N_1540,N_1190,N_1325);
or U1541 (N_1541,N_1081,N_1267);
or U1542 (N_1542,N_1339,N_1128);
xor U1543 (N_1543,N_1103,N_1002);
xnor U1544 (N_1544,N_1469,N_1042);
or U1545 (N_1545,N_1348,N_1273);
nand U1546 (N_1546,N_1416,N_1386);
nor U1547 (N_1547,N_1043,N_1396);
and U1548 (N_1548,N_1126,N_1491);
nand U1549 (N_1549,N_1129,N_1252);
and U1550 (N_1550,N_1323,N_1146);
xor U1551 (N_1551,N_1497,N_1182);
and U1552 (N_1552,N_1490,N_1020);
nand U1553 (N_1553,N_1347,N_1286);
nand U1554 (N_1554,N_1050,N_1245);
and U1555 (N_1555,N_1194,N_1242);
nor U1556 (N_1556,N_1188,N_1222);
nand U1557 (N_1557,N_1368,N_1333);
nand U1558 (N_1558,N_1147,N_1496);
xnor U1559 (N_1559,N_1375,N_1456);
xnor U1560 (N_1560,N_1397,N_1143);
or U1561 (N_1561,N_1055,N_1220);
and U1562 (N_1562,N_1407,N_1085);
or U1563 (N_1563,N_1107,N_1363);
nand U1564 (N_1564,N_1284,N_1074);
and U1565 (N_1565,N_1259,N_1178);
xnor U1566 (N_1566,N_1420,N_1319);
and U1567 (N_1567,N_1274,N_1299);
and U1568 (N_1568,N_1179,N_1172);
nor U1569 (N_1569,N_1295,N_1390);
nand U1570 (N_1570,N_1431,N_1216);
nor U1571 (N_1571,N_1095,N_1365);
nand U1572 (N_1572,N_1285,N_1251);
and U1573 (N_1573,N_1230,N_1461);
and U1574 (N_1574,N_1039,N_1340);
xnor U1575 (N_1575,N_1265,N_1385);
nand U1576 (N_1576,N_1485,N_1387);
nand U1577 (N_1577,N_1404,N_1080);
nor U1578 (N_1578,N_1200,N_1429);
and U1579 (N_1579,N_1183,N_1330);
nor U1580 (N_1580,N_1249,N_1291);
or U1581 (N_1581,N_1070,N_1254);
or U1582 (N_1582,N_1048,N_1093);
xor U1583 (N_1583,N_1059,N_1306);
and U1584 (N_1584,N_1239,N_1199);
xor U1585 (N_1585,N_1255,N_1040);
xor U1586 (N_1586,N_1495,N_1111);
nor U1587 (N_1587,N_1001,N_1352);
nor U1588 (N_1588,N_1403,N_1017);
or U1589 (N_1589,N_1433,N_1224);
nand U1590 (N_1590,N_1164,N_1296);
nand U1591 (N_1591,N_1214,N_1038);
or U1592 (N_1592,N_1448,N_1482);
nand U1593 (N_1593,N_1359,N_1241);
xor U1594 (N_1594,N_1405,N_1218);
nand U1595 (N_1595,N_1057,N_1135);
or U1596 (N_1596,N_1280,N_1498);
nand U1597 (N_1597,N_1444,N_1309);
nor U1598 (N_1598,N_1266,N_1409);
nand U1599 (N_1599,N_1116,N_1383);
and U1600 (N_1600,N_1314,N_1056);
nand U1601 (N_1601,N_1353,N_1374);
nand U1602 (N_1602,N_1140,N_1293);
and U1603 (N_1603,N_1003,N_1492);
nand U1604 (N_1604,N_1226,N_1455);
xor U1605 (N_1605,N_1238,N_1364);
and U1606 (N_1606,N_1228,N_1108);
xnor U1607 (N_1607,N_1428,N_1162);
or U1608 (N_1608,N_1424,N_1148);
nor U1609 (N_1609,N_1453,N_1237);
nor U1610 (N_1610,N_1082,N_1079);
and U1611 (N_1611,N_1392,N_1327);
and U1612 (N_1612,N_1225,N_1414);
or U1613 (N_1613,N_1227,N_1317);
nand U1614 (N_1614,N_1104,N_1153);
or U1615 (N_1615,N_1235,N_1212);
nor U1616 (N_1616,N_1380,N_1304);
and U1617 (N_1617,N_1271,N_1434);
xor U1618 (N_1618,N_1355,N_1247);
nor U1619 (N_1619,N_1278,N_1260);
xnor U1620 (N_1620,N_1217,N_1289);
or U1621 (N_1621,N_1195,N_1019);
and U1622 (N_1622,N_1337,N_1362);
or U1623 (N_1623,N_1058,N_1069);
xnor U1624 (N_1624,N_1290,N_1154);
nor U1625 (N_1625,N_1438,N_1012);
and U1626 (N_1626,N_1044,N_1134);
nand U1627 (N_1627,N_1145,N_1137);
xor U1628 (N_1628,N_1460,N_1471);
and U1629 (N_1629,N_1302,N_1136);
or U1630 (N_1630,N_1315,N_1294);
xnor U1631 (N_1631,N_1499,N_1096);
or U1632 (N_1632,N_1357,N_1269);
nand U1633 (N_1633,N_1467,N_1029);
nor U1634 (N_1634,N_1449,N_1360);
xnor U1635 (N_1635,N_1288,N_1150);
or U1636 (N_1636,N_1324,N_1031);
xnor U1637 (N_1637,N_1006,N_1268);
and U1638 (N_1638,N_1276,N_1394);
and U1639 (N_1639,N_1321,N_1168);
xor U1640 (N_1640,N_1076,N_1243);
xnor U1641 (N_1641,N_1110,N_1206);
and U1642 (N_1642,N_1435,N_1022);
or U1643 (N_1643,N_1275,N_1090);
and U1644 (N_1644,N_1087,N_1262);
nand U1645 (N_1645,N_1197,N_1287);
nand U1646 (N_1646,N_1332,N_1231);
or U1647 (N_1647,N_1421,N_1412);
or U1648 (N_1648,N_1106,N_1068);
nor U1649 (N_1649,N_1229,N_1341);
or U1650 (N_1650,N_1334,N_1257);
and U1651 (N_1651,N_1041,N_1361);
xor U1652 (N_1652,N_1077,N_1468);
or U1653 (N_1653,N_1459,N_1084);
nand U1654 (N_1654,N_1138,N_1026);
nor U1655 (N_1655,N_1311,N_1073);
nor U1656 (N_1656,N_1209,N_1349);
or U1657 (N_1657,N_1083,N_1481);
and U1658 (N_1658,N_1223,N_1253);
nand U1659 (N_1659,N_1078,N_1474);
or U1660 (N_1660,N_1487,N_1427);
or U1661 (N_1661,N_1205,N_1089);
and U1662 (N_1662,N_1091,N_1384);
or U1663 (N_1663,N_1398,N_1377);
nand U1664 (N_1664,N_1452,N_1114);
and U1665 (N_1665,N_1401,N_1475);
nor U1666 (N_1666,N_1023,N_1156);
nor U1667 (N_1667,N_1071,N_1066);
xnor U1668 (N_1668,N_1244,N_1410);
or U1669 (N_1669,N_1063,N_1447);
and U1670 (N_1670,N_1300,N_1149);
nand U1671 (N_1671,N_1035,N_1281);
and U1672 (N_1672,N_1356,N_1187);
or U1673 (N_1673,N_1417,N_1282);
or U1674 (N_1674,N_1478,N_1378);
nand U1675 (N_1675,N_1476,N_1120);
nor U1676 (N_1676,N_1258,N_1173);
and U1677 (N_1677,N_1232,N_1494);
xor U1678 (N_1678,N_1163,N_1328);
and U1679 (N_1679,N_1144,N_1130);
xnor U1680 (N_1680,N_1463,N_1439);
and U1681 (N_1681,N_1215,N_1075);
nand U1682 (N_1682,N_1142,N_1320);
and U1683 (N_1683,N_1010,N_1489);
nor U1684 (N_1684,N_1213,N_1008);
xnor U1685 (N_1685,N_1272,N_1366);
nand U1686 (N_1686,N_1322,N_1303);
and U1687 (N_1687,N_1307,N_1086);
nor U1688 (N_1688,N_1052,N_1312);
nand U1689 (N_1689,N_1064,N_1049);
nor U1690 (N_1690,N_1326,N_1113);
nand U1691 (N_1691,N_1443,N_1171);
nor U1692 (N_1692,N_1027,N_1277);
xnor U1693 (N_1693,N_1166,N_1053);
nand U1694 (N_1694,N_1264,N_1060);
xnor U1695 (N_1695,N_1458,N_1025);
xnor U1696 (N_1696,N_1045,N_1342);
xor U1697 (N_1697,N_1483,N_1234);
xnor U1698 (N_1698,N_1193,N_1298);
xor U1699 (N_1699,N_1488,N_1054);
nand U1700 (N_1700,N_1316,N_1432);
nand U1701 (N_1701,N_1100,N_1372);
or U1702 (N_1702,N_1151,N_1233);
or U1703 (N_1703,N_1159,N_1279);
and U1704 (N_1704,N_1301,N_1204);
and U1705 (N_1705,N_1167,N_1346);
xor U1706 (N_1706,N_1470,N_1371);
or U1707 (N_1707,N_1350,N_1013);
or U1708 (N_1708,N_1335,N_1102);
or U1709 (N_1709,N_1221,N_1201);
nand U1710 (N_1710,N_1192,N_1250);
and U1711 (N_1711,N_1331,N_1395);
xnor U1712 (N_1712,N_1210,N_1005);
or U1713 (N_1713,N_1132,N_1406);
nor U1714 (N_1714,N_1389,N_1441);
and U1715 (N_1715,N_1422,N_1036);
or U1716 (N_1716,N_1185,N_1014);
nand U1717 (N_1717,N_1408,N_1486);
nand U1718 (N_1718,N_1292,N_1236);
nor U1719 (N_1719,N_1160,N_1177);
nor U1720 (N_1720,N_1313,N_1033);
xnor U1721 (N_1721,N_1181,N_1169);
or U1722 (N_1722,N_1437,N_1440);
nor U1723 (N_1723,N_1016,N_1240);
xor U1724 (N_1724,N_1462,N_1047);
xnor U1725 (N_1725,N_1061,N_1133);
or U1726 (N_1726,N_1203,N_1094);
nand U1727 (N_1727,N_1098,N_1009);
nor U1728 (N_1728,N_1180,N_1139);
nand U1729 (N_1729,N_1370,N_1186);
nor U1730 (N_1730,N_1248,N_1308);
or U1731 (N_1731,N_1270,N_1464);
or U1732 (N_1732,N_1413,N_1121);
nand U1733 (N_1733,N_1436,N_1034);
and U1734 (N_1734,N_1032,N_1208);
nand U1735 (N_1735,N_1450,N_1305);
and U1736 (N_1736,N_1119,N_1161);
and U1737 (N_1737,N_1046,N_1115);
or U1738 (N_1738,N_1170,N_1430);
nand U1739 (N_1739,N_1477,N_1344);
and U1740 (N_1740,N_1457,N_1391);
and U1741 (N_1741,N_1297,N_1099);
xnor U1742 (N_1742,N_1004,N_1127);
and U1743 (N_1743,N_1175,N_1393);
nor U1744 (N_1744,N_1376,N_1480);
xnor U1745 (N_1745,N_1345,N_1024);
and U1746 (N_1746,N_1219,N_1152);
xor U1747 (N_1747,N_1493,N_1184);
or U1748 (N_1748,N_1117,N_1191);
and U1749 (N_1749,N_1028,N_1065);
and U1750 (N_1750,N_1242,N_1207);
nand U1751 (N_1751,N_1462,N_1378);
nand U1752 (N_1752,N_1427,N_1446);
nand U1753 (N_1753,N_1442,N_1276);
nor U1754 (N_1754,N_1269,N_1162);
nand U1755 (N_1755,N_1483,N_1241);
nand U1756 (N_1756,N_1272,N_1215);
or U1757 (N_1757,N_1339,N_1485);
and U1758 (N_1758,N_1154,N_1381);
xor U1759 (N_1759,N_1173,N_1223);
or U1760 (N_1760,N_1158,N_1257);
xor U1761 (N_1761,N_1228,N_1115);
or U1762 (N_1762,N_1124,N_1214);
xor U1763 (N_1763,N_1108,N_1441);
nor U1764 (N_1764,N_1494,N_1057);
or U1765 (N_1765,N_1137,N_1009);
or U1766 (N_1766,N_1426,N_1086);
nand U1767 (N_1767,N_1403,N_1112);
and U1768 (N_1768,N_1248,N_1142);
or U1769 (N_1769,N_1094,N_1271);
or U1770 (N_1770,N_1032,N_1254);
or U1771 (N_1771,N_1280,N_1208);
or U1772 (N_1772,N_1232,N_1103);
xor U1773 (N_1773,N_1297,N_1227);
xnor U1774 (N_1774,N_1169,N_1382);
xnor U1775 (N_1775,N_1216,N_1160);
nor U1776 (N_1776,N_1186,N_1176);
or U1777 (N_1777,N_1328,N_1307);
nor U1778 (N_1778,N_1088,N_1106);
xnor U1779 (N_1779,N_1024,N_1495);
nor U1780 (N_1780,N_1298,N_1072);
and U1781 (N_1781,N_1409,N_1462);
nand U1782 (N_1782,N_1275,N_1057);
and U1783 (N_1783,N_1059,N_1325);
nand U1784 (N_1784,N_1335,N_1186);
nand U1785 (N_1785,N_1425,N_1306);
or U1786 (N_1786,N_1062,N_1451);
and U1787 (N_1787,N_1170,N_1495);
nand U1788 (N_1788,N_1325,N_1307);
or U1789 (N_1789,N_1262,N_1437);
nor U1790 (N_1790,N_1373,N_1385);
nor U1791 (N_1791,N_1486,N_1077);
nor U1792 (N_1792,N_1336,N_1134);
nor U1793 (N_1793,N_1295,N_1139);
and U1794 (N_1794,N_1421,N_1370);
nand U1795 (N_1795,N_1499,N_1250);
xnor U1796 (N_1796,N_1141,N_1489);
and U1797 (N_1797,N_1259,N_1303);
nand U1798 (N_1798,N_1129,N_1204);
or U1799 (N_1799,N_1417,N_1378);
and U1800 (N_1800,N_1141,N_1086);
or U1801 (N_1801,N_1032,N_1316);
or U1802 (N_1802,N_1194,N_1377);
xor U1803 (N_1803,N_1287,N_1360);
nor U1804 (N_1804,N_1017,N_1147);
or U1805 (N_1805,N_1170,N_1475);
nor U1806 (N_1806,N_1288,N_1361);
and U1807 (N_1807,N_1183,N_1459);
nand U1808 (N_1808,N_1140,N_1480);
and U1809 (N_1809,N_1110,N_1198);
or U1810 (N_1810,N_1024,N_1251);
xor U1811 (N_1811,N_1381,N_1284);
nand U1812 (N_1812,N_1456,N_1273);
or U1813 (N_1813,N_1252,N_1355);
nand U1814 (N_1814,N_1425,N_1282);
xnor U1815 (N_1815,N_1392,N_1426);
and U1816 (N_1816,N_1284,N_1075);
xor U1817 (N_1817,N_1237,N_1027);
and U1818 (N_1818,N_1257,N_1284);
nor U1819 (N_1819,N_1376,N_1410);
and U1820 (N_1820,N_1083,N_1230);
and U1821 (N_1821,N_1376,N_1038);
nand U1822 (N_1822,N_1227,N_1005);
or U1823 (N_1823,N_1414,N_1363);
and U1824 (N_1824,N_1457,N_1328);
nand U1825 (N_1825,N_1241,N_1199);
xor U1826 (N_1826,N_1450,N_1036);
nand U1827 (N_1827,N_1210,N_1497);
nand U1828 (N_1828,N_1167,N_1446);
nand U1829 (N_1829,N_1021,N_1254);
xor U1830 (N_1830,N_1150,N_1092);
xor U1831 (N_1831,N_1030,N_1212);
or U1832 (N_1832,N_1378,N_1037);
or U1833 (N_1833,N_1058,N_1243);
nand U1834 (N_1834,N_1146,N_1043);
nand U1835 (N_1835,N_1005,N_1253);
and U1836 (N_1836,N_1124,N_1363);
or U1837 (N_1837,N_1319,N_1114);
nand U1838 (N_1838,N_1002,N_1366);
nor U1839 (N_1839,N_1497,N_1147);
or U1840 (N_1840,N_1457,N_1125);
nor U1841 (N_1841,N_1210,N_1077);
nor U1842 (N_1842,N_1204,N_1398);
nor U1843 (N_1843,N_1429,N_1425);
and U1844 (N_1844,N_1183,N_1185);
nor U1845 (N_1845,N_1119,N_1328);
nand U1846 (N_1846,N_1245,N_1377);
nor U1847 (N_1847,N_1111,N_1464);
xnor U1848 (N_1848,N_1359,N_1109);
or U1849 (N_1849,N_1136,N_1272);
nor U1850 (N_1850,N_1071,N_1324);
or U1851 (N_1851,N_1402,N_1288);
or U1852 (N_1852,N_1224,N_1288);
and U1853 (N_1853,N_1430,N_1192);
nand U1854 (N_1854,N_1183,N_1360);
or U1855 (N_1855,N_1287,N_1399);
or U1856 (N_1856,N_1409,N_1331);
or U1857 (N_1857,N_1418,N_1141);
xnor U1858 (N_1858,N_1447,N_1316);
xor U1859 (N_1859,N_1252,N_1216);
nor U1860 (N_1860,N_1312,N_1369);
or U1861 (N_1861,N_1131,N_1155);
or U1862 (N_1862,N_1042,N_1192);
nand U1863 (N_1863,N_1073,N_1321);
and U1864 (N_1864,N_1190,N_1155);
nand U1865 (N_1865,N_1306,N_1444);
xnor U1866 (N_1866,N_1057,N_1282);
and U1867 (N_1867,N_1068,N_1436);
nand U1868 (N_1868,N_1365,N_1175);
xor U1869 (N_1869,N_1435,N_1292);
nor U1870 (N_1870,N_1157,N_1352);
xnor U1871 (N_1871,N_1153,N_1480);
nand U1872 (N_1872,N_1100,N_1345);
nand U1873 (N_1873,N_1158,N_1347);
or U1874 (N_1874,N_1381,N_1397);
nor U1875 (N_1875,N_1344,N_1047);
xor U1876 (N_1876,N_1327,N_1254);
or U1877 (N_1877,N_1291,N_1447);
and U1878 (N_1878,N_1173,N_1211);
nand U1879 (N_1879,N_1192,N_1175);
and U1880 (N_1880,N_1425,N_1435);
xor U1881 (N_1881,N_1137,N_1055);
xor U1882 (N_1882,N_1085,N_1203);
and U1883 (N_1883,N_1008,N_1078);
or U1884 (N_1884,N_1273,N_1053);
and U1885 (N_1885,N_1358,N_1317);
nand U1886 (N_1886,N_1259,N_1130);
xnor U1887 (N_1887,N_1221,N_1175);
or U1888 (N_1888,N_1018,N_1202);
nand U1889 (N_1889,N_1038,N_1290);
nor U1890 (N_1890,N_1232,N_1019);
and U1891 (N_1891,N_1066,N_1416);
or U1892 (N_1892,N_1176,N_1090);
nor U1893 (N_1893,N_1077,N_1445);
and U1894 (N_1894,N_1424,N_1279);
nand U1895 (N_1895,N_1440,N_1275);
xnor U1896 (N_1896,N_1152,N_1012);
and U1897 (N_1897,N_1310,N_1153);
and U1898 (N_1898,N_1307,N_1221);
xnor U1899 (N_1899,N_1309,N_1402);
xnor U1900 (N_1900,N_1119,N_1138);
nand U1901 (N_1901,N_1201,N_1498);
or U1902 (N_1902,N_1272,N_1054);
nor U1903 (N_1903,N_1218,N_1024);
xor U1904 (N_1904,N_1307,N_1122);
and U1905 (N_1905,N_1312,N_1397);
nand U1906 (N_1906,N_1125,N_1365);
and U1907 (N_1907,N_1016,N_1091);
xnor U1908 (N_1908,N_1242,N_1460);
nor U1909 (N_1909,N_1197,N_1428);
and U1910 (N_1910,N_1272,N_1348);
nand U1911 (N_1911,N_1254,N_1065);
xnor U1912 (N_1912,N_1245,N_1127);
and U1913 (N_1913,N_1029,N_1020);
and U1914 (N_1914,N_1269,N_1390);
and U1915 (N_1915,N_1207,N_1043);
and U1916 (N_1916,N_1382,N_1189);
nand U1917 (N_1917,N_1125,N_1285);
nor U1918 (N_1918,N_1235,N_1220);
nand U1919 (N_1919,N_1081,N_1432);
or U1920 (N_1920,N_1109,N_1381);
nand U1921 (N_1921,N_1205,N_1066);
xor U1922 (N_1922,N_1444,N_1239);
nand U1923 (N_1923,N_1233,N_1384);
nor U1924 (N_1924,N_1056,N_1230);
nand U1925 (N_1925,N_1105,N_1283);
xnor U1926 (N_1926,N_1430,N_1358);
xnor U1927 (N_1927,N_1317,N_1385);
nand U1928 (N_1928,N_1023,N_1277);
nor U1929 (N_1929,N_1207,N_1354);
nand U1930 (N_1930,N_1433,N_1014);
nor U1931 (N_1931,N_1283,N_1033);
or U1932 (N_1932,N_1210,N_1141);
or U1933 (N_1933,N_1451,N_1310);
and U1934 (N_1934,N_1357,N_1389);
xor U1935 (N_1935,N_1031,N_1232);
xnor U1936 (N_1936,N_1068,N_1092);
and U1937 (N_1937,N_1201,N_1073);
nor U1938 (N_1938,N_1328,N_1079);
and U1939 (N_1939,N_1016,N_1097);
nor U1940 (N_1940,N_1178,N_1392);
nand U1941 (N_1941,N_1062,N_1226);
nor U1942 (N_1942,N_1136,N_1471);
xor U1943 (N_1943,N_1070,N_1340);
xnor U1944 (N_1944,N_1474,N_1476);
and U1945 (N_1945,N_1335,N_1292);
xor U1946 (N_1946,N_1072,N_1026);
and U1947 (N_1947,N_1012,N_1096);
or U1948 (N_1948,N_1464,N_1035);
nand U1949 (N_1949,N_1041,N_1140);
and U1950 (N_1950,N_1061,N_1066);
xnor U1951 (N_1951,N_1004,N_1307);
and U1952 (N_1952,N_1229,N_1126);
and U1953 (N_1953,N_1251,N_1165);
nor U1954 (N_1954,N_1140,N_1243);
nand U1955 (N_1955,N_1347,N_1017);
nor U1956 (N_1956,N_1360,N_1425);
and U1957 (N_1957,N_1250,N_1480);
xnor U1958 (N_1958,N_1463,N_1424);
or U1959 (N_1959,N_1468,N_1339);
nor U1960 (N_1960,N_1464,N_1452);
and U1961 (N_1961,N_1451,N_1296);
nand U1962 (N_1962,N_1377,N_1481);
or U1963 (N_1963,N_1423,N_1382);
xor U1964 (N_1964,N_1073,N_1384);
or U1965 (N_1965,N_1192,N_1124);
or U1966 (N_1966,N_1449,N_1209);
nand U1967 (N_1967,N_1036,N_1052);
xor U1968 (N_1968,N_1179,N_1362);
or U1969 (N_1969,N_1083,N_1255);
nand U1970 (N_1970,N_1014,N_1374);
nor U1971 (N_1971,N_1102,N_1174);
xor U1972 (N_1972,N_1311,N_1387);
or U1973 (N_1973,N_1431,N_1205);
xnor U1974 (N_1974,N_1146,N_1111);
and U1975 (N_1975,N_1217,N_1394);
and U1976 (N_1976,N_1091,N_1386);
and U1977 (N_1977,N_1080,N_1322);
nor U1978 (N_1978,N_1363,N_1411);
nor U1979 (N_1979,N_1260,N_1314);
and U1980 (N_1980,N_1129,N_1147);
xor U1981 (N_1981,N_1257,N_1385);
and U1982 (N_1982,N_1175,N_1088);
or U1983 (N_1983,N_1399,N_1006);
and U1984 (N_1984,N_1129,N_1109);
or U1985 (N_1985,N_1429,N_1178);
nand U1986 (N_1986,N_1174,N_1233);
or U1987 (N_1987,N_1316,N_1183);
or U1988 (N_1988,N_1127,N_1046);
xnor U1989 (N_1989,N_1232,N_1270);
xnor U1990 (N_1990,N_1185,N_1025);
nand U1991 (N_1991,N_1386,N_1380);
nor U1992 (N_1992,N_1071,N_1170);
nand U1993 (N_1993,N_1453,N_1330);
or U1994 (N_1994,N_1354,N_1106);
nor U1995 (N_1995,N_1296,N_1322);
or U1996 (N_1996,N_1026,N_1129);
nor U1997 (N_1997,N_1348,N_1342);
and U1998 (N_1998,N_1287,N_1067);
and U1999 (N_1999,N_1015,N_1028);
nand U2000 (N_2000,N_1637,N_1666);
nand U2001 (N_2001,N_1976,N_1567);
nor U2002 (N_2002,N_1574,N_1948);
nor U2003 (N_2003,N_1713,N_1578);
and U2004 (N_2004,N_1593,N_1876);
and U2005 (N_2005,N_1902,N_1670);
nand U2006 (N_2006,N_1965,N_1701);
nor U2007 (N_2007,N_1984,N_1907);
or U2008 (N_2008,N_1546,N_1805);
and U2009 (N_2009,N_1563,N_1904);
or U2010 (N_2010,N_1848,N_1630);
nor U2011 (N_2011,N_1814,N_1792);
xnor U2012 (N_2012,N_1505,N_1899);
or U2013 (N_2013,N_1828,N_1649);
nand U2014 (N_2014,N_1530,N_1872);
nor U2015 (N_2015,N_1524,N_1830);
xnor U2016 (N_2016,N_1529,N_1572);
and U2017 (N_2017,N_1536,N_1641);
nand U2018 (N_2018,N_1935,N_1757);
nor U2019 (N_2019,N_1929,N_1644);
nand U2020 (N_2020,N_1739,N_1879);
nor U2021 (N_2021,N_1681,N_1866);
nor U2022 (N_2022,N_1922,N_1581);
or U2023 (N_2023,N_1862,N_1527);
nor U2024 (N_2024,N_1895,N_1813);
xnor U2025 (N_2025,N_1843,N_1638);
or U2026 (N_2026,N_1588,N_1921);
or U2027 (N_2027,N_1610,N_1580);
nor U2028 (N_2028,N_1525,N_1779);
nor U2029 (N_2029,N_1963,N_1560);
xor U2030 (N_2030,N_1617,N_1582);
nand U2031 (N_2031,N_1806,N_1518);
and U2032 (N_2032,N_1770,N_1734);
nor U2033 (N_2033,N_1655,N_1717);
nand U2034 (N_2034,N_1869,N_1903);
nor U2035 (N_2035,N_1815,N_1503);
or U2036 (N_2036,N_1835,N_1928);
nor U2037 (N_2037,N_1595,N_1628);
nand U2038 (N_2038,N_1868,N_1554);
or U2039 (N_2039,N_1724,N_1817);
xor U2040 (N_2040,N_1931,N_1821);
xor U2041 (N_2041,N_1811,N_1614);
nand U2042 (N_2042,N_1715,N_1905);
nand U2043 (N_2043,N_1627,N_1732);
nor U2044 (N_2044,N_1592,N_1591);
nand U2045 (N_2045,N_1889,N_1620);
nor U2046 (N_2046,N_1647,N_1777);
nand U2047 (N_2047,N_1733,N_1771);
or U2048 (N_2048,N_1808,N_1744);
and U2049 (N_2049,N_1937,N_1776);
or U2050 (N_2050,N_1861,N_1601);
nor U2051 (N_2051,N_1507,N_1636);
or U2052 (N_2052,N_1690,N_1799);
and U2053 (N_2053,N_1616,N_1990);
nand U2054 (N_2054,N_1975,N_1542);
nand U2055 (N_2055,N_1962,N_1596);
or U2056 (N_2056,N_1716,N_1911);
nor U2057 (N_2057,N_1998,N_1726);
or U2058 (N_2058,N_1926,N_1521);
or U2059 (N_2059,N_1679,N_1762);
and U2060 (N_2060,N_1608,N_1668);
and U2061 (N_2061,N_1839,N_1634);
nor U2062 (N_2062,N_1730,N_1629);
xnor U2063 (N_2063,N_1740,N_1547);
nand U2064 (N_2064,N_1663,N_1988);
nor U2065 (N_2065,N_1852,N_1979);
or U2066 (N_2066,N_1781,N_1856);
and U2067 (N_2067,N_1896,N_1936);
and U2068 (N_2068,N_1619,N_1657);
nor U2069 (N_2069,N_1587,N_1515);
nor U2070 (N_2070,N_1583,N_1689);
and U2071 (N_2071,N_1892,N_1568);
xor U2072 (N_2072,N_1646,N_1800);
xnor U2073 (N_2073,N_1942,N_1873);
and U2074 (N_2074,N_1796,N_1709);
nor U2075 (N_2075,N_1841,N_1829);
or U2076 (N_2076,N_1812,N_1598);
nand U2077 (N_2077,N_1961,N_1842);
nor U2078 (N_2078,N_1924,N_1564);
nor U2079 (N_2079,N_1768,N_1901);
xnor U2080 (N_2080,N_1845,N_1803);
nand U2081 (N_2081,N_1957,N_1579);
or U2082 (N_2082,N_1923,N_1674);
xor U2083 (N_2083,N_1600,N_1971);
or U2084 (N_2084,N_1802,N_1658);
xor U2085 (N_2085,N_1985,N_1513);
or U2086 (N_2086,N_1898,N_1784);
or U2087 (N_2087,N_1589,N_1676);
nand U2088 (N_2088,N_1705,N_1913);
or U2089 (N_2089,N_1585,N_1718);
nand U2090 (N_2090,N_1712,N_1978);
nand U2091 (N_2091,N_1920,N_1544);
or U2092 (N_2092,N_1890,N_1840);
nor U2093 (N_2093,N_1767,N_1612);
or U2094 (N_2094,N_1682,N_1983);
nand U2095 (N_2095,N_1914,N_1720);
or U2096 (N_2096,N_1787,N_1838);
and U2097 (N_2097,N_1859,N_1523);
xnor U2098 (N_2098,N_1747,N_1837);
and U2099 (N_2099,N_1669,N_1539);
and U2100 (N_2100,N_1943,N_1946);
or U2101 (N_2101,N_1711,N_1827);
nand U2102 (N_2102,N_1754,N_1794);
and U2103 (N_2103,N_1695,N_1857);
and U2104 (N_2104,N_1750,N_1915);
and U2105 (N_2105,N_1611,N_1603);
or U2106 (N_2106,N_1789,N_1877);
nand U2107 (N_2107,N_1912,N_1995);
nand U2108 (N_2108,N_1742,N_1997);
nor U2109 (N_2109,N_1888,N_1729);
nor U2110 (N_2110,N_1570,N_1749);
xnor U2111 (N_2111,N_1652,N_1783);
or U2112 (N_2112,N_1508,N_1569);
and U2113 (N_2113,N_1916,N_1631);
nor U2114 (N_2114,N_1615,N_1633);
nor U2115 (N_2115,N_1751,N_1917);
or U2116 (N_2116,N_1675,N_1556);
or U2117 (N_2117,N_1645,N_1551);
nand U2118 (N_2118,N_1847,N_1906);
xnor U2119 (N_2119,N_1822,N_1723);
or U2120 (N_2120,N_1624,N_1999);
nor U2121 (N_2121,N_1584,N_1698);
or U2122 (N_2122,N_1894,N_1970);
and U2123 (N_2123,N_1502,N_1960);
nand U2124 (N_2124,N_1597,N_1565);
nor U2125 (N_2125,N_1782,N_1844);
nand U2126 (N_2126,N_1651,N_1989);
or U2127 (N_2127,N_1543,N_1826);
nor U2128 (N_2128,N_1662,N_1613);
and U2129 (N_2129,N_1793,N_1878);
and U2130 (N_2130,N_1531,N_1622);
or U2131 (N_2131,N_1553,N_1748);
or U2132 (N_2132,N_1552,N_1727);
or U2133 (N_2133,N_1558,N_1968);
and U2134 (N_2134,N_1953,N_1625);
nor U2135 (N_2135,N_1526,N_1540);
nor U2136 (N_2136,N_1606,N_1884);
and U2137 (N_2137,N_1632,N_1688);
nor U2138 (N_2138,N_1880,N_1927);
and U2139 (N_2139,N_1512,N_1846);
and U2140 (N_2140,N_1609,N_1667);
nand U2141 (N_2141,N_1501,N_1795);
and U2142 (N_2142,N_1656,N_1653);
or U2143 (N_2143,N_1506,N_1964);
nor U2144 (N_2144,N_1874,N_1939);
or U2145 (N_2145,N_1871,N_1764);
nand U2146 (N_2146,N_1678,N_1743);
nand U2147 (N_2147,N_1672,N_1714);
and U2148 (N_2148,N_1908,N_1725);
or U2149 (N_2149,N_1746,N_1825);
or U2150 (N_2150,N_1831,N_1532);
xor U2151 (N_2151,N_1900,N_1759);
nand U2152 (N_2152,N_1604,N_1893);
or U2153 (N_2153,N_1561,N_1575);
or U2154 (N_2154,N_1519,N_1548);
xnor U2155 (N_2155,N_1686,N_1954);
nor U2156 (N_2156,N_1664,N_1738);
xnor U2157 (N_2157,N_1977,N_1959);
and U2158 (N_2158,N_1791,N_1535);
xor U2159 (N_2159,N_1510,N_1685);
or U2160 (N_2160,N_1736,N_1973);
nor U2161 (N_2161,N_1760,N_1566);
or U2162 (N_2162,N_1755,N_1930);
xnor U2163 (N_2163,N_1801,N_1761);
or U2164 (N_2164,N_1680,N_1661);
xor U2165 (N_2165,N_1650,N_1981);
nand U2166 (N_2166,N_1993,N_1853);
xor U2167 (N_2167,N_1969,N_1721);
or U2168 (N_2168,N_1858,N_1867);
and U2169 (N_2169,N_1697,N_1819);
xor U2170 (N_2170,N_1778,N_1775);
or U2171 (N_2171,N_1504,N_1763);
and U2172 (N_2172,N_1780,N_1863);
nor U2173 (N_2173,N_1958,N_1735);
nor U2174 (N_2174,N_1991,N_1966);
nor U2175 (N_2175,N_1798,N_1882);
xnor U2176 (N_2176,N_1785,N_1992);
and U2177 (N_2177,N_1642,N_1511);
xnor U2178 (N_2178,N_1687,N_1618);
nor U2179 (N_2179,N_1623,N_1545);
and U2180 (N_2180,N_1648,N_1897);
nor U2181 (N_2181,N_1683,N_1945);
and U2182 (N_2182,N_1602,N_1941);
nor U2183 (N_2183,N_1952,N_1522);
and U2184 (N_2184,N_1691,N_1643);
xor U2185 (N_2185,N_1824,N_1797);
xor U2186 (N_2186,N_1707,N_1967);
xnor U2187 (N_2187,N_1708,N_1986);
nor U2188 (N_2188,N_1934,N_1944);
or U2189 (N_2189,N_1559,N_1719);
nor U2190 (N_2190,N_1883,N_1865);
or U2191 (N_2191,N_1639,N_1820);
xor U2192 (N_2192,N_1586,N_1854);
nor U2193 (N_2193,N_1537,N_1772);
and U2194 (N_2194,N_1753,N_1517);
or U2195 (N_2195,N_1520,N_1766);
and U2196 (N_2196,N_1832,N_1528);
nand U2197 (N_2197,N_1704,N_1710);
xnor U2198 (N_2198,N_1850,N_1509);
nand U2199 (N_2199,N_1816,N_1833);
xnor U2200 (N_2200,N_1980,N_1925);
nand U2201 (N_2201,N_1684,N_1982);
or U2202 (N_2202,N_1938,N_1919);
and U2203 (N_2203,N_1870,N_1550);
and U2204 (N_2204,N_1706,N_1809);
xnor U2205 (N_2205,N_1765,N_1702);
nand U2206 (N_2206,N_1541,N_1731);
nand U2207 (N_2207,N_1933,N_1594);
xnor U2208 (N_2208,N_1699,N_1660);
or U2209 (N_2209,N_1758,N_1790);
and U2210 (N_2210,N_1555,N_1500);
nor U2211 (N_2211,N_1956,N_1788);
and U2212 (N_2212,N_1804,N_1947);
nand U2213 (N_2213,N_1635,N_1786);
or U2214 (N_2214,N_1752,N_1576);
xnor U2215 (N_2215,N_1741,N_1640);
or U2216 (N_2216,N_1533,N_1703);
nand U2217 (N_2217,N_1972,N_1851);
xor U2218 (N_2218,N_1737,N_1855);
or U2219 (N_2219,N_1875,N_1756);
nand U2220 (N_2220,N_1955,N_1538);
xor U2221 (N_2221,N_1834,N_1951);
xor U2222 (N_2222,N_1864,N_1836);
and U2223 (N_2223,N_1692,N_1700);
nand U2224 (N_2224,N_1860,N_1810);
xor U2225 (N_2225,N_1849,N_1557);
xnor U2226 (N_2226,N_1696,N_1516);
nand U2227 (N_2227,N_1534,N_1549);
xnor U2228 (N_2228,N_1605,N_1693);
nand U2229 (N_2229,N_1886,N_1728);
or U2230 (N_2230,N_1818,N_1677);
nand U2231 (N_2231,N_1626,N_1773);
xor U2232 (N_2232,N_1774,N_1654);
xnor U2233 (N_2233,N_1909,N_1514);
xnor U2234 (N_2234,N_1823,N_1987);
or U2235 (N_2235,N_1885,N_1950);
nor U2236 (N_2236,N_1949,N_1974);
xor U2237 (N_2237,N_1745,N_1671);
nand U2238 (N_2238,N_1562,N_1918);
nor U2239 (N_2239,N_1571,N_1996);
nor U2240 (N_2240,N_1881,N_1673);
or U2241 (N_2241,N_1590,N_1573);
xor U2242 (N_2242,N_1577,N_1932);
nand U2243 (N_2243,N_1607,N_1807);
nor U2244 (N_2244,N_1887,N_1769);
and U2245 (N_2245,N_1910,N_1940);
nor U2246 (N_2246,N_1694,N_1599);
xnor U2247 (N_2247,N_1722,N_1659);
nor U2248 (N_2248,N_1994,N_1665);
nand U2249 (N_2249,N_1891,N_1621);
nand U2250 (N_2250,N_1577,N_1746);
xor U2251 (N_2251,N_1991,N_1807);
and U2252 (N_2252,N_1998,N_1879);
nand U2253 (N_2253,N_1712,N_1508);
nand U2254 (N_2254,N_1539,N_1597);
or U2255 (N_2255,N_1680,N_1967);
or U2256 (N_2256,N_1782,N_1860);
xnor U2257 (N_2257,N_1642,N_1841);
and U2258 (N_2258,N_1624,N_1793);
and U2259 (N_2259,N_1720,N_1837);
nand U2260 (N_2260,N_1541,N_1518);
nand U2261 (N_2261,N_1592,N_1501);
and U2262 (N_2262,N_1579,N_1615);
nand U2263 (N_2263,N_1734,N_1500);
and U2264 (N_2264,N_1718,N_1834);
nor U2265 (N_2265,N_1717,N_1951);
nor U2266 (N_2266,N_1808,N_1717);
or U2267 (N_2267,N_1565,N_1792);
xor U2268 (N_2268,N_1505,N_1682);
nor U2269 (N_2269,N_1587,N_1785);
xnor U2270 (N_2270,N_1929,N_1690);
and U2271 (N_2271,N_1896,N_1566);
xor U2272 (N_2272,N_1603,N_1702);
nand U2273 (N_2273,N_1789,N_1604);
and U2274 (N_2274,N_1501,N_1685);
or U2275 (N_2275,N_1716,N_1957);
xor U2276 (N_2276,N_1699,N_1976);
xor U2277 (N_2277,N_1580,N_1643);
nand U2278 (N_2278,N_1633,N_1973);
nand U2279 (N_2279,N_1888,N_1803);
nand U2280 (N_2280,N_1783,N_1584);
nor U2281 (N_2281,N_1704,N_1919);
xor U2282 (N_2282,N_1956,N_1531);
or U2283 (N_2283,N_1854,N_1760);
xor U2284 (N_2284,N_1687,N_1831);
xor U2285 (N_2285,N_1821,N_1928);
xnor U2286 (N_2286,N_1581,N_1958);
nor U2287 (N_2287,N_1884,N_1966);
and U2288 (N_2288,N_1521,N_1792);
and U2289 (N_2289,N_1932,N_1750);
and U2290 (N_2290,N_1883,N_1994);
nor U2291 (N_2291,N_1845,N_1899);
nor U2292 (N_2292,N_1590,N_1945);
nand U2293 (N_2293,N_1602,N_1785);
xnor U2294 (N_2294,N_1565,N_1534);
or U2295 (N_2295,N_1755,N_1866);
nor U2296 (N_2296,N_1847,N_1578);
nand U2297 (N_2297,N_1951,N_1981);
or U2298 (N_2298,N_1992,N_1520);
or U2299 (N_2299,N_1811,N_1781);
or U2300 (N_2300,N_1995,N_1990);
or U2301 (N_2301,N_1761,N_1522);
or U2302 (N_2302,N_1799,N_1866);
and U2303 (N_2303,N_1591,N_1547);
nand U2304 (N_2304,N_1516,N_1598);
nor U2305 (N_2305,N_1836,N_1571);
or U2306 (N_2306,N_1633,N_1533);
nand U2307 (N_2307,N_1973,N_1606);
xnor U2308 (N_2308,N_1968,N_1876);
nand U2309 (N_2309,N_1844,N_1820);
and U2310 (N_2310,N_1530,N_1615);
xnor U2311 (N_2311,N_1691,N_1623);
xnor U2312 (N_2312,N_1607,N_1564);
nor U2313 (N_2313,N_1581,N_1615);
and U2314 (N_2314,N_1821,N_1682);
nand U2315 (N_2315,N_1524,N_1561);
and U2316 (N_2316,N_1769,N_1537);
nor U2317 (N_2317,N_1657,N_1711);
xnor U2318 (N_2318,N_1582,N_1898);
and U2319 (N_2319,N_1624,N_1767);
or U2320 (N_2320,N_1925,N_1990);
nor U2321 (N_2321,N_1605,N_1766);
and U2322 (N_2322,N_1830,N_1512);
or U2323 (N_2323,N_1731,N_1745);
nor U2324 (N_2324,N_1892,N_1806);
nand U2325 (N_2325,N_1585,N_1824);
xor U2326 (N_2326,N_1913,N_1833);
nand U2327 (N_2327,N_1709,N_1810);
or U2328 (N_2328,N_1930,N_1913);
nor U2329 (N_2329,N_1982,N_1925);
nand U2330 (N_2330,N_1752,N_1554);
and U2331 (N_2331,N_1702,N_1596);
nor U2332 (N_2332,N_1707,N_1519);
nand U2333 (N_2333,N_1843,N_1974);
and U2334 (N_2334,N_1587,N_1791);
nand U2335 (N_2335,N_1603,N_1848);
xnor U2336 (N_2336,N_1674,N_1707);
xnor U2337 (N_2337,N_1842,N_1990);
nor U2338 (N_2338,N_1500,N_1960);
nor U2339 (N_2339,N_1568,N_1564);
and U2340 (N_2340,N_1601,N_1923);
xnor U2341 (N_2341,N_1557,N_1751);
xor U2342 (N_2342,N_1972,N_1959);
and U2343 (N_2343,N_1665,N_1575);
nor U2344 (N_2344,N_1530,N_1650);
nand U2345 (N_2345,N_1983,N_1931);
nor U2346 (N_2346,N_1638,N_1527);
xor U2347 (N_2347,N_1878,N_1520);
nand U2348 (N_2348,N_1901,N_1850);
nor U2349 (N_2349,N_1568,N_1577);
and U2350 (N_2350,N_1999,N_1758);
xor U2351 (N_2351,N_1874,N_1754);
xnor U2352 (N_2352,N_1825,N_1847);
xnor U2353 (N_2353,N_1935,N_1544);
nor U2354 (N_2354,N_1737,N_1928);
and U2355 (N_2355,N_1613,N_1503);
nor U2356 (N_2356,N_1835,N_1718);
nor U2357 (N_2357,N_1629,N_1887);
or U2358 (N_2358,N_1909,N_1522);
or U2359 (N_2359,N_1647,N_1970);
nor U2360 (N_2360,N_1605,N_1599);
nor U2361 (N_2361,N_1736,N_1551);
or U2362 (N_2362,N_1556,N_1930);
and U2363 (N_2363,N_1998,N_1674);
nand U2364 (N_2364,N_1613,N_1682);
nand U2365 (N_2365,N_1848,N_1740);
nand U2366 (N_2366,N_1500,N_1737);
and U2367 (N_2367,N_1508,N_1908);
nand U2368 (N_2368,N_1894,N_1986);
or U2369 (N_2369,N_1673,N_1571);
nor U2370 (N_2370,N_1664,N_1914);
nand U2371 (N_2371,N_1903,N_1762);
and U2372 (N_2372,N_1900,N_1630);
nor U2373 (N_2373,N_1808,N_1733);
nand U2374 (N_2374,N_1595,N_1835);
nor U2375 (N_2375,N_1804,N_1978);
and U2376 (N_2376,N_1780,N_1560);
xnor U2377 (N_2377,N_1697,N_1664);
and U2378 (N_2378,N_1915,N_1569);
and U2379 (N_2379,N_1501,N_1906);
and U2380 (N_2380,N_1612,N_1851);
and U2381 (N_2381,N_1622,N_1727);
nand U2382 (N_2382,N_1627,N_1686);
or U2383 (N_2383,N_1760,N_1961);
and U2384 (N_2384,N_1913,N_1542);
or U2385 (N_2385,N_1633,N_1502);
nand U2386 (N_2386,N_1792,N_1895);
and U2387 (N_2387,N_1913,N_1943);
nand U2388 (N_2388,N_1978,N_1888);
nand U2389 (N_2389,N_1504,N_1852);
nor U2390 (N_2390,N_1657,N_1732);
nand U2391 (N_2391,N_1687,N_1532);
or U2392 (N_2392,N_1530,N_1945);
nand U2393 (N_2393,N_1681,N_1885);
nor U2394 (N_2394,N_1962,N_1724);
nor U2395 (N_2395,N_1700,N_1610);
xnor U2396 (N_2396,N_1579,N_1681);
xor U2397 (N_2397,N_1714,N_1771);
nor U2398 (N_2398,N_1669,N_1963);
nand U2399 (N_2399,N_1737,N_1604);
nor U2400 (N_2400,N_1798,N_1569);
nor U2401 (N_2401,N_1635,N_1980);
and U2402 (N_2402,N_1517,N_1538);
or U2403 (N_2403,N_1589,N_1923);
nand U2404 (N_2404,N_1529,N_1975);
xor U2405 (N_2405,N_1517,N_1971);
nand U2406 (N_2406,N_1870,N_1850);
and U2407 (N_2407,N_1959,N_1777);
and U2408 (N_2408,N_1532,N_1883);
xnor U2409 (N_2409,N_1702,N_1534);
or U2410 (N_2410,N_1866,N_1978);
and U2411 (N_2411,N_1948,N_1629);
xnor U2412 (N_2412,N_1523,N_1769);
and U2413 (N_2413,N_1876,N_1825);
xor U2414 (N_2414,N_1916,N_1796);
and U2415 (N_2415,N_1987,N_1902);
and U2416 (N_2416,N_1818,N_1813);
nand U2417 (N_2417,N_1681,N_1687);
nor U2418 (N_2418,N_1525,N_1519);
nor U2419 (N_2419,N_1748,N_1732);
xnor U2420 (N_2420,N_1864,N_1640);
and U2421 (N_2421,N_1892,N_1931);
nor U2422 (N_2422,N_1594,N_1931);
xnor U2423 (N_2423,N_1787,N_1529);
and U2424 (N_2424,N_1538,N_1878);
nand U2425 (N_2425,N_1940,N_1992);
nor U2426 (N_2426,N_1699,N_1802);
or U2427 (N_2427,N_1553,N_1973);
nor U2428 (N_2428,N_1504,N_1762);
xnor U2429 (N_2429,N_1889,N_1903);
nand U2430 (N_2430,N_1588,N_1577);
and U2431 (N_2431,N_1904,N_1832);
or U2432 (N_2432,N_1950,N_1712);
xnor U2433 (N_2433,N_1517,N_1770);
nor U2434 (N_2434,N_1688,N_1805);
nor U2435 (N_2435,N_1934,N_1705);
or U2436 (N_2436,N_1865,N_1997);
nor U2437 (N_2437,N_1935,N_1616);
xor U2438 (N_2438,N_1567,N_1669);
or U2439 (N_2439,N_1964,N_1883);
or U2440 (N_2440,N_1715,N_1587);
or U2441 (N_2441,N_1704,N_1932);
or U2442 (N_2442,N_1768,N_1843);
xnor U2443 (N_2443,N_1649,N_1545);
nor U2444 (N_2444,N_1984,N_1972);
nor U2445 (N_2445,N_1583,N_1614);
nand U2446 (N_2446,N_1652,N_1872);
or U2447 (N_2447,N_1835,N_1596);
nand U2448 (N_2448,N_1524,N_1938);
xor U2449 (N_2449,N_1907,N_1599);
or U2450 (N_2450,N_1923,N_1847);
or U2451 (N_2451,N_1717,N_1866);
and U2452 (N_2452,N_1524,N_1688);
and U2453 (N_2453,N_1906,N_1694);
nand U2454 (N_2454,N_1711,N_1748);
nand U2455 (N_2455,N_1600,N_1617);
and U2456 (N_2456,N_1725,N_1514);
nand U2457 (N_2457,N_1967,N_1697);
nor U2458 (N_2458,N_1559,N_1604);
nand U2459 (N_2459,N_1907,N_1535);
xnor U2460 (N_2460,N_1815,N_1988);
and U2461 (N_2461,N_1981,N_1800);
xnor U2462 (N_2462,N_1883,N_1806);
and U2463 (N_2463,N_1658,N_1749);
xnor U2464 (N_2464,N_1619,N_1570);
nand U2465 (N_2465,N_1997,N_1922);
nor U2466 (N_2466,N_1642,N_1688);
xor U2467 (N_2467,N_1898,N_1709);
and U2468 (N_2468,N_1584,N_1933);
or U2469 (N_2469,N_1616,N_1785);
or U2470 (N_2470,N_1812,N_1813);
and U2471 (N_2471,N_1638,N_1522);
or U2472 (N_2472,N_1738,N_1856);
xor U2473 (N_2473,N_1743,N_1761);
or U2474 (N_2474,N_1560,N_1715);
nor U2475 (N_2475,N_1966,N_1982);
or U2476 (N_2476,N_1653,N_1543);
xor U2477 (N_2477,N_1555,N_1545);
xor U2478 (N_2478,N_1804,N_1502);
xor U2479 (N_2479,N_1743,N_1535);
nand U2480 (N_2480,N_1752,N_1522);
xnor U2481 (N_2481,N_1522,N_1735);
and U2482 (N_2482,N_1769,N_1760);
nor U2483 (N_2483,N_1617,N_1964);
nand U2484 (N_2484,N_1627,N_1577);
nand U2485 (N_2485,N_1824,N_1961);
nor U2486 (N_2486,N_1776,N_1798);
or U2487 (N_2487,N_1906,N_1833);
nor U2488 (N_2488,N_1736,N_1715);
or U2489 (N_2489,N_1526,N_1942);
nand U2490 (N_2490,N_1541,N_1776);
or U2491 (N_2491,N_1896,N_1549);
nor U2492 (N_2492,N_1770,N_1808);
or U2493 (N_2493,N_1901,N_1791);
xnor U2494 (N_2494,N_1834,N_1763);
nor U2495 (N_2495,N_1852,N_1795);
and U2496 (N_2496,N_1911,N_1977);
xor U2497 (N_2497,N_1879,N_1867);
nor U2498 (N_2498,N_1945,N_1772);
xnor U2499 (N_2499,N_1853,N_1878);
nor U2500 (N_2500,N_2423,N_2178);
nor U2501 (N_2501,N_2378,N_2375);
nor U2502 (N_2502,N_2055,N_2197);
and U2503 (N_2503,N_2456,N_2071);
or U2504 (N_2504,N_2437,N_2361);
or U2505 (N_2505,N_2426,N_2436);
and U2506 (N_2506,N_2447,N_2101);
or U2507 (N_2507,N_2179,N_2278);
nand U2508 (N_2508,N_2037,N_2255);
or U2509 (N_2509,N_2469,N_2427);
or U2510 (N_2510,N_2470,N_2247);
nor U2511 (N_2511,N_2339,N_2373);
and U2512 (N_2512,N_2085,N_2371);
and U2513 (N_2513,N_2160,N_2345);
and U2514 (N_2514,N_2200,N_2372);
or U2515 (N_2515,N_2177,N_2299);
xor U2516 (N_2516,N_2498,N_2098);
xnor U2517 (N_2517,N_2273,N_2430);
and U2518 (N_2518,N_2229,N_2496);
nand U2519 (N_2519,N_2390,N_2243);
nand U2520 (N_2520,N_2297,N_2306);
and U2521 (N_2521,N_2488,N_2047);
or U2522 (N_2522,N_2158,N_2333);
nor U2523 (N_2523,N_2418,N_2481);
and U2524 (N_2524,N_2164,N_2484);
nand U2525 (N_2525,N_2081,N_2352);
and U2526 (N_2526,N_2324,N_2052);
nor U2527 (N_2527,N_2076,N_2004);
and U2528 (N_2528,N_2425,N_2190);
nand U2529 (N_2529,N_2440,N_2281);
and U2530 (N_2530,N_2040,N_2277);
or U2531 (N_2531,N_2495,N_2079);
and U2532 (N_2532,N_2043,N_2143);
and U2533 (N_2533,N_2216,N_2261);
and U2534 (N_2534,N_2062,N_2473);
nand U2535 (N_2535,N_2414,N_2359);
or U2536 (N_2536,N_2051,N_2205);
nand U2537 (N_2537,N_2117,N_2235);
and U2538 (N_2538,N_2168,N_2432);
nand U2539 (N_2539,N_2335,N_2121);
nand U2540 (N_2540,N_2327,N_2018);
nor U2541 (N_2541,N_2446,N_2226);
and U2542 (N_2542,N_2492,N_2448);
nand U2543 (N_2543,N_2093,N_2035);
nand U2544 (N_2544,N_2321,N_2225);
and U2545 (N_2545,N_2242,N_2073);
nand U2546 (N_2546,N_2494,N_2467);
nand U2547 (N_2547,N_2312,N_2453);
nor U2548 (N_2548,N_2349,N_2258);
nor U2549 (N_2549,N_2465,N_2175);
nand U2550 (N_2550,N_2376,N_2106);
or U2551 (N_2551,N_2217,N_2387);
nand U2552 (N_2552,N_2296,N_2240);
nand U2553 (N_2553,N_2377,N_2162);
and U2554 (N_2554,N_2188,N_2320);
nand U2555 (N_2555,N_2254,N_2429);
nand U2556 (N_2556,N_2389,N_2183);
or U2557 (N_2557,N_2357,N_2346);
and U2558 (N_2558,N_2319,N_2186);
and U2559 (N_2559,N_2233,N_2248);
xor U2560 (N_2560,N_2410,N_2094);
nor U2561 (N_2561,N_2326,N_2443);
nor U2562 (N_2562,N_2238,N_2256);
and U2563 (N_2563,N_2066,N_2288);
xor U2564 (N_2564,N_2220,N_2356);
or U2565 (N_2565,N_2120,N_2141);
and U2566 (N_2566,N_2351,N_2218);
xnor U2567 (N_2567,N_2170,N_2274);
or U2568 (N_2568,N_2404,N_2185);
xor U2569 (N_2569,N_2148,N_2355);
nand U2570 (N_2570,N_2182,N_2207);
or U2571 (N_2571,N_2201,N_2097);
xnor U2572 (N_2572,N_2264,N_2123);
xnor U2573 (N_2573,N_2065,N_2084);
xor U2574 (N_2574,N_2336,N_2295);
xnor U2575 (N_2575,N_2080,N_2012);
xor U2576 (N_2576,N_2394,N_2290);
or U2577 (N_2577,N_2303,N_2228);
or U2578 (N_2578,N_2338,N_2060);
and U2579 (N_2579,N_2382,N_2452);
nand U2580 (N_2580,N_2455,N_2298);
nand U2581 (N_2581,N_2204,N_2330);
or U2582 (N_2582,N_2027,N_2034);
or U2583 (N_2583,N_2478,N_2195);
and U2584 (N_2584,N_2155,N_2310);
or U2585 (N_2585,N_2328,N_2102);
or U2586 (N_2586,N_2317,N_2476);
nand U2587 (N_2587,N_2294,N_2393);
xnor U2588 (N_2588,N_2116,N_2244);
and U2589 (N_2589,N_2156,N_2318);
nor U2590 (N_2590,N_2276,N_2139);
nor U2591 (N_2591,N_2161,N_2413);
nand U2592 (N_2592,N_2099,N_2189);
or U2593 (N_2593,N_2280,N_2347);
xor U2594 (N_2594,N_2301,N_2088);
nand U2595 (N_2595,N_2223,N_2114);
xor U2596 (N_2596,N_2285,N_2471);
nand U2597 (N_2597,N_2428,N_2454);
nand U2598 (N_2598,N_2165,N_2489);
or U2599 (N_2599,N_2323,N_2388);
nor U2600 (N_2600,N_2309,N_2030);
nor U2601 (N_2601,N_2344,N_2129);
nand U2602 (N_2602,N_2305,N_2096);
xnor U2603 (N_2603,N_2045,N_2462);
nor U2604 (N_2604,N_2077,N_2006);
nand U2605 (N_2605,N_2300,N_2210);
xor U2606 (N_2606,N_2013,N_2314);
and U2607 (N_2607,N_2209,N_2271);
nand U2608 (N_2608,N_2211,N_2472);
nor U2609 (N_2609,N_2458,N_2202);
and U2610 (N_2610,N_2486,N_2463);
and U2611 (N_2611,N_2016,N_2444);
nor U2612 (N_2612,N_2400,N_2251);
or U2613 (N_2613,N_2451,N_2268);
or U2614 (N_2614,N_2024,N_2491);
or U2615 (N_2615,N_2212,N_2022);
xor U2616 (N_2616,N_2343,N_2194);
nor U2617 (N_2617,N_2137,N_2151);
nand U2618 (N_2618,N_2107,N_2086);
nor U2619 (N_2619,N_2246,N_2125);
nand U2620 (N_2620,N_2459,N_2411);
nand U2621 (N_2621,N_2287,N_2293);
xor U2622 (N_2622,N_2399,N_2157);
nand U2623 (N_2623,N_2069,N_2493);
nand U2624 (N_2624,N_2142,N_2431);
xor U2625 (N_2625,N_2193,N_2070);
nand U2626 (N_2626,N_2227,N_2395);
and U2627 (N_2627,N_2083,N_2128);
or U2628 (N_2628,N_2224,N_2033);
xor U2629 (N_2629,N_2474,N_2480);
and U2630 (N_2630,N_2307,N_2017);
xnor U2631 (N_2631,N_2483,N_2442);
nand U2632 (N_2632,N_2457,N_2350);
and U2633 (N_2633,N_2245,N_2331);
xnor U2634 (N_2634,N_2213,N_2416);
or U2635 (N_2635,N_2239,N_2103);
nor U2636 (N_2636,N_2119,N_2449);
or U2637 (N_2637,N_2075,N_2265);
and U2638 (N_2638,N_2174,N_2325);
and U2639 (N_2639,N_2180,N_2020);
nand U2640 (N_2640,N_2417,N_2384);
nand U2641 (N_2641,N_2140,N_2074);
nor U2642 (N_2642,N_2360,N_2134);
or U2643 (N_2643,N_2398,N_2270);
nand U2644 (N_2644,N_2401,N_2001);
and U2645 (N_2645,N_2391,N_2154);
xnor U2646 (N_2646,N_2313,N_2068);
and U2647 (N_2647,N_2253,N_2214);
nor U2648 (N_2648,N_2215,N_2292);
or U2649 (N_2649,N_2445,N_2208);
nand U2650 (N_2650,N_2172,N_2259);
xor U2651 (N_2651,N_2072,N_2127);
or U2652 (N_2652,N_2438,N_2367);
and U2653 (N_2653,N_2039,N_2184);
or U2654 (N_2654,N_2147,N_2311);
nor U2655 (N_2655,N_2230,N_2424);
and U2656 (N_2656,N_2358,N_2435);
or U2657 (N_2657,N_2383,N_2386);
or U2658 (N_2658,N_2056,N_2064);
nor U2659 (N_2659,N_2362,N_2434);
nor U2660 (N_2660,N_2196,N_2135);
nor U2661 (N_2661,N_2421,N_2231);
nor U2662 (N_2662,N_2354,N_2028);
and U2663 (N_2663,N_2091,N_2025);
nor U2664 (N_2664,N_2136,N_2152);
xor U2665 (N_2665,N_2366,N_2053);
and U2666 (N_2666,N_2023,N_2031);
or U2667 (N_2667,N_2221,N_2460);
nor U2668 (N_2668,N_2192,N_2497);
or U2669 (N_2669,N_2029,N_2009);
and U2670 (N_2670,N_2181,N_2171);
or U2671 (N_2671,N_2420,N_2061);
xor U2672 (N_2672,N_2409,N_2499);
nand U2673 (N_2673,N_2237,N_2441);
and U2674 (N_2674,N_2021,N_2252);
nor U2675 (N_2675,N_2124,N_2402);
xnor U2676 (N_2676,N_2477,N_2450);
nor U2677 (N_2677,N_2109,N_2087);
xor U2678 (N_2678,N_2063,N_2092);
nor U2679 (N_2679,N_2041,N_2090);
xnor U2680 (N_2680,N_2032,N_2369);
nor U2681 (N_2681,N_2115,N_2104);
nor U2682 (N_2682,N_2167,N_2396);
and U2683 (N_2683,N_2010,N_2475);
nor U2684 (N_2684,N_2379,N_2187);
nand U2685 (N_2685,N_2342,N_2126);
and U2686 (N_2686,N_2219,N_2007);
nand U2687 (N_2687,N_2408,N_2433);
nand U2688 (N_2688,N_2365,N_2110);
nor U2689 (N_2689,N_2370,N_2487);
or U2690 (N_2690,N_2019,N_2132);
xnor U2691 (N_2691,N_2466,N_2003);
and U2692 (N_2692,N_2011,N_2406);
nor U2693 (N_2693,N_2163,N_2439);
or U2694 (N_2694,N_2415,N_2112);
nand U2695 (N_2695,N_2059,N_2348);
nand U2696 (N_2696,N_2464,N_2078);
nor U2697 (N_2697,N_2262,N_2008);
nor U2698 (N_2698,N_2304,N_2048);
or U2699 (N_2699,N_2340,N_2149);
nand U2700 (N_2700,N_2257,N_2315);
or U2701 (N_2701,N_2364,N_2236);
or U2702 (N_2702,N_2014,N_2422);
or U2703 (N_2703,N_2329,N_2169);
xnor U2704 (N_2704,N_2234,N_2067);
nor U2705 (N_2705,N_2302,N_2279);
and U2706 (N_2706,N_2392,N_2150);
or U2707 (N_2707,N_2269,N_2490);
or U2708 (N_2708,N_2130,N_2203);
nand U2709 (N_2709,N_2334,N_2289);
nor U2710 (N_2710,N_2206,N_2108);
or U2711 (N_2711,N_2241,N_2198);
and U2712 (N_2712,N_2046,N_2385);
nor U2713 (N_2713,N_2026,N_2267);
nand U2714 (N_2714,N_2353,N_2322);
and U2715 (N_2715,N_2468,N_2049);
nor U2716 (N_2716,N_2250,N_2222);
and U2717 (N_2717,N_2118,N_2005);
nand U2718 (N_2718,N_2479,N_2397);
nor U2719 (N_2719,N_2266,N_2100);
or U2720 (N_2720,N_2095,N_2332);
and U2721 (N_2721,N_2284,N_2461);
xor U2722 (N_2722,N_2000,N_2368);
and U2723 (N_2723,N_2363,N_2381);
nor U2724 (N_2724,N_2146,N_2419);
or U2725 (N_2725,N_2038,N_2485);
and U2726 (N_2726,N_2407,N_2002);
xor U2727 (N_2727,N_2036,N_2403);
xor U2728 (N_2728,N_2272,N_2166);
nand U2729 (N_2729,N_2405,N_2232);
and U2730 (N_2730,N_2113,N_2131);
and U2731 (N_2731,N_2050,N_2341);
nor U2732 (N_2732,N_2054,N_2144);
and U2733 (N_2733,N_2316,N_2412);
xor U2734 (N_2734,N_2058,N_2145);
nand U2735 (N_2735,N_2260,N_2286);
or U2736 (N_2736,N_2275,N_2138);
nor U2737 (N_2737,N_2282,N_2380);
and U2738 (N_2738,N_2176,N_2082);
nand U2739 (N_2739,N_2199,N_2263);
xor U2740 (N_2740,N_2374,N_2249);
nor U2741 (N_2741,N_2042,N_2133);
and U2742 (N_2742,N_2159,N_2191);
nand U2743 (N_2743,N_2111,N_2153);
nand U2744 (N_2744,N_2173,N_2482);
nand U2745 (N_2745,N_2089,N_2308);
or U2746 (N_2746,N_2057,N_2044);
or U2747 (N_2747,N_2105,N_2337);
xnor U2748 (N_2748,N_2122,N_2283);
nor U2749 (N_2749,N_2015,N_2291);
nand U2750 (N_2750,N_2158,N_2136);
xor U2751 (N_2751,N_2156,N_2404);
nor U2752 (N_2752,N_2119,N_2015);
or U2753 (N_2753,N_2090,N_2204);
and U2754 (N_2754,N_2152,N_2431);
nor U2755 (N_2755,N_2114,N_2267);
or U2756 (N_2756,N_2134,N_2297);
and U2757 (N_2757,N_2179,N_2001);
and U2758 (N_2758,N_2086,N_2412);
or U2759 (N_2759,N_2198,N_2144);
and U2760 (N_2760,N_2125,N_2466);
and U2761 (N_2761,N_2369,N_2205);
nor U2762 (N_2762,N_2177,N_2376);
or U2763 (N_2763,N_2258,N_2055);
and U2764 (N_2764,N_2230,N_2387);
nor U2765 (N_2765,N_2124,N_2186);
xnor U2766 (N_2766,N_2180,N_2346);
or U2767 (N_2767,N_2405,N_2106);
and U2768 (N_2768,N_2215,N_2494);
and U2769 (N_2769,N_2238,N_2082);
xor U2770 (N_2770,N_2397,N_2263);
nand U2771 (N_2771,N_2497,N_2167);
or U2772 (N_2772,N_2460,N_2127);
nor U2773 (N_2773,N_2497,N_2183);
nand U2774 (N_2774,N_2168,N_2213);
nand U2775 (N_2775,N_2391,N_2492);
xnor U2776 (N_2776,N_2329,N_2006);
or U2777 (N_2777,N_2214,N_2383);
nand U2778 (N_2778,N_2017,N_2451);
nand U2779 (N_2779,N_2449,N_2046);
xor U2780 (N_2780,N_2201,N_2214);
nand U2781 (N_2781,N_2103,N_2438);
and U2782 (N_2782,N_2272,N_2183);
nand U2783 (N_2783,N_2352,N_2393);
xnor U2784 (N_2784,N_2468,N_2204);
and U2785 (N_2785,N_2466,N_2228);
xnor U2786 (N_2786,N_2167,N_2071);
nand U2787 (N_2787,N_2315,N_2461);
nand U2788 (N_2788,N_2196,N_2021);
nor U2789 (N_2789,N_2414,N_2302);
nand U2790 (N_2790,N_2474,N_2410);
xnor U2791 (N_2791,N_2438,N_2124);
and U2792 (N_2792,N_2047,N_2371);
xor U2793 (N_2793,N_2223,N_2124);
or U2794 (N_2794,N_2081,N_2457);
nand U2795 (N_2795,N_2315,N_2327);
and U2796 (N_2796,N_2056,N_2051);
nand U2797 (N_2797,N_2052,N_2193);
xor U2798 (N_2798,N_2071,N_2340);
nand U2799 (N_2799,N_2445,N_2004);
or U2800 (N_2800,N_2391,N_2121);
or U2801 (N_2801,N_2090,N_2444);
and U2802 (N_2802,N_2181,N_2497);
nand U2803 (N_2803,N_2416,N_2313);
nor U2804 (N_2804,N_2112,N_2217);
or U2805 (N_2805,N_2119,N_2117);
nand U2806 (N_2806,N_2020,N_2279);
nor U2807 (N_2807,N_2424,N_2124);
nand U2808 (N_2808,N_2285,N_2457);
xor U2809 (N_2809,N_2031,N_2177);
xor U2810 (N_2810,N_2431,N_2002);
xnor U2811 (N_2811,N_2044,N_2281);
or U2812 (N_2812,N_2207,N_2081);
and U2813 (N_2813,N_2285,N_2472);
nor U2814 (N_2814,N_2158,N_2252);
xor U2815 (N_2815,N_2403,N_2226);
and U2816 (N_2816,N_2451,N_2465);
and U2817 (N_2817,N_2430,N_2459);
nor U2818 (N_2818,N_2270,N_2018);
or U2819 (N_2819,N_2461,N_2493);
xnor U2820 (N_2820,N_2386,N_2172);
or U2821 (N_2821,N_2313,N_2469);
nor U2822 (N_2822,N_2354,N_2365);
nand U2823 (N_2823,N_2363,N_2266);
and U2824 (N_2824,N_2444,N_2066);
and U2825 (N_2825,N_2173,N_2263);
nor U2826 (N_2826,N_2154,N_2258);
or U2827 (N_2827,N_2036,N_2155);
xnor U2828 (N_2828,N_2332,N_2067);
and U2829 (N_2829,N_2248,N_2134);
or U2830 (N_2830,N_2190,N_2334);
nor U2831 (N_2831,N_2399,N_2014);
nand U2832 (N_2832,N_2394,N_2087);
or U2833 (N_2833,N_2231,N_2427);
xor U2834 (N_2834,N_2087,N_2026);
nor U2835 (N_2835,N_2042,N_2491);
and U2836 (N_2836,N_2422,N_2446);
xnor U2837 (N_2837,N_2271,N_2354);
xor U2838 (N_2838,N_2065,N_2282);
and U2839 (N_2839,N_2392,N_2415);
nor U2840 (N_2840,N_2275,N_2001);
nor U2841 (N_2841,N_2452,N_2295);
nand U2842 (N_2842,N_2361,N_2462);
and U2843 (N_2843,N_2152,N_2155);
or U2844 (N_2844,N_2078,N_2297);
or U2845 (N_2845,N_2185,N_2109);
nor U2846 (N_2846,N_2420,N_2223);
nand U2847 (N_2847,N_2051,N_2490);
xor U2848 (N_2848,N_2288,N_2226);
and U2849 (N_2849,N_2220,N_2063);
and U2850 (N_2850,N_2366,N_2155);
nand U2851 (N_2851,N_2252,N_2324);
nand U2852 (N_2852,N_2370,N_2107);
nor U2853 (N_2853,N_2247,N_2442);
nand U2854 (N_2854,N_2369,N_2467);
xor U2855 (N_2855,N_2223,N_2033);
and U2856 (N_2856,N_2318,N_2018);
or U2857 (N_2857,N_2037,N_2220);
nor U2858 (N_2858,N_2126,N_2491);
nor U2859 (N_2859,N_2272,N_2211);
and U2860 (N_2860,N_2202,N_2188);
or U2861 (N_2861,N_2467,N_2034);
and U2862 (N_2862,N_2245,N_2420);
nand U2863 (N_2863,N_2140,N_2132);
xor U2864 (N_2864,N_2233,N_2231);
nor U2865 (N_2865,N_2060,N_2373);
and U2866 (N_2866,N_2464,N_2295);
nor U2867 (N_2867,N_2434,N_2257);
xor U2868 (N_2868,N_2240,N_2415);
and U2869 (N_2869,N_2087,N_2203);
nor U2870 (N_2870,N_2466,N_2386);
nand U2871 (N_2871,N_2205,N_2392);
nor U2872 (N_2872,N_2200,N_2439);
or U2873 (N_2873,N_2430,N_2012);
xor U2874 (N_2874,N_2323,N_2381);
or U2875 (N_2875,N_2105,N_2358);
and U2876 (N_2876,N_2491,N_2090);
nand U2877 (N_2877,N_2245,N_2377);
xor U2878 (N_2878,N_2136,N_2365);
and U2879 (N_2879,N_2038,N_2220);
xor U2880 (N_2880,N_2188,N_2000);
xnor U2881 (N_2881,N_2306,N_2154);
nor U2882 (N_2882,N_2279,N_2469);
or U2883 (N_2883,N_2416,N_2275);
nor U2884 (N_2884,N_2197,N_2207);
nor U2885 (N_2885,N_2079,N_2219);
nor U2886 (N_2886,N_2385,N_2308);
or U2887 (N_2887,N_2290,N_2474);
or U2888 (N_2888,N_2024,N_2224);
and U2889 (N_2889,N_2146,N_2156);
nor U2890 (N_2890,N_2354,N_2289);
nand U2891 (N_2891,N_2448,N_2144);
xnor U2892 (N_2892,N_2329,N_2101);
nor U2893 (N_2893,N_2418,N_2013);
nor U2894 (N_2894,N_2265,N_2415);
and U2895 (N_2895,N_2061,N_2451);
or U2896 (N_2896,N_2163,N_2203);
and U2897 (N_2897,N_2437,N_2176);
nor U2898 (N_2898,N_2424,N_2479);
nand U2899 (N_2899,N_2379,N_2302);
nor U2900 (N_2900,N_2146,N_2278);
xor U2901 (N_2901,N_2305,N_2339);
nor U2902 (N_2902,N_2150,N_2249);
or U2903 (N_2903,N_2012,N_2449);
nor U2904 (N_2904,N_2153,N_2478);
nand U2905 (N_2905,N_2380,N_2307);
and U2906 (N_2906,N_2114,N_2175);
nand U2907 (N_2907,N_2062,N_2259);
or U2908 (N_2908,N_2077,N_2124);
nor U2909 (N_2909,N_2395,N_2408);
nor U2910 (N_2910,N_2111,N_2389);
xor U2911 (N_2911,N_2404,N_2459);
xor U2912 (N_2912,N_2044,N_2047);
or U2913 (N_2913,N_2254,N_2146);
nor U2914 (N_2914,N_2016,N_2296);
nand U2915 (N_2915,N_2278,N_2238);
xnor U2916 (N_2916,N_2283,N_2479);
xor U2917 (N_2917,N_2407,N_2074);
xor U2918 (N_2918,N_2265,N_2076);
nor U2919 (N_2919,N_2289,N_2234);
and U2920 (N_2920,N_2203,N_2043);
xor U2921 (N_2921,N_2110,N_2147);
and U2922 (N_2922,N_2419,N_2180);
or U2923 (N_2923,N_2206,N_2006);
xor U2924 (N_2924,N_2366,N_2151);
and U2925 (N_2925,N_2427,N_2431);
nand U2926 (N_2926,N_2126,N_2403);
nor U2927 (N_2927,N_2429,N_2487);
xor U2928 (N_2928,N_2268,N_2124);
xor U2929 (N_2929,N_2214,N_2439);
xor U2930 (N_2930,N_2040,N_2394);
nor U2931 (N_2931,N_2379,N_2341);
and U2932 (N_2932,N_2062,N_2031);
nor U2933 (N_2933,N_2261,N_2442);
nor U2934 (N_2934,N_2003,N_2074);
nand U2935 (N_2935,N_2344,N_2493);
xor U2936 (N_2936,N_2230,N_2087);
and U2937 (N_2937,N_2222,N_2171);
or U2938 (N_2938,N_2383,N_2008);
nand U2939 (N_2939,N_2360,N_2226);
or U2940 (N_2940,N_2144,N_2291);
or U2941 (N_2941,N_2081,N_2169);
or U2942 (N_2942,N_2050,N_2381);
nand U2943 (N_2943,N_2176,N_2081);
and U2944 (N_2944,N_2298,N_2282);
or U2945 (N_2945,N_2371,N_2176);
and U2946 (N_2946,N_2348,N_2044);
or U2947 (N_2947,N_2372,N_2055);
or U2948 (N_2948,N_2002,N_2080);
xnor U2949 (N_2949,N_2395,N_2066);
xnor U2950 (N_2950,N_2165,N_2340);
or U2951 (N_2951,N_2198,N_2477);
or U2952 (N_2952,N_2003,N_2159);
nor U2953 (N_2953,N_2423,N_2186);
nand U2954 (N_2954,N_2373,N_2318);
and U2955 (N_2955,N_2470,N_2395);
xnor U2956 (N_2956,N_2097,N_2486);
xor U2957 (N_2957,N_2110,N_2334);
xor U2958 (N_2958,N_2232,N_2053);
nor U2959 (N_2959,N_2018,N_2421);
and U2960 (N_2960,N_2420,N_2375);
xor U2961 (N_2961,N_2237,N_2069);
nand U2962 (N_2962,N_2145,N_2316);
xor U2963 (N_2963,N_2139,N_2353);
nand U2964 (N_2964,N_2040,N_2331);
and U2965 (N_2965,N_2455,N_2374);
nor U2966 (N_2966,N_2341,N_2331);
or U2967 (N_2967,N_2380,N_2253);
nand U2968 (N_2968,N_2468,N_2061);
nand U2969 (N_2969,N_2032,N_2051);
or U2970 (N_2970,N_2470,N_2259);
nor U2971 (N_2971,N_2252,N_2153);
and U2972 (N_2972,N_2211,N_2413);
and U2973 (N_2973,N_2070,N_2448);
nor U2974 (N_2974,N_2372,N_2380);
or U2975 (N_2975,N_2418,N_2389);
or U2976 (N_2976,N_2493,N_2429);
xor U2977 (N_2977,N_2284,N_2424);
xnor U2978 (N_2978,N_2461,N_2458);
or U2979 (N_2979,N_2298,N_2131);
nand U2980 (N_2980,N_2443,N_2210);
nor U2981 (N_2981,N_2148,N_2210);
and U2982 (N_2982,N_2225,N_2214);
nor U2983 (N_2983,N_2044,N_2194);
or U2984 (N_2984,N_2241,N_2411);
nor U2985 (N_2985,N_2265,N_2159);
xnor U2986 (N_2986,N_2226,N_2216);
or U2987 (N_2987,N_2249,N_2446);
nor U2988 (N_2988,N_2224,N_2427);
and U2989 (N_2989,N_2377,N_2246);
nand U2990 (N_2990,N_2199,N_2012);
or U2991 (N_2991,N_2115,N_2217);
nor U2992 (N_2992,N_2329,N_2395);
nor U2993 (N_2993,N_2296,N_2129);
or U2994 (N_2994,N_2014,N_2060);
or U2995 (N_2995,N_2017,N_2032);
nand U2996 (N_2996,N_2056,N_2426);
and U2997 (N_2997,N_2163,N_2386);
nor U2998 (N_2998,N_2265,N_2166);
or U2999 (N_2999,N_2103,N_2480);
xnor U3000 (N_3000,N_2943,N_2941);
nor U3001 (N_3001,N_2779,N_2935);
or U3002 (N_3002,N_2755,N_2684);
nor U3003 (N_3003,N_2663,N_2853);
xnor U3004 (N_3004,N_2759,N_2963);
nand U3005 (N_3005,N_2511,N_2770);
or U3006 (N_3006,N_2714,N_2506);
or U3007 (N_3007,N_2629,N_2903);
or U3008 (N_3008,N_2665,N_2966);
nor U3009 (N_3009,N_2564,N_2682);
and U3010 (N_3010,N_2879,N_2653);
xnor U3011 (N_3011,N_2995,N_2842);
xnor U3012 (N_3012,N_2911,N_2525);
nand U3013 (N_3013,N_2891,N_2922);
and U3014 (N_3014,N_2570,N_2819);
nor U3015 (N_3015,N_2633,N_2860);
nor U3016 (N_3016,N_2672,N_2946);
and U3017 (N_3017,N_2915,N_2652);
or U3018 (N_3018,N_2863,N_2975);
xnor U3019 (N_3019,N_2613,N_2698);
or U3020 (N_3020,N_2658,N_2587);
nor U3021 (N_3021,N_2961,N_2523);
nor U3022 (N_3022,N_2909,N_2902);
nand U3023 (N_3023,N_2960,N_2777);
nand U3024 (N_3024,N_2548,N_2631);
nand U3025 (N_3025,N_2816,N_2542);
or U3026 (N_3026,N_2557,N_2515);
or U3027 (N_3027,N_2594,N_2917);
nand U3028 (N_3028,N_2888,N_2823);
and U3029 (N_3029,N_2827,N_2883);
nor U3030 (N_3030,N_2899,N_2924);
and U3031 (N_3031,N_2581,N_2651);
or U3032 (N_3032,N_2826,N_2711);
xor U3033 (N_3033,N_2710,N_2640);
and U3034 (N_3034,N_2723,N_2942);
xnor U3035 (N_3035,N_2618,N_2959);
xnor U3036 (N_3036,N_2781,N_2931);
or U3037 (N_3037,N_2691,N_2906);
xor U3038 (N_3038,N_2894,N_2654);
xnor U3039 (N_3039,N_2828,N_2969);
and U3040 (N_3040,N_2914,N_2592);
nand U3041 (N_3041,N_2739,N_2986);
or U3042 (N_3042,N_2921,N_2549);
or U3043 (N_3043,N_2799,N_2807);
nor U3044 (N_3044,N_2859,N_2765);
xnor U3045 (N_3045,N_2784,N_2747);
and U3046 (N_3046,N_2760,N_2604);
xor U3047 (N_3047,N_2718,N_2687);
or U3048 (N_3048,N_2940,N_2662);
and U3049 (N_3049,N_2937,N_2996);
and U3050 (N_3050,N_2553,N_2624);
xnor U3051 (N_3051,N_2639,N_2571);
xor U3052 (N_3052,N_2843,N_2870);
nor U3053 (N_3053,N_2708,N_2797);
or U3054 (N_3054,N_2666,N_2775);
and U3055 (N_3055,N_2670,N_2575);
or U3056 (N_3056,N_2637,N_2838);
nand U3057 (N_3057,N_2674,N_2527);
and U3058 (N_3058,N_2832,N_2988);
or U3059 (N_3059,N_2659,N_2928);
and U3060 (N_3060,N_2861,N_2840);
nand U3061 (N_3061,N_2586,N_2676);
and U3062 (N_3062,N_2808,N_2881);
nor U3063 (N_3063,N_2751,N_2599);
nand U3064 (N_3064,N_2641,N_2721);
and U3065 (N_3065,N_2905,N_2907);
xor U3066 (N_3066,N_2731,N_2820);
xor U3067 (N_3067,N_2611,N_2593);
nand U3068 (N_3068,N_2858,N_2869);
or U3069 (N_3069,N_2873,N_2688);
or U3070 (N_3070,N_2713,N_2788);
or U3071 (N_3071,N_2795,N_2709);
xor U3072 (N_3072,N_2715,N_2836);
xor U3073 (N_3073,N_2780,N_2528);
or U3074 (N_3074,N_2706,N_2885);
nor U3075 (N_3075,N_2978,N_2776);
or U3076 (N_3076,N_2763,N_2729);
nand U3077 (N_3077,N_2783,N_2648);
xor U3078 (N_3078,N_2675,N_2771);
or U3079 (N_3079,N_2690,N_2892);
nand U3080 (N_3080,N_2513,N_2806);
nand U3081 (N_3081,N_2981,N_2634);
nor U3082 (N_3082,N_2635,N_2973);
nor U3083 (N_3083,N_2952,N_2574);
xor U3084 (N_3084,N_2678,N_2768);
xnor U3085 (N_3085,N_2578,N_2868);
xnor U3086 (N_3086,N_2554,N_2502);
and U3087 (N_3087,N_2520,N_2603);
xor U3088 (N_3088,N_2612,N_2617);
nand U3089 (N_3089,N_2880,N_2530);
xor U3090 (N_3090,N_2556,N_2671);
nand U3091 (N_3091,N_2796,N_2737);
or U3092 (N_3092,N_2991,N_2749);
xnor U3093 (N_3093,N_2752,N_2947);
xnor U3094 (N_3094,N_2601,N_2539);
or U3095 (N_3095,N_2644,N_2839);
xnor U3096 (N_3096,N_2786,N_2529);
nand U3097 (N_3097,N_2569,N_2918);
xor U3098 (N_3098,N_2757,N_2583);
nor U3099 (N_3099,N_2753,N_2893);
nor U3100 (N_3100,N_2756,N_2865);
nand U3101 (N_3101,N_2913,N_2983);
or U3102 (N_3102,N_2916,N_2792);
and U3103 (N_3103,N_2730,N_2598);
nor U3104 (N_3104,N_2805,N_2887);
or U3105 (N_3105,N_2833,N_2512);
or U3106 (N_3106,N_2615,N_2831);
nand U3107 (N_3107,N_2636,N_2811);
or U3108 (N_3108,N_2532,N_2862);
nand U3109 (N_3109,N_2874,N_2908);
xor U3110 (N_3110,N_2814,N_2974);
xnor U3111 (N_3111,N_2545,N_2938);
nor U3112 (N_3112,N_2519,N_2734);
nor U3113 (N_3113,N_2616,N_2886);
or U3114 (N_3114,N_2817,N_2929);
xnor U3115 (N_3115,N_2979,N_2877);
xor U3116 (N_3116,N_2504,N_2769);
nand U3117 (N_3117,N_2650,N_2852);
nor U3118 (N_3118,N_2610,N_2681);
nor U3119 (N_3119,N_2793,N_2965);
nand U3120 (N_3120,N_2912,N_2898);
xor U3121 (N_3121,N_2626,N_2851);
or U3122 (N_3122,N_2534,N_2732);
nor U3123 (N_3123,N_2638,N_2725);
and U3124 (N_3124,N_2901,N_2761);
nor U3125 (N_3125,N_2584,N_2565);
nor U3126 (N_3126,N_2503,N_2660);
nor U3127 (N_3127,N_2772,N_2850);
xor U3128 (N_3128,N_2518,N_2701);
or U3129 (N_3129,N_2856,N_2726);
and U3130 (N_3130,N_2944,N_2716);
or U3131 (N_3131,N_2794,N_2778);
or U3132 (N_3132,N_2516,N_2589);
nor U3133 (N_3133,N_2632,N_2742);
xnor U3134 (N_3134,N_2945,N_2841);
nand U3135 (N_3135,N_2573,N_2926);
nor U3136 (N_3136,N_2727,N_2904);
nor U3137 (N_3137,N_2724,N_2750);
nand U3138 (N_3138,N_2910,N_2738);
and U3139 (N_3139,N_2668,N_2608);
xnor U3140 (N_3140,N_2538,N_2889);
and U3141 (N_3141,N_2773,N_2971);
and U3142 (N_3142,N_2667,N_2628);
nor U3143 (N_3143,N_2657,N_2700);
and U3144 (N_3144,N_2656,N_2607);
nor U3145 (N_3145,N_2623,N_2925);
and U3146 (N_3146,N_2704,N_2890);
nand U3147 (N_3147,N_2955,N_2782);
nand U3148 (N_3148,N_2736,N_2767);
xor U3149 (N_3149,N_2720,N_2577);
or U3150 (N_3150,N_2923,N_2696);
nand U3151 (N_3151,N_2576,N_2968);
nand U3152 (N_3152,N_2933,N_2719);
nor U3153 (N_3153,N_2596,N_2643);
and U3154 (N_3154,N_2649,N_2982);
or U3155 (N_3155,N_2977,N_2537);
or U3156 (N_3156,N_2697,N_2563);
and U3157 (N_3157,N_2789,N_2551);
nand U3158 (N_3158,N_2661,N_2544);
or U3159 (N_3159,N_2962,N_2785);
nand U3160 (N_3160,N_2787,N_2740);
and U3161 (N_3161,N_2543,N_2998);
xnor U3162 (N_3162,N_2804,N_2680);
or U3163 (N_3163,N_2882,N_2600);
xor U3164 (N_3164,N_2694,N_2733);
or U3165 (N_3165,N_2837,N_2997);
or U3166 (N_3166,N_2572,N_2762);
xor U3167 (N_3167,N_2625,N_2531);
and U3168 (N_3168,N_2830,N_2939);
nor U3169 (N_3169,N_2602,N_2932);
xnor U3170 (N_3170,N_2541,N_2872);
and U3171 (N_3171,N_2683,N_2812);
xnor U3172 (N_3172,N_2620,N_2895);
and U3173 (N_3173,N_2825,N_2866);
nand U3174 (N_3174,N_2989,N_2993);
xor U3175 (N_3175,N_2536,N_2510);
and U3176 (N_3176,N_2951,N_2835);
xor U3177 (N_3177,N_2844,N_2848);
or U3178 (N_3178,N_2845,N_2588);
nor U3179 (N_3179,N_2521,N_2864);
nor U3180 (N_3180,N_2994,N_2744);
nor U3181 (N_3181,N_2818,N_2619);
nand U3182 (N_3182,N_2976,N_2514);
and U3183 (N_3183,N_2758,N_2802);
nor U3184 (N_3184,N_2559,N_2790);
nand U3185 (N_3185,N_2707,N_2934);
and U3186 (N_3186,N_2535,N_2524);
and U3187 (N_3187,N_2582,N_2717);
xor U3188 (N_3188,N_2505,N_2500);
nor U3189 (N_3189,N_2614,N_2702);
xnor U3190 (N_3190,N_2927,N_2950);
and U3191 (N_3191,N_2930,N_2810);
nand U3192 (N_3192,N_2957,N_2590);
and U3193 (N_3193,N_2948,N_2689);
or U3194 (N_3194,N_2692,N_2878);
nand U3195 (N_3195,N_2655,N_2875);
or U3196 (N_3196,N_2936,N_2630);
and U3197 (N_3197,N_2800,N_2550);
nor U3198 (N_3198,N_2646,N_2897);
xor U3199 (N_3199,N_2669,N_2693);
nand U3200 (N_3200,N_2546,N_2958);
or U3201 (N_3201,N_2728,N_2900);
xnor U3202 (N_3202,N_2754,N_2642);
nand U3203 (N_3203,N_2561,N_2647);
or U3204 (N_3204,N_2555,N_2849);
nor U3205 (N_3205,N_2741,N_2972);
or U3206 (N_3206,N_2985,N_2722);
nand U3207 (N_3207,N_2507,N_2798);
nand U3208 (N_3208,N_2580,N_2547);
xnor U3209 (N_3209,N_2954,N_2956);
nor U3210 (N_3210,N_2829,N_2645);
xor U3211 (N_3211,N_2522,N_2774);
xor U3212 (N_3212,N_2664,N_2801);
nand U3213 (N_3213,N_2766,N_2597);
xnor U3214 (N_3214,N_2834,N_2552);
xnor U3215 (N_3215,N_2533,N_2705);
nand U3216 (N_3216,N_2813,N_2871);
and U3217 (N_3217,N_2920,N_2857);
nand U3218 (N_3218,N_2606,N_2867);
and U3219 (N_3219,N_2745,N_2846);
and U3220 (N_3220,N_2703,N_2896);
nand U3221 (N_3221,N_2560,N_2558);
nand U3222 (N_3222,N_2695,N_2677);
nor U3223 (N_3223,N_2679,N_2517);
and U3224 (N_3224,N_2568,N_2579);
nor U3225 (N_3225,N_2824,N_2953);
and U3226 (N_3226,N_2764,N_2990);
nand U3227 (N_3227,N_2855,N_2595);
xor U3228 (N_3228,N_2743,N_2999);
nor U3229 (N_3229,N_2746,N_2919);
or U3230 (N_3230,N_2992,N_2673);
nor U3231 (N_3231,N_2627,N_2876);
xnor U3232 (N_3232,N_2622,N_2949);
nand U3233 (N_3233,N_2822,N_2585);
nor U3234 (N_3234,N_2567,N_2854);
xor U3235 (N_3235,N_2847,N_2540);
nand U3236 (N_3236,N_2609,N_2699);
or U3237 (N_3237,N_2685,N_2712);
or U3238 (N_3238,N_2591,N_2884);
nor U3239 (N_3239,N_2967,N_2735);
and U3240 (N_3240,N_2803,N_2686);
nand U3241 (N_3241,N_2980,N_2809);
nand U3242 (N_3242,N_2970,N_2621);
or U3243 (N_3243,N_2526,N_2605);
xor U3244 (N_3244,N_2987,N_2508);
and U3245 (N_3245,N_2964,N_2748);
or U3246 (N_3246,N_2984,N_2791);
nor U3247 (N_3247,N_2821,N_2562);
xnor U3248 (N_3248,N_2566,N_2509);
xnor U3249 (N_3249,N_2501,N_2815);
xnor U3250 (N_3250,N_2925,N_2551);
and U3251 (N_3251,N_2738,N_2736);
nand U3252 (N_3252,N_2737,N_2500);
nor U3253 (N_3253,N_2605,N_2711);
and U3254 (N_3254,N_2547,N_2627);
xor U3255 (N_3255,N_2702,N_2722);
or U3256 (N_3256,N_2761,N_2667);
or U3257 (N_3257,N_2616,N_2599);
nand U3258 (N_3258,N_2673,N_2614);
nand U3259 (N_3259,N_2555,N_2816);
nor U3260 (N_3260,N_2791,N_2593);
nand U3261 (N_3261,N_2735,N_2639);
xnor U3262 (N_3262,N_2987,N_2863);
nor U3263 (N_3263,N_2922,N_2993);
and U3264 (N_3264,N_2725,N_2971);
nand U3265 (N_3265,N_2691,N_2586);
or U3266 (N_3266,N_2789,N_2655);
or U3267 (N_3267,N_2979,N_2974);
xnor U3268 (N_3268,N_2711,N_2563);
nand U3269 (N_3269,N_2805,N_2765);
and U3270 (N_3270,N_2970,N_2743);
and U3271 (N_3271,N_2623,N_2621);
or U3272 (N_3272,N_2667,N_2915);
xor U3273 (N_3273,N_2504,N_2515);
nand U3274 (N_3274,N_2914,N_2698);
and U3275 (N_3275,N_2749,N_2519);
nand U3276 (N_3276,N_2803,N_2976);
nand U3277 (N_3277,N_2855,N_2530);
nand U3278 (N_3278,N_2768,N_2780);
and U3279 (N_3279,N_2825,N_2742);
and U3280 (N_3280,N_2879,N_2582);
nand U3281 (N_3281,N_2597,N_2907);
nor U3282 (N_3282,N_2560,N_2960);
or U3283 (N_3283,N_2887,N_2673);
xnor U3284 (N_3284,N_2711,N_2951);
nor U3285 (N_3285,N_2819,N_2662);
nor U3286 (N_3286,N_2735,N_2624);
or U3287 (N_3287,N_2766,N_2995);
and U3288 (N_3288,N_2986,N_2747);
nor U3289 (N_3289,N_2803,N_2850);
nor U3290 (N_3290,N_2901,N_2944);
nand U3291 (N_3291,N_2959,N_2680);
or U3292 (N_3292,N_2704,N_2721);
nor U3293 (N_3293,N_2548,N_2972);
xnor U3294 (N_3294,N_2840,N_2991);
xor U3295 (N_3295,N_2845,N_2896);
nand U3296 (N_3296,N_2516,N_2876);
xnor U3297 (N_3297,N_2674,N_2788);
nor U3298 (N_3298,N_2998,N_2656);
nand U3299 (N_3299,N_2627,N_2614);
xor U3300 (N_3300,N_2724,N_2826);
xnor U3301 (N_3301,N_2565,N_2988);
nor U3302 (N_3302,N_2966,N_2710);
or U3303 (N_3303,N_2579,N_2678);
or U3304 (N_3304,N_2644,N_2842);
nand U3305 (N_3305,N_2676,N_2985);
nor U3306 (N_3306,N_2560,N_2660);
and U3307 (N_3307,N_2816,N_2926);
xnor U3308 (N_3308,N_2664,N_2835);
and U3309 (N_3309,N_2804,N_2507);
nor U3310 (N_3310,N_2842,N_2715);
xnor U3311 (N_3311,N_2772,N_2966);
xor U3312 (N_3312,N_2707,N_2834);
or U3313 (N_3313,N_2803,N_2936);
and U3314 (N_3314,N_2892,N_2744);
and U3315 (N_3315,N_2795,N_2502);
and U3316 (N_3316,N_2848,N_2531);
xor U3317 (N_3317,N_2926,N_2993);
xor U3318 (N_3318,N_2512,N_2855);
or U3319 (N_3319,N_2525,N_2575);
or U3320 (N_3320,N_2741,N_2904);
xor U3321 (N_3321,N_2866,N_2580);
nor U3322 (N_3322,N_2802,N_2591);
and U3323 (N_3323,N_2866,N_2508);
or U3324 (N_3324,N_2998,N_2712);
nand U3325 (N_3325,N_2900,N_2989);
and U3326 (N_3326,N_2774,N_2532);
xor U3327 (N_3327,N_2558,N_2620);
or U3328 (N_3328,N_2692,N_2854);
or U3329 (N_3329,N_2692,N_2546);
nor U3330 (N_3330,N_2949,N_2609);
or U3331 (N_3331,N_2728,N_2603);
xnor U3332 (N_3332,N_2561,N_2588);
or U3333 (N_3333,N_2896,N_2646);
and U3334 (N_3334,N_2651,N_2950);
xor U3335 (N_3335,N_2807,N_2572);
xor U3336 (N_3336,N_2625,N_2887);
and U3337 (N_3337,N_2663,N_2857);
and U3338 (N_3338,N_2918,N_2951);
or U3339 (N_3339,N_2781,N_2605);
nand U3340 (N_3340,N_2553,N_2636);
nand U3341 (N_3341,N_2676,N_2775);
and U3342 (N_3342,N_2633,N_2961);
nor U3343 (N_3343,N_2574,N_2583);
and U3344 (N_3344,N_2777,N_2801);
and U3345 (N_3345,N_2651,N_2763);
nor U3346 (N_3346,N_2792,N_2544);
and U3347 (N_3347,N_2990,N_2994);
and U3348 (N_3348,N_2554,N_2833);
and U3349 (N_3349,N_2741,N_2690);
or U3350 (N_3350,N_2727,N_2870);
nand U3351 (N_3351,N_2898,N_2529);
nor U3352 (N_3352,N_2526,N_2988);
or U3353 (N_3353,N_2967,N_2554);
or U3354 (N_3354,N_2961,N_2987);
or U3355 (N_3355,N_2716,N_2768);
or U3356 (N_3356,N_2624,N_2669);
and U3357 (N_3357,N_2581,N_2591);
nor U3358 (N_3358,N_2780,N_2589);
and U3359 (N_3359,N_2984,N_2944);
nand U3360 (N_3360,N_2780,N_2599);
nor U3361 (N_3361,N_2915,N_2965);
nor U3362 (N_3362,N_2687,N_2933);
nor U3363 (N_3363,N_2947,N_2650);
xor U3364 (N_3364,N_2601,N_2873);
nor U3365 (N_3365,N_2763,N_2832);
xor U3366 (N_3366,N_2774,N_2650);
and U3367 (N_3367,N_2570,N_2676);
or U3368 (N_3368,N_2892,N_2755);
and U3369 (N_3369,N_2608,N_2981);
xor U3370 (N_3370,N_2961,N_2630);
xnor U3371 (N_3371,N_2892,N_2990);
or U3372 (N_3372,N_2585,N_2707);
or U3373 (N_3373,N_2999,N_2706);
and U3374 (N_3374,N_2760,N_2906);
nor U3375 (N_3375,N_2905,N_2704);
nor U3376 (N_3376,N_2780,N_2502);
and U3377 (N_3377,N_2950,N_2514);
xnor U3378 (N_3378,N_2922,N_2520);
xor U3379 (N_3379,N_2934,N_2824);
nor U3380 (N_3380,N_2712,N_2654);
and U3381 (N_3381,N_2979,N_2579);
xnor U3382 (N_3382,N_2531,N_2855);
and U3383 (N_3383,N_2536,N_2801);
or U3384 (N_3384,N_2614,N_2666);
nor U3385 (N_3385,N_2877,N_2977);
and U3386 (N_3386,N_2985,N_2790);
xnor U3387 (N_3387,N_2852,N_2854);
nand U3388 (N_3388,N_2713,N_2699);
nand U3389 (N_3389,N_2699,N_2869);
nor U3390 (N_3390,N_2682,N_2833);
nand U3391 (N_3391,N_2836,N_2872);
nor U3392 (N_3392,N_2584,N_2890);
nand U3393 (N_3393,N_2779,N_2720);
xor U3394 (N_3394,N_2621,N_2915);
and U3395 (N_3395,N_2880,N_2765);
nand U3396 (N_3396,N_2515,N_2682);
xor U3397 (N_3397,N_2833,N_2980);
or U3398 (N_3398,N_2607,N_2856);
and U3399 (N_3399,N_2596,N_2893);
xnor U3400 (N_3400,N_2692,N_2681);
xor U3401 (N_3401,N_2934,N_2560);
nor U3402 (N_3402,N_2913,N_2865);
nor U3403 (N_3403,N_2789,N_2898);
or U3404 (N_3404,N_2847,N_2839);
or U3405 (N_3405,N_2576,N_2962);
or U3406 (N_3406,N_2575,N_2972);
or U3407 (N_3407,N_2879,N_2851);
or U3408 (N_3408,N_2555,N_2791);
nor U3409 (N_3409,N_2996,N_2596);
and U3410 (N_3410,N_2766,N_2596);
and U3411 (N_3411,N_2936,N_2642);
and U3412 (N_3412,N_2695,N_2675);
xnor U3413 (N_3413,N_2881,N_2642);
nand U3414 (N_3414,N_2947,N_2846);
xnor U3415 (N_3415,N_2973,N_2942);
nand U3416 (N_3416,N_2646,N_2975);
nand U3417 (N_3417,N_2903,N_2934);
nand U3418 (N_3418,N_2571,N_2703);
or U3419 (N_3419,N_2834,N_2699);
or U3420 (N_3420,N_2645,N_2986);
or U3421 (N_3421,N_2765,N_2981);
nand U3422 (N_3422,N_2834,N_2545);
nor U3423 (N_3423,N_2910,N_2600);
nand U3424 (N_3424,N_2598,N_2571);
nor U3425 (N_3425,N_2701,N_2647);
or U3426 (N_3426,N_2638,N_2570);
xnor U3427 (N_3427,N_2965,N_2541);
nand U3428 (N_3428,N_2773,N_2812);
or U3429 (N_3429,N_2606,N_2600);
and U3430 (N_3430,N_2969,N_2741);
nand U3431 (N_3431,N_2585,N_2579);
nor U3432 (N_3432,N_2503,N_2510);
or U3433 (N_3433,N_2513,N_2895);
and U3434 (N_3434,N_2634,N_2857);
nor U3435 (N_3435,N_2998,N_2851);
nand U3436 (N_3436,N_2979,N_2704);
and U3437 (N_3437,N_2792,N_2705);
or U3438 (N_3438,N_2832,N_2887);
and U3439 (N_3439,N_2796,N_2999);
nand U3440 (N_3440,N_2795,N_2747);
or U3441 (N_3441,N_2581,N_2674);
and U3442 (N_3442,N_2838,N_2771);
nor U3443 (N_3443,N_2623,N_2773);
xnor U3444 (N_3444,N_2759,N_2556);
or U3445 (N_3445,N_2936,N_2699);
and U3446 (N_3446,N_2647,N_2973);
xor U3447 (N_3447,N_2831,N_2855);
nand U3448 (N_3448,N_2986,N_2709);
and U3449 (N_3449,N_2763,N_2631);
or U3450 (N_3450,N_2516,N_2926);
or U3451 (N_3451,N_2795,N_2608);
nand U3452 (N_3452,N_2560,N_2616);
nor U3453 (N_3453,N_2592,N_2769);
nor U3454 (N_3454,N_2969,N_2943);
nand U3455 (N_3455,N_2719,N_2948);
nor U3456 (N_3456,N_2755,N_2932);
and U3457 (N_3457,N_2900,N_2867);
or U3458 (N_3458,N_2844,N_2974);
nand U3459 (N_3459,N_2743,N_2974);
and U3460 (N_3460,N_2783,N_2546);
and U3461 (N_3461,N_2749,N_2560);
xnor U3462 (N_3462,N_2582,N_2670);
nand U3463 (N_3463,N_2574,N_2736);
and U3464 (N_3464,N_2810,N_2888);
and U3465 (N_3465,N_2523,N_2686);
nand U3466 (N_3466,N_2509,N_2523);
and U3467 (N_3467,N_2555,N_2800);
or U3468 (N_3468,N_2844,N_2973);
nor U3469 (N_3469,N_2788,N_2980);
xor U3470 (N_3470,N_2665,N_2597);
xor U3471 (N_3471,N_2658,N_2642);
and U3472 (N_3472,N_2622,N_2872);
nor U3473 (N_3473,N_2634,N_2879);
or U3474 (N_3474,N_2829,N_2572);
nor U3475 (N_3475,N_2974,N_2876);
xnor U3476 (N_3476,N_2628,N_2961);
nand U3477 (N_3477,N_2915,N_2887);
xnor U3478 (N_3478,N_2939,N_2648);
nand U3479 (N_3479,N_2862,N_2604);
nand U3480 (N_3480,N_2862,N_2990);
xor U3481 (N_3481,N_2755,N_2503);
nor U3482 (N_3482,N_2588,N_2635);
and U3483 (N_3483,N_2898,N_2961);
nor U3484 (N_3484,N_2509,N_2758);
nand U3485 (N_3485,N_2932,N_2642);
nand U3486 (N_3486,N_2568,N_2654);
nor U3487 (N_3487,N_2954,N_2664);
or U3488 (N_3488,N_2856,N_2640);
and U3489 (N_3489,N_2707,N_2665);
or U3490 (N_3490,N_2614,N_2861);
xor U3491 (N_3491,N_2959,N_2842);
nand U3492 (N_3492,N_2830,N_2631);
xor U3493 (N_3493,N_2885,N_2979);
or U3494 (N_3494,N_2902,N_2896);
and U3495 (N_3495,N_2971,N_2844);
xnor U3496 (N_3496,N_2878,N_2671);
and U3497 (N_3497,N_2562,N_2916);
or U3498 (N_3498,N_2603,N_2562);
xnor U3499 (N_3499,N_2755,N_2694);
or U3500 (N_3500,N_3465,N_3112);
xnor U3501 (N_3501,N_3092,N_3481);
xnor U3502 (N_3502,N_3312,N_3137);
nand U3503 (N_3503,N_3439,N_3352);
nor U3504 (N_3504,N_3059,N_3080);
and U3505 (N_3505,N_3339,N_3159);
or U3506 (N_3506,N_3042,N_3030);
nor U3507 (N_3507,N_3102,N_3258);
or U3508 (N_3508,N_3161,N_3143);
nand U3509 (N_3509,N_3006,N_3195);
xnor U3510 (N_3510,N_3445,N_3153);
xnor U3511 (N_3511,N_3200,N_3387);
or U3512 (N_3512,N_3244,N_3437);
xnor U3513 (N_3513,N_3331,N_3118);
and U3514 (N_3514,N_3045,N_3093);
xor U3515 (N_3515,N_3271,N_3172);
or U3516 (N_3516,N_3182,N_3377);
xnor U3517 (N_3517,N_3127,N_3069);
or U3518 (N_3518,N_3193,N_3212);
nand U3519 (N_3519,N_3178,N_3084);
xnor U3520 (N_3520,N_3297,N_3255);
nor U3521 (N_3521,N_3061,N_3156);
and U3522 (N_3522,N_3241,N_3369);
nor U3523 (N_3523,N_3476,N_3317);
nand U3524 (N_3524,N_3236,N_3231);
and U3525 (N_3525,N_3348,N_3459);
xor U3526 (N_3526,N_3315,N_3417);
nand U3527 (N_3527,N_3014,N_3431);
xor U3528 (N_3528,N_3499,N_3247);
and U3529 (N_3529,N_3217,N_3456);
nand U3530 (N_3530,N_3229,N_3207);
xor U3531 (N_3531,N_3373,N_3254);
xor U3532 (N_3532,N_3467,N_3239);
nor U3533 (N_3533,N_3432,N_3211);
nor U3534 (N_3534,N_3380,N_3027);
and U3535 (N_3535,N_3349,N_3150);
and U3536 (N_3536,N_3337,N_3371);
and U3537 (N_3537,N_3085,N_3302);
xnor U3538 (N_3538,N_3443,N_3232);
xnor U3539 (N_3539,N_3206,N_3238);
and U3540 (N_3540,N_3145,N_3123);
and U3541 (N_3541,N_3363,N_3198);
xor U3542 (N_3542,N_3131,N_3062);
xnor U3543 (N_3543,N_3100,N_3497);
nor U3544 (N_3544,N_3215,N_3414);
and U3545 (N_3545,N_3350,N_3287);
and U3546 (N_3546,N_3097,N_3181);
nand U3547 (N_3547,N_3139,N_3026);
nor U3548 (N_3548,N_3205,N_3036);
nor U3549 (N_3549,N_3457,N_3032);
or U3550 (N_3550,N_3202,N_3233);
and U3551 (N_3551,N_3282,N_3372);
and U3552 (N_3552,N_3281,N_3398);
or U3553 (N_3553,N_3487,N_3356);
nand U3554 (N_3554,N_3473,N_3248);
xor U3555 (N_3555,N_3213,N_3051);
nor U3556 (N_3556,N_3025,N_3035);
xor U3557 (N_3557,N_3422,N_3055);
nand U3558 (N_3558,N_3291,N_3355);
and U3559 (N_3559,N_3306,N_3015);
or U3560 (N_3560,N_3031,N_3184);
or U3561 (N_3561,N_3223,N_3171);
nand U3562 (N_3562,N_3338,N_3053);
nor U3563 (N_3563,N_3319,N_3274);
xnor U3564 (N_3564,N_3068,N_3196);
xor U3565 (N_3565,N_3086,N_3276);
nand U3566 (N_3566,N_3109,N_3428);
and U3567 (N_3567,N_3107,N_3169);
and U3568 (N_3568,N_3225,N_3144);
nand U3569 (N_3569,N_3477,N_3469);
nor U3570 (N_3570,N_3191,N_3095);
xor U3571 (N_3571,N_3135,N_3288);
or U3572 (N_3572,N_3447,N_3440);
xnor U3573 (N_3573,N_3074,N_3484);
xor U3574 (N_3574,N_3448,N_3420);
or U3575 (N_3575,N_3050,N_3077);
nor U3576 (N_3576,N_3168,N_3383);
or U3577 (N_3577,N_3300,N_3021);
nor U3578 (N_3578,N_3266,N_3090);
xnor U3579 (N_3579,N_3256,N_3376);
and U3580 (N_3580,N_3115,N_3237);
xor U3581 (N_3581,N_3192,N_3220);
or U3582 (N_3582,N_3165,N_3267);
nand U3583 (N_3583,N_3048,N_3060);
nand U3584 (N_3584,N_3190,N_3265);
and U3585 (N_3585,N_3136,N_3179);
and U3586 (N_3586,N_3052,N_3429);
xnor U3587 (N_3587,N_3466,N_3088);
xnor U3588 (N_3588,N_3038,N_3240);
nand U3589 (N_3589,N_3000,N_3367);
or U3590 (N_3590,N_3341,N_3284);
nand U3591 (N_3591,N_3263,N_3275);
or U3592 (N_3592,N_3007,N_3158);
xnor U3593 (N_3593,N_3189,N_3455);
nor U3594 (N_3594,N_3351,N_3180);
xor U3595 (N_3595,N_3132,N_3146);
nor U3596 (N_3596,N_3289,N_3301);
xnor U3597 (N_3597,N_3299,N_3359);
xnor U3598 (N_3598,N_3264,N_3313);
nand U3599 (N_3599,N_3280,N_3416);
or U3600 (N_3600,N_3490,N_3029);
nor U3601 (N_3601,N_3012,N_3444);
xor U3602 (N_3602,N_3020,N_3468);
xnor U3603 (N_3603,N_3047,N_3452);
nand U3604 (N_3604,N_3460,N_3270);
and U3605 (N_3605,N_3470,N_3216);
nor U3606 (N_3606,N_3201,N_3333);
xnor U3607 (N_3607,N_3250,N_3126);
and U3608 (N_3608,N_3324,N_3483);
nand U3609 (N_3609,N_3292,N_3357);
nand U3610 (N_3610,N_3391,N_3122);
or U3611 (N_3611,N_3296,N_3413);
xor U3612 (N_3612,N_3408,N_3147);
or U3613 (N_3613,N_3407,N_3128);
nor U3614 (N_3614,N_3471,N_3480);
nor U3615 (N_3615,N_3187,N_3049);
nand U3616 (N_3616,N_3204,N_3218);
nand U3617 (N_3617,N_3498,N_3058);
or U3618 (N_3618,N_3024,N_3425);
or U3619 (N_3619,N_3261,N_3342);
xnor U3620 (N_3620,N_3041,N_3016);
and U3621 (N_3621,N_3234,N_3091);
xor U3622 (N_3622,N_3082,N_3485);
xnor U3623 (N_3623,N_3174,N_3170);
nor U3624 (N_3624,N_3116,N_3382);
or U3625 (N_3625,N_3017,N_3397);
nand U3626 (N_3626,N_3406,N_3396);
nand U3627 (N_3627,N_3110,N_3298);
xor U3628 (N_3628,N_3451,N_3489);
xnor U3629 (N_3629,N_3354,N_3257);
nor U3630 (N_3630,N_3305,N_3418);
nor U3631 (N_3631,N_3098,N_3273);
nor U3632 (N_3632,N_3423,N_3076);
nor U3633 (N_3633,N_3404,N_3384);
nor U3634 (N_3634,N_3405,N_3308);
and U3635 (N_3635,N_3286,N_3065);
nand U3636 (N_3636,N_3303,N_3002);
or U3637 (N_3637,N_3424,N_3221);
xnor U3638 (N_3638,N_3124,N_3430);
nor U3639 (N_3639,N_3072,N_3004);
or U3640 (N_3640,N_3323,N_3328);
and U3641 (N_3641,N_3493,N_3379);
nand U3642 (N_3642,N_3119,N_3375);
nor U3643 (N_3643,N_3415,N_3009);
nand U3644 (N_3644,N_3067,N_3117);
nor U3645 (N_3645,N_3311,N_3409);
nand U3646 (N_3646,N_3314,N_3295);
nor U3647 (N_3647,N_3152,N_3399);
or U3648 (N_3648,N_3013,N_3066);
nor U3649 (N_3649,N_3166,N_3491);
nand U3650 (N_3650,N_3160,N_3173);
and U3651 (N_3651,N_3113,N_3043);
nand U3652 (N_3652,N_3054,N_3458);
nand U3653 (N_3653,N_3370,N_3336);
nand U3654 (N_3654,N_3148,N_3344);
and U3655 (N_3655,N_3070,N_3268);
and U3656 (N_3656,N_3393,N_3495);
or U3657 (N_3657,N_3079,N_3157);
nor U3658 (N_3658,N_3134,N_3394);
xor U3659 (N_3659,N_3434,N_3304);
nor U3660 (N_3660,N_3108,N_3056);
nor U3661 (N_3661,N_3167,N_3378);
nand U3662 (N_3662,N_3343,N_3366);
or U3663 (N_3663,N_3120,N_3099);
xor U3664 (N_3664,N_3492,N_3463);
and U3665 (N_3665,N_3154,N_3441);
or U3666 (N_3666,N_3037,N_3253);
or U3667 (N_3667,N_3353,N_3246);
or U3668 (N_3668,N_3033,N_3329);
or U3669 (N_3669,N_3224,N_3475);
or U3670 (N_3670,N_3358,N_3129);
or U3671 (N_3671,N_3316,N_3245);
or U3672 (N_3672,N_3081,N_3094);
nand U3673 (N_3673,N_3039,N_3411);
or U3674 (N_3674,N_3389,N_3242);
or U3675 (N_3675,N_3326,N_3044);
nor U3676 (N_3676,N_3103,N_3163);
or U3677 (N_3677,N_3449,N_3096);
or U3678 (N_3678,N_3386,N_3005);
or U3679 (N_3679,N_3461,N_3175);
and U3680 (N_3680,N_3340,N_3488);
and U3681 (N_3681,N_3071,N_3421);
nand U3682 (N_3682,N_3309,N_3410);
and U3683 (N_3683,N_3034,N_3142);
xor U3684 (N_3684,N_3307,N_3426);
nand U3685 (N_3685,N_3496,N_3023);
or U3686 (N_3686,N_3140,N_3427);
and U3687 (N_3687,N_3381,N_3008);
and U3688 (N_3688,N_3111,N_3046);
or U3689 (N_3689,N_3330,N_3272);
xnor U3690 (N_3690,N_3310,N_3176);
xor U3691 (N_3691,N_3073,N_3374);
or U3692 (N_3692,N_3327,N_3199);
xor U3693 (N_3693,N_3210,N_3285);
and U3694 (N_3694,N_3228,N_3064);
nand U3695 (N_3695,N_3089,N_3482);
nor U3696 (N_3696,N_3362,N_3105);
and U3697 (N_3697,N_3262,N_3278);
or U3698 (N_3698,N_3320,N_3104);
nand U3699 (N_3699,N_3325,N_3486);
xor U3700 (N_3700,N_3269,N_3345);
nand U3701 (N_3701,N_3087,N_3040);
and U3702 (N_3702,N_3293,N_3474);
or U3703 (N_3703,N_3186,N_3260);
nand U3704 (N_3704,N_3332,N_3322);
or U3705 (N_3705,N_3235,N_3003);
xnor U3706 (N_3706,N_3318,N_3462);
nor U3707 (N_3707,N_3130,N_3395);
nor U3708 (N_3708,N_3436,N_3290);
nand U3709 (N_3709,N_3230,N_3114);
xor U3710 (N_3710,N_3412,N_3203);
or U3711 (N_3711,N_3197,N_3226);
or U3712 (N_3712,N_3209,N_3106);
nand U3713 (N_3713,N_3419,N_3361);
or U3714 (N_3714,N_3011,N_3346);
xor U3715 (N_3715,N_3001,N_3151);
or U3716 (N_3716,N_3075,N_3185);
xnor U3717 (N_3717,N_3249,N_3149);
and U3718 (N_3718,N_3010,N_3022);
nand U3719 (N_3719,N_3368,N_3222);
nor U3720 (N_3720,N_3464,N_3155);
xnor U3721 (N_3721,N_3121,N_3438);
or U3722 (N_3722,N_3259,N_3435);
nor U3723 (N_3723,N_3450,N_3433);
xor U3724 (N_3724,N_3446,N_3294);
xnor U3725 (N_3725,N_3365,N_3183);
xor U3726 (N_3726,N_3133,N_3188);
xor U3727 (N_3727,N_3019,N_3057);
nor U3728 (N_3728,N_3388,N_3472);
and U3729 (N_3729,N_3227,N_3219);
or U3730 (N_3730,N_3283,N_3385);
and U3731 (N_3731,N_3208,N_3279);
or U3732 (N_3732,N_3194,N_3141);
nand U3733 (N_3733,N_3125,N_3400);
nor U3734 (N_3734,N_3494,N_3162);
xnor U3735 (N_3735,N_3214,N_3138);
or U3736 (N_3736,N_3478,N_3252);
or U3737 (N_3737,N_3453,N_3018);
xnor U3738 (N_3738,N_3028,N_3083);
nand U3739 (N_3739,N_3334,N_3277);
xor U3740 (N_3740,N_3335,N_3360);
and U3741 (N_3741,N_3442,N_3401);
and U3742 (N_3742,N_3101,N_3390);
nand U3743 (N_3743,N_3063,N_3164);
xnor U3744 (N_3744,N_3392,N_3402);
and U3745 (N_3745,N_3251,N_3321);
and U3746 (N_3746,N_3347,N_3403);
or U3747 (N_3747,N_3243,N_3454);
nor U3748 (N_3748,N_3479,N_3078);
xnor U3749 (N_3749,N_3364,N_3177);
xor U3750 (N_3750,N_3495,N_3342);
nand U3751 (N_3751,N_3046,N_3323);
nand U3752 (N_3752,N_3139,N_3292);
nand U3753 (N_3753,N_3056,N_3421);
nand U3754 (N_3754,N_3141,N_3309);
and U3755 (N_3755,N_3118,N_3000);
nand U3756 (N_3756,N_3326,N_3323);
xor U3757 (N_3757,N_3063,N_3430);
nor U3758 (N_3758,N_3060,N_3305);
or U3759 (N_3759,N_3208,N_3374);
nor U3760 (N_3760,N_3494,N_3204);
xor U3761 (N_3761,N_3009,N_3320);
nor U3762 (N_3762,N_3084,N_3118);
nor U3763 (N_3763,N_3437,N_3125);
nand U3764 (N_3764,N_3071,N_3268);
nor U3765 (N_3765,N_3287,N_3354);
nor U3766 (N_3766,N_3419,N_3489);
xnor U3767 (N_3767,N_3065,N_3248);
or U3768 (N_3768,N_3394,N_3129);
xnor U3769 (N_3769,N_3377,N_3338);
nand U3770 (N_3770,N_3458,N_3180);
and U3771 (N_3771,N_3148,N_3472);
or U3772 (N_3772,N_3076,N_3029);
nor U3773 (N_3773,N_3294,N_3329);
nand U3774 (N_3774,N_3359,N_3085);
xnor U3775 (N_3775,N_3234,N_3228);
nand U3776 (N_3776,N_3460,N_3413);
or U3777 (N_3777,N_3329,N_3356);
or U3778 (N_3778,N_3143,N_3154);
and U3779 (N_3779,N_3408,N_3215);
nand U3780 (N_3780,N_3370,N_3337);
nand U3781 (N_3781,N_3286,N_3424);
or U3782 (N_3782,N_3097,N_3290);
or U3783 (N_3783,N_3406,N_3463);
nand U3784 (N_3784,N_3398,N_3121);
nor U3785 (N_3785,N_3397,N_3179);
nor U3786 (N_3786,N_3181,N_3176);
and U3787 (N_3787,N_3272,N_3374);
xor U3788 (N_3788,N_3056,N_3425);
and U3789 (N_3789,N_3234,N_3055);
or U3790 (N_3790,N_3320,N_3027);
or U3791 (N_3791,N_3384,N_3498);
and U3792 (N_3792,N_3448,N_3041);
or U3793 (N_3793,N_3129,N_3145);
xnor U3794 (N_3794,N_3412,N_3316);
xnor U3795 (N_3795,N_3336,N_3374);
and U3796 (N_3796,N_3239,N_3409);
or U3797 (N_3797,N_3148,N_3242);
or U3798 (N_3798,N_3199,N_3093);
xor U3799 (N_3799,N_3097,N_3420);
nor U3800 (N_3800,N_3358,N_3300);
or U3801 (N_3801,N_3188,N_3041);
or U3802 (N_3802,N_3314,N_3419);
nand U3803 (N_3803,N_3265,N_3187);
nand U3804 (N_3804,N_3180,N_3034);
or U3805 (N_3805,N_3139,N_3302);
nor U3806 (N_3806,N_3110,N_3199);
and U3807 (N_3807,N_3115,N_3270);
nand U3808 (N_3808,N_3153,N_3340);
nand U3809 (N_3809,N_3365,N_3103);
nor U3810 (N_3810,N_3470,N_3242);
xnor U3811 (N_3811,N_3161,N_3247);
nand U3812 (N_3812,N_3432,N_3302);
and U3813 (N_3813,N_3416,N_3224);
and U3814 (N_3814,N_3221,N_3239);
and U3815 (N_3815,N_3266,N_3208);
nor U3816 (N_3816,N_3104,N_3018);
or U3817 (N_3817,N_3471,N_3057);
nor U3818 (N_3818,N_3341,N_3331);
xor U3819 (N_3819,N_3115,N_3483);
or U3820 (N_3820,N_3215,N_3080);
nor U3821 (N_3821,N_3035,N_3480);
nand U3822 (N_3822,N_3349,N_3170);
nor U3823 (N_3823,N_3388,N_3211);
nor U3824 (N_3824,N_3221,N_3122);
nor U3825 (N_3825,N_3453,N_3310);
and U3826 (N_3826,N_3266,N_3262);
xor U3827 (N_3827,N_3450,N_3251);
and U3828 (N_3828,N_3495,N_3260);
nor U3829 (N_3829,N_3303,N_3312);
and U3830 (N_3830,N_3148,N_3160);
or U3831 (N_3831,N_3009,N_3036);
nand U3832 (N_3832,N_3015,N_3056);
xor U3833 (N_3833,N_3291,N_3311);
and U3834 (N_3834,N_3495,N_3450);
nor U3835 (N_3835,N_3013,N_3157);
nor U3836 (N_3836,N_3216,N_3172);
or U3837 (N_3837,N_3485,N_3355);
or U3838 (N_3838,N_3322,N_3232);
xor U3839 (N_3839,N_3004,N_3210);
nand U3840 (N_3840,N_3253,N_3186);
nand U3841 (N_3841,N_3092,N_3380);
or U3842 (N_3842,N_3425,N_3017);
xnor U3843 (N_3843,N_3378,N_3454);
and U3844 (N_3844,N_3198,N_3223);
nor U3845 (N_3845,N_3167,N_3411);
or U3846 (N_3846,N_3392,N_3433);
nor U3847 (N_3847,N_3492,N_3257);
nand U3848 (N_3848,N_3181,N_3378);
or U3849 (N_3849,N_3314,N_3206);
nor U3850 (N_3850,N_3057,N_3311);
nor U3851 (N_3851,N_3121,N_3260);
and U3852 (N_3852,N_3423,N_3093);
nand U3853 (N_3853,N_3100,N_3449);
xor U3854 (N_3854,N_3102,N_3345);
nor U3855 (N_3855,N_3287,N_3098);
and U3856 (N_3856,N_3460,N_3221);
xor U3857 (N_3857,N_3027,N_3004);
or U3858 (N_3858,N_3427,N_3232);
nand U3859 (N_3859,N_3223,N_3057);
nand U3860 (N_3860,N_3489,N_3452);
nand U3861 (N_3861,N_3065,N_3124);
xnor U3862 (N_3862,N_3249,N_3490);
and U3863 (N_3863,N_3463,N_3400);
nand U3864 (N_3864,N_3484,N_3267);
nand U3865 (N_3865,N_3092,N_3465);
nand U3866 (N_3866,N_3348,N_3458);
nand U3867 (N_3867,N_3274,N_3453);
xor U3868 (N_3868,N_3108,N_3306);
or U3869 (N_3869,N_3203,N_3249);
and U3870 (N_3870,N_3057,N_3491);
nand U3871 (N_3871,N_3101,N_3132);
xnor U3872 (N_3872,N_3130,N_3265);
or U3873 (N_3873,N_3139,N_3118);
nor U3874 (N_3874,N_3089,N_3470);
nor U3875 (N_3875,N_3266,N_3085);
nand U3876 (N_3876,N_3046,N_3010);
and U3877 (N_3877,N_3118,N_3218);
nand U3878 (N_3878,N_3399,N_3394);
xnor U3879 (N_3879,N_3199,N_3340);
or U3880 (N_3880,N_3438,N_3004);
nor U3881 (N_3881,N_3270,N_3447);
and U3882 (N_3882,N_3465,N_3413);
nand U3883 (N_3883,N_3350,N_3081);
xor U3884 (N_3884,N_3323,N_3411);
nand U3885 (N_3885,N_3158,N_3321);
or U3886 (N_3886,N_3321,N_3095);
xor U3887 (N_3887,N_3176,N_3263);
xor U3888 (N_3888,N_3366,N_3494);
xor U3889 (N_3889,N_3106,N_3332);
nand U3890 (N_3890,N_3465,N_3372);
and U3891 (N_3891,N_3300,N_3401);
nor U3892 (N_3892,N_3323,N_3192);
nor U3893 (N_3893,N_3364,N_3220);
nor U3894 (N_3894,N_3039,N_3478);
nor U3895 (N_3895,N_3459,N_3333);
or U3896 (N_3896,N_3053,N_3336);
xor U3897 (N_3897,N_3132,N_3364);
xor U3898 (N_3898,N_3475,N_3191);
xor U3899 (N_3899,N_3133,N_3169);
xor U3900 (N_3900,N_3003,N_3063);
xor U3901 (N_3901,N_3464,N_3094);
xor U3902 (N_3902,N_3469,N_3271);
or U3903 (N_3903,N_3344,N_3328);
nor U3904 (N_3904,N_3060,N_3273);
and U3905 (N_3905,N_3343,N_3141);
or U3906 (N_3906,N_3431,N_3280);
nand U3907 (N_3907,N_3270,N_3122);
or U3908 (N_3908,N_3297,N_3048);
xnor U3909 (N_3909,N_3251,N_3037);
and U3910 (N_3910,N_3015,N_3322);
nand U3911 (N_3911,N_3121,N_3227);
or U3912 (N_3912,N_3092,N_3062);
or U3913 (N_3913,N_3282,N_3206);
xor U3914 (N_3914,N_3065,N_3255);
nand U3915 (N_3915,N_3362,N_3274);
xnor U3916 (N_3916,N_3189,N_3239);
and U3917 (N_3917,N_3115,N_3472);
nand U3918 (N_3918,N_3459,N_3078);
or U3919 (N_3919,N_3011,N_3484);
nand U3920 (N_3920,N_3328,N_3229);
and U3921 (N_3921,N_3336,N_3319);
nand U3922 (N_3922,N_3157,N_3466);
or U3923 (N_3923,N_3107,N_3299);
and U3924 (N_3924,N_3215,N_3122);
nor U3925 (N_3925,N_3348,N_3086);
and U3926 (N_3926,N_3355,N_3116);
and U3927 (N_3927,N_3489,N_3186);
xor U3928 (N_3928,N_3493,N_3399);
or U3929 (N_3929,N_3137,N_3437);
xor U3930 (N_3930,N_3282,N_3462);
nor U3931 (N_3931,N_3294,N_3466);
xor U3932 (N_3932,N_3420,N_3237);
and U3933 (N_3933,N_3401,N_3250);
nor U3934 (N_3934,N_3467,N_3088);
xor U3935 (N_3935,N_3094,N_3449);
and U3936 (N_3936,N_3452,N_3279);
nor U3937 (N_3937,N_3291,N_3239);
nand U3938 (N_3938,N_3026,N_3138);
and U3939 (N_3939,N_3495,N_3285);
or U3940 (N_3940,N_3179,N_3409);
xnor U3941 (N_3941,N_3290,N_3177);
nand U3942 (N_3942,N_3034,N_3302);
nand U3943 (N_3943,N_3495,N_3119);
nand U3944 (N_3944,N_3266,N_3265);
and U3945 (N_3945,N_3166,N_3275);
or U3946 (N_3946,N_3212,N_3131);
and U3947 (N_3947,N_3371,N_3488);
or U3948 (N_3948,N_3286,N_3077);
nand U3949 (N_3949,N_3155,N_3220);
nor U3950 (N_3950,N_3059,N_3079);
xnor U3951 (N_3951,N_3457,N_3478);
and U3952 (N_3952,N_3411,N_3208);
xnor U3953 (N_3953,N_3368,N_3119);
nor U3954 (N_3954,N_3429,N_3290);
nand U3955 (N_3955,N_3135,N_3292);
nand U3956 (N_3956,N_3246,N_3251);
or U3957 (N_3957,N_3391,N_3409);
nor U3958 (N_3958,N_3440,N_3116);
or U3959 (N_3959,N_3030,N_3418);
and U3960 (N_3960,N_3320,N_3278);
xnor U3961 (N_3961,N_3000,N_3396);
xnor U3962 (N_3962,N_3237,N_3361);
nor U3963 (N_3963,N_3284,N_3285);
or U3964 (N_3964,N_3047,N_3233);
and U3965 (N_3965,N_3402,N_3298);
or U3966 (N_3966,N_3106,N_3396);
nand U3967 (N_3967,N_3357,N_3229);
and U3968 (N_3968,N_3308,N_3228);
nand U3969 (N_3969,N_3329,N_3425);
xor U3970 (N_3970,N_3124,N_3078);
nor U3971 (N_3971,N_3349,N_3075);
and U3972 (N_3972,N_3007,N_3137);
nor U3973 (N_3973,N_3098,N_3343);
and U3974 (N_3974,N_3040,N_3318);
or U3975 (N_3975,N_3387,N_3299);
or U3976 (N_3976,N_3094,N_3096);
xnor U3977 (N_3977,N_3387,N_3169);
or U3978 (N_3978,N_3156,N_3167);
xor U3979 (N_3979,N_3291,N_3317);
xor U3980 (N_3980,N_3211,N_3032);
nand U3981 (N_3981,N_3202,N_3061);
or U3982 (N_3982,N_3048,N_3351);
or U3983 (N_3983,N_3043,N_3445);
xor U3984 (N_3984,N_3228,N_3272);
nor U3985 (N_3985,N_3449,N_3182);
and U3986 (N_3986,N_3423,N_3103);
and U3987 (N_3987,N_3274,N_3433);
nand U3988 (N_3988,N_3491,N_3170);
xnor U3989 (N_3989,N_3496,N_3453);
xor U3990 (N_3990,N_3328,N_3381);
nor U3991 (N_3991,N_3326,N_3483);
or U3992 (N_3992,N_3499,N_3140);
and U3993 (N_3993,N_3233,N_3173);
xor U3994 (N_3994,N_3401,N_3341);
and U3995 (N_3995,N_3149,N_3267);
nor U3996 (N_3996,N_3287,N_3347);
and U3997 (N_3997,N_3018,N_3094);
xor U3998 (N_3998,N_3370,N_3212);
xor U3999 (N_3999,N_3258,N_3020);
nor U4000 (N_4000,N_3939,N_3629);
xor U4001 (N_4001,N_3616,N_3908);
nor U4002 (N_4002,N_3950,N_3678);
nor U4003 (N_4003,N_3749,N_3690);
or U4004 (N_4004,N_3539,N_3587);
nor U4005 (N_4005,N_3988,N_3788);
nand U4006 (N_4006,N_3958,N_3681);
nor U4007 (N_4007,N_3898,N_3660);
xor U4008 (N_4008,N_3849,N_3882);
and U4009 (N_4009,N_3918,N_3821);
nand U4010 (N_4010,N_3506,N_3633);
nor U4011 (N_4011,N_3568,N_3626);
nand U4012 (N_4012,N_3507,N_3881);
or U4013 (N_4013,N_3528,N_3500);
and U4014 (N_4014,N_3793,N_3770);
xor U4015 (N_4015,N_3566,N_3783);
or U4016 (N_4016,N_3724,N_3924);
and U4017 (N_4017,N_3533,N_3986);
and U4018 (N_4018,N_3916,N_3923);
or U4019 (N_4019,N_3598,N_3571);
and U4020 (N_4020,N_3864,N_3611);
or U4021 (N_4021,N_3930,N_3897);
nor U4022 (N_4022,N_3818,N_3708);
and U4023 (N_4023,N_3888,N_3730);
xor U4024 (N_4024,N_3985,N_3640);
nand U4025 (N_4025,N_3789,N_3805);
and U4026 (N_4026,N_3826,N_3917);
or U4027 (N_4027,N_3523,N_3512);
and U4028 (N_4028,N_3602,N_3767);
nor U4029 (N_4029,N_3734,N_3860);
xor U4030 (N_4030,N_3847,N_3997);
or U4031 (N_4031,N_3573,N_3871);
nand U4032 (N_4032,N_3763,N_3675);
nor U4033 (N_4033,N_3710,N_3713);
and U4034 (N_4034,N_3804,N_3764);
xor U4035 (N_4035,N_3746,N_3726);
nand U4036 (N_4036,N_3612,N_3685);
xor U4037 (N_4037,N_3813,N_3731);
nand U4038 (N_4038,N_3522,N_3578);
nor U4039 (N_4039,N_3559,N_3910);
nand U4040 (N_4040,N_3853,N_3830);
nor U4041 (N_4041,N_3527,N_3901);
and U4042 (N_4042,N_3778,N_3779);
nor U4043 (N_4043,N_3814,N_3927);
or U4044 (N_4044,N_3773,N_3891);
xor U4045 (N_4045,N_3874,N_3683);
nand U4046 (N_4046,N_3838,N_3504);
nand U4047 (N_4047,N_3782,N_3766);
or U4048 (N_4048,N_3628,N_3510);
nor U4049 (N_4049,N_3593,N_3739);
nor U4050 (N_4050,N_3791,N_3857);
or U4051 (N_4051,N_3514,N_3712);
nand U4052 (N_4052,N_3900,N_3801);
and U4053 (N_4053,N_3803,N_3666);
xor U4054 (N_4054,N_3702,N_3921);
nor U4055 (N_4055,N_3638,N_3876);
nand U4056 (N_4056,N_3544,N_3561);
and U4057 (N_4057,N_3785,N_3933);
and U4058 (N_4058,N_3603,N_3934);
xor U4059 (N_4059,N_3648,N_3639);
xor U4060 (N_4060,N_3757,N_3920);
and U4061 (N_4061,N_3862,N_3787);
xnor U4062 (N_4062,N_3831,N_3643);
nand U4063 (N_4063,N_3955,N_3592);
and U4064 (N_4064,N_3932,N_3896);
and U4065 (N_4065,N_3966,N_3905);
and U4066 (N_4066,N_3972,N_3756);
nand U4067 (N_4067,N_3546,N_3954);
xnor U4068 (N_4068,N_3542,N_3919);
nand U4069 (N_4069,N_3599,N_3925);
nand U4070 (N_4070,N_3961,N_3852);
or U4071 (N_4071,N_3517,N_3680);
or U4072 (N_4072,N_3790,N_3851);
nand U4073 (N_4073,N_3704,N_3875);
and U4074 (N_4074,N_3995,N_3984);
and U4075 (N_4075,N_3644,N_3859);
xor U4076 (N_4076,N_3637,N_3562);
xor U4077 (N_4077,N_3904,N_3740);
nor U4078 (N_4078,N_3569,N_3550);
or U4079 (N_4079,N_3635,N_3662);
or U4080 (N_4080,N_3677,N_3866);
or U4081 (N_4081,N_3722,N_3840);
xnor U4082 (N_4082,N_3736,N_3889);
nor U4083 (N_4083,N_3647,N_3590);
nor U4084 (N_4084,N_3846,N_3560);
or U4085 (N_4085,N_3953,N_3714);
xnor U4086 (N_4086,N_3880,N_3511);
nor U4087 (N_4087,N_3607,N_3907);
xor U4088 (N_4088,N_3516,N_3946);
xor U4089 (N_4089,N_3980,N_3537);
xor U4090 (N_4090,N_3794,N_3679);
or U4091 (N_4091,N_3753,N_3684);
nand U4092 (N_4092,N_3868,N_3776);
xor U4093 (N_4093,N_3665,N_3654);
nor U4094 (N_4094,N_3822,N_3604);
nand U4095 (N_4095,N_3941,N_3957);
nand U4096 (N_4096,N_3892,N_3886);
nor U4097 (N_4097,N_3890,N_3543);
or U4098 (N_4098,N_3692,N_3716);
and U4099 (N_4099,N_3858,N_3781);
and U4100 (N_4100,N_3548,N_3720);
nor U4101 (N_4101,N_3585,N_3777);
and U4102 (N_4102,N_3952,N_3557);
or U4103 (N_4103,N_3993,N_3747);
xnor U4104 (N_4104,N_3536,N_3855);
nand U4105 (N_4105,N_3622,N_3715);
nor U4106 (N_4106,N_3872,N_3613);
xnor U4107 (N_4107,N_3834,N_3700);
or U4108 (N_4108,N_3967,N_3661);
nand U4109 (N_4109,N_3620,N_3706);
xnor U4110 (N_4110,N_3646,N_3761);
nor U4111 (N_4111,N_3922,N_3832);
xnor U4112 (N_4112,N_3579,N_3623);
nor U4113 (N_4113,N_3558,N_3796);
xnor U4114 (N_4114,N_3589,N_3601);
and U4115 (N_4115,N_3944,N_3549);
nand U4116 (N_4116,N_3937,N_3828);
and U4117 (N_4117,N_3538,N_3733);
nor U4118 (N_4118,N_3540,N_3745);
nand U4119 (N_4119,N_3621,N_3656);
xnor U4120 (N_4120,N_3884,N_3564);
or U4121 (N_4121,N_3845,N_3689);
nand U4122 (N_4122,N_3664,N_3938);
and U4123 (N_4123,N_3636,N_3861);
and U4124 (N_4124,N_3948,N_3998);
nand U4125 (N_4125,N_3928,N_3951);
nand U4126 (N_4126,N_3624,N_3674);
xor U4127 (N_4127,N_3659,N_3554);
nand U4128 (N_4128,N_3987,N_3841);
nand U4129 (N_4129,N_3594,N_3615);
nand U4130 (N_4130,N_3574,N_3869);
xor U4131 (N_4131,N_3591,N_3863);
nor U4132 (N_4132,N_3608,N_3996);
and U4133 (N_4133,N_3619,N_3669);
and U4134 (N_4134,N_3772,N_3755);
and U4135 (N_4135,N_3727,N_3581);
and U4136 (N_4136,N_3645,N_3529);
and U4137 (N_4137,N_3798,N_3673);
or U4138 (N_4138,N_3978,N_3894);
nor U4139 (N_4139,N_3973,N_3837);
nand U4140 (N_4140,N_3505,N_3947);
or U4141 (N_4141,N_3563,N_3926);
or U4142 (N_4142,N_3989,N_3545);
xor U4143 (N_4143,N_3848,N_3617);
nor U4144 (N_4144,N_3784,N_3650);
xnor U4145 (N_4145,N_3600,N_3555);
xor U4146 (N_4146,N_3899,N_3525);
nand U4147 (N_4147,N_3509,N_3597);
xor U4148 (N_4148,N_3760,N_3502);
xor U4149 (N_4149,N_3632,N_3565);
and U4150 (N_4150,N_3748,N_3812);
nor U4151 (N_4151,N_3968,N_3931);
and U4152 (N_4152,N_3588,N_3976);
nor U4153 (N_4153,N_3771,N_3694);
nor U4154 (N_4154,N_3752,N_3780);
xor U4155 (N_4155,N_3945,N_3503);
xor U4156 (N_4156,N_3914,N_3839);
nor U4157 (N_4157,N_3797,N_3895);
nor U4158 (N_4158,N_3580,N_3663);
xnor U4159 (N_4159,N_3556,N_3833);
or U4160 (N_4160,N_3802,N_3721);
nor U4161 (N_4161,N_3641,N_3824);
xnor U4162 (N_4162,N_3906,N_3768);
xor U4163 (N_4163,N_3552,N_3974);
xor U4164 (N_4164,N_3728,N_3935);
and U4165 (N_4165,N_3586,N_3701);
nand U4166 (N_4166,N_3759,N_3775);
or U4167 (N_4167,N_3829,N_3835);
nor U4168 (N_4168,N_3657,N_3792);
or U4169 (N_4169,N_3651,N_3809);
nand U4170 (N_4170,N_3572,N_3810);
nor U4171 (N_4171,N_3642,N_3977);
and U4172 (N_4172,N_3668,N_3762);
xor U4173 (N_4173,N_3524,N_3795);
xor U4174 (N_4174,N_3703,N_3606);
xnor U4175 (N_4175,N_3634,N_3983);
or U4176 (N_4176,N_3960,N_3649);
and U4177 (N_4177,N_3738,N_3769);
or U4178 (N_4178,N_3725,N_3671);
or U4179 (N_4179,N_3965,N_3823);
xor U4180 (N_4180,N_3553,N_3723);
nor U4181 (N_4181,N_3531,N_3969);
xor U4182 (N_4182,N_3705,N_3820);
nand U4183 (N_4183,N_3742,N_3521);
nand U4184 (N_4184,N_3885,N_3691);
or U4185 (N_4185,N_3902,N_3686);
nand U4186 (N_4186,N_3991,N_3879);
xnor U4187 (N_4187,N_3915,N_3609);
nor U4188 (N_4188,N_3854,N_3843);
and U4189 (N_4189,N_3658,N_3867);
nand U4190 (N_4190,N_3670,N_3741);
xor U4191 (N_4191,N_3672,N_3584);
nand U4192 (N_4192,N_3750,N_3903);
and U4193 (N_4193,N_3631,N_3799);
nand U4194 (N_4194,N_3518,N_3732);
nand U4195 (N_4195,N_3825,N_3817);
nand U4196 (N_4196,N_3964,N_3975);
nor U4197 (N_4197,N_3695,N_3811);
nor U4198 (N_4198,N_3744,N_3719);
and U4199 (N_4199,N_3717,N_3567);
nand U4200 (N_4200,N_3614,N_3520);
and U4201 (N_4201,N_3743,N_3956);
xnor U4202 (N_4202,N_3981,N_3942);
xnor U4203 (N_4203,N_3519,N_3627);
and U4204 (N_4204,N_3711,N_3577);
nor U4205 (N_4205,N_3751,N_3815);
nand U4206 (N_4206,N_3735,N_3786);
and U4207 (N_4207,N_3990,N_3625);
or U4208 (N_4208,N_3844,N_3707);
nand U4209 (N_4209,N_3570,N_3541);
xnor U4210 (N_4210,N_3827,N_3576);
and U4211 (N_4211,N_3575,N_3909);
or U4212 (N_4212,N_3992,N_3929);
xor U4213 (N_4213,N_3501,N_3936);
nand U4214 (N_4214,N_3605,N_3819);
xor U4215 (N_4215,N_3963,N_3718);
or U4216 (N_4216,N_3696,N_3582);
nand U4217 (N_4217,N_3940,N_3532);
xor U4218 (N_4218,N_3729,N_3816);
xor U4219 (N_4219,N_3911,N_3682);
xnor U4220 (N_4220,N_3962,N_3667);
or U4221 (N_4221,N_3893,N_3508);
nor U4222 (N_4222,N_3971,N_3865);
nor U4223 (N_4223,N_3610,N_3535);
and U4224 (N_4224,N_3551,N_3547);
nand U4225 (N_4225,N_3530,N_3836);
xnor U4226 (N_4226,N_3515,N_3806);
xnor U4227 (N_4227,N_3583,N_3687);
or U4228 (N_4228,N_3883,N_3737);
nand U4229 (N_4229,N_3800,N_3970);
xnor U4230 (N_4230,N_3758,N_3887);
or U4231 (N_4231,N_3877,N_3842);
or U4232 (N_4232,N_3688,N_3698);
or U4233 (N_4233,N_3676,N_3913);
and U4234 (N_4234,N_3870,N_3912);
and U4235 (N_4235,N_3513,N_3754);
xor U4236 (N_4236,N_3807,N_3697);
nand U4237 (N_4237,N_3534,N_3709);
nand U4238 (N_4238,N_3873,N_3982);
or U4239 (N_4239,N_3774,N_3526);
nand U4240 (N_4240,N_3699,N_3959);
or U4241 (N_4241,N_3979,N_3850);
nor U4242 (N_4242,N_3999,N_3765);
or U4243 (N_4243,N_3595,N_3878);
nand U4244 (N_4244,N_3653,N_3808);
nor U4245 (N_4245,N_3943,N_3655);
nor U4246 (N_4246,N_3994,N_3618);
and U4247 (N_4247,N_3856,N_3630);
nor U4248 (N_4248,N_3949,N_3596);
and U4249 (N_4249,N_3652,N_3693);
xor U4250 (N_4250,N_3972,N_3598);
nor U4251 (N_4251,N_3871,N_3636);
and U4252 (N_4252,N_3716,N_3950);
and U4253 (N_4253,N_3797,N_3556);
nor U4254 (N_4254,N_3769,N_3794);
or U4255 (N_4255,N_3879,N_3888);
xnor U4256 (N_4256,N_3669,N_3690);
and U4257 (N_4257,N_3918,N_3561);
nand U4258 (N_4258,N_3571,N_3785);
and U4259 (N_4259,N_3807,N_3862);
or U4260 (N_4260,N_3824,N_3757);
and U4261 (N_4261,N_3906,N_3807);
nor U4262 (N_4262,N_3506,N_3776);
or U4263 (N_4263,N_3815,N_3588);
or U4264 (N_4264,N_3521,N_3605);
xnor U4265 (N_4265,N_3571,N_3721);
xnor U4266 (N_4266,N_3895,N_3949);
xnor U4267 (N_4267,N_3596,N_3837);
xnor U4268 (N_4268,N_3643,N_3905);
and U4269 (N_4269,N_3697,N_3524);
and U4270 (N_4270,N_3520,N_3610);
nand U4271 (N_4271,N_3799,N_3751);
xnor U4272 (N_4272,N_3620,N_3793);
nand U4273 (N_4273,N_3603,N_3930);
nand U4274 (N_4274,N_3714,N_3878);
or U4275 (N_4275,N_3740,N_3932);
and U4276 (N_4276,N_3867,N_3670);
xnor U4277 (N_4277,N_3884,N_3809);
xnor U4278 (N_4278,N_3520,N_3828);
or U4279 (N_4279,N_3501,N_3675);
and U4280 (N_4280,N_3707,N_3653);
nand U4281 (N_4281,N_3827,N_3630);
nand U4282 (N_4282,N_3722,N_3989);
nand U4283 (N_4283,N_3826,N_3775);
nand U4284 (N_4284,N_3876,N_3931);
nand U4285 (N_4285,N_3750,N_3684);
and U4286 (N_4286,N_3732,N_3799);
or U4287 (N_4287,N_3975,N_3578);
or U4288 (N_4288,N_3887,N_3895);
nor U4289 (N_4289,N_3919,N_3870);
xnor U4290 (N_4290,N_3891,N_3678);
xor U4291 (N_4291,N_3698,N_3885);
and U4292 (N_4292,N_3998,N_3719);
xnor U4293 (N_4293,N_3756,N_3606);
nand U4294 (N_4294,N_3986,N_3502);
xor U4295 (N_4295,N_3568,N_3563);
and U4296 (N_4296,N_3805,N_3874);
nand U4297 (N_4297,N_3531,N_3611);
nor U4298 (N_4298,N_3543,N_3538);
nand U4299 (N_4299,N_3667,N_3929);
and U4300 (N_4300,N_3744,N_3684);
nand U4301 (N_4301,N_3650,N_3539);
or U4302 (N_4302,N_3838,N_3908);
nor U4303 (N_4303,N_3521,N_3856);
and U4304 (N_4304,N_3814,N_3674);
nand U4305 (N_4305,N_3512,N_3670);
nand U4306 (N_4306,N_3820,N_3993);
nand U4307 (N_4307,N_3583,N_3924);
nand U4308 (N_4308,N_3686,N_3565);
xnor U4309 (N_4309,N_3561,N_3797);
and U4310 (N_4310,N_3710,N_3591);
nand U4311 (N_4311,N_3607,N_3504);
xnor U4312 (N_4312,N_3527,N_3969);
nor U4313 (N_4313,N_3791,N_3750);
nand U4314 (N_4314,N_3533,N_3594);
nor U4315 (N_4315,N_3531,N_3824);
and U4316 (N_4316,N_3627,N_3969);
nor U4317 (N_4317,N_3615,N_3628);
and U4318 (N_4318,N_3967,N_3509);
nand U4319 (N_4319,N_3533,N_3829);
xnor U4320 (N_4320,N_3598,N_3674);
xor U4321 (N_4321,N_3519,N_3536);
nand U4322 (N_4322,N_3714,N_3601);
or U4323 (N_4323,N_3951,N_3755);
nor U4324 (N_4324,N_3595,N_3572);
and U4325 (N_4325,N_3561,N_3781);
and U4326 (N_4326,N_3580,N_3679);
or U4327 (N_4327,N_3626,N_3690);
and U4328 (N_4328,N_3957,N_3933);
xnor U4329 (N_4329,N_3864,N_3709);
and U4330 (N_4330,N_3919,N_3831);
or U4331 (N_4331,N_3515,N_3766);
xnor U4332 (N_4332,N_3755,N_3785);
xor U4333 (N_4333,N_3793,N_3802);
nor U4334 (N_4334,N_3513,N_3849);
and U4335 (N_4335,N_3858,N_3607);
nor U4336 (N_4336,N_3765,N_3997);
nor U4337 (N_4337,N_3879,N_3526);
or U4338 (N_4338,N_3908,N_3612);
and U4339 (N_4339,N_3795,N_3518);
nand U4340 (N_4340,N_3726,N_3722);
and U4341 (N_4341,N_3710,N_3947);
or U4342 (N_4342,N_3681,N_3835);
nor U4343 (N_4343,N_3861,N_3522);
and U4344 (N_4344,N_3528,N_3572);
xor U4345 (N_4345,N_3583,N_3657);
nand U4346 (N_4346,N_3619,N_3798);
and U4347 (N_4347,N_3991,N_3869);
nor U4348 (N_4348,N_3739,N_3810);
and U4349 (N_4349,N_3984,N_3660);
or U4350 (N_4350,N_3509,N_3637);
and U4351 (N_4351,N_3955,N_3919);
nor U4352 (N_4352,N_3567,N_3500);
xor U4353 (N_4353,N_3552,N_3575);
and U4354 (N_4354,N_3702,N_3931);
and U4355 (N_4355,N_3575,N_3661);
nand U4356 (N_4356,N_3648,N_3963);
nand U4357 (N_4357,N_3685,N_3564);
or U4358 (N_4358,N_3508,N_3694);
xnor U4359 (N_4359,N_3773,N_3642);
nand U4360 (N_4360,N_3929,N_3750);
nor U4361 (N_4361,N_3574,N_3839);
or U4362 (N_4362,N_3846,N_3576);
and U4363 (N_4363,N_3695,N_3787);
and U4364 (N_4364,N_3715,N_3882);
xnor U4365 (N_4365,N_3685,N_3871);
nor U4366 (N_4366,N_3693,N_3833);
nand U4367 (N_4367,N_3612,N_3620);
nand U4368 (N_4368,N_3518,N_3828);
nor U4369 (N_4369,N_3530,N_3834);
nor U4370 (N_4370,N_3993,N_3642);
nand U4371 (N_4371,N_3956,N_3981);
xor U4372 (N_4372,N_3707,N_3532);
xnor U4373 (N_4373,N_3508,N_3838);
xor U4374 (N_4374,N_3932,N_3769);
nor U4375 (N_4375,N_3776,N_3869);
or U4376 (N_4376,N_3633,N_3972);
nor U4377 (N_4377,N_3894,N_3682);
or U4378 (N_4378,N_3658,N_3852);
nand U4379 (N_4379,N_3760,N_3939);
or U4380 (N_4380,N_3625,N_3886);
or U4381 (N_4381,N_3730,N_3671);
and U4382 (N_4382,N_3915,N_3887);
nand U4383 (N_4383,N_3503,N_3906);
nand U4384 (N_4384,N_3960,N_3876);
nand U4385 (N_4385,N_3689,N_3869);
or U4386 (N_4386,N_3646,N_3534);
or U4387 (N_4387,N_3612,N_3555);
and U4388 (N_4388,N_3836,N_3558);
nand U4389 (N_4389,N_3625,N_3908);
nand U4390 (N_4390,N_3695,N_3915);
nand U4391 (N_4391,N_3957,N_3627);
nor U4392 (N_4392,N_3743,N_3616);
nand U4393 (N_4393,N_3529,N_3842);
nor U4394 (N_4394,N_3753,N_3773);
and U4395 (N_4395,N_3931,N_3709);
nand U4396 (N_4396,N_3980,N_3739);
and U4397 (N_4397,N_3709,N_3977);
xnor U4398 (N_4398,N_3824,N_3762);
nand U4399 (N_4399,N_3694,N_3913);
nand U4400 (N_4400,N_3805,N_3523);
nand U4401 (N_4401,N_3634,N_3803);
nor U4402 (N_4402,N_3922,N_3880);
nor U4403 (N_4403,N_3561,N_3648);
nand U4404 (N_4404,N_3617,N_3922);
and U4405 (N_4405,N_3758,N_3532);
and U4406 (N_4406,N_3970,N_3807);
or U4407 (N_4407,N_3933,N_3831);
xor U4408 (N_4408,N_3579,N_3606);
and U4409 (N_4409,N_3885,N_3947);
nor U4410 (N_4410,N_3898,N_3987);
and U4411 (N_4411,N_3933,N_3500);
xor U4412 (N_4412,N_3776,N_3733);
or U4413 (N_4413,N_3941,N_3600);
xor U4414 (N_4414,N_3576,N_3987);
or U4415 (N_4415,N_3697,N_3844);
or U4416 (N_4416,N_3774,N_3896);
and U4417 (N_4417,N_3710,N_3977);
xor U4418 (N_4418,N_3792,N_3731);
nand U4419 (N_4419,N_3902,N_3630);
or U4420 (N_4420,N_3706,N_3660);
xor U4421 (N_4421,N_3853,N_3931);
nand U4422 (N_4422,N_3936,N_3514);
and U4423 (N_4423,N_3635,N_3667);
or U4424 (N_4424,N_3554,N_3760);
xor U4425 (N_4425,N_3674,N_3558);
xnor U4426 (N_4426,N_3521,N_3633);
xnor U4427 (N_4427,N_3533,N_3703);
nand U4428 (N_4428,N_3913,N_3956);
nor U4429 (N_4429,N_3528,N_3535);
and U4430 (N_4430,N_3947,N_3529);
nand U4431 (N_4431,N_3649,N_3548);
xnor U4432 (N_4432,N_3761,N_3857);
and U4433 (N_4433,N_3992,N_3616);
nand U4434 (N_4434,N_3829,N_3975);
xnor U4435 (N_4435,N_3731,N_3974);
nand U4436 (N_4436,N_3679,N_3561);
nor U4437 (N_4437,N_3919,N_3733);
xor U4438 (N_4438,N_3901,N_3996);
and U4439 (N_4439,N_3600,N_3568);
nor U4440 (N_4440,N_3644,N_3790);
or U4441 (N_4441,N_3582,N_3720);
or U4442 (N_4442,N_3615,N_3766);
and U4443 (N_4443,N_3986,N_3767);
xor U4444 (N_4444,N_3928,N_3572);
nand U4445 (N_4445,N_3834,N_3783);
and U4446 (N_4446,N_3907,N_3835);
and U4447 (N_4447,N_3905,N_3753);
xnor U4448 (N_4448,N_3852,N_3735);
nand U4449 (N_4449,N_3535,N_3991);
and U4450 (N_4450,N_3646,N_3874);
or U4451 (N_4451,N_3764,N_3767);
xor U4452 (N_4452,N_3603,N_3598);
nand U4453 (N_4453,N_3895,N_3765);
and U4454 (N_4454,N_3587,N_3600);
or U4455 (N_4455,N_3916,N_3581);
nand U4456 (N_4456,N_3814,N_3745);
xor U4457 (N_4457,N_3770,N_3805);
xor U4458 (N_4458,N_3954,N_3576);
and U4459 (N_4459,N_3527,N_3783);
and U4460 (N_4460,N_3864,N_3841);
xor U4461 (N_4461,N_3656,N_3509);
or U4462 (N_4462,N_3744,N_3511);
nand U4463 (N_4463,N_3899,N_3965);
and U4464 (N_4464,N_3828,N_3892);
xor U4465 (N_4465,N_3565,N_3895);
nand U4466 (N_4466,N_3749,N_3805);
nor U4467 (N_4467,N_3922,N_3924);
nor U4468 (N_4468,N_3949,N_3761);
xnor U4469 (N_4469,N_3900,N_3754);
xnor U4470 (N_4470,N_3902,N_3943);
nand U4471 (N_4471,N_3756,N_3746);
and U4472 (N_4472,N_3811,N_3648);
nor U4473 (N_4473,N_3543,N_3882);
or U4474 (N_4474,N_3718,N_3953);
and U4475 (N_4475,N_3537,N_3669);
nor U4476 (N_4476,N_3979,N_3560);
xor U4477 (N_4477,N_3665,N_3525);
nand U4478 (N_4478,N_3581,N_3532);
xnor U4479 (N_4479,N_3577,N_3893);
nand U4480 (N_4480,N_3845,N_3549);
or U4481 (N_4481,N_3976,N_3879);
xor U4482 (N_4482,N_3664,N_3939);
and U4483 (N_4483,N_3515,N_3635);
and U4484 (N_4484,N_3685,N_3770);
or U4485 (N_4485,N_3743,N_3858);
or U4486 (N_4486,N_3960,N_3766);
nand U4487 (N_4487,N_3947,N_3935);
xor U4488 (N_4488,N_3630,N_3759);
nor U4489 (N_4489,N_3527,N_3502);
nand U4490 (N_4490,N_3864,N_3557);
and U4491 (N_4491,N_3644,N_3969);
nor U4492 (N_4492,N_3906,N_3668);
or U4493 (N_4493,N_3591,N_3771);
nand U4494 (N_4494,N_3862,N_3953);
nor U4495 (N_4495,N_3526,N_3898);
xnor U4496 (N_4496,N_3534,N_3655);
nand U4497 (N_4497,N_3706,N_3749);
or U4498 (N_4498,N_3963,N_3594);
nor U4499 (N_4499,N_3676,N_3886);
nor U4500 (N_4500,N_4062,N_4485);
or U4501 (N_4501,N_4070,N_4229);
nand U4502 (N_4502,N_4367,N_4429);
or U4503 (N_4503,N_4279,N_4009);
or U4504 (N_4504,N_4152,N_4327);
nor U4505 (N_4505,N_4054,N_4226);
nand U4506 (N_4506,N_4449,N_4460);
nand U4507 (N_4507,N_4237,N_4117);
nand U4508 (N_4508,N_4334,N_4476);
nand U4509 (N_4509,N_4042,N_4256);
nand U4510 (N_4510,N_4242,N_4058);
and U4511 (N_4511,N_4266,N_4398);
and U4512 (N_4512,N_4369,N_4496);
nor U4513 (N_4513,N_4383,N_4265);
xnor U4514 (N_4514,N_4444,N_4345);
nor U4515 (N_4515,N_4132,N_4257);
nor U4516 (N_4516,N_4119,N_4074);
nor U4517 (N_4517,N_4232,N_4135);
nor U4518 (N_4518,N_4436,N_4061);
nor U4519 (N_4519,N_4362,N_4461);
or U4520 (N_4520,N_4254,N_4106);
or U4521 (N_4521,N_4238,N_4354);
or U4522 (N_4522,N_4252,N_4101);
and U4523 (N_4523,N_4373,N_4419);
or U4524 (N_4524,N_4183,N_4481);
nor U4525 (N_4525,N_4015,N_4191);
nand U4526 (N_4526,N_4044,N_4283);
xor U4527 (N_4527,N_4415,N_4071);
nor U4528 (N_4528,N_4236,N_4432);
and U4529 (N_4529,N_4091,N_4378);
or U4530 (N_4530,N_4418,N_4055);
or U4531 (N_4531,N_4017,N_4412);
nand U4532 (N_4532,N_4231,N_4239);
and U4533 (N_4533,N_4249,N_4387);
nor U4534 (N_4534,N_4394,N_4255);
xnor U4535 (N_4535,N_4338,N_4423);
xnor U4536 (N_4536,N_4080,N_4483);
and U4537 (N_4537,N_4172,N_4308);
and U4538 (N_4538,N_4114,N_4408);
nor U4539 (N_4539,N_4318,N_4205);
nor U4540 (N_4540,N_4303,N_4122);
nor U4541 (N_4541,N_4220,N_4227);
and U4542 (N_4542,N_4385,N_4014);
nand U4543 (N_4543,N_4068,N_4079);
or U4544 (N_4544,N_4355,N_4134);
nand U4545 (N_4545,N_4399,N_4243);
nor U4546 (N_4546,N_4098,N_4032);
and U4547 (N_4547,N_4007,N_4493);
nand U4548 (N_4548,N_4333,N_4420);
nor U4549 (N_4549,N_4397,N_4435);
nand U4550 (N_4550,N_4371,N_4075);
or U4551 (N_4551,N_4196,N_4351);
nand U4552 (N_4552,N_4182,N_4206);
nor U4553 (N_4553,N_4212,N_4314);
nor U4554 (N_4554,N_4190,N_4088);
nand U4555 (N_4555,N_4467,N_4041);
nor U4556 (N_4556,N_4057,N_4019);
or U4557 (N_4557,N_4407,N_4111);
nor U4558 (N_4558,N_4443,N_4011);
xor U4559 (N_4559,N_4001,N_4305);
xor U4560 (N_4560,N_4386,N_4171);
nand U4561 (N_4561,N_4459,N_4175);
or U4562 (N_4562,N_4343,N_4274);
nand U4563 (N_4563,N_4250,N_4286);
and U4564 (N_4564,N_4102,N_4374);
nor U4565 (N_4565,N_4275,N_4324);
or U4566 (N_4566,N_4277,N_4160);
nand U4567 (N_4567,N_4458,N_4240);
and U4568 (N_4568,N_4006,N_4293);
nor U4569 (N_4569,N_4472,N_4320);
and U4570 (N_4570,N_4203,N_4187);
nor U4571 (N_4571,N_4377,N_4225);
nor U4572 (N_4572,N_4086,N_4000);
or U4573 (N_4573,N_4368,N_4005);
and U4574 (N_4574,N_4149,N_4004);
or U4575 (N_4575,N_4451,N_4163);
nor U4576 (N_4576,N_4141,N_4161);
and U4577 (N_4577,N_4494,N_4211);
xnor U4578 (N_4578,N_4213,N_4395);
and U4579 (N_4579,N_4440,N_4341);
nand U4580 (N_4580,N_4356,N_4261);
or U4581 (N_4581,N_4193,N_4025);
and U4582 (N_4582,N_4270,N_4137);
nand U4583 (N_4583,N_4123,N_4477);
xor U4584 (N_4584,N_4108,N_4046);
nor U4585 (N_4585,N_4309,N_4468);
nand U4586 (N_4586,N_4448,N_4072);
xor U4587 (N_4587,N_4221,N_4142);
nor U4588 (N_4588,N_4370,N_4234);
xnor U4589 (N_4589,N_4124,N_4159);
or U4590 (N_4590,N_4082,N_4428);
nand U4591 (N_4591,N_4083,N_4092);
xor U4592 (N_4592,N_4131,N_4487);
and U4593 (N_4593,N_4499,N_4260);
xor U4594 (N_4594,N_4329,N_4197);
or U4595 (N_4595,N_4396,N_4118);
and U4596 (N_4596,N_4437,N_4405);
nor U4597 (N_4597,N_4267,N_4363);
xnor U4598 (N_4598,N_4013,N_4328);
and U4599 (N_4599,N_4120,N_4115);
nor U4600 (N_4600,N_4099,N_4352);
nand U4601 (N_4601,N_4392,N_4199);
or U4602 (N_4602,N_4219,N_4188);
nor U4603 (N_4603,N_4390,N_4282);
or U4604 (N_4604,N_4349,N_4488);
or U4605 (N_4605,N_4174,N_4288);
and U4606 (N_4606,N_4301,N_4469);
or U4607 (N_4607,N_4204,N_4002);
xor U4608 (N_4608,N_4143,N_4400);
and U4609 (N_4609,N_4081,N_4276);
nor U4610 (N_4610,N_4186,N_4248);
nor U4611 (N_4611,N_4037,N_4184);
and U4612 (N_4612,N_4312,N_4381);
xor U4613 (N_4613,N_4416,N_4410);
and U4614 (N_4614,N_4284,N_4421);
and U4615 (N_4615,N_4112,N_4452);
xnor U4616 (N_4616,N_4090,N_4136);
and U4617 (N_4617,N_4166,N_4024);
xor U4618 (N_4618,N_4036,N_4030);
nor U4619 (N_4619,N_4358,N_4097);
and U4620 (N_4620,N_4455,N_4273);
nor U4621 (N_4621,N_4315,N_4127);
and U4622 (N_4622,N_4235,N_4389);
and U4623 (N_4623,N_4475,N_4100);
nand U4624 (N_4624,N_4375,N_4177);
and U4625 (N_4625,N_4218,N_4294);
xor U4626 (N_4626,N_4317,N_4291);
and U4627 (N_4627,N_4129,N_4048);
xnor U4628 (N_4628,N_4052,N_4382);
xor U4629 (N_4629,N_4128,N_4150);
nor U4630 (N_4630,N_4020,N_4178);
or U4631 (N_4631,N_4484,N_4165);
nand U4632 (N_4632,N_4035,N_4209);
nor U4633 (N_4633,N_4325,N_4495);
nor U4634 (N_4634,N_4195,N_4216);
or U4635 (N_4635,N_4430,N_4332);
nor U4636 (N_4636,N_4262,N_4189);
nand U4637 (N_4637,N_4076,N_4147);
nand U4638 (N_4638,N_4372,N_4393);
or U4639 (N_4639,N_4158,N_4326);
nand U4640 (N_4640,N_4380,N_4350);
xor U4641 (N_4641,N_4346,N_4245);
nand U4642 (N_4642,N_4034,N_4466);
nand U4643 (N_4643,N_4210,N_4446);
or U4644 (N_4644,N_4154,N_4425);
nand U4645 (N_4645,N_4482,N_4281);
xor U4646 (N_4646,N_4008,N_4029);
or U4647 (N_4647,N_4251,N_4295);
nor U4648 (N_4648,N_4296,N_4103);
nand U4649 (N_4649,N_4464,N_4157);
or U4650 (N_4650,N_4010,N_4463);
nand U4651 (N_4651,N_4321,N_4357);
or U4652 (N_4652,N_4489,N_4116);
nor U4653 (N_4653,N_4376,N_4202);
or U4654 (N_4654,N_4109,N_4066);
or U4655 (N_4655,N_4170,N_4162);
nand U4656 (N_4656,N_4126,N_4297);
xor U4657 (N_4657,N_4271,N_4322);
nand U4658 (N_4658,N_4268,N_4050);
nand U4659 (N_4659,N_4300,N_4223);
and U4660 (N_4660,N_4105,N_4285);
xnor U4661 (N_4661,N_4307,N_4454);
and U4662 (N_4662,N_4292,N_4038);
xor U4663 (N_4663,N_4094,N_4153);
xnor U4664 (N_4664,N_4304,N_4053);
nand U4665 (N_4665,N_4330,N_4089);
xor U4666 (N_4666,N_4471,N_4391);
xnor U4667 (N_4667,N_4156,N_4388);
and U4668 (N_4668,N_4096,N_4201);
nor U4669 (N_4669,N_4028,N_4169);
xor U4670 (N_4670,N_4125,N_4479);
or U4671 (N_4671,N_4104,N_4043);
xor U4672 (N_4672,N_4364,N_4138);
nand U4673 (N_4673,N_4168,N_4264);
or U4674 (N_4674,N_4133,N_4215);
and U4675 (N_4675,N_4272,N_4491);
nand U4676 (N_4676,N_4474,N_4478);
nor U4677 (N_4677,N_4045,N_4176);
xor U4678 (N_4678,N_4480,N_4064);
nand U4679 (N_4679,N_4319,N_4462);
or U4680 (N_4680,N_4185,N_4450);
and U4681 (N_4681,N_4414,N_4016);
or U4682 (N_4682,N_4077,N_4051);
xor U4683 (N_4683,N_4148,N_4340);
xnor U4684 (N_4684,N_4253,N_4442);
nor U4685 (N_4685,N_4078,N_4224);
and U4686 (N_4686,N_4409,N_4208);
xnor U4687 (N_4687,N_4031,N_4233);
nor U4688 (N_4688,N_4289,N_4490);
or U4689 (N_4689,N_4084,N_4198);
nor U4690 (N_4690,N_4039,N_4403);
xnor U4691 (N_4691,N_4003,N_4060);
xor U4692 (N_4692,N_4151,N_4207);
nand U4693 (N_4693,N_4263,N_4228);
nor U4694 (N_4694,N_4447,N_4331);
nor U4695 (N_4695,N_4366,N_4306);
or U4696 (N_4696,N_4402,N_4427);
xor U4697 (N_4697,N_4336,N_4180);
xnor U4698 (N_4698,N_4313,N_4217);
or U4699 (N_4699,N_4085,N_4269);
or U4700 (N_4700,N_4335,N_4379);
nand U4701 (N_4701,N_4069,N_4065);
and U4702 (N_4702,N_4087,N_4200);
or U4703 (N_4703,N_4145,N_4107);
xor U4704 (N_4704,N_4047,N_4438);
or U4705 (N_4705,N_4139,N_4167);
nand U4706 (N_4706,N_4498,N_4337);
or U4707 (N_4707,N_4040,N_4339);
xor U4708 (N_4708,N_4113,N_4347);
xor U4709 (N_4709,N_4173,N_4130);
and U4710 (N_4710,N_4473,N_4018);
xor U4711 (N_4711,N_4311,N_4302);
nor U4712 (N_4712,N_4348,N_4280);
or U4713 (N_4713,N_4023,N_4144);
and U4714 (N_4714,N_4146,N_4365);
xnor U4715 (N_4715,N_4049,N_4056);
nand U4716 (N_4716,N_4359,N_4310);
nand U4717 (N_4717,N_4456,N_4194);
and U4718 (N_4718,N_4299,N_4422);
nor U4719 (N_4719,N_4492,N_4093);
or U4720 (N_4720,N_4360,N_4067);
nor U4721 (N_4721,N_4246,N_4431);
xor U4722 (N_4722,N_4247,N_4214);
xnor U4723 (N_4723,N_4445,N_4095);
or U4724 (N_4724,N_4278,N_4316);
nor U4725 (N_4725,N_4026,N_4441);
nand U4726 (N_4726,N_4424,N_4433);
nand U4727 (N_4727,N_4063,N_4298);
nor U4728 (N_4728,N_4027,N_4406);
or U4729 (N_4729,N_4073,N_4259);
nor U4730 (N_4730,N_4439,N_4486);
nand U4731 (N_4731,N_4401,N_4110);
or U4732 (N_4732,N_4192,N_4155);
and U4733 (N_4733,N_4059,N_4465);
xnor U4734 (N_4734,N_4434,N_4497);
nand U4735 (N_4735,N_4344,N_4384);
nand U4736 (N_4736,N_4222,N_4164);
nand U4737 (N_4737,N_4353,N_4413);
xnor U4738 (N_4738,N_4181,N_4258);
and U4739 (N_4739,N_4121,N_4033);
nor U4740 (N_4740,N_4290,N_4342);
nor U4741 (N_4741,N_4417,N_4426);
and U4742 (N_4742,N_4241,N_4140);
or U4743 (N_4743,N_4012,N_4361);
and U4744 (N_4744,N_4022,N_4470);
nor U4745 (N_4745,N_4287,N_4404);
or U4746 (N_4746,N_4453,N_4323);
nand U4747 (N_4747,N_4411,N_4230);
or U4748 (N_4748,N_4244,N_4457);
and U4749 (N_4749,N_4021,N_4179);
and U4750 (N_4750,N_4459,N_4333);
xor U4751 (N_4751,N_4135,N_4035);
nand U4752 (N_4752,N_4208,N_4473);
and U4753 (N_4753,N_4469,N_4085);
nor U4754 (N_4754,N_4248,N_4387);
nor U4755 (N_4755,N_4270,N_4460);
xnor U4756 (N_4756,N_4282,N_4333);
nand U4757 (N_4757,N_4205,N_4053);
nand U4758 (N_4758,N_4007,N_4413);
or U4759 (N_4759,N_4078,N_4207);
or U4760 (N_4760,N_4075,N_4413);
and U4761 (N_4761,N_4234,N_4191);
xnor U4762 (N_4762,N_4088,N_4150);
or U4763 (N_4763,N_4478,N_4436);
and U4764 (N_4764,N_4122,N_4128);
and U4765 (N_4765,N_4086,N_4282);
xor U4766 (N_4766,N_4128,N_4287);
and U4767 (N_4767,N_4340,N_4385);
and U4768 (N_4768,N_4414,N_4063);
xnor U4769 (N_4769,N_4455,N_4206);
nor U4770 (N_4770,N_4309,N_4066);
or U4771 (N_4771,N_4460,N_4327);
or U4772 (N_4772,N_4145,N_4104);
nand U4773 (N_4773,N_4076,N_4433);
and U4774 (N_4774,N_4280,N_4386);
nor U4775 (N_4775,N_4051,N_4097);
and U4776 (N_4776,N_4184,N_4436);
nand U4777 (N_4777,N_4275,N_4184);
xor U4778 (N_4778,N_4302,N_4361);
xnor U4779 (N_4779,N_4213,N_4264);
or U4780 (N_4780,N_4369,N_4171);
nand U4781 (N_4781,N_4311,N_4171);
nor U4782 (N_4782,N_4167,N_4013);
or U4783 (N_4783,N_4460,N_4310);
nand U4784 (N_4784,N_4111,N_4388);
nor U4785 (N_4785,N_4486,N_4000);
or U4786 (N_4786,N_4495,N_4351);
nor U4787 (N_4787,N_4164,N_4284);
and U4788 (N_4788,N_4133,N_4082);
nand U4789 (N_4789,N_4482,N_4264);
xor U4790 (N_4790,N_4420,N_4099);
xor U4791 (N_4791,N_4441,N_4196);
xnor U4792 (N_4792,N_4321,N_4346);
nor U4793 (N_4793,N_4097,N_4147);
or U4794 (N_4794,N_4478,N_4292);
or U4795 (N_4795,N_4324,N_4447);
nor U4796 (N_4796,N_4463,N_4065);
or U4797 (N_4797,N_4223,N_4492);
and U4798 (N_4798,N_4397,N_4483);
or U4799 (N_4799,N_4423,N_4210);
or U4800 (N_4800,N_4357,N_4225);
nor U4801 (N_4801,N_4491,N_4215);
and U4802 (N_4802,N_4363,N_4196);
or U4803 (N_4803,N_4026,N_4216);
xnor U4804 (N_4804,N_4358,N_4174);
and U4805 (N_4805,N_4244,N_4407);
xor U4806 (N_4806,N_4248,N_4490);
or U4807 (N_4807,N_4026,N_4365);
and U4808 (N_4808,N_4498,N_4315);
or U4809 (N_4809,N_4190,N_4413);
nand U4810 (N_4810,N_4183,N_4057);
and U4811 (N_4811,N_4281,N_4083);
xnor U4812 (N_4812,N_4334,N_4262);
or U4813 (N_4813,N_4347,N_4373);
xor U4814 (N_4814,N_4358,N_4018);
nand U4815 (N_4815,N_4452,N_4093);
nand U4816 (N_4816,N_4280,N_4225);
xor U4817 (N_4817,N_4382,N_4296);
and U4818 (N_4818,N_4189,N_4135);
xor U4819 (N_4819,N_4368,N_4002);
and U4820 (N_4820,N_4414,N_4067);
and U4821 (N_4821,N_4337,N_4077);
nand U4822 (N_4822,N_4273,N_4014);
or U4823 (N_4823,N_4368,N_4364);
or U4824 (N_4824,N_4499,N_4254);
and U4825 (N_4825,N_4431,N_4172);
nor U4826 (N_4826,N_4441,N_4334);
and U4827 (N_4827,N_4185,N_4334);
or U4828 (N_4828,N_4223,N_4097);
or U4829 (N_4829,N_4447,N_4454);
nor U4830 (N_4830,N_4436,N_4236);
and U4831 (N_4831,N_4138,N_4473);
nand U4832 (N_4832,N_4317,N_4085);
nor U4833 (N_4833,N_4098,N_4352);
nor U4834 (N_4834,N_4355,N_4299);
and U4835 (N_4835,N_4086,N_4380);
xnor U4836 (N_4836,N_4104,N_4401);
nor U4837 (N_4837,N_4298,N_4385);
nor U4838 (N_4838,N_4306,N_4084);
nor U4839 (N_4839,N_4498,N_4063);
nand U4840 (N_4840,N_4098,N_4048);
and U4841 (N_4841,N_4481,N_4383);
xor U4842 (N_4842,N_4467,N_4293);
and U4843 (N_4843,N_4492,N_4072);
nor U4844 (N_4844,N_4470,N_4041);
nor U4845 (N_4845,N_4477,N_4300);
and U4846 (N_4846,N_4253,N_4326);
and U4847 (N_4847,N_4336,N_4331);
nor U4848 (N_4848,N_4324,N_4492);
and U4849 (N_4849,N_4115,N_4221);
nand U4850 (N_4850,N_4052,N_4193);
xor U4851 (N_4851,N_4207,N_4005);
and U4852 (N_4852,N_4108,N_4448);
xnor U4853 (N_4853,N_4005,N_4091);
and U4854 (N_4854,N_4236,N_4305);
nor U4855 (N_4855,N_4443,N_4020);
nor U4856 (N_4856,N_4325,N_4193);
nor U4857 (N_4857,N_4402,N_4406);
or U4858 (N_4858,N_4094,N_4390);
and U4859 (N_4859,N_4406,N_4477);
xor U4860 (N_4860,N_4382,N_4290);
xnor U4861 (N_4861,N_4216,N_4365);
nand U4862 (N_4862,N_4437,N_4418);
or U4863 (N_4863,N_4121,N_4407);
xor U4864 (N_4864,N_4089,N_4357);
nor U4865 (N_4865,N_4428,N_4200);
xor U4866 (N_4866,N_4463,N_4202);
or U4867 (N_4867,N_4086,N_4144);
and U4868 (N_4868,N_4101,N_4468);
nor U4869 (N_4869,N_4461,N_4474);
or U4870 (N_4870,N_4006,N_4074);
nand U4871 (N_4871,N_4256,N_4268);
nor U4872 (N_4872,N_4258,N_4175);
nor U4873 (N_4873,N_4298,N_4133);
nor U4874 (N_4874,N_4459,N_4141);
nand U4875 (N_4875,N_4453,N_4205);
and U4876 (N_4876,N_4231,N_4480);
nand U4877 (N_4877,N_4426,N_4339);
or U4878 (N_4878,N_4233,N_4431);
xnor U4879 (N_4879,N_4306,N_4221);
and U4880 (N_4880,N_4089,N_4208);
nand U4881 (N_4881,N_4260,N_4108);
or U4882 (N_4882,N_4009,N_4291);
xnor U4883 (N_4883,N_4290,N_4194);
xnor U4884 (N_4884,N_4135,N_4456);
nor U4885 (N_4885,N_4288,N_4488);
and U4886 (N_4886,N_4009,N_4207);
and U4887 (N_4887,N_4481,N_4240);
xnor U4888 (N_4888,N_4481,N_4052);
or U4889 (N_4889,N_4496,N_4120);
or U4890 (N_4890,N_4132,N_4479);
nor U4891 (N_4891,N_4438,N_4347);
or U4892 (N_4892,N_4434,N_4144);
and U4893 (N_4893,N_4045,N_4289);
and U4894 (N_4894,N_4326,N_4050);
nor U4895 (N_4895,N_4188,N_4379);
and U4896 (N_4896,N_4099,N_4027);
and U4897 (N_4897,N_4426,N_4095);
xor U4898 (N_4898,N_4489,N_4238);
nand U4899 (N_4899,N_4283,N_4499);
and U4900 (N_4900,N_4331,N_4204);
or U4901 (N_4901,N_4423,N_4296);
nand U4902 (N_4902,N_4059,N_4247);
nor U4903 (N_4903,N_4245,N_4325);
and U4904 (N_4904,N_4458,N_4064);
xnor U4905 (N_4905,N_4458,N_4183);
nand U4906 (N_4906,N_4028,N_4208);
nand U4907 (N_4907,N_4224,N_4414);
and U4908 (N_4908,N_4470,N_4149);
or U4909 (N_4909,N_4459,N_4177);
xor U4910 (N_4910,N_4356,N_4191);
and U4911 (N_4911,N_4271,N_4277);
nand U4912 (N_4912,N_4333,N_4161);
xor U4913 (N_4913,N_4371,N_4233);
and U4914 (N_4914,N_4319,N_4302);
nor U4915 (N_4915,N_4426,N_4110);
or U4916 (N_4916,N_4108,N_4128);
nor U4917 (N_4917,N_4071,N_4237);
and U4918 (N_4918,N_4483,N_4090);
and U4919 (N_4919,N_4258,N_4058);
nand U4920 (N_4920,N_4227,N_4131);
nor U4921 (N_4921,N_4135,N_4155);
and U4922 (N_4922,N_4015,N_4473);
xor U4923 (N_4923,N_4267,N_4026);
nand U4924 (N_4924,N_4133,N_4420);
or U4925 (N_4925,N_4269,N_4243);
nor U4926 (N_4926,N_4453,N_4479);
and U4927 (N_4927,N_4018,N_4289);
or U4928 (N_4928,N_4336,N_4472);
and U4929 (N_4929,N_4114,N_4363);
nand U4930 (N_4930,N_4113,N_4438);
nand U4931 (N_4931,N_4162,N_4447);
and U4932 (N_4932,N_4232,N_4449);
or U4933 (N_4933,N_4078,N_4476);
or U4934 (N_4934,N_4211,N_4398);
xnor U4935 (N_4935,N_4432,N_4253);
nand U4936 (N_4936,N_4326,N_4144);
or U4937 (N_4937,N_4405,N_4186);
nand U4938 (N_4938,N_4278,N_4370);
and U4939 (N_4939,N_4343,N_4485);
xor U4940 (N_4940,N_4355,N_4047);
xor U4941 (N_4941,N_4271,N_4360);
nor U4942 (N_4942,N_4220,N_4002);
or U4943 (N_4943,N_4090,N_4156);
xor U4944 (N_4944,N_4328,N_4182);
xor U4945 (N_4945,N_4489,N_4218);
xor U4946 (N_4946,N_4409,N_4440);
nor U4947 (N_4947,N_4435,N_4292);
nor U4948 (N_4948,N_4493,N_4322);
nor U4949 (N_4949,N_4346,N_4359);
or U4950 (N_4950,N_4250,N_4481);
nor U4951 (N_4951,N_4115,N_4194);
xor U4952 (N_4952,N_4160,N_4366);
or U4953 (N_4953,N_4495,N_4247);
or U4954 (N_4954,N_4088,N_4485);
and U4955 (N_4955,N_4038,N_4240);
and U4956 (N_4956,N_4017,N_4420);
nand U4957 (N_4957,N_4242,N_4409);
nor U4958 (N_4958,N_4141,N_4421);
nand U4959 (N_4959,N_4054,N_4376);
nor U4960 (N_4960,N_4302,N_4212);
or U4961 (N_4961,N_4331,N_4366);
or U4962 (N_4962,N_4001,N_4387);
nand U4963 (N_4963,N_4290,N_4287);
nor U4964 (N_4964,N_4312,N_4109);
nor U4965 (N_4965,N_4247,N_4434);
xor U4966 (N_4966,N_4170,N_4378);
and U4967 (N_4967,N_4301,N_4256);
nor U4968 (N_4968,N_4445,N_4098);
or U4969 (N_4969,N_4279,N_4415);
xor U4970 (N_4970,N_4189,N_4432);
nand U4971 (N_4971,N_4052,N_4293);
nand U4972 (N_4972,N_4178,N_4246);
xor U4973 (N_4973,N_4084,N_4385);
nand U4974 (N_4974,N_4476,N_4280);
and U4975 (N_4975,N_4122,N_4447);
and U4976 (N_4976,N_4241,N_4118);
and U4977 (N_4977,N_4346,N_4110);
and U4978 (N_4978,N_4159,N_4224);
nor U4979 (N_4979,N_4197,N_4300);
nand U4980 (N_4980,N_4200,N_4316);
and U4981 (N_4981,N_4231,N_4497);
xor U4982 (N_4982,N_4072,N_4134);
or U4983 (N_4983,N_4240,N_4313);
or U4984 (N_4984,N_4364,N_4230);
and U4985 (N_4985,N_4474,N_4287);
nand U4986 (N_4986,N_4335,N_4117);
nand U4987 (N_4987,N_4051,N_4168);
and U4988 (N_4988,N_4398,N_4179);
nor U4989 (N_4989,N_4438,N_4408);
nor U4990 (N_4990,N_4228,N_4332);
or U4991 (N_4991,N_4245,N_4049);
or U4992 (N_4992,N_4397,N_4127);
or U4993 (N_4993,N_4266,N_4052);
xor U4994 (N_4994,N_4224,N_4184);
and U4995 (N_4995,N_4043,N_4151);
nand U4996 (N_4996,N_4186,N_4470);
xnor U4997 (N_4997,N_4134,N_4170);
or U4998 (N_4998,N_4279,N_4416);
nand U4999 (N_4999,N_4038,N_4471);
xnor UO_0 (O_0,N_4558,N_4738);
nor UO_1 (O_1,N_4735,N_4579);
nor UO_2 (O_2,N_4870,N_4863);
nand UO_3 (O_3,N_4981,N_4925);
and UO_4 (O_4,N_4764,N_4915);
nand UO_5 (O_5,N_4512,N_4517);
xor UO_6 (O_6,N_4903,N_4884);
nor UO_7 (O_7,N_4799,N_4922);
or UO_8 (O_8,N_4840,N_4741);
nor UO_9 (O_9,N_4580,N_4762);
nand UO_10 (O_10,N_4742,N_4541);
nor UO_11 (O_11,N_4706,N_4542);
or UO_12 (O_12,N_4530,N_4511);
and UO_13 (O_13,N_4792,N_4958);
and UO_14 (O_14,N_4613,N_4784);
xor UO_15 (O_15,N_4631,N_4749);
or UO_16 (O_16,N_4565,N_4848);
and UO_17 (O_17,N_4534,N_4798);
xor UO_18 (O_18,N_4937,N_4805);
nand UO_19 (O_19,N_4596,N_4666);
nor UO_20 (O_20,N_4837,N_4747);
nand UO_21 (O_21,N_4627,N_4624);
and UO_22 (O_22,N_4868,N_4797);
xor UO_23 (O_23,N_4985,N_4947);
or UO_24 (O_24,N_4800,N_4990);
nand UO_25 (O_25,N_4639,N_4948);
or UO_26 (O_26,N_4982,N_4707);
and UO_27 (O_27,N_4543,N_4731);
and UO_28 (O_28,N_4720,N_4873);
or UO_29 (O_29,N_4655,N_4615);
or UO_30 (O_30,N_4779,N_4643);
xor UO_31 (O_31,N_4778,N_4519);
nor UO_32 (O_32,N_4700,N_4507);
or UO_33 (O_33,N_4988,N_4653);
nor UO_34 (O_34,N_4960,N_4644);
xor UO_35 (O_35,N_4630,N_4864);
or UO_36 (O_36,N_4516,N_4824);
or UO_37 (O_37,N_4629,N_4583);
nand UO_38 (O_38,N_4818,N_4640);
and UO_39 (O_39,N_4575,N_4692);
or UO_40 (O_40,N_4743,N_4756);
nor UO_41 (O_41,N_4670,N_4833);
nor UO_42 (O_42,N_4772,N_4637);
and UO_43 (O_43,N_4992,N_4725);
xnor UO_44 (O_44,N_4536,N_4621);
xnor UO_45 (O_45,N_4967,N_4562);
and UO_46 (O_46,N_4814,N_4683);
xnor UO_47 (O_47,N_4758,N_4578);
and UO_48 (O_48,N_4610,N_4500);
nand UO_49 (O_49,N_4964,N_4769);
xnor UO_50 (O_50,N_4813,N_4946);
xor UO_51 (O_51,N_4774,N_4592);
xnor UO_52 (O_52,N_4828,N_4972);
nand UO_53 (O_53,N_4574,N_4654);
or UO_54 (O_54,N_4667,N_4970);
and UO_55 (O_55,N_4938,N_4866);
and UO_56 (O_56,N_4555,N_4577);
xor UO_57 (O_57,N_4665,N_4770);
nor UO_58 (O_58,N_4994,N_4690);
or UO_59 (O_59,N_4913,N_4663);
or UO_60 (O_60,N_4538,N_4609);
and UO_61 (O_61,N_4673,N_4727);
xor UO_62 (O_62,N_4572,N_4573);
nand UO_63 (O_63,N_4827,N_4664);
and UO_64 (O_64,N_4995,N_4755);
nand UO_65 (O_65,N_4595,N_4636);
nor UO_66 (O_66,N_4715,N_4693);
and UO_67 (O_67,N_4851,N_4879);
nor UO_68 (O_68,N_4688,N_4872);
xor UO_69 (O_69,N_4569,N_4528);
or UO_70 (O_70,N_4689,N_4954);
or UO_71 (O_71,N_4899,N_4953);
or UO_72 (O_72,N_4815,N_4904);
nor UO_73 (O_73,N_4944,N_4829);
nand UO_74 (O_74,N_4976,N_4788);
or UO_75 (O_75,N_4561,N_4767);
nand UO_76 (O_76,N_4750,N_4748);
nor UO_77 (O_77,N_4614,N_4880);
and UO_78 (O_78,N_4980,N_4826);
xnor UO_79 (O_79,N_4998,N_4895);
or UO_80 (O_80,N_4724,N_4751);
nor UO_81 (O_81,N_4810,N_4878);
nor UO_82 (O_82,N_4726,N_4957);
or UO_83 (O_83,N_4783,N_4612);
xnor UO_84 (O_84,N_4794,N_4765);
xor UO_85 (O_85,N_4618,N_4539);
nor UO_86 (O_86,N_4703,N_4856);
nor UO_87 (O_87,N_4785,N_4682);
and UO_88 (O_88,N_4926,N_4917);
nor UO_89 (O_89,N_4734,N_4606);
nor UO_90 (O_90,N_4941,N_4846);
xnor UO_91 (O_91,N_4674,N_4831);
xor UO_92 (O_92,N_4527,N_4849);
nand UO_93 (O_93,N_4969,N_4563);
or UO_94 (O_94,N_4820,N_4696);
nand UO_95 (O_95,N_4597,N_4713);
nor UO_96 (O_96,N_4545,N_4830);
nor UO_97 (O_97,N_4845,N_4628);
nand UO_98 (O_98,N_4657,N_4656);
nor UO_99 (O_99,N_4716,N_4625);
xnor UO_100 (O_100,N_4699,N_4920);
or UO_101 (O_101,N_4841,N_4648);
or UO_102 (O_102,N_4590,N_4931);
or UO_103 (O_103,N_4984,N_4997);
or UO_104 (O_104,N_4855,N_4681);
nand UO_105 (O_105,N_4897,N_4679);
and UO_106 (O_106,N_4649,N_4701);
xnor UO_107 (O_107,N_4901,N_4651);
and UO_108 (O_108,N_4921,N_4705);
and UO_109 (O_109,N_4836,N_4605);
nand UO_110 (O_110,N_4773,N_4568);
or UO_111 (O_111,N_4822,N_4717);
nor UO_112 (O_112,N_4996,N_4671);
xor UO_113 (O_113,N_4812,N_4927);
or UO_114 (O_114,N_4566,N_4601);
nor UO_115 (O_115,N_4801,N_4771);
or UO_116 (O_116,N_4887,N_4702);
xnor UO_117 (O_117,N_4659,N_4504);
and UO_118 (O_118,N_4619,N_4515);
nand UO_119 (O_119,N_4554,N_4632);
nand UO_120 (O_120,N_4675,N_4687);
nor UO_121 (O_121,N_4802,N_4510);
and UO_122 (O_122,N_4875,N_4952);
nor UO_123 (O_123,N_4842,N_4730);
or UO_124 (O_124,N_4900,N_4834);
xor UO_125 (O_125,N_4823,N_4647);
xnor UO_126 (O_126,N_4959,N_4684);
xnor UO_127 (O_127,N_4962,N_4835);
nand UO_128 (O_128,N_4571,N_4932);
xor UO_129 (O_129,N_4719,N_4739);
or UO_130 (O_130,N_4943,N_4852);
xnor UO_131 (O_131,N_4733,N_4753);
xor UO_132 (O_132,N_4839,N_4916);
xnor UO_133 (O_133,N_4965,N_4894);
xor UO_134 (O_134,N_4918,N_4718);
xor UO_135 (O_135,N_4806,N_4677);
and UO_136 (O_136,N_4781,N_4514);
nand UO_137 (O_137,N_4914,N_4808);
or UO_138 (O_138,N_4503,N_4560);
or UO_139 (O_139,N_4722,N_4923);
nand UO_140 (O_140,N_4660,N_4961);
nand UO_141 (O_141,N_4721,N_4971);
and UO_142 (O_142,N_4912,N_4591);
xnor UO_143 (O_143,N_4593,N_4567);
and UO_144 (O_144,N_4782,N_4939);
and UO_145 (O_145,N_4861,N_4668);
and UO_146 (O_146,N_4803,N_4929);
nor UO_147 (O_147,N_4680,N_4844);
and UO_148 (O_148,N_4518,N_4807);
xnor UO_149 (O_149,N_4646,N_4607);
nor UO_150 (O_150,N_4854,N_4620);
nor UO_151 (O_151,N_4874,N_4711);
nand UO_152 (O_152,N_4871,N_4935);
nor UO_153 (O_153,N_4529,N_4780);
nand UO_154 (O_154,N_4626,N_4608);
nor UO_155 (O_155,N_4600,N_4816);
and UO_156 (O_156,N_4850,N_4505);
xor UO_157 (O_157,N_4987,N_4790);
xnor UO_158 (O_158,N_4676,N_4535);
and UO_159 (O_159,N_4736,N_4945);
xnor UO_160 (O_160,N_4732,N_4936);
nor UO_161 (O_161,N_4796,N_4532);
or UO_162 (O_162,N_4513,N_4766);
or UO_163 (O_163,N_4757,N_4893);
and UO_164 (O_164,N_4544,N_4754);
nor UO_165 (O_165,N_4832,N_4847);
nand UO_166 (O_166,N_4956,N_4729);
nand UO_167 (O_167,N_4641,N_4763);
nand UO_168 (O_168,N_4973,N_4890);
and UO_169 (O_169,N_4979,N_4645);
nor UO_170 (O_170,N_4672,N_4570);
nand UO_171 (O_171,N_4942,N_4599);
nor UO_172 (O_172,N_4502,N_4556);
nor UO_173 (O_173,N_4533,N_4564);
nor UO_174 (O_174,N_4709,N_4885);
and UO_175 (O_175,N_4869,N_4553);
nor UO_176 (O_176,N_4587,N_4616);
and UO_177 (O_177,N_4865,N_4652);
or UO_178 (O_178,N_4883,N_4905);
xor UO_179 (O_179,N_4949,N_4602);
and UO_180 (O_180,N_4603,N_4902);
or UO_181 (O_181,N_4858,N_4506);
nor UO_182 (O_182,N_4698,N_4522);
nand UO_183 (O_183,N_4633,N_4975);
nand UO_184 (O_184,N_4623,N_4910);
xnor UO_185 (O_185,N_4557,N_4898);
and UO_186 (O_186,N_4737,N_4746);
nor UO_187 (O_187,N_4789,N_4867);
xor UO_188 (O_188,N_4617,N_4886);
or UO_189 (O_189,N_4584,N_4907);
or UO_190 (O_190,N_4552,N_4974);
nor UO_191 (O_191,N_4508,N_4793);
xnor UO_192 (O_192,N_4691,N_4551);
xnor UO_193 (O_193,N_4638,N_4896);
nor UO_194 (O_194,N_4892,N_4550);
or UO_195 (O_195,N_4838,N_4786);
nand UO_196 (O_196,N_4882,N_4744);
and UO_197 (O_197,N_4585,N_4678);
nand UO_198 (O_198,N_4991,N_4752);
and UO_199 (O_199,N_4740,N_4582);
and UO_200 (O_200,N_4951,N_4549);
or UO_201 (O_201,N_4540,N_4934);
and UO_202 (O_202,N_4642,N_4804);
xnor UO_203 (O_203,N_4586,N_4876);
xnor UO_204 (O_204,N_4889,N_4968);
nor UO_205 (O_205,N_4695,N_4581);
or UO_206 (O_206,N_4776,N_4686);
or UO_207 (O_207,N_4548,N_4859);
nor UO_208 (O_208,N_4598,N_4594);
and UO_209 (O_209,N_4694,N_4999);
nor UO_210 (O_210,N_4635,N_4661);
nand UO_211 (O_211,N_4761,N_4930);
and UO_212 (O_212,N_4919,N_4521);
or UO_213 (O_213,N_4768,N_4817);
and UO_214 (O_214,N_4611,N_4723);
xor UO_215 (O_215,N_4860,N_4993);
nor UO_216 (O_216,N_4821,N_4714);
and UO_217 (O_217,N_4881,N_4911);
nor UO_218 (O_218,N_4650,N_4977);
nand UO_219 (O_219,N_4950,N_4728);
nor UO_220 (O_220,N_4523,N_4588);
xor UO_221 (O_221,N_4509,N_4819);
and UO_222 (O_222,N_4986,N_4685);
nand UO_223 (O_223,N_4966,N_4546);
nand UO_224 (O_224,N_4877,N_4760);
nand UO_225 (O_225,N_4908,N_4940);
nand UO_226 (O_226,N_4704,N_4983);
nor UO_227 (O_227,N_4775,N_4928);
nand UO_228 (O_228,N_4891,N_4909);
and UO_229 (O_229,N_4634,N_4759);
nor UO_230 (O_230,N_4525,N_4787);
xnor UO_231 (O_231,N_4888,N_4501);
xor UO_232 (O_232,N_4933,N_4537);
and UO_233 (O_233,N_4955,N_4710);
nand UO_234 (O_234,N_4531,N_4924);
and UO_235 (O_235,N_4658,N_4989);
nor UO_236 (O_236,N_4520,N_4604);
nand UO_237 (O_237,N_4547,N_4795);
nand UO_238 (O_238,N_4524,N_4669);
xor UO_239 (O_239,N_4589,N_4662);
nor UO_240 (O_240,N_4862,N_4745);
and UO_241 (O_241,N_4825,N_4712);
nand UO_242 (O_242,N_4843,N_4853);
and UO_243 (O_243,N_4708,N_4791);
or UO_244 (O_244,N_4978,N_4526);
and UO_245 (O_245,N_4777,N_4811);
nor UO_246 (O_246,N_4963,N_4622);
xnor UO_247 (O_247,N_4906,N_4559);
nand UO_248 (O_248,N_4697,N_4576);
or UO_249 (O_249,N_4809,N_4857);
and UO_250 (O_250,N_4833,N_4567);
xnor UO_251 (O_251,N_4597,N_4951);
or UO_252 (O_252,N_4645,N_4550);
or UO_253 (O_253,N_4756,N_4904);
nor UO_254 (O_254,N_4635,N_4652);
nor UO_255 (O_255,N_4698,N_4918);
nor UO_256 (O_256,N_4773,N_4686);
xnor UO_257 (O_257,N_4727,N_4703);
and UO_258 (O_258,N_4517,N_4581);
nor UO_259 (O_259,N_4986,N_4930);
nand UO_260 (O_260,N_4629,N_4979);
or UO_261 (O_261,N_4635,N_4951);
and UO_262 (O_262,N_4560,N_4575);
and UO_263 (O_263,N_4911,N_4728);
nor UO_264 (O_264,N_4805,N_4801);
and UO_265 (O_265,N_4778,N_4885);
xor UO_266 (O_266,N_4912,N_4938);
nand UO_267 (O_267,N_4580,N_4817);
nor UO_268 (O_268,N_4988,N_4513);
nor UO_269 (O_269,N_4692,N_4563);
nand UO_270 (O_270,N_4982,N_4757);
nand UO_271 (O_271,N_4830,N_4896);
nor UO_272 (O_272,N_4999,N_4523);
nor UO_273 (O_273,N_4999,N_4589);
nor UO_274 (O_274,N_4987,N_4989);
or UO_275 (O_275,N_4505,N_4989);
xor UO_276 (O_276,N_4733,N_4887);
xor UO_277 (O_277,N_4919,N_4740);
or UO_278 (O_278,N_4609,N_4887);
nand UO_279 (O_279,N_4652,N_4950);
nand UO_280 (O_280,N_4551,N_4956);
or UO_281 (O_281,N_4799,N_4530);
or UO_282 (O_282,N_4850,N_4963);
and UO_283 (O_283,N_4534,N_4665);
and UO_284 (O_284,N_4613,N_4843);
nand UO_285 (O_285,N_4639,N_4869);
nand UO_286 (O_286,N_4817,N_4937);
and UO_287 (O_287,N_4883,N_4918);
nor UO_288 (O_288,N_4547,N_4503);
nor UO_289 (O_289,N_4984,N_4937);
nor UO_290 (O_290,N_4904,N_4531);
and UO_291 (O_291,N_4747,N_4943);
or UO_292 (O_292,N_4995,N_4780);
nand UO_293 (O_293,N_4825,N_4692);
xnor UO_294 (O_294,N_4869,N_4889);
nand UO_295 (O_295,N_4793,N_4629);
nor UO_296 (O_296,N_4533,N_4529);
or UO_297 (O_297,N_4508,N_4539);
or UO_298 (O_298,N_4840,N_4983);
or UO_299 (O_299,N_4518,N_4575);
and UO_300 (O_300,N_4605,N_4612);
nand UO_301 (O_301,N_4601,N_4616);
and UO_302 (O_302,N_4559,N_4998);
or UO_303 (O_303,N_4947,N_4920);
nor UO_304 (O_304,N_4745,N_4943);
xor UO_305 (O_305,N_4983,N_4961);
nand UO_306 (O_306,N_4896,N_4813);
and UO_307 (O_307,N_4975,N_4968);
and UO_308 (O_308,N_4536,N_4748);
xor UO_309 (O_309,N_4624,N_4930);
and UO_310 (O_310,N_4745,N_4948);
nor UO_311 (O_311,N_4519,N_4686);
and UO_312 (O_312,N_4648,N_4616);
nand UO_313 (O_313,N_4583,N_4740);
nand UO_314 (O_314,N_4915,N_4627);
nor UO_315 (O_315,N_4544,N_4617);
nor UO_316 (O_316,N_4693,N_4626);
nand UO_317 (O_317,N_4734,N_4961);
nor UO_318 (O_318,N_4729,N_4845);
xnor UO_319 (O_319,N_4734,N_4663);
and UO_320 (O_320,N_4579,N_4607);
or UO_321 (O_321,N_4952,N_4579);
xnor UO_322 (O_322,N_4852,N_4634);
and UO_323 (O_323,N_4668,N_4743);
nand UO_324 (O_324,N_4784,N_4533);
or UO_325 (O_325,N_4660,N_4796);
nor UO_326 (O_326,N_4830,N_4584);
and UO_327 (O_327,N_4719,N_4668);
and UO_328 (O_328,N_4876,N_4991);
and UO_329 (O_329,N_4741,N_4691);
or UO_330 (O_330,N_4567,N_4621);
and UO_331 (O_331,N_4816,N_4713);
nor UO_332 (O_332,N_4511,N_4597);
and UO_333 (O_333,N_4737,N_4599);
or UO_334 (O_334,N_4502,N_4908);
nor UO_335 (O_335,N_4878,N_4539);
nor UO_336 (O_336,N_4809,N_4656);
xor UO_337 (O_337,N_4727,N_4640);
nor UO_338 (O_338,N_4597,N_4835);
nor UO_339 (O_339,N_4527,N_4953);
xnor UO_340 (O_340,N_4692,N_4643);
nor UO_341 (O_341,N_4707,N_4534);
xor UO_342 (O_342,N_4745,N_4758);
or UO_343 (O_343,N_4692,N_4842);
nor UO_344 (O_344,N_4846,N_4654);
xnor UO_345 (O_345,N_4543,N_4771);
and UO_346 (O_346,N_4665,N_4805);
and UO_347 (O_347,N_4662,N_4615);
nand UO_348 (O_348,N_4873,N_4880);
and UO_349 (O_349,N_4685,N_4776);
nand UO_350 (O_350,N_4628,N_4591);
nand UO_351 (O_351,N_4672,N_4912);
nor UO_352 (O_352,N_4747,N_4822);
or UO_353 (O_353,N_4997,N_4741);
and UO_354 (O_354,N_4748,N_4577);
nor UO_355 (O_355,N_4694,N_4652);
nand UO_356 (O_356,N_4868,N_4672);
xnor UO_357 (O_357,N_4799,N_4788);
and UO_358 (O_358,N_4840,N_4555);
xor UO_359 (O_359,N_4777,N_4923);
and UO_360 (O_360,N_4746,N_4780);
and UO_361 (O_361,N_4724,N_4683);
nand UO_362 (O_362,N_4540,N_4563);
nand UO_363 (O_363,N_4902,N_4786);
and UO_364 (O_364,N_4528,N_4580);
and UO_365 (O_365,N_4949,N_4851);
and UO_366 (O_366,N_4545,N_4988);
nor UO_367 (O_367,N_4537,N_4988);
xnor UO_368 (O_368,N_4827,N_4870);
nor UO_369 (O_369,N_4866,N_4946);
nor UO_370 (O_370,N_4834,N_4624);
nor UO_371 (O_371,N_4749,N_4958);
and UO_372 (O_372,N_4799,N_4932);
and UO_373 (O_373,N_4720,N_4729);
nor UO_374 (O_374,N_4739,N_4525);
or UO_375 (O_375,N_4771,N_4663);
xor UO_376 (O_376,N_4624,N_4553);
nand UO_377 (O_377,N_4658,N_4896);
nand UO_378 (O_378,N_4652,N_4610);
and UO_379 (O_379,N_4680,N_4688);
or UO_380 (O_380,N_4833,N_4649);
or UO_381 (O_381,N_4970,N_4977);
or UO_382 (O_382,N_4776,N_4757);
nor UO_383 (O_383,N_4693,N_4772);
and UO_384 (O_384,N_4883,N_4719);
nand UO_385 (O_385,N_4709,N_4510);
nor UO_386 (O_386,N_4769,N_4923);
nand UO_387 (O_387,N_4920,N_4791);
nand UO_388 (O_388,N_4661,N_4717);
nand UO_389 (O_389,N_4518,N_4910);
or UO_390 (O_390,N_4740,N_4796);
nand UO_391 (O_391,N_4544,N_4542);
and UO_392 (O_392,N_4508,N_4826);
xor UO_393 (O_393,N_4610,N_4626);
xnor UO_394 (O_394,N_4985,N_4952);
and UO_395 (O_395,N_4658,N_4909);
nor UO_396 (O_396,N_4607,N_4604);
or UO_397 (O_397,N_4533,N_4527);
or UO_398 (O_398,N_4951,N_4858);
xnor UO_399 (O_399,N_4690,N_4525);
nor UO_400 (O_400,N_4638,N_4777);
nor UO_401 (O_401,N_4647,N_4773);
xnor UO_402 (O_402,N_4985,N_4745);
nand UO_403 (O_403,N_4529,N_4787);
nor UO_404 (O_404,N_4735,N_4759);
and UO_405 (O_405,N_4595,N_4708);
nor UO_406 (O_406,N_4809,N_4727);
and UO_407 (O_407,N_4646,N_4726);
and UO_408 (O_408,N_4622,N_4900);
xnor UO_409 (O_409,N_4995,N_4736);
nand UO_410 (O_410,N_4741,N_4664);
nor UO_411 (O_411,N_4931,N_4909);
and UO_412 (O_412,N_4633,N_4589);
or UO_413 (O_413,N_4965,N_4847);
and UO_414 (O_414,N_4548,N_4667);
nand UO_415 (O_415,N_4701,N_4502);
and UO_416 (O_416,N_4986,N_4739);
xor UO_417 (O_417,N_4760,N_4561);
nor UO_418 (O_418,N_4796,N_4717);
nand UO_419 (O_419,N_4787,N_4877);
nand UO_420 (O_420,N_4773,N_4561);
xor UO_421 (O_421,N_4686,N_4623);
or UO_422 (O_422,N_4509,N_4541);
or UO_423 (O_423,N_4703,N_4936);
nor UO_424 (O_424,N_4570,N_4552);
xnor UO_425 (O_425,N_4761,N_4765);
nand UO_426 (O_426,N_4772,N_4508);
nand UO_427 (O_427,N_4823,N_4775);
nor UO_428 (O_428,N_4981,N_4857);
nor UO_429 (O_429,N_4720,N_4763);
or UO_430 (O_430,N_4563,N_4983);
xnor UO_431 (O_431,N_4640,N_4715);
xnor UO_432 (O_432,N_4668,N_4966);
and UO_433 (O_433,N_4940,N_4902);
nand UO_434 (O_434,N_4968,N_4846);
or UO_435 (O_435,N_4936,N_4756);
and UO_436 (O_436,N_4627,N_4913);
or UO_437 (O_437,N_4842,N_4883);
nand UO_438 (O_438,N_4725,N_4618);
or UO_439 (O_439,N_4790,N_4757);
xnor UO_440 (O_440,N_4981,N_4980);
nor UO_441 (O_441,N_4516,N_4983);
or UO_442 (O_442,N_4638,N_4582);
nor UO_443 (O_443,N_4839,N_4927);
or UO_444 (O_444,N_4638,N_4698);
or UO_445 (O_445,N_4577,N_4756);
or UO_446 (O_446,N_4837,N_4762);
and UO_447 (O_447,N_4770,N_4840);
nor UO_448 (O_448,N_4763,N_4597);
nor UO_449 (O_449,N_4912,N_4731);
nor UO_450 (O_450,N_4890,N_4814);
xnor UO_451 (O_451,N_4692,N_4844);
or UO_452 (O_452,N_4718,N_4867);
xor UO_453 (O_453,N_4722,N_4615);
nand UO_454 (O_454,N_4729,N_4866);
nand UO_455 (O_455,N_4500,N_4667);
or UO_456 (O_456,N_4862,N_4677);
nand UO_457 (O_457,N_4502,N_4934);
or UO_458 (O_458,N_4551,N_4778);
xor UO_459 (O_459,N_4981,N_4538);
xnor UO_460 (O_460,N_4562,N_4949);
and UO_461 (O_461,N_4887,N_4730);
xnor UO_462 (O_462,N_4939,N_4739);
xor UO_463 (O_463,N_4525,N_4693);
nor UO_464 (O_464,N_4826,N_4683);
xnor UO_465 (O_465,N_4700,N_4646);
nand UO_466 (O_466,N_4811,N_4604);
nand UO_467 (O_467,N_4609,N_4701);
nand UO_468 (O_468,N_4972,N_4801);
nor UO_469 (O_469,N_4816,N_4972);
nor UO_470 (O_470,N_4798,N_4980);
nand UO_471 (O_471,N_4874,N_4649);
nand UO_472 (O_472,N_4531,N_4602);
and UO_473 (O_473,N_4550,N_4911);
nor UO_474 (O_474,N_4921,N_4819);
or UO_475 (O_475,N_4989,N_4695);
and UO_476 (O_476,N_4588,N_4706);
nand UO_477 (O_477,N_4777,N_4906);
nor UO_478 (O_478,N_4549,N_4556);
nor UO_479 (O_479,N_4736,N_4737);
nor UO_480 (O_480,N_4817,N_4702);
or UO_481 (O_481,N_4642,N_4864);
nor UO_482 (O_482,N_4512,N_4794);
nor UO_483 (O_483,N_4572,N_4957);
and UO_484 (O_484,N_4845,N_4533);
and UO_485 (O_485,N_4702,N_4778);
and UO_486 (O_486,N_4525,N_4905);
or UO_487 (O_487,N_4921,N_4898);
nor UO_488 (O_488,N_4910,N_4967);
nor UO_489 (O_489,N_4579,N_4957);
and UO_490 (O_490,N_4847,N_4530);
xor UO_491 (O_491,N_4572,N_4662);
or UO_492 (O_492,N_4903,N_4604);
and UO_493 (O_493,N_4820,N_4658);
and UO_494 (O_494,N_4716,N_4794);
or UO_495 (O_495,N_4607,N_4631);
and UO_496 (O_496,N_4509,N_4961);
nand UO_497 (O_497,N_4684,N_4545);
or UO_498 (O_498,N_4750,N_4736);
and UO_499 (O_499,N_4759,N_4873);
nand UO_500 (O_500,N_4663,N_4557);
nor UO_501 (O_501,N_4685,N_4801);
xnor UO_502 (O_502,N_4816,N_4539);
and UO_503 (O_503,N_4536,N_4732);
and UO_504 (O_504,N_4825,N_4517);
nor UO_505 (O_505,N_4623,N_4896);
xnor UO_506 (O_506,N_4501,N_4817);
nor UO_507 (O_507,N_4969,N_4713);
or UO_508 (O_508,N_4623,N_4845);
xnor UO_509 (O_509,N_4667,N_4816);
xor UO_510 (O_510,N_4968,N_4770);
nand UO_511 (O_511,N_4622,N_4897);
and UO_512 (O_512,N_4835,N_4849);
or UO_513 (O_513,N_4746,N_4602);
xor UO_514 (O_514,N_4672,N_4801);
nor UO_515 (O_515,N_4847,N_4840);
or UO_516 (O_516,N_4592,N_4957);
nand UO_517 (O_517,N_4972,N_4583);
xnor UO_518 (O_518,N_4567,N_4695);
and UO_519 (O_519,N_4603,N_4727);
and UO_520 (O_520,N_4699,N_4716);
or UO_521 (O_521,N_4792,N_4919);
and UO_522 (O_522,N_4630,N_4567);
xor UO_523 (O_523,N_4573,N_4654);
xor UO_524 (O_524,N_4716,N_4534);
nor UO_525 (O_525,N_4794,N_4790);
and UO_526 (O_526,N_4604,N_4551);
nor UO_527 (O_527,N_4531,N_4677);
xor UO_528 (O_528,N_4507,N_4889);
nand UO_529 (O_529,N_4682,N_4743);
nor UO_530 (O_530,N_4565,N_4705);
nand UO_531 (O_531,N_4587,N_4550);
nor UO_532 (O_532,N_4800,N_4892);
nor UO_533 (O_533,N_4724,N_4564);
xnor UO_534 (O_534,N_4894,N_4529);
nor UO_535 (O_535,N_4515,N_4770);
nand UO_536 (O_536,N_4665,N_4945);
nor UO_537 (O_537,N_4892,N_4844);
nand UO_538 (O_538,N_4949,N_4618);
or UO_539 (O_539,N_4997,N_4687);
nand UO_540 (O_540,N_4959,N_4505);
nand UO_541 (O_541,N_4889,N_4823);
nand UO_542 (O_542,N_4795,N_4988);
nor UO_543 (O_543,N_4671,N_4833);
or UO_544 (O_544,N_4552,N_4501);
or UO_545 (O_545,N_4622,N_4831);
nand UO_546 (O_546,N_4835,N_4938);
nor UO_547 (O_547,N_4823,N_4642);
nor UO_548 (O_548,N_4828,N_4701);
xnor UO_549 (O_549,N_4782,N_4960);
xnor UO_550 (O_550,N_4747,N_4918);
nand UO_551 (O_551,N_4582,N_4533);
nor UO_552 (O_552,N_4784,N_4939);
nand UO_553 (O_553,N_4689,N_4927);
xnor UO_554 (O_554,N_4817,N_4608);
or UO_555 (O_555,N_4671,N_4755);
nor UO_556 (O_556,N_4953,N_4672);
or UO_557 (O_557,N_4540,N_4822);
xnor UO_558 (O_558,N_4695,N_4786);
nor UO_559 (O_559,N_4998,N_4638);
or UO_560 (O_560,N_4667,N_4894);
nor UO_561 (O_561,N_4924,N_4502);
nand UO_562 (O_562,N_4662,N_4811);
and UO_563 (O_563,N_4954,N_4734);
nor UO_564 (O_564,N_4581,N_4682);
xor UO_565 (O_565,N_4772,N_4784);
or UO_566 (O_566,N_4566,N_4709);
nand UO_567 (O_567,N_4590,N_4528);
and UO_568 (O_568,N_4658,N_4903);
xnor UO_569 (O_569,N_4753,N_4583);
nor UO_570 (O_570,N_4769,N_4612);
nor UO_571 (O_571,N_4816,N_4959);
or UO_572 (O_572,N_4858,N_4966);
and UO_573 (O_573,N_4746,N_4730);
xnor UO_574 (O_574,N_4854,N_4574);
or UO_575 (O_575,N_4572,N_4871);
nor UO_576 (O_576,N_4981,N_4524);
and UO_577 (O_577,N_4567,N_4635);
nor UO_578 (O_578,N_4740,N_4640);
or UO_579 (O_579,N_4730,N_4963);
nor UO_580 (O_580,N_4846,N_4605);
and UO_581 (O_581,N_4689,N_4743);
xor UO_582 (O_582,N_4523,N_4668);
or UO_583 (O_583,N_4875,N_4903);
nor UO_584 (O_584,N_4528,N_4677);
and UO_585 (O_585,N_4876,N_4957);
nor UO_586 (O_586,N_4797,N_4638);
nand UO_587 (O_587,N_4824,N_4899);
nand UO_588 (O_588,N_4998,N_4805);
xor UO_589 (O_589,N_4749,N_4501);
xor UO_590 (O_590,N_4750,N_4709);
or UO_591 (O_591,N_4773,N_4692);
xor UO_592 (O_592,N_4979,N_4959);
and UO_593 (O_593,N_4883,N_4788);
nor UO_594 (O_594,N_4599,N_4909);
nand UO_595 (O_595,N_4796,N_4634);
and UO_596 (O_596,N_4627,N_4514);
xnor UO_597 (O_597,N_4750,N_4866);
and UO_598 (O_598,N_4849,N_4571);
or UO_599 (O_599,N_4863,N_4577);
nand UO_600 (O_600,N_4749,N_4946);
xor UO_601 (O_601,N_4818,N_4658);
nand UO_602 (O_602,N_4669,N_4889);
xnor UO_603 (O_603,N_4869,N_4600);
nor UO_604 (O_604,N_4800,N_4684);
nand UO_605 (O_605,N_4782,N_4929);
xor UO_606 (O_606,N_4585,N_4946);
and UO_607 (O_607,N_4763,N_4854);
nand UO_608 (O_608,N_4560,N_4986);
nand UO_609 (O_609,N_4787,N_4973);
nand UO_610 (O_610,N_4725,N_4957);
or UO_611 (O_611,N_4907,N_4928);
nor UO_612 (O_612,N_4905,N_4793);
nor UO_613 (O_613,N_4752,N_4533);
xor UO_614 (O_614,N_4551,N_4726);
or UO_615 (O_615,N_4731,N_4940);
nor UO_616 (O_616,N_4741,N_4752);
and UO_617 (O_617,N_4896,N_4966);
and UO_618 (O_618,N_4924,N_4645);
and UO_619 (O_619,N_4740,N_4900);
xnor UO_620 (O_620,N_4815,N_4819);
or UO_621 (O_621,N_4758,N_4858);
and UO_622 (O_622,N_4515,N_4858);
xnor UO_623 (O_623,N_4515,N_4974);
or UO_624 (O_624,N_4717,N_4653);
and UO_625 (O_625,N_4705,N_4550);
nand UO_626 (O_626,N_4652,N_4510);
nor UO_627 (O_627,N_4957,N_4583);
or UO_628 (O_628,N_4521,N_4833);
and UO_629 (O_629,N_4649,N_4591);
nor UO_630 (O_630,N_4527,N_4686);
or UO_631 (O_631,N_4739,N_4785);
or UO_632 (O_632,N_4873,N_4519);
and UO_633 (O_633,N_4940,N_4796);
or UO_634 (O_634,N_4862,N_4994);
nand UO_635 (O_635,N_4506,N_4753);
and UO_636 (O_636,N_4784,N_4501);
and UO_637 (O_637,N_4773,N_4945);
or UO_638 (O_638,N_4735,N_4633);
and UO_639 (O_639,N_4540,N_4898);
or UO_640 (O_640,N_4582,N_4915);
and UO_641 (O_641,N_4633,N_4946);
or UO_642 (O_642,N_4646,N_4691);
and UO_643 (O_643,N_4786,N_4897);
nor UO_644 (O_644,N_4594,N_4892);
nand UO_645 (O_645,N_4509,N_4698);
nor UO_646 (O_646,N_4986,N_4766);
and UO_647 (O_647,N_4961,N_4584);
xnor UO_648 (O_648,N_4812,N_4568);
and UO_649 (O_649,N_4937,N_4806);
nor UO_650 (O_650,N_4845,N_4722);
and UO_651 (O_651,N_4930,N_4602);
or UO_652 (O_652,N_4651,N_4824);
nand UO_653 (O_653,N_4833,N_4921);
and UO_654 (O_654,N_4738,N_4600);
and UO_655 (O_655,N_4757,N_4861);
nor UO_656 (O_656,N_4927,N_4760);
or UO_657 (O_657,N_4703,N_4901);
nand UO_658 (O_658,N_4820,N_4643);
xnor UO_659 (O_659,N_4581,N_4837);
or UO_660 (O_660,N_4692,N_4976);
nand UO_661 (O_661,N_4692,N_4838);
nor UO_662 (O_662,N_4741,N_4888);
nand UO_663 (O_663,N_4727,N_4786);
or UO_664 (O_664,N_4810,N_4792);
nand UO_665 (O_665,N_4557,N_4612);
xor UO_666 (O_666,N_4543,N_4878);
nand UO_667 (O_667,N_4517,N_4849);
or UO_668 (O_668,N_4873,N_4814);
nand UO_669 (O_669,N_4685,N_4631);
or UO_670 (O_670,N_4903,N_4665);
nand UO_671 (O_671,N_4536,N_4702);
nand UO_672 (O_672,N_4650,N_4974);
nand UO_673 (O_673,N_4717,N_4631);
xor UO_674 (O_674,N_4720,N_4917);
or UO_675 (O_675,N_4592,N_4899);
and UO_676 (O_676,N_4568,N_4728);
and UO_677 (O_677,N_4991,N_4903);
nor UO_678 (O_678,N_4994,N_4610);
or UO_679 (O_679,N_4984,N_4850);
and UO_680 (O_680,N_4576,N_4503);
and UO_681 (O_681,N_4721,N_4935);
or UO_682 (O_682,N_4744,N_4747);
nor UO_683 (O_683,N_4700,N_4996);
or UO_684 (O_684,N_4975,N_4583);
nor UO_685 (O_685,N_4969,N_4503);
or UO_686 (O_686,N_4943,N_4639);
and UO_687 (O_687,N_4632,N_4711);
or UO_688 (O_688,N_4585,N_4625);
and UO_689 (O_689,N_4630,N_4575);
nand UO_690 (O_690,N_4553,N_4699);
and UO_691 (O_691,N_4615,N_4640);
nor UO_692 (O_692,N_4974,N_4857);
and UO_693 (O_693,N_4549,N_4667);
or UO_694 (O_694,N_4922,N_4730);
and UO_695 (O_695,N_4758,N_4888);
xor UO_696 (O_696,N_4659,N_4792);
and UO_697 (O_697,N_4978,N_4568);
xor UO_698 (O_698,N_4799,N_4779);
nor UO_699 (O_699,N_4554,N_4797);
or UO_700 (O_700,N_4815,N_4990);
nand UO_701 (O_701,N_4658,N_4971);
xor UO_702 (O_702,N_4588,N_4894);
xnor UO_703 (O_703,N_4579,N_4688);
or UO_704 (O_704,N_4509,N_4612);
nor UO_705 (O_705,N_4716,N_4999);
or UO_706 (O_706,N_4782,N_4771);
nand UO_707 (O_707,N_4741,N_4514);
xnor UO_708 (O_708,N_4591,N_4968);
or UO_709 (O_709,N_4520,N_4807);
or UO_710 (O_710,N_4669,N_4973);
and UO_711 (O_711,N_4714,N_4642);
and UO_712 (O_712,N_4543,N_4581);
xnor UO_713 (O_713,N_4693,N_4586);
or UO_714 (O_714,N_4727,N_4719);
or UO_715 (O_715,N_4661,N_4594);
xor UO_716 (O_716,N_4834,N_4843);
nand UO_717 (O_717,N_4930,N_4910);
xor UO_718 (O_718,N_4522,N_4724);
and UO_719 (O_719,N_4951,N_4555);
or UO_720 (O_720,N_4827,N_4532);
or UO_721 (O_721,N_4742,N_4826);
and UO_722 (O_722,N_4691,N_4605);
or UO_723 (O_723,N_4602,N_4794);
and UO_724 (O_724,N_4641,N_4879);
and UO_725 (O_725,N_4658,N_4861);
nor UO_726 (O_726,N_4857,N_4956);
nand UO_727 (O_727,N_4872,N_4567);
xnor UO_728 (O_728,N_4637,N_4562);
and UO_729 (O_729,N_4913,N_4743);
nand UO_730 (O_730,N_4666,N_4965);
or UO_731 (O_731,N_4514,N_4868);
xnor UO_732 (O_732,N_4869,N_4506);
nor UO_733 (O_733,N_4517,N_4688);
or UO_734 (O_734,N_4605,N_4891);
or UO_735 (O_735,N_4641,N_4750);
nor UO_736 (O_736,N_4770,N_4702);
nor UO_737 (O_737,N_4547,N_4587);
or UO_738 (O_738,N_4948,N_4705);
nor UO_739 (O_739,N_4744,N_4981);
and UO_740 (O_740,N_4697,N_4827);
or UO_741 (O_741,N_4805,N_4707);
nor UO_742 (O_742,N_4681,N_4560);
xnor UO_743 (O_743,N_4818,N_4650);
nand UO_744 (O_744,N_4720,N_4550);
or UO_745 (O_745,N_4991,N_4840);
and UO_746 (O_746,N_4602,N_4772);
xnor UO_747 (O_747,N_4509,N_4975);
and UO_748 (O_748,N_4534,N_4620);
and UO_749 (O_749,N_4871,N_4531);
nor UO_750 (O_750,N_4996,N_4749);
nor UO_751 (O_751,N_4766,N_4664);
nor UO_752 (O_752,N_4976,N_4839);
xor UO_753 (O_753,N_4835,N_4733);
nor UO_754 (O_754,N_4569,N_4996);
nand UO_755 (O_755,N_4849,N_4750);
nor UO_756 (O_756,N_4975,N_4780);
xnor UO_757 (O_757,N_4942,N_4889);
nor UO_758 (O_758,N_4557,N_4833);
nor UO_759 (O_759,N_4612,N_4653);
nand UO_760 (O_760,N_4633,N_4849);
and UO_761 (O_761,N_4736,N_4954);
nand UO_762 (O_762,N_4851,N_4893);
nor UO_763 (O_763,N_4577,N_4722);
nand UO_764 (O_764,N_4896,N_4812);
nand UO_765 (O_765,N_4732,N_4793);
or UO_766 (O_766,N_4964,N_4793);
or UO_767 (O_767,N_4947,N_4594);
nor UO_768 (O_768,N_4619,N_4511);
nor UO_769 (O_769,N_4781,N_4768);
xor UO_770 (O_770,N_4589,N_4759);
xnor UO_771 (O_771,N_4507,N_4796);
and UO_772 (O_772,N_4512,N_4960);
nand UO_773 (O_773,N_4939,N_4865);
nor UO_774 (O_774,N_4594,N_4823);
or UO_775 (O_775,N_4958,N_4837);
or UO_776 (O_776,N_4910,N_4854);
or UO_777 (O_777,N_4617,N_4818);
xnor UO_778 (O_778,N_4574,N_4575);
nor UO_779 (O_779,N_4750,N_4692);
nor UO_780 (O_780,N_4777,N_4551);
nand UO_781 (O_781,N_4616,N_4892);
nand UO_782 (O_782,N_4564,N_4615);
and UO_783 (O_783,N_4624,N_4618);
nand UO_784 (O_784,N_4886,N_4764);
nor UO_785 (O_785,N_4573,N_4583);
and UO_786 (O_786,N_4673,N_4627);
or UO_787 (O_787,N_4966,N_4580);
and UO_788 (O_788,N_4942,N_4754);
and UO_789 (O_789,N_4968,N_4586);
xor UO_790 (O_790,N_4845,N_4869);
nand UO_791 (O_791,N_4850,N_4532);
nand UO_792 (O_792,N_4533,N_4509);
xor UO_793 (O_793,N_4991,N_4757);
or UO_794 (O_794,N_4760,N_4677);
or UO_795 (O_795,N_4768,N_4969);
xor UO_796 (O_796,N_4681,N_4624);
and UO_797 (O_797,N_4979,N_4837);
nand UO_798 (O_798,N_4512,N_4605);
and UO_799 (O_799,N_4760,N_4934);
or UO_800 (O_800,N_4707,N_4745);
and UO_801 (O_801,N_4879,N_4747);
or UO_802 (O_802,N_4992,N_4870);
xor UO_803 (O_803,N_4553,N_4908);
nor UO_804 (O_804,N_4716,N_4909);
xor UO_805 (O_805,N_4857,N_4654);
nand UO_806 (O_806,N_4864,N_4879);
and UO_807 (O_807,N_4975,N_4627);
and UO_808 (O_808,N_4639,N_4989);
nor UO_809 (O_809,N_4979,N_4539);
or UO_810 (O_810,N_4642,N_4663);
xor UO_811 (O_811,N_4957,N_4640);
and UO_812 (O_812,N_4621,N_4508);
nor UO_813 (O_813,N_4849,N_4968);
and UO_814 (O_814,N_4799,N_4762);
xor UO_815 (O_815,N_4749,N_4736);
xor UO_816 (O_816,N_4578,N_4597);
and UO_817 (O_817,N_4556,N_4925);
nor UO_818 (O_818,N_4517,N_4607);
xnor UO_819 (O_819,N_4521,N_4676);
or UO_820 (O_820,N_4567,N_4738);
and UO_821 (O_821,N_4872,N_4960);
nand UO_822 (O_822,N_4963,N_4747);
nor UO_823 (O_823,N_4851,N_4843);
and UO_824 (O_824,N_4853,N_4503);
nor UO_825 (O_825,N_4840,N_4579);
nand UO_826 (O_826,N_4796,N_4811);
nand UO_827 (O_827,N_4947,N_4521);
and UO_828 (O_828,N_4627,N_4899);
nand UO_829 (O_829,N_4848,N_4798);
and UO_830 (O_830,N_4580,N_4521);
xnor UO_831 (O_831,N_4629,N_4513);
or UO_832 (O_832,N_4500,N_4664);
and UO_833 (O_833,N_4891,N_4595);
xor UO_834 (O_834,N_4851,N_4732);
nand UO_835 (O_835,N_4643,N_4920);
and UO_836 (O_836,N_4567,N_4704);
or UO_837 (O_837,N_4542,N_4936);
xnor UO_838 (O_838,N_4856,N_4824);
or UO_839 (O_839,N_4571,N_4822);
nand UO_840 (O_840,N_4683,N_4856);
nor UO_841 (O_841,N_4757,N_4598);
nor UO_842 (O_842,N_4617,N_4910);
xor UO_843 (O_843,N_4515,N_4917);
or UO_844 (O_844,N_4967,N_4959);
nand UO_845 (O_845,N_4869,N_4727);
nand UO_846 (O_846,N_4687,N_4757);
and UO_847 (O_847,N_4693,N_4998);
xor UO_848 (O_848,N_4698,N_4704);
xnor UO_849 (O_849,N_4751,N_4615);
or UO_850 (O_850,N_4729,N_4521);
and UO_851 (O_851,N_4566,N_4795);
xnor UO_852 (O_852,N_4646,N_4550);
nand UO_853 (O_853,N_4934,N_4962);
nand UO_854 (O_854,N_4503,N_4569);
xor UO_855 (O_855,N_4744,N_4924);
or UO_856 (O_856,N_4946,N_4777);
nand UO_857 (O_857,N_4764,N_4762);
and UO_858 (O_858,N_4941,N_4800);
or UO_859 (O_859,N_4804,N_4912);
xnor UO_860 (O_860,N_4601,N_4733);
and UO_861 (O_861,N_4857,N_4533);
or UO_862 (O_862,N_4878,N_4986);
or UO_863 (O_863,N_4981,N_4736);
nand UO_864 (O_864,N_4813,N_4609);
or UO_865 (O_865,N_4772,N_4653);
or UO_866 (O_866,N_4943,N_4530);
or UO_867 (O_867,N_4834,N_4524);
and UO_868 (O_868,N_4991,N_4786);
or UO_869 (O_869,N_4618,N_4718);
and UO_870 (O_870,N_4544,N_4512);
nor UO_871 (O_871,N_4679,N_4554);
nor UO_872 (O_872,N_4892,N_4906);
or UO_873 (O_873,N_4589,N_4876);
or UO_874 (O_874,N_4829,N_4895);
nand UO_875 (O_875,N_4946,N_4776);
or UO_876 (O_876,N_4996,N_4822);
xnor UO_877 (O_877,N_4701,N_4724);
xnor UO_878 (O_878,N_4630,N_4928);
and UO_879 (O_879,N_4783,N_4684);
or UO_880 (O_880,N_4848,N_4863);
or UO_881 (O_881,N_4689,N_4675);
nand UO_882 (O_882,N_4846,N_4703);
and UO_883 (O_883,N_4774,N_4500);
xnor UO_884 (O_884,N_4909,N_4779);
or UO_885 (O_885,N_4906,N_4618);
and UO_886 (O_886,N_4726,N_4843);
or UO_887 (O_887,N_4598,N_4875);
nand UO_888 (O_888,N_4944,N_4674);
or UO_889 (O_889,N_4693,N_4847);
nand UO_890 (O_890,N_4624,N_4570);
nor UO_891 (O_891,N_4557,N_4501);
nor UO_892 (O_892,N_4640,N_4838);
nor UO_893 (O_893,N_4648,N_4775);
nor UO_894 (O_894,N_4553,N_4745);
or UO_895 (O_895,N_4980,N_4742);
and UO_896 (O_896,N_4683,N_4726);
nor UO_897 (O_897,N_4555,N_4960);
nand UO_898 (O_898,N_4934,N_4859);
or UO_899 (O_899,N_4789,N_4858);
xor UO_900 (O_900,N_4788,N_4778);
nand UO_901 (O_901,N_4871,N_4760);
nand UO_902 (O_902,N_4935,N_4576);
and UO_903 (O_903,N_4759,N_4600);
nand UO_904 (O_904,N_4798,N_4613);
nand UO_905 (O_905,N_4834,N_4732);
nand UO_906 (O_906,N_4955,N_4756);
xor UO_907 (O_907,N_4546,N_4633);
and UO_908 (O_908,N_4655,N_4880);
nor UO_909 (O_909,N_4662,N_4614);
xnor UO_910 (O_910,N_4626,N_4789);
and UO_911 (O_911,N_4503,N_4812);
xnor UO_912 (O_912,N_4818,N_4559);
and UO_913 (O_913,N_4973,N_4561);
nor UO_914 (O_914,N_4869,N_4535);
nor UO_915 (O_915,N_4640,N_4835);
nor UO_916 (O_916,N_4806,N_4827);
nand UO_917 (O_917,N_4751,N_4960);
nand UO_918 (O_918,N_4826,N_4859);
nor UO_919 (O_919,N_4668,N_4635);
nand UO_920 (O_920,N_4546,N_4587);
nor UO_921 (O_921,N_4829,N_4989);
nor UO_922 (O_922,N_4825,N_4873);
or UO_923 (O_923,N_4722,N_4710);
nand UO_924 (O_924,N_4811,N_4729);
nor UO_925 (O_925,N_4694,N_4779);
nand UO_926 (O_926,N_4639,N_4722);
and UO_927 (O_927,N_4509,N_4758);
nor UO_928 (O_928,N_4986,N_4871);
nand UO_929 (O_929,N_4554,N_4580);
and UO_930 (O_930,N_4531,N_4565);
and UO_931 (O_931,N_4999,N_4676);
or UO_932 (O_932,N_4976,N_4891);
nor UO_933 (O_933,N_4642,N_4582);
xor UO_934 (O_934,N_4546,N_4670);
xnor UO_935 (O_935,N_4853,N_4615);
nand UO_936 (O_936,N_4832,N_4703);
xor UO_937 (O_937,N_4525,N_4661);
nor UO_938 (O_938,N_4659,N_4530);
nor UO_939 (O_939,N_4640,N_4613);
nand UO_940 (O_940,N_4705,N_4534);
or UO_941 (O_941,N_4606,N_4870);
nor UO_942 (O_942,N_4650,N_4601);
and UO_943 (O_943,N_4550,N_4559);
xnor UO_944 (O_944,N_4908,N_4923);
and UO_945 (O_945,N_4804,N_4566);
and UO_946 (O_946,N_4601,N_4992);
xor UO_947 (O_947,N_4813,N_4789);
nand UO_948 (O_948,N_4709,N_4786);
xor UO_949 (O_949,N_4970,N_4682);
nor UO_950 (O_950,N_4519,N_4982);
nor UO_951 (O_951,N_4974,N_4701);
nand UO_952 (O_952,N_4904,N_4626);
nor UO_953 (O_953,N_4890,N_4984);
nand UO_954 (O_954,N_4613,N_4946);
nand UO_955 (O_955,N_4872,N_4656);
nand UO_956 (O_956,N_4590,N_4830);
or UO_957 (O_957,N_4742,N_4510);
xnor UO_958 (O_958,N_4849,N_4891);
and UO_959 (O_959,N_4773,N_4573);
nor UO_960 (O_960,N_4847,N_4861);
and UO_961 (O_961,N_4941,N_4578);
nand UO_962 (O_962,N_4624,N_4648);
nand UO_963 (O_963,N_4790,N_4625);
and UO_964 (O_964,N_4815,N_4681);
nor UO_965 (O_965,N_4981,N_4996);
nand UO_966 (O_966,N_4891,N_4779);
nor UO_967 (O_967,N_4999,N_4753);
xor UO_968 (O_968,N_4752,N_4805);
and UO_969 (O_969,N_4637,N_4663);
or UO_970 (O_970,N_4724,N_4996);
nand UO_971 (O_971,N_4704,N_4574);
or UO_972 (O_972,N_4775,N_4695);
nand UO_973 (O_973,N_4602,N_4907);
nand UO_974 (O_974,N_4788,N_4834);
nor UO_975 (O_975,N_4848,N_4684);
or UO_976 (O_976,N_4609,N_4543);
and UO_977 (O_977,N_4906,N_4810);
xnor UO_978 (O_978,N_4778,N_4767);
and UO_979 (O_979,N_4930,N_4608);
or UO_980 (O_980,N_4898,N_4940);
nand UO_981 (O_981,N_4672,N_4548);
nand UO_982 (O_982,N_4719,N_4726);
and UO_983 (O_983,N_4860,N_4822);
and UO_984 (O_984,N_4954,N_4570);
and UO_985 (O_985,N_4777,N_4501);
xnor UO_986 (O_986,N_4836,N_4972);
or UO_987 (O_987,N_4510,N_4589);
or UO_988 (O_988,N_4713,N_4701);
and UO_989 (O_989,N_4676,N_4883);
or UO_990 (O_990,N_4937,N_4705);
nand UO_991 (O_991,N_4898,N_4846);
and UO_992 (O_992,N_4750,N_4893);
nor UO_993 (O_993,N_4561,N_4616);
and UO_994 (O_994,N_4706,N_4900);
nand UO_995 (O_995,N_4996,N_4998);
nor UO_996 (O_996,N_4590,N_4988);
nor UO_997 (O_997,N_4722,N_4657);
and UO_998 (O_998,N_4892,N_4621);
nor UO_999 (O_999,N_4555,N_4819);
endmodule