module basic_3000_30000_3500_10_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_608,In_52);
nor U1 (N_1,In_2848,In_2343);
and U2 (N_2,In_2682,In_2843);
nand U3 (N_3,In_292,In_2192);
nand U4 (N_4,In_1745,In_2536);
nand U5 (N_5,In_2052,In_1475);
or U6 (N_6,In_129,In_253);
xnor U7 (N_7,In_2406,In_2038);
xnor U8 (N_8,In_1092,In_28);
xnor U9 (N_9,In_1012,In_2508);
nor U10 (N_10,In_2598,In_540);
and U11 (N_11,In_3,In_640);
nor U12 (N_12,In_2278,In_2102);
nor U13 (N_13,In_1235,In_869);
or U14 (N_14,In_87,In_2417);
nand U15 (N_15,In_2518,In_2894);
nand U16 (N_16,In_1304,In_2451);
nand U17 (N_17,In_1287,In_128);
or U18 (N_18,In_837,In_242);
and U19 (N_19,In_1638,In_1705);
nand U20 (N_20,In_152,In_2607);
nand U21 (N_21,In_2074,In_537);
nand U22 (N_22,In_2004,In_1900);
and U23 (N_23,In_2198,In_962);
or U24 (N_24,In_2551,In_2630);
or U25 (N_25,In_2832,In_114);
nor U26 (N_26,In_2206,In_420);
and U27 (N_27,In_660,In_1898);
and U28 (N_28,In_1251,In_543);
xnor U29 (N_29,In_697,In_131);
or U30 (N_30,In_1759,In_1465);
and U31 (N_31,In_15,In_743);
xnor U32 (N_32,In_1102,In_567);
and U33 (N_33,In_2288,In_410);
nor U34 (N_34,In_1083,In_397);
nor U35 (N_35,In_388,In_1044);
or U36 (N_36,In_1780,In_1138);
nor U37 (N_37,In_2683,In_2071);
nor U38 (N_38,In_1355,In_555);
or U39 (N_39,In_429,In_744);
xor U40 (N_40,In_1764,In_2898);
nor U41 (N_41,In_447,In_463);
nand U42 (N_42,In_965,In_186);
nand U43 (N_43,In_1103,In_2575);
nor U44 (N_44,In_2538,In_2549);
or U45 (N_45,In_930,In_1207);
or U46 (N_46,In_1196,In_2594);
or U47 (N_47,In_623,In_2083);
nor U48 (N_48,In_2305,In_343);
or U49 (N_49,In_1294,In_38);
nand U50 (N_50,In_165,In_1698);
or U51 (N_51,In_589,In_2766);
xnor U52 (N_52,In_1484,In_2027);
xnor U53 (N_53,In_1988,In_2797);
xor U54 (N_54,In_1661,In_2972);
and U55 (N_55,In_2232,In_1811);
xnor U56 (N_56,In_526,In_1219);
nand U57 (N_57,In_2642,In_1527);
or U58 (N_58,In_2204,In_1299);
or U59 (N_59,In_1758,In_2907);
and U60 (N_60,In_32,In_405);
nand U61 (N_61,In_1576,In_1603);
and U62 (N_62,In_446,In_355);
and U63 (N_63,In_2916,In_1589);
nand U64 (N_64,In_2123,In_2046);
nor U65 (N_65,In_549,In_2981);
and U66 (N_66,In_2162,In_80);
and U67 (N_67,In_2474,In_1627);
nand U68 (N_68,In_278,In_1959);
and U69 (N_69,In_2971,In_2635);
xnor U70 (N_70,In_952,In_2928);
nor U71 (N_71,In_2895,In_1094);
nor U72 (N_72,In_34,In_988);
xnor U73 (N_73,In_126,In_2560);
nand U74 (N_74,In_2872,In_2869);
nand U75 (N_75,In_1806,In_195);
xor U76 (N_76,In_1167,In_286);
and U77 (N_77,In_1282,In_2116);
nand U78 (N_78,In_1503,In_307);
or U79 (N_79,In_2180,In_935);
nand U80 (N_80,In_839,In_448);
and U81 (N_81,In_1075,In_629);
xnor U82 (N_82,In_856,In_654);
and U83 (N_83,In_2571,In_2314);
xor U84 (N_84,In_1420,In_2212);
and U85 (N_85,In_320,In_1542);
nor U86 (N_86,In_2859,In_2727);
nand U87 (N_87,In_1560,In_1699);
or U88 (N_88,In_2955,In_1701);
or U89 (N_89,In_1155,In_2721);
or U90 (N_90,In_298,In_301);
nand U91 (N_91,In_1781,In_2193);
and U92 (N_92,In_634,In_1091);
nand U93 (N_93,In_2262,In_742);
xor U94 (N_94,In_1424,In_846);
xor U95 (N_95,In_1752,In_2735);
or U96 (N_96,In_2320,In_668);
nor U97 (N_97,In_2374,In_518);
and U98 (N_98,In_1021,In_2325);
nand U99 (N_99,In_2017,In_875);
or U100 (N_100,In_805,In_2281);
xor U101 (N_101,In_135,In_1966);
nand U102 (N_102,In_973,In_2677);
and U103 (N_103,In_1876,In_1389);
nand U104 (N_104,In_185,In_1418);
or U105 (N_105,In_490,In_1053);
xor U106 (N_106,In_525,In_917);
nor U107 (N_107,In_542,In_949);
nor U108 (N_108,In_1778,In_2029);
nand U109 (N_109,In_1857,In_529);
and U110 (N_110,In_519,In_2650);
xor U111 (N_111,In_1894,In_2030);
nor U112 (N_112,In_1881,In_2962);
or U113 (N_113,In_1830,In_2513);
and U114 (N_114,In_1571,In_2725);
or U115 (N_115,In_256,In_1556);
xor U116 (N_116,In_1800,In_2941);
nor U117 (N_117,In_2203,In_2758);
xor U118 (N_118,In_1559,In_2930);
or U119 (N_119,In_2499,In_2426);
and U120 (N_120,In_2570,In_2681);
nor U121 (N_121,In_1283,In_1112);
nand U122 (N_122,In_2590,In_1303);
or U123 (N_123,In_802,In_2656);
nand U124 (N_124,In_2864,In_581);
nor U125 (N_125,In_1650,In_1869);
or U126 (N_126,In_2333,In_2459);
nor U127 (N_127,In_16,In_819);
nor U128 (N_128,In_2697,In_1085);
nand U129 (N_129,In_572,In_348);
nand U130 (N_130,In_427,In_2121);
and U131 (N_131,In_808,In_1770);
nand U132 (N_132,In_622,In_1851);
nor U133 (N_133,In_2479,In_1909);
nor U134 (N_134,In_512,In_2960);
nand U135 (N_135,In_1049,In_645);
xor U136 (N_136,In_2050,In_104);
or U137 (N_137,In_67,In_167);
xor U138 (N_138,In_2384,In_1105);
and U139 (N_139,In_1651,In_360);
and U140 (N_140,In_1911,In_643);
nand U141 (N_141,In_2435,In_1330);
xor U142 (N_142,In_539,In_2668);
nor U143 (N_143,In_803,In_1170);
and U144 (N_144,In_2803,In_1314);
nand U145 (N_145,In_2833,In_2628);
and U146 (N_146,In_1369,In_2040);
nor U147 (N_147,In_306,In_2574);
and U148 (N_148,In_748,In_842);
nor U149 (N_149,In_1662,In_2910);
nor U150 (N_150,In_302,In_174);
nor U151 (N_151,In_50,In_2126);
xor U152 (N_152,In_2866,In_73);
nor U153 (N_153,In_2937,In_1610);
nand U154 (N_154,In_1042,In_1288);
nand U155 (N_155,In_2863,In_996);
nor U156 (N_156,In_1835,In_2517);
or U157 (N_157,In_2616,In_1690);
and U158 (N_158,In_2090,In_905);
or U159 (N_159,In_788,In_1691);
nor U160 (N_160,In_250,In_1244);
and U161 (N_161,In_2063,In_433);
or U162 (N_162,In_1865,In_644);
xor U163 (N_163,In_1351,In_2425);
and U164 (N_164,In_1118,In_800);
nand U165 (N_165,In_107,In_797);
nor U166 (N_166,In_1510,In_2658);
nand U167 (N_167,In_1718,In_477);
xor U168 (N_168,In_254,In_1216);
or U169 (N_169,In_2336,In_1229);
or U170 (N_170,In_127,In_828);
nand U171 (N_171,In_557,In_2068);
nor U172 (N_172,In_456,In_1407);
nand U173 (N_173,In_245,In_662);
nand U174 (N_174,In_2839,In_2334);
and U175 (N_175,In_2316,In_2657);
nand U176 (N_176,In_2057,In_2362);
and U177 (N_177,In_49,In_657);
nand U178 (N_178,In_934,In_1144);
nand U179 (N_179,In_2613,In_786);
xnor U180 (N_180,In_288,In_471);
nor U181 (N_181,In_1967,In_173);
xor U182 (N_182,In_1276,In_2034);
xnor U183 (N_183,In_78,In_179);
nand U184 (N_184,In_1408,In_1957);
or U185 (N_185,In_1686,In_1008);
nand U186 (N_186,In_1061,In_1514);
or U187 (N_187,In_1300,In_926);
nor U188 (N_188,In_494,In_1179);
and U189 (N_189,In_1356,In_2619);
and U190 (N_190,In_1275,In_2825);
or U191 (N_191,In_208,In_403);
and U192 (N_192,In_690,In_637);
nor U193 (N_193,In_508,In_1723);
and U194 (N_194,In_1913,In_2404);
nor U195 (N_195,In_1625,In_2263);
nand U196 (N_196,In_2395,In_833);
or U197 (N_197,In_1297,In_1863);
nand U198 (N_198,In_2828,In_1187);
nand U199 (N_199,In_2265,In_19);
xnor U200 (N_200,In_1847,In_2606);
nand U201 (N_201,In_2147,In_2414);
nor U202 (N_202,In_2544,In_2423);
nor U203 (N_203,In_1469,In_2678);
xnor U204 (N_204,In_338,In_514);
nand U205 (N_205,In_100,In_2500);
nand U206 (N_206,In_145,In_1132);
xor U207 (N_207,In_2101,In_1979);
xnor U208 (N_208,In_1535,In_2372);
or U209 (N_209,In_2795,In_2502);
nor U210 (N_210,In_492,In_2956);
nand U211 (N_211,In_1995,In_773);
or U212 (N_212,In_1726,In_2900);
and U213 (N_213,In_2279,In_2850);
xnor U214 (N_214,In_2891,In_2009);
nand U215 (N_215,In_2511,In_215);
nor U216 (N_216,In_2061,In_878);
and U217 (N_217,In_1230,In_264);
nand U218 (N_218,In_491,In_202);
nand U219 (N_219,In_2586,In_462);
nor U220 (N_220,In_1551,In_1357);
and U221 (N_221,In_2951,In_1016);
nor U222 (N_222,In_451,In_2327);
and U223 (N_223,In_455,In_896);
xor U224 (N_224,In_2533,In_1277);
or U225 (N_225,In_2213,In_2318);
or U226 (N_226,In_2383,In_801);
or U227 (N_227,In_2566,In_982);
xnor U228 (N_228,In_1816,In_2564);
nand U229 (N_229,In_1078,In_280);
xor U230 (N_230,In_575,In_1512);
xnor U231 (N_231,In_1295,In_231);
and U232 (N_232,In_1626,In_1520);
or U233 (N_233,In_1779,In_1984);
xor U234 (N_234,In_1433,In_130);
nand U235 (N_235,In_864,In_1963);
nand U236 (N_236,In_1710,In_2645);
nand U237 (N_237,In_2600,In_2707);
and U238 (N_238,In_1896,In_2800);
nand U239 (N_239,In_554,In_1978);
nor U240 (N_240,In_628,In_719);
xor U241 (N_241,In_597,In_1255);
and U242 (N_242,In_1753,In_1573);
xnor U243 (N_243,In_260,In_2983);
nand U244 (N_244,In_1647,In_2664);
and U245 (N_245,In_2494,In_2750);
and U246 (N_246,In_614,In_586);
xnor U247 (N_247,In_1635,In_733);
nand U248 (N_248,In_1598,In_2802);
or U249 (N_249,In_340,In_1343);
and U250 (N_250,In_2182,In_1073);
nor U251 (N_251,In_1126,In_1954);
and U252 (N_252,In_2249,In_2632);
or U253 (N_253,In_2884,In_2641);
and U254 (N_254,In_585,In_2779);
or U255 (N_255,In_672,In_2969);
nand U256 (N_256,In_2274,In_386);
nor U257 (N_257,In_2811,In_2610);
and U258 (N_258,In_787,In_2103);
nand U259 (N_259,In_170,In_204);
or U260 (N_260,In_2453,In_2836);
xnor U261 (N_261,In_40,In_2798);
and U262 (N_262,In_761,In_1256);
xor U263 (N_263,In_2056,In_545);
nand U264 (N_264,In_2791,In_578);
or U265 (N_265,In_793,In_2088);
and U266 (N_266,In_1501,In_576);
and U267 (N_267,In_1172,In_794);
nor U268 (N_268,In_734,In_2926);
nand U269 (N_269,In_1956,In_872);
or U270 (N_270,In_2873,In_62);
xor U271 (N_271,In_1413,In_2749);
xor U272 (N_272,In_2243,In_756);
and U273 (N_273,In_2411,In_1768);
nor U274 (N_274,In_1225,In_1458);
nor U275 (N_275,In_346,In_2447);
nor U276 (N_276,In_45,In_238);
and U277 (N_277,In_2143,In_1428);
and U278 (N_278,In_2757,In_1238);
or U279 (N_279,In_2122,In_2692);
xnor U280 (N_280,In_2420,In_2060);
or U281 (N_281,In_2695,In_2136);
nand U282 (N_282,In_979,In_1495);
nor U283 (N_283,In_826,In_1301);
nand U284 (N_284,In_992,In_978);
or U285 (N_285,In_1050,In_1921);
nand U286 (N_286,In_2977,In_975);
and U287 (N_287,In_2118,In_841);
or U288 (N_288,In_2033,In_2099);
xor U289 (N_289,In_1064,In_123);
or U290 (N_290,In_956,In_1532);
xnor U291 (N_291,In_2441,In_1862);
xnor U292 (N_292,In_550,In_1613);
xnor U293 (N_293,In_1245,In_497);
nand U294 (N_294,In_2301,In_387);
nor U295 (N_295,In_1853,In_2064);
nor U296 (N_296,In_2280,In_2031);
or U297 (N_297,In_1115,In_2671);
nand U298 (N_298,In_2106,In_2312);
or U299 (N_299,In_2706,In_1237);
xor U300 (N_300,In_1586,In_2845);
nor U301 (N_301,In_2261,In_2821);
nor U302 (N_302,In_2649,In_2646);
nand U303 (N_303,In_1893,In_893);
xnor U304 (N_304,In_619,In_860);
nor U305 (N_305,In_770,In_2541);
nor U306 (N_306,In_698,In_2504);
nand U307 (N_307,In_1374,In_1926);
nor U308 (N_308,In_1574,In_311);
xor U309 (N_309,In_1421,In_2174);
and U310 (N_310,In_579,In_1797);
nor U311 (N_311,In_2818,In_2231);
or U312 (N_312,In_1649,In_300);
and U313 (N_313,In_2718,In_2455);
xor U314 (N_314,In_1941,In_2584);
nand U315 (N_315,In_323,In_1051);
or U316 (N_316,In_2273,In_2939);
nor U317 (N_317,In_2719,In_1708);
and U318 (N_318,In_440,In_1695);
nor U319 (N_319,In_488,In_1669);
nand U320 (N_320,In_653,In_20);
nand U321 (N_321,In_580,In_1606);
nor U322 (N_322,In_641,In_769);
nor U323 (N_323,In_1620,In_1526);
or U324 (N_324,In_2108,In_1224);
and U325 (N_325,In_1034,In_99);
and U326 (N_326,In_1702,In_482);
or U327 (N_327,In_1292,In_2705);
or U328 (N_328,In_2660,In_857);
and U329 (N_329,In_1942,In_2189);
nand U330 (N_330,In_1960,In_331);
nor U331 (N_331,In_1788,In_2440);
nor U332 (N_332,In_1386,In_2558);
or U333 (N_333,In_2633,In_2239);
or U334 (N_334,In_274,In_725);
and U335 (N_335,In_468,In_1633);
xnor U336 (N_336,In_1339,In_2117);
xnor U337 (N_337,In_1192,In_2188);
nand U338 (N_338,In_959,In_618);
xnor U339 (N_339,In_2378,In_2742);
xor U340 (N_340,In_2653,In_1767);
or U341 (N_341,In_796,In_2562);
nand U342 (N_342,In_758,In_443);
xor U343 (N_343,In_1871,In_1757);
nand U344 (N_344,In_1082,In_1741);
nor U345 (N_345,In_785,In_520);
or U346 (N_346,In_1221,In_196);
xor U347 (N_347,In_381,In_2892);
or U348 (N_348,In_1246,In_2018);
nand U349 (N_349,In_1210,In_92);
or U350 (N_350,In_1630,In_275);
or U351 (N_351,In_141,In_1490);
nand U352 (N_352,In_2950,In_2287);
xnor U353 (N_353,In_2065,In_1149);
and U354 (N_354,In_1657,In_2023);
xnor U355 (N_355,In_2732,In_1499);
or U356 (N_356,In_1372,In_1150);
and U357 (N_357,In_1266,In_2556);
nor U358 (N_358,In_1344,In_1880);
xnor U359 (N_359,In_776,In_1859);
nand U360 (N_360,In_66,In_983);
nor U361 (N_361,In_188,In_664);
nor U362 (N_362,In_2792,In_2043);
nor U363 (N_363,In_2585,In_1837);
nand U364 (N_364,In_315,In_953);
xnor U365 (N_365,In_849,In_2882);
or U366 (N_366,In_2861,In_2953);
and U367 (N_367,In_1823,In_2942);
nand U368 (N_368,In_2991,In_2840);
and U369 (N_369,In_1310,In_2929);
nor U370 (N_370,In_1243,In_316);
xor U371 (N_371,In_824,In_898);
or U372 (N_372,In_2858,In_705);
and U373 (N_373,In_639,In_2002);
and U374 (N_374,In_2819,In_2183);
nand U375 (N_375,In_2925,In_122);
or U376 (N_376,In_333,In_884);
nand U377 (N_377,In_84,In_1493);
nand U378 (N_378,In_1687,In_564);
or U379 (N_379,In_2380,In_2238);
nor U380 (N_380,In_1653,In_43);
or U381 (N_381,In_2669,In_2125);
or U382 (N_382,In_1572,In_2466);
or U383 (N_383,In_1383,In_1366);
nor U384 (N_384,In_2724,In_1990);
and U385 (N_385,In_1041,In_299);
xnor U386 (N_386,In_1636,In_714);
nand U387 (N_387,In_1872,In_2006);
or U388 (N_388,In_2460,In_1089);
xnor U389 (N_389,In_913,In_2392);
nor U390 (N_390,In_2245,In_2734);
or U391 (N_391,In_265,In_1482);
or U392 (N_392,In_1934,In_2659);
xor U393 (N_393,In_2992,In_217);
and U394 (N_394,In_1460,In_2089);
xnor U395 (N_395,In_2949,In_604);
or U396 (N_396,In_2651,In_2485);
nand U397 (N_397,In_1066,In_506);
nand U398 (N_398,In_2979,In_453);
nor U399 (N_399,In_2783,In_2297);
nor U400 (N_400,In_1498,In_434);
nand U401 (N_401,In_859,In_2568);
xor U402 (N_402,In_58,In_1239);
xor U403 (N_403,In_817,In_2230);
nor U404 (N_404,In_2717,In_2473);
nor U405 (N_405,In_2587,In_1202);
nor U406 (N_406,In_1592,In_2654);
xnor U407 (N_407,In_1511,In_738);
nand U408 (N_408,In_1810,In_2247);
and U409 (N_409,In_2005,In_544);
xor U410 (N_410,In_351,In_2207);
xor U411 (N_411,In_1766,In_1733);
nand U412 (N_412,In_1973,In_2067);
nor U413 (N_413,In_1867,In_2912);
or U414 (N_414,In_2744,In_2110);
nand U415 (N_415,In_432,In_1109);
nand U416 (N_416,In_1378,In_2923);
nand U417 (N_417,In_2529,In_224);
or U418 (N_418,In_2290,In_1380);
and U419 (N_419,In_1284,In_1644);
and U420 (N_420,In_1792,In_2532);
and U421 (N_421,In_1502,In_1664);
nor U422 (N_422,In_2581,In_2856);
and U423 (N_423,In_687,In_1203);
xnor U424 (N_424,In_374,In_2772);
nor U425 (N_425,In_693,In_1208);
and U426 (N_426,In_1481,In_228);
nor U427 (N_427,In_1595,In_772);
nand U428 (N_428,In_1147,In_1432);
nand U429 (N_429,In_1516,In_2405);
and U430 (N_430,In_454,In_1152);
or U431 (N_431,In_2728,In_1974);
nand U432 (N_432,In_1795,In_2258);
or U433 (N_433,In_2543,In_2793);
nand U434 (N_434,In_2927,In_1176);
nand U435 (N_435,In_2531,In_30);
or U436 (N_436,In_1060,In_2947);
nand U437 (N_437,In_1370,In_1430);
nor U438 (N_438,In_1782,In_2629);
nor U439 (N_439,In_2233,In_1404);
nor U440 (N_440,In_2255,In_2346);
nand U441 (N_441,In_312,In_1685);
and U442 (N_442,In_108,In_44);
or U443 (N_443,In_861,In_1528);
or U444 (N_444,In_2070,In_1204);
nand U445 (N_445,In_2191,In_1769);
nor U446 (N_446,In_23,In_1254);
xor U447 (N_447,In_460,In_1437);
and U448 (N_448,In_1477,In_1807);
nand U449 (N_449,In_584,In_1897);
nand U450 (N_450,In_418,In_363);
nand U451 (N_451,In_920,In_2899);
xor U452 (N_452,In_507,In_1715);
and U453 (N_453,In_1232,In_2307);
or U454 (N_454,In_2185,In_168);
nor U455 (N_455,In_1994,In_696);
xnor U456 (N_456,In_303,In_349);
xnor U457 (N_457,In_1488,In_600);
xor U458 (N_458,In_1213,In_33);
nor U459 (N_459,In_1734,In_792);
and U460 (N_460,In_2583,In_2865);
or U461 (N_461,In_2661,In_2835);
or U462 (N_462,In_2386,In_815);
and U463 (N_463,In_1371,In_144);
and U464 (N_464,In_1340,In_465);
xnor U465 (N_465,In_1448,In_18);
nor U466 (N_466,In_206,In_2084);
or U467 (N_467,In_1923,In_330);
nor U468 (N_468,In_1611,In_383);
nand U469 (N_469,In_2331,In_879);
and U470 (N_470,In_2617,In_1107);
or U471 (N_471,In_244,In_928);
xor U472 (N_472,In_1285,In_2519);
xnor U473 (N_473,In_2170,In_1240);
and U474 (N_474,In_835,In_2234);
and U475 (N_475,In_726,In_1434);
or U476 (N_476,In_203,In_1728);
nor U477 (N_477,In_799,In_1891);
nor U478 (N_478,In_2369,In_677);
or U479 (N_479,In_2410,In_2155);
or U480 (N_480,In_2827,In_1177);
and U481 (N_481,In_395,In_421);
and U482 (N_482,In_1729,In_1032);
nand U483 (N_483,In_1604,In_493);
or U484 (N_484,In_2418,In_272);
nor U485 (N_485,In_1308,In_1958);
nor U486 (N_486,In_1451,In_269);
or U487 (N_487,In_1583,In_2228);
nand U488 (N_488,In_1773,In_716);
and U489 (N_489,In_277,In_172);
nand U490 (N_490,In_906,In_1154);
nand U491 (N_491,In_1272,In_176);
or U492 (N_492,In_2085,In_1322);
and U493 (N_493,In_1569,In_1250);
or U494 (N_494,In_1642,In_2545);
nand U495 (N_495,In_1289,In_1335);
and U496 (N_496,In_1870,In_995);
and U497 (N_497,In_1674,In_1623);
nand U498 (N_498,In_207,In_1619);
or U499 (N_499,In_1027,In_183);
and U500 (N_500,In_1223,In_1918);
or U501 (N_501,In_1220,In_2407);
nor U502 (N_502,In_1833,In_2810);
or U503 (N_503,In_2311,In_2432);
nor U504 (N_504,In_359,In_1929);
nor U505 (N_505,In_505,In_220);
and U506 (N_506,In_782,In_936);
and U507 (N_507,In_1098,In_2495);
nor U508 (N_508,In_858,In_2094);
nor U509 (N_509,In_1824,In_593);
and U510 (N_510,In_2112,In_691);
and U511 (N_511,In_1124,In_458);
and U512 (N_512,In_399,In_247);
or U513 (N_513,In_241,In_1987);
nor U514 (N_514,In_2528,In_943);
xnor U515 (N_515,In_2552,In_504);
nand U516 (N_516,In_1280,In_101);
nor U517 (N_517,In_1321,In_2208);
and U518 (N_518,In_2419,In_1403);
and U519 (N_519,In_1843,In_137);
xor U520 (N_520,In_2163,In_2431);
nor U521 (N_521,In_510,In_484);
nor U522 (N_522,In_1410,In_1052);
xor U523 (N_523,In_781,In_1394);
xor U524 (N_524,In_591,In_2284);
and U525 (N_525,In_807,In_921);
or U526 (N_526,In_46,In_541);
and U527 (N_527,In_2723,In_1496);
or U528 (N_528,In_2250,In_449);
or U529 (N_529,In_767,In_931);
or U530 (N_530,In_72,In_1682);
nand U531 (N_531,In_225,In_2394);
or U532 (N_532,In_2799,In_2636);
and U533 (N_533,In_1039,In_485);
nand U534 (N_534,In_14,In_2472);
or U535 (N_535,In_2730,In_1992);
and U536 (N_536,In_2524,In_2291);
nor U537 (N_537,In_2780,In_96);
nor U538 (N_538,In_2157,In_753);
and U539 (N_539,In_2756,In_362);
nor U540 (N_540,In_1566,In_877);
and U541 (N_541,In_2244,In_1474);
nand U542 (N_542,In_2876,In_751);
and U543 (N_543,In_1507,In_2361);
or U544 (N_544,In_442,In_527);
nor U545 (N_545,In_972,In_2521);
and U546 (N_546,In_2323,In_132);
nor U547 (N_547,In_160,In_2622);
nand U548 (N_548,In_113,In_192);
nand U549 (N_549,In_2690,In_1043);
nor U550 (N_550,In_813,In_683);
nor U551 (N_551,In_230,In_2371);
and U552 (N_552,In_2236,In_1784);
nor U553 (N_553,In_838,In_2154);
nor U554 (N_554,In_2366,In_1236);
xnor U555 (N_555,In_790,In_295);
and U556 (N_556,In_2345,In_940);
xnor U557 (N_557,In_1261,In_1002);
or U558 (N_558,In_1151,In_1141);
xor U559 (N_559,In_2142,In_1858);
nand U560 (N_560,In_556,In_70);
xor U561 (N_561,In_1655,In_2767);
and U562 (N_562,In_876,In_85);
or U563 (N_563,In_111,In_1739);
or U564 (N_564,In_987,In_1054);
nor U565 (N_565,In_1828,In_36);
nand U566 (N_566,In_2842,In_1159);
nor U567 (N_567,In_2051,In_2464);
nor U568 (N_568,In_2988,In_1654);
nand U569 (N_569,In_951,In_2826);
xor U570 (N_570,In_396,In_341);
nand U571 (N_571,In_2364,In_2382);
nor U572 (N_572,In_2202,In_1658);
nor U573 (N_573,In_2011,In_2857);
or U574 (N_574,In_944,In_2561);
xnor U575 (N_575,In_2144,In_243);
or U576 (N_576,In_2809,In_1790);
nand U577 (N_577,In_2901,In_627);
nor U578 (N_578,In_2920,In_435);
nor U579 (N_579,In_1873,In_310);
or U580 (N_580,In_852,In_2313);
or U581 (N_581,In_1065,In_1819);
xnor U582 (N_582,In_1128,In_1011);
or U583 (N_583,In_335,In_804);
and U584 (N_584,In_13,In_2938);
nand U585 (N_585,In_1787,In_379);
nand U586 (N_586,In_1709,In_2269);
nand U587 (N_587,In_428,In_1209);
or U588 (N_588,In_2919,In_1917);
and U589 (N_589,In_1742,In_406);
and U590 (N_590,In_121,In_1345);
nand U591 (N_591,In_609,In_1412);
nor U592 (N_592,In_2643,In_2129);
or U593 (N_593,In_154,In_469);
or U594 (N_594,In_1173,In_1494);
nor U595 (N_595,In_2458,In_1948);
nand U596 (N_596,In_109,In_1489);
xor U597 (N_597,In_2789,In_318);
nor U598 (N_598,In_475,In_1640);
xnor U599 (N_599,In_2999,In_1462);
and U600 (N_600,In_2693,In_2665);
and U601 (N_601,In_197,In_1628);
and U602 (N_602,In_1665,In_862);
and U603 (N_603,In_2775,In_939);
or U604 (N_604,In_694,In_2375);
nand U605 (N_605,In_661,In_236);
and U606 (N_606,In_1750,In_1148);
xnor U607 (N_607,In_82,In_2430);
or U608 (N_608,In_777,In_2762);
xor U609 (N_609,In_1895,In_882);
nand U610 (N_610,In_1143,In_457);
and U611 (N_611,In_2181,In_117);
nand U612 (N_612,In_899,In_2438);
nand U613 (N_613,In_1930,In_1385);
xor U614 (N_614,In_436,In_970);
nor U615 (N_615,In_1470,In_2548);
nor U616 (N_616,In_613,In_1142);
and U617 (N_617,In_732,In_138);
xor U618 (N_618,In_1643,In_1373);
nor U619 (N_619,In_1890,In_843);
and U620 (N_620,In_147,In_2086);
and U621 (N_621,In_1471,In_746);
xnor U622 (N_622,In_55,In_1317);
xor U623 (N_623,In_248,In_907);
and U624 (N_624,In_1774,In_259);
or U625 (N_625,In_499,In_2021);
and U626 (N_626,In_2354,In_1360);
nand U627 (N_627,In_1456,In_2350);
nand U628 (N_628,In_528,In_2214);
nand U629 (N_629,In_2829,In_1003);
nor U630 (N_630,In_1309,In_136);
xor U631 (N_631,In_94,In_2019);
nor U632 (N_632,In_133,In_81);
or U633 (N_633,In_412,In_2921);
xor U634 (N_634,In_1717,In_750);
nor U635 (N_635,In_706,In_2978);
xnor U636 (N_636,In_2525,In_148);
and U637 (N_637,In_1892,In_385);
nor U638 (N_638,In_1467,In_2535);
and U639 (N_639,In_2761,In_2079);
xor U640 (N_640,In_1641,In_830);
xor U641 (N_641,In_2837,In_91);
xor U642 (N_642,In_42,In_1171);
or U643 (N_643,In_1731,In_885);
xor U644 (N_644,In_1775,In_1980);
or U645 (N_645,In_2624,In_2270);
nor U646 (N_646,In_2077,In_2755);
nand U647 (N_647,In_1889,In_1762);
nand U648 (N_648,In_616,In_2078);
or U649 (N_649,In_2764,In_1609);
nand U650 (N_650,In_1928,In_1536);
or U651 (N_651,In_93,In_2648);
or U652 (N_652,In_897,In_2264);
or U653 (N_653,In_2639,In_2520);
nor U654 (N_654,In_2463,In_938);
and U655 (N_655,In_780,In_1540);
or U656 (N_656,In_679,In_730);
or U657 (N_657,In_1931,In_2412);
and U658 (N_658,In_2542,In_676);
xor U659 (N_659,In_1333,In_1348);
xnor U660 (N_660,In_279,In_737);
and U661 (N_661,In_1307,In_2082);
or U662 (N_662,In_2769,In_2493);
and U663 (N_663,In_293,In_1316);
xnor U664 (N_664,In_12,In_2553);
xor U665 (N_665,In_2347,In_2852);
or U666 (N_666,In_473,In_2398);
or U667 (N_667,In_287,In_1392);
and U668 (N_668,In_2997,In_213);
and U669 (N_669,In_2315,In_2816);
nand U670 (N_670,In_522,In_1727);
and U671 (N_671,In_1384,In_1312);
or U672 (N_672,In_2601,In_2467);
nor U673 (N_673,In_916,In_1468);
xor U674 (N_674,In_1671,In_177);
nor U675 (N_675,In_2177,In_1);
or U676 (N_676,In_211,In_2137);
and U677 (N_677,In_1821,In_735);
nand U678 (N_678,In_459,In_866);
nor U679 (N_679,In_2888,In_642);
xor U680 (N_680,In_404,In_146);
nor U681 (N_681,In_2439,In_384);
nor U682 (N_682,In_370,In_2626);
nor U683 (N_683,In_560,In_2299);
nor U684 (N_684,In_980,In_724);
or U685 (N_685,In_1563,In_2186);
nand U686 (N_686,In_2904,In_1329);
xnor U687 (N_687,In_2001,In_1084);
nand U688 (N_688,In_1755,In_212);
xnor U689 (N_689,In_1884,In_888);
and U690 (N_690,In_1004,In_371);
xor U691 (N_691,In_2573,In_445);
xnor U692 (N_692,In_1305,In_2781);
nand U693 (N_693,In_1125,In_699);
nand U694 (N_694,In_649,In_1205);
nor U695 (N_695,In_35,In_1740);
and U696 (N_696,In_500,In_1443);
or U697 (N_697,In_1480,In_961);
and U698 (N_698,In_2946,In_143);
nor U699 (N_699,In_1817,In_483);
nor U700 (N_700,In_1252,In_2267);
nand U701 (N_701,In_2149,In_1666);
or U702 (N_702,In_1183,In_2954);
xnor U703 (N_703,In_881,In_2111);
or U704 (N_704,In_1692,In_2662);
or U705 (N_705,In_2621,In_2647);
nor U706 (N_706,In_83,In_1110);
and U707 (N_707,In_1161,In_2874);
nand U708 (N_708,In_729,In_1274);
xor U709 (N_709,In_297,In_1262);
or U710 (N_710,In_1269,In_1046);
nand U711 (N_711,In_1153,In_741);
nor U712 (N_712,In_2187,In_308);
nor U713 (N_713,In_883,In_89);
and U714 (N_714,In_919,In_1694);
nor U715 (N_715,In_968,In_97);
or U716 (N_716,In_1441,In_1681);
nand U717 (N_717,In_2266,In_1804);
nand U718 (N_718,In_357,In_2670);
or U719 (N_719,In_2746,In_2409);
and U720 (N_720,In_1146,In_2340);
or U721 (N_721,In_2069,In_736);
nand U722 (N_722,In_398,In_2168);
xor U723 (N_723,In_2020,In_1972);
or U724 (N_724,In_2634,In_317);
nor U725 (N_725,In_1538,In_2259);
xor U726 (N_726,In_2385,In_865);
nand U727 (N_727,In_670,In_1877);
and U728 (N_728,In_752,In_352);
nand U729 (N_729,In_890,In_559);
or U730 (N_730,In_1358,In_2054);
xnor U731 (N_731,In_517,In_2804);
nand U732 (N_732,In_1582,In_601);
or U733 (N_733,In_450,In_1561);
and U734 (N_734,In_1622,In_1273);
and U735 (N_735,In_2422,In_844);
nand U736 (N_736,In_189,In_908);
nand U737 (N_737,In_1794,In_912);
or U738 (N_738,In_2696,In_1749);
xor U739 (N_739,In_1185,In_2817);
nand U740 (N_740,In_2160,In_1916);
nor U741 (N_741,In_2415,In_2546);
nand U742 (N_742,In_867,In_239);
nor U743 (N_743,In_1947,In_2302);
nand U744 (N_744,In_831,In_163);
nand U745 (N_745,In_2968,In_2537);
and U746 (N_746,In_2365,In_285);
xnor U747 (N_747,In_1646,In_1070);
xor U748 (N_748,In_414,In_1555);
nor U749 (N_749,In_1368,In_2032);
or U750 (N_750,In_1964,In_2666);
or U751 (N_751,In_709,In_2221);
or U752 (N_752,In_325,In_621);
and U753 (N_753,In_665,In_2776);
and U754 (N_754,In_1668,In_10);
nand U755 (N_755,In_2436,In_759);
xnor U756 (N_756,In_155,In_924);
nor U757 (N_757,In_1445,In_1175);
nand U758 (N_758,In_2523,In_2765);
nor U759 (N_759,In_376,In_1751);
nand U760 (N_760,In_2689,In_1211);
nor U761 (N_761,In_1772,In_2304);
nand U762 (N_762,In_2093,In_2293);
and U763 (N_763,In_201,In_2785);
nand U764 (N_764,In_2726,In_2446);
nand U765 (N_765,In_547,In_647);
or U766 (N_766,In_1568,In_562);
nand U767 (N_767,In_1594,In_1062);
nand U768 (N_768,In_2289,In_345);
xor U769 (N_769,In_1139,In_1400);
or U770 (N_770,In_1095,In_1045);
and U771 (N_771,In_2915,In_1940);
xnor U772 (N_772,In_2738,In_237);
nand U773 (N_773,In_715,In_2733);
xnor U774 (N_774,In_1885,In_911);
nor U775 (N_775,In_818,In_234);
or U776 (N_776,In_1976,In_106);
xor U777 (N_777,In_328,In_1607);
and U778 (N_778,In_2171,In_1776);
xor U779 (N_779,In_1564,In_1157);
xor U780 (N_780,In_632,In_2480);
xnor U781 (N_781,In_974,In_903);
xnor U782 (N_782,In_1901,In_2507);
nor U783 (N_783,In_2184,In_1842);
nor U784 (N_784,In_1111,In_969);
nor U785 (N_785,In_1416,In_2853);
nor U786 (N_786,In_667,In_51);
nor U787 (N_787,In_2875,In_2699);
nor U788 (N_788,In_2478,In_116);
nand U789 (N_789,In_2740,In_1088);
and U790 (N_790,In_2638,In_2860);
xnor U791 (N_791,In_1521,In_1121);
nand U792 (N_792,In_1998,In_1985);
nand U793 (N_793,In_1349,In_1200);
xor U794 (N_794,In_1022,In_1659);
xor U795 (N_795,In_2000,In_2748);
xnor U796 (N_796,In_119,In_235);
or U797 (N_797,In_2175,In_6);
xor U798 (N_798,In_1519,In_692);
and U799 (N_799,In_5,In_950);
nand U800 (N_800,In_2625,In_266);
nand U801 (N_801,In_198,In_2563);
xnor U802 (N_802,In_2914,In_2475);
xnor U803 (N_803,In_563,In_495);
xnor U804 (N_804,In_56,In_2667);
nor U805 (N_805,In_2276,In_1543);
nand U806 (N_806,In_1131,In_452);
xor U807 (N_807,In_2510,In_1076);
xor U808 (N_808,In_1079,In_1689);
xor U809 (N_809,In_2702,In_2454);
and U810 (N_810,In_2353,In_401);
xnor U811 (N_811,In_1390,In_2608);
nor U812 (N_812,In_102,In_2477);
nor U813 (N_813,In_1575,In_423);
xor U814 (N_814,In_21,In_2035);
xnor U815 (N_815,In_1350,In_1048);
xor U816 (N_816,In_1080,In_2326);
nor U817 (N_817,In_2557,In_2107);
xnor U818 (N_818,In_480,In_1134);
nand U819 (N_819,In_1353,In_1440);
nor U820 (N_820,In_1459,In_1168);
xor U821 (N_821,In_947,In_2889);
and U822 (N_822,In_2497,In_1376);
xnor U823 (N_823,In_789,In_39);
nor U824 (N_824,In_309,In_666);
nand U825 (N_825,In_948,In_246);
and U826 (N_826,In_2555,In_868);
nand U827 (N_827,In_635,In_2961);
and U828 (N_828,In_1466,In_1518);
and U829 (N_829,In_626,In_565);
and U830 (N_830,In_927,In_2457);
or U831 (N_831,In_2703,In_1019);
nand U832 (N_832,In_960,In_2081);
and U833 (N_833,In_394,In_2012);
and U834 (N_834,In_1820,In_848);
and U835 (N_835,In_2016,In_2751);
and U836 (N_836,In_1968,In_631);
or U837 (N_837,In_282,In_1597);
nand U838 (N_838,In_1279,In_2309);
nor U839 (N_839,In_850,In_2924);
nand U840 (N_840,In_2308,In_2153);
or U841 (N_841,In_1160,In_184);
nand U842 (N_842,In_1035,In_2672);
xnor U843 (N_843,In_2044,In_538);
or U844 (N_844,In_1813,In_1228);
and U845 (N_845,In_2577,In_2743);
nor U846 (N_846,In_1886,In_587);
xnor U847 (N_847,In_703,In_993);
and U848 (N_848,In_2588,In_2759);
xor U849 (N_849,In_985,In_957);
xnor U850 (N_850,In_327,In_125);
nand U851 (N_851,In_958,In_892);
xor U852 (N_852,In_2335,In_2285);
and U853 (N_853,In_1001,In_1504);
or U854 (N_854,In_1090,In_2824);
or U855 (N_855,In_103,In_2540);
nor U856 (N_856,In_227,In_305);
nand U857 (N_857,In_1108,In_2959);
and U858 (N_858,In_1055,In_821);
nor U859 (N_859,In_1943,In_2694);
nor U860 (N_860,In_263,In_11);
xnor U861 (N_861,In_2580,In_2505);
and U862 (N_862,In_1530,In_764);
nor U863 (N_863,In_582,In_1531);
nand U864 (N_864,In_2911,In_1587);
xnor U865 (N_865,In_489,In_1713);
nand U866 (N_866,In_607,In_1639);
nand U867 (N_867,In_1315,In_675);
or U868 (N_868,In_795,In_219);
nor U869 (N_869,In_891,In_2512);
or U870 (N_870,In_832,In_524);
nand U871 (N_871,In_1818,In_1005);
and U872 (N_872,In_2403,In_2113);
nor U873 (N_873,In_827,In_2936);
xor U874 (N_874,In_2140,In_2130);
xor U875 (N_875,In_2260,In_118);
and U876 (N_876,In_1848,In_2922);
xnor U877 (N_877,In_1983,In_2770);
and U878 (N_878,In_1476,In_1401);
nand U879 (N_879,In_712,In_2823);
nor U880 (N_880,In_997,In_86);
or U881 (N_881,In_2138,In_461);
nor U882 (N_882,In_430,In_2332);
xnor U883 (N_883,In_2484,In_1874);
or U884 (N_884,In_1615,In_771);
and U885 (N_885,In_646,In_1841);
and U886 (N_886,In_1072,In_1922);
and U887 (N_887,In_2381,In_2087);
or U888 (N_888,In_112,In_1014);
and U889 (N_889,In_1361,In_1722);
nand U890 (N_890,In_181,In_1522);
nand U891 (N_891,In_895,In_2909);
nand U892 (N_892,In_1618,In_115);
and U893 (N_893,In_289,In_503);
nand U894 (N_894,In_990,In_1570);
or U895 (N_895,In_605,In_2197);
or U896 (N_896,In_2698,In_1730);
or U897 (N_897,In_2215,In_1938);
or U898 (N_898,In_1955,In_65);
xnor U899 (N_899,In_2970,In_400);
and U900 (N_900,In_1505,In_194);
nand U901 (N_901,In_2055,In_2169);
nor U902 (N_902,In_22,In_994);
nand U903 (N_903,In_2612,In_2676);
or U904 (N_904,In_438,In_791);
xnor U905 (N_905,In_1593,In_1267);
and U906 (N_906,In_1040,In_61);
and U907 (N_907,In_2526,In_1667);
or U908 (N_908,In_1379,In_516);
xnor U909 (N_909,In_1977,In_1866);
nor U910 (N_910,In_2402,In_1825);
nor U911 (N_911,In_249,In_1414);
or U912 (N_912,In_1347,In_2940);
nand U913 (N_913,In_1832,In_2674);
or U914 (N_914,In_2596,In_1181);
nand U915 (N_915,In_1508,In_954);
xor U916 (N_916,In_1007,In_1163);
nand U917 (N_917,In_946,In_845);
nor U918 (N_918,In_476,In_829);
nor U919 (N_919,In_2935,In_2753);
or U920 (N_920,In_910,In_651);
and U921 (N_921,In_41,In_1030);
nor U922 (N_922,In_617,In_1226);
nor U923 (N_923,In_276,In_2715);
nand U924 (N_924,In_1291,In_1325);
nand U925 (N_925,In_2547,In_2846);
or U926 (N_926,In_1737,In_1263);
or U927 (N_927,In_478,In_2902);
nor U928 (N_928,In_673,In_603);
nand U929 (N_929,In_1517,In_851);
nand U930 (N_930,In_2980,In_963);
or U931 (N_931,In_2134,In_2814);
xor U932 (N_932,In_2931,In_27);
nand U933 (N_933,In_2443,In_2768);
and U934 (N_934,In_2737,In_2834);
xnor U935 (N_935,In_389,In_1409);
xnor U936 (N_936,In_223,In_511);
or U937 (N_937,In_717,In_2073);
or U938 (N_938,In_1227,In_922);
and U939 (N_939,In_2468,In_1907);
and U940 (N_940,In_754,In_1396);
and U941 (N_941,In_2877,In_1588);
or U942 (N_942,In_2104,In_1799);
nor U943 (N_943,In_2042,In_2489);
or U944 (N_944,In_2408,In_558);
xnor U945 (N_945,In_798,In_684);
and U946 (N_946,In_610,In_1550);
nor U947 (N_947,In_2592,In_2173);
nand U948 (N_948,In_834,In_444);
xnor U949 (N_949,In_1803,In_2098);
xnor U950 (N_950,In_1796,In_825);
nor U951 (N_951,In_809,In_1217);
nor U952 (N_952,In_2368,In_2994);
nand U953 (N_953,In_1634,In_873);
or U954 (N_954,In_2602,In_966);
and U955 (N_955,In_2974,In_2879);
or U956 (N_956,In_1632,In_1802);
nand U957 (N_957,In_681,In_2373);
nor U958 (N_958,In_373,In_2248);
nor U959 (N_959,In_2722,In_1953);
nand U960 (N_960,In_1114,In_718);
or U961 (N_961,In_2847,In_467);
xnor U962 (N_962,In_2871,In_2897);
xor U963 (N_963,In_1123,In_1461);
xnor U964 (N_964,In_2491,In_1696);
xor U965 (N_965,In_2604,In_2855);
nand U966 (N_966,In_1975,In_366);
xnor U967 (N_967,In_2973,In_2567);
nor U968 (N_968,In_304,In_592);
or U969 (N_969,In_88,In_1241);
nor U970 (N_970,In_2774,In_925);
and U971 (N_971,In_1856,In_1018);
or U972 (N_972,In_1020,In_411);
and U973 (N_973,In_2752,In_2376);
nand U974 (N_974,In_296,In_1899);
or U975 (N_975,In_2148,In_1656);
nor U976 (N_976,In_680,In_1483);
nor U977 (N_977,In_1677,In_1982);
or U978 (N_978,In_1387,In_814);
or U979 (N_979,In_1069,In_1506);
or U980 (N_980,In_977,In_205);
and U981 (N_981,In_321,In_175);
nor U982 (N_982,In_561,In_191);
nor U983 (N_983,In_967,In_548);
xnor U984 (N_984,In_1919,In_2282);
nor U985 (N_985,In_2397,In_1961);
or U986 (N_986,In_532,In_2967);
or U987 (N_987,In_1056,In_1338);
nor U988 (N_988,In_2908,In_763);
nor U989 (N_989,In_2178,In_2786);
or U990 (N_990,In_854,In_886);
nor U991 (N_991,In_1523,In_1195);
xnor U992 (N_992,In_1194,In_2200);
nor U993 (N_993,In_1600,In_166);
nand U994 (N_994,In_1879,In_2605);
and U995 (N_995,In_2522,In_2355);
nor U996 (N_996,In_1524,In_2982);
or U997 (N_997,In_2092,In_2427);
nand U998 (N_998,In_60,In_2351);
or U999 (N_999,In_1479,In_369);
xor U1000 (N_1000,In_870,In_1473);
xnor U1001 (N_1001,In_1342,In_1439);
nand U1002 (N_1002,In_1327,In_1431);
and U1003 (N_1003,In_1720,In_1549);
and U1004 (N_1004,In_2167,In_1397);
nand U1005 (N_1005,In_2456,In_1605);
nor U1006 (N_1006,In_408,In_2841);
and U1007 (N_1007,In_1104,In_955);
and U1008 (N_1008,In_377,In_2179);
or U1009 (N_1009,In_900,In_2965);
and U1010 (N_1010,In_1215,In_1652);
or U1011 (N_1011,In_1993,In_648);
nand U1012 (N_1012,In_551,In_180);
xor U1013 (N_1013,In_1135,In_1673);
nor U1014 (N_1014,In_1025,In_1186);
and U1015 (N_1015,In_2984,In_2091);
nor U1016 (N_1016,In_2437,In_1743);
and U1017 (N_1017,In_1031,In_2152);
nor U1018 (N_1018,In_368,In_2461);
or U1019 (N_1019,In_1097,In_566);
and U1020 (N_1020,In_336,In_727);
or U1021 (N_1021,In_1074,In_2024);
nor U1022 (N_1022,In_466,In_1036);
nor U1023 (N_1023,In_2534,In_2773);
xnor U1024 (N_1024,In_390,In_2047);
and U1025 (N_1025,In_1399,In_1670);
nor U1026 (N_1026,In_2254,In_1785);
or U1027 (N_1027,In_1010,In_313);
xnor U1028 (N_1028,In_1855,In_2611);
or U1029 (N_1029,In_747,In_1354);
nand U1030 (N_1030,In_1253,In_602);
or U1031 (N_1031,In_464,In_1789);
or U1032 (N_1032,In_1086,In_1006);
and U1033 (N_1033,In_2310,In_2957);
or U1034 (N_1034,In_812,In_711);
or U1035 (N_1035,In_1071,In_1306);
nand U1036 (N_1036,In_775,In_1363);
and U1037 (N_1037,In_1944,In_270);
xor U1038 (N_1038,In_596,In_658);
or U1039 (N_1039,In_409,In_1331);
xnor U1040 (N_1040,In_2579,In_378);
or U1041 (N_1041,In_1047,In_2275);
xor U1042 (N_1042,In_2784,In_655);
xnor U1043 (N_1043,In_1286,In_1257);
nand U1044 (N_1044,In_1017,In_233);
and U1045 (N_1045,In_322,In_193);
nor U1046 (N_1046,In_437,In_2277);
or U1047 (N_1047,In_1405,In_1015);
nor U1048 (N_1048,In_1621,In_630);
xnor U1049 (N_1049,In_2813,In_1436);
and U1050 (N_1050,In_382,In_1365);
and U1051 (N_1051,In_569,In_871);
xnor U1052 (N_1052,In_1991,In_1544);
nor U1053 (N_1053,In_77,In_2490);
and U1054 (N_1054,In_1771,In_2849);
xnor U1055 (N_1055,In_1744,In_1472);
xnor U1056 (N_1056,In_2416,In_1732);
xor U1057 (N_1057,In_989,In_2039);
xnor U1058 (N_1058,In_1827,In_2713);
nor U1059 (N_1059,In_1234,In_2159);
nand U1060 (N_1060,In_17,In_1812);
xnor U1061 (N_1061,In_904,In_332);
or U1062 (N_1062,In_964,In_2442);
or U1063 (N_1063,In_1557,In_633);
nor U1064 (N_1064,In_999,In_1791);
and U1065 (N_1065,In_1914,In_2778);
xnor U1066 (N_1066,In_2048,In_2022);
and U1067 (N_1067,In_2015,In_2503);
or U1068 (N_1068,In_48,In_2448);
xnor U1069 (N_1069,In_778,In_71);
nand U1070 (N_1070,In_364,In_1596);
or U1071 (N_1071,In_2195,In_284);
nand U1072 (N_1072,In_2680,In_1545);
xnor U1073 (N_1073,In_2883,In_324);
nor U1074 (N_1074,In_187,In_2062);
xnor U1075 (N_1075,In_757,In_1116);
xor U1076 (N_1076,In_2509,In_1834);
xnor U1077 (N_1077,In_2352,In_329);
and U1078 (N_1078,In_2396,In_1122);
nand U1079 (N_1079,In_1700,In_9);
nand U1080 (N_1080,In_1935,In_1614);
nand U1081 (N_1081,In_1463,In_2007);
or U1082 (N_1082,In_1162,In_290);
nor U1083 (N_1083,In_695,In_1989);
xor U1084 (N_1084,In_2235,In_2161);
or U1085 (N_1085,In_1904,In_1537);
nand U1086 (N_1086,In_1912,In_481);
or U1087 (N_1087,In_1324,In_2286);
or U1088 (N_1088,In_2787,In_2471);
xor U1089 (N_1089,In_319,In_577);
nor U1090 (N_1090,In_342,In_574);
nand U1091 (N_1091,In_784,In_2298);
and U1092 (N_1092,In_678,In_2462);
or U1093 (N_1093,In_570,In_1539);
xor U1094 (N_1094,In_1839,In_986);
nand U1095 (N_1095,In_2492,In_1293);
and U1096 (N_1096,In_1814,In_1932);
and U1097 (N_1097,In_2686,In_1427);
nand U1098 (N_1098,In_2716,In_1182);
nor U1099 (N_1099,In_2218,In_140);
and U1100 (N_1100,In_2306,In_822);
and U1101 (N_1101,In_1395,In_2390);
and U1102 (N_1102,In_998,In_222);
nand U1103 (N_1103,In_314,In_2363);
and U1104 (N_1104,In_2433,In_2165);
nand U1105 (N_1105,In_2424,In_1164);
xnor U1106 (N_1106,In_2620,In_1738);
xnor U1107 (N_1107,In_2300,In_2003);
nand U1108 (N_1108,In_1883,In_69);
nor U1109 (N_1109,In_1965,In_2964);
or U1110 (N_1110,In_1826,In_612);
xnor U1111 (N_1111,In_1761,In_2317);
and U1112 (N_1112,In_199,In_2934);
nand U1113 (N_1113,In_615,In_2987);
or U1114 (N_1114,In_1346,In_1270);
nand U1115 (N_1115,In_1529,In_153);
nand U1116 (N_1116,In_749,In_1714);
xnor U1117 (N_1117,In_671,In_2296);
or U1118 (N_1118,In_2885,In_2944);
nand U1119 (N_1119,In_2905,In_2075);
xor U1120 (N_1120,In_2429,In_1631);
nor U1121 (N_1121,In_932,In_2711);
and U1122 (N_1122,In_887,In_2370);
and U1123 (N_1123,In_1534,In_232);
nor U1124 (N_1124,In_1844,In_1136);
xor U1125 (N_1125,In_271,In_535);
nand U1126 (N_1126,In_2614,In_252);
nand U1127 (N_1127,In_2515,In_2190);
or U1128 (N_1128,In_1707,In_1302);
nor U1129 (N_1129,In_1190,In_1815);
xor U1130 (N_1130,In_2388,In_2037);
or U1131 (N_1131,In_1735,In_1786);
xor U1132 (N_1132,In_164,In_536);
and U1133 (N_1133,In_90,In_1100);
xor U1134 (N_1134,In_1063,In_2771);
xor U1135 (N_1135,In_1326,In_1367);
nand U1136 (N_1136,In_1721,In_2133);
and U1137 (N_1137,In_2609,In_2229);
xor U1138 (N_1138,In_419,In_723);
and U1139 (N_1139,In_2603,In_1860);
nor U1140 (N_1140,In_2966,In_2867);
or U1141 (N_1141,In_251,In_380);
and U1142 (N_1142,In_1712,In_221);
nand U1143 (N_1143,In_501,In_281);
or U1144 (N_1144,In_1981,In_2337);
xnor U1145 (N_1145,In_1296,In_1313);
xnor U1146 (N_1146,In_2328,In_151);
and U1147 (N_1147,In_710,In_863);
or U1148 (N_1148,In_2013,In_2812);
nor U1149 (N_1149,In_1497,In_190);
or U1150 (N_1150,In_530,In_1233);
and U1151 (N_1151,In_1513,In_2139);
and U1152 (N_1152,In_1337,In_209);
nand U1153 (N_1153,In_178,In_1336);
or U1154 (N_1154,In_1311,In_1117);
and U1155 (N_1155,In_688,In_2597);
xor U1156 (N_1156,In_1584,In_1777);
and U1157 (N_1157,In_1903,In_1565);
or U1158 (N_1158,In_713,In_1119);
nand U1159 (N_1159,In_553,In_686);
or U1160 (N_1160,In_2488,In_139);
nand U1161 (N_1161,In_2880,In_407);
and U1162 (N_1162,In_1145,In_344);
xnor U1163 (N_1163,In_470,In_1996);
nor U1164 (N_1164,In_1029,In_902);
and U1165 (N_1165,In_2482,In_1426);
or U1166 (N_1166,In_2559,In_105);
xnor U1167 (N_1167,In_182,In_1318);
and U1168 (N_1168,In_59,In_1925);
xor U1169 (N_1169,In_1191,In_53);
nor U1170 (N_1170,In_1198,In_2);
nand U1171 (N_1171,In_595,In_2903);
xnor U1172 (N_1172,In_534,In_2256);
nor U1173 (N_1173,In_1096,In_8);
or U1174 (N_1174,In_820,In_1444);
or U1175 (N_1175,In_2582,In_2663);
nand U1176 (N_1176,In_2399,In_721);
and U1177 (N_1177,In_1268,In_161);
and U1178 (N_1178,In_1402,In_150);
nand U1179 (N_1179,In_2565,In_2319);
or U1180 (N_1180,In_2763,In_2224);
and U1181 (N_1181,In_1320,In_1485);
nand U1182 (N_1182,In_1158,In_439);
and U1183 (N_1183,In_156,In_2114);
and U1184 (N_1184,In_2806,In_1645);
or U1185 (N_1185,In_1375,In_1882);
or U1186 (N_1186,In_2708,In_945);
and U1187 (N_1187,In_24,In_1747);
and U1188 (N_1188,In_294,In_1945);
nand U1189 (N_1189,In_1793,In_257);
nor U1190 (N_1190,In_2747,In_2205);
or U1191 (N_1191,In_929,In_1579);
xor U1192 (N_1192,In_1875,In_1541);
nor U1193 (N_1193,In_2251,In_268);
and U1194 (N_1194,In_120,In_625);
nor U1195 (N_1195,In_76,In_2760);
nor U1196 (N_1196,In_1836,In_704);
nor U1197 (N_1197,In_422,In_2530);
xnor U1198 (N_1198,In_2913,In_2782);
and U1199 (N_1199,In_2120,In_1602);
xor U1200 (N_1200,In_755,In_2434);
nand U1201 (N_1201,In_1822,In_1763);
nor U1202 (N_1202,In_1000,In_361);
and U1203 (N_1203,In_2393,In_1137);
or U1204 (N_1204,In_728,In_1169);
or U1205 (N_1205,In_1242,In_2854);
and U1206 (N_1206,In_2906,In_1077);
nand U1207 (N_1207,In_533,In_158);
nor U1208 (N_1208,In_1736,In_75);
and U1209 (N_1209,In_2868,In_1214);
or U1210 (N_1210,In_984,In_2701);
nor U1211 (N_1211,In_1166,In_479);
nor U1212 (N_1212,In_1464,In_2652);
or U1213 (N_1213,In_598,In_1429);
xnor U1214 (N_1214,In_2358,In_1629);
xor U1215 (N_1215,In_2995,In_63);
nand U1216 (N_1216,In_2709,In_1783);
or U1217 (N_1217,In_765,In_2851);
nor U1218 (N_1218,In_157,In_2348);
nor U1219 (N_1219,In_1986,In_1888);
and U1220 (N_1220,In_1359,In_1260);
or U1221 (N_1221,In_1724,In_513);
xor U1222 (N_1222,In_909,In_1180);
xnor U1223 (N_1223,In_2710,In_1449);
nand U1224 (N_1224,In_1558,In_2058);
xnor U1225 (N_1225,In_2918,In_1415);
nor U1226 (N_1226,In_2295,In_2933);
or U1227 (N_1227,In_1660,In_2128);
nor U1228 (N_1228,In_2219,In_2593);
and U1229 (N_1229,In_1950,In_392);
nand U1230 (N_1230,In_2210,In_1962);
or U1231 (N_1231,In_2292,In_375);
xnor U1232 (N_1232,In_1756,In_1026);
or U1233 (N_1233,In_2387,In_1059);
xnor U1234 (N_1234,In_2008,In_2796);
xnor U1235 (N_1235,In_923,In_2822);
and U1236 (N_1236,In_2627,In_1997);
nor U1237 (N_1237,In_1406,In_739);
xor U1238 (N_1238,In_1578,In_1562);
and U1239 (N_1239,In_2986,In_1608);
or U1240 (N_1240,In_1648,In_1927);
xnor U1241 (N_1241,In_652,In_47);
or U1242 (N_1242,In_1999,In_1525);
nand U1243 (N_1243,In_2268,In_811);
nand U1244 (N_1244,In_334,In_2257);
and U1245 (N_1245,In_1258,In_2014);
and U1246 (N_1246,In_2241,In_1382);
or U1247 (N_1247,In_1679,In_663);
nand U1248 (N_1248,In_2623,In_1140);
and U1249 (N_1249,In_1068,In_1178);
nor U1250 (N_1250,In_262,In_1905);
or U1251 (N_1251,In_2237,In_1849);
xor U1252 (N_1252,In_441,In_2685);
xor U1253 (N_1253,In_981,In_2344);
or U1254 (N_1254,In_2862,In_2283);
nor U1255 (N_1255,In_1442,In_2391);
xnor U1256 (N_1256,In_707,In_1352);
nor U1257 (N_1257,In_656,In_1746);
nor U1258 (N_1258,In_74,In_26);
nor U1259 (N_1259,In_1013,In_1878);
nor U1260 (N_1260,In_1971,In_1946);
or U1261 (N_1261,In_2878,In_1798);
or U1262 (N_1262,In_413,In_2790);
or U1263 (N_1263,In_391,In_2356);
nand U1264 (N_1264,In_2729,In_487);
xor U1265 (N_1265,In_1748,In_531);
nor U1266 (N_1266,In_2996,In_2097);
and U1267 (N_1267,In_2127,In_515);
xnor U1268 (N_1268,In_2886,In_588);
nand U1269 (N_1269,In_731,In_2222);
or U1270 (N_1270,In_2049,In_1808);
or U1271 (N_1271,In_1676,In_840);
or U1272 (N_1272,In_1106,In_901);
and U1273 (N_1273,In_79,In_134);
or U1274 (N_1274,In_611,In_689);
and U1275 (N_1275,In_2993,In_1129);
and U1276 (N_1276,In_1093,In_149);
xnor U1277 (N_1277,In_1509,In_874);
xnor U1278 (N_1278,In_2041,In_1906);
nand U1279 (N_1279,In_1492,In_2516);
nor U1280 (N_1280,In_2514,In_918);
and U1281 (N_1281,In_2338,In_2788);
xnor U1282 (N_1282,In_415,In_337);
or U1283 (N_1283,In_2615,In_933);
nand U1284 (N_1284,In_474,In_2444);
nand U1285 (N_1285,In_1259,In_226);
nand U1286 (N_1286,In_2589,In_1937);
xor U1287 (N_1287,In_2989,In_1672);
nor U1288 (N_1288,In_2794,In_624);
xor U1289 (N_1289,In_1719,In_2360);
or U1290 (N_1290,In_2476,In_1487);
or U1291 (N_1291,In_95,In_124);
and U1292 (N_1292,In_1547,In_393);
and U1293 (N_1293,In_57,In_766);
or U1294 (N_1294,In_2119,In_2976);
nor U1295 (N_1295,In_2820,In_1601);
or U1296 (N_1296,In_1546,In_1067);
nand U1297 (N_1297,In_2952,In_416);
and U1298 (N_1298,In_638,In_2176);
and U1299 (N_1299,In_356,In_283);
nor U1300 (N_1300,In_762,In_240);
and U1301 (N_1301,In_779,In_1174);
nor U1302 (N_1302,In_1590,In_1033);
nor U1303 (N_1303,In_267,In_64);
nor U1304 (N_1304,In_2808,In_1697);
or U1305 (N_1305,In_229,In_1936);
and U1306 (N_1306,In_347,In_2109);
xor U1307 (N_1307,In_426,In_1809);
xor U1308 (N_1308,In_552,In_1425);
nor U1309 (N_1309,In_2303,In_2704);
nor U1310 (N_1310,In_2428,In_1624);
xnor U1311 (N_1311,In_1231,In_1612);
xnor U1312 (N_1312,In_1218,In_2329);
nor U1313 (N_1313,In_1533,In_1829);
xnor U1314 (N_1314,In_1127,In_1846);
nand U1315 (N_1315,In_1362,In_806);
and U1316 (N_1316,In_669,In_169);
nor U1317 (N_1317,In_2100,In_214);
nand U1318 (N_1318,In_1581,In_894);
or U1319 (N_1319,In_1332,In_1281);
or U1320 (N_1320,In_1915,In_142);
xnor U1321 (N_1321,In_1831,In_2754);
and U1322 (N_1322,In_2389,In_2675);
or U1323 (N_1323,In_1500,In_218);
or U1324 (N_1324,In_1688,In_2684);
xor U1325 (N_1325,In_2595,In_2539);
xnor U1326 (N_1326,In_1478,In_2945);
nand U1327 (N_1327,In_2483,In_1765);
xnor U1328 (N_1328,In_2066,In_1711);
and U1329 (N_1329,In_2341,In_98);
and U1330 (N_1330,In_2421,In_2322);
nand U1331 (N_1331,In_2550,In_1838);
or U1332 (N_1332,In_2599,In_590);
and U1333 (N_1333,In_720,In_2124);
and U1334 (N_1334,In_2379,In_823);
nand U1335 (N_1335,In_29,In_2449);
or U1336 (N_1336,In_1910,In_1417);
xnor U1337 (N_1337,In_1716,In_1081);
or U1338 (N_1338,In_1364,In_2096);
nand U1339 (N_1339,In_2893,In_2246);
xor U1340 (N_1340,In_1446,In_2324);
and U1341 (N_1341,In_1617,In_1599);
or U1342 (N_1342,In_2481,In_1845);
and U1343 (N_1343,In_2072,In_1908);
or U1344 (N_1344,In_701,In_971);
xor U1345 (N_1345,In_1165,In_599);
nor U1346 (N_1346,In_2357,In_425);
xor U1347 (N_1347,In_2655,In_2700);
and U1348 (N_1348,In_1264,In_1805);
nor U1349 (N_1349,In_1887,In_2036);
xnor U1350 (N_1350,In_2932,In_1933);
nand U1351 (N_1351,In_171,In_1704);
nor U1352 (N_1352,In_760,In_573);
xor U1353 (N_1353,In_2076,In_1852);
nor U1354 (N_1354,In_2209,In_1341);
xnor U1355 (N_1355,In_1278,In_2216);
xnor U1356 (N_1356,In_1038,In_496);
nand U1357 (N_1357,In_1099,In_2059);
nand U1358 (N_1358,In_2095,In_1024);
nor U1359 (N_1359,In_2470,In_2080);
and U1360 (N_1360,In_2943,In_365);
and U1361 (N_1361,In_2554,In_1952);
nor U1362 (N_1362,In_1113,In_2028);
nor U1363 (N_1363,In_2496,In_745);
nor U1364 (N_1364,In_1920,In_1457);
nand U1365 (N_1365,In_1553,In_1212);
and U1366 (N_1366,In_2807,In_1864);
or U1367 (N_1367,In_54,In_2687);
nor U1368 (N_1368,In_2131,In_1377);
xnor U1369 (N_1369,In_1247,In_1248);
nor U1370 (N_1370,In_1637,In_1391);
xnor U1371 (N_1371,In_486,In_2225);
nor U1372 (N_1372,In_1693,In_685);
xnor U1373 (N_1373,In_1591,In_1199);
or U1374 (N_1374,In_210,In_2272);
nor U1375 (N_1375,In_1381,In_1725);
or U1376 (N_1376,In_855,In_847);
nand U1377 (N_1377,In_1156,In_2105);
nand U1378 (N_1378,In_1577,In_2890);
and U1379 (N_1379,In_2211,In_2339);
nor U1380 (N_1380,In_2720,In_1101);
or U1381 (N_1381,In_4,In_2115);
or U1382 (N_1382,In_498,In_2025);
nor U1383 (N_1383,In_1678,In_1585);
or U1384 (N_1384,In_2166,In_1939);
and U1385 (N_1385,In_2527,In_1949);
or U1386 (N_1386,In_783,In_2132);
or U1387 (N_1387,In_1271,In_620);
or U1388 (N_1388,In_1057,In_1193);
or U1389 (N_1389,In_1840,In_1924);
xor U1390 (N_1390,In_2452,In_2240);
nand U1391 (N_1391,In_2815,In_502);
and U1392 (N_1392,In_2413,In_1393);
and U1393 (N_1393,In_0,In_2465);
xor U1394 (N_1394,In_889,In_740);
nand U1395 (N_1395,In_2691,In_2156);
and U1396 (N_1396,In_1548,In_1130);
or U1397 (N_1397,In_2640,In_1298);
xor U1398 (N_1398,In_1388,In_1249);
nor U1399 (N_1399,In_1435,In_2644);
or U1400 (N_1400,In_417,In_2196);
xor U1401 (N_1401,In_2164,In_708);
nor U1402 (N_1402,In_1450,In_1515);
nand U1403 (N_1403,In_1663,In_1120);
xor U1404 (N_1404,In_472,In_2958);
or U1405 (N_1405,In_2831,In_2217);
xor U1406 (N_1406,In_25,In_1970);
xor U1407 (N_1407,In_31,In_255);
or U1408 (N_1408,In_1703,In_2194);
nor U1409 (N_1409,In_702,In_1675);
nor U1410 (N_1410,In_915,In_2349);
nor U1411 (N_1411,In_2252,In_2739);
xor U1412 (N_1412,In_722,In_2801);
or U1413 (N_1413,In_402,In_2618);
nand U1414 (N_1414,In_2359,In_7);
nor U1415 (N_1415,In_659,In_1754);
and U1416 (N_1416,In_1222,In_2445);
nor U1417 (N_1417,In_571,In_2673);
and U1418 (N_1418,In_1189,In_273);
and U1419 (N_1419,In_2731,In_1491);
or U1420 (N_1420,In_1453,In_1028);
and U1421 (N_1421,In_2253,In_1037);
and U1422 (N_1422,In_1486,In_2220);
and U1423 (N_1423,In_1452,In_594);
xnor U1424 (N_1424,In_2271,In_1398);
xnor U1425 (N_1425,In_1087,In_2150);
and U1426 (N_1426,In_431,In_354);
nand U1427 (N_1427,In_2975,In_216);
xor U1428 (N_1428,In_2242,In_110);
xnor U1429 (N_1429,In_2010,In_1684);
xnor U1430 (N_1430,In_1454,In_2948);
xnor U1431 (N_1431,In_2844,In_2679);
and U1432 (N_1432,In_937,In_2330);
or U1433 (N_1433,In_162,In_991);
and U1434 (N_1434,In_2688,In_2591);
or U1435 (N_1435,In_2637,In_1265);
and U1436 (N_1436,In_2985,In_1411);
nand U1437 (N_1437,In_339,In_1133);
and U1438 (N_1438,In_2741,In_2631);
or U1439 (N_1439,In_37,In_1422);
or U1440 (N_1440,In_1680,In_261);
or U1441 (N_1441,In_2146,In_1009);
nor U1442 (N_1442,In_2736,In_1567);
xor U1443 (N_1443,In_636,In_606);
nand U1444 (N_1444,In_159,In_1455);
nor U1445 (N_1445,In_424,In_2053);
xor U1446 (N_1446,In_2501,In_367);
nor U1447 (N_1447,In_2401,In_2377);
nand U1448 (N_1448,In_2201,In_372);
or U1449 (N_1449,In_1706,In_291);
nor U1450 (N_1450,In_2450,In_2135);
or U1451 (N_1451,In_1423,In_650);
xnor U1452 (N_1452,In_1201,In_2887);
and U1453 (N_1453,In_914,In_2342);
or U1454 (N_1454,In_2223,In_583);
nand U1455 (N_1455,In_2777,In_2486);
nor U1456 (N_1456,In_682,In_509);
and U1457 (N_1457,In_1058,In_2870);
xnor U1458 (N_1458,In_1328,In_674);
and U1459 (N_1459,In_836,In_1801);
nand U1460 (N_1460,In_2294,In_1760);
xnor U1461 (N_1461,In_1951,In_2830);
nand U1462 (N_1462,In_353,In_2199);
nor U1463 (N_1463,In_2578,In_976);
and U1464 (N_1464,In_2572,In_1323);
and U1465 (N_1465,In_2226,In_358);
or U1466 (N_1466,In_853,In_700);
and U1467 (N_1467,In_2158,In_774);
xnor U1468 (N_1468,In_2498,In_1184);
nor U1469 (N_1469,In_768,In_2321);
nor U1470 (N_1470,In_1850,In_2712);
nor U1471 (N_1471,In_1290,In_1868);
or U1472 (N_1472,In_2367,In_258);
and U1473 (N_1473,In_1616,In_2896);
and U1474 (N_1474,In_2145,In_1902);
xor U1475 (N_1475,In_2917,In_1552);
xnor U1476 (N_1476,In_1969,In_2172);
and U1477 (N_1477,In_810,In_1554);
xnor U1478 (N_1478,In_1861,In_2745);
nor U1479 (N_1479,In_1580,In_568);
nor U1480 (N_1480,In_2141,In_941);
or U1481 (N_1481,In_1419,In_2151);
xnor U1482 (N_1482,In_2506,In_2998);
nand U1483 (N_1483,In_2400,In_1447);
and U1484 (N_1484,In_1023,In_942);
nor U1485 (N_1485,In_2838,In_2714);
xnor U1486 (N_1486,In_816,In_2569);
xnor U1487 (N_1487,In_200,In_1188);
and U1488 (N_1488,In_350,In_68);
and U1489 (N_1489,In_1206,In_1334);
nor U1490 (N_1490,In_2026,In_2227);
or U1491 (N_1491,In_2487,In_1319);
nand U1492 (N_1492,In_546,In_2805);
xnor U1493 (N_1493,In_1197,In_326);
nor U1494 (N_1494,In_2990,In_1854);
and U1495 (N_1495,In_1438,In_523);
or U1496 (N_1496,In_2045,In_2469);
or U1497 (N_1497,In_880,In_521);
and U1498 (N_1498,In_1683,In_2963);
xnor U1499 (N_1499,In_2576,In_2881);
nand U1500 (N_1500,In_1649,In_942);
nand U1501 (N_1501,In_1924,In_1301);
nand U1502 (N_1502,In_1800,In_2696);
or U1503 (N_1503,In_675,In_515);
and U1504 (N_1504,In_661,In_1991);
or U1505 (N_1505,In_2159,In_1916);
nand U1506 (N_1506,In_1531,In_647);
xnor U1507 (N_1507,In_1828,In_284);
xnor U1508 (N_1508,In_2499,In_814);
xor U1509 (N_1509,In_373,In_226);
and U1510 (N_1510,In_1976,In_1098);
nor U1511 (N_1511,In_2041,In_2437);
and U1512 (N_1512,In_1776,In_1497);
and U1513 (N_1513,In_725,In_1208);
and U1514 (N_1514,In_568,In_141);
nand U1515 (N_1515,In_297,In_1603);
nand U1516 (N_1516,In_2391,In_2887);
or U1517 (N_1517,In_2431,In_1113);
nand U1518 (N_1518,In_1830,In_1709);
xnor U1519 (N_1519,In_1011,In_1266);
xnor U1520 (N_1520,In_1785,In_2120);
nor U1521 (N_1521,In_614,In_2828);
xor U1522 (N_1522,In_1410,In_1783);
nor U1523 (N_1523,In_2770,In_2086);
nand U1524 (N_1524,In_1210,In_1452);
nand U1525 (N_1525,In_26,In_884);
nand U1526 (N_1526,In_1764,In_2482);
and U1527 (N_1527,In_1876,In_1576);
nor U1528 (N_1528,In_473,In_443);
xnor U1529 (N_1529,In_1598,In_1964);
nand U1530 (N_1530,In_1136,In_329);
or U1531 (N_1531,In_1426,In_1091);
nand U1532 (N_1532,In_2233,In_514);
and U1533 (N_1533,In_2509,In_126);
xnor U1534 (N_1534,In_2347,In_1406);
xor U1535 (N_1535,In_2750,In_1528);
nor U1536 (N_1536,In_172,In_1613);
nand U1537 (N_1537,In_2131,In_2373);
xor U1538 (N_1538,In_2225,In_2668);
nand U1539 (N_1539,In_1360,In_755);
xor U1540 (N_1540,In_2550,In_795);
nor U1541 (N_1541,In_515,In_2533);
or U1542 (N_1542,In_1700,In_1370);
and U1543 (N_1543,In_916,In_1314);
xor U1544 (N_1544,In_315,In_393);
nand U1545 (N_1545,In_1666,In_173);
nor U1546 (N_1546,In_229,In_1952);
and U1547 (N_1547,In_1048,In_1955);
or U1548 (N_1548,In_2095,In_1905);
xor U1549 (N_1549,In_2295,In_1578);
or U1550 (N_1550,In_1166,In_1503);
nand U1551 (N_1551,In_473,In_1635);
or U1552 (N_1552,In_1480,In_1193);
and U1553 (N_1553,In_1020,In_2714);
xnor U1554 (N_1554,In_30,In_2594);
nand U1555 (N_1555,In_1011,In_2217);
xor U1556 (N_1556,In_937,In_423);
nand U1557 (N_1557,In_732,In_2017);
nor U1558 (N_1558,In_1412,In_2732);
nand U1559 (N_1559,In_828,In_1649);
nand U1560 (N_1560,In_795,In_2369);
nand U1561 (N_1561,In_185,In_1459);
or U1562 (N_1562,In_2283,In_2617);
and U1563 (N_1563,In_408,In_2122);
nand U1564 (N_1564,In_2020,In_1558);
xnor U1565 (N_1565,In_169,In_331);
or U1566 (N_1566,In_233,In_2010);
nand U1567 (N_1567,In_2436,In_1176);
nor U1568 (N_1568,In_1082,In_1023);
nand U1569 (N_1569,In_2993,In_917);
xor U1570 (N_1570,In_1916,In_433);
and U1571 (N_1571,In_1389,In_1757);
and U1572 (N_1572,In_242,In_58);
nand U1573 (N_1573,In_2435,In_1122);
nand U1574 (N_1574,In_1805,In_1162);
and U1575 (N_1575,In_423,In_1474);
xor U1576 (N_1576,In_1724,In_1997);
or U1577 (N_1577,In_1567,In_393);
and U1578 (N_1578,In_244,In_448);
nor U1579 (N_1579,In_242,In_2014);
nor U1580 (N_1580,In_2753,In_371);
xnor U1581 (N_1581,In_1801,In_1912);
xnor U1582 (N_1582,In_2622,In_2035);
and U1583 (N_1583,In_1439,In_1799);
and U1584 (N_1584,In_2026,In_1625);
and U1585 (N_1585,In_609,In_2349);
nand U1586 (N_1586,In_1776,In_1263);
nor U1587 (N_1587,In_2811,In_1537);
and U1588 (N_1588,In_925,In_1308);
nand U1589 (N_1589,In_592,In_2106);
nand U1590 (N_1590,In_951,In_1865);
nor U1591 (N_1591,In_2495,In_2782);
or U1592 (N_1592,In_1633,In_2943);
xnor U1593 (N_1593,In_2451,In_548);
nand U1594 (N_1594,In_1837,In_25);
or U1595 (N_1595,In_1422,In_692);
nor U1596 (N_1596,In_2185,In_437);
xor U1597 (N_1597,In_2388,In_2838);
nor U1598 (N_1598,In_2745,In_442);
xnor U1599 (N_1599,In_1029,In_1300);
xor U1600 (N_1600,In_1609,In_2574);
and U1601 (N_1601,In_2388,In_1852);
nand U1602 (N_1602,In_657,In_847);
and U1603 (N_1603,In_2381,In_84);
and U1604 (N_1604,In_1810,In_1752);
or U1605 (N_1605,In_1837,In_2798);
and U1606 (N_1606,In_1538,In_1896);
nor U1607 (N_1607,In_2736,In_2486);
nor U1608 (N_1608,In_2462,In_896);
nor U1609 (N_1609,In_837,In_267);
and U1610 (N_1610,In_2452,In_819);
xor U1611 (N_1611,In_1598,In_2642);
nor U1612 (N_1612,In_2234,In_1445);
nand U1613 (N_1613,In_1585,In_889);
nand U1614 (N_1614,In_699,In_339);
nand U1615 (N_1615,In_816,In_1091);
nor U1616 (N_1616,In_1316,In_1769);
xnor U1617 (N_1617,In_84,In_887);
and U1618 (N_1618,In_1990,In_2131);
xnor U1619 (N_1619,In_502,In_1096);
and U1620 (N_1620,In_1815,In_2062);
and U1621 (N_1621,In_777,In_519);
nand U1622 (N_1622,In_95,In_2792);
nand U1623 (N_1623,In_2861,In_2302);
and U1624 (N_1624,In_2558,In_877);
nand U1625 (N_1625,In_2981,In_2887);
and U1626 (N_1626,In_203,In_1321);
nand U1627 (N_1627,In_1218,In_683);
nand U1628 (N_1628,In_1725,In_1078);
xnor U1629 (N_1629,In_2121,In_1315);
nand U1630 (N_1630,In_999,In_699);
or U1631 (N_1631,In_317,In_2418);
nand U1632 (N_1632,In_923,In_887);
and U1633 (N_1633,In_1370,In_875);
nand U1634 (N_1634,In_1530,In_2999);
and U1635 (N_1635,In_1895,In_373);
and U1636 (N_1636,In_2584,In_778);
and U1637 (N_1637,In_637,In_2804);
and U1638 (N_1638,In_837,In_2552);
or U1639 (N_1639,In_2705,In_1145);
and U1640 (N_1640,In_2276,In_1277);
nand U1641 (N_1641,In_49,In_1546);
nor U1642 (N_1642,In_1328,In_183);
nor U1643 (N_1643,In_956,In_1545);
or U1644 (N_1644,In_1546,In_497);
nor U1645 (N_1645,In_1268,In_577);
nand U1646 (N_1646,In_324,In_2672);
nor U1647 (N_1647,In_621,In_412);
and U1648 (N_1648,In_221,In_1250);
and U1649 (N_1649,In_2252,In_1675);
and U1650 (N_1650,In_489,In_2240);
xnor U1651 (N_1651,In_366,In_2529);
xor U1652 (N_1652,In_2431,In_562);
xnor U1653 (N_1653,In_715,In_2994);
nand U1654 (N_1654,In_432,In_1388);
and U1655 (N_1655,In_1070,In_104);
nor U1656 (N_1656,In_352,In_551);
xor U1657 (N_1657,In_823,In_1976);
or U1658 (N_1658,In_2561,In_2431);
or U1659 (N_1659,In_1764,In_2735);
nor U1660 (N_1660,In_9,In_1190);
xnor U1661 (N_1661,In_90,In_920);
nor U1662 (N_1662,In_2342,In_1534);
nor U1663 (N_1663,In_2426,In_605);
xor U1664 (N_1664,In_1898,In_481);
and U1665 (N_1665,In_1136,In_1149);
nor U1666 (N_1666,In_1061,In_832);
and U1667 (N_1667,In_2883,In_2495);
or U1668 (N_1668,In_1785,In_1897);
nor U1669 (N_1669,In_2830,In_2418);
and U1670 (N_1670,In_1815,In_2072);
nand U1671 (N_1671,In_635,In_1840);
or U1672 (N_1672,In_2074,In_1248);
nor U1673 (N_1673,In_685,In_2568);
nor U1674 (N_1674,In_1521,In_678);
or U1675 (N_1675,In_1300,In_2621);
nand U1676 (N_1676,In_1413,In_1981);
nand U1677 (N_1677,In_2652,In_608);
or U1678 (N_1678,In_2598,In_2488);
nand U1679 (N_1679,In_1933,In_270);
nand U1680 (N_1680,In_2821,In_722);
nor U1681 (N_1681,In_1983,In_580);
nor U1682 (N_1682,In_386,In_2189);
xor U1683 (N_1683,In_172,In_1841);
nand U1684 (N_1684,In_2985,In_2682);
xor U1685 (N_1685,In_752,In_2568);
nand U1686 (N_1686,In_73,In_1862);
and U1687 (N_1687,In_1988,In_1258);
or U1688 (N_1688,In_485,In_1521);
and U1689 (N_1689,In_480,In_547);
nor U1690 (N_1690,In_113,In_1101);
or U1691 (N_1691,In_2695,In_176);
xnor U1692 (N_1692,In_2433,In_537);
xor U1693 (N_1693,In_2829,In_517);
or U1694 (N_1694,In_504,In_688);
xnor U1695 (N_1695,In_2257,In_166);
nand U1696 (N_1696,In_2629,In_2530);
nand U1697 (N_1697,In_2321,In_2033);
and U1698 (N_1698,In_2630,In_427);
nor U1699 (N_1699,In_689,In_2780);
xor U1700 (N_1700,In_2145,In_990);
xnor U1701 (N_1701,In_1249,In_2852);
or U1702 (N_1702,In_97,In_2337);
and U1703 (N_1703,In_360,In_1414);
nor U1704 (N_1704,In_2886,In_619);
and U1705 (N_1705,In_653,In_2509);
xor U1706 (N_1706,In_1790,In_1014);
or U1707 (N_1707,In_955,In_1062);
and U1708 (N_1708,In_2602,In_288);
and U1709 (N_1709,In_2509,In_2975);
and U1710 (N_1710,In_2700,In_33);
or U1711 (N_1711,In_2941,In_2066);
xor U1712 (N_1712,In_2243,In_373);
and U1713 (N_1713,In_2486,In_563);
xor U1714 (N_1714,In_2542,In_1050);
xor U1715 (N_1715,In_826,In_898);
xnor U1716 (N_1716,In_2146,In_950);
or U1717 (N_1717,In_1377,In_194);
or U1718 (N_1718,In_619,In_2462);
nor U1719 (N_1719,In_989,In_1684);
or U1720 (N_1720,In_837,In_194);
or U1721 (N_1721,In_2100,In_1672);
xnor U1722 (N_1722,In_559,In_1742);
and U1723 (N_1723,In_2240,In_1512);
and U1724 (N_1724,In_833,In_1163);
nor U1725 (N_1725,In_1151,In_2282);
xnor U1726 (N_1726,In_113,In_2073);
and U1727 (N_1727,In_431,In_2235);
xor U1728 (N_1728,In_2466,In_2020);
or U1729 (N_1729,In_909,In_2364);
nor U1730 (N_1730,In_2358,In_532);
nand U1731 (N_1731,In_1912,In_1924);
nand U1732 (N_1732,In_2866,In_1019);
xor U1733 (N_1733,In_1764,In_1390);
and U1734 (N_1734,In_684,In_24);
xnor U1735 (N_1735,In_1099,In_2054);
xnor U1736 (N_1736,In_1397,In_1599);
nor U1737 (N_1737,In_285,In_1553);
xnor U1738 (N_1738,In_1624,In_2549);
and U1739 (N_1739,In_1181,In_803);
nor U1740 (N_1740,In_2961,In_1295);
xnor U1741 (N_1741,In_1653,In_639);
and U1742 (N_1742,In_1744,In_173);
nand U1743 (N_1743,In_1559,In_746);
or U1744 (N_1744,In_1815,In_2323);
nand U1745 (N_1745,In_370,In_1987);
nor U1746 (N_1746,In_617,In_1285);
and U1747 (N_1747,In_1576,In_1382);
or U1748 (N_1748,In_1697,In_2237);
nand U1749 (N_1749,In_50,In_1278);
nand U1750 (N_1750,In_782,In_1246);
nand U1751 (N_1751,In_2437,In_2465);
nand U1752 (N_1752,In_1494,In_837);
nand U1753 (N_1753,In_495,In_2806);
and U1754 (N_1754,In_69,In_864);
xnor U1755 (N_1755,In_1432,In_1845);
nor U1756 (N_1756,In_1230,In_2667);
nor U1757 (N_1757,In_1056,In_2777);
nand U1758 (N_1758,In_280,In_1064);
xnor U1759 (N_1759,In_1355,In_552);
or U1760 (N_1760,In_2097,In_1703);
nand U1761 (N_1761,In_952,In_2569);
or U1762 (N_1762,In_1737,In_2274);
nand U1763 (N_1763,In_2305,In_1969);
nor U1764 (N_1764,In_2276,In_2524);
nand U1765 (N_1765,In_1419,In_2841);
nor U1766 (N_1766,In_12,In_2808);
or U1767 (N_1767,In_512,In_833);
xnor U1768 (N_1768,In_2620,In_2561);
nand U1769 (N_1769,In_308,In_473);
and U1770 (N_1770,In_195,In_1658);
nor U1771 (N_1771,In_2762,In_1905);
or U1772 (N_1772,In_594,In_318);
or U1773 (N_1773,In_2516,In_471);
xor U1774 (N_1774,In_1930,In_1704);
nand U1775 (N_1775,In_2526,In_405);
and U1776 (N_1776,In_2007,In_51);
or U1777 (N_1777,In_179,In_75);
nor U1778 (N_1778,In_2067,In_2209);
nor U1779 (N_1779,In_2538,In_1209);
nor U1780 (N_1780,In_2132,In_1921);
or U1781 (N_1781,In_2508,In_2023);
xnor U1782 (N_1782,In_1767,In_1201);
nand U1783 (N_1783,In_1182,In_636);
nand U1784 (N_1784,In_2236,In_136);
xor U1785 (N_1785,In_654,In_2467);
and U1786 (N_1786,In_1834,In_2085);
nor U1787 (N_1787,In_2895,In_577);
or U1788 (N_1788,In_2639,In_2707);
nor U1789 (N_1789,In_1221,In_208);
and U1790 (N_1790,In_2289,In_2558);
and U1791 (N_1791,In_2756,In_574);
xnor U1792 (N_1792,In_2383,In_1589);
or U1793 (N_1793,In_2461,In_208);
xor U1794 (N_1794,In_612,In_751);
nor U1795 (N_1795,In_2815,In_1510);
or U1796 (N_1796,In_1400,In_2879);
or U1797 (N_1797,In_2720,In_1562);
xor U1798 (N_1798,In_2022,In_2266);
or U1799 (N_1799,In_2409,In_911);
and U1800 (N_1800,In_1893,In_797);
xnor U1801 (N_1801,In_2722,In_2293);
and U1802 (N_1802,In_2577,In_1841);
and U1803 (N_1803,In_33,In_1933);
xnor U1804 (N_1804,In_806,In_2268);
or U1805 (N_1805,In_1164,In_2952);
nand U1806 (N_1806,In_2429,In_1285);
and U1807 (N_1807,In_2761,In_1149);
nand U1808 (N_1808,In_2534,In_2630);
nand U1809 (N_1809,In_1592,In_865);
nand U1810 (N_1810,In_2046,In_2781);
xor U1811 (N_1811,In_226,In_575);
nand U1812 (N_1812,In_1639,In_1654);
nand U1813 (N_1813,In_2220,In_2520);
or U1814 (N_1814,In_1443,In_369);
and U1815 (N_1815,In_1441,In_775);
xnor U1816 (N_1816,In_1768,In_879);
nand U1817 (N_1817,In_2334,In_1556);
or U1818 (N_1818,In_684,In_60);
xor U1819 (N_1819,In_2300,In_564);
and U1820 (N_1820,In_2590,In_2172);
nor U1821 (N_1821,In_2870,In_2954);
or U1822 (N_1822,In_211,In_636);
xor U1823 (N_1823,In_2733,In_2888);
and U1824 (N_1824,In_2962,In_2469);
xor U1825 (N_1825,In_229,In_1696);
or U1826 (N_1826,In_2569,In_190);
xnor U1827 (N_1827,In_142,In_258);
and U1828 (N_1828,In_1762,In_1668);
nor U1829 (N_1829,In_1960,In_1655);
nor U1830 (N_1830,In_2321,In_1710);
and U1831 (N_1831,In_1687,In_2864);
nor U1832 (N_1832,In_2596,In_2418);
xor U1833 (N_1833,In_2260,In_1269);
and U1834 (N_1834,In_1696,In_1864);
xor U1835 (N_1835,In_1208,In_492);
nor U1836 (N_1836,In_2721,In_1667);
nand U1837 (N_1837,In_2393,In_2456);
and U1838 (N_1838,In_2692,In_1197);
and U1839 (N_1839,In_1207,In_1572);
or U1840 (N_1840,In_1353,In_2779);
and U1841 (N_1841,In_2890,In_2089);
nor U1842 (N_1842,In_536,In_783);
and U1843 (N_1843,In_657,In_687);
or U1844 (N_1844,In_580,In_1893);
or U1845 (N_1845,In_1537,In_1141);
or U1846 (N_1846,In_620,In_1681);
xor U1847 (N_1847,In_369,In_1111);
xnor U1848 (N_1848,In_2422,In_1967);
nand U1849 (N_1849,In_1770,In_597);
and U1850 (N_1850,In_44,In_1120);
or U1851 (N_1851,In_682,In_289);
or U1852 (N_1852,In_2088,In_1850);
or U1853 (N_1853,In_2318,In_1811);
xnor U1854 (N_1854,In_2020,In_913);
nor U1855 (N_1855,In_2958,In_21);
xnor U1856 (N_1856,In_1892,In_1781);
nor U1857 (N_1857,In_545,In_1215);
nand U1858 (N_1858,In_1366,In_2260);
or U1859 (N_1859,In_476,In_896);
xor U1860 (N_1860,In_210,In_1132);
nand U1861 (N_1861,In_2554,In_2698);
and U1862 (N_1862,In_1227,In_952);
nand U1863 (N_1863,In_2399,In_830);
nor U1864 (N_1864,In_1793,In_1735);
nand U1865 (N_1865,In_317,In_2802);
nor U1866 (N_1866,In_573,In_622);
and U1867 (N_1867,In_2738,In_1589);
xnor U1868 (N_1868,In_1380,In_2206);
nand U1869 (N_1869,In_2593,In_1207);
and U1870 (N_1870,In_2513,In_279);
or U1871 (N_1871,In_2045,In_1815);
or U1872 (N_1872,In_258,In_2038);
xor U1873 (N_1873,In_1375,In_917);
xor U1874 (N_1874,In_540,In_2100);
and U1875 (N_1875,In_1028,In_991);
xnor U1876 (N_1876,In_970,In_2809);
nand U1877 (N_1877,In_964,In_158);
xnor U1878 (N_1878,In_1007,In_230);
nand U1879 (N_1879,In_1586,In_278);
or U1880 (N_1880,In_1151,In_1436);
and U1881 (N_1881,In_2642,In_253);
or U1882 (N_1882,In_1847,In_357);
xnor U1883 (N_1883,In_979,In_103);
nor U1884 (N_1884,In_1533,In_1922);
or U1885 (N_1885,In_2493,In_1998);
nand U1886 (N_1886,In_1250,In_538);
nand U1887 (N_1887,In_1795,In_1127);
nor U1888 (N_1888,In_1786,In_798);
or U1889 (N_1889,In_679,In_2436);
nand U1890 (N_1890,In_236,In_2011);
nor U1891 (N_1891,In_360,In_1298);
or U1892 (N_1892,In_554,In_2843);
nor U1893 (N_1893,In_1922,In_323);
nand U1894 (N_1894,In_850,In_209);
xnor U1895 (N_1895,In_2400,In_2147);
nor U1896 (N_1896,In_272,In_772);
nand U1897 (N_1897,In_901,In_2120);
and U1898 (N_1898,In_2969,In_938);
and U1899 (N_1899,In_2785,In_1004);
nor U1900 (N_1900,In_1398,In_1767);
nor U1901 (N_1901,In_802,In_2245);
or U1902 (N_1902,In_1134,In_1723);
or U1903 (N_1903,In_1039,In_1013);
nor U1904 (N_1904,In_1479,In_145);
xnor U1905 (N_1905,In_118,In_1944);
or U1906 (N_1906,In_2602,In_2757);
or U1907 (N_1907,In_410,In_1768);
or U1908 (N_1908,In_1960,In_509);
nor U1909 (N_1909,In_2893,In_1428);
and U1910 (N_1910,In_2262,In_599);
nor U1911 (N_1911,In_2764,In_2239);
or U1912 (N_1912,In_2943,In_705);
or U1913 (N_1913,In_1429,In_1360);
xor U1914 (N_1914,In_2165,In_169);
or U1915 (N_1915,In_849,In_1239);
nor U1916 (N_1916,In_2717,In_2611);
xnor U1917 (N_1917,In_2493,In_2828);
or U1918 (N_1918,In_1760,In_158);
and U1919 (N_1919,In_1296,In_1900);
xnor U1920 (N_1920,In_2895,In_26);
or U1921 (N_1921,In_2122,In_428);
nand U1922 (N_1922,In_2193,In_2008);
xnor U1923 (N_1923,In_355,In_2138);
nor U1924 (N_1924,In_2448,In_1156);
xor U1925 (N_1925,In_1439,In_1174);
or U1926 (N_1926,In_58,In_2364);
or U1927 (N_1927,In_348,In_310);
nor U1928 (N_1928,In_1762,In_849);
or U1929 (N_1929,In_1109,In_422);
or U1930 (N_1930,In_989,In_8);
nor U1931 (N_1931,In_1669,In_620);
or U1932 (N_1932,In_377,In_1136);
or U1933 (N_1933,In_1848,In_2255);
and U1934 (N_1934,In_2760,In_1501);
and U1935 (N_1935,In_1907,In_1312);
xor U1936 (N_1936,In_1371,In_359);
or U1937 (N_1937,In_1730,In_2684);
or U1938 (N_1938,In_319,In_1776);
or U1939 (N_1939,In_2837,In_867);
xor U1940 (N_1940,In_1593,In_757);
nor U1941 (N_1941,In_1419,In_1788);
xor U1942 (N_1942,In_509,In_1360);
xnor U1943 (N_1943,In_596,In_1446);
nand U1944 (N_1944,In_2236,In_2538);
nand U1945 (N_1945,In_1102,In_1372);
nand U1946 (N_1946,In_873,In_474);
nor U1947 (N_1947,In_2370,In_324);
nand U1948 (N_1948,In_147,In_319);
and U1949 (N_1949,In_1812,In_179);
nor U1950 (N_1950,In_1823,In_1539);
and U1951 (N_1951,In_2508,In_341);
nand U1952 (N_1952,In_2829,In_1166);
or U1953 (N_1953,In_1161,In_1699);
and U1954 (N_1954,In_2127,In_1655);
or U1955 (N_1955,In_1522,In_2968);
xor U1956 (N_1956,In_68,In_550);
xnor U1957 (N_1957,In_820,In_2410);
xor U1958 (N_1958,In_2399,In_2592);
xnor U1959 (N_1959,In_573,In_2283);
nor U1960 (N_1960,In_2551,In_2890);
and U1961 (N_1961,In_1994,In_1735);
or U1962 (N_1962,In_1083,In_1594);
nor U1963 (N_1963,In_705,In_1757);
or U1964 (N_1964,In_773,In_817);
xnor U1965 (N_1965,In_1326,In_2605);
nor U1966 (N_1966,In_1018,In_2550);
nand U1967 (N_1967,In_1238,In_1756);
nor U1968 (N_1968,In_1754,In_2142);
xnor U1969 (N_1969,In_108,In_1087);
or U1970 (N_1970,In_881,In_273);
or U1971 (N_1971,In_161,In_719);
xor U1972 (N_1972,In_486,In_763);
xor U1973 (N_1973,In_1710,In_2817);
nand U1974 (N_1974,In_969,In_1734);
and U1975 (N_1975,In_1305,In_1228);
nor U1976 (N_1976,In_544,In_14);
and U1977 (N_1977,In_1390,In_2308);
nor U1978 (N_1978,In_1901,In_106);
nand U1979 (N_1979,In_1597,In_2062);
xor U1980 (N_1980,In_361,In_495);
and U1981 (N_1981,In_1851,In_2054);
nor U1982 (N_1982,In_2769,In_1037);
xnor U1983 (N_1983,In_15,In_2760);
nor U1984 (N_1984,In_1203,In_734);
and U1985 (N_1985,In_2066,In_2384);
nor U1986 (N_1986,In_668,In_1614);
nand U1987 (N_1987,In_2482,In_2044);
nor U1988 (N_1988,In_2710,In_2069);
or U1989 (N_1989,In_2425,In_1811);
nand U1990 (N_1990,In_2847,In_222);
and U1991 (N_1991,In_598,In_2655);
and U1992 (N_1992,In_2232,In_1110);
xor U1993 (N_1993,In_1075,In_2089);
xor U1994 (N_1994,In_2016,In_109);
or U1995 (N_1995,In_2060,In_1965);
xor U1996 (N_1996,In_2846,In_1651);
nand U1997 (N_1997,In_370,In_1714);
or U1998 (N_1998,In_823,In_2817);
nand U1999 (N_1999,In_595,In_2375);
xnor U2000 (N_2000,In_1904,In_2489);
nor U2001 (N_2001,In_1955,In_1294);
or U2002 (N_2002,In_1764,In_328);
or U2003 (N_2003,In_285,In_2077);
nor U2004 (N_2004,In_1921,In_536);
nor U2005 (N_2005,In_207,In_2823);
nand U2006 (N_2006,In_745,In_2081);
or U2007 (N_2007,In_2324,In_58);
and U2008 (N_2008,In_479,In_377);
nor U2009 (N_2009,In_2901,In_2655);
nand U2010 (N_2010,In_337,In_2953);
nor U2011 (N_2011,In_1222,In_19);
nand U2012 (N_2012,In_2247,In_949);
and U2013 (N_2013,In_600,In_2581);
xnor U2014 (N_2014,In_1306,In_2703);
xor U2015 (N_2015,In_1264,In_2522);
xor U2016 (N_2016,In_1631,In_1625);
nor U2017 (N_2017,In_1767,In_831);
and U2018 (N_2018,In_2606,In_1007);
and U2019 (N_2019,In_1447,In_2050);
and U2020 (N_2020,In_1142,In_2379);
and U2021 (N_2021,In_1001,In_446);
nand U2022 (N_2022,In_2638,In_345);
or U2023 (N_2023,In_1530,In_519);
and U2024 (N_2024,In_1921,In_1351);
nand U2025 (N_2025,In_2758,In_1064);
xnor U2026 (N_2026,In_1433,In_2699);
xor U2027 (N_2027,In_1458,In_99);
nand U2028 (N_2028,In_362,In_1075);
and U2029 (N_2029,In_2374,In_1929);
nand U2030 (N_2030,In_698,In_2305);
nor U2031 (N_2031,In_2769,In_549);
xnor U2032 (N_2032,In_95,In_2538);
nor U2033 (N_2033,In_2046,In_2975);
nand U2034 (N_2034,In_356,In_2272);
nand U2035 (N_2035,In_541,In_1333);
nor U2036 (N_2036,In_684,In_2193);
nor U2037 (N_2037,In_1281,In_2868);
nand U2038 (N_2038,In_530,In_577);
nor U2039 (N_2039,In_118,In_1508);
or U2040 (N_2040,In_2081,In_1268);
nand U2041 (N_2041,In_2808,In_1490);
and U2042 (N_2042,In_824,In_2814);
nor U2043 (N_2043,In_2115,In_1455);
nor U2044 (N_2044,In_1234,In_2542);
or U2045 (N_2045,In_1962,In_1806);
nor U2046 (N_2046,In_1972,In_879);
or U2047 (N_2047,In_1913,In_885);
xor U2048 (N_2048,In_2532,In_707);
and U2049 (N_2049,In_1297,In_2951);
xnor U2050 (N_2050,In_1973,In_1250);
nand U2051 (N_2051,In_1370,In_1979);
and U2052 (N_2052,In_1844,In_195);
and U2053 (N_2053,In_775,In_534);
or U2054 (N_2054,In_1305,In_1921);
nand U2055 (N_2055,In_1753,In_605);
nand U2056 (N_2056,In_2007,In_1312);
nor U2057 (N_2057,In_606,In_1288);
nand U2058 (N_2058,In_1869,In_343);
or U2059 (N_2059,In_2390,In_2688);
and U2060 (N_2060,In_589,In_1652);
nor U2061 (N_2061,In_912,In_2278);
nor U2062 (N_2062,In_2067,In_1281);
nand U2063 (N_2063,In_178,In_950);
xnor U2064 (N_2064,In_422,In_2660);
nand U2065 (N_2065,In_1087,In_1147);
nand U2066 (N_2066,In_1278,In_2002);
nor U2067 (N_2067,In_2592,In_1051);
and U2068 (N_2068,In_1362,In_1573);
xnor U2069 (N_2069,In_1431,In_1336);
nor U2070 (N_2070,In_1100,In_785);
xor U2071 (N_2071,In_901,In_2473);
nor U2072 (N_2072,In_2328,In_1017);
nor U2073 (N_2073,In_2907,In_2218);
xnor U2074 (N_2074,In_430,In_283);
or U2075 (N_2075,In_2255,In_2280);
nor U2076 (N_2076,In_1027,In_2371);
and U2077 (N_2077,In_387,In_619);
and U2078 (N_2078,In_2506,In_2241);
and U2079 (N_2079,In_1900,In_39);
and U2080 (N_2080,In_406,In_1646);
xnor U2081 (N_2081,In_961,In_2973);
and U2082 (N_2082,In_2663,In_2691);
or U2083 (N_2083,In_2721,In_1461);
xnor U2084 (N_2084,In_1298,In_862);
and U2085 (N_2085,In_585,In_2385);
xor U2086 (N_2086,In_803,In_1847);
or U2087 (N_2087,In_1199,In_2225);
and U2088 (N_2088,In_1211,In_2371);
and U2089 (N_2089,In_745,In_1626);
and U2090 (N_2090,In_68,In_2489);
and U2091 (N_2091,In_394,In_1271);
or U2092 (N_2092,In_1100,In_1788);
and U2093 (N_2093,In_2546,In_1569);
and U2094 (N_2094,In_975,In_2212);
or U2095 (N_2095,In_1812,In_1707);
nor U2096 (N_2096,In_2381,In_2824);
nand U2097 (N_2097,In_951,In_1134);
and U2098 (N_2098,In_2682,In_2154);
nor U2099 (N_2099,In_1502,In_2625);
and U2100 (N_2100,In_1548,In_386);
nor U2101 (N_2101,In_246,In_311);
nor U2102 (N_2102,In_2725,In_602);
xor U2103 (N_2103,In_2688,In_1552);
xor U2104 (N_2104,In_2467,In_183);
nor U2105 (N_2105,In_1752,In_714);
nand U2106 (N_2106,In_484,In_1564);
nor U2107 (N_2107,In_41,In_2185);
nor U2108 (N_2108,In_1629,In_758);
xnor U2109 (N_2109,In_2600,In_87);
and U2110 (N_2110,In_135,In_722);
xnor U2111 (N_2111,In_1717,In_1847);
and U2112 (N_2112,In_1074,In_2038);
or U2113 (N_2113,In_786,In_1738);
or U2114 (N_2114,In_729,In_165);
nor U2115 (N_2115,In_55,In_88);
and U2116 (N_2116,In_2326,In_265);
nor U2117 (N_2117,In_93,In_208);
and U2118 (N_2118,In_2152,In_1668);
or U2119 (N_2119,In_296,In_2509);
or U2120 (N_2120,In_831,In_896);
xor U2121 (N_2121,In_878,In_318);
xnor U2122 (N_2122,In_19,In_376);
nand U2123 (N_2123,In_2222,In_154);
nand U2124 (N_2124,In_963,In_2797);
or U2125 (N_2125,In_1450,In_945);
or U2126 (N_2126,In_1106,In_427);
nand U2127 (N_2127,In_1946,In_1489);
or U2128 (N_2128,In_2251,In_2200);
and U2129 (N_2129,In_2878,In_1535);
nor U2130 (N_2130,In_383,In_1859);
and U2131 (N_2131,In_2997,In_756);
nor U2132 (N_2132,In_1577,In_492);
nand U2133 (N_2133,In_2705,In_2840);
and U2134 (N_2134,In_1495,In_152);
nor U2135 (N_2135,In_1378,In_2696);
xor U2136 (N_2136,In_2527,In_228);
and U2137 (N_2137,In_531,In_1881);
nand U2138 (N_2138,In_2161,In_1144);
nand U2139 (N_2139,In_585,In_1705);
or U2140 (N_2140,In_93,In_2213);
nor U2141 (N_2141,In_1909,In_577);
xor U2142 (N_2142,In_1254,In_2241);
xnor U2143 (N_2143,In_1111,In_2467);
or U2144 (N_2144,In_15,In_1178);
nor U2145 (N_2145,In_805,In_1145);
nor U2146 (N_2146,In_1254,In_1596);
nor U2147 (N_2147,In_1640,In_2715);
nand U2148 (N_2148,In_2076,In_519);
nand U2149 (N_2149,In_1102,In_2932);
or U2150 (N_2150,In_2915,In_2660);
nor U2151 (N_2151,In_1399,In_2670);
xor U2152 (N_2152,In_971,In_1408);
or U2153 (N_2153,In_1959,In_384);
nand U2154 (N_2154,In_1967,In_760);
and U2155 (N_2155,In_1636,In_2005);
nor U2156 (N_2156,In_1120,In_1075);
nand U2157 (N_2157,In_2592,In_1695);
nor U2158 (N_2158,In_1585,In_1809);
xnor U2159 (N_2159,In_1391,In_2667);
or U2160 (N_2160,In_1102,In_261);
nand U2161 (N_2161,In_116,In_2427);
and U2162 (N_2162,In_1415,In_1270);
nand U2163 (N_2163,In_638,In_2764);
xnor U2164 (N_2164,In_2608,In_488);
or U2165 (N_2165,In_677,In_124);
xnor U2166 (N_2166,In_1853,In_257);
or U2167 (N_2167,In_2401,In_946);
nor U2168 (N_2168,In_395,In_2813);
xnor U2169 (N_2169,In_965,In_607);
nor U2170 (N_2170,In_636,In_1669);
and U2171 (N_2171,In_266,In_2308);
xor U2172 (N_2172,In_480,In_977);
and U2173 (N_2173,In_1622,In_2784);
nand U2174 (N_2174,In_2045,In_1387);
xnor U2175 (N_2175,In_1645,In_2179);
or U2176 (N_2176,In_194,In_763);
or U2177 (N_2177,In_1374,In_44);
nand U2178 (N_2178,In_2608,In_2554);
nand U2179 (N_2179,In_1153,In_1579);
nor U2180 (N_2180,In_2791,In_2459);
and U2181 (N_2181,In_2351,In_820);
or U2182 (N_2182,In_1250,In_104);
nand U2183 (N_2183,In_1498,In_1124);
nand U2184 (N_2184,In_2475,In_2048);
nor U2185 (N_2185,In_1612,In_1855);
or U2186 (N_2186,In_1887,In_1440);
or U2187 (N_2187,In_137,In_1387);
or U2188 (N_2188,In_1259,In_2032);
and U2189 (N_2189,In_1173,In_2697);
nor U2190 (N_2190,In_2173,In_105);
nand U2191 (N_2191,In_1470,In_121);
xor U2192 (N_2192,In_33,In_375);
and U2193 (N_2193,In_279,In_1599);
xor U2194 (N_2194,In_2700,In_2426);
xor U2195 (N_2195,In_2250,In_965);
xnor U2196 (N_2196,In_1448,In_1503);
xor U2197 (N_2197,In_2866,In_2405);
nor U2198 (N_2198,In_603,In_2891);
nand U2199 (N_2199,In_18,In_1464);
xnor U2200 (N_2200,In_2489,In_2506);
nand U2201 (N_2201,In_1349,In_224);
xor U2202 (N_2202,In_375,In_2841);
nor U2203 (N_2203,In_2620,In_349);
nor U2204 (N_2204,In_2367,In_707);
and U2205 (N_2205,In_2158,In_1581);
nand U2206 (N_2206,In_1128,In_769);
nor U2207 (N_2207,In_1011,In_456);
nand U2208 (N_2208,In_1206,In_1928);
nor U2209 (N_2209,In_648,In_2712);
xor U2210 (N_2210,In_411,In_1033);
nand U2211 (N_2211,In_2401,In_2071);
or U2212 (N_2212,In_1500,In_1678);
nand U2213 (N_2213,In_70,In_742);
nand U2214 (N_2214,In_2245,In_1332);
and U2215 (N_2215,In_696,In_1249);
nor U2216 (N_2216,In_1020,In_2955);
and U2217 (N_2217,In_2248,In_2552);
nand U2218 (N_2218,In_1128,In_1199);
nor U2219 (N_2219,In_249,In_2927);
nor U2220 (N_2220,In_1468,In_2371);
nor U2221 (N_2221,In_2047,In_2791);
nor U2222 (N_2222,In_357,In_2263);
and U2223 (N_2223,In_1919,In_1733);
or U2224 (N_2224,In_2209,In_620);
nor U2225 (N_2225,In_666,In_234);
nor U2226 (N_2226,In_1560,In_705);
nor U2227 (N_2227,In_1661,In_2585);
nand U2228 (N_2228,In_256,In_2245);
nand U2229 (N_2229,In_59,In_618);
and U2230 (N_2230,In_614,In_99);
nand U2231 (N_2231,In_648,In_2248);
and U2232 (N_2232,In_70,In_1600);
xor U2233 (N_2233,In_1094,In_8);
nand U2234 (N_2234,In_909,In_2403);
or U2235 (N_2235,In_1857,In_302);
nand U2236 (N_2236,In_1791,In_2787);
xor U2237 (N_2237,In_1344,In_2299);
or U2238 (N_2238,In_2704,In_2790);
and U2239 (N_2239,In_1647,In_756);
or U2240 (N_2240,In_1590,In_540);
nor U2241 (N_2241,In_1765,In_1713);
xnor U2242 (N_2242,In_2162,In_76);
or U2243 (N_2243,In_1848,In_2301);
nor U2244 (N_2244,In_1886,In_1522);
nor U2245 (N_2245,In_666,In_1559);
xor U2246 (N_2246,In_49,In_2067);
nor U2247 (N_2247,In_395,In_1760);
or U2248 (N_2248,In_2514,In_181);
xnor U2249 (N_2249,In_1954,In_2831);
nor U2250 (N_2250,In_1686,In_2174);
and U2251 (N_2251,In_203,In_802);
or U2252 (N_2252,In_978,In_194);
or U2253 (N_2253,In_291,In_953);
nor U2254 (N_2254,In_783,In_2228);
or U2255 (N_2255,In_1565,In_2347);
and U2256 (N_2256,In_756,In_385);
nand U2257 (N_2257,In_310,In_2324);
xor U2258 (N_2258,In_2848,In_1655);
nor U2259 (N_2259,In_1944,In_505);
xor U2260 (N_2260,In_783,In_769);
xnor U2261 (N_2261,In_2961,In_2705);
or U2262 (N_2262,In_2830,In_130);
and U2263 (N_2263,In_908,In_859);
and U2264 (N_2264,In_1341,In_2185);
nor U2265 (N_2265,In_627,In_1403);
nor U2266 (N_2266,In_429,In_1462);
and U2267 (N_2267,In_2960,In_546);
xor U2268 (N_2268,In_1197,In_1770);
nand U2269 (N_2269,In_2331,In_2538);
nor U2270 (N_2270,In_2826,In_902);
xnor U2271 (N_2271,In_782,In_415);
or U2272 (N_2272,In_314,In_1313);
nand U2273 (N_2273,In_907,In_1708);
nor U2274 (N_2274,In_1372,In_532);
nand U2275 (N_2275,In_1944,In_2394);
nand U2276 (N_2276,In_2087,In_2919);
or U2277 (N_2277,In_380,In_1452);
or U2278 (N_2278,In_423,In_199);
or U2279 (N_2279,In_2127,In_2438);
xor U2280 (N_2280,In_482,In_855);
nor U2281 (N_2281,In_2824,In_654);
or U2282 (N_2282,In_576,In_2701);
nor U2283 (N_2283,In_475,In_1796);
xnor U2284 (N_2284,In_1064,In_2720);
nand U2285 (N_2285,In_15,In_1128);
nand U2286 (N_2286,In_2691,In_377);
or U2287 (N_2287,In_2312,In_379);
nand U2288 (N_2288,In_1674,In_2501);
or U2289 (N_2289,In_1665,In_2628);
nor U2290 (N_2290,In_1186,In_1393);
nor U2291 (N_2291,In_932,In_2188);
or U2292 (N_2292,In_1941,In_2514);
nand U2293 (N_2293,In_2433,In_71);
xor U2294 (N_2294,In_1876,In_152);
nor U2295 (N_2295,In_51,In_675);
or U2296 (N_2296,In_1950,In_1962);
nand U2297 (N_2297,In_1301,In_2730);
nor U2298 (N_2298,In_1808,In_1223);
nor U2299 (N_2299,In_2210,In_2364);
xor U2300 (N_2300,In_1021,In_778);
nor U2301 (N_2301,In_941,In_818);
and U2302 (N_2302,In_2689,In_1220);
xnor U2303 (N_2303,In_2592,In_2252);
nand U2304 (N_2304,In_560,In_2885);
and U2305 (N_2305,In_1505,In_813);
xor U2306 (N_2306,In_827,In_2453);
nand U2307 (N_2307,In_2991,In_2928);
nand U2308 (N_2308,In_717,In_2794);
nand U2309 (N_2309,In_1870,In_558);
and U2310 (N_2310,In_1231,In_2286);
nand U2311 (N_2311,In_755,In_2211);
nand U2312 (N_2312,In_55,In_2238);
nor U2313 (N_2313,In_745,In_2316);
nand U2314 (N_2314,In_1911,In_2812);
xor U2315 (N_2315,In_729,In_1594);
and U2316 (N_2316,In_834,In_2919);
nor U2317 (N_2317,In_948,In_2999);
nor U2318 (N_2318,In_2762,In_2838);
and U2319 (N_2319,In_2315,In_276);
nand U2320 (N_2320,In_1772,In_2794);
nand U2321 (N_2321,In_596,In_2662);
and U2322 (N_2322,In_597,In_2966);
xor U2323 (N_2323,In_1943,In_696);
nor U2324 (N_2324,In_850,In_1625);
nand U2325 (N_2325,In_1169,In_2359);
or U2326 (N_2326,In_49,In_1663);
and U2327 (N_2327,In_1801,In_2152);
and U2328 (N_2328,In_2785,In_1985);
xnor U2329 (N_2329,In_143,In_2793);
and U2330 (N_2330,In_342,In_1141);
or U2331 (N_2331,In_415,In_2408);
xor U2332 (N_2332,In_981,In_2100);
nor U2333 (N_2333,In_782,In_449);
and U2334 (N_2334,In_1287,In_2243);
or U2335 (N_2335,In_584,In_381);
or U2336 (N_2336,In_2076,In_337);
xnor U2337 (N_2337,In_358,In_2740);
nand U2338 (N_2338,In_1407,In_1158);
xnor U2339 (N_2339,In_1296,In_1809);
nand U2340 (N_2340,In_55,In_523);
nand U2341 (N_2341,In_110,In_2524);
or U2342 (N_2342,In_962,In_1929);
and U2343 (N_2343,In_632,In_2865);
nor U2344 (N_2344,In_2705,In_568);
nand U2345 (N_2345,In_1058,In_1593);
or U2346 (N_2346,In_95,In_1449);
and U2347 (N_2347,In_2140,In_2127);
nand U2348 (N_2348,In_774,In_1682);
nor U2349 (N_2349,In_513,In_1784);
nand U2350 (N_2350,In_2927,In_1259);
xnor U2351 (N_2351,In_2124,In_796);
nand U2352 (N_2352,In_1773,In_1818);
nand U2353 (N_2353,In_2340,In_2930);
and U2354 (N_2354,In_3,In_731);
nand U2355 (N_2355,In_2348,In_79);
or U2356 (N_2356,In_527,In_2622);
or U2357 (N_2357,In_2155,In_2080);
nand U2358 (N_2358,In_56,In_1308);
and U2359 (N_2359,In_1715,In_2430);
xor U2360 (N_2360,In_2288,In_1747);
or U2361 (N_2361,In_718,In_1503);
and U2362 (N_2362,In_49,In_1372);
nand U2363 (N_2363,In_327,In_459);
and U2364 (N_2364,In_920,In_323);
nor U2365 (N_2365,In_713,In_638);
and U2366 (N_2366,In_515,In_993);
nand U2367 (N_2367,In_888,In_1594);
nor U2368 (N_2368,In_2644,In_2275);
xor U2369 (N_2369,In_2690,In_2098);
and U2370 (N_2370,In_2068,In_138);
xor U2371 (N_2371,In_1696,In_558);
nor U2372 (N_2372,In_546,In_481);
nand U2373 (N_2373,In_1638,In_1091);
xor U2374 (N_2374,In_1688,In_1720);
xnor U2375 (N_2375,In_1634,In_753);
xor U2376 (N_2376,In_2539,In_866);
or U2377 (N_2377,In_1899,In_720);
xor U2378 (N_2378,In_1436,In_541);
xor U2379 (N_2379,In_1235,In_2038);
and U2380 (N_2380,In_2526,In_410);
and U2381 (N_2381,In_1325,In_2947);
nor U2382 (N_2382,In_1010,In_50);
xnor U2383 (N_2383,In_983,In_1307);
and U2384 (N_2384,In_1543,In_422);
and U2385 (N_2385,In_343,In_62);
nor U2386 (N_2386,In_2462,In_378);
nand U2387 (N_2387,In_2157,In_1426);
nor U2388 (N_2388,In_842,In_22);
xnor U2389 (N_2389,In_2516,In_2460);
nor U2390 (N_2390,In_1226,In_367);
xnor U2391 (N_2391,In_2939,In_1292);
nand U2392 (N_2392,In_2827,In_2096);
or U2393 (N_2393,In_1919,In_2086);
and U2394 (N_2394,In_2133,In_2275);
or U2395 (N_2395,In_122,In_2244);
and U2396 (N_2396,In_741,In_2945);
xnor U2397 (N_2397,In_1945,In_272);
nand U2398 (N_2398,In_120,In_2541);
and U2399 (N_2399,In_2238,In_1780);
xnor U2400 (N_2400,In_2879,In_2554);
xnor U2401 (N_2401,In_2068,In_383);
and U2402 (N_2402,In_1763,In_1972);
or U2403 (N_2403,In_1978,In_1889);
nor U2404 (N_2404,In_1012,In_1754);
or U2405 (N_2405,In_529,In_2944);
nand U2406 (N_2406,In_1281,In_2429);
nor U2407 (N_2407,In_2031,In_897);
nor U2408 (N_2408,In_911,In_1088);
nor U2409 (N_2409,In_1346,In_1776);
xor U2410 (N_2410,In_2442,In_2085);
nand U2411 (N_2411,In_754,In_789);
or U2412 (N_2412,In_1289,In_2909);
and U2413 (N_2413,In_97,In_2214);
xnor U2414 (N_2414,In_464,In_1675);
nor U2415 (N_2415,In_242,In_1848);
and U2416 (N_2416,In_1760,In_2491);
and U2417 (N_2417,In_1755,In_85);
or U2418 (N_2418,In_2897,In_1606);
nand U2419 (N_2419,In_2618,In_683);
xor U2420 (N_2420,In_2675,In_337);
nor U2421 (N_2421,In_1728,In_1604);
xnor U2422 (N_2422,In_1690,In_1913);
and U2423 (N_2423,In_1375,In_1087);
and U2424 (N_2424,In_305,In_443);
nor U2425 (N_2425,In_2121,In_2915);
xnor U2426 (N_2426,In_1226,In_674);
nand U2427 (N_2427,In_1390,In_1165);
or U2428 (N_2428,In_2802,In_933);
xnor U2429 (N_2429,In_823,In_873);
and U2430 (N_2430,In_2183,In_691);
nor U2431 (N_2431,In_1016,In_1642);
nor U2432 (N_2432,In_2908,In_707);
or U2433 (N_2433,In_1904,In_2093);
xnor U2434 (N_2434,In_1160,In_1190);
and U2435 (N_2435,In_2850,In_1364);
nand U2436 (N_2436,In_1958,In_1849);
xnor U2437 (N_2437,In_1348,In_910);
xor U2438 (N_2438,In_2894,In_740);
nand U2439 (N_2439,In_2898,In_2941);
or U2440 (N_2440,In_1923,In_530);
nand U2441 (N_2441,In_1479,In_2179);
or U2442 (N_2442,In_1390,In_1497);
or U2443 (N_2443,In_618,In_435);
nand U2444 (N_2444,In_372,In_2745);
xnor U2445 (N_2445,In_2223,In_2387);
nor U2446 (N_2446,In_2166,In_2285);
nand U2447 (N_2447,In_279,In_442);
and U2448 (N_2448,In_870,In_2730);
nand U2449 (N_2449,In_1368,In_2821);
or U2450 (N_2450,In_2516,In_2151);
nor U2451 (N_2451,In_2418,In_496);
nand U2452 (N_2452,In_602,In_2502);
or U2453 (N_2453,In_1616,In_2395);
and U2454 (N_2454,In_1957,In_1137);
or U2455 (N_2455,In_458,In_1555);
nor U2456 (N_2456,In_2581,In_2627);
xor U2457 (N_2457,In_1703,In_433);
or U2458 (N_2458,In_1588,In_2311);
nor U2459 (N_2459,In_2579,In_2568);
xor U2460 (N_2460,In_10,In_155);
xnor U2461 (N_2461,In_73,In_342);
nor U2462 (N_2462,In_118,In_1953);
nor U2463 (N_2463,In_1059,In_1673);
nor U2464 (N_2464,In_1903,In_1522);
and U2465 (N_2465,In_2788,In_2954);
nand U2466 (N_2466,In_1350,In_2609);
and U2467 (N_2467,In_2369,In_2468);
nor U2468 (N_2468,In_2262,In_777);
or U2469 (N_2469,In_899,In_1922);
nor U2470 (N_2470,In_709,In_1518);
xnor U2471 (N_2471,In_2874,In_461);
nor U2472 (N_2472,In_290,In_2479);
nand U2473 (N_2473,In_371,In_226);
and U2474 (N_2474,In_1849,In_1905);
and U2475 (N_2475,In_2752,In_164);
or U2476 (N_2476,In_2232,In_2100);
nor U2477 (N_2477,In_1183,In_338);
nor U2478 (N_2478,In_1298,In_2701);
or U2479 (N_2479,In_1064,In_1927);
nand U2480 (N_2480,In_560,In_2995);
nand U2481 (N_2481,In_947,In_2545);
or U2482 (N_2482,In_2374,In_2648);
nand U2483 (N_2483,In_338,In_1738);
nor U2484 (N_2484,In_991,In_1018);
and U2485 (N_2485,In_539,In_1774);
xor U2486 (N_2486,In_2130,In_2014);
nand U2487 (N_2487,In_2980,In_310);
and U2488 (N_2488,In_1881,In_604);
xor U2489 (N_2489,In_2879,In_2065);
xnor U2490 (N_2490,In_1995,In_1742);
nor U2491 (N_2491,In_1033,In_625);
nand U2492 (N_2492,In_2110,In_2122);
nand U2493 (N_2493,In_1408,In_1823);
or U2494 (N_2494,In_2618,In_372);
nor U2495 (N_2495,In_1506,In_1397);
or U2496 (N_2496,In_1264,In_1646);
and U2497 (N_2497,In_2911,In_2600);
nor U2498 (N_2498,In_1245,In_1855);
or U2499 (N_2499,In_1491,In_2580);
xor U2500 (N_2500,In_2391,In_1500);
xor U2501 (N_2501,In_1754,In_1214);
nand U2502 (N_2502,In_1558,In_1337);
xor U2503 (N_2503,In_161,In_809);
and U2504 (N_2504,In_1264,In_366);
xor U2505 (N_2505,In_2979,In_786);
nand U2506 (N_2506,In_2557,In_327);
or U2507 (N_2507,In_1015,In_428);
nand U2508 (N_2508,In_1891,In_2035);
xor U2509 (N_2509,In_937,In_2129);
xnor U2510 (N_2510,In_2930,In_1866);
or U2511 (N_2511,In_848,In_780);
nor U2512 (N_2512,In_299,In_1095);
and U2513 (N_2513,In_1445,In_737);
nor U2514 (N_2514,In_2745,In_2204);
nor U2515 (N_2515,In_640,In_1398);
or U2516 (N_2516,In_1747,In_581);
and U2517 (N_2517,In_1881,In_2877);
nor U2518 (N_2518,In_1215,In_2244);
or U2519 (N_2519,In_1714,In_1395);
and U2520 (N_2520,In_2474,In_1004);
nand U2521 (N_2521,In_764,In_1050);
nand U2522 (N_2522,In_1028,In_835);
nand U2523 (N_2523,In_1674,In_322);
and U2524 (N_2524,In_2791,In_518);
xor U2525 (N_2525,In_2896,In_1087);
nand U2526 (N_2526,In_2908,In_2382);
xnor U2527 (N_2527,In_681,In_1913);
nand U2528 (N_2528,In_117,In_2855);
or U2529 (N_2529,In_1274,In_1495);
xnor U2530 (N_2530,In_852,In_847);
xor U2531 (N_2531,In_2906,In_2637);
nand U2532 (N_2532,In_745,In_1774);
and U2533 (N_2533,In_1034,In_909);
xor U2534 (N_2534,In_2874,In_36);
nand U2535 (N_2535,In_441,In_1183);
nand U2536 (N_2536,In_1191,In_2683);
nor U2537 (N_2537,In_1812,In_625);
nor U2538 (N_2538,In_2378,In_444);
nand U2539 (N_2539,In_360,In_1726);
and U2540 (N_2540,In_1741,In_38);
xor U2541 (N_2541,In_1933,In_152);
or U2542 (N_2542,In_2419,In_520);
or U2543 (N_2543,In_1341,In_1718);
xor U2544 (N_2544,In_1691,In_1517);
and U2545 (N_2545,In_1564,In_782);
nand U2546 (N_2546,In_1215,In_2785);
nor U2547 (N_2547,In_814,In_1469);
nand U2548 (N_2548,In_1938,In_1672);
nor U2549 (N_2549,In_1404,In_2560);
xnor U2550 (N_2550,In_1173,In_1520);
nor U2551 (N_2551,In_1364,In_77);
xor U2552 (N_2552,In_568,In_1650);
and U2553 (N_2553,In_481,In_1507);
or U2554 (N_2554,In_1108,In_2017);
nor U2555 (N_2555,In_2983,In_1917);
and U2556 (N_2556,In_1519,In_1343);
nand U2557 (N_2557,In_2026,In_354);
or U2558 (N_2558,In_964,In_360);
nand U2559 (N_2559,In_1711,In_880);
and U2560 (N_2560,In_949,In_352);
nand U2561 (N_2561,In_1899,In_94);
nor U2562 (N_2562,In_2552,In_1887);
nor U2563 (N_2563,In_956,In_208);
or U2564 (N_2564,In_662,In_469);
or U2565 (N_2565,In_2545,In_2692);
and U2566 (N_2566,In_1951,In_375);
and U2567 (N_2567,In_1356,In_1165);
and U2568 (N_2568,In_2254,In_1607);
and U2569 (N_2569,In_414,In_1333);
and U2570 (N_2570,In_2200,In_1517);
nand U2571 (N_2571,In_1052,In_2591);
xnor U2572 (N_2572,In_1408,In_1714);
or U2573 (N_2573,In_811,In_1141);
nand U2574 (N_2574,In_2083,In_2068);
nor U2575 (N_2575,In_1834,In_985);
nand U2576 (N_2576,In_1251,In_378);
nor U2577 (N_2577,In_2459,In_2131);
xor U2578 (N_2578,In_320,In_309);
and U2579 (N_2579,In_2521,In_335);
nand U2580 (N_2580,In_1795,In_1543);
and U2581 (N_2581,In_2412,In_342);
and U2582 (N_2582,In_2916,In_1115);
and U2583 (N_2583,In_2615,In_997);
or U2584 (N_2584,In_1458,In_2268);
or U2585 (N_2585,In_474,In_1190);
xor U2586 (N_2586,In_2962,In_1897);
nor U2587 (N_2587,In_2328,In_2575);
nand U2588 (N_2588,In_431,In_2427);
and U2589 (N_2589,In_339,In_1885);
or U2590 (N_2590,In_1790,In_2652);
nor U2591 (N_2591,In_653,In_1458);
nand U2592 (N_2592,In_284,In_1587);
xnor U2593 (N_2593,In_1981,In_2391);
or U2594 (N_2594,In_460,In_643);
xnor U2595 (N_2595,In_302,In_927);
nand U2596 (N_2596,In_2690,In_105);
nor U2597 (N_2597,In_2344,In_443);
xor U2598 (N_2598,In_1420,In_2332);
nand U2599 (N_2599,In_25,In_22);
or U2600 (N_2600,In_2402,In_181);
nand U2601 (N_2601,In_701,In_2911);
xor U2602 (N_2602,In_121,In_1043);
and U2603 (N_2603,In_2808,In_1679);
or U2604 (N_2604,In_272,In_73);
nand U2605 (N_2605,In_739,In_2875);
xnor U2606 (N_2606,In_1294,In_2641);
xnor U2607 (N_2607,In_1569,In_2708);
and U2608 (N_2608,In_582,In_1547);
nand U2609 (N_2609,In_1284,In_1662);
nand U2610 (N_2610,In_277,In_1721);
or U2611 (N_2611,In_1147,In_2635);
and U2612 (N_2612,In_1419,In_2560);
xnor U2613 (N_2613,In_1207,In_2714);
xnor U2614 (N_2614,In_1200,In_1247);
and U2615 (N_2615,In_696,In_1646);
and U2616 (N_2616,In_222,In_2972);
nor U2617 (N_2617,In_1000,In_2033);
and U2618 (N_2618,In_2271,In_1749);
nand U2619 (N_2619,In_2538,In_475);
or U2620 (N_2620,In_1667,In_712);
xor U2621 (N_2621,In_2454,In_2755);
nand U2622 (N_2622,In_2793,In_1233);
and U2623 (N_2623,In_512,In_1224);
nand U2624 (N_2624,In_931,In_2085);
or U2625 (N_2625,In_857,In_1512);
or U2626 (N_2626,In_1752,In_1391);
xnor U2627 (N_2627,In_592,In_66);
or U2628 (N_2628,In_541,In_1092);
xnor U2629 (N_2629,In_119,In_1892);
or U2630 (N_2630,In_2740,In_775);
or U2631 (N_2631,In_446,In_2388);
and U2632 (N_2632,In_1939,In_1739);
xor U2633 (N_2633,In_2275,In_219);
nand U2634 (N_2634,In_132,In_997);
nor U2635 (N_2635,In_2146,In_939);
nor U2636 (N_2636,In_2981,In_267);
nor U2637 (N_2637,In_2685,In_1499);
and U2638 (N_2638,In_1759,In_1189);
nand U2639 (N_2639,In_2474,In_755);
nor U2640 (N_2640,In_1751,In_2223);
and U2641 (N_2641,In_1695,In_1270);
xor U2642 (N_2642,In_1102,In_1182);
and U2643 (N_2643,In_2011,In_263);
nor U2644 (N_2644,In_2121,In_2892);
xor U2645 (N_2645,In_1663,In_1749);
nor U2646 (N_2646,In_2926,In_1644);
xnor U2647 (N_2647,In_1345,In_2173);
and U2648 (N_2648,In_2804,In_2105);
xnor U2649 (N_2649,In_1239,In_200);
xnor U2650 (N_2650,In_1912,In_1969);
or U2651 (N_2651,In_2421,In_2313);
or U2652 (N_2652,In_1828,In_1089);
and U2653 (N_2653,In_966,In_1148);
xor U2654 (N_2654,In_1967,In_382);
or U2655 (N_2655,In_2258,In_797);
or U2656 (N_2656,In_1954,In_2531);
xnor U2657 (N_2657,In_2819,In_348);
nand U2658 (N_2658,In_1570,In_1726);
and U2659 (N_2659,In_515,In_569);
xnor U2660 (N_2660,In_2707,In_2873);
and U2661 (N_2661,In_2091,In_1943);
xnor U2662 (N_2662,In_1943,In_604);
or U2663 (N_2663,In_2052,In_2468);
nor U2664 (N_2664,In_1844,In_1369);
xor U2665 (N_2665,In_1218,In_1945);
nor U2666 (N_2666,In_2136,In_2207);
xnor U2667 (N_2667,In_851,In_740);
or U2668 (N_2668,In_2400,In_2897);
or U2669 (N_2669,In_926,In_406);
nand U2670 (N_2670,In_1392,In_1039);
and U2671 (N_2671,In_1156,In_2142);
nor U2672 (N_2672,In_2480,In_1116);
or U2673 (N_2673,In_431,In_1457);
or U2674 (N_2674,In_682,In_2085);
and U2675 (N_2675,In_903,In_2947);
and U2676 (N_2676,In_1052,In_36);
nand U2677 (N_2677,In_12,In_546);
and U2678 (N_2678,In_1209,In_2365);
or U2679 (N_2679,In_2906,In_573);
and U2680 (N_2680,In_2655,In_2085);
and U2681 (N_2681,In_1919,In_358);
and U2682 (N_2682,In_2867,In_1059);
and U2683 (N_2683,In_1274,In_2127);
nor U2684 (N_2684,In_1703,In_865);
nand U2685 (N_2685,In_2232,In_354);
and U2686 (N_2686,In_1449,In_83);
nand U2687 (N_2687,In_1999,In_2148);
nor U2688 (N_2688,In_1837,In_272);
or U2689 (N_2689,In_444,In_2630);
or U2690 (N_2690,In_2478,In_503);
xor U2691 (N_2691,In_814,In_1686);
xor U2692 (N_2692,In_1959,In_2189);
and U2693 (N_2693,In_2359,In_577);
or U2694 (N_2694,In_520,In_1912);
nand U2695 (N_2695,In_211,In_495);
xor U2696 (N_2696,In_2015,In_289);
and U2697 (N_2697,In_2578,In_1058);
and U2698 (N_2698,In_1264,In_2661);
nand U2699 (N_2699,In_253,In_415);
nor U2700 (N_2700,In_2240,In_1593);
nor U2701 (N_2701,In_2371,In_640);
nor U2702 (N_2702,In_301,In_2504);
or U2703 (N_2703,In_1280,In_1377);
nand U2704 (N_2704,In_85,In_1430);
xor U2705 (N_2705,In_2058,In_335);
and U2706 (N_2706,In_1424,In_837);
nor U2707 (N_2707,In_2977,In_264);
xor U2708 (N_2708,In_1330,In_676);
xnor U2709 (N_2709,In_1301,In_2199);
or U2710 (N_2710,In_1027,In_1288);
nand U2711 (N_2711,In_2708,In_2554);
nor U2712 (N_2712,In_590,In_226);
xor U2713 (N_2713,In_2086,In_1738);
xor U2714 (N_2714,In_533,In_1399);
or U2715 (N_2715,In_71,In_1175);
xor U2716 (N_2716,In_827,In_1029);
nand U2717 (N_2717,In_2372,In_2915);
nand U2718 (N_2718,In_2079,In_1419);
nor U2719 (N_2719,In_107,In_166);
or U2720 (N_2720,In_2097,In_1776);
nand U2721 (N_2721,In_2930,In_2275);
nand U2722 (N_2722,In_2601,In_2402);
and U2723 (N_2723,In_2322,In_1105);
nand U2724 (N_2724,In_2578,In_425);
nor U2725 (N_2725,In_362,In_2378);
and U2726 (N_2726,In_667,In_736);
or U2727 (N_2727,In_1808,In_2173);
or U2728 (N_2728,In_2642,In_1865);
or U2729 (N_2729,In_915,In_2854);
nand U2730 (N_2730,In_2468,In_1844);
or U2731 (N_2731,In_1036,In_590);
and U2732 (N_2732,In_218,In_2089);
xor U2733 (N_2733,In_1511,In_381);
or U2734 (N_2734,In_932,In_2085);
xnor U2735 (N_2735,In_528,In_241);
xnor U2736 (N_2736,In_46,In_1391);
nor U2737 (N_2737,In_1803,In_2977);
nor U2738 (N_2738,In_1517,In_2168);
or U2739 (N_2739,In_908,In_2387);
and U2740 (N_2740,In_2393,In_1021);
nor U2741 (N_2741,In_2874,In_432);
nand U2742 (N_2742,In_577,In_265);
or U2743 (N_2743,In_561,In_1290);
or U2744 (N_2744,In_869,In_2880);
or U2745 (N_2745,In_1451,In_2392);
nand U2746 (N_2746,In_2310,In_2309);
or U2747 (N_2747,In_2899,In_340);
nor U2748 (N_2748,In_2744,In_2141);
nor U2749 (N_2749,In_2590,In_443);
and U2750 (N_2750,In_1735,In_634);
nand U2751 (N_2751,In_639,In_749);
and U2752 (N_2752,In_2338,In_840);
nor U2753 (N_2753,In_375,In_2684);
or U2754 (N_2754,In_1780,In_1793);
xor U2755 (N_2755,In_1757,In_614);
nand U2756 (N_2756,In_1557,In_1555);
nor U2757 (N_2757,In_2103,In_2112);
nor U2758 (N_2758,In_1875,In_2091);
xnor U2759 (N_2759,In_531,In_1416);
nor U2760 (N_2760,In_2994,In_2873);
xor U2761 (N_2761,In_2937,In_394);
nor U2762 (N_2762,In_2090,In_1702);
nand U2763 (N_2763,In_2911,In_877);
and U2764 (N_2764,In_659,In_310);
nand U2765 (N_2765,In_1071,In_2579);
nand U2766 (N_2766,In_1129,In_2600);
xnor U2767 (N_2767,In_2081,In_421);
nor U2768 (N_2768,In_354,In_82);
nand U2769 (N_2769,In_1750,In_2728);
nand U2770 (N_2770,In_1791,In_301);
and U2771 (N_2771,In_2508,In_2917);
and U2772 (N_2772,In_2238,In_1693);
xor U2773 (N_2773,In_2698,In_1736);
xor U2774 (N_2774,In_1965,In_47);
nor U2775 (N_2775,In_485,In_1662);
and U2776 (N_2776,In_2882,In_1260);
or U2777 (N_2777,In_2506,In_2708);
or U2778 (N_2778,In_2920,In_706);
xor U2779 (N_2779,In_917,In_1465);
xnor U2780 (N_2780,In_298,In_528);
nor U2781 (N_2781,In_405,In_1700);
or U2782 (N_2782,In_1443,In_436);
or U2783 (N_2783,In_1502,In_1158);
nor U2784 (N_2784,In_1125,In_1531);
nand U2785 (N_2785,In_2986,In_2680);
xnor U2786 (N_2786,In_1793,In_450);
and U2787 (N_2787,In_1602,In_1714);
xor U2788 (N_2788,In_1415,In_265);
or U2789 (N_2789,In_2521,In_2230);
or U2790 (N_2790,In_1251,In_2366);
and U2791 (N_2791,In_406,In_2459);
nand U2792 (N_2792,In_1658,In_1823);
nand U2793 (N_2793,In_2745,In_2485);
nor U2794 (N_2794,In_1868,In_1871);
xnor U2795 (N_2795,In_854,In_2774);
nor U2796 (N_2796,In_1153,In_637);
xor U2797 (N_2797,In_1084,In_1877);
and U2798 (N_2798,In_1920,In_2518);
xnor U2799 (N_2799,In_2558,In_2309);
nand U2800 (N_2800,In_754,In_475);
and U2801 (N_2801,In_563,In_373);
or U2802 (N_2802,In_2414,In_774);
nor U2803 (N_2803,In_2095,In_2878);
xnor U2804 (N_2804,In_857,In_547);
nor U2805 (N_2805,In_2741,In_2946);
nand U2806 (N_2806,In_125,In_1847);
xor U2807 (N_2807,In_1135,In_656);
nand U2808 (N_2808,In_137,In_202);
nor U2809 (N_2809,In_395,In_1460);
nand U2810 (N_2810,In_1630,In_2116);
or U2811 (N_2811,In_577,In_785);
xor U2812 (N_2812,In_751,In_2733);
nand U2813 (N_2813,In_720,In_246);
and U2814 (N_2814,In_147,In_1702);
xnor U2815 (N_2815,In_1116,In_811);
xnor U2816 (N_2816,In_1618,In_1530);
or U2817 (N_2817,In_1147,In_539);
nor U2818 (N_2818,In_1642,In_1710);
xor U2819 (N_2819,In_2039,In_185);
nor U2820 (N_2820,In_373,In_1016);
or U2821 (N_2821,In_196,In_98);
xnor U2822 (N_2822,In_1798,In_523);
or U2823 (N_2823,In_2117,In_2363);
nand U2824 (N_2824,In_2174,In_1809);
xor U2825 (N_2825,In_2909,In_1056);
xnor U2826 (N_2826,In_2645,In_1515);
and U2827 (N_2827,In_283,In_80);
nand U2828 (N_2828,In_193,In_2528);
nand U2829 (N_2829,In_2151,In_1486);
nand U2830 (N_2830,In_886,In_2190);
or U2831 (N_2831,In_1887,In_2006);
nor U2832 (N_2832,In_2919,In_2935);
and U2833 (N_2833,In_2470,In_1234);
or U2834 (N_2834,In_1355,In_2778);
xnor U2835 (N_2835,In_1763,In_2969);
xor U2836 (N_2836,In_2385,In_1310);
or U2837 (N_2837,In_1619,In_1595);
and U2838 (N_2838,In_2940,In_1233);
xnor U2839 (N_2839,In_2101,In_2487);
xor U2840 (N_2840,In_644,In_1803);
xor U2841 (N_2841,In_2889,In_2995);
nor U2842 (N_2842,In_1132,In_1049);
nor U2843 (N_2843,In_1187,In_1145);
xnor U2844 (N_2844,In_230,In_2894);
and U2845 (N_2845,In_466,In_1096);
nand U2846 (N_2846,In_2297,In_987);
xnor U2847 (N_2847,In_837,In_1926);
nor U2848 (N_2848,In_1124,In_1646);
and U2849 (N_2849,In_2332,In_331);
nor U2850 (N_2850,In_1533,In_620);
and U2851 (N_2851,In_1435,In_1219);
nor U2852 (N_2852,In_667,In_2937);
xnor U2853 (N_2853,In_473,In_1715);
and U2854 (N_2854,In_929,In_1603);
and U2855 (N_2855,In_1789,In_1571);
xnor U2856 (N_2856,In_2905,In_2833);
or U2857 (N_2857,In_2200,In_726);
nand U2858 (N_2858,In_1152,In_663);
nand U2859 (N_2859,In_1787,In_178);
xor U2860 (N_2860,In_133,In_2824);
xnor U2861 (N_2861,In_37,In_2424);
nor U2862 (N_2862,In_801,In_1515);
nor U2863 (N_2863,In_1221,In_2853);
and U2864 (N_2864,In_2713,In_422);
xor U2865 (N_2865,In_1112,In_452);
nand U2866 (N_2866,In_490,In_82);
nor U2867 (N_2867,In_831,In_2723);
and U2868 (N_2868,In_2934,In_651);
xor U2869 (N_2869,In_1648,In_997);
and U2870 (N_2870,In_2746,In_761);
and U2871 (N_2871,In_2205,In_2398);
nor U2872 (N_2872,In_1905,In_1265);
xor U2873 (N_2873,In_1926,In_2995);
or U2874 (N_2874,In_2718,In_2932);
nand U2875 (N_2875,In_2444,In_2728);
xor U2876 (N_2876,In_1241,In_2458);
nor U2877 (N_2877,In_676,In_2839);
nor U2878 (N_2878,In_202,In_1128);
or U2879 (N_2879,In_326,In_459);
nor U2880 (N_2880,In_1478,In_802);
and U2881 (N_2881,In_2666,In_2640);
nor U2882 (N_2882,In_1499,In_2761);
xnor U2883 (N_2883,In_1006,In_2102);
nand U2884 (N_2884,In_1802,In_1229);
and U2885 (N_2885,In_979,In_1728);
or U2886 (N_2886,In_871,In_2569);
nor U2887 (N_2887,In_1531,In_1515);
and U2888 (N_2888,In_1277,In_545);
xnor U2889 (N_2889,In_1600,In_2157);
and U2890 (N_2890,In_204,In_1286);
and U2891 (N_2891,In_455,In_1154);
and U2892 (N_2892,In_2699,In_1822);
and U2893 (N_2893,In_179,In_1428);
xor U2894 (N_2894,In_763,In_357);
or U2895 (N_2895,In_2912,In_1921);
nor U2896 (N_2896,In_2906,In_2241);
nand U2897 (N_2897,In_750,In_2024);
and U2898 (N_2898,In_725,In_203);
nand U2899 (N_2899,In_649,In_2385);
and U2900 (N_2900,In_2341,In_1374);
nor U2901 (N_2901,In_1579,In_1080);
nor U2902 (N_2902,In_556,In_2510);
nand U2903 (N_2903,In_358,In_138);
nor U2904 (N_2904,In_2146,In_1057);
xnor U2905 (N_2905,In_718,In_948);
nor U2906 (N_2906,In_1355,In_1023);
nand U2907 (N_2907,In_831,In_1906);
nand U2908 (N_2908,In_2496,In_1226);
or U2909 (N_2909,In_2423,In_754);
or U2910 (N_2910,In_634,In_2066);
and U2911 (N_2911,In_2572,In_1890);
and U2912 (N_2912,In_15,In_1873);
and U2913 (N_2913,In_706,In_1717);
nor U2914 (N_2914,In_974,In_2500);
or U2915 (N_2915,In_519,In_1271);
and U2916 (N_2916,In_608,In_2379);
nand U2917 (N_2917,In_1961,In_812);
nor U2918 (N_2918,In_2007,In_2512);
xor U2919 (N_2919,In_2119,In_1730);
nand U2920 (N_2920,In_1016,In_1210);
nand U2921 (N_2921,In_2748,In_1589);
xor U2922 (N_2922,In_1952,In_28);
or U2923 (N_2923,In_2212,In_15);
nor U2924 (N_2924,In_532,In_2870);
nor U2925 (N_2925,In_1637,In_2959);
and U2926 (N_2926,In_1492,In_1598);
nand U2927 (N_2927,In_1697,In_1187);
xnor U2928 (N_2928,In_1714,In_687);
nor U2929 (N_2929,In_2835,In_246);
nand U2930 (N_2930,In_2821,In_2393);
nor U2931 (N_2931,In_2311,In_1358);
and U2932 (N_2932,In_262,In_2139);
and U2933 (N_2933,In_1522,In_878);
nand U2934 (N_2934,In_161,In_2805);
and U2935 (N_2935,In_2732,In_2780);
xnor U2936 (N_2936,In_1806,In_279);
or U2937 (N_2937,In_1938,In_961);
or U2938 (N_2938,In_1709,In_877);
xnor U2939 (N_2939,In_88,In_235);
nor U2940 (N_2940,In_216,In_2324);
or U2941 (N_2941,In_1430,In_2126);
nand U2942 (N_2942,In_585,In_1142);
nand U2943 (N_2943,In_759,In_243);
nor U2944 (N_2944,In_2513,In_1462);
and U2945 (N_2945,In_240,In_1338);
or U2946 (N_2946,In_2391,In_155);
and U2947 (N_2947,In_1604,In_583);
nand U2948 (N_2948,In_2480,In_2018);
and U2949 (N_2949,In_485,In_660);
nand U2950 (N_2950,In_1584,In_1122);
xor U2951 (N_2951,In_1560,In_1086);
and U2952 (N_2952,In_1881,In_2180);
and U2953 (N_2953,In_2612,In_2908);
nand U2954 (N_2954,In_611,In_996);
and U2955 (N_2955,In_81,In_277);
nand U2956 (N_2956,In_1481,In_1787);
xnor U2957 (N_2957,In_1481,In_2087);
nand U2958 (N_2958,In_700,In_2733);
nor U2959 (N_2959,In_2444,In_561);
nor U2960 (N_2960,In_2994,In_1350);
or U2961 (N_2961,In_428,In_1736);
xor U2962 (N_2962,In_1245,In_523);
xor U2963 (N_2963,In_893,In_277);
nor U2964 (N_2964,In_1947,In_554);
and U2965 (N_2965,In_335,In_2925);
nand U2966 (N_2966,In_1146,In_923);
or U2967 (N_2967,In_2356,In_2655);
nand U2968 (N_2968,In_154,In_2196);
nor U2969 (N_2969,In_122,In_1714);
xor U2970 (N_2970,In_1036,In_2387);
and U2971 (N_2971,In_2212,In_2323);
nand U2972 (N_2972,In_349,In_865);
nor U2973 (N_2973,In_2594,In_2766);
nand U2974 (N_2974,In_2002,In_675);
xor U2975 (N_2975,In_2598,In_2294);
nor U2976 (N_2976,In_252,In_2563);
xnor U2977 (N_2977,In_2439,In_1093);
nand U2978 (N_2978,In_2024,In_2166);
xnor U2979 (N_2979,In_2651,In_1780);
nand U2980 (N_2980,In_2265,In_2292);
nand U2981 (N_2981,In_2414,In_154);
and U2982 (N_2982,In_444,In_2178);
and U2983 (N_2983,In_904,In_515);
nor U2984 (N_2984,In_670,In_2539);
nand U2985 (N_2985,In_1328,In_1926);
or U2986 (N_2986,In_1975,In_961);
nand U2987 (N_2987,In_544,In_1044);
and U2988 (N_2988,In_2986,In_835);
nor U2989 (N_2989,In_1183,In_1384);
xnor U2990 (N_2990,In_470,In_2375);
or U2991 (N_2991,In_2238,In_156);
xnor U2992 (N_2992,In_2220,In_2632);
or U2993 (N_2993,In_854,In_2993);
nor U2994 (N_2994,In_1281,In_585);
nor U2995 (N_2995,In_1675,In_1158);
or U2996 (N_2996,In_2807,In_61);
nor U2997 (N_2997,In_1541,In_2751);
nor U2998 (N_2998,In_75,In_607);
and U2999 (N_2999,In_2779,In_355);
xnor U3000 (N_3000,N_1067,N_2781);
and U3001 (N_3001,N_1682,N_532);
and U3002 (N_3002,N_1114,N_690);
nor U3003 (N_3003,N_1543,N_585);
nor U3004 (N_3004,N_1071,N_2310);
nor U3005 (N_3005,N_2034,N_137);
nor U3006 (N_3006,N_2428,N_1421);
nor U3007 (N_3007,N_1109,N_1342);
nand U3008 (N_3008,N_2268,N_892);
or U3009 (N_3009,N_799,N_1996);
xor U3010 (N_3010,N_903,N_1781);
xor U3011 (N_3011,N_2670,N_1378);
nand U3012 (N_3012,N_2157,N_1398);
and U3013 (N_3013,N_2945,N_164);
and U3014 (N_3014,N_2730,N_272);
xnor U3015 (N_3015,N_2165,N_473);
xnor U3016 (N_3016,N_407,N_901);
and U3017 (N_3017,N_295,N_2671);
or U3018 (N_3018,N_2590,N_27);
nand U3019 (N_3019,N_2028,N_1390);
xor U3020 (N_3020,N_2155,N_2546);
or U3021 (N_3021,N_1040,N_1498);
or U3022 (N_3022,N_2204,N_35);
or U3023 (N_3023,N_2626,N_689);
or U3024 (N_3024,N_1835,N_244);
xor U3025 (N_3025,N_949,N_2122);
nor U3026 (N_3026,N_2870,N_2996);
or U3027 (N_3027,N_933,N_2649);
nand U3028 (N_3028,N_1819,N_1135);
xor U3029 (N_3029,N_308,N_1286);
or U3030 (N_3030,N_2445,N_194);
xor U3031 (N_3031,N_2918,N_1671);
and U3032 (N_3032,N_577,N_1634);
nor U3033 (N_3033,N_2010,N_2568);
nand U3034 (N_3034,N_1593,N_962);
nand U3035 (N_3035,N_2968,N_2624);
or U3036 (N_3036,N_1408,N_2143);
or U3037 (N_3037,N_2422,N_1709);
or U3038 (N_3038,N_725,N_1055);
nand U3039 (N_3039,N_1441,N_2164);
nor U3040 (N_3040,N_876,N_742);
and U3041 (N_3041,N_1233,N_351);
nand U3042 (N_3042,N_78,N_2217);
xnor U3043 (N_3043,N_261,N_1480);
xnor U3044 (N_3044,N_1830,N_961);
or U3045 (N_3045,N_2934,N_2615);
nor U3046 (N_3046,N_1760,N_1504);
xor U3047 (N_3047,N_465,N_2196);
nor U3048 (N_3048,N_2186,N_1918);
xor U3049 (N_3049,N_1841,N_792);
nor U3050 (N_3050,N_824,N_58);
nor U3051 (N_3051,N_2916,N_2024);
or U3052 (N_3052,N_2860,N_1724);
nor U3053 (N_3053,N_2848,N_266);
or U3054 (N_3054,N_2978,N_664);
and U3055 (N_3055,N_1776,N_2255);
or U3056 (N_3056,N_1719,N_2987);
nor U3057 (N_3057,N_1644,N_2761);
and U3058 (N_3058,N_31,N_2766);
or U3059 (N_3059,N_441,N_109);
nor U3060 (N_3060,N_2912,N_2536);
nor U3061 (N_3061,N_663,N_1569);
xnor U3062 (N_3062,N_2777,N_586);
nand U3063 (N_3063,N_72,N_77);
xnor U3064 (N_3064,N_706,N_1096);
nor U3065 (N_3065,N_2844,N_2698);
nand U3066 (N_3066,N_536,N_457);
nand U3067 (N_3067,N_157,N_161);
or U3068 (N_3068,N_1159,N_1939);
and U3069 (N_3069,N_2956,N_2454);
and U3070 (N_3070,N_897,N_2304);
nand U3071 (N_3071,N_1586,N_2988);
nor U3072 (N_3072,N_2661,N_301);
or U3073 (N_3073,N_1991,N_788);
and U3074 (N_3074,N_406,N_1857);
xor U3075 (N_3075,N_2066,N_761);
xnor U3076 (N_3076,N_1374,N_1121);
and U3077 (N_3077,N_1777,N_1610);
or U3078 (N_3078,N_36,N_1276);
xnor U3079 (N_3079,N_2270,N_338);
nand U3080 (N_3080,N_2347,N_1497);
or U3081 (N_3081,N_181,N_2643);
nor U3082 (N_3082,N_1456,N_2829);
nor U3083 (N_3083,N_2940,N_100);
nor U3084 (N_3084,N_1426,N_2256);
xor U3085 (N_3085,N_2962,N_297);
xnor U3086 (N_3086,N_342,N_231);
xnor U3087 (N_3087,N_1530,N_1532);
and U3088 (N_3088,N_966,N_2434);
nand U3089 (N_3089,N_1962,N_1186);
nor U3090 (N_3090,N_1556,N_1546);
nand U3091 (N_3091,N_2764,N_1486);
nand U3092 (N_3092,N_1513,N_1050);
nand U3093 (N_3093,N_1507,N_1028);
or U3094 (N_3094,N_1411,N_293);
nand U3095 (N_3095,N_1791,N_1592);
and U3096 (N_3096,N_2461,N_2433);
nand U3097 (N_3097,N_1959,N_2498);
nand U3098 (N_3098,N_932,N_1372);
and U3099 (N_3099,N_873,N_1360);
xnor U3100 (N_3100,N_2647,N_2283);
nor U3101 (N_3101,N_737,N_271);
xnor U3102 (N_3102,N_2176,N_1927);
or U3103 (N_3103,N_1252,N_2107);
nand U3104 (N_3104,N_922,N_316);
and U3105 (N_3105,N_1044,N_131);
and U3106 (N_3106,N_1358,N_794);
nand U3107 (N_3107,N_2279,N_1492);
nand U3108 (N_3108,N_2343,N_505);
or U3109 (N_3109,N_813,N_1725);
or U3110 (N_3110,N_2148,N_2265);
and U3111 (N_3111,N_1163,N_2991);
nand U3112 (N_3112,N_436,N_1740);
xnor U3113 (N_3113,N_1578,N_2648);
nand U3114 (N_3114,N_485,N_1410);
or U3115 (N_3115,N_2384,N_1230);
or U3116 (N_3116,N_2150,N_699);
or U3117 (N_3117,N_2364,N_1713);
and U3118 (N_3118,N_1321,N_999);
xnor U3119 (N_3119,N_492,N_1161);
nand U3120 (N_3120,N_1314,N_1908);
and U3121 (N_3121,N_1455,N_1614);
xnor U3122 (N_3122,N_1836,N_1889);
or U3123 (N_3123,N_1750,N_628);
nor U3124 (N_3124,N_2017,N_479);
or U3125 (N_3125,N_2635,N_2064);
nand U3126 (N_3126,N_1559,N_1169);
xor U3127 (N_3127,N_1481,N_731);
xor U3128 (N_3128,N_387,N_1554);
and U3129 (N_3129,N_2409,N_2506);
xor U3130 (N_3130,N_1451,N_462);
nor U3131 (N_3131,N_599,N_2052);
nor U3132 (N_3132,N_2793,N_1417);
and U3133 (N_3133,N_2146,N_2241);
and U3134 (N_3134,N_2873,N_2533);
nand U3135 (N_3135,N_793,N_1662);
nor U3136 (N_3136,N_170,N_647);
or U3137 (N_3137,N_448,N_1926);
nor U3138 (N_3138,N_153,N_952);
nor U3139 (N_3139,N_2640,N_1132);
nand U3140 (N_3140,N_574,N_908);
xor U3141 (N_3141,N_629,N_20);
or U3142 (N_3142,N_2687,N_1903);
or U3143 (N_3143,N_1764,N_1771);
nor U3144 (N_3144,N_2926,N_870);
nand U3145 (N_3145,N_1412,N_2869);
and U3146 (N_3146,N_2208,N_2485);
nor U3147 (N_3147,N_984,N_1907);
xor U3148 (N_3148,N_209,N_790);
nor U3149 (N_3149,N_641,N_2654);
or U3150 (N_3150,N_1123,N_917);
nor U3151 (N_3151,N_214,N_1683);
xor U3152 (N_3152,N_2076,N_503);
or U3153 (N_3153,N_2920,N_885);
and U3154 (N_3154,N_1058,N_225);
and U3155 (N_3155,N_2380,N_259);
and U3156 (N_3156,N_847,N_1313);
nor U3157 (N_3157,N_2630,N_2469);
or U3158 (N_3158,N_2273,N_995);
xnor U3159 (N_3159,N_686,N_247);
or U3160 (N_3160,N_341,N_2866);
xnor U3161 (N_3161,N_958,N_1248);
xnor U3162 (N_3162,N_540,N_1236);
or U3163 (N_3163,N_1944,N_2980);
nand U3164 (N_3164,N_605,N_2048);
xnor U3165 (N_3165,N_1352,N_778);
or U3166 (N_3166,N_973,N_1381);
and U3167 (N_3167,N_1278,N_2377);
or U3168 (N_3168,N_1607,N_1029);
and U3169 (N_3169,N_1422,N_769);
nand U3170 (N_3170,N_2642,N_2449);
xor U3171 (N_3171,N_420,N_2111);
or U3172 (N_3172,N_2072,N_1665);
or U3173 (N_3173,N_2412,N_2252);
nand U3174 (N_3174,N_2922,N_1053);
or U3175 (N_3175,N_1880,N_782);
and U3176 (N_3176,N_1746,N_2705);
nand U3177 (N_3177,N_273,N_2303);
nor U3178 (N_3178,N_2727,N_235);
xor U3179 (N_3179,N_791,N_2877);
and U3180 (N_3180,N_1968,N_1883);
nand U3181 (N_3181,N_1967,N_57);
and U3182 (N_3182,N_1344,N_545);
nor U3183 (N_3183,N_911,N_2113);
nor U3184 (N_3184,N_1258,N_1183);
nor U3185 (N_3185,N_1453,N_718);
or U3186 (N_3186,N_1149,N_1871);
nor U3187 (N_3187,N_139,N_230);
and U3188 (N_3188,N_73,N_2801);
or U3189 (N_3189,N_287,N_352);
xor U3190 (N_3190,N_666,N_91);
xor U3191 (N_3191,N_893,N_413);
and U3192 (N_3192,N_395,N_290);
xor U3193 (N_3193,N_1717,N_2802);
and U3194 (N_3194,N_5,N_719);
nor U3195 (N_3195,N_1400,N_747);
nand U3196 (N_3196,N_2701,N_2058);
and U3197 (N_3197,N_192,N_696);
xnor U3198 (N_3198,N_1404,N_2979);
xnor U3199 (N_3199,N_2893,N_900);
xnor U3200 (N_3200,N_488,N_2995);
nor U3201 (N_3201,N_953,N_429);
or U3202 (N_3202,N_2846,N_590);
and U3203 (N_3203,N_1265,N_1171);
and U3204 (N_3204,N_1565,N_432);
nand U3205 (N_3205,N_2693,N_1917);
xor U3206 (N_3206,N_1282,N_375);
nor U3207 (N_3207,N_1484,N_2889);
nor U3208 (N_3208,N_80,N_621);
and U3209 (N_3209,N_2745,N_2309);
and U3210 (N_3210,N_1340,N_2240);
xor U3211 (N_3211,N_13,N_426);
xor U3212 (N_3212,N_2288,N_2599);
and U3213 (N_3213,N_631,N_840);
nor U3214 (N_3214,N_398,N_360);
or U3215 (N_3215,N_834,N_862);
xnor U3216 (N_3216,N_1605,N_2521);
xnor U3217 (N_3217,N_171,N_2732);
or U3218 (N_3218,N_668,N_2955);
and U3219 (N_3219,N_1524,N_1146);
or U3220 (N_3220,N_2621,N_2892);
nand U3221 (N_3221,N_1388,N_519);
nand U3222 (N_3222,N_2823,N_2441);
and U3223 (N_3223,N_1037,N_2612);
nor U3224 (N_3224,N_1778,N_159);
and U3225 (N_3225,N_2411,N_2410);
or U3226 (N_3226,N_1452,N_2733);
and U3227 (N_3227,N_2425,N_1443);
and U3228 (N_3228,N_2838,N_1158);
xnor U3229 (N_3229,N_2898,N_1879);
and U3230 (N_3230,N_1415,N_1221);
nand U3231 (N_3231,N_1304,N_475);
nand U3232 (N_3232,N_2426,N_2767);
and U3233 (N_3233,N_1487,N_1082);
nor U3234 (N_3234,N_292,N_1744);
xnor U3235 (N_3235,N_1743,N_1870);
and U3236 (N_3236,N_2708,N_1861);
or U3237 (N_3237,N_2937,N_1721);
nand U3238 (N_3238,N_1198,N_709);
nor U3239 (N_3239,N_1273,N_1268);
xor U3240 (N_3240,N_822,N_349);
nor U3241 (N_3241,N_1639,N_30);
or U3242 (N_3242,N_2952,N_2178);
nor U3243 (N_3243,N_638,N_2000);
nor U3244 (N_3244,N_2077,N_976);
nor U3245 (N_3245,N_120,N_374);
xor U3246 (N_3246,N_2378,N_2567);
xnor U3247 (N_3247,N_1303,N_526);
or U3248 (N_3248,N_2297,N_2110);
and U3249 (N_3249,N_2397,N_2826);
nor U3250 (N_3250,N_2785,N_2915);
nor U3251 (N_3251,N_299,N_2639);
and U3252 (N_3252,N_2637,N_289);
nand U3253 (N_3253,N_997,N_2651);
and U3254 (N_3254,N_204,N_1250);
xor U3255 (N_3255,N_2211,N_2133);
or U3256 (N_3256,N_2957,N_2774);
nand U3257 (N_3257,N_502,N_2120);
nor U3258 (N_3258,N_2261,N_1017);
or U3259 (N_3259,N_1667,N_1659);
nand U3260 (N_3260,N_783,N_2814);
xor U3261 (N_3261,N_927,N_625);
or U3262 (N_3262,N_2228,N_1444);
and U3263 (N_3263,N_1947,N_1025);
or U3264 (N_3264,N_948,N_2725);
or U3265 (N_3265,N_1450,N_2868);
or U3266 (N_3266,N_1018,N_1829);
and U3267 (N_3267,N_918,N_562);
nor U3268 (N_3268,N_370,N_1038);
nor U3269 (N_3269,N_45,N_2039);
xor U3270 (N_3270,N_2544,N_2570);
nand U3271 (N_3271,N_929,N_2750);
and U3272 (N_3272,N_2959,N_359);
nor U3273 (N_3273,N_1104,N_1978);
xnor U3274 (N_3274,N_2582,N_424);
nand U3275 (N_3275,N_1189,N_1601);
or U3276 (N_3276,N_1970,N_1020);
and U3277 (N_3277,N_566,N_2328);
xnor U3278 (N_3278,N_2719,N_2470);
nor U3279 (N_3279,N_2205,N_317);
nor U3280 (N_3280,N_2216,N_2247);
or U3281 (N_3281,N_2341,N_1157);
and U3282 (N_3282,N_1325,N_184);
nand U3283 (N_3283,N_1876,N_1235);
nor U3284 (N_3284,N_2529,N_487);
or U3285 (N_3285,N_2466,N_2147);
or U3286 (N_3286,N_1828,N_1603);
and U3287 (N_3287,N_2497,N_307);
xor U3288 (N_3288,N_372,N_1107);
and U3289 (N_3289,N_844,N_2910);
xnor U3290 (N_3290,N_1260,N_2234);
nor U3291 (N_3291,N_210,N_1723);
xnor U3292 (N_3292,N_336,N_2589);
nand U3293 (N_3293,N_2872,N_51);
xnor U3294 (N_3294,N_2320,N_1473);
xor U3295 (N_3295,N_2153,N_2723);
or U3296 (N_3296,N_882,N_1001);
or U3297 (N_3297,N_1211,N_854);
xor U3298 (N_3298,N_2562,N_1005);
or U3299 (N_3299,N_1172,N_1884);
xor U3300 (N_3300,N_1999,N_584);
or U3301 (N_3301,N_767,N_2843);
nor U3302 (N_3302,N_591,N_2748);
xnor U3303 (N_3303,N_1330,N_1936);
nand U3304 (N_3304,N_1886,N_2138);
nand U3305 (N_3305,N_187,N_996);
or U3306 (N_3306,N_2201,N_702);
or U3307 (N_3307,N_458,N_875);
xnor U3308 (N_3308,N_2789,N_859);
xor U3309 (N_3309,N_1941,N_1837);
xor U3310 (N_3310,N_333,N_2609);
or U3311 (N_3311,N_2997,N_1434);
or U3312 (N_3312,N_48,N_2728);
nand U3313 (N_3313,N_303,N_2931);
or U3314 (N_3314,N_283,N_814);
nor U3315 (N_3315,N_1653,N_2857);
nand U3316 (N_3316,N_820,N_1350);
or U3317 (N_3317,N_2419,N_2969);
or U3318 (N_3318,N_2260,N_2778);
nand U3319 (N_3319,N_1447,N_573);
or U3320 (N_3320,N_2689,N_2665);
nor U3321 (N_3321,N_888,N_1041);
nor U3322 (N_3322,N_1752,N_2597);
nand U3323 (N_3323,N_46,N_1262);
nand U3324 (N_3324,N_579,N_1222);
or U3325 (N_3325,N_2492,N_2462);
nand U3326 (N_3326,N_781,N_750);
nand U3327 (N_3327,N_2682,N_1162);
xor U3328 (N_3328,N_186,N_2853);
xnor U3329 (N_3329,N_228,N_1826);
nor U3330 (N_3330,N_653,N_328);
nand U3331 (N_3331,N_2999,N_1299);
nor U3332 (N_3332,N_2699,N_1858);
and U3333 (N_3333,N_1301,N_154);
nand U3334 (N_3334,N_275,N_142);
xor U3335 (N_3335,N_1580,N_2713);
or U3336 (N_3336,N_786,N_269);
and U3337 (N_3337,N_2439,N_2759);
or U3338 (N_3338,N_2876,N_2269);
or U3339 (N_3339,N_816,N_1094);
or U3340 (N_3340,N_1755,N_2653);
nor U3341 (N_3341,N_635,N_2115);
xor U3342 (N_3342,N_1166,N_1000);
nand U3343 (N_3343,N_945,N_1855);
xor U3344 (N_3344,N_1615,N_2958);
nand U3345 (N_3345,N_2510,N_821);
nor U3346 (N_3346,N_1868,N_1843);
or U3347 (N_3347,N_108,N_464);
nor U3348 (N_3348,N_2557,N_456);
nand U3349 (N_3349,N_648,N_2990);
nor U3350 (N_3350,N_193,N_1973);
or U3351 (N_3351,N_2137,N_1613);
xnor U3352 (N_3352,N_484,N_2007);
nand U3353 (N_3353,N_2266,N_44);
or U3354 (N_3354,N_1401,N_2209);
nor U3355 (N_3355,N_798,N_2734);
xnor U3356 (N_3356,N_601,N_697);
nand U3357 (N_3357,N_988,N_2928);
or U3358 (N_3358,N_1311,N_1496);
and U3359 (N_3359,N_1418,N_2587);
xnor U3360 (N_3360,N_1890,N_514);
nor U3361 (N_3361,N_1164,N_527);
and U3362 (N_3362,N_1462,N_1849);
nor U3363 (N_3363,N_580,N_288);
and U3364 (N_3364,N_1130,N_1328);
nand U3365 (N_3365,N_2029,N_1306);
nor U3366 (N_3366,N_2575,N_2079);
xnor U3367 (N_3367,N_2121,N_2856);
and U3368 (N_3368,N_872,N_1637);
xor U3369 (N_3369,N_832,N_1337);
nor U3370 (N_3370,N_646,N_2743);
and U3371 (N_3371,N_1284,N_974);
nor U3372 (N_3372,N_2951,N_2440);
nor U3373 (N_3373,N_373,N_1366);
or U3374 (N_3374,N_1478,N_2134);
or U3375 (N_3375,N_216,N_419);
nor U3376 (N_3376,N_238,N_1747);
or U3377 (N_3377,N_2967,N_313);
nand U3378 (N_3378,N_2360,N_2601);
nand U3379 (N_3379,N_1253,N_384);
xor U3380 (N_3380,N_695,N_1174);
nand U3381 (N_3381,N_2159,N_1520);
nor U3382 (N_3382,N_2755,N_1329);
xnor U3383 (N_3383,N_86,N_815);
or U3384 (N_3384,N_1924,N_2085);
and U3385 (N_3385,N_2396,N_2923);
or U3386 (N_3386,N_2301,N_2338);
or U3387 (N_3387,N_915,N_2527);
xor U3388 (N_3388,N_943,N_597);
xor U3389 (N_3389,N_2371,N_877);
nand U3390 (N_3390,N_2655,N_1477);
and U3391 (N_3391,N_1711,N_1463);
or U3392 (N_3392,N_1897,N_1553);
and U3393 (N_3393,N_40,N_364);
nor U3394 (N_3394,N_1729,N_1472);
nor U3395 (N_3395,N_1097,N_623);
nor U3396 (N_3396,N_2223,N_1255);
nand U3397 (N_3397,N_1681,N_2638);
and U3398 (N_3398,N_2238,N_2001);
and U3399 (N_3399,N_941,N_1825);
nor U3400 (N_3400,N_2264,N_1690);
or U3401 (N_3401,N_867,N_611);
or U3402 (N_3402,N_1618,N_2365);
and U3403 (N_3403,N_2057,N_1134);
and U3404 (N_3404,N_1502,N_2579);
and U3405 (N_3405,N_1748,N_765);
and U3406 (N_3406,N_2395,N_2129);
nor U3407 (N_3407,N_2156,N_807);
xor U3408 (N_3408,N_2489,N_809);
xor U3409 (N_3409,N_2592,N_970);
nor U3410 (N_3410,N_1234,N_763);
nor U3411 (N_3411,N_2030,N_1617);
and U3412 (N_3412,N_1628,N_1840);
nor U3413 (N_3413,N_2961,N_724);
or U3414 (N_3414,N_1034,N_1223);
xnor U3415 (N_3415,N_2796,N_1878);
nor U3416 (N_3416,N_476,N_2839);
xnor U3417 (N_3417,N_365,N_39);
or U3418 (N_3418,N_2359,N_1124);
and U3419 (N_3419,N_1790,N_11);
or U3420 (N_3420,N_2941,N_662);
or U3421 (N_3421,N_2971,N_222);
xor U3422 (N_3422,N_430,N_808);
nand U3423 (N_3423,N_2016,N_2722);
xnor U3424 (N_3424,N_2248,N_1591);
or U3425 (N_3425,N_1943,N_926);
and U3426 (N_3426,N_366,N_177);
or U3427 (N_3427,N_2037,N_1465);
nor U3428 (N_3428,N_951,N_2455);
nor U3429 (N_3429,N_2692,N_2082);
or U3430 (N_3430,N_1259,N_1458);
or U3431 (N_3431,N_609,N_0);
and U3432 (N_3432,N_797,N_136);
or U3433 (N_3433,N_2206,N_1431);
nand U3434 (N_3434,N_1669,N_2634);
nor U3435 (N_3435,N_1518,N_2964);
and U3436 (N_3436,N_963,N_1510);
and U3437 (N_3437,N_1851,N_2763);
nor U3438 (N_3438,N_2381,N_1092);
xnor U3439 (N_3439,N_2136,N_524);
and U3440 (N_3440,N_2667,N_1047);
or U3441 (N_3441,N_946,N_380);
xor U3442 (N_3442,N_2093,N_811);
and U3443 (N_3443,N_1049,N_1864);
nand U3444 (N_3444,N_1346,N_2986);
or U3445 (N_3445,N_2773,N_2909);
nor U3446 (N_3446,N_1244,N_2392);
xnor U3447 (N_3447,N_1676,N_2404);
or U3448 (N_3448,N_2513,N_323);
nand U3449 (N_3449,N_2098,N_169);
or U3450 (N_3450,N_2388,N_787);
nand U3451 (N_3451,N_2004,N_1127);
nand U3452 (N_3452,N_21,N_1229);
xnor U3453 (N_3453,N_2891,N_2935);
or U3454 (N_3454,N_1227,N_2859);
xor U3455 (N_3455,N_1904,N_2691);
nand U3456 (N_3456,N_1900,N_2549);
nand U3457 (N_3457,N_557,N_2018);
xor U3458 (N_3458,N_331,N_452);
xor U3459 (N_3459,N_1220,N_67);
nand U3460 (N_3460,N_425,N_2083);
nand U3461 (N_3461,N_2177,N_449);
nand U3462 (N_3462,N_1081,N_1293);
or U3463 (N_3463,N_296,N_418);
nor U3464 (N_3464,N_227,N_1606);
nor U3465 (N_3465,N_402,N_1948);
nor U3466 (N_3466,N_1738,N_1657);
and U3467 (N_3467,N_229,N_2363);
xnor U3468 (N_3468,N_508,N_1031);
nand U3469 (N_3469,N_1048,N_2191);
and U3470 (N_3470,N_2189,N_710);
xor U3471 (N_3471,N_1706,N_853);
and U3472 (N_3472,N_515,N_693);
and U3473 (N_3473,N_509,N_1439);
nor U3474 (N_3474,N_1865,N_890);
and U3475 (N_3475,N_1859,N_346);
nor U3476 (N_3476,N_2351,N_340);
and U3477 (N_3477,N_1254,N_1297);
nand U3478 (N_3478,N_1735,N_401);
nand U3479 (N_3479,N_2162,N_2812);
nand U3480 (N_3480,N_2685,N_930);
and U3481 (N_3481,N_764,N_1818);
nand U3482 (N_3482,N_1375,N_1188);
or U3483 (N_3483,N_1228,N_2031);
nand U3484 (N_3484,N_2942,N_127);
nor U3485 (N_3485,N_2550,N_546);
xor U3486 (N_3486,N_1789,N_55);
and U3487 (N_3487,N_2827,N_2379);
or U3488 (N_3488,N_2501,N_2580);
nand U3489 (N_3489,N_2342,N_1363);
nor U3490 (N_3490,N_1291,N_2711);
nand U3491 (N_3491,N_2901,N_144);
nor U3492 (N_3492,N_1869,N_431);
nand U3493 (N_3493,N_175,N_2011);
nand U3494 (N_3494,N_726,N_196);
nor U3495 (N_3495,N_382,N_1416);
nor U3496 (N_3496,N_1208,N_1195);
nor U3497 (N_3497,N_1645,N_85);
nand U3498 (N_3498,N_898,N_1193);
and U3499 (N_3499,N_749,N_347);
and U3500 (N_3500,N_2886,N_179);
xnor U3501 (N_3501,N_405,N_1517);
and U3502 (N_3502,N_490,N_1905);
and U3503 (N_3503,N_1799,N_2929);
xnor U3504 (N_3504,N_2628,N_1702);
xor U3505 (N_3505,N_463,N_1533);
xor U3506 (N_3506,N_1490,N_935);
xor U3507 (N_3507,N_2538,N_884);
xnor U3508 (N_3508,N_602,N_2278);
xnor U3509 (N_3509,N_1994,N_758);
and U3510 (N_3510,N_442,N_1584);
or U3511 (N_3511,N_2577,N_1787);
nand U3512 (N_3512,N_285,N_1457);
xnor U3513 (N_3513,N_2027,N_1577);
xor U3514 (N_3514,N_692,N_2374);
or U3515 (N_3515,N_1102,N_2245);
or U3516 (N_3516,N_2707,N_2576);
and U3517 (N_3517,N_2399,N_1112);
nand U3518 (N_3518,N_1289,N_2581);
and U3519 (N_3519,N_1379,N_1300);
nor U3520 (N_3520,N_1167,N_2075);
or U3521 (N_3521,N_149,N_1562);
xnor U3522 (N_3522,N_2906,N_1898);
or U3523 (N_3523,N_801,N_1547);
nor U3524 (N_3524,N_1633,N_2348);
and U3525 (N_3525,N_651,N_561);
xor U3526 (N_3526,N_134,N_2322);
and U3527 (N_3527,N_685,N_1989);
and U3528 (N_3528,N_2982,N_2946);
or U3529 (N_3529,N_746,N_239);
nor U3530 (N_3530,N_2476,N_391);
xor U3531 (N_3531,N_1277,N_459);
xor U3532 (N_3532,N_2175,N_2834);
xnor U3533 (N_3533,N_468,N_1945);
nor U3534 (N_3534,N_658,N_1338);
nor U3535 (N_3535,N_2571,N_649);
or U3536 (N_3536,N_679,N_2420);
nand U3537 (N_3537,N_477,N_1148);
nor U3538 (N_3538,N_2073,N_2067);
xnor U3539 (N_3539,N_881,N_26);
or U3540 (N_3540,N_8,N_274);
or U3541 (N_3541,N_1501,N_1213);
and U3542 (N_3542,N_1995,N_1763);
or U3543 (N_3543,N_1537,N_2171);
nor U3544 (N_3544,N_857,N_404);
and U3545 (N_3545,N_440,N_2593);
nor U3546 (N_3546,N_1640,N_886);
xor U3547 (N_3547,N_1024,N_525);
and U3548 (N_3548,N_708,N_2895);
nor U3549 (N_3549,N_1882,N_99);
nor U3550 (N_3550,N_803,N_1283);
and U3551 (N_3551,N_2788,N_1568);
and U3552 (N_3552,N_1448,N_2532);
or U3553 (N_3553,N_2284,N_451);
or U3554 (N_3554,N_2798,N_1611);
or U3555 (N_3555,N_1084,N_818);
xnor U3556 (N_3556,N_258,N_2094);
nor U3557 (N_3557,N_956,N_1602);
nand U3558 (N_3558,N_107,N_1680);
nor U3559 (N_3559,N_353,N_115);
or U3560 (N_3560,N_1971,N_2262);
xor U3561 (N_3561,N_332,N_215);
or U3562 (N_3562,N_1656,N_1712);
nand U3563 (N_3563,N_59,N_1575);
nor U3564 (N_3564,N_2717,N_1641);
xnor U3565 (N_3565,N_774,N_326);
xor U3566 (N_3566,N_1914,N_2421);
nand U3567 (N_3567,N_2046,N_2563);
xnor U3568 (N_3568,N_90,N_2035);
nand U3569 (N_3569,N_523,N_2180);
and U3570 (N_3570,N_1582,N_377);
and U3571 (N_3571,N_2765,N_1548);
and U3572 (N_3572,N_1022,N_252);
nand U3573 (N_3573,N_1332,N_1736);
or U3574 (N_3574,N_1428,N_1563);
nand U3575 (N_3575,N_1932,N_1915);
or U3576 (N_3576,N_2286,N_62);
or U3577 (N_3577,N_1780,N_446);
nor U3578 (N_3578,N_863,N_1011);
or U3579 (N_3579,N_1241,N_1946);
and U3580 (N_3580,N_1296,N_2145);
nand U3581 (N_3581,N_1931,N_626);
nor U3582 (N_3582,N_838,N_858);
nand U3583 (N_3583,N_233,N_2314);
and U3584 (N_3584,N_2307,N_439);
and U3585 (N_3585,N_1585,N_1626);
nand U3586 (N_3586,N_199,N_2787);
or U3587 (N_3587,N_964,N_433);
xnor U3588 (N_3588,N_990,N_738);
nor U3589 (N_3589,N_1197,N_114);
nor U3590 (N_3590,N_2407,N_2135);
xnor U3591 (N_3591,N_1010,N_2084);
nor U3592 (N_3592,N_49,N_369);
or U3593 (N_3593,N_1694,N_2158);
nor U3594 (N_3594,N_2070,N_1696);
or U3595 (N_3595,N_248,N_2989);
nor U3596 (N_3596,N_656,N_2611);
xor U3597 (N_3597,N_1437,N_2032);
nor U3598 (N_3598,N_2369,N_1212);
and U3599 (N_3599,N_2251,N_2970);
nand U3600 (N_3600,N_2981,N_2097);
or U3601 (N_3601,N_435,N_1187);
or U3602 (N_3602,N_1312,N_914);
and U3603 (N_3603,N_549,N_2747);
xnor U3604 (N_3604,N_2636,N_2966);
and U3605 (N_3605,N_2933,N_1089);
and U3606 (N_3606,N_2566,N_1466);
nand U3607 (N_3607,N_1891,N_936);
nand U3608 (N_3608,N_2810,N_2002);
and U3609 (N_3609,N_2361,N_1922);
nand U3610 (N_3610,N_1182,N_1803);
xor U3611 (N_3611,N_1521,N_571);
xnor U3612 (N_3612,N_2294,N_1673);
nor U3613 (N_3613,N_396,N_1015);
xnor U3614 (N_3614,N_2089,N_2675);
nor U3615 (N_3615,N_63,N_1459);
nor U3616 (N_3616,N_1820,N_2925);
xnor U3617 (N_3617,N_2108,N_1976);
and U3618 (N_3618,N_1270,N_1961);
or U3619 (N_3619,N_400,N_2398);
nand U3620 (N_3620,N_987,N_640);
nor U3621 (N_3621,N_2215,N_2296);
or U3622 (N_3622,N_306,N_1650);
or U3623 (N_3623,N_2806,N_129);
nand U3624 (N_3624,N_224,N_1608);
nand U3625 (N_3625,N_2973,N_2290);
nand U3626 (N_3626,N_1823,N_825);
xnor U3627 (N_3627,N_2233,N_1339);
nor U3628 (N_3628,N_606,N_219);
or U3629 (N_3629,N_280,N_2505);
nand U3630 (N_3630,N_344,N_1072);
and U3631 (N_3631,N_2974,N_1063);
or U3632 (N_3632,N_389,N_2662);
or U3633 (N_3633,N_1589,N_111);
and U3634 (N_3634,N_711,N_2169);
xor U3635 (N_3635,N_851,N_2867);
nor U3636 (N_3636,N_2519,N_2344);
xor U3637 (N_3637,N_2026,N_1753);
nand U3638 (N_3638,N_1509,N_734);
nand U3639 (N_3639,N_1739,N_1177);
or U3640 (N_3640,N_772,N_501);
nor U3641 (N_3641,N_661,N_2854);
xor U3642 (N_3642,N_2816,N_2190);
nand U3643 (N_3643,N_320,N_2317);
and U3644 (N_3644,N_2494,N_1414);
nand U3645 (N_3645,N_1847,N_1635);
or U3646 (N_3646,N_2845,N_3);
and U3647 (N_3647,N_1689,N_379);
and U3648 (N_3648,N_1489,N_957);
nor U3649 (N_3649,N_2850,N_1769);
nor U3650 (N_3650,N_539,N_2871);
nor U3651 (N_3651,N_1485,N_1986);
xnor U3652 (N_3652,N_2760,N_2038);
xnor U3653 (N_3653,N_2312,N_887);
nor U3654 (N_3654,N_104,N_2656);
xor U3655 (N_3655,N_1827,N_1506);
xor U3656 (N_3656,N_71,N_2424);
xor U3657 (N_3657,N_1245,N_2907);
or U3658 (N_3658,N_1955,N_1257);
and U3659 (N_3659,N_1376,N_2797);
nand U3660 (N_3660,N_1660,N_768);
or U3661 (N_3661,N_1974,N_1792);
nand U3662 (N_3662,N_455,N_1389);
or U3663 (N_3663,N_1016,N_250);
and U3664 (N_3664,N_2219,N_1596);
nor U3665 (N_3665,N_2694,N_2818);
or U3666 (N_3666,N_717,N_613);
nand U3667 (N_3667,N_2835,N_493);
nand U3668 (N_3668,N_1263,N_103);
or U3669 (N_3669,N_2194,N_560);
xnor U3670 (N_3670,N_2451,N_2585);
xnor U3671 (N_3671,N_2152,N_1077);
xnor U3672 (N_3672,N_2697,N_2402);
nor U3673 (N_3673,N_622,N_156);
and U3674 (N_3674,N_1632,N_1009);
nor U3675 (N_3675,N_291,N_771);
or U3676 (N_3676,N_198,N_1116);
xor U3677 (N_3677,N_2674,N_2700);
nand U3678 (N_3678,N_2275,N_1362);
xnor U3679 (N_3679,N_1137,N_1623);
xnor U3680 (N_3680,N_587,N_1579);
nor U3681 (N_3681,N_2913,N_1206);
and U3682 (N_3682,N_2021,N_1785);
and U3683 (N_3683,N_2684,N_2619);
nand U3684 (N_3684,N_1921,N_985);
nor U3685 (N_3685,N_2531,N_2828);
nand U3686 (N_3686,N_1734,N_645);
xor U3687 (N_3687,N_1409,N_1983);
nor U3688 (N_3688,N_217,N_1120);
nor U3689 (N_3689,N_1796,N_1549);
or U3690 (N_3690,N_1664,N_1745);
or U3691 (N_3691,N_1622,N_1292);
and U3692 (N_3692,N_1536,N_678);
and U3693 (N_3693,N_1742,N_855);
nor U3694 (N_3694,N_140,N_1901);
or U3695 (N_3695,N_902,N_833);
or U3696 (N_3696,N_1320,N_2977);
xnor U3697 (N_3697,N_2883,N_2013);
nand U3698 (N_3698,N_1209,N_2272);
or U3699 (N_3699,N_2358,N_279);
and U3700 (N_3700,N_2349,N_1138);
and U3701 (N_3701,N_1119,N_1805);
nand U3702 (N_3702,N_2334,N_1527);
xor U3703 (N_3703,N_2258,N_1555);
nand U3704 (N_3704,N_472,N_83);
nand U3705 (N_3705,N_2659,N_981);
nor U3706 (N_3706,N_173,N_2131);
or U3707 (N_3707,N_680,N_819);
and U3708 (N_3708,N_700,N_704);
nor U3709 (N_3709,N_652,N_251);
nor U3710 (N_3710,N_32,N_2340);
nor U3711 (N_3711,N_2230,N_1393);
nor U3712 (N_3712,N_2605,N_2811);
nor U3713 (N_3713,N_2202,N_2218);
nand U3714 (N_3714,N_42,N_2006);
nand U3715 (N_3715,N_1004,N_1954);
nor U3716 (N_3716,N_1526,N_2481);
xor U3717 (N_3717,N_1811,N_2504);
or U3718 (N_3718,N_2588,N_2095);
nand U3719 (N_3719,N_2851,N_1716);
xnor U3720 (N_3720,N_2043,N_2954);
nor U3721 (N_3721,N_2267,N_188);
nand U3722 (N_3722,N_371,N_1140);
or U3723 (N_3723,N_1373,N_1269);
nor U3724 (N_3724,N_2545,N_780);
and U3725 (N_3725,N_1911,N_1468);
xor U3726 (N_3726,N_1906,N_1136);
xor U3727 (N_3727,N_831,N_28);
and U3728 (N_3728,N_2770,N_1588);
nand U3729 (N_3729,N_1110,N_2435);
or U3730 (N_3730,N_618,N_1027);
or U3731 (N_3731,N_2650,N_2472);
nand U3732 (N_3732,N_2063,N_2775);
or U3733 (N_3733,N_1894,N_785);
or U3734 (N_3734,N_940,N_977);
xor U3735 (N_3735,N_2391,N_1666);
nor U3736 (N_3736,N_2373,N_1247);
and U3737 (N_3737,N_1951,N_839);
nand U3738 (N_3738,N_2271,N_762);
nand U3739 (N_3739,N_1272,N_2368);
or U3740 (N_3740,N_281,N_675);
xor U3741 (N_3741,N_756,N_2458);
xor U3742 (N_3742,N_2622,N_2274);
nand U3743 (N_3743,N_1280,N_276);
nor U3744 (N_3744,N_2329,N_409);
and U3745 (N_3745,N_616,N_634);
and U3746 (N_3746,N_52,N_1720);
nor U3747 (N_3747,N_1860,N_1942);
nor U3748 (N_3748,N_1105,N_773);
or U3749 (N_3749,N_1919,N_2905);
and U3750 (N_3750,N_2463,N_1560);
or U3751 (N_3751,N_2166,N_2712);
and U3752 (N_3752,N_256,N_547);
xnor U3753 (N_3753,N_92,N_720);
nor U3754 (N_3754,N_2080,N_1649);
and U3755 (N_3755,N_1392,N_1394);
or U3756 (N_3756,N_1493,N_294);
xnor U3757 (N_3757,N_2416,N_2474);
nand U3758 (N_3758,N_2862,N_1319);
xor U3759 (N_3759,N_33,N_2298);
xnor U3760 (N_3760,N_2151,N_2484);
or U3761 (N_3761,N_1202,N_2025);
and U3762 (N_3762,N_703,N_1505);
or U3763 (N_3763,N_356,N_112);
nor U3764 (N_3764,N_2511,N_2564);
xor U3765 (N_3765,N_683,N_979);
nor U3766 (N_3766,N_2491,N_2695);
or U3767 (N_3767,N_43,N_1570);
xnor U3768 (N_3768,N_23,N_924);
nor U3769 (N_3769,N_1108,N_1423);
nor U3770 (N_3770,N_2282,N_1176);
nand U3771 (N_3771,N_939,N_191);
xor U3772 (N_3772,N_1026,N_2277);
xnor U3773 (N_3773,N_1364,N_1774);
nor U3774 (N_3774,N_2594,N_670);
nand U3775 (N_3775,N_2060,N_278);
nor U3776 (N_3776,N_1080,N_117);
xnor U3777 (N_3777,N_2584,N_2880);
nor U3778 (N_3778,N_2528,N_553);
xor U3779 (N_3779,N_2413,N_1807);
or U3780 (N_3780,N_849,N_2771);
nand U3781 (N_3781,N_1117,N_2754);
or U3782 (N_3782,N_2450,N_2417);
nor U3783 (N_3783,N_1950,N_1677);
nor U3784 (N_3784,N_1875,N_2633);
xnor U3785 (N_3785,N_2401,N_1838);
nand U3786 (N_3786,N_1793,N_1698);
and U3787 (N_3787,N_752,N_2948);
nor U3788 (N_3788,N_1705,N_1599);
nor U3789 (N_3789,N_1581,N_1854);
or U3790 (N_3790,N_2704,N_604);
xor U3791 (N_3791,N_1678,N_1190);
xor U3792 (N_3792,N_1368,N_894);
nand U3793 (N_3793,N_1979,N_544);
and U3794 (N_3794,N_311,N_659);
xor U3795 (N_3795,N_2263,N_1175);
nand U3796 (N_3796,N_2112,N_2480);
xnor U3797 (N_3797,N_1113,N_106);
nand U3798 (N_3798,N_1531,N_2142);
nor U3799 (N_3799,N_934,N_118);
nor U3800 (N_3800,N_329,N_2221);
nand U3801 (N_3801,N_2244,N_2354);
nor U3802 (N_3802,N_1515,N_416);
or U3803 (N_3803,N_1651,N_138);
nand U3804 (N_3804,N_707,N_2617);
nand U3805 (N_3805,N_18,N_1564);
nor U3806 (N_3806,N_569,N_1087);
and U3807 (N_3807,N_2608,N_1893);
or U3808 (N_3808,N_2690,N_1043);
or U3809 (N_3809,N_2830,N_2832);
xnor U3810 (N_3810,N_116,N_1464);
and U3811 (N_3811,N_469,N_367);
or U3812 (N_3812,N_1060,N_1361);
and U3813 (N_3813,N_2173,N_1726);
xnor U3814 (N_3814,N_1207,N_2237);
xnor U3815 (N_3815,N_211,N_2346);
nor U3816 (N_3816,N_2858,N_1815);
nand U3817 (N_3817,N_2114,N_2899);
and U3818 (N_3818,N_928,N_2718);
nand U3819 (N_3819,N_17,N_1033);
xnor U3820 (N_3820,N_1775,N_1139);
nor U3821 (N_3821,N_612,N_980);
and U3822 (N_3822,N_208,N_2610);
nand U3823 (N_3823,N_2447,N_438);
or U3824 (N_3824,N_2005,N_1056);
and U3825 (N_3825,N_1305,N_2306);
nand U3826 (N_3826,N_1850,N_2672);
and U3827 (N_3827,N_2090,N_1757);
and U3828 (N_3828,N_1359,N_480);
nor U3829 (N_3829,N_1294,N_2311);
and U3830 (N_3830,N_592,N_190);
xor U3831 (N_3831,N_723,N_1324);
nor U3832 (N_3832,N_70,N_1151);
or U3833 (N_3833,N_1594,N_2197);
nor U3834 (N_3834,N_982,N_1103);
and U3835 (N_3835,N_810,N_1624);
xor U3836 (N_3836,N_856,N_1885);
xnor U3837 (N_3837,N_1156,N_828);
and U3838 (N_3838,N_1251,N_499);
or U3839 (N_3839,N_823,N_264);
nand U3840 (N_3840,N_516,N_2677);
nand U3841 (N_3841,N_2556,N_327);
nand U3842 (N_3842,N_1795,N_1476);
xor U3843 (N_3843,N_555,N_1511);
nor U3844 (N_3844,N_2714,N_2149);
and U3845 (N_3845,N_1956,N_1500);
nor U3846 (N_3846,N_254,N_2780);
xnor U3847 (N_3847,N_2976,N_2894);
nand U3848 (N_3848,N_868,N_1371);
xor U3849 (N_3849,N_619,N_1281);
nand U3850 (N_3850,N_2172,N_1647);
and U3851 (N_3851,N_2473,N_2356);
nor U3852 (N_3852,N_2953,N_1288);
xor U3853 (N_3853,N_125,N_2124);
nor U3854 (N_3854,N_121,N_357);
nor U3855 (N_3855,N_757,N_2716);
and U3856 (N_3856,N_2350,N_1298);
xor U3857 (N_3857,N_305,N_1470);
xor U3858 (N_3858,N_1934,N_2488);
nor U3859 (N_3859,N_1413,N_1981);
nand U3860 (N_3860,N_2362,N_1225);
or U3861 (N_3861,N_1406,N_1895);
nand U3862 (N_3862,N_1365,N_2543);
and U3863 (N_3863,N_920,N_2482);
nor U3864 (N_3864,N_2836,N_1544);
xnor U3865 (N_3865,N_2516,N_2551);
or U3866 (N_3866,N_1512,N_671);
xor U3867 (N_3867,N_1488,N_1714);
or U3868 (N_3868,N_1965,N_2448);
xnor U3869 (N_3869,N_1194,N_221);
or U3870 (N_3870,N_399,N_2772);
nor U3871 (N_3871,N_302,N_309);
nand U3872 (N_3872,N_2464,N_1913);
and U3873 (N_3873,N_603,N_1842);
or U3874 (N_3874,N_312,N_923);
nor U3875 (N_3875,N_1144,N_722);
xnor U3876 (N_3876,N_2993,N_65);
and U3877 (N_3877,N_350,N_361);
and U3878 (N_3878,N_145,N_537);
and U3879 (N_3879,N_842,N_1179);
xnor U3880 (N_3880,N_245,N_1661);
nand U3881 (N_3881,N_1810,N_2681);
xor U3882 (N_3882,N_989,N_620);
and U3883 (N_3883,N_681,N_860);
xnor U3884 (N_3884,N_1892,N_730);
nand U3885 (N_3885,N_2293,N_1732);
nor U3886 (N_3886,N_2471,N_2792);
nand U3887 (N_3887,N_1937,N_2613);
nor U3888 (N_3888,N_201,N_2749);
or U3889 (N_3889,N_2614,N_994);
nor U3890 (N_3890,N_1751,N_2243);
nor U3891 (N_3891,N_1285,N_2897);
nand U3892 (N_3892,N_2680,N_522);
xnor U3893 (N_3893,N_1844,N_1923);
and U3894 (N_3894,N_202,N_260);
xor U3895 (N_3895,N_2864,N_913);
xnor U3896 (N_3896,N_304,N_220);
nand U3897 (N_3897,N_68,N_1440);
and U3898 (N_3898,N_358,N_1178);
nand U3899 (N_3899,N_965,N_655);
nand U3900 (N_3900,N_2808,N_1261);
or U3901 (N_3901,N_2703,N_147);
nand U3902 (N_3902,N_991,N_348);
and U3903 (N_3903,N_60,N_1754);
or U3904 (N_3904,N_1435,N_2524);
nand U3905 (N_3905,N_410,N_253);
or U3906 (N_3906,N_1710,N_15);
nor U3907 (N_3907,N_1972,N_2071);
and U3908 (N_3908,N_1993,N_1066);
nand U3909 (N_3909,N_596,N_1032);
nand U3910 (N_3910,N_1012,N_2357);
xnor U3911 (N_3911,N_2824,N_2984);
or U3912 (N_3912,N_595,N_2752);
nor U3913 (N_3913,N_1483,N_50);
nand U3914 (N_3914,N_2526,N_2059);
nand U3915 (N_3915,N_826,N_2744);
xor U3916 (N_3916,N_113,N_2220);
and U3917 (N_3917,N_2720,N_2214);
nand U3918 (N_3918,N_2132,N_1929);
xor U3919 (N_3919,N_1953,N_1099);
xnor U3920 (N_3920,N_912,N_1808);
or U3921 (N_3921,N_2106,N_895);
and U3922 (N_3922,N_1881,N_2737);
nand U3923 (N_3923,N_1133,N_755);
and U3924 (N_3924,N_1975,N_130);
nor U3925 (N_3925,N_1318,N_2963);
and U3926 (N_3926,N_1987,N_921);
xor U3927 (N_3927,N_2586,N_2903);
nand U3928 (N_3928,N_343,N_1129);
nor U3929 (N_3929,N_575,N_2254);
or U3930 (N_3930,N_237,N_2768);
and U3931 (N_3931,N_2250,N_2805);
and U3932 (N_3932,N_950,N_1152);
nor U3933 (N_3933,N_189,N_1181);
nand U3934 (N_3934,N_879,N_411);
or U3935 (N_3935,N_2507,N_471);
xnor U3936 (N_3936,N_2739,N_1809);
xnor U3937 (N_3937,N_548,N_324);
nor U3938 (N_3938,N_1240,N_1006);
and U3939 (N_3939,N_1046,N_986);
nand U3940 (N_3940,N_421,N_1091);
xor U3941 (N_3941,N_2616,N_1687);
xnor U3942 (N_3942,N_830,N_2683);
xnor U3943 (N_3943,N_843,N_2795);
or U3944 (N_3944,N_1051,N_2257);
or U3945 (N_3945,N_1191,N_1749);
or U3946 (N_3946,N_2144,N_185);
nand U3947 (N_3947,N_1385,N_2606);
nor U3948 (N_3948,N_654,N_1595);
xnor U3949 (N_3949,N_1395,N_869);
nor U3950 (N_3950,N_2203,N_827);
xor U3951 (N_3951,N_1184,N_242);
nor U3952 (N_3952,N_124,N_511);
or U3953 (N_3953,N_2101,N_1557);
nand U3954 (N_3954,N_1343,N_1707);
and U3955 (N_3955,N_1315,N_1938);
nand U3956 (N_3956,N_883,N_1782);
nand U3957 (N_3957,N_972,N_745);
and U3958 (N_3958,N_87,N_1308);
xnor U3959 (N_3959,N_282,N_2193);
or U3960 (N_3960,N_759,N_1145);
nand U3961 (N_3961,N_146,N_674);
or U3962 (N_3962,N_2596,N_2436);
nand U3963 (N_3963,N_2569,N_263);
xor U3964 (N_3964,N_2390,N_2523);
or U3965 (N_3965,N_910,N_388);
xor U3966 (N_3966,N_415,N_2117);
and U3967 (N_3967,N_2813,N_12);
or U3968 (N_3968,N_88,N_2678);
and U3969 (N_3969,N_1522,N_899);
and U3970 (N_3970,N_2325,N_1957);
or U3971 (N_3971,N_1237,N_1523);
xnor U3972 (N_3972,N_2280,N_2299);
or U3973 (N_3973,N_2825,N_2087);
nand U3974 (N_3974,N_676,N_593);
and U3975 (N_3975,N_95,N_2849);
xnor U3976 (N_3976,N_1684,N_2295);
xnor U3977 (N_3977,N_394,N_2182);
xor U3978 (N_3978,N_2429,N_2442);
nand U3979 (N_3979,N_1170,N_2012);
xor U3980 (N_3980,N_632,N_2604);
nor U3981 (N_3981,N_1887,N_34);
xor U3982 (N_3982,N_2167,N_2042);
nor U3983 (N_3983,N_931,N_1290);
xnor U3984 (N_3984,N_583,N_265);
nor U3985 (N_3985,N_582,N_576);
or U3986 (N_3986,N_2375,N_2423);
or U3987 (N_3987,N_2200,N_2276);
and U3988 (N_3988,N_2726,N_581);
or U3989 (N_3989,N_2930,N_2305);
and U3990 (N_3990,N_2109,N_2927);
nand U3991 (N_3991,N_82,N_1214);
nand U3992 (N_3992,N_1246,N_2047);
xor U3993 (N_3993,N_2885,N_512);
nand U3994 (N_3994,N_1353,N_1571);
nor U3995 (N_3995,N_2735,N_1786);
nand U3996 (N_3996,N_1449,N_1609);
nor U3997 (N_3997,N_1076,N_1856);
nand U3998 (N_3998,N_408,N_1433);
and U3999 (N_3999,N_2607,N_207);
or U4000 (N_4000,N_846,N_2465);
nand U4001 (N_4001,N_1654,N_1770);
nand U4002 (N_4002,N_2467,N_1429);
or U4003 (N_4003,N_589,N_841);
or U4004 (N_4004,N_1218,N_1920);
nand U4005 (N_4005,N_467,N_2313);
or U4006 (N_4006,N_168,N_971);
nand U4007 (N_4007,N_1899,N_1573);
xnor U4008 (N_4008,N_24,N_2817);
xor U4009 (N_4009,N_1204,N_1703);
and U4010 (N_4010,N_1817,N_744);
nor U4011 (N_4011,N_1334,N_1761);
xor U4012 (N_4012,N_319,N_1215);
xor U4013 (N_4013,N_1370,N_1143);
xnor U4014 (N_4014,N_2645,N_93);
nor U4015 (N_4015,N_335,N_1039);
and U4016 (N_4016,N_174,N_1648);
or U4017 (N_4017,N_2809,N_165);
xor U4018 (N_4018,N_2669,N_1960);
nor U4019 (N_4019,N_2355,N_551);
and U4020 (N_4020,N_2231,N_1912);
or U4021 (N_4021,N_1367,N_2729);
or U4022 (N_4022,N_2323,N_172);
nand U4023 (N_4023,N_482,N_2352);
or U4024 (N_4024,N_983,N_2088);
nand U4025 (N_4025,N_2702,N_2292);
xnor U4026 (N_4026,N_1023,N_556);
nor U4027 (N_4027,N_1427,N_2125);
nor U4028 (N_4028,N_2213,N_2382);
nor U4029 (N_4029,N_1057,N_507);
nor U4030 (N_4030,N_1446,N_1335);
xor U4031 (N_4031,N_1154,N_1203);
xnor U4032 (N_4032,N_1839,N_1852);
xor U4033 (N_4033,N_2074,N_2092);
or U4034 (N_4034,N_1598,N_955);
or U4035 (N_4035,N_2139,N_2389);
nand U4036 (N_4036,N_535,N_559);
nor U4037 (N_4037,N_543,N_298);
xnor U4038 (N_4038,N_2847,N_1896);
nand U4039 (N_4039,N_1964,N_2947);
and U4040 (N_4040,N_2246,N_729);
xnor U4041 (N_4041,N_2068,N_152);
and U4042 (N_4042,N_64,N_2478);
nor U4043 (N_4043,N_552,N_2756);
and U4044 (N_4044,N_2520,N_2222);
xnor U4045 (N_4045,N_2123,N_1126);
and U4046 (N_4046,N_1192,N_2710);
or U4047 (N_4047,N_1788,N_1619);
nor U4048 (N_4048,N_904,N_1317);
nand U4049 (N_4049,N_1160,N_1668);
or U4050 (N_4050,N_2540,N_687);
nand U4051 (N_4051,N_325,N_1583);
and U4052 (N_4052,N_1122,N_1998);
xor U4053 (N_4053,N_1495,N_495);
or U4054 (N_4054,N_321,N_1045);
nand U4055 (N_4055,N_2281,N_1380);
nor U4056 (N_4056,N_2757,N_558);
and U4057 (N_4057,N_2518,N_2096);
or U4058 (N_4058,N_1958,N_246);
or U4059 (N_4059,N_607,N_567);
nor U4060 (N_4060,N_483,N_937);
nor U4061 (N_4061,N_2490,N_500);
xnor U4062 (N_4062,N_925,N_1733);
or U4063 (N_4063,N_197,N_1307);
xnor U4064 (N_4064,N_403,N_1567);
and U4065 (N_4065,N_2821,N_2336);
xor U4066 (N_4066,N_1088,N_2679);
nand U4067 (N_4067,N_300,N_2660);
and U4068 (N_4068,N_1862,N_386);
or U4069 (N_4069,N_2515,N_1863);
nand U4070 (N_4070,N_2881,N_1479);
or U4071 (N_4071,N_2509,N_1728);
or U4072 (N_4072,N_2020,N_1295);
or U4073 (N_4073,N_1106,N_128);
nor U4074 (N_4074,N_1545,N_2081);
xnor U4075 (N_4075,N_969,N_10);
or U4076 (N_4076,N_494,N_1727);
nand U4077 (N_4077,N_2443,N_240);
and U4078 (N_4078,N_705,N_615);
or U4079 (N_4079,N_1118,N_1405);
nor U4080 (N_4080,N_944,N_2170);
and U4081 (N_4081,N_1266,N_1333);
nor U4082 (N_4082,N_2658,N_2620);
nand U4083 (N_4083,N_1150,N_1783);
xnor U4084 (N_4084,N_270,N_481);
nand U4085 (N_4085,N_2315,N_392);
or U4086 (N_4086,N_1085,N_1111);
xor U4087 (N_4087,N_2179,N_2055);
nor U4088 (N_4088,N_2212,N_1201);
nand U4089 (N_4089,N_1316,N_497);
nor U4090 (N_4090,N_2430,N_1773);
nand U4091 (N_4091,N_1243,N_2924);
xor U4092 (N_4092,N_2803,N_166);
nand U4093 (N_4093,N_132,N_1357);
xor U4094 (N_4094,N_41,N_1013);
and U4095 (N_4095,N_1391,N_2242);
nand U4096 (N_4096,N_1093,N_698);
nor U4097 (N_4097,N_2333,N_1432);
nand U4098 (N_4098,N_1600,N_2875);
nand U4099 (N_4099,N_2863,N_1064);
nor U4100 (N_4100,N_330,N_2865);
xor U4101 (N_4101,N_2185,N_2688);
and U4102 (N_4102,N_66,N_2522);
or U4103 (N_4103,N_1984,N_817);
xor U4104 (N_4104,N_470,N_2721);
or U4105 (N_4105,N_1814,N_660);
nor U4106 (N_4106,N_2663,N_2065);
and U4107 (N_4107,N_891,N_1980);
nand U4108 (N_4108,N_2049,N_2);
nor U4109 (N_4109,N_1759,N_800);
nand U4110 (N_4110,N_143,N_1377);
nor U4111 (N_4111,N_1700,N_2100);
and U4112 (N_4112,N_748,N_938);
nand U4113 (N_4113,N_133,N_1274);
or U4114 (N_4114,N_1095,N_267);
or U4115 (N_4115,N_1069,N_2174);
nand U4116 (N_4116,N_1525,N_2161);
nor U4117 (N_4117,N_1442,N_397);
or U4118 (N_4118,N_1115,N_528);
and U4119 (N_4119,N_1,N_2130);
and U4120 (N_4120,N_180,N_2644);
or U4121 (N_4121,N_1242,N_2943);
nand U4122 (N_4122,N_14,N_25);
or U4123 (N_4123,N_2105,N_2331);
xnor U4124 (N_4124,N_1925,N_2444);
nand U4125 (N_4125,N_1302,N_2383);
nor U4126 (N_4126,N_2983,N_2069);
nor U4127 (N_4127,N_864,N_1848);
or U4128 (N_4128,N_2287,N_1436);
xor U4129 (N_4129,N_2226,N_2598);
nor U4130 (N_4130,N_286,N_414);
xnor U4131 (N_4131,N_1168,N_315);
or U4132 (N_4132,N_740,N_234);
or U4133 (N_4133,N_1165,N_2181);
xnor U4134 (N_4134,N_2842,N_1722);
xor U4135 (N_4135,N_1765,N_1652);
or U4136 (N_4136,N_1832,N_212);
and U4137 (N_4137,N_1219,N_802);
and U4138 (N_4138,N_2686,N_2253);
nor U4139 (N_4139,N_2794,N_672);
nand U4140 (N_4140,N_2192,N_624);
and U4141 (N_4141,N_1587,N_1322);
xnor U4142 (N_4142,N_751,N_1482);
xnor U4143 (N_4143,N_1216,N_2855);
and U4144 (N_4144,N_805,N_135);
and U4145 (N_4145,N_608,N_1210);
or U4146 (N_4146,N_1798,N_2499);
or U4147 (N_4147,N_959,N_614);
nand U4148 (N_4148,N_1877,N_1756);
nor U4149 (N_4149,N_520,N_443);
and U4150 (N_4150,N_691,N_1369);
nor U4151 (N_4151,N_1347,N_2078);
nand U4152 (N_4152,N_906,N_871);
or U4153 (N_4153,N_1816,N_665);
or U4154 (N_4154,N_205,N_2908);
nor U4155 (N_4155,N_2790,N_568);
xor U4156 (N_4156,N_1708,N_1949);
and U4157 (N_4157,N_1866,N_2841);
xnor U4158 (N_4158,N_1185,N_715);
nand U4159 (N_4159,N_2427,N_1155);
xor U4160 (N_4160,N_721,N_2554);
and U4161 (N_4161,N_2574,N_518);
nor U4162 (N_4162,N_1345,N_123);
nand U4163 (N_4163,N_1963,N_2512);
and U4164 (N_4164,N_474,N_2102);
nand U4165 (N_4165,N_354,N_2232);
or U4166 (N_4166,N_644,N_2385);
nand U4167 (N_4167,N_2188,N_954);
nor U4168 (N_4168,N_694,N_2911);
or U4169 (N_4169,N_1387,N_2345);
or U4170 (N_4170,N_368,N_998);
xnor U4171 (N_4171,N_1621,N_975);
xor U4172 (N_4172,N_1909,N_1762);
and U4173 (N_4173,N_1471,N_1813);
or U4174 (N_4174,N_1718,N_4);
and U4175 (N_4175,N_9,N_98);
nand U4176 (N_4176,N_673,N_2044);
nor U4177 (N_4177,N_155,N_728);
or U4178 (N_4178,N_2330,N_376);
xnor U4179 (N_4179,N_850,N_226);
xor U4180 (N_4180,N_2884,N_2541);
nand U4181 (N_4181,N_1519,N_2014);
nand U4182 (N_4182,N_2285,N_2033);
nor U4183 (N_4183,N_2731,N_1655);
xor U4184 (N_4184,N_496,N_2406);
nand U4185 (N_4185,N_2822,N_2840);
or U4186 (N_4186,N_942,N_262);
xnor U4187 (N_4187,N_2696,N_1693);
nor U4188 (N_4188,N_2210,N_2023);
nand U4189 (N_4189,N_2815,N_1399);
nand U4190 (N_4190,N_1199,N_249);
nor U4191 (N_4191,N_1574,N_412);
xor U4192 (N_4192,N_2904,N_2119);
or U4193 (N_4193,N_1348,N_53);
nor U4194 (N_4194,N_454,N_1355);
and U4195 (N_4195,N_909,N_1797);
nor U4196 (N_4196,N_1845,N_2335);
and U4197 (N_4197,N_2367,N_1491);
xnor U4198 (N_4198,N_2949,N_150);
xor U4199 (N_4199,N_1800,N_1128);
nor U4200 (N_4200,N_1576,N_2652);
or U4201 (N_4201,N_1691,N_2040);
or U4202 (N_4202,N_2353,N_1535);
or U4203 (N_4203,N_878,N_2668);
nor U4204 (N_4204,N_1445,N_504);
or U4205 (N_4205,N_2394,N_2932);
or U4206 (N_4206,N_2432,N_2289);
nor U4207 (N_4207,N_1407,N_866);
nor U4208 (N_4208,N_2537,N_754);
and U4209 (N_4209,N_1279,N_7);
nor U4210 (N_4210,N_541,N_578);
xor U4211 (N_4211,N_2558,N_2676);
and U4212 (N_4212,N_1062,N_2393);
nor U4213 (N_4213,N_2235,N_2861);
or U4214 (N_4214,N_1867,N_1935);
or U4215 (N_4215,N_775,N_633);
and U4216 (N_4216,N_1382,N_727);
or U4217 (N_4217,N_2641,N_1933);
nor U4218 (N_4218,N_2709,N_243);
or U4219 (N_4219,N_2742,N_2207);
xnor U4220 (N_4220,N_1977,N_1930);
or U4221 (N_4221,N_1420,N_2327);
nor U4222 (N_4222,N_1833,N_2583);
or U4223 (N_4223,N_1550,N_1310);
or U4224 (N_4224,N_2337,N_521);
or U4225 (N_4225,N_777,N_182);
xnor U4226 (N_4226,N_56,N_2479);
nor U4227 (N_4227,N_684,N_1054);
nand U4228 (N_4228,N_1438,N_2782);
and U4229 (N_4229,N_992,N_2632);
nor U4230 (N_4230,N_2800,N_947);
nor U4231 (N_4231,N_570,N_381);
or U4232 (N_4232,N_1083,N_1249);
or U4233 (N_4233,N_2459,N_2629);
nor U4234 (N_4234,N_1685,N_517);
and U4235 (N_4235,N_1822,N_2414);
and U4236 (N_4236,N_1853,N_2896);
nor U4237 (N_4237,N_1238,N_1686);
xnor U4238 (N_4238,N_1627,N_385);
nand U4239 (N_4239,N_2784,N_2530);
nand U4240 (N_4240,N_1098,N_461);
nand U4241 (N_4241,N_1078,N_1704);
xnor U4242 (N_4242,N_2116,N_1460);
nand U4243 (N_4243,N_1419,N_1309);
nor U4244 (N_4244,N_2483,N_2236);
xnor U4245 (N_4245,N_650,N_554);
or U4246 (N_4246,N_1147,N_534);
xor U4247 (N_4247,N_318,N_167);
xnor U4248 (N_4248,N_736,N_489);
xor U4249 (N_4249,N_322,N_2831);
and U4250 (N_4250,N_1534,N_2673);
or U4251 (N_4251,N_1699,N_2184);
nand U4252 (N_4252,N_1670,N_122);
xnor U4253 (N_4253,N_16,N_1231);
and U4254 (N_4254,N_2127,N_2852);
xor U4255 (N_4255,N_550,N_445);
nand U4256 (N_4256,N_2625,N_1323);
and U4257 (N_4257,N_735,N_1679);
and U4258 (N_4258,N_1824,N_363);
and U4259 (N_4259,N_1552,N_1638);
nor U4260 (N_4260,N_2163,N_2326);
and U4261 (N_4261,N_1821,N_2249);
or U4262 (N_4262,N_2050,N_1173);
nor U4263 (N_4263,N_1539,N_600);
and U4264 (N_4264,N_2086,N_594);
and U4265 (N_4265,N_1516,N_1036);
nor U4266 (N_4266,N_2724,N_1620);
nand U4267 (N_4267,N_1597,N_38);
xnor U4268 (N_4268,N_1916,N_1767);
nor U4269 (N_4269,N_2517,N_2738);
nor U4270 (N_4270,N_1341,N_1141);
and U4271 (N_4271,N_54,N_1153);
nor U4272 (N_4272,N_1643,N_1692);
or U4273 (N_4273,N_2199,N_2602);
nor U4274 (N_4274,N_1801,N_2552);
nand U4275 (N_4275,N_743,N_1061);
nand U4276 (N_4276,N_1068,N_2477);
nand U4277 (N_4277,N_236,N_466);
nor U4278 (N_4278,N_1616,N_2437);
or U4279 (N_4279,N_69,N_2036);
nand U4280 (N_4280,N_1019,N_2054);
nand U4281 (N_4281,N_1561,N_1572);
nor U4282 (N_4282,N_1672,N_2539);
or U4283 (N_4283,N_2104,N_2224);
xor U4284 (N_4284,N_390,N_1551);
or U4285 (N_4285,N_1794,N_889);
nor U4286 (N_4286,N_630,N_2239);
xor U4287 (N_4287,N_2936,N_1003);
xor U4288 (N_4288,N_284,N_1646);
and U4289 (N_4289,N_2453,N_1474);
xor U4290 (N_4290,N_2408,N_486);
or U4291 (N_4291,N_2939,N_119);
xor U4292 (N_4292,N_1475,N_1590);
nor U4293 (N_4293,N_1695,N_812);
nand U4294 (N_4294,N_1542,N_2319);
and U4295 (N_4295,N_2187,N_1079);
or U4296 (N_4296,N_848,N_779);
and U4297 (N_4297,N_126,N_2229);
nor U4298 (N_4298,N_96,N_203);
and U4299 (N_4299,N_1356,N_2561);
nand U4300 (N_4300,N_334,N_76);
nand U4301 (N_4301,N_533,N_2475);
and U4302 (N_4302,N_2992,N_776);
and U4303 (N_4303,N_572,N_1688);
nand U4304 (N_4304,N_2056,N_1779);
and U4305 (N_4305,N_564,N_2291);
nand U4306 (N_4306,N_2495,N_2741);
xnor U4307 (N_4307,N_2534,N_682);
and U4308 (N_4308,N_277,N_2799);
nor U4309 (N_4309,N_2888,N_2324);
nor U4310 (N_4310,N_1541,N_339);
and U4311 (N_4311,N_2618,N_1503);
or U4312 (N_4312,N_2657,N_739);
nand U4313 (N_4313,N_919,N_1874);
xnor U4314 (N_4314,N_75,N_1636);
or U4315 (N_4315,N_1674,N_183);
or U4316 (N_4316,N_2786,N_2503);
xor U4317 (N_4317,N_1997,N_257);
and U4318 (N_4318,N_2555,N_2666);
or U4319 (N_4319,N_2418,N_2751);
or U4320 (N_4320,N_1021,N_2820);
nor U4321 (N_4321,N_2882,N_701);
nand U4322 (N_4322,N_2372,N_160);
nand U4323 (N_4323,N_2791,N_2972);
nor U4324 (N_4324,N_2646,N_81);
xor U4325 (N_4325,N_2126,N_1070);
and U4326 (N_4326,N_2938,N_1030);
and U4327 (N_4327,N_1612,N_2460);
or U4328 (N_4328,N_2502,N_2195);
nand U4329 (N_4329,N_22,N_1514);
nand U4330 (N_4330,N_2051,N_657);
nor U4331 (N_4331,N_1180,N_1784);
nand U4332 (N_4332,N_2559,N_241);
and U4333 (N_4333,N_2456,N_1351);
xnor U4334 (N_4334,N_2452,N_1928);
and U4335 (N_4335,N_2446,N_2736);
nor U4336 (N_4336,N_538,N_47);
nand U4337 (N_4337,N_1768,N_2776);
and U4338 (N_4338,N_102,N_1226);
or U4339 (N_4339,N_2631,N_218);
and U4340 (N_4340,N_506,N_2405);
or U4341 (N_4341,N_2740,N_2819);
nor U4342 (N_4342,N_447,N_960);
xnor U4343 (N_4343,N_1675,N_2525);
or U4344 (N_4344,N_2573,N_2879);
and U4345 (N_4345,N_1125,N_1766);
or U4346 (N_4346,N_148,N_2887);
nand U4347 (N_4347,N_2141,N_491);
and U4348 (N_4348,N_1969,N_79);
or U4349 (N_4349,N_101,N_531);
and U4350 (N_4350,N_1642,N_345);
xor U4351 (N_4351,N_437,N_530);
nand U4352 (N_4352,N_1336,N_636);
or U4353 (N_4353,N_713,N_1425);
or U4354 (N_4354,N_223,N_2837);
nor U4355 (N_4355,N_176,N_105);
nor U4356 (N_4356,N_542,N_1873);
nand U4357 (N_4357,N_1403,N_766);
nand U4358 (N_4358,N_1090,N_1205);
nand U4359 (N_4359,N_627,N_795);
nor U4360 (N_4360,N_1424,N_637);
nand U4361 (N_4361,N_667,N_677);
nor U4362 (N_4362,N_1007,N_2664);
xnor U4363 (N_4363,N_2623,N_2508);
or U4364 (N_4364,N_1100,N_1383);
and U4365 (N_4365,N_2415,N_829);
or U4366 (N_4366,N_1074,N_688);
or U4367 (N_4367,N_163,N_2804);
nor U4368 (N_4368,N_2578,N_393);
xor U4369 (N_4369,N_1327,N_1469);
and U4370 (N_4370,N_1831,N_1910);
and U4371 (N_4371,N_2400,N_268);
xor U4372 (N_4372,N_1397,N_2758);
nor U4373 (N_4373,N_2386,N_1990);
and U4374 (N_4374,N_2154,N_1985);
and U4375 (N_4375,N_84,N_510);
nand U4376 (N_4376,N_789,N_907);
or U4377 (N_4377,N_1402,N_2548);
or U4378 (N_4378,N_1566,N_1540);
or U4379 (N_4379,N_880,N_460);
xor U4380 (N_4380,N_2431,N_498);
nor U4381 (N_4381,N_1065,N_617);
nor U4382 (N_4382,N_1629,N_2960);
nor U4383 (N_4383,N_337,N_2600);
nor U4384 (N_4384,N_1802,N_1631);
nor U4385 (N_4385,N_968,N_1002);
nand U4386 (N_4386,N_1558,N_2487);
or U4387 (N_4387,N_1326,N_2061);
or U4388 (N_4388,N_1604,N_1715);
xor U4389 (N_4389,N_967,N_1758);
xor U4390 (N_4390,N_2128,N_2591);
nor U4391 (N_4391,N_1200,N_2565);
or U4392 (N_4392,N_2753,N_151);
or U4393 (N_4393,N_450,N_1271);
nor U4394 (N_4394,N_1872,N_2950);
xnor U4395 (N_4395,N_1888,N_1059);
nand U4396 (N_4396,N_1529,N_716);
xor U4397 (N_4397,N_2493,N_2227);
nor U4398 (N_4398,N_453,N_732);
nand U4399 (N_4399,N_2975,N_1430);
nor U4400 (N_4400,N_141,N_89);
nor U4401 (N_4401,N_162,N_2008);
nor U4402 (N_4402,N_837,N_1384);
nand U4403 (N_4403,N_1982,N_29);
xor U4404 (N_4404,N_845,N_1275);
or U4405 (N_4405,N_206,N_434);
nor U4406 (N_4406,N_1052,N_796);
nand U4407 (N_4407,N_195,N_2168);
and U4408 (N_4408,N_2542,N_2900);
and U4409 (N_4409,N_255,N_1008);
nand U4410 (N_4410,N_1697,N_1940);
or U4411 (N_4411,N_2053,N_2919);
nand U4412 (N_4412,N_310,N_97);
and U4413 (N_4413,N_1494,N_1354);
nand U4414 (N_4414,N_2547,N_2890);
xor U4415 (N_4415,N_916,N_428);
nor U4416 (N_4416,N_2302,N_1349);
and U4417 (N_4417,N_760,N_874);
nand U4418 (N_4418,N_1846,N_2878);
nor U4419 (N_4419,N_563,N_770);
nand U4420 (N_4420,N_1467,N_423);
and U4421 (N_4421,N_2779,N_852);
xnor U4422 (N_4422,N_1952,N_2438);
nor U4423 (N_4423,N_1224,N_2140);
xor U4424 (N_4424,N_1196,N_2332);
xor U4425 (N_4425,N_2091,N_6);
or U4426 (N_4426,N_2486,N_2496);
and U4427 (N_4427,N_733,N_513);
and U4428 (N_4428,N_896,N_2339);
nor U4429 (N_4429,N_427,N_2225);
and U4430 (N_4430,N_2045,N_565);
xnor U4431 (N_4431,N_1630,N_2902);
nor U4432 (N_4432,N_200,N_1239);
xor U4433 (N_4433,N_2917,N_1142);
and U4434 (N_4434,N_2965,N_1086);
and U4435 (N_4435,N_478,N_2019);
and U4436 (N_4436,N_588,N_2944);
nand U4437 (N_4437,N_1101,N_1331);
xnor U4438 (N_4438,N_2387,N_178);
nand U4439 (N_4439,N_2783,N_1966);
xnor U4440 (N_4440,N_37,N_861);
xnor U4441 (N_4441,N_639,N_1461);
xor U4442 (N_4442,N_417,N_2627);
nand U4443 (N_4443,N_2041,N_712);
nand U4444 (N_4444,N_905,N_741);
and U4445 (N_4445,N_2595,N_2457);
or U4446 (N_4446,N_362,N_2572);
xnor U4447 (N_4447,N_865,N_2099);
and U4448 (N_4448,N_2833,N_642);
nor U4449 (N_4449,N_2009,N_1014);
nand U4450 (N_4450,N_314,N_2300);
and U4451 (N_4451,N_2985,N_1988);
nand U4452 (N_4452,N_2746,N_1538);
xnor U4453 (N_4453,N_2874,N_2022);
nor U4454 (N_4454,N_355,N_2198);
or U4455 (N_4455,N_669,N_2316);
or U4456 (N_4456,N_1804,N_1396);
and U4457 (N_4457,N_422,N_2403);
nand U4458 (N_4458,N_2535,N_2762);
or U4459 (N_4459,N_94,N_978);
nand U4460 (N_4460,N_444,N_2921);
or U4461 (N_4461,N_1902,N_1658);
or U4462 (N_4462,N_610,N_2500);
or U4463 (N_4463,N_2308,N_2914);
or U4464 (N_4464,N_643,N_1528);
or U4465 (N_4465,N_1663,N_1499);
xnor U4466 (N_4466,N_213,N_2603);
and U4467 (N_4467,N_806,N_1508);
and U4468 (N_4468,N_1267,N_2160);
xnor U4469 (N_4469,N_529,N_2321);
or U4470 (N_4470,N_2807,N_2118);
nor U4471 (N_4471,N_2706,N_2003);
and U4472 (N_4472,N_19,N_1217);
and U4473 (N_4473,N_1731,N_74);
or U4474 (N_4474,N_2183,N_993);
nor U4475 (N_4475,N_804,N_383);
nand U4476 (N_4476,N_753,N_2103);
nand U4477 (N_4477,N_1454,N_2769);
nand U4478 (N_4478,N_2715,N_836);
or U4479 (N_4479,N_1232,N_378);
xnor U4480 (N_4480,N_2468,N_784);
and U4481 (N_4481,N_1075,N_1772);
and U4482 (N_4482,N_835,N_2370);
xor U4483 (N_4483,N_1730,N_61);
nand U4484 (N_4484,N_2062,N_714);
and U4485 (N_4485,N_1701,N_1834);
nor U4486 (N_4486,N_1806,N_2318);
xnor U4487 (N_4487,N_2998,N_2015);
xnor U4488 (N_4488,N_598,N_158);
nor U4489 (N_4489,N_1042,N_1287);
nor U4490 (N_4490,N_1625,N_1264);
or U4491 (N_4491,N_1073,N_2514);
xor U4492 (N_4492,N_2366,N_1737);
nand U4493 (N_4493,N_1741,N_2259);
nand U4494 (N_4494,N_1386,N_110);
xnor U4495 (N_4495,N_1992,N_1256);
nor U4496 (N_4496,N_2560,N_232);
and U4497 (N_4497,N_1131,N_2994);
nand U4498 (N_4498,N_2553,N_1035);
nand U4499 (N_4499,N_1812,N_2376);
or U4500 (N_4500,N_1192,N_1725);
nor U4501 (N_4501,N_1877,N_119);
nor U4502 (N_4502,N_988,N_1107);
or U4503 (N_4503,N_768,N_1512);
nand U4504 (N_4504,N_1293,N_338);
xor U4505 (N_4505,N_597,N_1363);
xor U4506 (N_4506,N_566,N_1999);
or U4507 (N_4507,N_1057,N_957);
nand U4508 (N_4508,N_2306,N_115);
or U4509 (N_4509,N_2909,N_1570);
or U4510 (N_4510,N_1904,N_131);
xor U4511 (N_4511,N_1670,N_2112);
or U4512 (N_4512,N_1948,N_2738);
and U4513 (N_4513,N_1061,N_1045);
xnor U4514 (N_4514,N_1460,N_780);
or U4515 (N_4515,N_1304,N_2187);
or U4516 (N_4516,N_189,N_2392);
and U4517 (N_4517,N_117,N_1019);
nor U4518 (N_4518,N_644,N_264);
xnor U4519 (N_4519,N_2963,N_1073);
nor U4520 (N_4520,N_1787,N_1126);
nor U4521 (N_4521,N_1601,N_1927);
or U4522 (N_4522,N_360,N_1351);
or U4523 (N_4523,N_2503,N_2551);
and U4524 (N_4524,N_661,N_1988);
nor U4525 (N_4525,N_1982,N_1142);
or U4526 (N_4526,N_1735,N_663);
or U4527 (N_4527,N_882,N_1510);
nor U4528 (N_4528,N_956,N_2823);
or U4529 (N_4529,N_351,N_2);
nor U4530 (N_4530,N_2523,N_1158);
or U4531 (N_4531,N_2639,N_743);
xor U4532 (N_4532,N_2002,N_1633);
nor U4533 (N_4533,N_0,N_1062);
nor U4534 (N_4534,N_1546,N_666);
and U4535 (N_4535,N_2020,N_1790);
nor U4536 (N_4536,N_500,N_2543);
nand U4537 (N_4537,N_2223,N_2474);
xor U4538 (N_4538,N_2663,N_974);
nand U4539 (N_4539,N_1027,N_1474);
or U4540 (N_4540,N_1376,N_1198);
nand U4541 (N_4541,N_1002,N_92);
and U4542 (N_4542,N_1772,N_883);
or U4543 (N_4543,N_1366,N_1291);
xnor U4544 (N_4544,N_1377,N_1987);
or U4545 (N_4545,N_1543,N_2564);
nand U4546 (N_4546,N_902,N_251);
and U4547 (N_4547,N_584,N_532);
xnor U4548 (N_4548,N_1331,N_857);
or U4549 (N_4549,N_697,N_328);
xnor U4550 (N_4550,N_562,N_478);
xnor U4551 (N_4551,N_2203,N_2550);
nor U4552 (N_4552,N_2641,N_105);
nor U4553 (N_4553,N_1640,N_1060);
and U4554 (N_4554,N_465,N_2998);
nor U4555 (N_4555,N_1730,N_1830);
or U4556 (N_4556,N_1571,N_1086);
nand U4557 (N_4557,N_1628,N_2894);
xor U4558 (N_4558,N_2451,N_960);
or U4559 (N_4559,N_579,N_1496);
nand U4560 (N_4560,N_1331,N_1769);
xor U4561 (N_4561,N_998,N_658);
nand U4562 (N_4562,N_351,N_1165);
xnor U4563 (N_4563,N_1860,N_659);
nor U4564 (N_4564,N_684,N_1742);
and U4565 (N_4565,N_1715,N_2056);
xor U4566 (N_4566,N_834,N_79);
nand U4567 (N_4567,N_1309,N_2659);
xnor U4568 (N_4568,N_2392,N_2970);
or U4569 (N_4569,N_2509,N_2813);
nor U4570 (N_4570,N_1100,N_758);
or U4571 (N_4571,N_2549,N_1320);
and U4572 (N_4572,N_1182,N_919);
nor U4573 (N_4573,N_161,N_2709);
nand U4574 (N_4574,N_329,N_575);
nor U4575 (N_4575,N_198,N_1023);
xnor U4576 (N_4576,N_2617,N_1677);
xnor U4577 (N_4577,N_959,N_1452);
and U4578 (N_4578,N_1655,N_1942);
nand U4579 (N_4579,N_1817,N_2558);
and U4580 (N_4580,N_1916,N_971);
nor U4581 (N_4581,N_2273,N_1621);
nand U4582 (N_4582,N_1299,N_311);
and U4583 (N_4583,N_2632,N_1743);
or U4584 (N_4584,N_2442,N_1283);
nand U4585 (N_4585,N_2042,N_1033);
nor U4586 (N_4586,N_2978,N_2669);
xnor U4587 (N_4587,N_387,N_2598);
or U4588 (N_4588,N_1201,N_2370);
nor U4589 (N_4589,N_951,N_1621);
and U4590 (N_4590,N_1149,N_235);
or U4591 (N_4591,N_1329,N_2325);
and U4592 (N_4592,N_2094,N_2354);
nand U4593 (N_4593,N_1619,N_1061);
nor U4594 (N_4594,N_1971,N_650);
xnor U4595 (N_4595,N_1765,N_106);
or U4596 (N_4596,N_2485,N_1305);
nor U4597 (N_4597,N_2941,N_800);
or U4598 (N_4598,N_1903,N_78);
xor U4599 (N_4599,N_853,N_486);
and U4600 (N_4600,N_714,N_529);
xnor U4601 (N_4601,N_2324,N_660);
nand U4602 (N_4602,N_2528,N_573);
or U4603 (N_4603,N_204,N_1004);
nor U4604 (N_4604,N_260,N_2177);
or U4605 (N_4605,N_1187,N_915);
xnor U4606 (N_4606,N_892,N_1416);
nor U4607 (N_4607,N_1259,N_1707);
xor U4608 (N_4608,N_2042,N_1892);
nor U4609 (N_4609,N_1417,N_2843);
or U4610 (N_4610,N_1047,N_1436);
or U4611 (N_4611,N_2463,N_2134);
nor U4612 (N_4612,N_1731,N_2089);
nor U4613 (N_4613,N_305,N_2616);
nor U4614 (N_4614,N_249,N_1961);
and U4615 (N_4615,N_500,N_2178);
xnor U4616 (N_4616,N_1335,N_1774);
or U4617 (N_4617,N_2325,N_2109);
xor U4618 (N_4618,N_1468,N_2867);
nand U4619 (N_4619,N_2543,N_1593);
or U4620 (N_4620,N_2639,N_2605);
nor U4621 (N_4621,N_1830,N_2090);
nand U4622 (N_4622,N_1966,N_1932);
xor U4623 (N_4623,N_878,N_2520);
nand U4624 (N_4624,N_1082,N_2856);
xor U4625 (N_4625,N_293,N_155);
and U4626 (N_4626,N_1106,N_2580);
nor U4627 (N_4627,N_2545,N_249);
and U4628 (N_4628,N_2536,N_604);
nor U4629 (N_4629,N_2484,N_1370);
xnor U4630 (N_4630,N_1481,N_1490);
nor U4631 (N_4631,N_2392,N_2456);
and U4632 (N_4632,N_2531,N_393);
nand U4633 (N_4633,N_2218,N_1430);
and U4634 (N_4634,N_1009,N_1215);
or U4635 (N_4635,N_673,N_2567);
xor U4636 (N_4636,N_981,N_2938);
and U4637 (N_4637,N_2874,N_1043);
and U4638 (N_4638,N_1894,N_231);
and U4639 (N_4639,N_745,N_2511);
nor U4640 (N_4640,N_2637,N_1400);
nand U4641 (N_4641,N_336,N_260);
nor U4642 (N_4642,N_1364,N_2589);
nor U4643 (N_4643,N_2851,N_1613);
nand U4644 (N_4644,N_767,N_20);
or U4645 (N_4645,N_690,N_2824);
and U4646 (N_4646,N_1571,N_2805);
and U4647 (N_4647,N_1858,N_2353);
or U4648 (N_4648,N_2091,N_1022);
or U4649 (N_4649,N_1675,N_2565);
nand U4650 (N_4650,N_1201,N_1857);
or U4651 (N_4651,N_280,N_2749);
nand U4652 (N_4652,N_2974,N_1677);
nand U4653 (N_4653,N_684,N_1979);
nor U4654 (N_4654,N_1842,N_712);
and U4655 (N_4655,N_1980,N_1816);
xnor U4656 (N_4656,N_2390,N_1261);
and U4657 (N_4657,N_2096,N_63);
or U4658 (N_4658,N_716,N_876);
nor U4659 (N_4659,N_188,N_1482);
nand U4660 (N_4660,N_2490,N_2655);
nor U4661 (N_4661,N_241,N_1714);
or U4662 (N_4662,N_2684,N_732);
and U4663 (N_4663,N_544,N_2515);
and U4664 (N_4664,N_707,N_2927);
nand U4665 (N_4665,N_2876,N_2105);
nor U4666 (N_4666,N_1192,N_2266);
nor U4667 (N_4667,N_2972,N_643);
and U4668 (N_4668,N_2139,N_1795);
nand U4669 (N_4669,N_218,N_1951);
nand U4670 (N_4670,N_1607,N_1261);
and U4671 (N_4671,N_1006,N_1844);
and U4672 (N_4672,N_1533,N_1415);
nor U4673 (N_4673,N_1389,N_1727);
and U4674 (N_4674,N_2316,N_1650);
and U4675 (N_4675,N_2412,N_872);
or U4676 (N_4676,N_117,N_1614);
nand U4677 (N_4677,N_2335,N_1824);
nor U4678 (N_4678,N_959,N_432);
nor U4679 (N_4679,N_1497,N_86);
or U4680 (N_4680,N_2408,N_2651);
nand U4681 (N_4681,N_2859,N_89);
nor U4682 (N_4682,N_1552,N_1981);
or U4683 (N_4683,N_2747,N_1613);
nor U4684 (N_4684,N_1764,N_2474);
nor U4685 (N_4685,N_270,N_1558);
and U4686 (N_4686,N_2500,N_1894);
xnor U4687 (N_4687,N_1808,N_1413);
xnor U4688 (N_4688,N_2127,N_346);
nor U4689 (N_4689,N_2824,N_994);
xor U4690 (N_4690,N_1986,N_2740);
or U4691 (N_4691,N_783,N_2811);
nand U4692 (N_4692,N_1403,N_1874);
nor U4693 (N_4693,N_2890,N_948);
and U4694 (N_4694,N_2537,N_521);
xor U4695 (N_4695,N_2237,N_665);
and U4696 (N_4696,N_2145,N_798);
xor U4697 (N_4697,N_1478,N_312);
xnor U4698 (N_4698,N_2206,N_2348);
and U4699 (N_4699,N_1657,N_1889);
xor U4700 (N_4700,N_2417,N_2165);
nor U4701 (N_4701,N_862,N_1662);
or U4702 (N_4702,N_687,N_2289);
and U4703 (N_4703,N_639,N_1174);
xor U4704 (N_4704,N_1592,N_2532);
nand U4705 (N_4705,N_1581,N_2069);
and U4706 (N_4706,N_2822,N_532);
or U4707 (N_4707,N_1057,N_1818);
and U4708 (N_4708,N_2889,N_1307);
and U4709 (N_4709,N_2021,N_1333);
or U4710 (N_4710,N_1095,N_581);
or U4711 (N_4711,N_2678,N_2991);
nand U4712 (N_4712,N_398,N_1797);
and U4713 (N_4713,N_2147,N_1576);
nand U4714 (N_4714,N_464,N_296);
and U4715 (N_4715,N_2535,N_1109);
xor U4716 (N_4716,N_2738,N_1120);
xnor U4717 (N_4717,N_296,N_192);
xor U4718 (N_4718,N_2369,N_638);
nor U4719 (N_4719,N_910,N_1533);
xor U4720 (N_4720,N_1940,N_223);
xnor U4721 (N_4721,N_1613,N_1312);
xnor U4722 (N_4722,N_2328,N_16);
xor U4723 (N_4723,N_2757,N_1920);
nor U4724 (N_4724,N_2085,N_1181);
nand U4725 (N_4725,N_499,N_1993);
or U4726 (N_4726,N_321,N_826);
nor U4727 (N_4727,N_1130,N_2081);
nor U4728 (N_4728,N_82,N_1377);
xnor U4729 (N_4729,N_1615,N_1521);
and U4730 (N_4730,N_2201,N_407);
xnor U4731 (N_4731,N_353,N_1668);
nand U4732 (N_4732,N_845,N_1376);
nor U4733 (N_4733,N_1990,N_45);
nor U4734 (N_4734,N_541,N_2839);
or U4735 (N_4735,N_1388,N_1394);
and U4736 (N_4736,N_1476,N_2930);
nor U4737 (N_4737,N_2001,N_2546);
nand U4738 (N_4738,N_706,N_1412);
and U4739 (N_4739,N_2052,N_2142);
and U4740 (N_4740,N_1664,N_2610);
or U4741 (N_4741,N_184,N_2608);
nand U4742 (N_4742,N_2034,N_2708);
and U4743 (N_4743,N_813,N_699);
and U4744 (N_4744,N_560,N_1212);
xnor U4745 (N_4745,N_1211,N_2932);
nand U4746 (N_4746,N_2540,N_2092);
nor U4747 (N_4747,N_1247,N_674);
and U4748 (N_4748,N_2483,N_2025);
and U4749 (N_4749,N_639,N_1653);
and U4750 (N_4750,N_648,N_66);
or U4751 (N_4751,N_102,N_1804);
xor U4752 (N_4752,N_2927,N_2549);
and U4753 (N_4753,N_1033,N_637);
and U4754 (N_4754,N_2865,N_2861);
and U4755 (N_4755,N_1216,N_544);
nor U4756 (N_4756,N_2670,N_2306);
or U4757 (N_4757,N_1166,N_997);
nand U4758 (N_4758,N_872,N_1154);
xor U4759 (N_4759,N_313,N_1966);
nand U4760 (N_4760,N_1787,N_816);
nand U4761 (N_4761,N_2527,N_317);
or U4762 (N_4762,N_1635,N_2322);
nor U4763 (N_4763,N_160,N_2032);
or U4764 (N_4764,N_2193,N_1386);
xnor U4765 (N_4765,N_2912,N_1555);
and U4766 (N_4766,N_947,N_2356);
nor U4767 (N_4767,N_1132,N_557);
and U4768 (N_4768,N_1086,N_904);
nand U4769 (N_4769,N_1458,N_2821);
nor U4770 (N_4770,N_1198,N_1704);
nor U4771 (N_4771,N_707,N_2233);
nor U4772 (N_4772,N_1938,N_787);
or U4773 (N_4773,N_2212,N_194);
nor U4774 (N_4774,N_1529,N_1057);
nor U4775 (N_4775,N_2812,N_955);
xnor U4776 (N_4776,N_467,N_278);
or U4777 (N_4777,N_2288,N_1140);
xnor U4778 (N_4778,N_1250,N_192);
xnor U4779 (N_4779,N_1079,N_1888);
nand U4780 (N_4780,N_582,N_271);
or U4781 (N_4781,N_366,N_2052);
xor U4782 (N_4782,N_2403,N_2478);
xnor U4783 (N_4783,N_1498,N_1984);
and U4784 (N_4784,N_2255,N_877);
and U4785 (N_4785,N_2488,N_653);
xor U4786 (N_4786,N_1875,N_997);
xor U4787 (N_4787,N_37,N_1288);
and U4788 (N_4788,N_2038,N_2697);
nand U4789 (N_4789,N_221,N_714);
nand U4790 (N_4790,N_76,N_685);
nand U4791 (N_4791,N_2250,N_2320);
nor U4792 (N_4792,N_1649,N_633);
xnor U4793 (N_4793,N_1645,N_2324);
or U4794 (N_4794,N_2971,N_2700);
xnor U4795 (N_4795,N_658,N_2421);
or U4796 (N_4796,N_209,N_896);
nand U4797 (N_4797,N_802,N_286);
nand U4798 (N_4798,N_429,N_1830);
xnor U4799 (N_4799,N_1338,N_1871);
xnor U4800 (N_4800,N_575,N_2929);
or U4801 (N_4801,N_2035,N_1172);
and U4802 (N_4802,N_299,N_1829);
or U4803 (N_4803,N_1392,N_1606);
nor U4804 (N_4804,N_226,N_1071);
xor U4805 (N_4805,N_2050,N_2260);
or U4806 (N_4806,N_1157,N_2208);
xnor U4807 (N_4807,N_1141,N_955);
nand U4808 (N_4808,N_2239,N_2181);
nor U4809 (N_4809,N_492,N_502);
nor U4810 (N_4810,N_253,N_580);
or U4811 (N_4811,N_1255,N_1733);
or U4812 (N_4812,N_1133,N_1412);
nor U4813 (N_4813,N_419,N_2987);
and U4814 (N_4814,N_249,N_2883);
or U4815 (N_4815,N_1484,N_2317);
and U4816 (N_4816,N_2698,N_859);
or U4817 (N_4817,N_127,N_2838);
and U4818 (N_4818,N_898,N_1069);
xor U4819 (N_4819,N_2036,N_839);
and U4820 (N_4820,N_866,N_754);
xor U4821 (N_4821,N_2011,N_1685);
nor U4822 (N_4822,N_266,N_677);
or U4823 (N_4823,N_162,N_1880);
nor U4824 (N_4824,N_714,N_240);
nor U4825 (N_4825,N_1850,N_618);
nor U4826 (N_4826,N_566,N_2723);
nand U4827 (N_4827,N_270,N_1555);
and U4828 (N_4828,N_2095,N_988);
nor U4829 (N_4829,N_1633,N_2082);
xnor U4830 (N_4830,N_1964,N_1963);
nor U4831 (N_4831,N_256,N_2432);
nor U4832 (N_4832,N_884,N_2790);
nor U4833 (N_4833,N_1098,N_1360);
and U4834 (N_4834,N_995,N_51);
nand U4835 (N_4835,N_345,N_208);
and U4836 (N_4836,N_1348,N_1032);
nand U4837 (N_4837,N_758,N_1315);
or U4838 (N_4838,N_2538,N_405);
xor U4839 (N_4839,N_943,N_1014);
nand U4840 (N_4840,N_2199,N_2750);
xor U4841 (N_4841,N_922,N_1257);
nand U4842 (N_4842,N_82,N_2120);
nor U4843 (N_4843,N_1151,N_1815);
or U4844 (N_4844,N_2494,N_2572);
or U4845 (N_4845,N_1723,N_2858);
nand U4846 (N_4846,N_2285,N_2503);
and U4847 (N_4847,N_2161,N_2238);
xor U4848 (N_4848,N_2019,N_1969);
or U4849 (N_4849,N_588,N_126);
xnor U4850 (N_4850,N_2453,N_579);
nor U4851 (N_4851,N_1904,N_2642);
or U4852 (N_4852,N_1507,N_2385);
nand U4853 (N_4853,N_401,N_1671);
nand U4854 (N_4854,N_1384,N_2961);
nor U4855 (N_4855,N_1794,N_2299);
or U4856 (N_4856,N_694,N_905);
and U4857 (N_4857,N_2612,N_2830);
or U4858 (N_4858,N_154,N_1826);
xor U4859 (N_4859,N_2609,N_1527);
or U4860 (N_4860,N_146,N_1734);
nor U4861 (N_4861,N_1108,N_2527);
xnor U4862 (N_4862,N_1182,N_1993);
nand U4863 (N_4863,N_2291,N_1935);
or U4864 (N_4864,N_2849,N_1810);
nand U4865 (N_4865,N_2255,N_855);
or U4866 (N_4866,N_2106,N_122);
xor U4867 (N_4867,N_782,N_1320);
and U4868 (N_4868,N_1008,N_2592);
and U4869 (N_4869,N_759,N_2007);
and U4870 (N_4870,N_883,N_362);
or U4871 (N_4871,N_1705,N_3);
nor U4872 (N_4872,N_2640,N_1817);
and U4873 (N_4873,N_2385,N_579);
xnor U4874 (N_4874,N_2875,N_1426);
xor U4875 (N_4875,N_160,N_1648);
or U4876 (N_4876,N_1289,N_1);
xnor U4877 (N_4877,N_1468,N_2367);
xnor U4878 (N_4878,N_2169,N_2755);
and U4879 (N_4879,N_1930,N_1265);
nor U4880 (N_4880,N_1912,N_524);
and U4881 (N_4881,N_647,N_1795);
or U4882 (N_4882,N_752,N_2424);
nand U4883 (N_4883,N_1188,N_519);
or U4884 (N_4884,N_1083,N_1330);
and U4885 (N_4885,N_2384,N_1265);
nand U4886 (N_4886,N_356,N_2245);
and U4887 (N_4887,N_2104,N_2870);
and U4888 (N_4888,N_2737,N_2881);
xor U4889 (N_4889,N_1748,N_1361);
nand U4890 (N_4890,N_195,N_819);
nor U4891 (N_4891,N_2278,N_247);
or U4892 (N_4892,N_517,N_2113);
nand U4893 (N_4893,N_2764,N_917);
nand U4894 (N_4894,N_1230,N_1392);
nor U4895 (N_4895,N_1517,N_1804);
or U4896 (N_4896,N_2881,N_2594);
nand U4897 (N_4897,N_1681,N_1577);
nor U4898 (N_4898,N_1931,N_1725);
or U4899 (N_4899,N_2227,N_1130);
nor U4900 (N_4900,N_1669,N_1627);
xor U4901 (N_4901,N_630,N_608);
and U4902 (N_4902,N_1717,N_2660);
nor U4903 (N_4903,N_1891,N_2612);
xnor U4904 (N_4904,N_1879,N_1747);
nor U4905 (N_4905,N_95,N_2774);
and U4906 (N_4906,N_2931,N_2351);
nor U4907 (N_4907,N_321,N_869);
nand U4908 (N_4908,N_182,N_1635);
xnor U4909 (N_4909,N_286,N_475);
nand U4910 (N_4910,N_1010,N_1648);
or U4911 (N_4911,N_1567,N_687);
nor U4912 (N_4912,N_960,N_622);
nand U4913 (N_4913,N_2391,N_2170);
nor U4914 (N_4914,N_1690,N_430);
and U4915 (N_4915,N_243,N_2056);
nor U4916 (N_4916,N_1355,N_1408);
and U4917 (N_4917,N_1975,N_11);
xor U4918 (N_4918,N_433,N_2046);
or U4919 (N_4919,N_2701,N_2414);
and U4920 (N_4920,N_1150,N_1889);
or U4921 (N_4921,N_106,N_2994);
nor U4922 (N_4922,N_660,N_1271);
nor U4923 (N_4923,N_157,N_350);
nand U4924 (N_4924,N_2903,N_593);
or U4925 (N_4925,N_2833,N_558);
xor U4926 (N_4926,N_1061,N_1153);
xor U4927 (N_4927,N_1633,N_990);
or U4928 (N_4928,N_2839,N_1600);
and U4929 (N_4929,N_1465,N_609);
or U4930 (N_4930,N_328,N_1861);
or U4931 (N_4931,N_2255,N_1284);
or U4932 (N_4932,N_2194,N_2252);
nand U4933 (N_4933,N_1738,N_853);
and U4934 (N_4934,N_62,N_1274);
and U4935 (N_4935,N_1469,N_549);
xor U4936 (N_4936,N_2174,N_1710);
and U4937 (N_4937,N_2116,N_1381);
nand U4938 (N_4938,N_1790,N_68);
xnor U4939 (N_4939,N_1675,N_1058);
xor U4940 (N_4940,N_288,N_1875);
xnor U4941 (N_4941,N_2761,N_2233);
nor U4942 (N_4942,N_2155,N_274);
nand U4943 (N_4943,N_747,N_1940);
nor U4944 (N_4944,N_1071,N_2082);
nor U4945 (N_4945,N_2210,N_2307);
xnor U4946 (N_4946,N_1525,N_2135);
and U4947 (N_4947,N_578,N_2185);
or U4948 (N_4948,N_198,N_576);
and U4949 (N_4949,N_257,N_1427);
or U4950 (N_4950,N_2849,N_1363);
and U4951 (N_4951,N_2141,N_434);
xnor U4952 (N_4952,N_2070,N_1636);
nor U4953 (N_4953,N_2743,N_70);
or U4954 (N_4954,N_382,N_782);
xnor U4955 (N_4955,N_414,N_1826);
xnor U4956 (N_4956,N_2250,N_637);
nor U4957 (N_4957,N_2869,N_468);
or U4958 (N_4958,N_2162,N_1948);
or U4959 (N_4959,N_2690,N_854);
xor U4960 (N_4960,N_2252,N_2806);
nor U4961 (N_4961,N_569,N_1930);
nand U4962 (N_4962,N_840,N_1823);
and U4963 (N_4963,N_761,N_2476);
nor U4964 (N_4964,N_2098,N_2445);
xor U4965 (N_4965,N_185,N_293);
or U4966 (N_4966,N_803,N_1122);
or U4967 (N_4967,N_1561,N_2179);
nand U4968 (N_4968,N_2056,N_2250);
xnor U4969 (N_4969,N_1694,N_450);
nand U4970 (N_4970,N_1417,N_1126);
and U4971 (N_4971,N_1607,N_2815);
or U4972 (N_4972,N_1796,N_1021);
and U4973 (N_4973,N_1857,N_438);
xnor U4974 (N_4974,N_1988,N_721);
nand U4975 (N_4975,N_2836,N_2653);
nor U4976 (N_4976,N_2264,N_818);
and U4977 (N_4977,N_759,N_911);
nand U4978 (N_4978,N_2656,N_300);
and U4979 (N_4979,N_2325,N_2169);
or U4980 (N_4980,N_2195,N_1993);
or U4981 (N_4981,N_1475,N_1717);
nand U4982 (N_4982,N_391,N_2494);
xnor U4983 (N_4983,N_2404,N_2046);
xor U4984 (N_4984,N_203,N_2646);
nand U4985 (N_4985,N_2021,N_874);
or U4986 (N_4986,N_159,N_876);
or U4987 (N_4987,N_2794,N_989);
nand U4988 (N_4988,N_1136,N_2567);
nand U4989 (N_4989,N_1923,N_246);
xor U4990 (N_4990,N_1845,N_2827);
nor U4991 (N_4991,N_2529,N_1412);
or U4992 (N_4992,N_843,N_141);
or U4993 (N_4993,N_2082,N_2511);
xnor U4994 (N_4994,N_2473,N_333);
nor U4995 (N_4995,N_2945,N_972);
xnor U4996 (N_4996,N_1914,N_2075);
and U4997 (N_4997,N_2420,N_1452);
nand U4998 (N_4998,N_949,N_2127);
xor U4999 (N_4999,N_904,N_2638);
nand U5000 (N_5000,N_275,N_1957);
or U5001 (N_5001,N_2051,N_1954);
and U5002 (N_5002,N_1802,N_346);
and U5003 (N_5003,N_2467,N_562);
nand U5004 (N_5004,N_2952,N_1848);
xor U5005 (N_5005,N_489,N_809);
nor U5006 (N_5006,N_883,N_1217);
nand U5007 (N_5007,N_709,N_1233);
xnor U5008 (N_5008,N_817,N_2120);
or U5009 (N_5009,N_1238,N_933);
nand U5010 (N_5010,N_2658,N_1337);
nor U5011 (N_5011,N_994,N_2450);
nor U5012 (N_5012,N_2196,N_885);
xnor U5013 (N_5013,N_873,N_1977);
xnor U5014 (N_5014,N_2553,N_2991);
xor U5015 (N_5015,N_1165,N_286);
or U5016 (N_5016,N_996,N_943);
nor U5017 (N_5017,N_1601,N_2393);
and U5018 (N_5018,N_1550,N_2735);
xnor U5019 (N_5019,N_1443,N_2949);
nor U5020 (N_5020,N_1560,N_1948);
or U5021 (N_5021,N_2181,N_2818);
nor U5022 (N_5022,N_606,N_302);
xor U5023 (N_5023,N_827,N_1301);
nand U5024 (N_5024,N_699,N_879);
and U5025 (N_5025,N_1375,N_2912);
nand U5026 (N_5026,N_2081,N_905);
and U5027 (N_5027,N_1553,N_2020);
nor U5028 (N_5028,N_2139,N_2605);
or U5029 (N_5029,N_841,N_723);
or U5030 (N_5030,N_207,N_757);
nor U5031 (N_5031,N_876,N_1417);
or U5032 (N_5032,N_1140,N_192);
xor U5033 (N_5033,N_883,N_822);
xnor U5034 (N_5034,N_1456,N_284);
nor U5035 (N_5035,N_1967,N_95);
nor U5036 (N_5036,N_2999,N_1473);
or U5037 (N_5037,N_1736,N_2553);
nand U5038 (N_5038,N_2031,N_1696);
nor U5039 (N_5039,N_1857,N_2474);
nor U5040 (N_5040,N_1552,N_2254);
nor U5041 (N_5041,N_1384,N_2509);
and U5042 (N_5042,N_663,N_1911);
nor U5043 (N_5043,N_652,N_1844);
nor U5044 (N_5044,N_890,N_230);
nand U5045 (N_5045,N_1405,N_311);
or U5046 (N_5046,N_775,N_1362);
and U5047 (N_5047,N_360,N_1675);
xor U5048 (N_5048,N_1778,N_2707);
nor U5049 (N_5049,N_78,N_1005);
nand U5050 (N_5050,N_1089,N_1701);
and U5051 (N_5051,N_2614,N_2725);
nand U5052 (N_5052,N_2163,N_2751);
nor U5053 (N_5053,N_540,N_430);
nand U5054 (N_5054,N_1821,N_1130);
or U5055 (N_5055,N_340,N_1364);
or U5056 (N_5056,N_1030,N_510);
xnor U5057 (N_5057,N_945,N_1823);
nand U5058 (N_5058,N_125,N_2815);
nor U5059 (N_5059,N_1164,N_2990);
nand U5060 (N_5060,N_1471,N_526);
and U5061 (N_5061,N_2862,N_2538);
nor U5062 (N_5062,N_1953,N_1414);
and U5063 (N_5063,N_937,N_1973);
and U5064 (N_5064,N_948,N_471);
nor U5065 (N_5065,N_713,N_1133);
xor U5066 (N_5066,N_1226,N_690);
or U5067 (N_5067,N_498,N_2606);
nand U5068 (N_5068,N_1247,N_2678);
xor U5069 (N_5069,N_169,N_1942);
nand U5070 (N_5070,N_834,N_1795);
nor U5071 (N_5071,N_133,N_823);
nand U5072 (N_5072,N_2859,N_376);
nor U5073 (N_5073,N_2247,N_2439);
nor U5074 (N_5074,N_1953,N_2577);
and U5075 (N_5075,N_1096,N_2431);
or U5076 (N_5076,N_522,N_2082);
or U5077 (N_5077,N_157,N_1373);
nor U5078 (N_5078,N_300,N_1251);
and U5079 (N_5079,N_2536,N_436);
nand U5080 (N_5080,N_74,N_615);
or U5081 (N_5081,N_1042,N_2513);
or U5082 (N_5082,N_890,N_2727);
nand U5083 (N_5083,N_2813,N_233);
and U5084 (N_5084,N_1270,N_2522);
xnor U5085 (N_5085,N_2477,N_2481);
nand U5086 (N_5086,N_994,N_2954);
and U5087 (N_5087,N_577,N_948);
xnor U5088 (N_5088,N_2395,N_1606);
or U5089 (N_5089,N_1808,N_1407);
or U5090 (N_5090,N_2048,N_1026);
xnor U5091 (N_5091,N_1180,N_974);
xor U5092 (N_5092,N_1431,N_2436);
and U5093 (N_5093,N_1789,N_1599);
or U5094 (N_5094,N_534,N_1091);
and U5095 (N_5095,N_806,N_1935);
or U5096 (N_5096,N_1373,N_679);
or U5097 (N_5097,N_1385,N_219);
or U5098 (N_5098,N_1590,N_2350);
nand U5099 (N_5099,N_418,N_1727);
and U5100 (N_5100,N_886,N_2327);
or U5101 (N_5101,N_965,N_847);
or U5102 (N_5102,N_93,N_2255);
and U5103 (N_5103,N_2076,N_1708);
xor U5104 (N_5104,N_386,N_2584);
nor U5105 (N_5105,N_260,N_2820);
or U5106 (N_5106,N_1999,N_2491);
or U5107 (N_5107,N_1619,N_2531);
and U5108 (N_5108,N_2781,N_1634);
nor U5109 (N_5109,N_2491,N_2450);
and U5110 (N_5110,N_2009,N_204);
nor U5111 (N_5111,N_427,N_261);
xor U5112 (N_5112,N_782,N_571);
xor U5113 (N_5113,N_355,N_2002);
or U5114 (N_5114,N_1164,N_2188);
xnor U5115 (N_5115,N_869,N_271);
or U5116 (N_5116,N_73,N_204);
nor U5117 (N_5117,N_1525,N_2113);
and U5118 (N_5118,N_1384,N_660);
nand U5119 (N_5119,N_2217,N_1514);
nand U5120 (N_5120,N_1137,N_2675);
xor U5121 (N_5121,N_2878,N_110);
and U5122 (N_5122,N_2116,N_595);
nor U5123 (N_5123,N_131,N_2300);
and U5124 (N_5124,N_369,N_1167);
or U5125 (N_5125,N_1992,N_2171);
or U5126 (N_5126,N_2817,N_2621);
xnor U5127 (N_5127,N_1456,N_1052);
nor U5128 (N_5128,N_1760,N_1662);
and U5129 (N_5129,N_1805,N_2553);
and U5130 (N_5130,N_1460,N_1265);
nor U5131 (N_5131,N_2405,N_214);
nand U5132 (N_5132,N_1225,N_2115);
nor U5133 (N_5133,N_1169,N_1399);
xnor U5134 (N_5134,N_1863,N_254);
and U5135 (N_5135,N_2971,N_2518);
and U5136 (N_5136,N_1373,N_485);
xor U5137 (N_5137,N_2678,N_1936);
and U5138 (N_5138,N_1221,N_874);
or U5139 (N_5139,N_2600,N_837);
nor U5140 (N_5140,N_770,N_2468);
nor U5141 (N_5141,N_988,N_465);
xor U5142 (N_5142,N_2519,N_2896);
nor U5143 (N_5143,N_2624,N_1802);
nor U5144 (N_5144,N_1912,N_1745);
nor U5145 (N_5145,N_2584,N_1096);
xnor U5146 (N_5146,N_1309,N_51);
or U5147 (N_5147,N_1265,N_295);
nand U5148 (N_5148,N_1472,N_499);
nand U5149 (N_5149,N_2243,N_1799);
nor U5150 (N_5150,N_969,N_2817);
nor U5151 (N_5151,N_2101,N_104);
xnor U5152 (N_5152,N_2846,N_1889);
or U5153 (N_5153,N_2411,N_917);
xnor U5154 (N_5154,N_2414,N_161);
xor U5155 (N_5155,N_1046,N_1737);
nand U5156 (N_5156,N_1004,N_1000);
or U5157 (N_5157,N_1852,N_821);
nor U5158 (N_5158,N_1996,N_789);
nor U5159 (N_5159,N_2197,N_554);
and U5160 (N_5160,N_1407,N_1983);
xor U5161 (N_5161,N_1561,N_671);
or U5162 (N_5162,N_351,N_1841);
nor U5163 (N_5163,N_2586,N_2122);
and U5164 (N_5164,N_852,N_2813);
nor U5165 (N_5165,N_1363,N_199);
nor U5166 (N_5166,N_2754,N_453);
nor U5167 (N_5167,N_2569,N_2878);
nor U5168 (N_5168,N_2703,N_764);
and U5169 (N_5169,N_2023,N_1602);
nor U5170 (N_5170,N_2074,N_2431);
and U5171 (N_5171,N_1005,N_2147);
or U5172 (N_5172,N_508,N_1428);
nor U5173 (N_5173,N_1535,N_2424);
nand U5174 (N_5174,N_2719,N_983);
or U5175 (N_5175,N_2582,N_156);
nor U5176 (N_5176,N_2177,N_2568);
nor U5177 (N_5177,N_1983,N_1161);
nand U5178 (N_5178,N_191,N_1198);
xnor U5179 (N_5179,N_707,N_2096);
or U5180 (N_5180,N_2181,N_337);
nor U5181 (N_5181,N_1601,N_543);
xor U5182 (N_5182,N_2925,N_1346);
nor U5183 (N_5183,N_2653,N_2015);
xnor U5184 (N_5184,N_388,N_946);
nand U5185 (N_5185,N_2375,N_2984);
xnor U5186 (N_5186,N_1575,N_419);
xor U5187 (N_5187,N_2815,N_2857);
nor U5188 (N_5188,N_1816,N_480);
and U5189 (N_5189,N_144,N_2877);
and U5190 (N_5190,N_145,N_1384);
nor U5191 (N_5191,N_1297,N_1227);
nor U5192 (N_5192,N_1582,N_685);
or U5193 (N_5193,N_662,N_939);
nor U5194 (N_5194,N_1964,N_139);
nand U5195 (N_5195,N_271,N_720);
nor U5196 (N_5196,N_2561,N_1814);
xor U5197 (N_5197,N_912,N_372);
xor U5198 (N_5198,N_2967,N_880);
nand U5199 (N_5199,N_423,N_455);
nand U5200 (N_5200,N_936,N_588);
nor U5201 (N_5201,N_505,N_2042);
nand U5202 (N_5202,N_2724,N_2059);
xnor U5203 (N_5203,N_624,N_105);
nand U5204 (N_5204,N_2138,N_2678);
xnor U5205 (N_5205,N_2205,N_2088);
nor U5206 (N_5206,N_1756,N_412);
nor U5207 (N_5207,N_2149,N_1673);
xor U5208 (N_5208,N_2428,N_438);
nand U5209 (N_5209,N_595,N_1310);
or U5210 (N_5210,N_2961,N_911);
nand U5211 (N_5211,N_1812,N_492);
xnor U5212 (N_5212,N_1489,N_2290);
xnor U5213 (N_5213,N_2211,N_339);
nand U5214 (N_5214,N_1299,N_1673);
or U5215 (N_5215,N_868,N_1989);
xor U5216 (N_5216,N_1981,N_2529);
xnor U5217 (N_5217,N_849,N_1899);
nand U5218 (N_5218,N_1784,N_2092);
xnor U5219 (N_5219,N_1257,N_2158);
or U5220 (N_5220,N_162,N_1659);
nor U5221 (N_5221,N_996,N_1327);
nor U5222 (N_5222,N_2781,N_2454);
nor U5223 (N_5223,N_1195,N_2858);
or U5224 (N_5224,N_1356,N_1564);
xnor U5225 (N_5225,N_24,N_454);
nor U5226 (N_5226,N_1436,N_2957);
or U5227 (N_5227,N_237,N_1148);
and U5228 (N_5228,N_1925,N_661);
nand U5229 (N_5229,N_2194,N_2556);
xor U5230 (N_5230,N_2586,N_2718);
nor U5231 (N_5231,N_2833,N_1109);
or U5232 (N_5232,N_1295,N_1466);
nor U5233 (N_5233,N_1868,N_515);
or U5234 (N_5234,N_1702,N_1467);
xor U5235 (N_5235,N_958,N_993);
nand U5236 (N_5236,N_622,N_2579);
nand U5237 (N_5237,N_1540,N_2915);
and U5238 (N_5238,N_2387,N_1927);
xnor U5239 (N_5239,N_2922,N_1594);
and U5240 (N_5240,N_436,N_1595);
or U5241 (N_5241,N_548,N_2771);
nand U5242 (N_5242,N_1604,N_1427);
or U5243 (N_5243,N_925,N_1090);
xor U5244 (N_5244,N_1124,N_1894);
nor U5245 (N_5245,N_595,N_575);
xnor U5246 (N_5246,N_2364,N_1674);
xnor U5247 (N_5247,N_1772,N_847);
xor U5248 (N_5248,N_25,N_2959);
or U5249 (N_5249,N_1308,N_2649);
and U5250 (N_5250,N_813,N_2537);
and U5251 (N_5251,N_725,N_2005);
xor U5252 (N_5252,N_614,N_1167);
xnor U5253 (N_5253,N_331,N_328);
nor U5254 (N_5254,N_1921,N_1611);
xnor U5255 (N_5255,N_1554,N_2235);
nor U5256 (N_5256,N_2678,N_1288);
nand U5257 (N_5257,N_2646,N_1857);
or U5258 (N_5258,N_2512,N_23);
and U5259 (N_5259,N_476,N_2734);
xnor U5260 (N_5260,N_1512,N_2867);
nand U5261 (N_5261,N_2752,N_544);
nand U5262 (N_5262,N_754,N_1081);
or U5263 (N_5263,N_2242,N_315);
and U5264 (N_5264,N_954,N_199);
nor U5265 (N_5265,N_1351,N_1216);
nor U5266 (N_5266,N_2332,N_2990);
xnor U5267 (N_5267,N_2103,N_1397);
nor U5268 (N_5268,N_2134,N_1731);
xor U5269 (N_5269,N_2974,N_1803);
nand U5270 (N_5270,N_1037,N_2636);
nor U5271 (N_5271,N_950,N_766);
nor U5272 (N_5272,N_2290,N_2662);
xor U5273 (N_5273,N_1486,N_762);
or U5274 (N_5274,N_548,N_141);
nand U5275 (N_5275,N_2611,N_1434);
nand U5276 (N_5276,N_778,N_1288);
nand U5277 (N_5277,N_2644,N_2954);
nand U5278 (N_5278,N_2672,N_976);
and U5279 (N_5279,N_2840,N_1773);
nand U5280 (N_5280,N_2681,N_1273);
xnor U5281 (N_5281,N_2458,N_1231);
nand U5282 (N_5282,N_2726,N_715);
xnor U5283 (N_5283,N_291,N_423);
xnor U5284 (N_5284,N_1434,N_2666);
xnor U5285 (N_5285,N_2404,N_425);
nand U5286 (N_5286,N_1172,N_2389);
and U5287 (N_5287,N_1387,N_2718);
nor U5288 (N_5288,N_2325,N_1544);
and U5289 (N_5289,N_1989,N_834);
or U5290 (N_5290,N_2860,N_182);
nand U5291 (N_5291,N_1249,N_960);
nand U5292 (N_5292,N_798,N_2718);
and U5293 (N_5293,N_1072,N_1839);
nor U5294 (N_5294,N_1804,N_360);
and U5295 (N_5295,N_2715,N_2696);
nand U5296 (N_5296,N_415,N_2543);
nand U5297 (N_5297,N_134,N_361);
xor U5298 (N_5298,N_291,N_2388);
nand U5299 (N_5299,N_2417,N_2005);
nand U5300 (N_5300,N_406,N_628);
or U5301 (N_5301,N_1382,N_275);
and U5302 (N_5302,N_1256,N_716);
xor U5303 (N_5303,N_2100,N_285);
and U5304 (N_5304,N_1540,N_2491);
nor U5305 (N_5305,N_1324,N_1206);
and U5306 (N_5306,N_2935,N_1805);
or U5307 (N_5307,N_2372,N_2773);
nand U5308 (N_5308,N_2261,N_787);
and U5309 (N_5309,N_1405,N_495);
nand U5310 (N_5310,N_1085,N_1743);
nor U5311 (N_5311,N_2451,N_267);
xor U5312 (N_5312,N_1308,N_416);
xor U5313 (N_5313,N_387,N_1659);
nor U5314 (N_5314,N_405,N_113);
xor U5315 (N_5315,N_197,N_2776);
nand U5316 (N_5316,N_372,N_470);
xnor U5317 (N_5317,N_2210,N_1496);
nand U5318 (N_5318,N_2509,N_2174);
and U5319 (N_5319,N_1631,N_945);
or U5320 (N_5320,N_2441,N_2415);
nand U5321 (N_5321,N_681,N_927);
or U5322 (N_5322,N_1274,N_856);
and U5323 (N_5323,N_1681,N_2869);
nand U5324 (N_5324,N_1066,N_327);
xnor U5325 (N_5325,N_237,N_221);
nor U5326 (N_5326,N_2436,N_2073);
xnor U5327 (N_5327,N_2528,N_2875);
nand U5328 (N_5328,N_1914,N_446);
xnor U5329 (N_5329,N_2560,N_1975);
nand U5330 (N_5330,N_2526,N_1306);
or U5331 (N_5331,N_283,N_1653);
xor U5332 (N_5332,N_2648,N_1549);
nor U5333 (N_5333,N_298,N_124);
nand U5334 (N_5334,N_1696,N_2790);
and U5335 (N_5335,N_2736,N_2391);
nand U5336 (N_5336,N_368,N_2585);
nand U5337 (N_5337,N_2997,N_1517);
nor U5338 (N_5338,N_2064,N_1472);
and U5339 (N_5339,N_2398,N_556);
nor U5340 (N_5340,N_1943,N_1276);
xor U5341 (N_5341,N_1772,N_720);
nand U5342 (N_5342,N_1745,N_865);
or U5343 (N_5343,N_250,N_973);
or U5344 (N_5344,N_1979,N_2541);
xnor U5345 (N_5345,N_2677,N_987);
nand U5346 (N_5346,N_2001,N_2209);
xor U5347 (N_5347,N_2988,N_1683);
or U5348 (N_5348,N_418,N_1765);
and U5349 (N_5349,N_437,N_1601);
nand U5350 (N_5350,N_1769,N_2828);
or U5351 (N_5351,N_1090,N_1923);
xnor U5352 (N_5352,N_1638,N_1425);
and U5353 (N_5353,N_1438,N_72);
xor U5354 (N_5354,N_1751,N_216);
xor U5355 (N_5355,N_1927,N_1199);
nor U5356 (N_5356,N_1202,N_2157);
nor U5357 (N_5357,N_1058,N_1928);
and U5358 (N_5358,N_974,N_2144);
or U5359 (N_5359,N_994,N_2799);
nand U5360 (N_5360,N_1401,N_1028);
nand U5361 (N_5361,N_41,N_2014);
or U5362 (N_5362,N_1898,N_2102);
or U5363 (N_5363,N_862,N_1715);
and U5364 (N_5364,N_1534,N_1761);
xnor U5365 (N_5365,N_2379,N_463);
and U5366 (N_5366,N_2344,N_223);
xor U5367 (N_5367,N_318,N_772);
nor U5368 (N_5368,N_2890,N_1904);
nand U5369 (N_5369,N_2417,N_860);
and U5370 (N_5370,N_852,N_2140);
nor U5371 (N_5371,N_1817,N_743);
and U5372 (N_5372,N_449,N_2885);
or U5373 (N_5373,N_1259,N_905);
nor U5374 (N_5374,N_1182,N_2069);
nand U5375 (N_5375,N_2302,N_1747);
or U5376 (N_5376,N_2571,N_1762);
nand U5377 (N_5377,N_241,N_2405);
nor U5378 (N_5378,N_1306,N_2573);
nand U5379 (N_5379,N_982,N_2321);
xor U5380 (N_5380,N_351,N_582);
and U5381 (N_5381,N_2415,N_2717);
nor U5382 (N_5382,N_1144,N_2463);
nor U5383 (N_5383,N_2074,N_1166);
nand U5384 (N_5384,N_1049,N_193);
nor U5385 (N_5385,N_1594,N_2683);
and U5386 (N_5386,N_289,N_1565);
nand U5387 (N_5387,N_184,N_177);
or U5388 (N_5388,N_1981,N_2440);
and U5389 (N_5389,N_497,N_2453);
and U5390 (N_5390,N_2900,N_1317);
or U5391 (N_5391,N_2328,N_2511);
nand U5392 (N_5392,N_2904,N_2643);
nor U5393 (N_5393,N_1410,N_954);
nand U5394 (N_5394,N_916,N_2236);
and U5395 (N_5395,N_1076,N_2717);
or U5396 (N_5396,N_2414,N_2800);
xor U5397 (N_5397,N_2913,N_2434);
nand U5398 (N_5398,N_459,N_2172);
and U5399 (N_5399,N_2450,N_2938);
or U5400 (N_5400,N_1590,N_1143);
nor U5401 (N_5401,N_327,N_882);
or U5402 (N_5402,N_2253,N_46);
and U5403 (N_5403,N_1093,N_1820);
nand U5404 (N_5404,N_1653,N_2348);
xor U5405 (N_5405,N_2042,N_2003);
nand U5406 (N_5406,N_2505,N_465);
or U5407 (N_5407,N_1503,N_1291);
and U5408 (N_5408,N_1435,N_2087);
and U5409 (N_5409,N_2309,N_571);
nand U5410 (N_5410,N_1803,N_563);
and U5411 (N_5411,N_2665,N_2165);
xor U5412 (N_5412,N_296,N_719);
xor U5413 (N_5413,N_1561,N_1107);
nand U5414 (N_5414,N_910,N_2398);
or U5415 (N_5415,N_1729,N_2069);
xnor U5416 (N_5416,N_1278,N_279);
or U5417 (N_5417,N_2539,N_2633);
nand U5418 (N_5418,N_263,N_467);
nor U5419 (N_5419,N_2189,N_554);
xor U5420 (N_5420,N_2836,N_1661);
xor U5421 (N_5421,N_531,N_2957);
xor U5422 (N_5422,N_2615,N_257);
xor U5423 (N_5423,N_2320,N_213);
and U5424 (N_5424,N_1109,N_2890);
and U5425 (N_5425,N_570,N_808);
xor U5426 (N_5426,N_941,N_2330);
xnor U5427 (N_5427,N_1935,N_2456);
and U5428 (N_5428,N_865,N_498);
and U5429 (N_5429,N_346,N_1316);
and U5430 (N_5430,N_531,N_844);
nand U5431 (N_5431,N_2503,N_1553);
nand U5432 (N_5432,N_491,N_2026);
xor U5433 (N_5433,N_974,N_2029);
xor U5434 (N_5434,N_2878,N_1373);
nand U5435 (N_5435,N_1553,N_152);
xnor U5436 (N_5436,N_2910,N_784);
nor U5437 (N_5437,N_2503,N_69);
and U5438 (N_5438,N_2038,N_2834);
and U5439 (N_5439,N_2089,N_2058);
and U5440 (N_5440,N_1754,N_1881);
and U5441 (N_5441,N_2471,N_2745);
and U5442 (N_5442,N_104,N_1074);
and U5443 (N_5443,N_1837,N_2487);
xor U5444 (N_5444,N_725,N_2223);
nor U5445 (N_5445,N_1656,N_382);
or U5446 (N_5446,N_2924,N_996);
xnor U5447 (N_5447,N_946,N_2834);
or U5448 (N_5448,N_2527,N_1982);
xor U5449 (N_5449,N_2585,N_714);
nand U5450 (N_5450,N_2550,N_1126);
nand U5451 (N_5451,N_1778,N_1780);
nand U5452 (N_5452,N_694,N_478);
xnor U5453 (N_5453,N_846,N_1049);
or U5454 (N_5454,N_685,N_1117);
or U5455 (N_5455,N_2425,N_2052);
nor U5456 (N_5456,N_445,N_2279);
nand U5457 (N_5457,N_231,N_1526);
nor U5458 (N_5458,N_2209,N_1290);
xnor U5459 (N_5459,N_2152,N_2822);
nor U5460 (N_5460,N_170,N_478);
and U5461 (N_5461,N_2003,N_307);
nand U5462 (N_5462,N_651,N_450);
or U5463 (N_5463,N_2984,N_817);
xnor U5464 (N_5464,N_1782,N_2915);
xor U5465 (N_5465,N_406,N_1274);
or U5466 (N_5466,N_804,N_2671);
and U5467 (N_5467,N_1341,N_2737);
and U5468 (N_5468,N_1946,N_272);
and U5469 (N_5469,N_1199,N_772);
xor U5470 (N_5470,N_1624,N_41);
nor U5471 (N_5471,N_1646,N_734);
and U5472 (N_5472,N_159,N_2898);
xnor U5473 (N_5473,N_2624,N_2596);
nand U5474 (N_5474,N_1301,N_2536);
and U5475 (N_5475,N_1620,N_1270);
nor U5476 (N_5476,N_2292,N_2328);
and U5477 (N_5477,N_2138,N_1845);
nand U5478 (N_5478,N_303,N_2236);
or U5479 (N_5479,N_68,N_1091);
and U5480 (N_5480,N_2610,N_148);
and U5481 (N_5481,N_2371,N_1729);
xor U5482 (N_5482,N_972,N_276);
nor U5483 (N_5483,N_246,N_168);
and U5484 (N_5484,N_1274,N_965);
and U5485 (N_5485,N_1241,N_2886);
nand U5486 (N_5486,N_907,N_2599);
and U5487 (N_5487,N_2825,N_690);
xor U5488 (N_5488,N_1511,N_1118);
or U5489 (N_5489,N_2687,N_1662);
xor U5490 (N_5490,N_1040,N_940);
xnor U5491 (N_5491,N_2502,N_1426);
and U5492 (N_5492,N_2660,N_718);
nor U5493 (N_5493,N_2864,N_786);
xor U5494 (N_5494,N_1120,N_1609);
or U5495 (N_5495,N_2788,N_1202);
xor U5496 (N_5496,N_2761,N_753);
and U5497 (N_5497,N_198,N_2953);
or U5498 (N_5498,N_409,N_179);
nand U5499 (N_5499,N_2790,N_2333);
and U5500 (N_5500,N_1126,N_2667);
nor U5501 (N_5501,N_189,N_1701);
nand U5502 (N_5502,N_693,N_2925);
xor U5503 (N_5503,N_354,N_745);
and U5504 (N_5504,N_2055,N_742);
nand U5505 (N_5505,N_1582,N_2735);
and U5506 (N_5506,N_700,N_2131);
xnor U5507 (N_5507,N_788,N_1259);
nand U5508 (N_5508,N_1935,N_890);
and U5509 (N_5509,N_1879,N_138);
and U5510 (N_5510,N_1208,N_1244);
or U5511 (N_5511,N_210,N_1614);
nor U5512 (N_5512,N_1564,N_2416);
or U5513 (N_5513,N_1770,N_2629);
and U5514 (N_5514,N_2210,N_2304);
nand U5515 (N_5515,N_1160,N_997);
and U5516 (N_5516,N_641,N_990);
nand U5517 (N_5517,N_1128,N_2208);
xor U5518 (N_5518,N_2186,N_1397);
nand U5519 (N_5519,N_788,N_2406);
xor U5520 (N_5520,N_2777,N_1053);
xor U5521 (N_5521,N_312,N_206);
nor U5522 (N_5522,N_336,N_2081);
xor U5523 (N_5523,N_2362,N_2539);
nand U5524 (N_5524,N_2337,N_279);
or U5525 (N_5525,N_795,N_425);
and U5526 (N_5526,N_1345,N_2994);
nor U5527 (N_5527,N_406,N_198);
nor U5528 (N_5528,N_2557,N_2951);
and U5529 (N_5529,N_541,N_9);
and U5530 (N_5530,N_2799,N_116);
nand U5531 (N_5531,N_1490,N_680);
nand U5532 (N_5532,N_493,N_1286);
nand U5533 (N_5533,N_547,N_607);
or U5534 (N_5534,N_2364,N_1935);
and U5535 (N_5535,N_2744,N_2950);
and U5536 (N_5536,N_907,N_1907);
and U5537 (N_5537,N_367,N_1720);
nor U5538 (N_5538,N_976,N_1448);
nor U5539 (N_5539,N_2064,N_1371);
xor U5540 (N_5540,N_2593,N_1043);
or U5541 (N_5541,N_587,N_1687);
and U5542 (N_5542,N_779,N_1553);
nand U5543 (N_5543,N_662,N_426);
or U5544 (N_5544,N_2068,N_77);
or U5545 (N_5545,N_2977,N_539);
xor U5546 (N_5546,N_1327,N_2297);
nand U5547 (N_5547,N_2275,N_69);
nand U5548 (N_5548,N_1682,N_2911);
xor U5549 (N_5549,N_2839,N_2598);
xnor U5550 (N_5550,N_270,N_2288);
xor U5551 (N_5551,N_90,N_165);
or U5552 (N_5552,N_1703,N_2475);
xor U5553 (N_5553,N_2442,N_1869);
xnor U5554 (N_5554,N_2308,N_878);
nand U5555 (N_5555,N_2039,N_1626);
nand U5556 (N_5556,N_2981,N_1264);
nor U5557 (N_5557,N_2306,N_1310);
xor U5558 (N_5558,N_1910,N_1440);
and U5559 (N_5559,N_2178,N_2819);
xnor U5560 (N_5560,N_2741,N_140);
nor U5561 (N_5561,N_1149,N_939);
and U5562 (N_5562,N_2731,N_2231);
and U5563 (N_5563,N_646,N_232);
xnor U5564 (N_5564,N_811,N_1534);
or U5565 (N_5565,N_1111,N_2106);
nand U5566 (N_5566,N_1350,N_1977);
or U5567 (N_5567,N_241,N_260);
or U5568 (N_5568,N_1650,N_2487);
or U5569 (N_5569,N_1187,N_453);
nand U5570 (N_5570,N_79,N_2268);
xor U5571 (N_5571,N_2273,N_132);
nor U5572 (N_5572,N_1206,N_2948);
xnor U5573 (N_5573,N_1399,N_449);
nor U5574 (N_5574,N_868,N_1983);
or U5575 (N_5575,N_2749,N_367);
nor U5576 (N_5576,N_1735,N_1169);
xor U5577 (N_5577,N_2448,N_2663);
xor U5578 (N_5578,N_1229,N_2175);
nand U5579 (N_5579,N_2556,N_1276);
or U5580 (N_5580,N_1743,N_2044);
and U5581 (N_5581,N_1509,N_2376);
or U5582 (N_5582,N_2122,N_156);
or U5583 (N_5583,N_2507,N_2114);
and U5584 (N_5584,N_2338,N_2380);
nor U5585 (N_5585,N_1437,N_2113);
nand U5586 (N_5586,N_1428,N_2616);
and U5587 (N_5587,N_2808,N_1568);
or U5588 (N_5588,N_2544,N_2819);
nor U5589 (N_5589,N_2686,N_1887);
nand U5590 (N_5590,N_2280,N_2920);
and U5591 (N_5591,N_2451,N_2015);
or U5592 (N_5592,N_1885,N_2615);
xnor U5593 (N_5593,N_792,N_1198);
nor U5594 (N_5594,N_2212,N_1415);
nor U5595 (N_5595,N_2944,N_278);
nand U5596 (N_5596,N_1157,N_2666);
nand U5597 (N_5597,N_643,N_2700);
nor U5598 (N_5598,N_178,N_1287);
or U5599 (N_5599,N_328,N_1139);
and U5600 (N_5600,N_841,N_1153);
nand U5601 (N_5601,N_1997,N_2934);
nand U5602 (N_5602,N_580,N_2026);
nor U5603 (N_5603,N_1848,N_350);
nor U5604 (N_5604,N_2462,N_2065);
xnor U5605 (N_5605,N_105,N_313);
nand U5606 (N_5606,N_2324,N_2735);
xor U5607 (N_5607,N_2751,N_2726);
nor U5608 (N_5608,N_845,N_1496);
and U5609 (N_5609,N_2147,N_1992);
nor U5610 (N_5610,N_300,N_442);
nand U5611 (N_5611,N_2801,N_1357);
nor U5612 (N_5612,N_1558,N_2082);
xnor U5613 (N_5613,N_466,N_1345);
nand U5614 (N_5614,N_1204,N_2329);
and U5615 (N_5615,N_1476,N_1999);
xor U5616 (N_5616,N_851,N_307);
and U5617 (N_5617,N_487,N_1670);
and U5618 (N_5618,N_653,N_1106);
xor U5619 (N_5619,N_2279,N_1632);
or U5620 (N_5620,N_697,N_2001);
and U5621 (N_5621,N_179,N_1629);
nand U5622 (N_5622,N_2659,N_10);
nand U5623 (N_5623,N_2493,N_1143);
nor U5624 (N_5624,N_48,N_1350);
and U5625 (N_5625,N_449,N_891);
xor U5626 (N_5626,N_407,N_2652);
xnor U5627 (N_5627,N_1116,N_1918);
nor U5628 (N_5628,N_1052,N_2939);
nand U5629 (N_5629,N_755,N_524);
nand U5630 (N_5630,N_2661,N_2285);
xnor U5631 (N_5631,N_2743,N_77);
nand U5632 (N_5632,N_2565,N_511);
and U5633 (N_5633,N_63,N_2210);
nor U5634 (N_5634,N_1007,N_2716);
nor U5635 (N_5635,N_2701,N_435);
nand U5636 (N_5636,N_1748,N_2775);
nand U5637 (N_5637,N_1821,N_2767);
or U5638 (N_5638,N_1507,N_2673);
or U5639 (N_5639,N_2138,N_2109);
nor U5640 (N_5640,N_208,N_2864);
nor U5641 (N_5641,N_413,N_2545);
nand U5642 (N_5642,N_950,N_937);
nor U5643 (N_5643,N_2371,N_1857);
nor U5644 (N_5644,N_1959,N_1361);
nor U5645 (N_5645,N_940,N_1037);
xnor U5646 (N_5646,N_976,N_2580);
xnor U5647 (N_5647,N_2315,N_313);
xnor U5648 (N_5648,N_1333,N_947);
nor U5649 (N_5649,N_1274,N_2813);
nand U5650 (N_5650,N_1960,N_1395);
nand U5651 (N_5651,N_80,N_534);
and U5652 (N_5652,N_1062,N_1116);
or U5653 (N_5653,N_1713,N_1971);
or U5654 (N_5654,N_68,N_623);
xnor U5655 (N_5655,N_2317,N_2592);
or U5656 (N_5656,N_2889,N_2239);
nor U5657 (N_5657,N_1189,N_2352);
xnor U5658 (N_5658,N_2846,N_2849);
nand U5659 (N_5659,N_2434,N_1847);
or U5660 (N_5660,N_912,N_568);
and U5661 (N_5661,N_34,N_1696);
nor U5662 (N_5662,N_2092,N_1093);
or U5663 (N_5663,N_631,N_391);
or U5664 (N_5664,N_2892,N_1525);
or U5665 (N_5665,N_114,N_535);
xor U5666 (N_5666,N_2844,N_2251);
nand U5667 (N_5667,N_1465,N_2176);
nand U5668 (N_5668,N_2725,N_1620);
or U5669 (N_5669,N_1675,N_179);
nand U5670 (N_5670,N_1345,N_267);
and U5671 (N_5671,N_356,N_979);
nand U5672 (N_5672,N_530,N_1156);
xnor U5673 (N_5673,N_1246,N_187);
nand U5674 (N_5674,N_1239,N_845);
and U5675 (N_5675,N_1045,N_2115);
and U5676 (N_5676,N_882,N_1909);
xor U5677 (N_5677,N_777,N_100);
and U5678 (N_5678,N_2531,N_2093);
or U5679 (N_5679,N_1628,N_2536);
nor U5680 (N_5680,N_2966,N_2329);
and U5681 (N_5681,N_2153,N_1927);
xnor U5682 (N_5682,N_186,N_1796);
and U5683 (N_5683,N_2558,N_2591);
or U5684 (N_5684,N_1896,N_2711);
xor U5685 (N_5685,N_1735,N_1090);
xnor U5686 (N_5686,N_135,N_555);
nand U5687 (N_5687,N_2589,N_91);
or U5688 (N_5688,N_2870,N_2551);
nand U5689 (N_5689,N_2173,N_1210);
or U5690 (N_5690,N_2865,N_2518);
nor U5691 (N_5691,N_2579,N_917);
xnor U5692 (N_5692,N_342,N_1444);
nor U5693 (N_5693,N_1018,N_2633);
xor U5694 (N_5694,N_1297,N_2031);
and U5695 (N_5695,N_710,N_400);
or U5696 (N_5696,N_1607,N_688);
and U5697 (N_5697,N_852,N_1784);
and U5698 (N_5698,N_1816,N_96);
or U5699 (N_5699,N_486,N_2746);
nor U5700 (N_5700,N_602,N_574);
or U5701 (N_5701,N_1290,N_2960);
and U5702 (N_5702,N_2038,N_961);
nor U5703 (N_5703,N_1238,N_2394);
nor U5704 (N_5704,N_909,N_2140);
xor U5705 (N_5705,N_1515,N_1141);
and U5706 (N_5706,N_1163,N_579);
or U5707 (N_5707,N_1794,N_303);
nand U5708 (N_5708,N_1890,N_1882);
nand U5709 (N_5709,N_1970,N_1838);
xnor U5710 (N_5710,N_441,N_2311);
or U5711 (N_5711,N_2460,N_1827);
and U5712 (N_5712,N_2048,N_696);
nor U5713 (N_5713,N_1030,N_1195);
and U5714 (N_5714,N_571,N_2787);
xor U5715 (N_5715,N_640,N_2989);
or U5716 (N_5716,N_2301,N_1347);
or U5717 (N_5717,N_2886,N_1492);
nand U5718 (N_5718,N_2719,N_809);
or U5719 (N_5719,N_2344,N_2388);
xor U5720 (N_5720,N_1214,N_1094);
xor U5721 (N_5721,N_1929,N_748);
xor U5722 (N_5722,N_1866,N_1579);
nor U5723 (N_5723,N_2637,N_151);
xor U5724 (N_5724,N_1582,N_401);
nor U5725 (N_5725,N_400,N_2834);
nand U5726 (N_5726,N_2913,N_699);
nand U5727 (N_5727,N_136,N_2041);
nand U5728 (N_5728,N_1584,N_1895);
and U5729 (N_5729,N_103,N_732);
xnor U5730 (N_5730,N_2199,N_548);
nor U5731 (N_5731,N_296,N_1745);
xnor U5732 (N_5732,N_379,N_1289);
xnor U5733 (N_5733,N_1954,N_1792);
and U5734 (N_5734,N_55,N_2916);
and U5735 (N_5735,N_1391,N_1126);
nand U5736 (N_5736,N_1856,N_1760);
nor U5737 (N_5737,N_994,N_1304);
or U5738 (N_5738,N_972,N_2112);
or U5739 (N_5739,N_1769,N_288);
and U5740 (N_5740,N_2423,N_737);
or U5741 (N_5741,N_2900,N_1947);
nor U5742 (N_5742,N_1367,N_60);
and U5743 (N_5743,N_2358,N_1886);
nor U5744 (N_5744,N_1719,N_531);
xnor U5745 (N_5745,N_2894,N_2126);
and U5746 (N_5746,N_59,N_1485);
nor U5747 (N_5747,N_1671,N_749);
nand U5748 (N_5748,N_405,N_2785);
and U5749 (N_5749,N_1309,N_1196);
or U5750 (N_5750,N_2466,N_929);
nor U5751 (N_5751,N_2387,N_2326);
or U5752 (N_5752,N_1934,N_2547);
nand U5753 (N_5753,N_734,N_518);
and U5754 (N_5754,N_804,N_1858);
or U5755 (N_5755,N_677,N_852);
nand U5756 (N_5756,N_2703,N_1557);
and U5757 (N_5757,N_2982,N_1903);
nand U5758 (N_5758,N_2110,N_2802);
or U5759 (N_5759,N_1711,N_2244);
or U5760 (N_5760,N_2454,N_953);
nand U5761 (N_5761,N_2129,N_142);
nand U5762 (N_5762,N_1719,N_2681);
xor U5763 (N_5763,N_1705,N_468);
nor U5764 (N_5764,N_881,N_2776);
and U5765 (N_5765,N_1323,N_2983);
and U5766 (N_5766,N_1096,N_1691);
xnor U5767 (N_5767,N_1449,N_2344);
nand U5768 (N_5768,N_710,N_1);
nand U5769 (N_5769,N_1280,N_2205);
nor U5770 (N_5770,N_36,N_2014);
nand U5771 (N_5771,N_899,N_225);
nor U5772 (N_5772,N_2310,N_2431);
and U5773 (N_5773,N_1433,N_1030);
nor U5774 (N_5774,N_2880,N_1811);
or U5775 (N_5775,N_1080,N_535);
nand U5776 (N_5776,N_2310,N_1058);
or U5777 (N_5777,N_1912,N_934);
or U5778 (N_5778,N_1738,N_954);
and U5779 (N_5779,N_435,N_2821);
and U5780 (N_5780,N_997,N_1512);
xor U5781 (N_5781,N_1166,N_1047);
xnor U5782 (N_5782,N_2122,N_2046);
nor U5783 (N_5783,N_2516,N_853);
nor U5784 (N_5784,N_2102,N_2828);
xnor U5785 (N_5785,N_483,N_1805);
xnor U5786 (N_5786,N_559,N_2927);
nand U5787 (N_5787,N_632,N_8);
nor U5788 (N_5788,N_1307,N_2956);
xnor U5789 (N_5789,N_451,N_967);
or U5790 (N_5790,N_246,N_2536);
nand U5791 (N_5791,N_2729,N_2799);
or U5792 (N_5792,N_1711,N_329);
and U5793 (N_5793,N_369,N_1263);
or U5794 (N_5794,N_760,N_588);
nand U5795 (N_5795,N_28,N_816);
nand U5796 (N_5796,N_1289,N_1857);
xnor U5797 (N_5797,N_363,N_605);
nor U5798 (N_5798,N_2215,N_2524);
or U5799 (N_5799,N_2455,N_1500);
and U5800 (N_5800,N_1581,N_2232);
or U5801 (N_5801,N_1558,N_46);
nor U5802 (N_5802,N_757,N_2988);
nand U5803 (N_5803,N_1637,N_706);
or U5804 (N_5804,N_2423,N_648);
and U5805 (N_5805,N_634,N_2652);
xor U5806 (N_5806,N_791,N_2168);
nand U5807 (N_5807,N_808,N_643);
and U5808 (N_5808,N_2327,N_1048);
nand U5809 (N_5809,N_2066,N_1811);
or U5810 (N_5810,N_62,N_1937);
nor U5811 (N_5811,N_1149,N_722);
or U5812 (N_5812,N_1648,N_1608);
or U5813 (N_5813,N_1610,N_1655);
or U5814 (N_5814,N_2742,N_450);
and U5815 (N_5815,N_2365,N_783);
or U5816 (N_5816,N_2640,N_299);
and U5817 (N_5817,N_1677,N_2635);
and U5818 (N_5818,N_2876,N_1549);
and U5819 (N_5819,N_549,N_1512);
and U5820 (N_5820,N_2800,N_890);
nor U5821 (N_5821,N_1272,N_1553);
nand U5822 (N_5822,N_1302,N_160);
xnor U5823 (N_5823,N_2407,N_656);
and U5824 (N_5824,N_2017,N_558);
or U5825 (N_5825,N_1394,N_1872);
or U5826 (N_5826,N_983,N_731);
nor U5827 (N_5827,N_1297,N_220);
nor U5828 (N_5828,N_2237,N_1824);
nor U5829 (N_5829,N_2948,N_1125);
xor U5830 (N_5830,N_837,N_285);
and U5831 (N_5831,N_1551,N_2492);
xnor U5832 (N_5832,N_759,N_772);
and U5833 (N_5833,N_943,N_1677);
and U5834 (N_5834,N_1358,N_1887);
or U5835 (N_5835,N_1576,N_2615);
or U5836 (N_5836,N_423,N_1654);
nor U5837 (N_5837,N_1347,N_2023);
and U5838 (N_5838,N_1040,N_2748);
nor U5839 (N_5839,N_344,N_449);
and U5840 (N_5840,N_1844,N_2692);
xnor U5841 (N_5841,N_2670,N_431);
and U5842 (N_5842,N_823,N_1588);
nor U5843 (N_5843,N_1058,N_1277);
or U5844 (N_5844,N_2597,N_2949);
and U5845 (N_5845,N_2181,N_201);
or U5846 (N_5846,N_2469,N_228);
nor U5847 (N_5847,N_1169,N_2427);
or U5848 (N_5848,N_2447,N_458);
nor U5849 (N_5849,N_817,N_59);
nor U5850 (N_5850,N_1872,N_1515);
and U5851 (N_5851,N_12,N_1247);
xor U5852 (N_5852,N_870,N_1423);
nor U5853 (N_5853,N_738,N_1063);
or U5854 (N_5854,N_1413,N_121);
nand U5855 (N_5855,N_1282,N_1434);
nor U5856 (N_5856,N_117,N_425);
nor U5857 (N_5857,N_1297,N_576);
xor U5858 (N_5858,N_972,N_368);
xnor U5859 (N_5859,N_522,N_2186);
nor U5860 (N_5860,N_1060,N_353);
xor U5861 (N_5861,N_1185,N_560);
xor U5862 (N_5862,N_2320,N_1502);
xnor U5863 (N_5863,N_210,N_649);
xor U5864 (N_5864,N_2305,N_2764);
nor U5865 (N_5865,N_1953,N_1692);
and U5866 (N_5866,N_162,N_2009);
or U5867 (N_5867,N_1872,N_2481);
nor U5868 (N_5868,N_523,N_2081);
nor U5869 (N_5869,N_1270,N_200);
nor U5870 (N_5870,N_501,N_2962);
nor U5871 (N_5871,N_613,N_748);
or U5872 (N_5872,N_932,N_931);
or U5873 (N_5873,N_1335,N_543);
and U5874 (N_5874,N_2873,N_1957);
xnor U5875 (N_5875,N_2023,N_881);
xnor U5876 (N_5876,N_939,N_2779);
nor U5877 (N_5877,N_2177,N_410);
nor U5878 (N_5878,N_388,N_2695);
nand U5879 (N_5879,N_1290,N_763);
or U5880 (N_5880,N_884,N_10);
and U5881 (N_5881,N_1605,N_2386);
nand U5882 (N_5882,N_1111,N_2450);
or U5883 (N_5883,N_2692,N_1021);
nor U5884 (N_5884,N_1534,N_373);
nor U5885 (N_5885,N_1692,N_1482);
and U5886 (N_5886,N_1180,N_802);
or U5887 (N_5887,N_2450,N_408);
nor U5888 (N_5888,N_1643,N_2005);
or U5889 (N_5889,N_1297,N_1308);
xnor U5890 (N_5890,N_1627,N_2043);
nand U5891 (N_5891,N_412,N_1858);
nand U5892 (N_5892,N_114,N_622);
nand U5893 (N_5893,N_1040,N_204);
nand U5894 (N_5894,N_411,N_1767);
xnor U5895 (N_5895,N_432,N_1292);
and U5896 (N_5896,N_2943,N_2552);
nor U5897 (N_5897,N_1625,N_1464);
xor U5898 (N_5898,N_35,N_601);
xnor U5899 (N_5899,N_2998,N_1880);
and U5900 (N_5900,N_1598,N_2952);
nor U5901 (N_5901,N_1735,N_2771);
or U5902 (N_5902,N_544,N_671);
or U5903 (N_5903,N_1891,N_2943);
nor U5904 (N_5904,N_779,N_1164);
nand U5905 (N_5905,N_1267,N_2583);
or U5906 (N_5906,N_536,N_1750);
xor U5907 (N_5907,N_268,N_2807);
nand U5908 (N_5908,N_1739,N_1357);
and U5909 (N_5909,N_94,N_1932);
or U5910 (N_5910,N_664,N_2576);
nor U5911 (N_5911,N_409,N_1857);
or U5912 (N_5912,N_1589,N_513);
nand U5913 (N_5913,N_1913,N_2059);
nor U5914 (N_5914,N_1101,N_579);
nand U5915 (N_5915,N_1689,N_2998);
and U5916 (N_5916,N_2551,N_177);
and U5917 (N_5917,N_2964,N_1736);
xnor U5918 (N_5918,N_2656,N_2987);
or U5919 (N_5919,N_2387,N_1376);
or U5920 (N_5920,N_2225,N_930);
xor U5921 (N_5921,N_300,N_2455);
nor U5922 (N_5922,N_2257,N_634);
nand U5923 (N_5923,N_1628,N_593);
or U5924 (N_5924,N_2025,N_1130);
nor U5925 (N_5925,N_2097,N_1313);
and U5926 (N_5926,N_497,N_1391);
or U5927 (N_5927,N_1276,N_2322);
xnor U5928 (N_5928,N_1881,N_1145);
and U5929 (N_5929,N_854,N_1848);
nor U5930 (N_5930,N_884,N_1689);
xor U5931 (N_5931,N_1870,N_2620);
nor U5932 (N_5932,N_2755,N_16);
nand U5933 (N_5933,N_1318,N_2089);
and U5934 (N_5934,N_1999,N_1920);
nand U5935 (N_5935,N_2465,N_1510);
or U5936 (N_5936,N_2522,N_262);
xor U5937 (N_5937,N_265,N_260);
or U5938 (N_5938,N_2446,N_2471);
and U5939 (N_5939,N_2122,N_1473);
or U5940 (N_5940,N_841,N_638);
or U5941 (N_5941,N_1487,N_1647);
xor U5942 (N_5942,N_360,N_1233);
xor U5943 (N_5943,N_575,N_2913);
nor U5944 (N_5944,N_1077,N_696);
or U5945 (N_5945,N_1300,N_2112);
xnor U5946 (N_5946,N_1797,N_1834);
xnor U5947 (N_5947,N_2491,N_752);
or U5948 (N_5948,N_2207,N_655);
and U5949 (N_5949,N_2875,N_280);
and U5950 (N_5950,N_2432,N_176);
nor U5951 (N_5951,N_1799,N_526);
nor U5952 (N_5952,N_2029,N_426);
xor U5953 (N_5953,N_2011,N_1303);
xor U5954 (N_5954,N_760,N_616);
nor U5955 (N_5955,N_769,N_1609);
nand U5956 (N_5956,N_167,N_264);
and U5957 (N_5957,N_2955,N_1356);
nor U5958 (N_5958,N_271,N_1388);
or U5959 (N_5959,N_2829,N_773);
nand U5960 (N_5960,N_2982,N_132);
or U5961 (N_5961,N_2722,N_267);
nor U5962 (N_5962,N_2403,N_34);
nand U5963 (N_5963,N_1422,N_1915);
and U5964 (N_5964,N_788,N_603);
and U5965 (N_5965,N_2344,N_1193);
xnor U5966 (N_5966,N_1278,N_2227);
xnor U5967 (N_5967,N_1153,N_726);
and U5968 (N_5968,N_1536,N_1838);
or U5969 (N_5969,N_169,N_598);
nor U5970 (N_5970,N_660,N_2496);
xor U5971 (N_5971,N_1427,N_1553);
nor U5972 (N_5972,N_1495,N_2064);
nor U5973 (N_5973,N_996,N_179);
nand U5974 (N_5974,N_2076,N_1580);
xor U5975 (N_5975,N_500,N_2431);
nor U5976 (N_5976,N_1374,N_2734);
nand U5977 (N_5977,N_1210,N_408);
nand U5978 (N_5978,N_986,N_1906);
and U5979 (N_5979,N_1314,N_1306);
nor U5980 (N_5980,N_2321,N_66);
nand U5981 (N_5981,N_1572,N_1312);
nor U5982 (N_5982,N_1987,N_2050);
xnor U5983 (N_5983,N_2887,N_1266);
nand U5984 (N_5984,N_924,N_2482);
xor U5985 (N_5985,N_567,N_1714);
nor U5986 (N_5986,N_1781,N_2153);
xnor U5987 (N_5987,N_1942,N_35);
xor U5988 (N_5988,N_2236,N_254);
or U5989 (N_5989,N_2877,N_2551);
and U5990 (N_5990,N_1822,N_1234);
or U5991 (N_5991,N_1352,N_258);
nor U5992 (N_5992,N_2702,N_1030);
and U5993 (N_5993,N_1677,N_2343);
or U5994 (N_5994,N_281,N_2436);
nor U5995 (N_5995,N_987,N_795);
or U5996 (N_5996,N_2030,N_1976);
or U5997 (N_5997,N_1111,N_2923);
or U5998 (N_5998,N_842,N_343);
or U5999 (N_5999,N_853,N_2275);
nand U6000 (N_6000,N_3750,N_3777);
nand U6001 (N_6001,N_5993,N_5737);
xor U6002 (N_6002,N_5782,N_3797);
nand U6003 (N_6003,N_4664,N_5657);
and U6004 (N_6004,N_3746,N_5276);
nor U6005 (N_6005,N_5919,N_5923);
and U6006 (N_6006,N_5749,N_5365);
xnor U6007 (N_6007,N_3424,N_4108);
and U6008 (N_6008,N_5921,N_5128);
nand U6009 (N_6009,N_3780,N_5186);
nand U6010 (N_6010,N_3430,N_5174);
and U6011 (N_6011,N_4437,N_5475);
xnor U6012 (N_6012,N_5030,N_5658);
nor U6013 (N_6013,N_4005,N_3858);
and U6014 (N_6014,N_3158,N_5525);
or U6015 (N_6015,N_5953,N_3282);
or U6016 (N_6016,N_5252,N_3370);
or U6017 (N_6017,N_5383,N_3016);
and U6018 (N_6018,N_4349,N_4762);
or U6019 (N_6019,N_5247,N_5136);
xor U6020 (N_6020,N_3119,N_3264);
and U6021 (N_6021,N_5862,N_3725);
nand U6022 (N_6022,N_3206,N_3606);
and U6023 (N_6023,N_4298,N_4281);
xnor U6024 (N_6024,N_5514,N_3917);
xnor U6025 (N_6025,N_5499,N_3267);
or U6026 (N_6026,N_3703,N_4732);
xor U6027 (N_6027,N_3798,N_5332);
nor U6028 (N_6028,N_5971,N_5780);
or U6029 (N_6029,N_5967,N_3838);
nand U6030 (N_6030,N_3859,N_4378);
or U6031 (N_6031,N_4653,N_3031);
and U6032 (N_6032,N_5369,N_5717);
nor U6033 (N_6033,N_3680,N_4011);
nor U6034 (N_6034,N_3927,N_4561);
nand U6035 (N_6035,N_3566,N_3658);
xnor U6036 (N_6036,N_3467,N_3181);
or U6037 (N_6037,N_5185,N_5129);
nand U6038 (N_6038,N_4700,N_4498);
and U6039 (N_6039,N_3835,N_5445);
nand U6040 (N_6040,N_3591,N_5668);
xnor U6041 (N_6041,N_3537,N_5502);
or U6042 (N_6042,N_3716,N_3135);
or U6043 (N_6043,N_3827,N_5533);
or U6044 (N_6044,N_3749,N_3509);
and U6045 (N_6045,N_4646,N_5883);
nand U6046 (N_6046,N_5501,N_3241);
nand U6047 (N_6047,N_3333,N_5507);
nor U6048 (N_6048,N_3454,N_5856);
or U6049 (N_6049,N_4279,N_4450);
nor U6050 (N_6050,N_3253,N_3484);
or U6051 (N_6051,N_3695,N_3588);
nand U6052 (N_6052,N_3783,N_3775);
nand U6053 (N_6053,N_5567,N_3375);
and U6054 (N_6054,N_4726,N_4181);
nand U6055 (N_6055,N_5382,N_5672);
or U6056 (N_6056,N_3195,N_5891);
or U6057 (N_6057,N_3672,N_3573);
or U6058 (N_6058,N_3490,N_5178);
nand U6059 (N_6059,N_5064,N_4858);
nand U6060 (N_6060,N_4176,N_5554);
nand U6061 (N_6061,N_3882,N_5970);
xnor U6062 (N_6062,N_4363,N_3470);
nand U6063 (N_6063,N_5958,N_4409);
nor U6064 (N_6064,N_4477,N_5646);
nand U6065 (N_6065,N_3739,N_4737);
nand U6066 (N_6066,N_4185,N_5745);
or U6067 (N_6067,N_3022,N_5298);
nor U6068 (N_6068,N_4854,N_4074);
nand U6069 (N_6069,N_4585,N_3431);
and U6070 (N_6070,N_3975,N_4616);
and U6071 (N_6071,N_4900,N_5900);
nand U6072 (N_6072,N_4972,N_4875);
nand U6073 (N_6073,N_5860,N_5779);
nor U6074 (N_6074,N_5506,N_4420);
nand U6075 (N_6075,N_3069,N_4271);
nor U6076 (N_6076,N_5476,N_5652);
xor U6077 (N_6077,N_3621,N_5527);
or U6078 (N_6078,N_5463,N_4845);
xnor U6079 (N_6079,N_3203,N_4643);
and U6080 (N_6080,N_5297,N_5725);
nor U6081 (N_6081,N_4636,N_3209);
or U6082 (N_6082,N_5179,N_3717);
and U6083 (N_6083,N_3003,N_3698);
xnor U6084 (N_6084,N_3788,N_3929);
xor U6085 (N_6085,N_3021,N_4556);
nor U6086 (N_6086,N_4178,N_5778);
or U6087 (N_6087,N_3440,N_3543);
nor U6088 (N_6088,N_5182,N_3262);
or U6089 (N_6089,N_4496,N_4464);
or U6090 (N_6090,N_4621,N_5394);
nor U6091 (N_6091,N_5444,N_3968);
nor U6092 (N_6092,N_4177,N_5903);
xor U6093 (N_6093,N_5894,N_5569);
and U6094 (N_6094,N_5612,N_4567);
nor U6095 (N_6095,N_4473,N_4175);
or U6096 (N_6096,N_3937,N_3715);
or U6097 (N_6097,N_5158,N_3562);
xor U6098 (N_6098,N_5131,N_5884);
nor U6099 (N_6099,N_4043,N_4186);
or U6100 (N_6100,N_3026,N_3057);
xor U6101 (N_6101,N_5156,N_5774);
nor U6102 (N_6102,N_3930,N_5340);
and U6103 (N_6103,N_4961,N_3112);
nor U6104 (N_6104,N_4432,N_3417);
nor U6105 (N_6105,N_4276,N_4617);
nor U6106 (N_6106,N_3252,N_3995);
and U6107 (N_6107,N_3028,N_4256);
or U6108 (N_6108,N_3459,N_5814);
nor U6109 (N_6109,N_4428,N_4361);
and U6110 (N_6110,N_5270,N_3477);
xnor U6111 (N_6111,N_4038,N_4704);
xor U6112 (N_6112,N_4046,N_4358);
or U6113 (N_6113,N_5807,N_4212);
and U6114 (N_6114,N_4321,N_5283);
nor U6115 (N_6115,N_3906,N_4441);
or U6116 (N_6116,N_3125,N_3318);
or U6117 (N_6117,N_5052,N_4916);
nand U6118 (N_6118,N_3913,N_3399);
and U6119 (N_6119,N_5722,N_4575);
and U6120 (N_6120,N_5162,N_3527);
nor U6121 (N_6121,N_4215,N_3786);
and U6122 (N_6122,N_3974,N_5886);
xnor U6123 (N_6123,N_4828,N_5975);
xor U6124 (N_6124,N_5126,N_5102);
nor U6125 (N_6125,N_3166,N_5834);
and U6126 (N_6126,N_4397,N_5074);
xnor U6127 (N_6127,N_5763,N_3244);
or U6128 (N_6128,N_5543,N_4796);
or U6129 (N_6129,N_4105,N_3885);
and U6130 (N_6130,N_4752,N_3668);
or U6131 (N_6131,N_4385,N_4323);
or U6132 (N_6132,N_3579,N_3455);
nor U6133 (N_6133,N_3789,N_5644);
or U6134 (N_6134,N_5330,N_4093);
nor U6135 (N_6135,N_4873,N_4287);
nand U6136 (N_6136,N_5755,N_3067);
xor U6137 (N_6137,N_5107,N_3505);
and U6138 (N_6138,N_3380,N_5209);
and U6139 (N_6139,N_3912,N_4742);
or U6140 (N_6140,N_4334,N_5123);
nor U6141 (N_6141,N_4770,N_5704);
nand U6142 (N_6142,N_3321,N_3486);
and U6143 (N_6143,N_5248,N_5690);
xor U6144 (N_6144,N_5824,N_4656);
nand U6145 (N_6145,N_5464,N_4623);
nand U6146 (N_6146,N_4063,N_3952);
nand U6147 (N_6147,N_3903,N_4446);
or U6148 (N_6148,N_5676,N_3113);
or U6149 (N_6149,N_3934,N_3935);
nand U6150 (N_6150,N_3463,N_4172);
nor U6151 (N_6151,N_3977,N_5594);
and U6152 (N_6152,N_5944,N_3524);
xnor U6153 (N_6153,N_4896,N_4722);
and U6154 (N_6154,N_4768,N_5647);
and U6155 (N_6155,N_3785,N_3270);
nand U6156 (N_6156,N_3178,N_4891);
and U6157 (N_6157,N_3354,N_5399);
or U6158 (N_6158,N_3171,N_5998);
nand U6159 (N_6159,N_5603,N_3192);
and U6160 (N_6160,N_4760,N_3973);
or U6161 (N_6161,N_5733,N_3652);
xnor U6162 (N_6162,N_4535,N_5537);
and U6163 (N_6163,N_3612,N_3920);
nand U6164 (N_6164,N_4850,N_5304);
or U6165 (N_6165,N_3218,N_4200);
nor U6166 (N_6166,N_3950,N_3110);
nand U6167 (N_6167,N_5640,N_3081);
and U6168 (N_6168,N_3475,N_3724);
or U6169 (N_6169,N_4090,N_4534);
nand U6170 (N_6170,N_5928,N_3010);
or U6171 (N_6171,N_5593,N_5138);
or U6172 (N_6172,N_3711,N_4136);
or U6173 (N_6173,N_3767,N_4257);
or U6174 (N_6174,N_3942,N_4673);
nand U6175 (N_6175,N_5922,N_3465);
nand U6176 (N_6176,N_5563,N_4937);
and U6177 (N_6177,N_5380,N_4179);
xnor U6178 (N_6178,N_4784,N_3800);
nor U6179 (N_6179,N_3774,N_4309);
xnor U6180 (N_6180,N_5301,N_4982);
nand U6181 (N_6181,N_3522,N_5762);
xnor U6182 (N_6182,N_5326,N_5319);
or U6183 (N_6183,N_4746,N_4092);
and U6184 (N_6184,N_3288,N_4552);
or U6185 (N_6185,N_5266,N_4262);
and U6186 (N_6186,N_4343,N_5081);
and U6187 (N_6187,N_5582,N_3759);
xnor U6188 (N_6188,N_4702,N_3275);
nor U6189 (N_6189,N_4007,N_3544);
nor U6190 (N_6190,N_3024,N_5941);
and U6191 (N_6191,N_4774,N_3598);
nand U6192 (N_6192,N_4431,N_5237);
and U6193 (N_6193,N_3384,N_3994);
nand U6194 (N_6194,N_3329,N_5153);
or U6195 (N_6195,N_4275,N_4674);
nand U6196 (N_6196,N_5911,N_3602);
or U6197 (N_6197,N_3678,N_3681);
xor U6198 (N_6198,N_3837,N_3462);
nor U6199 (N_6199,N_5068,N_5288);
nor U6200 (N_6200,N_3418,N_3614);
xnor U6201 (N_6201,N_4675,N_5295);
nor U6202 (N_6202,N_5478,N_4138);
nand U6203 (N_6203,N_3271,N_3359);
nand U6204 (N_6204,N_3856,N_5187);
nand U6205 (N_6205,N_4439,N_4749);
xor U6206 (N_6206,N_3550,N_5936);
and U6207 (N_6207,N_3325,N_4504);
or U6208 (N_6208,N_4569,N_5830);
nand U6209 (N_6209,N_4268,N_5191);
nor U6210 (N_6210,N_4261,N_3823);
xnor U6211 (N_6211,N_3972,N_3266);
nand U6212 (N_6212,N_4015,N_5093);
or U6213 (N_6213,N_5265,N_5094);
and U6214 (N_6214,N_3029,N_4347);
nor U6215 (N_6215,N_3491,N_5157);
or U6216 (N_6216,N_5351,N_3223);
and U6217 (N_6217,N_4618,N_5566);
nand U6218 (N_6218,N_4506,N_3938);
or U6219 (N_6219,N_3768,N_4541);
nand U6220 (N_6220,N_4910,N_3033);
nand U6221 (N_6221,N_4427,N_4599);
nor U6222 (N_6222,N_4696,N_5318);
nor U6223 (N_6223,N_5665,N_5707);
xnor U6224 (N_6224,N_5151,N_3686);
or U6225 (N_6225,N_4307,N_4260);
nand U6226 (N_6226,N_5561,N_5576);
xor U6227 (N_6227,N_3257,N_4490);
xor U6228 (N_6228,N_4947,N_3915);
nor U6229 (N_6229,N_4255,N_3133);
nor U6230 (N_6230,N_3970,N_4786);
nor U6231 (N_6231,N_4503,N_5986);
xnor U6232 (N_6232,N_5496,N_3082);
nor U6233 (N_6233,N_5879,N_5255);
or U6234 (N_6234,N_3630,N_4229);
or U6235 (N_6235,N_5739,N_4266);
nor U6236 (N_6236,N_3956,N_3408);
or U6237 (N_6237,N_3613,N_5401);
or U6238 (N_6238,N_3758,N_5540);
nor U6239 (N_6239,N_5244,N_5144);
and U6240 (N_6240,N_3084,N_4830);
or U6241 (N_6241,N_3526,N_3852);
and U6242 (N_6242,N_3820,N_4035);
or U6243 (N_6243,N_3712,N_5504);
and U6244 (N_6244,N_5217,N_4151);
xor U6245 (N_6245,N_5435,N_3000);
and U6246 (N_6246,N_5724,N_3093);
nand U6247 (N_6247,N_4205,N_4198);
or U6248 (N_6248,N_3991,N_3908);
nor U6249 (N_6249,N_5979,N_4203);
nand U6250 (N_6250,N_5044,N_5654);
nand U6251 (N_6251,N_5536,N_3572);
or U6252 (N_6252,N_5099,N_5411);
nand U6253 (N_6253,N_5267,N_5379);
and U6254 (N_6254,N_5988,N_4750);
nor U6255 (N_6255,N_3762,N_3701);
and U6256 (N_6256,N_3626,N_4064);
nand U6257 (N_6257,N_5359,N_5441);
and U6258 (N_6258,N_4027,N_4348);
nand U6259 (N_6259,N_5345,N_4977);
nand U6260 (N_6260,N_4613,N_5173);
nand U6261 (N_6261,N_4544,N_4714);
nand U6262 (N_6262,N_4611,N_4848);
xnor U6263 (N_6263,N_5663,N_4707);
xnor U6264 (N_6264,N_3233,N_4153);
nand U6265 (N_6265,N_5368,N_5338);
or U6266 (N_6266,N_5405,N_3346);
nand U6267 (N_6267,N_3276,N_4282);
nand U6268 (N_6268,N_5089,N_3056);
xor U6269 (N_6269,N_4944,N_4115);
xor U6270 (N_6270,N_5494,N_4856);
nand U6271 (N_6271,N_3078,N_3434);
and U6272 (N_6272,N_5969,N_4157);
and U6273 (N_6273,N_3302,N_4512);
nor U6274 (N_6274,N_3374,N_3517);
nor U6275 (N_6275,N_3568,N_4975);
nor U6276 (N_6276,N_5296,N_4829);
xnor U6277 (N_6277,N_5788,N_4059);
and U6278 (N_6278,N_4332,N_5145);
xor U6279 (N_6279,N_5876,N_3412);
xor U6280 (N_6280,N_5051,N_4640);
and U6281 (N_6281,N_5920,N_5216);
nor U6282 (N_6282,N_5550,N_5208);
nand U6283 (N_6283,N_5624,N_3575);
nor U6284 (N_6284,N_5560,N_3261);
nand U6285 (N_6285,N_4487,N_5336);
nor U6286 (N_6286,N_4720,N_4016);
nor U6287 (N_6287,N_3175,N_4641);
or U6288 (N_6288,N_5959,N_3998);
nand U6289 (N_6289,N_3340,N_4839);
nand U6290 (N_6290,N_4558,N_4124);
xor U6291 (N_6291,N_3368,N_3848);
xor U6292 (N_6292,N_3707,N_3098);
xnor U6293 (N_6293,N_3255,N_5811);
nand U6294 (N_6294,N_5042,N_3733);
nor U6295 (N_6295,N_5512,N_3516);
xnor U6296 (N_6296,N_3087,N_4993);
nand U6297 (N_6297,N_4061,N_5034);
xnor U6298 (N_6298,N_3290,N_5135);
or U6299 (N_6299,N_4037,N_3729);
xor U6300 (N_6300,N_3202,N_3283);
and U6301 (N_6301,N_3892,N_5931);
nor U6302 (N_6302,N_3872,N_4422);
nor U6303 (N_6303,N_4773,N_5578);
or U6304 (N_6304,N_4394,N_4740);
nand U6305 (N_6305,N_5451,N_4531);
xnor U6306 (N_6306,N_3311,N_3895);
nand U6307 (N_6307,N_3458,N_4293);
and U6308 (N_6308,N_5628,N_3644);
xnor U6309 (N_6309,N_4958,N_5005);
xor U6310 (N_6310,N_5754,N_3461);
or U6311 (N_6311,N_3349,N_4497);
xnor U6312 (N_6312,N_4099,N_4761);
or U6313 (N_6313,N_5013,N_3336);
nor U6314 (N_6314,N_5987,N_5954);
xor U6315 (N_6315,N_3850,N_3460);
or U6316 (N_6316,N_5822,N_3179);
and U6317 (N_6317,N_5930,N_4793);
nand U6318 (N_6318,N_4912,N_3182);
nand U6319 (N_6319,N_4258,N_3273);
xnor U6320 (N_6320,N_5212,N_3803);
and U6321 (N_6321,N_4126,N_3291);
xor U6322 (N_6322,N_3577,N_4683);
or U6323 (N_6323,N_3249,N_5181);
nor U6324 (N_6324,N_5293,N_5282);
xor U6325 (N_6325,N_3664,N_3979);
and U6326 (N_6326,N_5027,N_5500);
and U6327 (N_6327,N_5025,N_4608);
xor U6328 (N_6328,N_5759,N_4973);
nand U6329 (N_6329,N_4026,N_3306);
and U6330 (N_6330,N_3445,N_3293);
nor U6331 (N_6331,N_5568,N_5992);
and U6332 (N_6332,N_3471,N_3685);
nor U6333 (N_6333,N_3190,N_5033);
or U6334 (N_6334,N_3294,N_4393);
nand U6335 (N_6335,N_3365,N_4083);
nand U6336 (N_6336,N_4204,N_3165);
nand U6337 (N_6337,N_3933,N_5870);
xor U6338 (N_6338,N_3634,N_4344);
or U6339 (N_6339,N_3594,N_4637);
nor U6340 (N_6340,N_3073,N_3511);
xnor U6341 (N_6341,N_3832,N_3450);
and U6342 (N_6342,N_3744,N_5564);
or U6343 (N_6343,N_5402,N_3221);
or U6344 (N_6344,N_5671,N_5610);
and U6345 (N_6345,N_4291,N_4501);
nor U6346 (N_6346,N_5516,N_3828);
nor U6347 (N_6347,N_5939,N_5080);
xor U6348 (N_6348,N_4933,N_3563);
nor U6349 (N_6349,N_5758,N_5542);
nand U6350 (N_6350,N_3435,N_5426);
nand U6351 (N_6351,N_3651,N_4491);
xnor U6352 (N_6352,N_3714,N_5466);
and U6353 (N_6353,N_4071,N_4076);
and U6354 (N_6354,N_5623,N_4466);
xor U6355 (N_6355,N_3694,N_4087);
nor U6356 (N_6356,N_5331,N_4406);
nand U6357 (N_6357,N_4580,N_4096);
xor U6358 (N_6358,N_5598,N_5448);
and U6359 (N_6359,N_5257,N_4008);
nor U6360 (N_6360,N_3008,N_3773);
and U6361 (N_6361,N_3414,N_4222);
nand U6362 (N_6362,N_5712,N_3530);
xnor U6363 (N_6363,N_5661,N_3231);
nor U6364 (N_6364,N_4816,N_4017);
nand U6365 (N_6365,N_4955,N_3019);
xor U6366 (N_6366,N_4967,N_4141);
xor U6367 (N_6367,N_4069,N_3388);
and U6368 (N_6368,N_4805,N_3383);
and U6369 (N_6369,N_4818,N_3600);
or U6370 (N_6370,N_5170,N_4474);
and U6371 (N_6371,N_4996,N_5125);
xnor U6372 (N_6372,N_5505,N_3020);
nand U6373 (N_6373,N_4607,N_5557);
or U6374 (N_6374,N_3831,N_3967);
or U6375 (N_6375,N_3628,N_5716);
nor U6376 (N_6376,N_5231,N_5750);
and U6377 (N_6377,N_5802,N_3951);
and U6378 (N_6378,N_5076,N_4926);
or U6379 (N_6379,N_4392,N_5087);
nand U6380 (N_6380,N_5881,N_3210);
and U6381 (N_6381,N_5680,N_5279);
or U6382 (N_6382,N_5997,N_3616);
or U6383 (N_6383,N_5146,N_4274);
and U6384 (N_6384,N_4682,N_4382);
or U6385 (N_6385,N_5510,N_5227);
xnor U6386 (N_6386,N_5434,N_4920);
nor U6387 (N_6387,N_5960,N_3839);
and U6388 (N_6388,N_4555,N_4002);
and U6389 (N_6389,N_4680,N_3319);
and U6390 (N_6390,N_5866,N_4615);
nor U6391 (N_6391,N_4359,N_3295);
and U6392 (N_6392,N_3204,N_4815);
nand U6393 (N_6393,N_5417,N_5458);
xnor U6394 (N_6394,N_5784,N_4187);
and U6395 (N_6395,N_4863,N_3313);
xnor U6396 (N_6396,N_4859,N_4666);
xor U6397 (N_6397,N_4218,N_4834);
xnor U6398 (N_6398,N_5357,N_4219);
and U6399 (N_6399,N_4907,N_5674);
or U6400 (N_6400,N_3234,N_5539);
and U6401 (N_6401,N_5271,N_3411);
and U6402 (N_6402,N_4368,N_4938);
nand U6403 (N_6403,N_4644,N_3999);
xor U6404 (N_6404,N_5343,N_3541);
xor U6405 (N_6405,N_5608,N_3143);
or U6406 (N_6406,N_5139,N_4190);
or U6407 (N_6407,N_3196,N_5120);
and U6408 (N_6408,N_5354,N_3356);
nor U6409 (N_6409,N_3809,N_3919);
nand U6410 (N_6410,N_3407,N_3617);
or U6411 (N_6411,N_4509,N_5078);
nor U6412 (N_6412,N_5946,N_3629);
and U6413 (N_6413,N_4651,N_4265);
or U6414 (N_6414,N_4073,N_3055);
xnor U6415 (N_6415,N_4983,N_3043);
or U6416 (N_6416,N_4542,N_5645);
and U6417 (N_6417,N_3801,N_3753);
xor U6418 (N_6418,N_4459,N_3960);
and U6419 (N_6419,N_3840,N_3259);
and U6420 (N_6420,N_4241,N_5022);
nand U6421 (N_6421,N_4711,N_3529);
or U6422 (N_6422,N_3647,N_4436);
nor U6423 (N_6423,N_3369,N_4870);
and U6424 (N_6424,N_4950,N_5334);
nand U6425 (N_6425,N_4117,N_3360);
nor U6426 (N_6426,N_4520,N_4905);
xor U6427 (N_6427,N_4857,N_4620);
xnor U6428 (N_6428,N_3147,N_5377);
xor U6429 (N_6429,N_5897,N_5703);
or U6430 (N_6430,N_5235,N_3921);
or U6431 (N_6431,N_4741,N_5233);
and U6432 (N_6432,N_5075,N_4012);
or U6433 (N_6433,N_5112,N_5934);
or U6434 (N_6434,N_3845,N_4080);
nor U6435 (N_6435,N_3317,N_3766);
and U6436 (N_6436,N_3362,N_4295);
nand U6437 (N_6437,N_5105,N_4744);
nor U6438 (N_6438,N_3954,N_3656);
xor U6439 (N_6439,N_4692,N_4192);
or U6440 (N_6440,N_5277,N_5698);
nor U6441 (N_6441,N_3492,N_5036);
nor U6442 (N_6442,N_3278,N_4244);
or U6443 (N_6443,N_3625,N_4990);
and U6444 (N_6444,N_3909,N_4954);
xnor U6445 (N_6445,N_3870,N_4051);
nor U6446 (N_6446,N_4039,N_4791);
nand U6447 (N_6447,N_4979,N_3274);
and U6448 (N_6448,N_3071,N_4988);
or U6449 (N_6449,N_3323,N_5721);
and U6450 (N_6450,N_4697,N_3141);
nand U6451 (N_6451,N_4871,N_4549);
or U6452 (N_6452,N_3833,N_5590);
xor U6453 (N_6453,N_5529,N_3565);
nor U6454 (N_6454,N_3401,N_4612);
nor U6455 (N_6455,N_4661,N_3500);
and U6456 (N_6456,N_4524,N_3756);
nor U6457 (N_6457,N_3654,N_5240);
xnor U6458 (N_6458,N_3394,N_3343);
nor U6459 (N_6459,N_3778,N_3790);
nand U6460 (N_6460,N_3889,N_5468);
nand U6461 (N_6461,N_5281,N_5307);
xnor U6462 (N_6462,N_4671,N_3692);
xnor U6463 (N_6463,N_3946,N_5771);
xnor U6464 (N_6464,N_4247,N_4718);
or U6465 (N_6465,N_3605,N_5898);
and U6466 (N_6466,N_3802,N_3199);
xnor U6467 (N_6467,N_4354,N_3727);
xnor U6468 (N_6468,N_5781,N_5404);
xnor U6469 (N_6469,N_5337,N_5692);
or U6470 (N_6470,N_5427,N_4047);
xnor U6471 (N_6471,N_4934,N_3564);
nand U6472 (N_6472,N_3873,N_3826);
and U6473 (N_6473,N_3704,N_3094);
nor U6474 (N_6474,N_4778,N_5290);
or U6475 (N_6475,N_3106,N_5858);
or U6476 (N_6476,N_5073,N_4230);
nor U6477 (N_6477,N_3219,N_3637);
nand U6478 (N_6478,N_3978,N_5333);
nor U6479 (N_6479,N_4594,N_3111);
nor U6480 (N_6480,N_5364,N_4438);
xor U6481 (N_6481,N_4029,N_5039);
or U6482 (N_6482,N_4862,N_3806);
nand U6483 (N_6483,N_4031,N_4688);
xnor U6484 (N_6484,N_4478,N_3497);
and U6485 (N_6485,N_4327,N_5804);
or U6486 (N_6486,N_5109,N_3552);
nor U6487 (N_6487,N_3339,N_5118);
xnor U6488 (N_6488,N_5026,N_3240);
xor U6489 (N_6489,N_4107,N_3145);
nand U6490 (N_6490,N_4943,N_3627);
or U6491 (N_6491,N_4018,N_3482);
nand U6492 (N_6492,N_4889,N_3367);
nor U6493 (N_6493,N_5308,N_5605);
or U6494 (N_6494,N_5278,N_4433);
and U6495 (N_6495,N_4654,N_3322);
or U6496 (N_6496,N_4925,N_5857);
nand U6497 (N_6497,N_4525,N_3398);
and U6498 (N_6498,N_5286,N_3229);
nor U6499 (N_6499,N_5189,N_4233);
nor U6500 (N_6500,N_4103,N_4122);
nand U6501 (N_6501,N_5601,N_4906);
nor U6502 (N_6502,N_5816,N_3897);
xnor U6503 (N_6503,N_5250,N_3693);
xnor U6504 (N_6504,N_4831,N_4162);
xnor U6505 (N_6505,N_5609,N_3796);
nor U6506 (N_6506,N_4553,N_4030);
and U6507 (N_6507,N_5890,N_5339);
and U6508 (N_6508,N_5432,N_5016);
or U6509 (N_6509,N_3597,N_4299);
xnor U6510 (N_6510,N_4060,N_3246);
xor U6511 (N_6511,N_4710,N_3580);
or U6512 (N_6512,N_3423,N_5362);
nor U6513 (N_6513,N_5061,N_5989);
xor U6514 (N_6514,N_4777,N_5453);
xnor U6515 (N_6515,N_4927,N_3854);
nand U6516 (N_6516,N_5965,N_4743);
and U6517 (N_6517,N_4170,N_3957);
nand U6518 (N_6518,N_3515,N_3393);
and U6519 (N_6519,N_3345,N_5655);
or U6520 (N_6520,N_3172,N_5764);
or U6521 (N_6521,N_3453,N_4475);
nor U6522 (N_6522,N_4984,N_3713);
or U6523 (N_6523,N_3574,N_5360);
nor U6524 (N_6524,N_5905,N_5159);
and U6525 (N_6525,N_4738,N_3121);
and U6526 (N_6526,N_5889,N_4649);
xnor U6527 (N_6527,N_5744,N_4263);
nor U6528 (N_6528,N_3162,N_5855);
xnor U6529 (N_6529,N_3129,N_3269);
or U6530 (N_6530,N_4224,N_4998);
nor U6531 (N_6531,N_3437,N_3761);
xnor U6532 (N_6532,N_5581,N_3225);
or U6533 (N_6533,N_5234,N_5648);
or U6534 (N_6534,N_4166,N_4540);
xor U6535 (N_6535,N_4689,N_4853);
and U6536 (N_6536,N_5373,N_4902);
and U6537 (N_6537,N_4284,N_3260);
nor U6538 (N_6538,N_3070,N_4981);
or U6539 (N_6539,N_4072,N_3409);
or U6540 (N_6540,N_5913,N_3256);
and U6541 (N_6541,N_3723,N_5116);
and U6542 (N_6542,N_3296,N_4855);
and U6543 (N_6543,N_3105,N_3478);
nor U6544 (N_6544,N_4267,N_3865);
xor U6545 (N_6545,N_3232,N_4285);
xor U6546 (N_6546,N_3097,N_3787);
nor U6547 (N_6547,N_5893,N_3242);
nand U6548 (N_6548,N_3151,N_5847);
and U6549 (N_6549,N_4333,N_3381);
xor U6550 (N_6550,N_3235,N_3396);
nor U6551 (N_6551,N_3277,N_4997);
or U6552 (N_6552,N_5768,N_5371);
nor U6553 (N_6553,N_4144,N_5400);
nor U6554 (N_6554,N_3485,N_4822);
nand U6555 (N_6555,N_3925,N_5571);
and U6556 (N_6556,N_5132,N_3188);
and U6557 (N_6557,N_4313,N_3546);
or U6558 (N_6558,N_5642,N_4619);
and U6559 (N_6559,N_3377,N_5794);
and U6560 (N_6560,N_4515,N_3142);
xor U6561 (N_6561,N_3551,N_5115);
xnor U6562 (N_6562,N_5455,N_5607);
nor U6563 (N_6563,N_5066,N_3997);
or U6564 (N_6564,N_5565,N_4301);
nor U6565 (N_6565,N_3305,N_3899);
or U6566 (N_6566,N_5192,N_5994);
or U6567 (N_6567,N_5752,N_4444);
xor U6568 (N_6568,N_5790,N_5710);
nor U6569 (N_6569,N_4754,N_4452);
or U6570 (N_6570,N_4604,N_3289);
xnor U6571 (N_6571,N_4706,N_4040);
nand U6572 (N_6572,N_4131,N_3085);
nand U6573 (N_6573,N_3441,N_5416);
or U6574 (N_6574,N_4451,N_4974);
and U6575 (N_6575,N_3320,N_3825);
nor U6576 (N_6576,N_5786,N_5896);
and U6577 (N_6577,N_5656,N_3054);
nor U6578 (N_6578,N_3018,N_4399);
nand U6579 (N_6579,N_4893,N_3631);
nand U6580 (N_6580,N_5361,N_3817);
xnor U6581 (N_6581,N_5808,N_5742);
and U6582 (N_6582,N_3444,N_5403);
or U6583 (N_6583,N_3357,N_3083);
xor U6584 (N_6584,N_5917,N_4365);
and U6585 (N_6585,N_5347,N_5580);
and U6586 (N_6586,N_3648,N_4457);
and U6587 (N_6587,N_4766,N_5161);
or U6588 (N_6588,N_5431,N_4118);
or U6589 (N_6589,N_4199,N_4339);
xor U6590 (N_6590,N_5682,N_3353);
nor U6591 (N_6591,N_5702,N_5981);
or U6592 (N_6592,N_5374,N_5264);
nand U6593 (N_6593,N_3567,N_3705);
xor U6594 (N_6594,N_3438,N_5517);
xnor U6595 (N_6595,N_3867,N_4603);
nor U6596 (N_6596,N_5638,N_3122);
nand U6597 (N_6597,N_3996,N_5760);
xor U6598 (N_6598,N_3883,N_5848);
and U6599 (N_6599,N_4976,N_3638);
or U6600 (N_6600,N_5439,N_4374);
xor U6601 (N_6601,N_5038,N_4331);
and U6602 (N_6602,N_4277,N_3023);
or U6603 (N_6603,N_5242,N_5910);
nor U6604 (N_6604,N_5526,N_3187);
and U6605 (N_6605,N_3312,N_4447);
or U6606 (N_6606,N_4724,N_4248);
or U6607 (N_6607,N_4573,N_5961);
nand U6608 (N_6608,N_4899,N_5035);
xor U6609 (N_6609,N_3428,N_3748);
or U6610 (N_6610,N_5222,N_3585);
nor U6611 (N_6611,N_4625,N_3507);
or U6612 (N_6612,N_3690,N_4771);
nor U6613 (N_6613,N_4201,N_4312);
nor U6614 (N_6614,N_3760,N_4196);
nand U6615 (N_6615,N_3035,N_3379);
xnor U6616 (N_6616,N_3843,N_4058);
and U6617 (N_6617,N_4208,N_4054);
and U6618 (N_6618,N_4191,N_3769);
or U6619 (N_6619,N_4662,N_3126);
and U6620 (N_6620,N_4111,N_4811);
nor U6621 (N_6621,N_5101,N_4813);
nor U6622 (N_6622,N_4160,N_4174);
or U6623 (N_6623,N_5221,N_5619);
nand U6624 (N_6624,N_5599,N_4290);
or U6625 (N_6625,N_5211,N_4171);
and U6626 (N_6626,N_4453,N_3072);
nand U6627 (N_6627,N_5835,N_5206);
or U6628 (N_6628,N_3108,N_3265);
nand U6629 (N_6629,N_5363,N_3646);
xor U6630 (N_6630,N_5425,N_3764);
or U6631 (N_6631,N_4079,N_5874);
nor U6632 (N_6632,N_5490,N_4865);
nor U6633 (N_6633,N_4242,N_5086);
nor U6634 (N_6634,N_4329,N_5552);
or U6635 (N_6635,N_4991,N_5714);
and U6636 (N_6636,N_4592,N_5167);
nand U6637 (N_6637,N_4147,N_4288);
xor U6638 (N_6638,N_3347,N_4837);
xnor U6639 (N_6639,N_3898,N_5544);
and U6640 (N_6640,N_5583,N_5632);
xor U6641 (N_6641,N_5480,N_5878);
and U6642 (N_6642,N_3689,N_3747);
xnor U6643 (N_6643,N_5538,N_4006);
or U6644 (N_6644,N_5367,N_3560);
and U6645 (N_6645,N_5829,N_3137);
nor U6646 (N_6646,N_4946,N_4253);
nor U6647 (N_6647,N_4657,N_3963);
or U6648 (N_6648,N_4532,N_5772);
nor U6649 (N_6649,N_4234,N_4598);
and U6650 (N_6650,N_4189,N_3197);
nor U6651 (N_6651,N_4519,N_4584);
or U6652 (N_6652,N_3609,N_3815);
xnor U6653 (N_6653,N_5701,N_4775);
and U6654 (N_6654,N_4250,N_4941);
or U6655 (N_6655,N_5513,N_5777);
and U6656 (N_6656,N_5324,N_3239);
xnor U6657 (N_6657,N_3706,N_3738);
nor U6658 (N_6658,N_4658,N_5767);
or U6659 (N_6659,N_3052,N_4765);
xnor U6660 (N_6660,N_3479,N_3593);
xor U6661 (N_6661,N_5549,N_4132);
xnor U6662 (N_6662,N_4799,N_5524);
or U6663 (N_6663,N_5108,N_5637);
nand U6664 (N_6664,N_4056,N_4089);
and U6665 (N_6665,N_4684,N_5684);
and U6666 (N_6666,N_4094,N_5643);
and U6667 (N_6667,N_3433,N_3037);
nand U6668 (N_6668,N_5957,N_4969);
and U6669 (N_6669,N_5868,N_4713);
or U6670 (N_6670,N_3861,N_4560);
nor U6671 (N_6671,N_4860,N_3062);
xor U6672 (N_6672,N_3120,N_5045);
nand U6673 (N_6673,N_3350,N_4352);
nor U6674 (N_6674,N_4316,N_4879);
xor U6675 (N_6675,N_5223,N_5292);
xor U6676 (N_6676,N_4479,N_3004);
or U6677 (N_6677,N_4463,N_3781);
xnor U6678 (N_6678,N_3510,N_3918);
nand U6679 (N_6679,N_3251,N_5828);
nor U6680 (N_6680,N_4470,N_4824);
nor U6681 (N_6681,N_5462,N_3669);
and U6682 (N_6682,N_3272,N_3948);
nor U6683 (N_6683,N_4578,N_5287);
or U6684 (N_6684,N_4426,N_3059);
and U6685 (N_6685,N_3096,N_3641);
and U6686 (N_6686,N_3822,N_3639);
and U6687 (N_6687,N_5412,N_5972);
nand U6688 (N_6688,N_4838,N_4819);
or U6689 (N_6689,N_5017,N_5523);
xnor U6690 (N_6690,N_3468,N_5812);
nand U6691 (N_6691,N_4465,N_5888);
xnor U6692 (N_6692,N_3160,N_3015);
or U6693 (N_6693,N_3080,N_3503);
nand U6694 (N_6694,N_4589,N_4717);
xor U6695 (N_6695,N_3115,N_3287);
or U6696 (N_6696,N_4728,N_5815);
and U6697 (N_6697,N_3599,N_5955);
nand U6698 (N_6698,N_4493,N_5924);
xnor U6699 (N_6699,N_5914,N_3534);
nor U6700 (N_6700,N_4894,N_4574);
and U6701 (N_6701,N_4134,N_5872);
or U6702 (N_6702,N_4401,N_5110);
xor U6703 (N_6703,N_3687,N_5050);
or U6704 (N_6704,N_5346,N_4053);
nand U6705 (N_6705,N_3540,N_3039);
nor U6706 (N_6706,N_3696,N_3213);
nor U6707 (N_6707,N_4486,N_3238);
nand U6708 (N_6708,N_4091,N_4237);
and U6709 (N_6709,N_5322,N_3653);
xnor U6710 (N_6710,N_3429,N_4476);
nand U6711 (N_6711,N_5335,N_5831);
or U6712 (N_6712,N_4404,N_5509);
nor U6713 (N_6713,N_5687,N_5681);
nand U6714 (N_6714,N_4395,N_4844);
xor U6715 (N_6715,N_4652,N_5428);
or U6716 (N_6716,N_4622,N_3215);
nand U6717 (N_6717,N_4715,N_5761);
and U6718 (N_6718,N_4596,N_3793);
xnor U6719 (N_6719,N_4808,N_5621);
nor U6720 (N_6720,N_4232,N_3857);
nand U6721 (N_6721,N_5948,N_5024);
nand U6722 (N_6722,N_5452,N_3871);
or U6723 (N_6723,N_5810,N_3508);
nor U6724 (N_6724,N_3812,N_4570);
nor U6725 (N_6725,N_3523,N_4514);
or U6726 (N_6726,N_3344,N_4482);
or U6727 (N_6727,N_4308,N_5636);
or U6728 (N_6728,N_5515,N_5918);
nand U6729 (N_6729,N_3887,N_3391);
or U6730 (N_6730,N_3940,N_4411);
and U6731 (N_6731,N_5691,N_4669);
xor U6732 (N_6732,N_5184,N_5356);
nor U6733 (N_6733,N_4795,N_4957);
nand U6734 (N_6734,N_4351,N_3068);
nand U6735 (N_6735,N_3807,N_5689);
nor U6736 (N_6736,N_4812,N_3326);
xnor U6737 (N_6737,N_3549,N_3358);
and U6738 (N_6738,N_5547,N_4782);
nor U6739 (N_6739,N_3177,N_5773);
xor U6740 (N_6740,N_5467,N_3144);
nor U6741 (N_6741,N_5572,N_5908);
nand U6742 (N_6742,N_5597,N_4787);
and U6743 (N_6743,N_3632,N_4959);
and U6744 (N_6744,N_5459,N_4082);
nand U6745 (N_6745,N_5111,N_4881);
nand U6746 (N_6746,N_3811,N_4690);
xnor U6747 (N_6747,N_3341,N_4121);
xor U6748 (N_6748,N_3752,N_3496);
or U6749 (N_6749,N_3114,N_5902);
nand U6750 (N_6750,N_4686,N_3012);
or U6751 (N_6751,N_5555,N_5747);
nand U6752 (N_6752,N_5633,N_5190);
nand U6753 (N_6753,N_4455,N_5349);
xor U6754 (N_6754,N_3436,N_3911);
xor U6755 (N_6755,N_5015,N_5454);
xor U6756 (N_6756,N_3426,N_5699);
or U6757 (N_6757,N_3456,N_4500);
nor U6758 (N_6758,N_5697,N_5203);
xnor U6759 (N_6759,N_5397,N_4207);
or U6760 (N_6760,N_5700,N_4897);
and U6761 (N_6761,N_4042,N_3299);
xnor U6762 (N_6762,N_4936,N_5826);
nor U6763 (N_6763,N_3134,N_3076);
or U6764 (N_6764,N_4694,N_3824);
nor U6765 (N_6765,N_3813,N_5096);
nor U6766 (N_6766,N_3164,N_3372);
xnor U6767 (N_6767,N_5312,N_4472);
nand U6768 (N_6768,N_3618,N_4693);
nand U6769 (N_6769,N_3844,N_5059);
nor U6770 (N_6770,N_5272,N_3136);
nand U6771 (N_6771,N_3237,N_5818);
nand U6772 (N_6772,N_3308,N_3732);
nand U6773 (N_6773,N_5009,N_5103);
nand U6774 (N_6774,N_4747,N_4507);
nor U6775 (N_6775,N_4919,N_5589);
nor U6776 (N_6776,N_4488,N_3064);
or U6777 (N_6777,N_3794,N_3371);
or U6778 (N_6778,N_3730,N_3006);
or U6779 (N_6779,N_4032,N_4730);
xnor U6780 (N_6780,N_5262,N_3559);
and U6781 (N_6781,N_5836,N_4045);
or U6782 (N_6782,N_5325,N_3487);
or U6783 (N_6783,N_5885,N_4371);
nand U6784 (N_6784,N_5031,N_5696);
nand U6785 (N_6785,N_5877,N_5775);
nand U6786 (N_6786,N_5303,N_3734);
xnor U6787 (N_6787,N_5229,N_5546);
or U6788 (N_6788,N_4642,N_5200);
nor U6789 (N_6789,N_4565,N_4769);
and U6790 (N_6790,N_5871,N_4235);
nor U6791 (N_6791,N_5302,N_4956);
nand U6792 (N_6792,N_3513,N_3584);
nand U6793 (N_6793,N_4370,N_3481);
or U6794 (N_6794,N_4759,N_3254);
or U6795 (N_6795,N_5489,N_5314);
xnor U6796 (N_6796,N_4214,N_4685);
or U6797 (N_6797,N_4025,N_5795);
nand U6798 (N_6798,N_5469,N_4877);
xor U6799 (N_6799,N_3818,N_5393);
or U6800 (N_6800,N_5556,N_4562);
nand U6801 (N_6801,N_5952,N_3611);
or U6802 (N_6802,N_5048,N_3720);
nor U6803 (N_6803,N_4878,N_4419);
xor U6804 (N_6804,N_4511,N_3902);
or U6805 (N_6805,N_4734,N_5825);
nor U6806 (N_6806,N_3124,N_3851);
nand U6807 (N_6807,N_4821,N_5757);
xor U6808 (N_6808,N_4876,N_3662);
or U6809 (N_6809,N_3555,N_5983);
and U6810 (N_6810,N_3860,N_4101);
nor U6811 (N_6811,N_3697,N_5586);
or U6812 (N_6812,N_5695,N_3765);
nand U6813 (N_6813,N_4273,N_4505);
nor U6814 (N_6814,N_4128,N_4135);
xnor U6815 (N_6815,N_5406,N_3446);
or U6816 (N_6816,N_5713,N_3091);
nand U6817 (N_6817,N_5062,N_4003);
and U6818 (N_6818,N_5321,N_4745);
nor U6819 (N_6819,N_3645,N_4341);
or U6820 (N_6820,N_3674,N_3180);
nor U6821 (N_6821,N_3532,N_5753);
and U6822 (N_6822,N_4629,N_5418);
nand U6823 (N_6823,N_3309,N_5508);
nand U6824 (N_6824,N_4792,N_3499);
nand U6825 (N_6825,N_4882,N_3866);
nor U6826 (N_6826,N_4086,N_3205);
xnor U6827 (N_6827,N_3303,N_4480);
nand U6828 (N_6828,N_5008,N_5999);
or U6829 (N_6829,N_4319,N_4336);
nor U6830 (N_6830,N_4659,N_5670);
nor U6831 (N_6831,N_4914,N_5029);
or U6832 (N_6832,N_3846,N_4156);
and U6833 (N_6833,N_5414,N_4676);
nand U6834 (N_6834,N_3556,N_4609);
xor U6835 (N_6835,N_3819,N_3622);
and U6836 (N_6836,N_4048,N_5968);
nor U6837 (N_6837,N_5328,N_5631);
or U6838 (N_6838,N_4922,N_4402);
xnor U6839 (N_6839,N_5820,N_3047);
or U6840 (N_6840,N_5092,N_4687);
and U6841 (N_6841,N_5320,N_4326);
nand U6842 (N_6842,N_3044,N_5708);
or U6843 (N_6843,N_5797,N_5348);
xor U6844 (N_6844,N_5591,N_5783);
nor U6845 (N_6845,N_3901,N_5875);
nand U6846 (N_6846,N_3214,N_4735);
and U6847 (N_6847,N_5018,N_4942);
and U6848 (N_6848,N_5491,N_4495);
nand U6849 (N_6849,N_3285,N_4469);
nand U6850 (N_6850,N_4415,N_5522);
and U6851 (N_6851,N_4545,N_3439);
nor U6852 (N_6852,N_3220,N_3884);
nand U6853 (N_6853,N_5766,N_5196);
or U6854 (N_6854,N_3677,N_4709);
and U6855 (N_6855,N_4648,N_4345);
nand U6856 (N_6856,N_5477,N_4065);
nand U6857 (N_6857,N_4161,N_5728);
and U6858 (N_6858,N_3161,N_3893);
nand U6859 (N_6859,N_3208,N_4167);
xor U6860 (N_6860,N_5933,N_3236);
or U6861 (N_6861,N_5669,N_5437);
nor U6862 (N_6862,N_4626,N_4753);
and U6863 (N_6863,N_3791,N_5904);
xor U6864 (N_6864,N_3335,N_3736);
nand U6865 (N_6865,N_3905,N_5892);
xor U6866 (N_6866,N_5573,N_5084);
and U6867 (N_6867,N_5869,N_5859);
or U6868 (N_6868,N_3331,N_5551);
nor U6869 (N_6869,N_5800,N_3587);
nor U6870 (N_6870,N_4112,N_5041);
and U6871 (N_6871,N_4194,N_3879);
xnor U6872 (N_6872,N_3660,N_3615);
or U6873 (N_6873,N_3663,N_5990);
nor U6874 (N_6874,N_4429,N_3949);
nor U6875 (N_6875,N_5424,N_3422);
xor U6876 (N_6876,N_5584,N_4842);
or U6877 (N_6877,N_4872,N_5641);
nor U6878 (N_6878,N_5629,N_4213);
xnor U6879 (N_6879,N_4240,N_4405);
nand U6880 (N_6880,N_4106,N_4909);
or U6881 (N_6881,N_4139,N_3667);
or U6882 (N_6882,N_4962,N_3604);
or U6883 (N_6883,N_5389,N_5218);
and U6884 (N_6884,N_5241,N_5863);
nor U6885 (N_6885,N_4994,N_3799);
or U6886 (N_6886,N_4013,N_5852);
or U6887 (N_6887,N_3966,N_5164);
xnor U6888 (N_6888,N_3965,N_4867);
nand U6889 (N_6889,N_5001,N_3980);
or U6890 (N_6890,N_4445,N_4931);
and U6891 (N_6891,N_4130,N_5943);
and U6892 (N_6892,N_4739,N_3910);
nand U6893 (N_6893,N_4989,N_5730);
nand U6894 (N_6894,N_5207,N_5152);
nand U6895 (N_6895,N_3874,N_5666);
xnor U6896 (N_6896,N_4183,N_3066);
and U6897 (N_6897,N_5995,N_5082);
and U6898 (N_6898,N_4547,N_5532);
nand U6899 (N_6899,N_3226,N_3065);
and U6900 (N_6900,N_4283,N_5077);
or U6901 (N_6901,N_5047,N_4297);
nor U6902 (N_6902,N_3168,N_3268);
xnor U6903 (N_6903,N_4462,N_4785);
xor U6904 (N_6904,N_3007,N_4953);
nand U6905 (N_6905,N_4986,N_5493);
nor U6906 (N_6906,N_5613,N_4550);
nand U6907 (N_6907,N_5246,N_4206);
nand U6908 (N_6908,N_5756,N_4987);
or U6909 (N_6909,N_5011,N_5043);
and U6910 (N_6910,N_4650,N_4968);
nand U6911 (N_6911,N_3581,N_4731);
nor U6912 (N_6912,N_5531,N_3061);
nor U6913 (N_6913,N_3476,N_4100);
xnor U6914 (N_6914,N_4537,N_5720);
xnor U6915 (N_6915,N_5067,N_5776);
nand U6916 (N_6916,N_5376,N_3876);
and U6917 (N_6917,N_3684,N_4606);
xnor U6918 (N_6918,N_4806,N_3636);
or U6919 (N_6919,N_3814,N_3842);
nor U6920 (N_6920,N_3366,N_5065);
xnor U6921 (N_6921,N_4369,N_4388);
or U6922 (N_6922,N_5901,N_3148);
xor U6923 (N_6923,N_3364,N_5664);
nand U6924 (N_6924,N_3034,N_5127);
nand U6925 (N_6925,N_3014,N_5150);
and U6926 (N_6926,N_3976,N_4751);
xnor U6927 (N_6927,N_5023,N_4081);
and U6928 (N_6928,N_3038,N_5440);
nand U6929 (N_6929,N_3964,N_4670);
nand U6930 (N_6930,N_5950,N_3880);
xor U6931 (N_6931,N_4435,N_3472);
nor U6932 (N_6932,N_4320,N_4803);
nor U6933 (N_6933,N_3156,N_5966);
nand U6934 (N_6934,N_5028,N_4418);
or U6935 (N_6935,N_4668,N_3452);
or U6936 (N_6936,N_4999,N_5137);
nor U6937 (N_6937,N_3709,N_4756);
and U6938 (N_6938,N_4846,N_5419);
nor U6939 (N_6939,N_5090,N_3971);
xnor U6940 (N_6940,N_3448,N_3387);
nor U6941 (N_6941,N_3578,N_5163);
nor U6942 (N_6942,N_5473,N_4062);
xor U6943 (N_6943,N_4951,N_4800);
xnor U6944 (N_6944,N_3425,N_3457);
nand U6945 (N_6945,N_5787,N_4407);
nand U6946 (N_6946,N_5626,N_4066);
or U6947 (N_6947,N_5442,N_5423);
nor U6948 (N_6948,N_5254,N_5938);
nor U6949 (N_6949,N_4930,N_4843);
or U6950 (N_6950,N_4430,N_5639);
and U6951 (N_6951,N_5726,N_4180);
nor U6952 (N_6952,N_5471,N_3228);
or U6953 (N_6953,N_5169,N_5932);
xnor U6954 (N_6954,N_5350,N_5600);
or U6955 (N_6955,N_4965,N_5269);
and U6956 (N_6956,N_4639,N_3017);
and U6957 (N_6957,N_4917,N_4471);
nand U6958 (N_6958,N_3217,N_3258);
nand U6959 (N_6959,N_4454,N_5195);
nand U6960 (N_6960,N_3708,N_4033);
or U6961 (N_6961,N_5188,N_4386);
or U6962 (N_6962,N_4725,N_3691);
nand U6963 (N_6963,N_4583,N_4034);
nand U6964 (N_6964,N_4067,N_3413);
and U6965 (N_6965,N_3488,N_4789);
nor U6966 (N_6966,N_3936,N_5675);
nor U6967 (N_6967,N_3623,N_5479);
xor U6968 (N_6968,N_3710,N_5706);
nor U6969 (N_6969,N_3506,N_3784);
nand U6970 (N_6970,N_4913,N_5789);
nand U6971 (N_6971,N_4755,N_3334);
xnor U6972 (N_6972,N_3128,N_3649);
xnor U6973 (N_6973,N_3466,N_3875);
nor U6974 (N_6974,N_3109,N_4403);
nand U6975 (N_6975,N_5770,N_4587);
xnor U6976 (N_6976,N_5355,N_4518);
or U6977 (N_6977,N_4695,N_4055);
xnor U6978 (N_6978,N_4373,N_3792);
nand U6979 (N_6979,N_4849,N_5678);
xor U6980 (N_6980,N_3742,N_5143);
or U6981 (N_6981,N_4460,N_3655);
or U6982 (N_6982,N_5095,N_3174);
xor U6983 (N_6983,N_4679,N_4217);
or U6984 (N_6984,N_4510,N_5650);
nor U6985 (N_6985,N_5677,N_5548);
nand U6986 (N_6986,N_4548,N_5980);
nor U6987 (N_6987,N_5765,N_4836);
and U6988 (N_6988,N_5446,N_3740);
nand U6989 (N_6989,N_4353,N_4226);
xor U6990 (N_6990,N_4239,N_3138);
or U6991 (N_6991,N_3077,N_3571);
or U6992 (N_6992,N_4952,N_4776);
nor U6993 (N_6993,N_5198,N_4057);
nor U6994 (N_6994,N_4315,N_3036);
nand U6995 (N_6995,N_5735,N_5106);
xor U6996 (N_6996,N_5072,N_3855);
nand U6997 (N_6997,N_3212,N_5488);
nor U6998 (N_6998,N_4527,N_3184);
nor U6999 (N_6999,N_5625,N_4380);
xnor U7000 (N_7000,N_3688,N_5003);
nand U7001 (N_7001,N_3200,N_4489);
nor U7002 (N_7002,N_4932,N_4424);
xnor U7003 (N_7003,N_3805,N_3728);
xor U7004 (N_7004,N_4494,N_5268);
or U7005 (N_7005,N_4150,N_5006);
nor U7006 (N_7006,N_5055,N_4579);
nand U7007 (N_7007,N_3103,N_5553);
and U7008 (N_7008,N_5991,N_5054);
and U7009 (N_7009,N_4384,N_5738);
xnor U7010 (N_7010,N_3107,N_4508);
and U7011 (N_7011,N_3619,N_5309);
nand U7012 (N_7012,N_3955,N_4159);
or U7013 (N_7013,N_5253,N_4523);
and U7014 (N_7014,N_5785,N_4554);
nor U7015 (N_7015,N_3836,N_3222);
or U7016 (N_7016,N_5915,N_4322);
and U7017 (N_7017,N_5149,N_4699);
and U7018 (N_7018,N_5104,N_5407);
or U7019 (N_7019,N_5792,N_4410);
xnor U7020 (N_7020,N_5521,N_5004);
and U7021 (N_7021,N_3853,N_4939);
xnor U7022 (N_7022,N_5134,N_3013);
nand U7023 (N_7023,N_5197,N_4278);
or U7024 (N_7024,N_5718,N_3045);
xnor U7025 (N_7025,N_3675,N_4929);
nor U7026 (N_7026,N_3421,N_5385);
or U7027 (N_7027,N_3608,N_4243);
or U7028 (N_7028,N_4884,N_3868);
nand U7029 (N_7029,N_4772,N_4851);
or U7030 (N_7030,N_3130,N_4663);
or U7031 (N_7031,N_5996,N_4387);
nor U7032 (N_7032,N_5220,N_3316);
nor U7033 (N_7033,N_4588,N_5585);
xnor U7034 (N_7034,N_3131,N_3504);
xor U7035 (N_7035,N_5854,N_5370);
xnor U7036 (N_7036,N_5342,N_3620);
nor U7037 (N_7037,N_3498,N_4633);
nand U7038 (N_7038,N_3570,N_5317);
and U7039 (N_7039,N_5088,N_4456);
nor U7040 (N_7040,N_3250,N_3159);
and U7041 (N_7041,N_4325,N_3351);
and U7042 (N_7042,N_3307,N_3985);
and U7043 (N_7043,N_4814,N_4024);
nand U7044 (N_7044,N_4992,N_3201);
xor U7045 (N_7045,N_3330,N_5387);
nor U7046 (N_7046,N_5060,N_5899);
xor U7047 (N_7047,N_4645,N_4097);
and U7048 (N_7048,N_5275,N_4605);
or U7049 (N_7049,N_5481,N_5398);
xor U7050 (N_7050,N_3040,N_3395);
xnor U7051 (N_7051,N_5937,N_3301);
nand U7052 (N_7052,N_5422,N_5746);
and U7053 (N_7053,N_3650,N_4978);
and U7054 (N_7054,N_5239,N_4667);
and U7055 (N_7055,N_5562,N_4543);
nand U7056 (N_7056,N_4362,N_4360);
and U7057 (N_7057,N_3643,N_3888);
nor U7058 (N_7058,N_3886,N_3743);
xor U7059 (N_7059,N_4908,N_4202);
and U7060 (N_7060,N_5263,N_4533);
nand U7061 (N_7061,N_5358,N_4140);
and U7062 (N_7062,N_4142,N_3001);
nand U7063 (N_7063,N_5201,N_4832);
xnor U7064 (N_7064,N_4330,N_4634);
or U7065 (N_7065,N_3890,N_3342);
nand U7066 (N_7066,N_4314,N_4492);
xor U7067 (N_7067,N_3771,N_4538);
or U7068 (N_7068,N_4238,N_4627);
nand U7069 (N_7069,N_4077,N_3869);
xor U7070 (N_7070,N_5942,N_5978);
and U7071 (N_7071,N_5723,N_3224);
nand U7072 (N_7072,N_4915,N_4835);
nor U7073 (N_7073,N_4483,N_5408);
nand U7074 (N_7074,N_4306,N_4346);
nand U7075 (N_7075,N_5511,N_5461);
nand U7076 (N_7076,N_5935,N_5956);
nor U7077 (N_7077,N_4182,N_3536);
nand U7078 (N_7078,N_3735,N_4337);
or U7079 (N_7079,N_5037,N_4148);
xor U7080 (N_7080,N_4557,N_3483);
nand U7081 (N_7081,N_3961,N_5731);
nor U7082 (N_7082,N_5839,N_3048);
nand U7083 (N_7083,N_5803,N_5410);
and U7084 (N_7084,N_4582,N_3447);
nand U7085 (N_7085,N_3092,N_3154);
xnor U7086 (N_7086,N_3442,N_5659);
nor U7087 (N_7087,N_3539,N_4600);
or U7088 (N_7088,N_3157,N_3558);
and U7089 (N_7089,N_4023,N_4416);
or U7090 (N_7090,N_5243,N_3194);
nand U7091 (N_7091,N_4158,N_4443);
nand U7092 (N_7092,N_5274,N_4516);
or U7093 (N_7093,N_5483,N_5313);
xor U7094 (N_7094,N_4169,N_5575);
nand U7095 (N_7095,N_3722,N_3419);
nor U7096 (N_7096,N_4109,N_3877);
and U7097 (N_7097,N_3060,N_3416);
xor U7098 (N_7098,N_4367,N_4197);
nor U7099 (N_7099,N_5492,N_5219);
nand U7100 (N_7100,N_4921,N_3327);
and U7101 (N_7101,N_4110,N_3495);
nand U7102 (N_7102,N_3596,N_4885);
nor U7103 (N_7103,N_3962,N_4528);
and U7104 (N_7104,N_3146,N_5160);
nor U7105 (N_7105,N_4586,N_3173);
or U7106 (N_7106,N_5117,N_4980);
nor U7107 (N_7107,N_4895,N_4366);
or U7108 (N_7108,N_3300,N_4923);
or U7109 (N_7109,N_3553,N_5947);
xnor U7110 (N_7110,N_5409,N_5819);
xnor U7111 (N_7111,N_3400,N_3404);
xor U7112 (N_7112,N_3216,N_5249);
nor U7113 (N_7113,N_5693,N_3169);
nand U7114 (N_7114,N_5559,N_4940);
xnor U7115 (N_7115,N_4289,N_4338);
and U7116 (N_7116,N_5443,N_4809);
xnor U7117 (N_7117,N_5940,N_5821);
nand U7118 (N_7118,N_3878,N_3263);
xor U7119 (N_7119,N_3198,N_3586);
and U7120 (N_7120,N_3700,N_5210);
xor U7121 (N_7121,N_5705,N_3002);
xnor U7122 (N_7122,N_3063,N_5230);
nor U7123 (N_7123,N_4892,N_5844);
nand U7124 (N_7124,N_3569,N_3464);
nand U7125 (N_7125,N_3731,N_4269);
and U7126 (N_7126,N_3443,N_4448);
nand U7127 (N_7127,N_5012,N_4521);
and U7128 (N_7128,N_3881,N_4155);
nor U7129 (N_7129,N_4798,N_4225);
and U7130 (N_7130,N_5113,N_3834);
nand U7131 (N_7131,N_4245,N_5497);
or U7132 (N_7132,N_4716,N_3958);
xor U7133 (N_7133,N_4184,N_4467);
nor U7134 (N_7134,N_4014,N_3589);
xnor U7135 (N_7135,N_4631,N_4566);
or U7136 (N_7136,N_5791,N_5316);
xnor U7137 (N_7137,N_4964,N_4381);
nor U7138 (N_7138,N_5864,N_5019);
xor U7139 (N_7139,N_5711,N_5806);
nand U7140 (N_7140,N_4231,N_3741);
xor U7141 (N_7141,N_5727,N_5294);
nand U7142 (N_7142,N_5977,N_4502);
nand U7143 (N_7143,N_3953,N_5436);
or U7144 (N_7144,N_3361,N_4292);
nor U7145 (N_7145,N_4678,N_3163);
xor U7146 (N_7146,N_5449,N_4810);
nor U7147 (N_7147,N_3610,N_3284);
xnor U7148 (N_7148,N_5388,N_4526);
and U7149 (N_7149,N_3348,N_5851);
nor U7150 (N_7150,N_3982,N_3922);
nand U7151 (N_7151,N_5202,N_4075);
xnor U7152 (N_7152,N_3332,N_4970);
or U7153 (N_7153,N_3779,N_3907);
nand U7154 (N_7154,N_4041,N_5183);
xor U7155 (N_7155,N_4044,N_5175);
or U7156 (N_7156,N_4723,N_4227);
nand U7157 (N_7157,N_4137,N_4068);
nand U7158 (N_7158,N_4701,N_5058);
nor U7159 (N_7159,N_4010,N_4904);
xnor U7160 (N_7160,N_3721,N_4396);
or U7161 (N_7161,N_5215,N_3102);
nor U7162 (N_7162,N_5740,N_3449);
nor U7163 (N_7163,N_5535,N_4272);
or U7164 (N_7164,N_3932,N_5395);
nand U7165 (N_7165,N_5519,N_5799);
xor U7166 (N_7166,N_4591,N_5390);
or U7167 (N_7167,N_4022,N_4841);
or U7168 (N_7168,N_4948,N_4529);
and U7169 (N_7169,N_4249,N_5114);
nand U7170 (N_7170,N_5238,N_3127);
or U7171 (N_7171,N_4223,N_4305);
xnor U7172 (N_7172,N_4389,N_3104);
and U7173 (N_7173,N_5155,N_5285);
and U7174 (N_7174,N_3501,N_3095);
nand U7175 (N_7175,N_5245,N_3150);
or U7176 (N_7176,N_5984,N_5384);
nand U7177 (N_7177,N_3385,N_3051);
nor U7178 (N_7178,N_4571,N_5622);
xor U7179 (N_7179,N_3337,N_5827);
or U7180 (N_7180,N_3751,N_5258);
and U7181 (N_7181,N_5865,N_4294);
nand U7182 (N_7182,N_4767,N_4729);
xor U7183 (N_7183,N_5833,N_4681);
xnor U7184 (N_7184,N_3027,N_3100);
nor U7185 (N_7185,N_3373,N_5194);
nand U7186 (N_7186,N_3896,N_5867);
and U7187 (N_7187,N_4049,N_3657);
nand U7188 (N_7188,N_5306,N_4807);
xor U7189 (N_7189,N_3451,N_4391);
and U7190 (N_7190,N_3041,N_5457);
xnor U7191 (N_7191,N_4708,N_4660);
and U7192 (N_7192,N_5311,N_4357);
and U7193 (N_7193,N_5873,N_3661);
or U7194 (N_7194,N_5056,N_4748);
or U7195 (N_7195,N_5817,N_4513);
nand U7196 (N_7196,N_4960,N_3382);
nor U7197 (N_7197,N_3770,N_4736);
nor U7198 (N_7198,N_3583,N_3405);
nor U7199 (N_7199,N_5945,N_3520);
xnor U7200 (N_7200,N_4861,N_4719);
nand U7201 (N_7201,N_4154,N_4481);
xnor U7202 (N_7202,N_5840,N_4085);
or U7203 (N_7203,N_4691,N_5142);
or U7204 (N_7204,N_3659,N_3590);
nand U7205 (N_7205,N_5130,N_4246);
nand U7206 (N_7206,N_3782,N_5344);
nor U7207 (N_7207,N_3230,N_4677);
and U7208 (N_7208,N_4340,N_4372);
and U7209 (N_7209,N_4009,N_5100);
or U7210 (N_7210,N_4318,N_5205);
xnor U7211 (N_7211,N_5694,N_3944);
and U7212 (N_7212,N_3519,N_3904);
xnor U7213 (N_7213,N_5651,N_5798);
nand U7214 (N_7214,N_4125,N_3576);
nand U7215 (N_7215,N_4098,N_5204);
and U7216 (N_7216,N_4209,N_4078);
nor U7217 (N_7217,N_5579,N_3410);
nand U7218 (N_7218,N_4423,N_4133);
nand U7219 (N_7219,N_5057,N_5261);
nand U7220 (N_7220,N_3086,N_3718);
or U7221 (N_7221,N_4577,N_3049);
or U7222 (N_7222,N_5224,N_3891);
nand U7223 (N_7223,N_4020,N_4781);
nand U7224 (N_7224,N_3679,N_5541);
nand U7225 (N_7225,N_4168,N_3554);
nor U7226 (N_7226,N_5140,N_4635);
or U7227 (N_7227,N_4304,N_4593);
or U7228 (N_7228,N_5683,N_3864);
or U7229 (N_7229,N_5040,N_4966);
nor U7230 (N_7230,N_4001,N_4342);
nand U7231 (N_7231,N_4887,N_4116);
or U7232 (N_7232,N_4442,N_3117);
xnor U7233 (N_7233,N_3227,N_5846);
nand U7234 (N_7234,N_3191,N_5420);
xor U7235 (N_7235,N_5251,N_5534);
nor U7236 (N_7236,N_4376,N_3328);
xor U7237 (N_7237,N_5225,N_3603);
and U7238 (N_7238,N_5378,N_5843);
nand U7239 (N_7239,N_3642,N_5046);
xor U7240 (N_7240,N_3011,N_5615);
or U7241 (N_7241,N_5520,N_4647);
nor U7242 (N_7242,N_5973,N_5310);
xor U7243 (N_7243,N_3829,N_3757);
xor U7244 (N_7244,N_5375,N_3582);
or U7245 (N_7245,N_5154,N_4146);
and U7246 (N_7246,N_5021,N_5121);
nor U7247 (N_7247,N_4804,N_3521);
nor U7248 (N_7248,N_5014,N_4601);
nand U7249 (N_7249,N_4840,N_5495);
nand U7250 (N_7250,N_4335,N_4779);
nand U7251 (N_7251,N_3640,N_3518);
xor U7252 (N_7252,N_5098,N_5259);
nor U7253 (N_7253,N_3601,N_4355);
or U7254 (N_7254,N_3841,N_5352);
and U7255 (N_7255,N_3183,N_5097);
and U7256 (N_7256,N_5032,N_3376);
nand U7257 (N_7257,N_5976,N_5805);
nand U7258 (N_7258,N_4576,N_5341);
nand U7259 (N_7259,N_5982,N_3981);
nand U7260 (N_7260,N_5649,N_5635);
or U7261 (N_7261,N_5391,N_4825);
or U7262 (N_7262,N_5686,N_5729);
nor U7263 (N_7263,N_3118,N_5653);
and U7264 (N_7264,N_5193,N_4252);
nor U7265 (N_7265,N_3538,N_3830);
or U7266 (N_7266,N_4398,N_3185);
and U7267 (N_7267,N_4780,N_3139);
and U7268 (N_7268,N_4356,N_5232);
xor U7269 (N_7269,N_3959,N_3849);
nand U7270 (N_7270,N_3099,N_3525);
and U7271 (N_7271,N_5213,N_5850);
nand U7272 (N_7272,N_4568,N_5472);
xor U7273 (N_7273,N_3248,N_4303);
or U7274 (N_7274,N_4390,N_3916);
nand U7275 (N_7275,N_5236,N_5574);
nor U7276 (N_7276,N_3514,N_3561);
nor U7277 (N_7277,N_4665,N_5743);
or U7278 (N_7278,N_3132,N_5122);
or U7279 (N_7279,N_3804,N_4727);
nor U7280 (N_7280,N_3474,N_5071);
and U7281 (N_7281,N_4945,N_4572);
nor U7282 (N_7282,N_3390,N_3155);
nor U7283 (N_7283,N_5837,N_3992);
nand U7284 (N_7284,N_3297,N_4536);
xnor U7285 (N_7285,N_5133,N_4864);
xnor U7286 (N_7286,N_4935,N_3315);
xor U7287 (N_7287,N_3863,N_3847);
nor U7288 (N_7288,N_3635,N_5063);
or U7289 (N_7289,N_3324,N_3378);
nor U7290 (N_7290,N_4383,N_4296);
nand U7291 (N_7291,N_5912,N_5484);
nand U7292 (N_7292,N_5214,N_4425);
and U7293 (N_7293,N_4417,N_5845);
xnor U7294 (N_7294,N_3531,N_4918);
nand U7295 (N_7295,N_4546,N_4236);
xor U7296 (N_7296,N_3355,N_4129);
nor U7297 (N_7297,N_4632,N_4949);
nand U7298 (N_7298,N_3984,N_3469);
and U7299 (N_7299,N_3494,N_4499);
and U7300 (N_7300,N_5177,N_3207);
and U7301 (N_7301,N_3298,N_3928);
nand U7302 (N_7302,N_4794,N_5715);
nor U7303 (N_7303,N_5172,N_5985);
xor U7304 (N_7304,N_3005,N_5882);
xor U7305 (N_7305,N_3512,N_4551);
nor U7306 (N_7306,N_5486,N_4826);
nor U7307 (N_7307,N_3914,N_4564);
xnor U7308 (N_7308,N_5381,N_4324);
nand U7309 (N_7309,N_5091,N_3772);
or U7310 (N_7310,N_3557,N_3862);
nor U7311 (N_7311,N_3900,N_4004);
nand U7312 (N_7312,N_5604,N_3665);
or U7313 (N_7313,N_4434,N_4421);
or U7314 (N_7314,N_4590,N_4120);
nor U7315 (N_7315,N_5570,N_4264);
nand U7316 (N_7316,N_5256,N_3502);
xnor U7317 (N_7317,N_4084,N_5429);
xnor U7318 (N_7318,N_3943,N_4328);
nand U7319 (N_7319,N_3719,N_5180);
nor U7320 (N_7320,N_5962,N_5558);
and U7321 (N_7321,N_4847,N_4300);
nor U7322 (N_7322,N_5853,N_3186);
or U7323 (N_7323,N_3699,N_4901);
or U7324 (N_7324,N_5530,N_3397);
and U7325 (N_7325,N_3988,N_5528);
nor U7326 (N_7326,N_4104,N_4852);
xnor U7327 (N_7327,N_4221,N_3247);
nor U7328 (N_7328,N_4216,N_4070);
and U7329 (N_7329,N_5002,N_5880);
nand U7330 (N_7330,N_3046,N_3633);
and U7331 (N_7331,N_4364,N_3280);
xnor U7332 (N_7332,N_4485,N_4705);
or U7333 (N_7333,N_5085,N_3683);
or U7334 (N_7334,N_3755,N_3432);
nand U7335 (N_7335,N_4375,N_3281);
nand U7336 (N_7336,N_4254,N_3211);
and U7337 (N_7337,N_3624,N_4123);
nor U7338 (N_7338,N_5450,N_4880);
xor U7339 (N_7339,N_3402,N_3671);
nor U7340 (N_7340,N_4883,N_5166);
nand U7341 (N_7341,N_3245,N_3987);
nand U7342 (N_7342,N_3042,N_3542);
and U7343 (N_7343,N_4377,N_4119);
nand U7344 (N_7344,N_5456,N_3149);
xor U7345 (N_7345,N_4757,N_5020);
and U7346 (N_7346,N_5679,N_5618);
nor U7347 (N_7347,N_3926,N_4672);
or U7348 (N_7348,N_3726,N_3545);
xnor U7349 (N_7349,N_3304,N_4703);
nor U7350 (N_7350,N_5000,N_4597);
and U7351 (N_7351,N_5577,N_3924);
xnor U7352 (N_7352,N_5260,N_3673);
nor U7353 (N_7353,N_4302,N_4286);
nand U7354 (N_7354,N_3030,N_4259);
nand U7355 (N_7355,N_4408,N_3403);
xor U7356 (N_7356,N_5291,N_4088);
nand U7357 (N_7357,N_5433,N_5887);
or U7358 (N_7358,N_5611,N_3535);
nand U7359 (N_7359,N_3025,N_5503);
nor U7360 (N_7360,N_4127,N_3279);
xor U7361 (N_7361,N_4414,N_4036);
or U7362 (N_7362,N_5280,N_3745);
and U7363 (N_7363,N_4164,N_3170);
and U7364 (N_7364,N_4280,N_5849);
xnor U7365 (N_7365,N_5895,N_5719);
xnor U7366 (N_7366,N_5660,N_3990);
nor U7367 (N_7367,N_4888,N_4440);
or U7368 (N_7368,N_5796,N_4251);
or U7369 (N_7369,N_4874,N_5353);
or U7370 (N_7370,N_3737,N_3592);
nand U7371 (N_7371,N_4050,N_4866);
nor U7372 (N_7372,N_5487,N_4413);
and U7373 (N_7373,N_5518,N_5620);
and U7374 (N_7374,N_4721,N_4820);
nor U7375 (N_7375,N_4468,N_3682);
nand U7376 (N_7376,N_3314,N_5300);
nand U7377 (N_7377,N_3009,N_3989);
and U7378 (N_7378,N_5430,N_4484);
and U7379 (N_7379,N_5732,N_3406);
xor U7380 (N_7380,N_5284,N_5736);
xor U7381 (N_7381,N_3821,N_3116);
and U7382 (N_7382,N_4102,N_5470);
and U7383 (N_7383,N_5438,N_4581);
nand U7384 (N_7384,N_3363,N_5662);
or U7385 (N_7385,N_5832,N_5176);
nor U7386 (N_7386,N_4113,N_5329);
nand U7387 (N_7387,N_5305,N_3493);
nor U7388 (N_7388,N_5916,N_5396);
xor U7389 (N_7389,N_4028,N_5949);
or U7390 (N_7390,N_4802,N_3776);
nand U7391 (N_7391,N_4152,N_5685);
xnor U7392 (N_7392,N_4698,N_5734);
and U7393 (N_7393,N_4610,N_5465);
or U7394 (N_7394,N_5485,N_5751);
xnor U7395 (N_7395,N_3140,N_4911);
xnor U7396 (N_7396,N_5323,N_3352);
and U7397 (N_7397,N_5083,N_3189);
or U7398 (N_7398,N_3123,N_4317);
nand U7399 (N_7399,N_3810,N_5974);
and U7400 (N_7400,N_3931,N_4559);
or U7401 (N_7401,N_4995,N_4114);
nor U7402 (N_7402,N_4971,N_3153);
nor U7403 (N_7403,N_5327,N_5793);
nor U7404 (N_7404,N_5053,N_5299);
or U7405 (N_7405,N_5630,N_3547);
and U7406 (N_7406,N_5165,N_3089);
or U7407 (N_7407,N_3939,N_3941);
nand U7408 (N_7408,N_4019,N_4461);
nor U7409 (N_7409,N_4868,N_4458);
nor U7410 (N_7410,N_4655,N_3415);
xnor U7411 (N_7411,N_5124,N_4052);
or U7412 (N_7412,N_4733,N_3894);
nand U7413 (N_7413,N_3053,N_3595);
and U7414 (N_7414,N_3754,N_5315);
nor U7415 (N_7415,N_5606,N_5141);
nand U7416 (N_7416,N_5906,N_4783);
nand U7417 (N_7417,N_3338,N_3243);
nand U7418 (N_7418,N_4614,N_3079);
nand U7419 (N_7419,N_4095,N_4890);
nor U7420 (N_7420,N_3528,N_3480);
xnor U7421 (N_7421,N_3763,N_5049);
or U7422 (N_7422,N_5809,N_5010);
and U7423 (N_7423,N_3702,N_4624);
nand U7424 (N_7424,N_5171,N_3993);
or U7425 (N_7425,N_5007,N_4165);
nand U7426 (N_7426,N_3292,N_4143);
nand U7427 (N_7427,N_4595,N_3816);
nor U7428 (N_7428,N_5069,N_4400);
and U7429 (N_7429,N_4539,N_4000);
nand U7430 (N_7430,N_4758,N_4220);
nand U7431 (N_7431,N_5627,N_5616);
xor U7432 (N_7432,N_5907,N_5148);
or U7433 (N_7433,N_4563,N_5841);
nand U7434 (N_7434,N_5614,N_4801);
and U7435 (N_7435,N_3386,N_4228);
xor U7436 (N_7436,N_5801,N_4379);
nor U7437 (N_7437,N_3670,N_3607);
xnor U7438 (N_7438,N_3050,N_4193);
nand U7439 (N_7439,N_4963,N_4788);
and U7440 (N_7440,N_5634,N_5366);
or U7441 (N_7441,N_4712,N_5447);
xnor U7442 (N_7442,N_5813,N_5748);
or U7443 (N_7443,N_5587,N_5460);
and U7444 (N_7444,N_3489,N_5199);
or U7445 (N_7445,N_4311,N_5929);
nor U7446 (N_7446,N_3923,N_3075);
nor U7447 (N_7447,N_3427,N_3969);
nand U7448 (N_7448,N_5228,N_5421);
or U7449 (N_7449,N_4145,N_5842);
nand U7450 (N_7450,N_4021,N_4602);
nor U7451 (N_7451,N_5963,N_4310);
xnor U7452 (N_7452,N_4903,N_4638);
nor U7453 (N_7453,N_5741,N_5119);
nand U7454 (N_7454,N_5147,N_3090);
or U7455 (N_7455,N_4797,N_3983);
nand U7456 (N_7456,N_3088,N_3193);
and U7457 (N_7457,N_4928,N_5595);
or U7458 (N_7458,N_4790,N_3058);
nand U7459 (N_7459,N_5386,N_5498);
nor U7460 (N_7460,N_4149,N_4163);
nor U7461 (N_7461,N_3420,N_5070);
nor U7462 (N_7462,N_3808,N_3310);
nor U7463 (N_7463,N_3947,N_5926);
nor U7464 (N_7464,N_5588,N_3101);
nand U7465 (N_7465,N_4173,N_4270);
and U7466 (N_7466,N_5673,N_5226);
xnor U7467 (N_7467,N_5415,N_5823);
and U7468 (N_7468,N_4898,N_3986);
nand U7469 (N_7469,N_4630,N_5709);
xnor U7470 (N_7470,N_3548,N_5168);
or U7471 (N_7471,N_4869,N_4188);
or U7472 (N_7472,N_5769,N_4985);
xor U7473 (N_7473,N_4763,N_3795);
and U7474 (N_7474,N_5927,N_4924);
xor U7475 (N_7475,N_3176,N_5289);
or U7476 (N_7476,N_3032,N_4823);
xor U7477 (N_7477,N_5602,N_3676);
and U7478 (N_7478,N_5964,N_4522);
and U7479 (N_7479,N_4195,N_5925);
and U7480 (N_7480,N_5482,N_5079);
nor U7481 (N_7481,N_3533,N_3286);
nand U7482 (N_7482,N_5372,N_3473);
nor U7483 (N_7483,N_3392,N_5667);
nor U7484 (N_7484,N_4817,N_4517);
nand U7485 (N_7485,N_4350,N_5545);
nor U7486 (N_7486,N_4628,N_3389);
nand U7487 (N_7487,N_3666,N_4886);
nor U7488 (N_7488,N_4827,N_4412);
and U7489 (N_7489,N_3167,N_5617);
or U7490 (N_7490,N_4833,N_5592);
and U7491 (N_7491,N_4211,N_5909);
nor U7492 (N_7492,N_3152,N_5413);
or U7493 (N_7493,N_5951,N_4530);
xnor U7494 (N_7494,N_5273,N_4764);
and U7495 (N_7495,N_3074,N_5596);
xnor U7496 (N_7496,N_5838,N_5688);
or U7497 (N_7497,N_4210,N_5861);
nand U7498 (N_7498,N_5392,N_4449);
nand U7499 (N_7499,N_5474,N_3945);
xor U7500 (N_7500,N_5966,N_5717);
or U7501 (N_7501,N_5405,N_5221);
xor U7502 (N_7502,N_4673,N_5533);
xor U7503 (N_7503,N_5574,N_5381);
or U7504 (N_7504,N_5129,N_5881);
and U7505 (N_7505,N_3644,N_4246);
nor U7506 (N_7506,N_4269,N_4773);
and U7507 (N_7507,N_4373,N_3333);
nand U7508 (N_7508,N_3580,N_3138);
xnor U7509 (N_7509,N_4476,N_3309);
or U7510 (N_7510,N_3675,N_4603);
or U7511 (N_7511,N_3739,N_5458);
xor U7512 (N_7512,N_3384,N_4008);
nand U7513 (N_7513,N_4971,N_3505);
and U7514 (N_7514,N_5285,N_4442);
and U7515 (N_7515,N_5877,N_5037);
nor U7516 (N_7516,N_3830,N_5847);
xor U7517 (N_7517,N_5888,N_4652);
or U7518 (N_7518,N_5317,N_3179);
and U7519 (N_7519,N_3869,N_3379);
or U7520 (N_7520,N_4468,N_5979);
and U7521 (N_7521,N_4453,N_5399);
nand U7522 (N_7522,N_4219,N_5099);
or U7523 (N_7523,N_5405,N_4617);
nor U7524 (N_7524,N_3139,N_5690);
nor U7525 (N_7525,N_3237,N_3490);
nand U7526 (N_7526,N_3019,N_3202);
and U7527 (N_7527,N_4727,N_5529);
and U7528 (N_7528,N_5134,N_3456);
or U7529 (N_7529,N_4636,N_5891);
and U7530 (N_7530,N_5060,N_5081);
xnor U7531 (N_7531,N_3669,N_3243);
and U7532 (N_7532,N_4127,N_4024);
and U7533 (N_7533,N_4523,N_4315);
nor U7534 (N_7534,N_4598,N_3065);
or U7535 (N_7535,N_3429,N_4321);
nor U7536 (N_7536,N_4087,N_5959);
and U7537 (N_7537,N_5296,N_3052);
nor U7538 (N_7538,N_3899,N_3527);
nor U7539 (N_7539,N_4131,N_3357);
xnor U7540 (N_7540,N_4090,N_4432);
and U7541 (N_7541,N_3494,N_3985);
xor U7542 (N_7542,N_4063,N_5753);
xor U7543 (N_7543,N_3489,N_5165);
nor U7544 (N_7544,N_4802,N_4535);
xor U7545 (N_7545,N_4119,N_3011);
nor U7546 (N_7546,N_5858,N_3679);
nor U7547 (N_7547,N_3505,N_5951);
or U7548 (N_7548,N_3656,N_5808);
nand U7549 (N_7549,N_3045,N_3587);
or U7550 (N_7550,N_5723,N_3143);
or U7551 (N_7551,N_4535,N_5532);
nor U7552 (N_7552,N_5385,N_3617);
nand U7553 (N_7553,N_5424,N_3091);
xor U7554 (N_7554,N_4508,N_4707);
or U7555 (N_7555,N_4412,N_5531);
xnor U7556 (N_7556,N_5314,N_3974);
and U7557 (N_7557,N_4639,N_3872);
and U7558 (N_7558,N_5998,N_3709);
nor U7559 (N_7559,N_4254,N_5560);
or U7560 (N_7560,N_4957,N_3610);
xor U7561 (N_7561,N_3583,N_4738);
and U7562 (N_7562,N_4451,N_3735);
nor U7563 (N_7563,N_3690,N_4429);
or U7564 (N_7564,N_4598,N_4276);
or U7565 (N_7565,N_3320,N_5337);
and U7566 (N_7566,N_4224,N_3925);
xnor U7567 (N_7567,N_5663,N_3324);
nor U7568 (N_7568,N_4272,N_4437);
xor U7569 (N_7569,N_4912,N_3153);
and U7570 (N_7570,N_3578,N_5434);
nor U7571 (N_7571,N_3407,N_4939);
or U7572 (N_7572,N_5173,N_5836);
nand U7573 (N_7573,N_3825,N_3806);
nand U7574 (N_7574,N_4481,N_4045);
and U7575 (N_7575,N_4908,N_4824);
nand U7576 (N_7576,N_3554,N_3731);
or U7577 (N_7577,N_4321,N_3865);
and U7578 (N_7578,N_5359,N_4021);
or U7579 (N_7579,N_4281,N_5730);
or U7580 (N_7580,N_3074,N_4059);
xor U7581 (N_7581,N_5636,N_4543);
or U7582 (N_7582,N_5342,N_5891);
or U7583 (N_7583,N_4592,N_3960);
or U7584 (N_7584,N_5973,N_5530);
xor U7585 (N_7585,N_4836,N_5508);
xor U7586 (N_7586,N_3662,N_4683);
and U7587 (N_7587,N_5980,N_4974);
or U7588 (N_7588,N_3319,N_4801);
nor U7589 (N_7589,N_4779,N_3826);
nor U7590 (N_7590,N_5798,N_4042);
or U7591 (N_7591,N_4134,N_5335);
nand U7592 (N_7592,N_5307,N_4128);
xnor U7593 (N_7593,N_3910,N_3932);
and U7594 (N_7594,N_5629,N_4250);
nand U7595 (N_7595,N_4798,N_5518);
xor U7596 (N_7596,N_4589,N_5141);
or U7597 (N_7597,N_5438,N_4708);
nand U7598 (N_7598,N_4883,N_5102);
or U7599 (N_7599,N_5559,N_5946);
or U7600 (N_7600,N_4029,N_3396);
nor U7601 (N_7601,N_4075,N_4396);
or U7602 (N_7602,N_4755,N_3457);
nand U7603 (N_7603,N_3654,N_4825);
and U7604 (N_7604,N_4901,N_3289);
or U7605 (N_7605,N_3234,N_4891);
xnor U7606 (N_7606,N_3416,N_5187);
nor U7607 (N_7607,N_3830,N_4186);
xnor U7608 (N_7608,N_4891,N_3479);
nand U7609 (N_7609,N_3376,N_3295);
xnor U7610 (N_7610,N_5378,N_3329);
or U7611 (N_7611,N_5690,N_4149);
or U7612 (N_7612,N_3110,N_3091);
xor U7613 (N_7613,N_3402,N_3946);
or U7614 (N_7614,N_5329,N_4617);
nand U7615 (N_7615,N_5007,N_3929);
nand U7616 (N_7616,N_3560,N_5679);
nand U7617 (N_7617,N_4960,N_4558);
nand U7618 (N_7618,N_3111,N_4304);
nor U7619 (N_7619,N_3627,N_5948);
xnor U7620 (N_7620,N_3255,N_5873);
or U7621 (N_7621,N_4490,N_5111);
and U7622 (N_7622,N_5087,N_3765);
nand U7623 (N_7623,N_3678,N_5581);
xor U7624 (N_7624,N_4966,N_3232);
xor U7625 (N_7625,N_4370,N_5003);
xor U7626 (N_7626,N_4262,N_4550);
or U7627 (N_7627,N_4269,N_4091);
xnor U7628 (N_7628,N_5092,N_5336);
xor U7629 (N_7629,N_5610,N_3198);
nor U7630 (N_7630,N_3361,N_4876);
and U7631 (N_7631,N_5849,N_4261);
xor U7632 (N_7632,N_3485,N_4211);
or U7633 (N_7633,N_5490,N_4554);
nor U7634 (N_7634,N_4150,N_3068);
xnor U7635 (N_7635,N_3905,N_3591);
nand U7636 (N_7636,N_5921,N_5929);
nand U7637 (N_7637,N_3856,N_3297);
and U7638 (N_7638,N_5043,N_3969);
xor U7639 (N_7639,N_3097,N_3889);
xnor U7640 (N_7640,N_5279,N_4379);
or U7641 (N_7641,N_5324,N_4725);
or U7642 (N_7642,N_3168,N_3721);
nand U7643 (N_7643,N_4070,N_5369);
nor U7644 (N_7644,N_4200,N_3290);
xor U7645 (N_7645,N_5392,N_4895);
nand U7646 (N_7646,N_5325,N_3186);
nand U7647 (N_7647,N_5208,N_3924);
nor U7648 (N_7648,N_5701,N_3242);
and U7649 (N_7649,N_3772,N_3915);
and U7650 (N_7650,N_5375,N_4045);
nand U7651 (N_7651,N_5638,N_3503);
nand U7652 (N_7652,N_5874,N_4429);
or U7653 (N_7653,N_5366,N_5395);
and U7654 (N_7654,N_5884,N_3393);
xnor U7655 (N_7655,N_5938,N_3750);
or U7656 (N_7656,N_5306,N_5901);
nor U7657 (N_7657,N_3133,N_4924);
nand U7658 (N_7658,N_4282,N_5705);
or U7659 (N_7659,N_3211,N_4740);
or U7660 (N_7660,N_5608,N_5319);
nand U7661 (N_7661,N_4576,N_4739);
nand U7662 (N_7662,N_4063,N_4822);
nor U7663 (N_7663,N_4538,N_3277);
and U7664 (N_7664,N_5322,N_3608);
xnor U7665 (N_7665,N_5696,N_5827);
and U7666 (N_7666,N_3793,N_4765);
xnor U7667 (N_7667,N_3502,N_4581);
or U7668 (N_7668,N_3044,N_3323);
and U7669 (N_7669,N_4959,N_4659);
or U7670 (N_7670,N_3636,N_4894);
nor U7671 (N_7671,N_4254,N_5482);
and U7672 (N_7672,N_5931,N_5533);
nor U7673 (N_7673,N_4287,N_3415);
nor U7674 (N_7674,N_4445,N_5937);
nor U7675 (N_7675,N_5565,N_4130);
nand U7676 (N_7676,N_4500,N_4123);
nand U7677 (N_7677,N_4387,N_5146);
nand U7678 (N_7678,N_3429,N_3069);
nor U7679 (N_7679,N_5313,N_3897);
nand U7680 (N_7680,N_4524,N_5946);
nand U7681 (N_7681,N_3103,N_5020);
and U7682 (N_7682,N_4954,N_4183);
nand U7683 (N_7683,N_3511,N_5678);
nand U7684 (N_7684,N_5211,N_5505);
and U7685 (N_7685,N_5819,N_3821);
nand U7686 (N_7686,N_3626,N_3143);
nor U7687 (N_7687,N_4496,N_4098);
and U7688 (N_7688,N_5403,N_5656);
or U7689 (N_7689,N_5363,N_4767);
nor U7690 (N_7690,N_5560,N_3573);
xor U7691 (N_7691,N_5507,N_3937);
or U7692 (N_7692,N_4577,N_4983);
and U7693 (N_7693,N_4403,N_3367);
nor U7694 (N_7694,N_5550,N_3342);
nand U7695 (N_7695,N_5676,N_3199);
nand U7696 (N_7696,N_4476,N_5454);
xor U7697 (N_7697,N_4374,N_3101);
nand U7698 (N_7698,N_5051,N_5277);
and U7699 (N_7699,N_3340,N_5207);
nand U7700 (N_7700,N_5785,N_5680);
or U7701 (N_7701,N_3860,N_5370);
and U7702 (N_7702,N_4301,N_3907);
nand U7703 (N_7703,N_4003,N_5677);
xor U7704 (N_7704,N_4216,N_4626);
or U7705 (N_7705,N_4241,N_4319);
or U7706 (N_7706,N_5152,N_4985);
or U7707 (N_7707,N_3302,N_5700);
or U7708 (N_7708,N_4324,N_3835);
xnor U7709 (N_7709,N_5137,N_4323);
or U7710 (N_7710,N_4423,N_5557);
and U7711 (N_7711,N_4311,N_4096);
and U7712 (N_7712,N_5499,N_5318);
xnor U7713 (N_7713,N_3964,N_3237);
or U7714 (N_7714,N_4629,N_5518);
nor U7715 (N_7715,N_4884,N_5177);
xor U7716 (N_7716,N_4465,N_5739);
or U7717 (N_7717,N_4761,N_3021);
nand U7718 (N_7718,N_4902,N_3146);
or U7719 (N_7719,N_5971,N_4923);
and U7720 (N_7720,N_5023,N_3786);
or U7721 (N_7721,N_3489,N_3398);
xnor U7722 (N_7722,N_4981,N_3888);
or U7723 (N_7723,N_4291,N_4519);
xor U7724 (N_7724,N_4014,N_3488);
nand U7725 (N_7725,N_3647,N_5654);
nor U7726 (N_7726,N_5848,N_3452);
and U7727 (N_7727,N_5470,N_5314);
or U7728 (N_7728,N_5834,N_3567);
or U7729 (N_7729,N_5315,N_5404);
and U7730 (N_7730,N_5065,N_5000);
nor U7731 (N_7731,N_4715,N_5164);
and U7732 (N_7732,N_5416,N_3016);
xor U7733 (N_7733,N_3416,N_3121);
or U7734 (N_7734,N_4918,N_3971);
nand U7735 (N_7735,N_4107,N_4248);
xnor U7736 (N_7736,N_4392,N_4756);
nand U7737 (N_7737,N_4736,N_4485);
xor U7738 (N_7738,N_5159,N_5086);
nor U7739 (N_7739,N_3389,N_5099);
xnor U7740 (N_7740,N_5764,N_4281);
and U7741 (N_7741,N_3246,N_4388);
nor U7742 (N_7742,N_3525,N_4962);
xor U7743 (N_7743,N_3714,N_3847);
nor U7744 (N_7744,N_4515,N_5083);
and U7745 (N_7745,N_3865,N_3433);
xor U7746 (N_7746,N_3900,N_5435);
nor U7747 (N_7747,N_5260,N_5179);
and U7748 (N_7748,N_5918,N_4450);
nand U7749 (N_7749,N_3764,N_3858);
nand U7750 (N_7750,N_5300,N_4648);
or U7751 (N_7751,N_5491,N_3183);
xor U7752 (N_7752,N_4243,N_4783);
nand U7753 (N_7753,N_4607,N_3171);
nand U7754 (N_7754,N_4116,N_5952);
or U7755 (N_7755,N_3824,N_5338);
xor U7756 (N_7756,N_5420,N_5166);
or U7757 (N_7757,N_4782,N_5561);
nor U7758 (N_7758,N_5483,N_4700);
nand U7759 (N_7759,N_4948,N_3474);
and U7760 (N_7760,N_3010,N_5943);
xor U7761 (N_7761,N_3108,N_5998);
and U7762 (N_7762,N_3279,N_5136);
nor U7763 (N_7763,N_3805,N_3795);
nand U7764 (N_7764,N_5433,N_4974);
and U7765 (N_7765,N_3073,N_4819);
and U7766 (N_7766,N_4117,N_5292);
xor U7767 (N_7767,N_4313,N_5831);
xor U7768 (N_7768,N_3889,N_5364);
and U7769 (N_7769,N_5151,N_4846);
nor U7770 (N_7770,N_4080,N_5529);
and U7771 (N_7771,N_3373,N_3047);
and U7772 (N_7772,N_5018,N_5124);
xnor U7773 (N_7773,N_3776,N_3877);
and U7774 (N_7774,N_5243,N_4517);
and U7775 (N_7775,N_3155,N_5385);
xor U7776 (N_7776,N_3753,N_4131);
xnor U7777 (N_7777,N_3799,N_5605);
nor U7778 (N_7778,N_5372,N_5592);
nand U7779 (N_7779,N_3235,N_3696);
xnor U7780 (N_7780,N_3151,N_3083);
and U7781 (N_7781,N_5528,N_5363);
xor U7782 (N_7782,N_5099,N_4018);
or U7783 (N_7783,N_4341,N_3127);
xnor U7784 (N_7784,N_4752,N_5500);
and U7785 (N_7785,N_3464,N_4074);
nand U7786 (N_7786,N_3841,N_5856);
and U7787 (N_7787,N_5766,N_5970);
or U7788 (N_7788,N_5985,N_5396);
nand U7789 (N_7789,N_5385,N_3215);
nor U7790 (N_7790,N_4485,N_4523);
xnor U7791 (N_7791,N_5451,N_3917);
and U7792 (N_7792,N_4822,N_5810);
and U7793 (N_7793,N_5810,N_5159);
or U7794 (N_7794,N_3084,N_3901);
and U7795 (N_7795,N_5328,N_3478);
nor U7796 (N_7796,N_5751,N_3180);
xor U7797 (N_7797,N_5783,N_5538);
xor U7798 (N_7798,N_3887,N_3314);
and U7799 (N_7799,N_3826,N_3241);
or U7800 (N_7800,N_5350,N_3038);
xnor U7801 (N_7801,N_5195,N_4731);
xor U7802 (N_7802,N_3751,N_3076);
and U7803 (N_7803,N_5966,N_3088);
nor U7804 (N_7804,N_3524,N_3325);
and U7805 (N_7805,N_3572,N_5265);
xor U7806 (N_7806,N_3013,N_5459);
nor U7807 (N_7807,N_4294,N_5015);
or U7808 (N_7808,N_3769,N_3210);
xnor U7809 (N_7809,N_3348,N_4666);
and U7810 (N_7810,N_4732,N_5642);
or U7811 (N_7811,N_4550,N_4659);
nand U7812 (N_7812,N_3095,N_5327);
nand U7813 (N_7813,N_5990,N_4944);
or U7814 (N_7814,N_5283,N_4352);
or U7815 (N_7815,N_3810,N_3014);
or U7816 (N_7816,N_4455,N_3746);
and U7817 (N_7817,N_4798,N_5843);
xor U7818 (N_7818,N_4109,N_5474);
or U7819 (N_7819,N_5485,N_3110);
xnor U7820 (N_7820,N_3720,N_5758);
nor U7821 (N_7821,N_5286,N_3821);
xnor U7822 (N_7822,N_4090,N_5470);
or U7823 (N_7823,N_5302,N_5413);
nor U7824 (N_7824,N_3385,N_5151);
or U7825 (N_7825,N_5040,N_5319);
nand U7826 (N_7826,N_5168,N_5096);
nor U7827 (N_7827,N_5683,N_4145);
xnor U7828 (N_7828,N_4046,N_3935);
and U7829 (N_7829,N_5966,N_5336);
nand U7830 (N_7830,N_4682,N_5190);
nor U7831 (N_7831,N_5623,N_3087);
xnor U7832 (N_7832,N_5229,N_5077);
xnor U7833 (N_7833,N_5751,N_3272);
nor U7834 (N_7834,N_4421,N_3605);
nor U7835 (N_7835,N_5172,N_4694);
nor U7836 (N_7836,N_4498,N_5920);
nor U7837 (N_7837,N_4066,N_5545);
and U7838 (N_7838,N_4279,N_5218);
xor U7839 (N_7839,N_3703,N_4007);
nand U7840 (N_7840,N_3107,N_3857);
and U7841 (N_7841,N_3262,N_3043);
and U7842 (N_7842,N_3272,N_5771);
nand U7843 (N_7843,N_3656,N_3064);
nand U7844 (N_7844,N_4190,N_3685);
xnor U7845 (N_7845,N_5617,N_3715);
or U7846 (N_7846,N_5899,N_4536);
nand U7847 (N_7847,N_5587,N_5665);
or U7848 (N_7848,N_3075,N_4308);
or U7849 (N_7849,N_3889,N_3863);
and U7850 (N_7850,N_4847,N_4489);
nand U7851 (N_7851,N_5573,N_3384);
xnor U7852 (N_7852,N_3853,N_3989);
nand U7853 (N_7853,N_5384,N_5163);
nand U7854 (N_7854,N_3092,N_5378);
xnor U7855 (N_7855,N_5751,N_4153);
nand U7856 (N_7856,N_3084,N_4377);
nand U7857 (N_7857,N_3691,N_4484);
nor U7858 (N_7858,N_5172,N_3404);
nand U7859 (N_7859,N_3577,N_5256);
xnor U7860 (N_7860,N_3120,N_3270);
xor U7861 (N_7861,N_5694,N_5966);
xor U7862 (N_7862,N_4334,N_3684);
xnor U7863 (N_7863,N_4131,N_3542);
or U7864 (N_7864,N_5539,N_5124);
or U7865 (N_7865,N_4651,N_5222);
xnor U7866 (N_7866,N_3541,N_3995);
xor U7867 (N_7867,N_3959,N_5526);
or U7868 (N_7868,N_5924,N_4304);
nor U7869 (N_7869,N_3181,N_4334);
nor U7870 (N_7870,N_3727,N_5559);
and U7871 (N_7871,N_4251,N_4668);
and U7872 (N_7872,N_4738,N_5442);
nor U7873 (N_7873,N_3793,N_5308);
nor U7874 (N_7874,N_5534,N_3377);
nor U7875 (N_7875,N_3317,N_3909);
and U7876 (N_7876,N_5510,N_4755);
xor U7877 (N_7877,N_4246,N_4216);
or U7878 (N_7878,N_4688,N_3056);
or U7879 (N_7879,N_4646,N_3850);
or U7880 (N_7880,N_4418,N_4768);
nor U7881 (N_7881,N_3337,N_3496);
or U7882 (N_7882,N_4963,N_3356);
xnor U7883 (N_7883,N_4712,N_3871);
and U7884 (N_7884,N_4167,N_5968);
xor U7885 (N_7885,N_4909,N_3366);
or U7886 (N_7886,N_3947,N_3137);
nor U7887 (N_7887,N_4643,N_4584);
and U7888 (N_7888,N_4577,N_5331);
xor U7889 (N_7889,N_3884,N_4383);
xnor U7890 (N_7890,N_4216,N_5751);
and U7891 (N_7891,N_4603,N_5656);
and U7892 (N_7892,N_5388,N_3622);
nor U7893 (N_7893,N_3316,N_5912);
and U7894 (N_7894,N_4855,N_3652);
nand U7895 (N_7895,N_5542,N_4110);
nand U7896 (N_7896,N_5353,N_5943);
or U7897 (N_7897,N_4419,N_4332);
nor U7898 (N_7898,N_4929,N_5605);
and U7899 (N_7899,N_3789,N_3583);
or U7900 (N_7900,N_5084,N_5300);
nor U7901 (N_7901,N_4364,N_4171);
and U7902 (N_7902,N_5538,N_5222);
or U7903 (N_7903,N_5979,N_3895);
nor U7904 (N_7904,N_4927,N_5022);
xnor U7905 (N_7905,N_4595,N_3473);
and U7906 (N_7906,N_5441,N_4169);
xnor U7907 (N_7907,N_4442,N_3432);
nor U7908 (N_7908,N_3520,N_3625);
xor U7909 (N_7909,N_3146,N_5228);
xnor U7910 (N_7910,N_3037,N_3579);
nor U7911 (N_7911,N_5440,N_4455);
and U7912 (N_7912,N_5262,N_5071);
nor U7913 (N_7913,N_5699,N_3017);
or U7914 (N_7914,N_4565,N_5688);
nor U7915 (N_7915,N_3191,N_3919);
nand U7916 (N_7916,N_3033,N_5523);
nand U7917 (N_7917,N_5837,N_4256);
nor U7918 (N_7918,N_4550,N_4004);
xor U7919 (N_7919,N_3743,N_4111);
nor U7920 (N_7920,N_4456,N_4359);
nand U7921 (N_7921,N_3187,N_5589);
or U7922 (N_7922,N_3793,N_5432);
and U7923 (N_7923,N_5647,N_4492);
nor U7924 (N_7924,N_3146,N_5126);
nand U7925 (N_7925,N_5319,N_5835);
and U7926 (N_7926,N_3407,N_3793);
xnor U7927 (N_7927,N_4046,N_5707);
and U7928 (N_7928,N_3659,N_4011);
xor U7929 (N_7929,N_5699,N_5595);
nand U7930 (N_7930,N_3919,N_3641);
nand U7931 (N_7931,N_5113,N_5661);
and U7932 (N_7932,N_3678,N_3032);
xnor U7933 (N_7933,N_5832,N_4206);
or U7934 (N_7934,N_3967,N_5518);
and U7935 (N_7935,N_4053,N_5524);
xnor U7936 (N_7936,N_5202,N_3402);
and U7937 (N_7937,N_5693,N_4123);
and U7938 (N_7938,N_3500,N_3238);
nand U7939 (N_7939,N_3828,N_4140);
and U7940 (N_7940,N_4387,N_5041);
nand U7941 (N_7941,N_3716,N_3568);
or U7942 (N_7942,N_4694,N_3741);
nor U7943 (N_7943,N_4228,N_3288);
or U7944 (N_7944,N_5359,N_4877);
nor U7945 (N_7945,N_4690,N_3343);
and U7946 (N_7946,N_5008,N_3282);
or U7947 (N_7947,N_3408,N_3617);
or U7948 (N_7948,N_4995,N_4522);
xnor U7949 (N_7949,N_4282,N_5396);
xnor U7950 (N_7950,N_5544,N_5946);
nand U7951 (N_7951,N_5580,N_3198);
and U7952 (N_7952,N_3097,N_3481);
and U7953 (N_7953,N_3635,N_3708);
or U7954 (N_7954,N_3136,N_5636);
xor U7955 (N_7955,N_5065,N_4230);
nand U7956 (N_7956,N_4472,N_3239);
nor U7957 (N_7957,N_3875,N_3793);
nor U7958 (N_7958,N_4331,N_4422);
xor U7959 (N_7959,N_4686,N_5524);
nor U7960 (N_7960,N_4928,N_3710);
and U7961 (N_7961,N_4029,N_4970);
and U7962 (N_7962,N_4574,N_5833);
xnor U7963 (N_7963,N_3333,N_4015);
xnor U7964 (N_7964,N_5013,N_4770);
or U7965 (N_7965,N_4488,N_5173);
xnor U7966 (N_7966,N_3296,N_4595);
xnor U7967 (N_7967,N_5855,N_5812);
nor U7968 (N_7968,N_4553,N_4659);
nor U7969 (N_7969,N_5976,N_4157);
nand U7970 (N_7970,N_3025,N_5807);
nor U7971 (N_7971,N_4418,N_3978);
nor U7972 (N_7972,N_3772,N_3115);
or U7973 (N_7973,N_5744,N_4415);
xor U7974 (N_7974,N_4996,N_5533);
or U7975 (N_7975,N_4570,N_4736);
or U7976 (N_7976,N_4479,N_3806);
or U7977 (N_7977,N_5161,N_5915);
nand U7978 (N_7978,N_3162,N_3236);
or U7979 (N_7979,N_4822,N_4815);
nand U7980 (N_7980,N_3478,N_4618);
nand U7981 (N_7981,N_4146,N_4696);
xor U7982 (N_7982,N_4231,N_3241);
nor U7983 (N_7983,N_4778,N_4324);
xor U7984 (N_7984,N_4324,N_4644);
or U7985 (N_7985,N_4835,N_5378);
nor U7986 (N_7986,N_5137,N_4893);
xnor U7987 (N_7987,N_3297,N_4545);
and U7988 (N_7988,N_5002,N_3208);
and U7989 (N_7989,N_4674,N_4970);
nand U7990 (N_7990,N_5653,N_3078);
and U7991 (N_7991,N_5026,N_5451);
xor U7992 (N_7992,N_5499,N_4193);
xnor U7993 (N_7993,N_4049,N_3242);
and U7994 (N_7994,N_4338,N_3316);
nor U7995 (N_7995,N_5605,N_4196);
or U7996 (N_7996,N_3990,N_5929);
xnor U7997 (N_7997,N_4446,N_3834);
xnor U7998 (N_7998,N_4656,N_3612);
nor U7999 (N_7999,N_4912,N_3742);
and U8000 (N_8000,N_5934,N_4204);
nand U8001 (N_8001,N_5370,N_4533);
xor U8002 (N_8002,N_5320,N_4875);
or U8003 (N_8003,N_5599,N_4107);
xor U8004 (N_8004,N_3008,N_3281);
and U8005 (N_8005,N_3702,N_4904);
xor U8006 (N_8006,N_4781,N_3742);
xnor U8007 (N_8007,N_4502,N_5470);
xor U8008 (N_8008,N_4273,N_5178);
nand U8009 (N_8009,N_4408,N_5820);
nor U8010 (N_8010,N_4625,N_5896);
nor U8011 (N_8011,N_4756,N_5513);
nand U8012 (N_8012,N_4636,N_4373);
xnor U8013 (N_8013,N_3605,N_5566);
nand U8014 (N_8014,N_4022,N_5222);
nand U8015 (N_8015,N_4119,N_3504);
nor U8016 (N_8016,N_4273,N_5527);
xor U8017 (N_8017,N_5027,N_3278);
nand U8018 (N_8018,N_3733,N_5547);
xor U8019 (N_8019,N_3934,N_4773);
xor U8020 (N_8020,N_3426,N_4858);
and U8021 (N_8021,N_3602,N_4299);
nor U8022 (N_8022,N_5789,N_3763);
xor U8023 (N_8023,N_4337,N_3581);
and U8024 (N_8024,N_5414,N_3948);
nor U8025 (N_8025,N_3450,N_3915);
and U8026 (N_8026,N_4436,N_5743);
nand U8027 (N_8027,N_5456,N_3612);
and U8028 (N_8028,N_4112,N_4015);
or U8029 (N_8029,N_5323,N_4832);
nand U8030 (N_8030,N_5573,N_5451);
xor U8031 (N_8031,N_5139,N_3955);
nand U8032 (N_8032,N_5221,N_4486);
xnor U8033 (N_8033,N_4915,N_3624);
xor U8034 (N_8034,N_4586,N_4958);
or U8035 (N_8035,N_3850,N_3527);
and U8036 (N_8036,N_4796,N_5920);
xor U8037 (N_8037,N_5113,N_5420);
and U8038 (N_8038,N_3725,N_3695);
nand U8039 (N_8039,N_5857,N_3533);
and U8040 (N_8040,N_3972,N_4397);
nand U8041 (N_8041,N_4346,N_5944);
or U8042 (N_8042,N_4566,N_3853);
xor U8043 (N_8043,N_3046,N_3376);
and U8044 (N_8044,N_5300,N_5649);
nor U8045 (N_8045,N_3103,N_5238);
nand U8046 (N_8046,N_4609,N_5516);
nor U8047 (N_8047,N_5202,N_5449);
nor U8048 (N_8048,N_3960,N_3400);
nand U8049 (N_8049,N_3736,N_4276);
nand U8050 (N_8050,N_4577,N_3352);
nor U8051 (N_8051,N_5044,N_4555);
nand U8052 (N_8052,N_4573,N_5438);
xnor U8053 (N_8053,N_5223,N_4795);
nor U8054 (N_8054,N_5630,N_4888);
and U8055 (N_8055,N_4091,N_4757);
xor U8056 (N_8056,N_4353,N_3968);
nor U8057 (N_8057,N_4496,N_5466);
and U8058 (N_8058,N_5448,N_4324);
and U8059 (N_8059,N_3332,N_5648);
xor U8060 (N_8060,N_5475,N_4142);
xor U8061 (N_8061,N_5877,N_5063);
and U8062 (N_8062,N_5790,N_5753);
or U8063 (N_8063,N_4015,N_5015);
and U8064 (N_8064,N_5094,N_5241);
xnor U8065 (N_8065,N_5418,N_3719);
and U8066 (N_8066,N_3496,N_4913);
nor U8067 (N_8067,N_3536,N_5991);
and U8068 (N_8068,N_4627,N_4223);
nand U8069 (N_8069,N_4314,N_3788);
xnor U8070 (N_8070,N_4171,N_4697);
and U8071 (N_8071,N_3365,N_5527);
xnor U8072 (N_8072,N_5867,N_3850);
and U8073 (N_8073,N_4791,N_5153);
xor U8074 (N_8074,N_4761,N_4190);
xnor U8075 (N_8075,N_4094,N_4352);
nor U8076 (N_8076,N_3014,N_4830);
and U8077 (N_8077,N_3499,N_3673);
and U8078 (N_8078,N_3009,N_4594);
xor U8079 (N_8079,N_3228,N_5686);
or U8080 (N_8080,N_4241,N_5822);
nand U8081 (N_8081,N_4724,N_3043);
nand U8082 (N_8082,N_5329,N_4234);
or U8083 (N_8083,N_4255,N_4920);
nand U8084 (N_8084,N_3961,N_5410);
and U8085 (N_8085,N_5935,N_5864);
and U8086 (N_8086,N_3130,N_3251);
or U8087 (N_8087,N_4601,N_5645);
nand U8088 (N_8088,N_5060,N_3904);
or U8089 (N_8089,N_4151,N_5475);
and U8090 (N_8090,N_3746,N_5154);
xnor U8091 (N_8091,N_5481,N_5229);
nor U8092 (N_8092,N_4578,N_4869);
nor U8093 (N_8093,N_3735,N_3845);
nor U8094 (N_8094,N_5183,N_4813);
and U8095 (N_8095,N_5009,N_5586);
xnor U8096 (N_8096,N_5088,N_4523);
xnor U8097 (N_8097,N_5087,N_5459);
nand U8098 (N_8098,N_4338,N_3097);
nor U8099 (N_8099,N_5639,N_4141);
xnor U8100 (N_8100,N_4535,N_4613);
xor U8101 (N_8101,N_4361,N_5990);
xor U8102 (N_8102,N_5721,N_4865);
nand U8103 (N_8103,N_5768,N_4892);
nor U8104 (N_8104,N_5044,N_4681);
nor U8105 (N_8105,N_4980,N_4775);
and U8106 (N_8106,N_4382,N_4486);
nand U8107 (N_8107,N_4734,N_4011);
xor U8108 (N_8108,N_3165,N_3647);
or U8109 (N_8109,N_5580,N_3273);
nand U8110 (N_8110,N_3485,N_3553);
nor U8111 (N_8111,N_5954,N_5538);
nand U8112 (N_8112,N_4535,N_5063);
or U8113 (N_8113,N_3858,N_3152);
nor U8114 (N_8114,N_3070,N_4925);
nor U8115 (N_8115,N_4218,N_5602);
and U8116 (N_8116,N_4157,N_3433);
and U8117 (N_8117,N_5892,N_3232);
or U8118 (N_8118,N_3291,N_4000);
nand U8119 (N_8119,N_3234,N_4332);
nor U8120 (N_8120,N_4211,N_4789);
xnor U8121 (N_8121,N_5640,N_5100);
nand U8122 (N_8122,N_4384,N_4520);
nand U8123 (N_8123,N_3826,N_4120);
or U8124 (N_8124,N_4841,N_5863);
nor U8125 (N_8125,N_3193,N_4082);
and U8126 (N_8126,N_5926,N_5637);
xor U8127 (N_8127,N_5823,N_5517);
nor U8128 (N_8128,N_5061,N_3879);
or U8129 (N_8129,N_3034,N_4239);
nand U8130 (N_8130,N_5418,N_4189);
and U8131 (N_8131,N_5316,N_3662);
nor U8132 (N_8132,N_5478,N_3209);
xor U8133 (N_8133,N_3744,N_3724);
nor U8134 (N_8134,N_5117,N_5751);
nor U8135 (N_8135,N_4328,N_5146);
xor U8136 (N_8136,N_4180,N_3494);
or U8137 (N_8137,N_5157,N_5109);
and U8138 (N_8138,N_4318,N_4734);
xnor U8139 (N_8139,N_3453,N_5315);
and U8140 (N_8140,N_5954,N_4690);
nor U8141 (N_8141,N_3122,N_3011);
xor U8142 (N_8142,N_4306,N_5137);
nand U8143 (N_8143,N_4801,N_4133);
or U8144 (N_8144,N_3156,N_5346);
or U8145 (N_8145,N_4370,N_5552);
nand U8146 (N_8146,N_5024,N_4747);
or U8147 (N_8147,N_3865,N_4765);
xor U8148 (N_8148,N_3913,N_4433);
and U8149 (N_8149,N_3139,N_5207);
nand U8150 (N_8150,N_5791,N_3975);
nand U8151 (N_8151,N_3417,N_5543);
nand U8152 (N_8152,N_3120,N_5917);
nand U8153 (N_8153,N_5542,N_5711);
or U8154 (N_8154,N_4156,N_4239);
nor U8155 (N_8155,N_5802,N_4676);
and U8156 (N_8156,N_5098,N_4543);
nand U8157 (N_8157,N_5553,N_3027);
and U8158 (N_8158,N_3109,N_5598);
nand U8159 (N_8159,N_5867,N_5298);
xor U8160 (N_8160,N_5545,N_5791);
xor U8161 (N_8161,N_4076,N_3481);
nor U8162 (N_8162,N_3696,N_5224);
and U8163 (N_8163,N_4621,N_5330);
or U8164 (N_8164,N_4340,N_3030);
xor U8165 (N_8165,N_4894,N_4275);
or U8166 (N_8166,N_4597,N_3595);
or U8167 (N_8167,N_5521,N_3760);
xor U8168 (N_8168,N_5947,N_5585);
and U8169 (N_8169,N_4059,N_4910);
and U8170 (N_8170,N_4453,N_5331);
nor U8171 (N_8171,N_3943,N_5816);
and U8172 (N_8172,N_4537,N_5657);
and U8173 (N_8173,N_4851,N_5755);
nor U8174 (N_8174,N_4796,N_5155);
nor U8175 (N_8175,N_4654,N_3668);
and U8176 (N_8176,N_4017,N_4070);
and U8177 (N_8177,N_3878,N_3261);
and U8178 (N_8178,N_4994,N_4561);
xor U8179 (N_8179,N_5030,N_4327);
or U8180 (N_8180,N_3716,N_4142);
and U8181 (N_8181,N_5561,N_5778);
or U8182 (N_8182,N_4060,N_5720);
and U8183 (N_8183,N_5948,N_4256);
xor U8184 (N_8184,N_4530,N_3208);
xor U8185 (N_8185,N_5190,N_5948);
or U8186 (N_8186,N_4650,N_3171);
xnor U8187 (N_8187,N_5456,N_3051);
and U8188 (N_8188,N_4414,N_5890);
and U8189 (N_8189,N_3714,N_3822);
nor U8190 (N_8190,N_4149,N_5108);
nand U8191 (N_8191,N_4307,N_3115);
nand U8192 (N_8192,N_3603,N_3351);
and U8193 (N_8193,N_5026,N_5520);
xor U8194 (N_8194,N_4062,N_5266);
nor U8195 (N_8195,N_3837,N_3641);
and U8196 (N_8196,N_3875,N_3332);
nor U8197 (N_8197,N_4129,N_4130);
or U8198 (N_8198,N_3166,N_4243);
or U8199 (N_8199,N_5866,N_3853);
xnor U8200 (N_8200,N_4220,N_5600);
and U8201 (N_8201,N_4187,N_5143);
or U8202 (N_8202,N_3565,N_5737);
and U8203 (N_8203,N_3992,N_3762);
nand U8204 (N_8204,N_5352,N_3558);
nand U8205 (N_8205,N_3083,N_5825);
nor U8206 (N_8206,N_3724,N_5940);
or U8207 (N_8207,N_3842,N_5716);
or U8208 (N_8208,N_4302,N_3572);
nand U8209 (N_8209,N_4290,N_5139);
nand U8210 (N_8210,N_5553,N_3713);
nor U8211 (N_8211,N_5390,N_3522);
and U8212 (N_8212,N_4638,N_3361);
xor U8213 (N_8213,N_3252,N_3007);
and U8214 (N_8214,N_3661,N_5028);
or U8215 (N_8215,N_3561,N_4733);
xnor U8216 (N_8216,N_4409,N_3886);
xor U8217 (N_8217,N_5842,N_5953);
or U8218 (N_8218,N_5721,N_4367);
or U8219 (N_8219,N_3298,N_3688);
nor U8220 (N_8220,N_3801,N_5610);
or U8221 (N_8221,N_5530,N_5406);
xnor U8222 (N_8222,N_3750,N_5106);
nor U8223 (N_8223,N_4678,N_3250);
or U8224 (N_8224,N_5052,N_5283);
or U8225 (N_8225,N_4480,N_4325);
and U8226 (N_8226,N_3052,N_3684);
nand U8227 (N_8227,N_5746,N_4045);
or U8228 (N_8228,N_3782,N_5174);
or U8229 (N_8229,N_5992,N_5833);
xor U8230 (N_8230,N_4495,N_5725);
xnor U8231 (N_8231,N_5036,N_4228);
nor U8232 (N_8232,N_4048,N_4664);
or U8233 (N_8233,N_3610,N_4419);
and U8234 (N_8234,N_4201,N_4821);
and U8235 (N_8235,N_3013,N_3798);
nor U8236 (N_8236,N_5255,N_4402);
and U8237 (N_8237,N_4090,N_3839);
xnor U8238 (N_8238,N_5361,N_3600);
nor U8239 (N_8239,N_4242,N_4954);
nor U8240 (N_8240,N_3686,N_4304);
nor U8241 (N_8241,N_4208,N_3234);
nand U8242 (N_8242,N_4046,N_3777);
or U8243 (N_8243,N_5291,N_4164);
or U8244 (N_8244,N_4708,N_4643);
and U8245 (N_8245,N_5798,N_5857);
and U8246 (N_8246,N_3221,N_3844);
or U8247 (N_8247,N_5093,N_3454);
or U8248 (N_8248,N_5708,N_3021);
or U8249 (N_8249,N_5910,N_3491);
or U8250 (N_8250,N_5775,N_4319);
nor U8251 (N_8251,N_3241,N_4584);
nand U8252 (N_8252,N_5642,N_4077);
xor U8253 (N_8253,N_3216,N_5402);
and U8254 (N_8254,N_5793,N_3171);
nand U8255 (N_8255,N_5544,N_4464);
or U8256 (N_8256,N_4807,N_5874);
or U8257 (N_8257,N_5137,N_3624);
nand U8258 (N_8258,N_5920,N_5974);
xnor U8259 (N_8259,N_4692,N_3565);
nand U8260 (N_8260,N_3660,N_3386);
or U8261 (N_8261,N_4254,N_3643);
nand U8262 (N_8262,N_5323,N_4614);
and U8263 (N_8263,N_3665,N_3040);
or U8264 (N_8264,N_4630,N_3438);
nor U8265 (N_8265,N_5884,N_5085);
and U8266 (N_8266,N_4990,N_3544);
xnor U8267 (N_8267,N_5001,N_5195);
nor U8268 (N_8268,N_4338,N_4845);
nor U8269 (N_8269,N_3903,N_4857);
and U8270 (N_8270,N_4743,N_5312);
nand U8271 (N_8271,N_5227,N_5598);
nor U8272 (N_8272,N_5162,N_3236);
nor U8273 (N_8273,N_3783,N_4375);
nand U8274 (N_8274,N_4641,N_4986);
and U8275 (N_8275,N_4384,N_5396);
or U8276 (N_8276,N_3909,N_3316);
xor U8277 (N_8277,N_4943,N_5199);
nor U8278 (N_8278,N_4638,N_3090);
or U8279 (N_8279,N_5085,N_3328);
or U8280 (N_8280,N_4418,N_4469);
and U8281 (N_8281,N_3449,N_3736);
nand U8282 (N_8282,N_5135,N_5107);
or U8283 (N_8283,N_3736,N_3789);
nor U8284 (N_8284,N_4310,N_5887);
or U8285 (N_8285,N_5726,N_3774);
nor U8286 (N_8286,N_5151,N_4456);
nor U8287 (N_8287,N_4160,N_5517);
nor U8288 (N_8288,N_3792,N_5922);
xor U8289 (N_8289,N_3486,N_4414);
xor U8290 (N_8290,N_5073,N_3634);
nand U8291 (N_8291,N_3596,N_4432);
nand U8292 (N_8292,N_3668,N_5891);
nor U8293 (N_8293,N_5444,N_3444);
xor U8294 (N_8294,N_4750,N_3382);
xnor U8295 (N_8295,N_5944,N_3860);
and U8296 (N_8296,N_3245,N_5186);
nand U8297 (N_8297,N_4589,N_4899);
and U8298 (N_8298,N_5514,N_4271);
xnor U8299 (N_8299,N_3198,N_4872);
nor U8300 (N_8300,N_3373,N_4311);
or U8301 (N_8301,N_5115,N_4064);
nand U8302 (N_8302,N_3987,N_4254);
nand U8303 (N_8303,N_3038,N_3727);
and U8304 (N_8304,N_5828,N_4035);
nor U8305 (N_8305,N_3641,N_4482);
and U8306 (N_8306,N_4006,N_4055);
nand U8307 (N_8307,N_5532,N_4666);
or U8308 (N_8308,N_4264,N_3041);
and U8309 (N_8309,N_4569,N_3702);
xnor U8310 (N_8310,N_4029,N_4056);
or U8311 (N_8311,N_4079,N_4455);
and U8312 (N_8312,N_4174,N_5204);
or U8313 (N_8313,N_3721,N_4244);
xnor U8314 (N_8314,N_5931,N_3379);
nor U8315 (N_8315,N_4530,N_5756);
nor U8316 (N_8316,N_4088,N_4545);
xor U8317 (N_8317,N_3246,N_5276);
nand U8318 (N_8318,N_4444,N_4510);
and U8319 (N_8319,N_4936,N_5498);
nor U8320 (N_8320,N_5203,N_3931);
nand U8321 (N_8321,N_4306,N_5972);
nand U8322 (N_8322,N_5207,N_3402);
and U8323 (N_8323,N_4369,N_5165);
and U8324 (N_8324,N_5680,N_3757);
or U8325 (N_8325,N_4129,N_4229);
and U8326 (N_8326,N_5788,N_4857);
or U8327 (N_8327,N_5193,N_3436);
and U8328 (N_8328,N_5088,N_5608);
xor U8329 (N_8329,N_3784,N_5351);
xnor U8330 (N_8330,N_5364,N_5267);
nor U8331 (N_8331,N_5150,N_3129);
and U8332 (N_8332,N_5336,N_5955);
nor U8333 (N_8333,N_3259,N_3077);
and U8334 (N_8334,N_5655,N_5399);
nand U8335 (N_8335,N_5858,N_5125);
nor U8336 (N_8336,N_3744,N_4983);
nand U8337 (N_8337,N_4822,N_5903);
nand U8338 (N_8338,N_5301,N_4256);
and U8339 (N_8339,N_4616,N_4391);
and U8340 (N_8340,N_3434,N_4158);
or U8341 (N_8341,N_4054,N_4868);
or U8342 (N_8342,N_3628,N_4826);
nor U8343 (N_8343,N_5313,N_3537);
or U8344 (N_8344,N_5018,N_3375);
and U8345 (N_8345,N_5125,N_3804);
xor U8346 (N_8346,N_4084,N_3027);
or U8347 (N_8347,N_5842,N_3158);
nand U8348 (N_8348,N_4780,N_3918);
nor U8349 (N_8349,N_3264,N_3024);
nor U8350 (N_8350,N_3459,N_4606);
nor U8351 (N_8351,N_5860,N_5622);
and U8352 (N_8352,N_5026,N_5146);
nand U8353 (N_8353,N_3136,N_4337);
nand U8354 (N_8354,N_5820,N_5141);
nor U8355 (N_8355,N_3231,N_5680);
nand U8356 (N_8356,N_5088,N_3552);
nor U8357 (N_8357,N_4212,N_5827);
and U8358 (N_8358,N_4643,N_4163);
or U8359 (N_8359,N_4667,N_3946);
nand U8360 (N_8360,N_4741,N_4434);
and U8361 (N_8361,N_3821,N_3061);
and U8362 (N_8362,N_4513,N_3153);
and U8363 (N_8363,N_4809,N_3286);
nand U8364 (N_8364,N_4103,N_3955);
xor U8365 (N_8365,N_4463,N_3967);
nand U8366 (N_8366,N_5959,N_5729);
xor U8367 (N_8367,N_5519,N_5783);
nor U8368 (N_8368,N_4252,N_4870);
nor U8369 (N_8369,N_5071,N_3604);
nor U8370 (N_8370,N_5553,N_3328);
nor U8371 (N_8371,N_4706,N_4407);
nor U8372 (N_8372,N_3602,N_4926);
or U8373 (N_8373,N_5902,N_3515);
nand U8374 (N_8374,N_3863,N_5488);
and U8375 (N_8375,N_3960,N_4706);
or U8376 (N_8376,N_5276,N_4236);
xor U8377 (N_8377,N_5367,N_3878);
xor U8378 (N_8378,N_3350,N_3669);
xor U8379 (N_8379,N_4493,N_5350);
xor U8380 (N_8380,N_4120,N_5130);
and U8381 (N_8381,N_4690,N_4945);
xor U8382 (N_8382,N_3947,N_5851);
xor U8383 (N_8383,N_5046,N_4468);
or U8384 (N_8384,N_4642,N_4325);
xnor U8385 (N_8385,N_4410,N_3287);
and U8386 (N_8386,N_3392,N_3688);
nand U8387 (N_8387,N_5017,N_5043);
nand U8388 (N_8388,N_5676,N_5742);
xnor U8389 (N_8389,N_4467,N_4102);
xor U8390 (N_8390,N_4654,N_4415);
nand U8391 (N_8391,N_5584,N_5000);
and U8392 (N_8392,N_3825,N_5478);
or U8393 (N_8393,N_5155,N_3673);
xor U8394 (N_8394,N_4587,N_4981);
and U8395 (N_8395,N_5713,N_4998);
or U8396 (N_8396,N_3335,N_3332);
and U8397 (N_8397,N_5829,N_3731);
nor U8398 (N_8398,N_4978,N_5743);
and U8399 (N_8399,N_4569,N_4756);
or U8400 (N_8400,N_4321,N_4294);
xnor U8401 (N_8401,N_4836,N_5644);
and U8402 (N_8402,N_3612,N_4836);
nand U8403 (N_8403,N_4637,N_5040);
nand U8404 (N_8404,N_4463,N_3498);
or U8405 (N_8405,N_5714,N_4373);
or U8406 (N_8406,N_5452,N_5783);
or U8407 (N_8407,N_5672,N_3542);
or U8408 (N_8408,N_3645,N_4546);
or U8409 (N_8409,N_3729,N_3683);
xnor U8410 (N_8410,N_3268,N_4325);
or U8411 (N_8411,N_5973,N_3883);
xnor U8412 (N_8412,N_5356,N_5634);
xnor U8413 (N_8413,N_3450,N_3498);
nor U8414 (N_8414,N_4797,N_3015);
xnor U8415 (N_8415,N_5453,N_3235);
or U8416 (N_8416,N_3490,N_3954);
or U8417 (N_8417,N_3578,N_5886);
or U8418 (N_8418,N_3040,N_3413);
nand U8419 (N_8419,N_4304,N_5096);
or U8420 (N_8420,N_4386,N_3785);
nand U8421 (N_8421,N_5542,N_5916);
nor U8422 (N_8422,N_5714,N_3646);
nand U8423 (N_8423,N_4962,N_3204);
and U8424 (N_8424,N_5361,N_4002);
xnor U8425 (N_8425,N_4063,N_4230);
nand U8426 (N_8426,N_5589,N_5609);
and U8427 (N_8427,N_4401,N_3743);
or U8428 (N_8428,N_5454,N_5621);
xnor U8429 (N_8429,N_5175,N_4047);
xor U8430 (N_8430,N_4180,N_5521);
nor U8431 (N_8431,N_3796,N_5447);
or U8432 (N_8432,N_5445,N_5986);
nand U8433 (N_8433,N_5608,N_3761);
nand U8434 (N_8434,N_5170,N_4223);
or U8435 (N_8435,N_5944,N_3534);
xor U8436 (N_8436,N_5267,N_5509);
xnor U8437 (N_8437,N_4527,N_3540);
nand U8438 (N_8438,N_3366,N_5579);
xor U8439 (N_8439,N_3109,N_4333);
and U8440 (N_8440,N_3510,N_4650);
nand U8441 (N_8441,N_4569,N_4539);
nor U8442 (N_8442,N_5930,N_4719);
nand U8443 (N_8443,N_5271,N_3819);
xnor U8444 (N_8444,N_4937,N_3510);
and U8445 (N_8445,N_3587,N_4048);
nand U8446 (N_8446,N_3052,N_5871);
nor U8447 (N_8447,N_4898,N_4656);
nand U8448 (N_8448,N_5300,N_5821);
and U8449 (N_8449,N_4931,N_4875);
and U8450 (N_8450,N_3187,N_3548);
or U8451 (N_8451,N_4656,N_5075);
xnor U8452 (N_8452,N_3155,N_4018);
xor U8453 (N_8453,N_4590,N_3454);
or U8454 (N_8454,N_5943,N_4350);
nand U8455 (N_8455,N_5760,N_5381);
xor U8456 (N_8456,N_3021,N_5844);
and U8457 (N_8457,N_4092,N_4687);
or U8458 (N_8458,N_5707,N_5857);
and U8459 (N_8459,N_5795,N_3248);
or U8460 (N_8460,N_4509,N_4830);
nor U8461 (N_8461,N_5528,N_4255);
xnor U8462 (N_8462,N_3693,N_3097);
nor U8463 (N_8463,N_4324,N_5736);
xnor U8464 (N_8464,N_5424,N_5920);
nor U8465 (N_8465,N_4586,N_3295);
xor U8466 (N_8466,N_4890,N_4047);
and U8467 (N_8467,N_3791,N_3132);
nor U8468 (N_8468,N_4776,N_3480);
xor U8469 (N_8469,N_3017,N_3245);
nor U8470 (N_8470,N_4555,N_4167);
nand U8471 (N_8471,N_4681,N_3497);
xor U8472 (N_8472,N_3930,N_5870);
xnor U8473 (N_8473,N_5017,N_3677);
nand U8474 (N_8474,N_4831,N_4239);
and U8475 (N_8475,N_4521,N_4644);
xor U8476 (N_8476,N_3464,N_4658);
xor U8477 (N_8477,N_3163,N_4484);
nor U8478 (N_8478,N_3055,N_4413);
xnor U8479 (N_8479,N_5892,N_4354);
nor U8480 (N_8480,N_4187,N_5773);
nand U8481 (N_8481,N_3184,N_4861);
or U8482 (N_8482,N_4129,N_5067);
nand U8483 (N_8483,N_5312,N_3938);
nor U8484 (N_8484,N_3368,N_5757);
nand U8485 (N_8485,N_4748,N_3287);
and U8486 (N_8486,N_4076,N_4852);
nor U8487 (N_8487,N_5781,N_5202);
xor U8488 (N_8488,N_4404,N_4050);
nor U8489 (N_8489,N_4707,N_3146);
nand U8490 (N_8490,N_4904,N_4246);
nor U8491 (N_8491,N_3469,N_3397);
nand U8492 (N_8492,N_3917,N_5101);
nand U8493 (N_8493,N_3579,N_3729);
nand U8494 (N_8494,N_5009,N_3145);
or U8495 (N_8495,N_4605,N_4866);
xnor U8496 (N_8496,N_4757,N_3510);
or U8497 (N_8497,N_4129,N_3947);
nor U8498 (N_8498,N_5885,N_5519);
and U8499 (N_8499,N_4179,N_5338);
or U8500 (N_8500,N_3049,N_3966);
nor U8501 (N_8501,N_5387,N_3778);
and U8502 (N_8502,N_4690,N_3919);
xor U8503 (N_8503,N_3955,N_3699);
and U8504 (N_8504,N_3941,N_4701);
nand U8505 (N_8505,N_3498,N_4632);
xnor U8506 (N_8506,N_4167,N_5905);
nor U8507 (N_8507,N_4516,N_5583);
and U8508 (N_8508,N_4778,N_3877);
and U8509 (N_8509,N_4907,N_3133);
xor U8510 (N_8510,N_4558,N_3616);
xnor U8511 (N_8511,N_3390,N_4245);
nor U8512 (N_8512,N_5741,N_5225);
and U8513 (N_8513,N_3686,N_3480);
nor U8514 (N_8514,N_3253,N_4012);
and U8515 (N_8515,N_3189,N_3546);
xnor U8516 (N_8516,N_3023,N_4772);
or U8517 (N_8517,N_5376,N_5668);
nor U8518 (N_8518,N_3837,N_3591);
nor U8519 (N_8519,N_3162,N_3160);
nand U8520 (N_8520,N_3990,N_4007);
and U8521 (N_8521,N_3048,N_5495);
nand U8522 (N_8522,N_4279,N_5510);
or U8523 (N_8523,N_5029,N_5220);
nand U8524 (N_8524,N_3348,N_4841);
or U8525 (N_8525,N_5019,N_4754);
xor U8526 (N_8526,N_4532,N_3974);
or U8527 (N_8527,N_4993,N_4467);
nor U8528 (N_8528,N_3133,N_5856);
nand U8529 (N_8529,N_4863,N_3173);
and U8530 (N_8530,N_4519,N_5297);
nand U8531 (N_8531,N_5215,N_3989);
and U8532 (N_8532,N_5282,N_4767);
and U8533 (N_8533,N_4841,N_3261);
nor U8534 (N_8534,N_4868,N_3410);
and U8535 (N_8535,N_3929,N_3813);
nor U8536 (N_8536,N_5895,N_5151);
nand U8537 (N_8537,N_4039,N_5536);
xnor U8538 (N_8538,N_3832,N_4511);
or U8539 (N_8539,N_4673,N_4802);
nand U8540 (N_8540,N_3838,N_3899);
nand U8541 (N_8541,N_4723,N_3878);
and U8542 (N_8542,N_5446,N_4471);
and U8543 (N_8543,N_3180,N_3266);
nor U8544 (N_8544,N_5397,N_5611);
and U8545 (N_8545,N_3304,N_5169);
nor U8546 (N_8546,N_4542,N_3023);
and U8547 (N_8547,N_3626,N_3934);
xnor U8548 (N_8548,N_5327,N_3517);
nor U8549 (N_8549,N_3295,N_4999);
nor U8550 (N_8550,N_5809,N_4707);
nand U8551 (N_8551,N_5731,N_4904);
nor U8552 (N_8552,N_4383,N_4292);
and U8553 (N_8553,N_5755,N_4740);
xnor U8554 (N_8554,N_3325,N_5263);
or U8555 (N_8555,N_3702,N_5278);
xor U8556 (N_8556,N_3473,N_5218);
xnor U8557 (N_8557,N_4286,N_3275);
xor U8558 (N_8558,N_5025,N_5410);
or U8559 (N_8559,N_3674,N_3268);
or U8560 (N_8560,N_3435,N_5683);
xor U8561 (N_8561,N_3037,N_3057);
and U8562 (N_8562,N_4487,N_4599);
and U8563 (N_8563,N_4157,N_4320);
nand U8564 (N_8564,N_5541,N_3171);
nor U8565 (N_8565,N_3424,N_4151);
and U8566 (N_8566,N_4527,N_3126);
nor U8567 (N_8567,N_4475,N_4612);
or U8568 (N_8568,N_5108,N_3673);
or U8569 (N_8569,N_4754,N_4936);
and U8570 (N_8570,N_3808,N_5364);
nand U8571 (N_8571,N_5665,N_3687);
and U8572 (N_8572,N_3494,N_5368);
nand U8573 (N_8573,N_4360,N_3182);
nor U8574 (N_8574,N_3277,N_3699);
or U8575 (N_8575,N_4750,N_5553);
and U8576 (N_8576,N_3233,N_4042);
or U8577 (N_8577,N_3112,N_5731);
nand U8578 (N_8578,N_4538,N_4561);
or U8579 (N_8579,N_5272,N_4748);
and U8580 (N_8580,N_3316,N_5390);
nand U8581 (N_8581,N_4355,N_4984);
or U8582 (N_8582,N_5494,N_5567);
and U8583 (N_8583,N_3011,N_4806);
nor U8584 (N_8584,N_5162,N_3580);
nor U8585 (N_8585,N_4100,N_3353);
nand U8586 (N_8586,N_5683,N_5305);
and U8587 (N_8587,N_5774,N_4012);
nor U8588 (N_8588,N_3867,N_3766);
xor U8589 (N_8589,N_3818,N_3833);
xor U8590 (N_8590,N_3228,N_4551);
and U8591 (N_8591,N_3985,N_5808);
xor U8592 (N_8592,N_5661,N_4213);
or U8593 (N_8593,N_5669,N_3329);
nor U8594 (N_8594,N_3245,N_5728);
nand U8595 (N_8595,N_3307,N_4736);
nand U8596 (N_8596,N_4403,N_5293);
nand U8597 (N_8597,N_3474,N_4543);
or U8598 (N_8598,N_4384,N_4371);
xor U8599 (N_8599,N_4049,N_3879);
or U8600 (N_8600,N_5244,N_4462);
and U8601 (N_8601,N_4504,N_4128);
nand U8602 (N_8602,N_3043,N_5633);
or U8603 (N_8603,N_5730,N_5138);
nand U8604 (N_8604,N_5597,N_3837);
xnor U8605 (N_8605,N_5184,N_5814);
nand U8606 (N_8606,N_5226,N_5368);
nor U8607 (N_8607,N_3221,N_3197);
nor U8608 (N_8608,N_3149,N_5314);
xnor U8609 (N_8609,N_3498,N_3293);
and U8610 (N_8610,N_3473,N_3343);
nand U8611 (N_8611,N_3014,N_4169);
nor U8612 (N_8612,N_4479,N_3227);
and U8613 (N_8613,N_4557,N_4181);
xor U8614 (N_8614,N_4569,N_3902);
xor U8615 (N_8615,N_5119,N_4071);
or U8616 (N_8616,N_5389,N_5824);
and U8617 (N_8617,N_5869,N_3116);
xor U8618 (N_8618,N_5815,N_4854);
nand U8619 (N_8619,N_4210,N_4352);
xnor U8620 (N_8620,N_4253,N_4841);
nand U8621 (N_8621,N_3002,N_3724);
and U8622 (N_8622,N_4707,N_3590);
nand U8623 (N_8623,N_3035,N_5895);
and U8624 (N_8624,N_3064,N_4646);
nor U8625 (N_8625,N_3571,N_5892);
xor U8626 (N_8626,N_4659,N_5225);
and U8627 (N_8627,N_3445,N_5410);
xnor U8628 (N_8628,N_5017,N_3561);
nand U8629 (N_8629,N_3496,N_4140);
and U8630 (N_8630,N_3314,N_3188);
xor U8631 (N_8631,N_5495,N_3199);
xor U8632 (N_8632,N_3569,N_5549);
nand U8633 (N_8633,N_4091,N_5131);
nor U8634 (N_8634,N_3824,N_3315);
nor U8635 (N_8635,N_5415,N_5332);
nand U8636 (N_8636,N_5983,N_5330);
xnor U8637 (N_8637,N_5658,N_5708);
nor U8638 (N_8638,N_5291,N_5679);
xor U8639 (N_8639,N_5604,N_3932);
and U8640 (N_8640,N_4660,N_3056);
xor U8641 (N_8641,N_4477,N_4203);
or U8642 (N_8642,N_4672,N_5272);
xor U8643 (N_8643,N_5180,N_5872);
xor U8644 (N_8644,N_3888,N_5902);
and U8645 (N_8645,N_4239,N_4876);
nand U8646 (N_8646,N_5576,N_4671);
or U8647 (N_8647,N_4048,N_5542);
or U8648 (N_8648,N_5129,N_5908);
xor U8649 (N_8649,N_3467,N_4560);
or U8650 (N_8650,N_5924,N_3770);
xnor U8651 (N_8651,N_5297,N_5707);
nand U8652 (N_8652,N_4740,N_3290);
nand U8653 (N_8653,N_3413,N_3385);
nand U8654 (N_8654,N_3191,N_5290);
xor U8655 (N_8655,N_3273,N_3789);
nor U8656 (N_8656,N_3128,N_3984);
and U8657 (N_8657,N_4680,N_4175);
xor U8658 (N_8658,N_4599,N_4856);
or U8659 (N_8659,N_5215,N_5176);
nor U8660 (N_8660,N_4177,N_4505);
xnor U8661 (N_8661,N_4520,N_3374);
or U8662 (N_8662,N_4228,N_3597);
xnor U8663 (N_8663,N_4148,N_3547);
and U8664 (N_8664,N_4068,N_4338);
or U8665 (N_8665,N_3461,N_5587);
and U8666 (N_8666,N_3813,N_4414);
and U8667 (N_8667,N_4614,N_5272);
or U8668 (N_8668,N_3177,N_3154);
nor U8669 (N_8669,N_3065,N_5024);
nor U8670 (N_8670,N_4141,N_3866);
nor U8671 (N_8671,N_4189,N_4972);
nand U8672 (N_8672,N_3638,N_4568);
xor U8673 (N_8673,N_5900,N_3353);
or U8674 (N_8674,N_4468,N_4065);
xnor U8675 (N_8675,N_3522,N_3521);
xor U8676 (N_8676,N_4450,N_4122);
and U8677 (N_8677,N_3433,N_5389);
or U8678 (N_8678,N_3220,N_5981);
or U8679 (N_8679,N_4846,N_3184);
or U8680 (N_8680,N_5414,N_3413);
xnor U8681 (N_8681,N_4605,N_3136);
nand U8682 (N_8682,N_4450,N_4073);
nand U8683 (N_8683,N_5878,N_5813);
and U8684 (N_8684,N_4323,N_4447);
xor U8685 (N_8685,N_5698,N_5950);
and U8686 (N_8686,N_5683,N_4271);
nor U8687 (N_8687,N_5185,N_5145);
xnor U8688 (N_8688,N_3471,N_5566);
nand U8689 (N_8689,N_3826,N_5698);
and U8690 (N_8690,N_3872,N_5231);
xnor U8691 (N_8691,N_5823,N_4083);
xnor U8692 (N_8692,N_5219,N_5091);
and U8693 (N_8693,N_3254,N_4146);
and U8694 (N_8694,N_4794,N_3580);
nand U8695 (N_8695,N_3560,N_5647);
or U8696 (N_8696,N_4317,N_5743);
xnor U8697 (N_8697,N_5324,N_5750);
and U8698 (N_8698,N_4369,N_5315);
nor U8699 (N_8699,N_3418,N_4932);
nor U8700 (N_8700,N_4902,N_4121);
xnor U8701 (N_8701,N_3221,N_5984);
nor U8702 (N_8702,N_5265,N_5994);
and U8703 (N_8703,N_5574,N_5268);
nor U8704 (N_8704,N_5794,N_5627);
and U8705 (N_8705,N_3197,N_4681);
xnor U8706 (N_8706,N_4189,N_4123);
xor U8707 (N_8707,N_4748,N_5107);
nand U8708 (N_8708,N_5214,N_3498);
and U8709 (N_8709,N_5625,N_4610);
nand U8710 (N_8710,N_3497,N_5863);
nand U8711 (N_8711,N_5072,N_5086);
and U8712 (N_8712,N_3640,N_4760);
xnor U8713 (N_8713,N_5692,N_3346);
nand U8714 (N_8714,N_4600,N_5898);
and U8715 (N_8715,N_3976,N_3826);
and U8716 (N_8716,N_3213,N_4927);
nand U8717 (N_8717,N_4143,N_5455);
nor U8718 (N_8718,N_5797,N_3385);
and U8719 (N_8719,N_3941,N_3109);
nand U8720 (N_8720,N_3999,N_5729);
xnor U8721 (N_8721,N_5512,N_3577);
and U8722 (N_8722,N_3768,N_3164);
and U8723 (N_8723,N_5412,N_5963);
or U8724 (N_8724,N_5287,N_4566);
or U8725 (N_8725,N_5405,N_3901);
xor U8726 (N_8726,N_3299,N_3670);
nor U8727 (N_8727,N_4575,N_5900);
xnor U8728 (N_8728,N_4239,N_4515);
and U8729 (N_8729,N_3041,N_3061);
and U8730 (N_8730,N_4124,N_5589);
nor U8731 (N_8731,N_5062,N_5128);
and U8732 (N_8732,N_5715,N_5135);
nand U8733 (N_8733,N_5294,N_3128);
and U8734 (N_8734,N_3533,N_5903);
nor U8735 (N_8735,N_3285,N_4624);
or U8736 (N_8736,N_4640,N_3735);
and U8737 (N_8737,N_4464,N_4757);
nor U8738 (N_8738,N_5879,N_4905);
nor U8739 (N_8739,N_3570,N_4132);
nand U8740 (N_8740,N_5401,N_3156);
nor U8741 (N_8741,N_3437,N_5876);
nand U8742 (N_8742,N_4179,N_5310);
nor U8743 (N_8743,N_5532,N_3691);
nor U8744 (N_8744,N_4139,N_5737);
nand U8745 (N_8745,N_3229,N_4915);
nor U8746 (N_8746,N_4403,N_4738);
nor U8747 (N_8747,N_4189,N_4454);
xnor U8748 (N_8748,N_3411,N_3936);
nand U8749 (N_8749,N_4807,N_5073);
xor U8750 (N_8750,N_5429,N_5124);
xnor U8751 (N_8751,N_5715,N_3639);
xnor U8752 (N_8752,N_5567,N_4580);
xor U8753 (N_8753,N_3537,N_3849);
or U8754 (N_8754,N_5894,N_4125);
nor U8755 (N_8755,N_3702,N_3140);
nor U8756 (N_8756,N_4464,N_5250);
or U8757 (N_8757,N_4113,N_3198);
xnor U8758 (N_8758,N_5256,N_5807);
nand U8759 (N_8759,N_4040,N_5400);
nor U8760 (N_8760,N_3348,N_5095);
nor U8761 (N_8761,N_5497,N_5682);
or U8762 (N_8762,N_4319,N_5931);
or U8763 (N_8763,N_3105,N_3942);
nand U8764 (N_8764,N_3647,N_4205);
nand U8765 (N_8765,N_4597,N_5510);
nand U8766 (N_8766,N_5282,N_3394);
nor U8767 (N_8767,N_5395,N_5178);
nand U8768 (N_8768,N_4266,N_3281);
nand U8769 (N_8769,N_5425,N_3051);
nor U8770 (N_8770,N_5058,N_4491);
xor U8771 (N_8771,N_3280,N_5010);
or U8772 (N_8772,N_4466,N_3133);
xnor U8773 (N_8773,N_5069,N_4744);
and U8774 (N_8774,N_5935,N_4184);
xor U8775 (N_8775,N_3727,N_5039);
or U8776 (N_8776,N_3744,N_3332);
xor U8777 (N_8777,N_4213,N_4707);
nand U8778 (N_8778,N_5043,N_5383);
and U8779 (N_8779,N_4343,N_5554);
or U8780 (N_8780,N_3133,N_3372);
nand U8781 (N_8781,N_5174,N_3755);
xnor U8782 (N_8782,N_3926,N_3947);
xor U8783 (N_8783,N_3500,N_4670);
nor U8784 (N_8784,N_3674,N_4575);
xor U8785 (N_8785,N_3473,N_3933);
or U8786 (N_8786,N_5740,N_5439);
or U8787 (N_8787,N_5656,N_4760);
nor U8788 (N_8788,N_4598,N_4432);
or U8789 (N_8789,N_5438,N_5215);
or U8790 (N_8790,N_4794,N_3583);
xor U8791 (N_8791,N_5123,N_4772);
xnor U8792 (N_8792,N_4874,N_5448);
nor U8793 (N_8793,N_3750,N_3580);
nand U8794 (N_8794,N_5782,N_3101);
nor U8795 (N_8795,N_4155,N_5051);
nand U8796 (N_8796,N_3260,N_4012);
or U8797 (N_8797,N_4710,N_4544);
and U8798 (N_8798,N_3333,N_5078);
nor U8799 (N_8799,N_3068,N_3242);
nor U8800 (N_8800,N_4838,N_5703);
or U8801 (N_8801,N_5930,N_3199);
xor U8802 (N_8802,N_3589,N_4974);
nor U8803 (N_8803,N_3360,N_3445);
or U8804 (N_8804,N_4426,N_3821);
or U8805 (N_8805,N_3157,N_4978);
or U8806 (N_8806,N_4257,N_4628);
nor U8807 (N_8807,N_4632,N_3758);
nor U8808 (N_8808,N_5953,N_4971);
nor U8809 (N_8809,N_4913,N_5540);
nand U8810 (N_8810,N_3898,N_4214);
xor U8811 (N_8811,N_4731,N_3177);
and U8812 (N_8812,N_3293,N_3685);
nor U8813 (N_8813,N_4416,N_4034);
xor U8814 (N_8814,N_3189,N_3648);
nand U8815 (N_8815,N_3893,N_3281);
and U8816 (N_8816,N_5376,N_4285);
and U8817 (N_8817,N_4373,N_5073);
or U8818 (N_8818,N_4319,N_5119);
or U8819 (N_8819,N_3670,N_3988);
nand U8820 (N_8820,N_3548,N_3391);
nor U8821 (N_8821,N_4097,N_5439);
nand U8822 (N_8822,N_5986,N_5997);
and U8823 (N_8823,N_4792,N_3511);
xor U8824 (N_8824,N_3738,N_4938);
nor U8825 (N_8825,N_3102,N_5226);
xor U8826 (N_8826,N_5340,N_3449);
nor U8827 (N_8827,N_4130,N_5250);
xor U8828 (N_8828,N_4949,N_3346);
or U8829 (N_8829,N_5823,N_4636);
xor U8830 (N_8830,N_5855,N_5029);
and U8831 (N_8831,N_4645,N_5890);
and U8832 (N_8832,N_4220,N_4818);
or U8833 (N_8833,N_5611,N_3229);
xor U8834 (N_8834,N_3871,N_4421);
xor U8835 (N_8835,N_4816,N_4421);
or U8836 (N_8836,N_4723,N_5651);
or U8837 (N_8837,N_4659,N_3521);
xor U8838 (N_8838,N_4733,N_4374);
and U8839 (N_8839,N_3765,N_4380);
or U8840 (N_8840,N_3597,N_4083);
nand U8841 (N_8841,N_3943,N_4931);
nand U8842 (N_8842,N_4053,N_4273);
or U8843 (N_8843,N_5531,N_3965);
and U8844 (N_8844,N_5907,N_3869);
and U8845 (N_8845,N_3147,N_3313);
and U8846 (N_8846,N_4481,N_5873);
and U8847 (N_8847,N_3084,N_3266);
xnor U8848 (N_8848,N_3424,N_4425);
or U8849 (N_8849,N_5933,N_4964);
nor U8850 (N_8850,N_3271,N_5663);
and U8851 (N_8851,N_3688,N_3859);
nor U8852 (N_8852,N_3905,N_5108);
nor U8853 (N_8853,N_5798,N_3548);
nor U8854 (N_8854,N_5487,N_5099);
nor U8855 (N_8855,N_3463,N_5099);
or U8856 (N_8856,N_5053,N_5282);
nand U8857 (N_8857,N_4985,N_5226);
xor U8858 (N_8858,N_4840,N_4727);
or U8859 (N_8859,N_4444,N_4312);
nand U8860 (N_8860,N_4944,N_5306);
nand U8861 (N_8861,N_3665,N_5317);
or U8862 (N_8862,N_3828,N_3510);
nand U8863 (N_8863,N_5646,N_3389);
nor U8864 (N_8864,N_4814,N_3167);
or U8865 (N_8865,N_5311,N_3946);
xnor U8866 (N_8866,N_4114,N_5704);
nor U8867 (N_8867,N_3293,N_4290);
nand U8868 (N_8868,N_5773,N_5319);
and U8869 (N_8869,N_4009,N_4895);
and U8870 (N_8870,N_5291,N_3182);
nor U8871 (N_8871,N_5209,N_3962);
xor U8872 (N_8872,N_5974,N_4097);
xor U8873 (N_8873,N_4476,N_5639);
nand U8874 (N_8874,N_5607,N_3623);
nor U8875 (N_8875,N_4542,N_4321);
or U8876 (N_8876,N_5268,N_5262);
and U8877 (N_8877,N_3780,N_4462);
nor U8878 (N_8878,N_3088,N_5864);
and U8879 (N_8879,N_3735,N_4115);
or U8880 (N_8880,N_3730,N_4342);
nor U8881 (N_8881,N_4507,N_5092);
or U8882 (N_8882,N_5920,N_5664);
and U8883 (N_8883,N_5768,N_4986);
nand U8884 (N_8884,N_4344,N_4922);
and U8885 (N_8885,N_4680,N_4722);
and U8886 (N_8886,N_4598,N_4918);
or U8887 (N_8887,N_4373,N_3204);
or U8888 (N_8888,N_5968,N_3323);
nor U8889 (N_8889,N_4809,N_3723);
nor U8890 (N_8890,N_4416,N_3154);
and U8891 (N_8891,N_3914,N_5121);
or U8892 (N_8892,N_4017,N_4259);
xnor U8893 (N_8893,N_5175,N_3574);
and U8894 (N_8894,N_3209,N_5949);
and U8895 (N_8895,N_5309,N_3145);
nand U8896 (N_8896,N_3250,N_3388);
or U8897 (N_8897,N_5011,N_4316);
xnor U8898 (N_8898,N_4854,N_4483);
nand U8899 (N_8899,N_3177,N_4974);
nor U8900 (N_8900,N_5809,N_5785);
nor U8901 (N_8901,N_5632,N_4967);
nor U8902 (N_8902,N_3204,N_4758);
and U8903 (N_8903,N_3172,N_3761);
or U8904 (N_8904,N_4170,N_3047);
nand U8905 (N_8905,N_4560,N_4148);
nand U8906 (N_8906,N_3734,N_4640);
or U8907 (N_8907,N_3330,N_4404);
nor U8908 (N_8908,N_4565,N_3020);
xnor U8909 (N_8909,N_5179,N_3134);
xor U8910 (N_8910,N_4396,N_4311);
nor U8911 (N_8911,N_4551,N_5123);
or U8912 (N_8912,N_4405,N_5682);
or U8913 (N_8913,N_5299,N_4202);
nand U8914 (N_8914,N_3378,N_4181);
nand U8915 (N_8915,N_4845,N_5751);
xnor U8916 (N_8916,N_5714,N_3513);
nand U8917 (N_8917,N_4969,N_3598);
or U8918 (N_8918,N_3798,N_5069);
nor U8919 (N_8919,N_4113,N_3879);
xor U8920 (N_8920,N_5755,N_4102);
xnor U8921 (N_8921,N_4605,N_3630);
or U8922 (N_8922,N_3060,N_5052);
nand U8923 (N_8923,N_3904,N_3954);
xor U8924 (N_8924,N_5507,N_3088);
or U8925 (N_8925,N_3721,N_4729);
nand U8926 (N_8926,N_4498,N_3487);
xor U8927 (N_8927,N_5993,N_5846);
xnor U8928 (N_8928,N_3552,N_3674);
or U8929 (N_8929,N_4514,N_5632);
or U8930 (N_8930,N_3698,N_3364);
nor U8931 (N_8931,N_5264,N_5234);
nand U8932 (N_8932,N_3559,N_4373);
or U8933 (N_8933,N_5571,N_4446);
or U8934 (N_8934,N_3397,N_3442);
xor U8935 (N_8935,N_4675,N_5201);
nand U8936 (N_8936,N_3636,N_4838);
xor U8937 (N_8937,N_4313,N_4676);
and U8938 (N_8938,N_3727,N_5818);
nand U8939 (N_8939,N_5318,N_5056);
or U8940 (N_8940,N_3816,N_5409);
and U8941 (N_8941,N_4035,N_3645);
nor U8942 (N_8942,N_3732,N_3026);
and U8943 (N_8943,N_5226,N_4295);
xnor U8944 (N_8944,N_4049,N_3767);
nor U8945 (N_8945,N_4455,N_4093);
and U8946 (N_8946,N_3696,N_3311);
nor U8947 (N_8947,N_4439,N_4009);
xnor U8948 (N_8948,N_5658,N_5352);
xor U8949 (N_8949,N_3671,N_3122);
nand U8950 (N_8950,N_4962,N_5689);
or U8951 (N_8951,N_4965,N_5442);
or U8952 (N_8952,N_5229,N_5273);
nand U8953 (N_8953,N_3318,N_5316);
xnor U8954 (N_8954,N_3953,N_5719);
and U8955 (N_8955,N_4919,N_5682);
xnor U8956 (N_8956,N_5721,N_3282);
and U8957 (N_8957,N_4507,N_4792);
and U8958 (N_8958,N_4060,N_4669);
nand U8959 (N_8959,N_5678,N_4211);
xor U8960 (N_8960,N_3880,N_5419);
xnor U8961 (N_8961,N_5956,N_3368);
nor U8962 (N_8962,N_5403,N_4927);
xnor U8963 (N_8963,N_5904,N_5390);
nand U8964 (N_8964,N_5044,N_3899);
xor U8965 (N_8965,N_5419,N_5120);
or U8966 (N_8966,N_3383,N_5263);
nor U8967 (N_8967,N_3191,N_5432);
xnor U8968 (N_8968,N_4512,N_5382);
and U8969 (N_8969,N_4280,N_4635);
nand U8970 (N_8970,N_5544,N_3142);
nor U8971 (N_8971,N_5132,N_3683);
nand U8972 (N_8972,N_5796,N_5281);
or U8973 (N_8973,N_4487,N_4905);
and U8974 (N_8974,N_5805,N_5609);
nand U8975 (N_8975,N_4588,N_5963);
nor U8976 (N_8976,N_4714,N_4449);
nor U8977 (N_8977,N_4921,N_5365);
nand U8978 (N_8978,N_3183,N_4241);
nor U8979 (N_8979,N_5368,N_4240);
and U8980 (N_8980,N_5178,N_5955);
and U8981 (N_8981,N_5066,N_4641);
nand U8982 (N_8982,N_3573,N_5465);
nand U8983 (N_8983,N_3773,N_5039);
nor U8984 (N_8984,N_4342,N_4011);
nand U8985 (N_8985,N_5562,N_3023);
xor U8986 (N_8986,N_3941,N_3358);
or U8987 (N_8987,N_4767,N_4792);
and U8988 (N_8988,N_4852,N_3496);
and U8989 (N_8989,N_3924,N_4841);
and U8990 (N_8990,N_4062,N_4194);
xnor U8991 (N_8991,N_3554,N_5520);
nor U8992 (N_8992,N_5571,N_5334);
and U8993 (N_8993,N_3369,N_5896);
nor U8994 (N_8994,N_3071,N_4528);
and U8995 (N_8995,N_3406,N_4501);
or U8996 (N_8996,N_3105,N_3078);
xor U8997 (N_8997,N_4165,N_4400);
and U8998 (N_8998,N_5164,N_4585);
nor U8999 (N_8999,N_5503,N_4584);
xor U9000 (N_9000,N_8350,N_8250);
or U9001 (N_9001,N_7229,N_6054);
nor U9002 (N_9002,N_7576,N_8451);
and U9003 (N_9003,N_8269,N_6277);
or U9004 (N_9004,N_6032,N_8032);
or U9005 (N_9005,N_6100,N_6015);
xor U9006 (N_9006,N_7345,N_6504);
and U9007 (N_9007,N_7362,N_8105);
nand U9008 (N_9008,N_8114,N_8015);
nand U9009 (N_9009,N_7269,N_8467);
nor U9010 (N_9010,N_8500,N_7129);
nand U9011 (N_9011,N_7389,N_7766);
and U9012 (N_9012,N_8836,N_8283);
or U9013 (N_9013,N_7147,N_6025);
and U9014 (N_9014,N_6718,N_8327);
xnor U9015 (N_9015,N_6543,N_7690);
nand U9016 (N_9016,N_8479,N_6669);
xnor U9017 (N_9017,N_6686,N_7169);
or U9018 (N_9018,N_6722,N_7500);
or U9019 (N_9019,N_7802,N_8165);
or U9020 (N_9020,N_7781,N_7672);
or U9021 (N_9021,N_7971,N_6119);
or U9022 (N_9022,N_7009,N_8781);
or U9023 (N_9023,N_8865,N_8139);
nand U9024 (N_9024,N_7928,N_8496);
and U9025 (N_9025,N_7652,N_6252);
xnor U9026 (N_9026,N_8773,N_7546);
and U9027 (N_9027,N_7022,N_6327);
xnor U9028 (N_9028,N_8675,N_8756);
xnor U9029 (N_9029,N_8529,N_6339);
and U9030 (N_9030,N_6187,N_7028);
nor U9031 (N_9031,N_6217,N_8372);
nor U9032 (N_9032,N_6180,N_6205);
and U9033 (N_9033,N_8875,N_6532);
nand U9034 (N_9034,N_6192,N_6797);
nand U9035 (N_9035,N_7912,N_7883);
nor U9036 (N_9036,N_7869,N_6198);
xnor U9037 (N_9037,N_6679,N_7836);
nor U9038 (N_9038,N_7418,N_6535);
nor U9039 (N_9039,N_6261,N_6745);
and U9040 (N_9040,N_6943,N_6562);
and U9041 (N_9041,N_7972,N_6492);
nor U9042 (N_9042,N_8866,N_8960);
and U9043 (N_9043,N_6442,N_7918);
and U9044 (N_9044,N_7800,N_8971);
nand U9045 (N_9045,N_7906,N_6857);
xnor U9046 (N_9046,N_6823,N_8491);
nor U9047 (N_9047,N_8279,N_7155);
nand U9048 (N_9048,N_8825,N_7215);
nor U9049 (N_9049,N_7102,N_7320);
nand U9050 (N_9050,N_6421,N_6378);
or U9051 (N_9051,N_8562,N_7412);
nor U9052 (N_9052,N_8889,N_6037);
nand U9053 (N_9053,N_8317,N_8024);
xnor U9054 (N_9054,N_6239,N_7748);
and U9055 (N_9055,N_6077,N_8134);
or U9056 (N_9056,N_7183,N_7166);
nand U9057 (N_9057,N_8962,N_6462);
and U9058 (N_9058,N_8247,N_6559);
or U9059 (N_9059,N_8427,N_8457);
xor U9060 (N_9060,N_7553,N_7054);
and U9061 (N_9061,N_6073,N_6185);
nor U9062 (N_9062,N_8205,N_6634);
nand U9063 (N_9063,N_8603,N_8633);
or U9064 (N_9064,N_7019,N_6507);
nand U9065 (N_9065,N_7644,N_7325);
nor U9066 (N_9066,N_7646,N_6712);
and U9067 (N_9067,N_7816,N_8109);
nor U9068 (N_9068,N_8840,N_6747);
or U9069 (N_9069,N_6542,N_6994);
nor U9070 (N_9070,N_7667,N_7225);
nor U9071 (N_9071,N_8503,N_6652);
and U9072 (N_9072,N_7932,N_6092);
or U9073 (N_9073,N_8371,N_6461);
nor U9074 (N_9074,N_8623,N_8740);
or U9075 (N_9075,N_8156,N_7421);
and U9076 (N_9076,N_7894,N_7872);
or U9077 (N_9077,N_7350,N_6911);
and U9078 (N_9078,N_6232,N_6915);
and U9079 (N_9079,N_8657,N_7235);
xnor U9080 (N_9080,N_6995,N_7167);
and U9081 (N_9081,N_8604,N_8648);
or U9082 (N_9082,N_8295,N_6183);
nand U9083 (N_9083,N_7643,N_8915);
or U9084 (N_9084,N_6146,N_8449);
nand U9085 (N_9085,N_6643,N_7112);
or U9086 (N_9086,N_6052,N_7823);
xor U9087 (N_9087,N_8418,N_8509);
and U9088 (N_9088,N_7631,N_6017);
nor U9089 (N_9089,N_8460,N_7964);
or U9090 (N_9090,N_8140,N_6453);
nand U9091 (N_9091,N_8937,N_6431);
nand U9092 (N_9092,N_8454,N_6880);
or U9093 (N_9093,N_6364,N_6821);
xnor U9094 (N_9094,N_7346,N_6330);
nor U9095 (N_9095,N_7716,N_6288);
nand U9096 (N_9096,N_6499,N_6920);
nand U9097 (N_9097,N_8211,N_6649);
xor U9098 (N_9098,N_8301,N_8616);
xor U9099 (N_9099,N_7388,N_8017);
nand U9100 (N_9100,N_8796,N_7550);
and U9101 (N_9101,N_6233,N_7228);
nor U9102 (N_9102,N_8123,N_7387);
or U9103 (N_9103,N_8369,N_6979);
xor U9104 (N_9104,N_6237,N_8887);
nand U9105 (N_9105,N_8396,N_8334);
xnor U9106 (N_9106,N_6897,N_7923);
or U9107 (N_9107,N_7444,N_7568);
nand U9108 (N_9108,N_6637,N_8236);
xnor U9109 (N_9109,N_6043,N_6283);
or U9110 (N_9110,N_8606,N_6488);
and U9111 (N_9111,N_8760,N_6206);
nor U9112 (N_9112,N_8768,N_7980);
and U9113 (N_9113,N_8929,N_8989);
nor U9114 (N_9114,N_6020,N_6827);
and U9115 (N_9115,N_6791,N_8585);
nand U9116 (N_9116,N_8986,N_8353);
nand U9117 (N_9117,N_8904,N_8444);
or U9118 (N_9118,N_7740,N_7828);
nor U9119 (N_9119,N_6299,N_6901);
xnor U9120 (N_9120,N_7523,N_8080);
xnor U9121 (N_9121,N_6810,N_8203);
or U9122 (N_9122,N_6362,N_8908);
or U9123 (N_9123,N_7011,N_6876);
nand U9124 (N_9124,N_7601,N_6298);
nor U9125 (N_9125,N_7850,N_6370);
xor U9126 (N_9126,N_8160,N_8905);
nand U9127 (N_9127,N_7124,N_8854);
nor U9128 (N_9128,N_6296,N_8034);
or U9129 (N_9129,N_8046,N_6372);
and U9130 (N_9130,N_7001,N_8645);
nand U9131 (N_9131,N_6270,N_8378);
and U9132 (N_9132,N_6227,N_8423);
xnor U9133 (N_9133,N_6272,N_8763);
nand U9134 (N_9134,N_6204,N_7283);
and U9135 (N_9135,N_8748,N_6142);
nand U9136 (N_9136,N_7603,N_6764);
xor U9137 (N_9137,N_6411,N_7571);
and U9138 (N_9138,N_7381,N_6965);
and U9139 (N_9139,N_6934,N_7433);
and U9140 (N_9140,N_6361,N_6385);
nor U9141 (N_9141,N_6700,N_6799);
xor U9142 (N_9142,N_6127,N_6717);
nor U9143 (N_9143,N_8726,N_8697);
nor U9144 (N_9144,N_6026,N_7371);
and U9145 (N_9145,N_7954,N_7795);
nand U9146 (N_9146,N_6804,N_6075);
or U9147 (N_9147,N_6592,N_8992);
nor U9148 (N_9148,N_8701,N_7525);
nor U9149 (N_9149,N_6910,N_8827);
nor U9150 (N_9150,N_7236,N_8425);
xnor U9151 (N_9151,N_8492,N_6567);
or U9152 (N_9152,N_8924,N_8856);
and U9153 (N_9153,N_7989,N_6016);
nand U9154 (N_9154,N_8389,N_6891);
xnor U9155 (N_9155,N_6523,N_8534);
and U9156 (N_9156,N_8043,N_8448);
nand U9157 (N_9157,N_6003,N_8931);
nand U9158 (N_9158,N_8344,N_7605);
nor U9159 (N_9159,N_7488,N_6501);
nand U9160 (N_9160,N_8366,N_7046);
and U9161 (N_9161,N_7521,N_6159);
or U9162 (N_9162,N_7319,N_7509);
and U9163 (N_9163,N_8209,N_8558);
xor U9164 (N_9164,N_8006,N_7351);
and U9165 (N_9165,N_7223,N_7305);
and U9166 (N_9166,N_7889,N_6993);
xnor U9167 (N_9167,N_8852,N_7222);
and U9168 (N_9168,N_8035,N_8438);
and U9169 (N_9169,N_6096,N_7151);
xnor U9170 (N_9170,N_7255,N_7335);
or U9171 (N_9171,N_7272,N_7837);
nand U9172 (N_9172,N_8195,N_8627);
or U9173 (N_9173,N_8437,N_6220);
nor U9174 (N_9174,N_6692,N_8517);
or U9175 (N_9175,N_6030,N_6400);
xnor U9176 (N_9176,N_8741,N_6992);
and U9177 (N_9177,N_8108,N_6269);
or U9178 (N_9178,N_8288,N_6267);
nand U9179 (N_9179,N_8498,N_6439);
nand U9180 (N_9180,N_8587,N_7678);
nor U9181 (N_9181,N_6463,N_7149);
or U9182 (N_9182,N_8672,N_6295);
xnor U9183 (N_9183,N_8646,N_6693);
xor U9184 (N_9184,N_7237,N_8253);
and U9185 (N_9185,N_8490,N_8619);
or U9186 (N_9186,N_7031,N_7827);
or U9187 (N_9187,N_7432,N_7710);
xnor U9188 (N_9188,N_6447,N_6755);
xor U9189 (N_9189,N_8696,N_8494);
and U9190 (N_9190,N_8313,N_7990);
nand U9191 (N_9191,N_6561,N_7522);
xor U9192 (N_9192,N_6308,N_8365);
nand U9193 (N_9193,N_6964,N_6599);
nor U9194 (N_9194,N_7718,N_7400);
xor U9195 (N_9195,N_6815,N_8663);
and U9196 (N_9196,N_7734,N_8167);
or U9197 (N_9197,N_8636,N_6218);
and U9198 (N_9198,N_7688,N_8426);
xor U9199 (N_9199,N_8308,N_7231);
nand U9200 (N_9200,N_7640,N_6028);
and U9201 (N_9201,N_6429,N_8634);
and U9202 (N_9202,N_8470,N_7664);
xor U9203 (N_9203,N_8319,N_7306);
nand U9204 (N_9204,N_8343,N_8475);
or U9205 (N_9205,N_7462,N_8596);
xor U9206 (N_9206,N_6707,N_8182);
and U9207 (N_9207,N_8694,N_7778);
nand U9208 (N_9208,N_8801,N_7287);
and U9209 (N_9209,N_8306,N_6107);
nand U9210 (N_9210,N_6551,N_7704);
nor U9211 (N_9211,N_8216,N_8525);
nand U9212 (N_9212,N_8590,N_7103);
nand U9213 (N_9213,N_6161,N_6770);
nor U9214 (N_9214,N_7693,N_6841);
nor U9215 (N_9215,N_8972,N_7020);
nor U9216 (N_9216,N_7244,N_7238);
nor U9217 (N_9217,N_7402,N_7949);
nor U9218 (N_9218,N_8477,N_6657);
nor U9219 (N_9219,N_8333,N_6720);
nand U9220 (N_9220,N_6319,N_8745);
or U9221 (N_9221,N_8413,N_6777);
and U9222 (N_9222,N_6397,N_7891);
and U9223 (N_9223,N_8499,N_7963);
nand U9224 (N_9224,N_7468,N_6409);
xor U9225 (N_9225,N_6489,N_6642);
and U9226 (N_9226,N_8052,N_6552);
nor U9227 (N_9227,N_6200,N_6886);
nand U9228 (N_9228,N_7006,N_7145);
nor U9229 (N_9229,N_6578,N_8917);
nor U9230 (N_9230,N_6487,N_7116);
nand U9231 (N_9231,N_8092,N_6098);
and U9232 (N_9232,N_8169,N_6022);
nand U9233 (N_9233,N_8660,N_8450);
nor U9234 (N_9234,N_7526,N_6219);
nand U9235 (N_9235,N_8273,N_7880);
and U9236 (N_9236,N_8664,N_7556);
or U9237 (N_9237,N_7258,N_6105);
xor U9238 (N_9238,N_7761,N_7623);
xnor U9239 (N_9239,N_6293,N_8898);
nand U9240 (N_9240,N_8286,N_7896);
or U9241 (N_9241,N_7334,N_7398);
or U9242 (N_9242,N_7057,N_6033);
or U9243 (N_9243,N_8967,N_6544);
xnor U9244 (N_9244,N_8089,N_7240);
and U9245 (N_9245,N_7375,N_7015);
nand U9246 (N_9246,N_6511,N_6613);
xor U9247 (N_9247,N_8508,N_7437);
nand U9248 (N_9248,N_8227,N_8051);
or U9249 (N_9249,N_8601,N_6338);
and U9250 (N_9250,N_6665,N_7774);
xor U9251 (N_9251,N_6224,N_6611);
xor U9252 (N_9252,N_7327,N_8897);
nor U9253 (N_9253,N_8806,N_8863);
or U9254 (N_9254,N_7679,N_8647);
xnor U9255 (N_9255,N_8462,N_7805);
xor U9256 (N_9256,N_7190,N_8443);
xor U9257 (N_9257,N_7796,N_8698);
nand U9258 (N_9258,N_8709,N_6469);
or U9259 (N_9259,N_7731,N_7074);
xnor U9260 (N_9260,N_8030,N_7227);
or U9261 (N_9261,N_7380,N_7430);
nor U9262 (N_9262,N_6318,N_6721);
nand U9263 (N_9263,N_7898,N_6001);
nand U9264 (N_9264,N_7621,N_7807);
and U9265 (N_9265,N_6460,N_8982);
or U9266 (N_9266,N_8932,N_6816);
or U9267 (N_9267,N_7379,N_6866);
and U9268 (N_9268,N_7144,N_6667);
nand U9269 (N_9269,N_7461,N_8577);
xor U9270 (N_9270,N_8691,N_7752);
xor U9271 (N_9271,N_7048,N_7728);
nor U9272 (N_9272,N_8082,N_7552);
and U9273 (N_9273,N_8000,N_6769);
and U9274 (N_9274,N_6622,N_8703);
xnor U9275 (N_9275,N_8560,N_7174);
nor U9276 (N_9276,N_7133,N_8859);
xor U9277 (N_9277,N_7966,N_8374);
xnor U9278 (N_9278,N_8686,N_6007);
xnor U9279 (N_9279,N_8210,N_6486);
nand U9280 (N_9280,N_7797,N_8652);
nor U9281 (N_9281,N_7573,N_8925);
xor U9282 (N_9282,N_6112,N_6768);
and U9283 (N_9283,N_7098,N_6527);
nor U9284 (N_9284,N_7447,N_8916);
or U9285 (N_9285,N_6434,N_6849);
nand U9286 (N_9286,N_8465,N_6895);
nor U9287 (N_9287,N_8593,N_6870);
nor U9288 (N_9288,N_8910,N_8208);
and U9289 (N_9289,N_8202,N_8348);
nor U9290 (N_9290,N_6675,N_6343);
or U9291 (N_9291,N_7114,N_6391);
nand U9292 (N_9292,N_7329,N_6059);
nor U9293 (N_9293,N_6687,N_8324);
and U9294 (N_9294,N_8695,N_6312);
xnor U9295 (N_9295,N_7354,N_8455);
nand U9296 (N_9296,N_7535,N_8817);
or U9297 (N_9297,N_6354,N_8018);
and U9298 (N_9298,N_8441,N_8835);
nand U9299 (N_9299,N_7405,N_7036);
nand U9300 (N_9300,N_8752,N_7777);
and U9301 (N_9301,N_8799,N_7602);
and U9302 (N_9302,N_8487,N_6305);
nand U9303 (N_9303,N_8435,N_8482);
or U9304 (N_9304,N_6458,N_8255);
nor U9305 (N_9305,N_6207,N_7051);
or U9306 (N_9306,N_6249,N_7491);
xor U9307 (N_9307,N_8238,N_8757);
and U9308 (N_9308,N_6909,N_6145);
and U9309 (N_9309,N_7886,N_7042);
xnor U9310 (N_9310,N_6210,N_6347);
nor U9311 (N_9311,N_8037,N_7876);
or U9312 (N_9312,N_6526,N_7452);
and U9313 (N_9313,N_6733,N_7451);
xor U9314 (N_9314,N_7780,N_6348);
and U9315 (N_9315,N_7624,N_7703);
or U9316 (N_9316,N_8977,N_6749);
and U9317 (N_9317,N_6229,N_8519);
or U9318 (N_9318,N_6684,N_8784);
xor U9319 (N_9319,N_8922,N_8266);
nand U9320 (N_9320,N_6029,N_6147);
nand U9321 (N_9321,N_7086,N_8407);
nor U9322 (N_9322,N_6111,N_8416);
nand U9323 (N_9323,N_7698,N_6872);
and U9324 (N_9324,N_6211,N_8053);
nand U9325 (N_9325,N_7749,N_6231);
nand U9326 (N_9326,N_6472,N_7120);
nor U9327 (N_9327,N_7712,N_8010);
or U9328 (N_9328,N_7392,N_6774);
nand U9329 (N_9329,N_6408,N_6548);
and U9330 (N_9330,N_7077,N_8004);
and U9331 (N_9331,N_6282,N_6120);
or U9332 (N_9332,N_6573,N_8552);
nand U9333 (N_9333,N_7296,N_8822);
and U9334 (N_9334,N_8063,N_6809);
nand U9335 (N_9335,N_7295,N_6844);
nand U9336 (N_9336,N_6351,N_6925);
nor U9337 (N_9337,N_8678,N_6129);
nand U9338 (N_9338,N_8945,N_8328);
nand U9339 (N_9339,N_7594,N_7927);
nand U9340 (N_9340,N_7733,N_7950);
nor U9341 (N_9341,N_6094,N_6949);
xor U9342 (N_9342,N_7600,N_6663);
or U9343 (N_9343,N_6625,N_6457);
and U9344 (N_9344,N_7300,N_7165);
nand U9345 (N_9345,N_6672,N_8064);
nor U9346 (N_9346,N_6884,N_6475);
and U9347 (N_9347,N_6176,N_6802);
or U9348 (N_9348,N_6572,N_8198);
xor U9349 (N_9349,N_8440,N_7383);
and U9350 (N_9350,N_7441,N_8339);
xnor U9351 (N_9351,N_7221,N_8829);
and U9352 (N_9352,N_6750,N_7656);
xor U9353 (N_9353,N_8938,N_7588);
or U9354 (N_9354,N_6440,N_6403);
nand U9355 (N_9355,N_6654,N_6290);
xnor U9356 (N_9356,N_8260,N_7899);
and U9357 (N_9357,N_8088,N_7315);
xnor U9358 (N_9358,N_6832,N_7847);
xor U9359 (N_9359,N_7391,N_6130);
nand U9360 (N_9360,N_6728,N_7176);
xnor U9361 (N_9361,N_7921,N_7893);
nand U9362 (N_9362,N_7291,N_6826);
nor U9363 (N_9363,N_7328,N_6375);
nor U9364 (N_9364,N_7649,N_7497);
xnor U9365 (N_9365,N_7393,N_6365);
and U9366 (N_9366,N_8567,N_8191);
xnor U9367 (N_9367,N_6328,N_7413);
nand U9368 (N_9368,N_8254,N_8857);
xnor U9369 (N_9369,N_8252,N_7996);
xnor U9370 (N_9370,N_7479,N_7445);
or U9371 (N_9371,N_6240,N_7423);
nand U9372 (N_9372,N_8087,N_6795);
and U9373 (N_9373,N_8300,N_8666);
or U9374 (N_9374,N_8595,N_6674);
xnor U9375 (N_9375,N_7615,N_8941);
xor U9376 (N_9376,N_7070,N_7720);
or U9377 (N_9377,N_6436,N_8096);
xor U9378 (N_9378,N_8436,N_7513);
and U9379 (N_9379,N_8994,N_8656);
nor U9380 (N_9380,N_8239,N_6739);
and U9381 (N_9381,N_7657,N_8766);
nor U9382 (N_9382,N_7763,N_6326);
and U9383 (N_9383,N_7881,N_6174);
nor U9384 (N_9384,N_6301,N_7349);
or U9385 (N_9385,N_7211,N_6279);
xnor U9386 (N_9386,N_8862,N_8998);
xor U9387 (N_9387,N_6478,N_6182);
or U9388 (N_9388,N_7955,N_8262);
xnor U9389 (N_9389,N_6208,N_8136);
xor U9390 (N_9390,N_6697,N_8544);
and U9391 (N_9391,N_8589,N_7463);
or U9392 (N_9392,N_8345,N_8535);
or U9393 (N_9393,N_7845,N_7683);
nor U9394 (N_9394,N_8047,N_6968);
nand U9395 (N_9395,N_8207,N_7822);
nor U9396 (N_9396,N_8023,N_6345);
or U9397 (N_9397,N_6757,N_7887);
or U9398 (N_9398,N_8119,N_7115);
and U9399 (N_9399,N_8618,N_6215);
xnor U9400 (N_9400,N_7093,N_8846);
nor U9401 (N_9401,N_8272,N_7981);
or U9402 (N_9402,N_7788,N_7355);
nand U9403 (N_9403,N_6248,N_7076);
xnor U9404 (N_9404,N_7161,N_8145);
and U9405 (N_9405,N_6137,N_8753);
and U9406 (N_9406,N_6256,N_8081);
and U9407 (N_9407,N_8890,N_7162);
xnor U9408 (N_9408,N_8810,N_6353);
and U9409 (N_9409,N_6243,N_6648);
or U9410 (N_9410,N_7685,N_8735);
xor U9411 (N_9411,N_7204,N_6601);
nor U9412 (N_9412,N_8742,N_6235);
xnor U9413 (N_9413,N_8453,N_6678);
and U9414 (N_9414,N_6761,N_7849);
xnor U9415 (N_9415,N_8923,N_6683);
or U9416 (N_9416,N_8800,N_8321);
and U9417 (N_9417,N_8097,N_6735);
nand U9418 (N_9418,N_6989,N_8659);
nand U9419 (N_9419,N_8993,N_7330);
xnor U9420 (N_9420,N_7681,N_7750);
nand U9421 (N_9421,N_6406,N_6039);
and U9422 (N_9422,N_7201,N_8724);
nor U9423 (N_9423,N_7234,N_7986);
or U9424 (N_9424,N_8429,N_7455);
nand U9425 (N_9425,N_6709,N_7559);
nor U9426 (N_9426,N_8792,N_7755);
or U9427 (N_9427,N_8683,N_7722);
and U9428 (N_9428,N_6134,N_8804);
or U9429 (N_9429,N_6333,N_8232);
or U9430 (N_9430,N_6024,N_6845);
nand U9431 (N_9431,N_7052,N_7645);
or U9432 (N_9432,N_7261,N_7713);
nor U9433 (N_9433,N_7738,N_8902);
and U9434 (N_9434,N_8758,N_6976);
nor U9435 (N_9435,N_8653,N_8011);
nand U9436 (N_9436,N_8769,N_6814);
or U9437 (N_9437,N_6600,N_7439);
nand U9438 (N_9438,N_8845,N_6784);
or U9439 (N_9439,N_8040,N_6263);
nand U9440 (N_9440,N_8555,N_7040);
nand U9441 (N_9441,N_8877,N_6947);
nand U9442 (N_9442,N_7002,N_8775);
nand U9443 (N_9443,N_6432,N_6099);
or U9444 (N_9444,N_7721,N_6490);
and U9445 (N_9445,N_7801,N_8391);
nand U9446 (N_9446,N_6853,N_6035);
or U9447 (N_9447,N_8473,N_8793);
and U9448 (N_9448,N_7630,N_6698);
nand U9449 (N_9449,N_8716,N_7266);
nor U9450 (N_9450,N_6074,N_8033);
or U9451 (N_9451,N_6012,N_8154);
or U9452 (N_9452,N_8281,N_6042);
and U9453 (N_9453,N_8688,N_6919);
and U9454 (N_9454,N_7436,N_7316);
nor U9455 (N_9455,N_7473,N_6155);
xnor U9456 (N_9456,N_7582,N_6538);
nor U9457 (N_9457,N_7264,N_8631);
nand U9458 (N_9458,N_7873,N_8003);
nand U9459 (N_9459,N_6172,N_8315);
nand U9460 (N_9460,N_8561,N_7792);
nor U9461 (N_9461,N_8539,N_8497);
xor U9462 (N_9462,N_7516,N_6723);
xor U9463 (N_9463,N_8914,N_8028);
nor U9464 (N_9464,N_6050,N_8293);
xor U9465 (N_9465,N_6286,N_8881);
xor U9466 (N_9466,N_8714,N_8007);
xor U9467 (N_9467,N_7613,N_7933);
xnor U9468 (N_9468,N_6671,N_8084);
nor U9469 (N_9469,N_6332,N_8488);
nand U9470 (N_9470,N_7081,N_8540);
nor U9471 (N_9471,N_6801,N_6602);
nand U9472 (N_9472,N_6324,N_6662);
xnor U9473 (N_9473,N_8186,N_7045);
nor U9474 (N_9474,N_8029,N_6556);
and U9475 (N_9475,N_8409,N_7608);
or U9476 (N_9476,N_8831,N_6067);
nor U9477 (N_9477,N_8067,N_8624);
or U9478 (N_9478,N_8248,N_6313);
or U9479 (N_9479,N_6615,N_8050);
or U9480 (N_9480,N_7126,N_6889);
nand U9481 (N_9481,N_6771,N_8942);
xnor U9482 (N_9482,N_7317,N_7596);
and U9483 (N_9483,N_7271,N_6702);
or U9484 (N_9484,N_8602,N_7428);
or U9485 (N_9485,N_7188,N_6000);
or U9486 (N_9486,N_7367,N_7882);
nor U9487 (N_9487,N_6874,N_7245);
nor U9488 (N_9488,N_7094,N_6846);
or U9489 (N_9489,N_7648,N_8091);
or U9490 (N_9490,N_7926,N_8858);
xor U9491 (N_9491,N_8715,N_7995);
xnor U9492 (N_9492,N_7851,N_8133);
nor U9493 (N_9493,N_6459,N_8307);
nand U9494 (N_9494,N_7771,N_6082);
nor U9495 (N_9495,N_8385,N_8352);
and U9496 (N_9496,N_8299,N_8641);
nand U9497 (N_9497,N_8711,N_7230);
or U9498 (N_9498,N_7534,N_8005);
nand U9499 (N_9499,N_7395,N_6878);
xnor U9500 (N_9500,N_7619,N_8422);
or U9501 (N_9501,N_6604,N_6464);
or U9502 (N_9502,N_8837,N_7974);
nand U9503 (N_9503,N_7024,N_6255);
and U9504 (N_9504,N_6725,N_6363);
nor U9505 (N_9505,N_8117,N_7732);
nor U9506 (N_9506,N_8122,N_8532);
and U9507 (N_9507,N_7212,N_7173);
or U9508 (N_9508,N_7617,N_6818);
or U9509 (N_9509,N_8755,N_7298);
and U9510 (N_9510,N_8412,N_8892);
xnor U9511 (N_9511,N_6392,N_6307);
nand U9512 (N_9512,N_7110,N_8330);
xnor U9513 (N_9513,N_6558,N_8673);
and U9514 (N_9514,N_7247,N_6640);
and U9515 (N_9515,N_8692,N_7419);
nand U9516 (N_9516,N_8405,N_6883);
and U9517 (N_9517,N_8903,N_7164);
nor U9518 (N_9518,N_8553,N_6083);
xnor U9519 (N_9519,N_6990,N_6850);
or U9520 (N_9520,N_8183,N_8644);
nand U9521 (N_9521,N_8605,N_6658);
xor U9522 (N_9522,N_8361,N_8403);
xor U9523 (N_9523,N_6423,N_8581);
nor U9524 (N_9524,N_6917,N_7875);
or U9525 (N_9525,N_8906,N_6923);
and U9526 (N_9526,N_8100,N_8580);
or U9527 (N_9527,N_7348,N_7310);
or U9528 (N_9528,N_6935,N_6273);
and U9529 (N_9529,N_7066,N_6482);
or U9530 (N_9530,N_6399,N_6317);
or U9531 (N_9531,N_8394,N_6581);
nand U9532 (N_9532,N_6356,N_8984);
and U9533 (N_9533,N_6216,N_6101);
nand U9534 (N_9534,N_6377,N_7224);
xor U9535 (N_9535,N_7030,N_8075);
nor U9536 (N_9536,N_8516,N_7560);
nor U9537 (N_9537,N_8276,N_6430);
or U9538 (N_9538,N_6586,N_8682);
or U9539 (N_9539,N_8316,N_7746);
xor U9540 (N_9540,N_8027,N_7342);
nand U9541 (N_9541,N_6767,N_6450);
nand U9542 (N_9542,N_6711,N_7194);
or U9543 (N_9543,N_7088,N_8341);
and U9544 (N_9544,N_7756,N_6321);
nor U9545 (N_9545,N_8264,N_8927);
and U9546 (N_9546,N_8098,N_6579);
nand U9547 (N_9547,N_7632,N_6892);
nor U9548 (N_9548,N_7214,N_7219);
nand U9549 (N_9549,N_6388,N_7113);
xor U9550 (N_9550,N_6407,N_6189);
or U9551 (N_9551,N_7533,N_6837);
xor U9552 (N_9552,N_7865,N_7820);
nand U9553 (N_9553,N_6038,N_6153);
or U9554 (N_9554,N_6575,N_6238);
and U9555 (N_9555,N_8340,N_8515);
and U9556 (N_9556,N_7590,N_7512);
nand U9557 (N_9557,N_8918,N_8446);
nand U9558 (N_9558,N_6956,N_8812);
nor U9559 (N_9559,N_8586,N_6121);
nand U9560 (N_9560,N_6420,N_6933);
or U9561 (N_9561,N_8813,N_8041);
nor U9562 (N_9562,N_7123,N_6115);
or U9563 (N_9563,N_7941,N_7530);
nor U9564 (N_9564,N_8823,N_8036);
nor U9565 (N_9565,N_7665,N_8231);
or U9566 (N_9566,N_7016,N_8731);
and U9567 (N_9567,N_7727,N_6287);
or U9568 (N_9568,N_6194,N_7140);
nor U9569 (N_9569,N_7486,N_6618);
xor U9570 (N_9570,N_8790,N_6031);
or U9571 (N_9571,N_7130,N_6230);
and U9572 (N_9572,N_8390,N_8421);
nor U9573 (N_9573,N_7242,N_6653);
nand U9574 (N_9574,N_7911,N_6619);
xnor U9575 (N_9575,N_8528,N_6806);
nor U9576 (N_9576,N_8042,N_7409);
or U9577 (N_9577,N_6743,N_8289);
nand U9578 (N_9578,N_6323,N_6419);
or U9579 (N_9579,N_7861,N_7984);
nand U9580 (N_9580,N_8669,N_8163);
nor U9581 (N_9581,N_6873,N_8830);
and U9582 (N_9582,N_6580,N_6513);
nand U9583 (N_9583,N_8550,N_8235);
nand U9584 (N_9584,N_7163,N_6843);
xnor U9585 (N_9585,N_6106,N_6617);
or U9586 (N_9586,N_8009,N_6595);
or U9587 (N_9587,N_6123,N_6792);
and U9588 (N_9588,N_7866,N_6914);
nand U9589 (N_9589,N_7729,N_8776);
xor U9590 (N_9590,N_8188,N_7067);
or U9591 (N_9591,N_8290,N_8305);
nor U9592 (N_9592,N_6632,N_8318);
xnor U9593 (N_9593,N_8076,N_6359);
and U9594 (N_9594,N_7131,N_6131);
nand U9595 (N_9595,N_7914,N_8142);
xor U9596 (N_9596,N_8975,N_6341);
or U9597 (N_9597,N_6537,N_7426);
nand U9598 (N_9598,N_6445,N_7386);
or U9599 (N_9599,N_8842,N_8548);
and U9600 (N_9600,N_7532,N_6004);
xor U9601 (N_9601,N_6636,N_8474);
and U9602 (N_9602,N_7940,N_8132);
xor U9603 (N_9603,N_7256,N_7691);
nor U9604 (N_9604,N_6446,N_7870);
xnor U9605 (N_9605,N_6582,N_6719);
nand U9606 (N_9606,N_7246,N_6703);
nand U9607 (N_9607,N_6201,N_7096);
or U9608 (N_9608,N_8054,N_8456);
nor U9609 (N_9609,N_6162,N_8401);
and U9610 (N_9610,N_8883,N_8157);
xnor U9611 (N_9611,N_7368,N_6890);
nand U9612 (N_9612,N_8536,N_6002);
nand U9613 (N_9613,N_6688,N_8707);
xor U9614 (N_9614,N_7385,N_7567);
nor U9615 (N_9615,N_7026,N_7121);
xnor U9616 (N_9616,N_8630,N_7730);
nor U9617 (N_9617,N_8357,N_8251);
nand U9618 (N_9618,N_7370,N_6803);
or U9619 (N_9619,N_8066,N_6474);
xor U9620 (N_9620,N_7769,N_6412);
xor U9621 (N_9621,N_8928,N_7945);
xnor U9622 (N_9622,N_8684,N_7829);
nor U9623 (N_9623,N_7154,N_7216);
xor U9624 (N_9624,N_8650,N_6737);
or U9625 (N_9625,N_6676,N_7988);
or U9626 (N_9626,N_8950,N_6009);
and U9627 (N_9627,N_8404,N_7498);
nand U9628 (N_9628,N_8234,N_7079);
nor U9629 (N_9629,N_7243,N_7003);
and U9630 (N_9630,N_6141,N_8223);
nand U9631 (N_9631,N_7090,N_6550);
and U9632 (N_9632,N_7099,N_8654);
and U9633 (N_9633,N_7674,N_6053);
nor U9634 (N_9634,N_8665,N_6729);
or U9635 (N_9635,N_7708,N_7700);
nor U9636 (N_9636,N_8569,N_8988);
nand U9637 (N_9637,N_6281,N_7699);
and U9638 (N_9638,N_7336,N_7959);
and U9639 (N_9639,N_8710,N_6898);
or U9640 (N_9640,N_7789,N_7055);
nor U9641 (N_9641,N_8346,N_6315);
xor U9642 (N_9642,N_7199,N_7737);
and U9643 (N_9643,N_8070,N_7936);
and U9644 (N_9644,N_8206,N_7318);
nor U9645 (N_9645,N_6927,N_8048);
nand U9646 (N_9646,N_6659,N_7815);
nor U9647 (N_9647,N_8417,N_8746);
xor U9648 (N_9648,N_6008,N_8481);
and U9649 (N_9649,N_7706,N_8947);
and U9650 (N_9650,N_6875,N_7799);
or U9651 (N_9651,N_6306,N_7662);
xnor U9652 (N_9652,N_8190,N_7858);
and U9653 (N_9653,N_7935,N_7411);
or U9654 (N_9654,N_6627,N_6334);
nor U9655 (N_9655,N_7852,N_6953);
nand U9656 (N_9656,N_6742,N_6930);
or U9657 (N_9657,N_8297,N_6854);
xor U9658 (N_9658,N_6967,N_7181);
or U9659 (N_9659,N_6999,N_8944);
or U9660 (N_9660,N_8818,N_8062);
and U9661 (N_9661,N_6851,N_6371);
or U9662 (N_9662,N_7041,N_8094);
nor U9663 (N_9663,N_8331,N_6405);
nand U9664 (N_9664,N_7951,N_7969);
xnor U9665 (N_9665,N_8575,N_7947);
and U9666 (N_9666,N_7584,N_8166);
or U9667 (N_9667,N_7268,N_6734);
and U9668 (N_9668,N_7651,N_6541);
xnor U9669 (N_9669,N_8116,N_8311);
nor U9670 (N_9670,N_7817,N_8323);
and U9671 (N_9671,N_8135,N_7857);
nand U9672 (N_9672,N_8192,N_7279);
and U9673 (N_9673,N_8257,N_7999);
nor U9674 (N_9674,N_6576,N_6950);
xor U9675 (N_9675,N_6292,N_8717);
nand U9676 (N_9676,N_8778,N_6531);
and U9677 (N_9677,N_7343,N_8658);
nand U9678 (N_9678,N_7146,N_7448);
or U9679 (N_9679,N_7340,N_6515);
xnor U9680 (N_9680,N_8538,N_8936);
or U9681 (N_9681,N_7930,N_7459);
nand U9682 (N_9682,N_6894,N_6242);
nor U9683 (N_9683,N_6116,N_8523);
or U9684 (N_9684,N_7396,N_6051);
xnor U9685 (N_9685,N_8640,N_8439);
xor U9686 (N_9686,N_6275,N_6553);
and U9687 (N_9687,N_7548,N_6612);
xnor U9688 (N_9688,N_8452,N_7347);
or U9689 (N_9689,N_7153,N_6754);
nor U9690 (N_9690,N_6078,N_8670);
and U9691 (N_9691,N_7958,N_8356);
xor U9692 (N_9692,N_6554,N_6565);
nor U9693 (N_9693,N_8787,N_8489);
or U9694 (N_9694,N_7825,N_8151);
or U9695 (N_9695,N_7929,N_6178);
and U9696 (N_9696,N_6505,N_7735);
or U9697 (N_9697,N_7005,N_6110);
or U9698 (N_9698,N_8798,N_8243);
or U9699 (N_9699,N_8526,N_8184);
nand U9700 (N_9700,N_6705,N_6380);
and U9701 (N_9701,N_6848,N_8582);
and U9702 (N_9702,N_7075,N_6190);
nor U9703 (N_9703,N_6262,N_8280);
nand U9704 (N_9704,N_6960,N_8973);
or U9705 (N_9705,N_6971,N_7676);
and U9706 (N_9706,N_6660,N_7824);
nand U9707 (N_9707,N_8959,N_7082);
nor U9708 (N_9708,N_6437,N_6109);
and U9709 (N_9709,N_7431,N_7132);
nor U9710 (N_9710,N_8628,N_6680);
or U9711 (N_9711,N_8976,N_7504);
nand U9712 (N_9712,N_7561,N_8621);
and U9713 (N_9713,N_8466,N_6794);
and U9714 (N_9714,N_7366,N_7931);
or U9715 (N_9715,N_6047,N_6069);
nor U9716 (N_9716,N_8485,N_8828);
or U9717 (N_9717,N_7854,N_7843);
and U9718 (N_9718,N_7290,N_8376);
nor U9719 (N_9719,N_6836,N_7018);
xnor U9720 (N_9720,N_6124,N_8901);
and U9721 (N_9721,N_8337,N_6415);
xor U9722 (N_9722,N_6885,N_7604);
xnor U9723 (N_9723,N_6689,N_8073);
nor U9724 (N_9724,N_6163,N_7814);
or U9725 (N_9725,N_6591,N_7360);
nor U9726 (N_9726,N_8113,N_8882);
xnor U9727 (N_9727,N_8551,N_7537);
or U9728 (N_9728,N_7302,N_7538);
nor U9729 (N_9729,N_6916,N_7118);
or U9730 (N_9730,N_6509,N_6793);
xor U9731 (N_9731,N_7280,N_8629);
nand U9732 (N_9732,N_7956,N_7864);
xor U9733 (N_9733,N_6144,N_8214);
nor U9734 (N_9734,N_6664,N_8314);
and U9735 (N_9735,N_6808,N_8049);
nor U9736 (N_9736,N_6644,N_7254);
and U9737 (N_9737,N_8322,N_7285);
nor U9738 (N_9738,N_8229,N_8326);
nor U9739 (N_9739,N_8219,N_7804);
or U9740 (N_9740,N_6122,N_8808);
or U9741 (N_9741,N_6329,N_8549);
xnor U9742 (N_9742,N_6954,N_7484);
nand U9743 (N_9743,N_8213,N_7819);
and U9744 (N_9744,N_7884,N_6495);
xnor U9745 (N_9745,N_6468,N_6508);
nor U9746 (N_9746,N_6340,N_7519);
and U9747 (N_9747,N_8127,N_8957);
or U9748 (N_9748,N_7709,N_6963);
nand U9749 (N_9749,N_6188,N_7610);
or U9750 (N_9750,N_7791,N_7058);
or U9751 (N_9751,N_6331,N_7528);
or U9752 (N_9752,N_7288,N_8705);
or U9753 (N_9753,N_8095,N_6448);
or U9754 (N_9754,N_8990,N_7092);
nand U9755 (N_9755,N_7831,N_6731);
nand U9756 (N_9756,N_7650,N_7175);
or U9757 (N_9757,N_7475,N_8021);
nand U9758 (N_9758,N_6090,N_6424);
or U9759 (N_9759,N_7495,N_7037);
or U9760 (N_9760,N_6781,N_7764);
nor U9761 (N_9761,N_6300,N_7407);
xnor U9762 (N_9762,N_8985,N_7524);
or U9763 (N_9763,N_7027,N_8690);
and U9764 (N_9764,N_7180,N_7661);
xor U9765 (N_9765,N_6197,N_6902);
nand U9766 (N_9766,N_6104,N_7868);
nor U9767 (N_9767,N_8564,N_8131);
and U9768 (N_9768,N_7477,N_6496);
or U9769 (N_9769,N_8949,N_6477);
xnor U9770 (N_9770,N_6108,N_8834);
or U9771 (N_9771,N_6699,N_7299);
and U9772 (N_9772,N_7493,N_6427);
or U9773 (N_9773,N_7905,N_6250);
or U9774 (N_9774,N_8933,N_7087);
nand U9775 (N_9775,N_8563,N_7108);
xor U9776 (N_9776,N_7633,N_7714);
and U9777 (N_9777,N_8193,N_6861);
xor U9778 (N_9778,N_6822,N_6212);
xnor U9779 (N_9779,N_7808,N_6946);
nand U9780 (N_9780,N_6539,N_8635);
xor U9781 (N_9781,N_7531,N_7365);
or U9782 (N_9782,N_6465,N_7136);
nor U9783 (N_9783,N_6588,N_6825);
and U9784 (N_9784,N_8981,N_7626);
and U9785 (N_9785,N_7372,N_6179);
xnor U9786 (N_9786,N_6998,N_8175);
or U9787 (N_9787,N_7304,N_8873);
nor U9788 (N_9788,N_8442,N_7913);
nand U9789 (N_9789,N_8533,N_6975);
xor U9790 (N_9790,N_7558,N_6246);
nor U9791 (N_9791,N_7527,N_7472);
or U9792 (N_9792,N_7186,N_6322);
nor U9793 (N_9793,N_8958,N_6214);
or U9794 (N_9794,N_7511,N_8224);
nor U9795 (N_9795,N_6639,N_7707);
xnor U9796 (N_9796,N_7374,N_6812);
nor U9797 (N_9797,N_7414,N_8736);
xnor U9798 (N_9798,N_8632,N_8411);
nand U9799 (N_9799,N_8871,N_6422);
nor U9800 (N_9800,N_6715,N_6368);
and U9801 (N_9801,N_6019,N_8643);
xnor U9802 (N_9802,N_6713,N_7073);
xor U9803 (N_9803,N_7638,N_8428);
nand U9804 (N_9804,N_8777,N_7776);
and U9805 (N_9805,N_6540,N_6855);
and U9806 (N_9806,N_7207,N_7510);
nor U9807 (N_9807,N_6969,N_8469);
nand U9808 (N_9808,N_7485,N_8230);
xor U9809 (N_9809,N_7390,N_8101);
nand U9810 (N_9810,N_8725,N_8708);
and U9811 (N_9811,N_8642,N_8107);
nor U9812 (N_9812,N_7458,N_7987);
xor U9813 (N_9813,N_6726,N_8565);
nand U9814 (N_9814,N_7038,N_8045);
and U9815 (N_9815,N_7000,N_6386);
or U9816 (N_9816,N_7599,N_7470);
nand U9817 (N_9817,N_8598,N_8689);
or U9818 (N_9818,N_7938,N_7265);
nand U9819 (N_9819,N_8430,N_6352);
nand U9820 (N_9820,N_7168,N_6048);
nand U9821 (N_9821,N_8008,N_7119);
xor U9822 (N_9822,N_6498,N_6813);
nor U9823 (N_9823,N_8338,N_8592);
nand U9824 (N_9824,N_8970,N_8068);
or U9825 (N_9825,N_7117,N_8200);
nand U9826 (N_9826,N_6650,N_8920);
and U9827 (N_9827,N_6160,N_8304);
xor U9828 (N_9828,N_7200,N_6151);
xor U9829 (N_9829,N_7301,N_6080);
or U9830 (N_9830,N_8637,N_8571);
xor U9831 (N_9831,N_6574,N_6139);
or U9832 (N_9832,N_6521,N_7892);
xor U9833 (N_9833,N_8744,N_6524);
and U9834 (N_9834,N_6906,N_6228);
or U9835 (N_9835,N_6807,N_6103);
xnor U9836 (N_9836,N_7897,N_8591);
nor U9837 (N_9837,N_7677,N_6708);
and U9838 (N_9838,N_8974,N_7583);
and U9839 (N_9839,N_6900,N_6265);
and U9840 (N_9840,N_6234,N_8486);
and U9841 (N_9841,N_7471,N_8747);
xor U9842 (N_9842,N_6881,N_7359);
xor U9843 (N_9843,N_7425,N_8754);
and U9844 (N_9844,N_6714,N_6606);
nor U9845 (N_9845,N_6589,N_7575);
or U9846 (N_9846,N_7877,N_7326);
nor U9847 (N_9847,N_8588,N_6603);
or U9848 (N_9848,N_6357,N_8913);
nand U9849 (N_9849,N_6549,N_7137);
nor U9850 (N_9850,N_7293,N_8025);
xnor U9851 (N_9851,N_8468,N_7692);
or U9852 (N_9852,N_8099,N_7203);
or U9853 (N_9853,N_8625,N_8556);
or U9854 (N_9854,N_7435,N_6959);
xnor U9855 (N_9855,N_8584,N_6221);
nand U9856 (N_9856,N_8722,N_7639);
and U9857 (N_9857,N_8242,N_8583);
and U9858 (N_9858,N_6451,N_7724);
nor U9859 (N_9859,N_7962,N_7033);
or U9860 (N_9860,N_7620,N_8980);
xnor U9861 (N_9861,N_8820,N_8267);
xnor U9862 (N_9862,N_8860,N_6921);
and U9863 (N_9863,N_7806,N_7106);
and U9864 (N_9864,N_6982,N_7341);
or U9865 (N_9865,N_7467,N_6961);
and U9866 (N_9866,N_8121,N_7078);
xor U9867 (N_9867,N_7991,N_6128);
and U9868 (N_9868,N_7182,N_7961);
and U9869 (N_9869,N_8074,N_7128);
nand U9870 (N_9870,N_7465,N_6046);
xor U9871 (N_9871,N_8302,N_8351);
xor U9872 (N_9872,N_7107,N_7775);
nand U9873 (N_9873,N_8743,N_6931);
xnor U9874 (N_9874,N_7464,N_8573);
xnor U9875 (N_9875,N_7239,N_6593);
nand U9876 (N_9876,N_6908,N_8240);
and U9877 (N_9877,N_8360,N_7547);
or U9878 (N_9878,N_6778,N_8118);
nand U9879 (N_9879,N_6858,N_7612);
nand U9880 (N_9880,N_6071,N_7754);
and U9881 (N_9881,N_7192,N_6677);
xor U9882 (N_9882,N_6633,N_8419);
xor U9883 (N_9883,N_7314,N_7501);
xnor U9884 (N_9884,N_8617,N_6690);
xnor U9885 (N_9885,N_6091,N_7357);
nand U9886 (N_9886,N_7697,N_6519);
nor U9887 (N_9887,N_7148,N_6125);
or U9888 (N_9888,N_6972,N_6597);
nand U9889 (N_9889,N_8071,N_6186);
xor U9890 (N_9890,N_6398,N_8639);
nor U9891 (N_9891,N_6268,N_7469);
nand U9892 (N_9892,N_6966,N_6089);
xnor U9893 (N_9893,N_7143,N_6608);
and U9894 (N_9894,N_6005,N_8864);
nor U9895 (N_9895,N_8622,N_7069);
nand U9896 (N_9896,N_7862,N_8612);
xnor U9897 (N_9897,N_6303,N_6241);
nor U9898 (N_9898,N_7021,N_7636);
and U9899 (N_9899,N_8072,N_6765);
xnor U9900 (N_9900,N_8298,N_6940);
nor U9901 (N_9901,N_8397,N_7517);
xnor U9902 (N_9902,N_8415,N_6730);
or U9903 (N_9903,N_7044,N_7627);
nand U9904 (N_9904,N_6752,N_6833);
or U9905 (N_9905,N_6547,N_6502);
and U9906 (N_9906,N_7297,N_6736);
nand U9907 (N_9907,N_6258,N_7562);
or U9908 (N_9908,N_7953,N_8364);
xor U9909 (N_9909,N_8838,N_6102);
nor U9910 (N_9910,N_8868,N_8178);
xor U9911 (N_9911,N_8867,N_7397);
nor U9912 (N_9912,N_7032,N_8410);
xor U9913 (N_9913,N_8739,N_8484);
xor U9914 (N_9914,N_7813,N_7609);
or U9915 (N_9915,N_7408,N_8278);
or U9916 (N_9916,N_6010,N_6863);
and U9917 (N_9917,N_8059,N_8187);
nor U9918 (N_9918,N_7993,N_7097);
nor U9919 (N_9919,N_7570,N_6503);
xor U9920 (N_9920,N_6247,N_8249);
nor U9921 (N_9921,N_6057,N_6596);
nor U9922 (N_9922,N_7480,N_8020);
nand U9923 (N_9923,N_7111,N_7536);
nand U9924 (N_9924,N_7196,N_6656);
nand U9925 (N_9925,N_7946,N_6014);
nor U9926 (N_9926,N_7821,N_7859);
and U9927 (N_9927,N_8706,N_8172);
and U9928 (N_9928,N_8044,N_7014);
nand U9929 (N_9929,N_8355,N_6304);
and U9930 (N_9930,N_8226,N_7925);
or U9931 (N_9931,N_6945,N_8170);
and U9932 (N_9932,N_7220,N_7917);
xnor U9933 (N_9933,N_8676,N_8844);
nand U9934 (N_9934,N_8016,N_6133);
nor U9935 (N_9935,N_6831,N_6476);
nor U9936 (N_9936,N_6607,N_8554);
or U9937 (N_9937,N_6018,N_7839);
or U9938 (N_9938,N_7460,N_6616);
and U9939 (N_9939,N_8543,N_7324);
nor U9940 (N_9940,N_8274,N_7686);
or U9941 (N_9941,N_6986,N_7010);
or U9942 (N_9942,N_8277,N_8685);
nand U9943 (N_9943,N_6516,N_8143);
or U9944 (N_9944,N_7919,N_7382);
nor U9945 (N_9945,N_7520,N_7968);
xor U9946 (N_9946,N_8847,N_8431);
and U9947 (N_9947,N_8853,N_7434);
nand U9948 (N_9948,N_8610,N_6951);
and U9949 (N_9949,N_8733,N_6170);
xnor U9950 (N_9950,N_6585,N_7680);
nand U9951 (N_9951,N_6510,N_7798);
nand U9952 (N_9952,N_7053,N_8342);
nor U9953 (N_9953,N_7233,N_8537);
xor U9954 (N_9954,N_8861,N_7344);
or U9955 (N_9955,N_7543,N_7895);
and U9956 (N_9956,N_7767,N_7127);
nand U9957 (N_9957,N_7848,N_8559);
and U9958 (N_9958,N_8943,N_7770);
xnor U9959 (N_9959,N_8770,N_7273);
nor U9960 (N_9960,N_6630,N_7952);
nor U9961 (N_9961,N_7779,N_8649);
nor U9962 (N_9962,N_6988,N_8785);
and U9963 (N_9963,N_7910,N_8668);
nor U9964 (N_9964,N_8258,N_6783);
and U9965 (N_9965,N_6181,N_7025);
xnor U9966 (N_9966,N_7675,N_6467);
or U9967 (N_9967,N_6040,N_6013);
xor U9968 (N_9968,N_7404,N_7618);
or U9969 (N_9969,N_8961,N_8507);
nor U9970 (N_9970,N_8730,N_8292);
nand U9971 (N_9971,N_8921,N_7508);
nor U9972 (N_9972,N_8530,N_6746);
or U9973 (N_9973,N_7179,N_6564);
or U9974 (N_9974,N_8699,N_8420);
nor U9975 (N_9975,N_7983,N_6254);
and U9976 (N_9976,N_6493,N_8125);
nand U9977 (N_9977,N_7879,N_8991);
nor U9978 (N_9978,N_8948,N_6418);
or U9979 (N_9979,N_6063,N_6609);
nor U9980 (N_9980,N_8721,N_7210);
and U9981 (N_9981,N_6980,N_7104);
and U9982 (N_9982,N_7654,N_6862);
nor U9983 (N_9983,N_8031,N_8729);
and U9984 (N_9984,N_6087,N_7308);
xnor U9985 (N_9985,N_6213,N_6529);
and U9986 (N_9986,N_6195,N_6973);
or U9987 (N_9987,N_6847,N_6389);
nand U9988 (N_9988,N_8146,N_7977);
nand U9989 (N_9989,N_7642,N_6320);
nor U9990 (N_9990,N_6879,N_6670);
nor U9991 (N_9991,N_6166,N_7262);
or U9992 (N_9992,N_6150,N_6379);
and U9993 (N_9993,N_6773,N_7427);
nor U9994 (N_9994,N_8805,N_8570);
nand U9995 (N_9995,N_7625,N_8291);
xor U9996 (N_9996,N_7101,N_7924);
nor U9997 (N_9997,N_8370,N_7035);
or U9998 (N_9998,N_6049,N_6114);
or U9999 (N_9999,N_8911,N_6830);
or U10000 (N_10000,N_8899,N_6584);
xnor U10001 (N_10001,N_6454,N_7753);
or U10002 (N_10002,N_6867,N_8150);
nor U10003 (N_10003,N_8174,N_6904);
nor U10004 (N_10004,N_8935,N_7967);
xor U10005 (N_10005,N_8383,N_6838);
and U10006 (N_10006,N_6748,N_6701);
nor U10007 (N_10007,N_8542,N_6274);
and U10008 (N_10008,N_7920,N_7515);
nor U10009 (N_10009,N_8951,N_8019);
nor U10010 (N_10010,N_6785,N_8874);
xor U10011 (N_10011,N_7581,N_8424);
xor U10012 (N_10012,N_7768,N_6533);
or U10013 (N_10013,N_7363,N_6673);
and U10014 (N_10014,N_7312,N_6426);
xnor U10015 (N_10015,N_7809,N_7138);
or U10016 (N_10016,N_6337,N_8271);
xor U10017 (N_10017,N_6751,N_7856);
or U10018 (N_10018,N_8952,N_7466);
nor U10019 (N_10019,N_7376,N_7563);
and U10020 (N_10020,N_8261,N_8782);
or U10021 (N_10021,N_8919,N_7846);
nor U10022 (N_10022,N_6629,N_7641);
xnor U10023 (N_10023,N_8814,N_8106);
xnor U10024 (N_10024,N_6763,N_6819);
and U10025 (N_10025,N_6860,N_6587);
nand U10026 (N_10026,N_6716,N_8309);
xor U10027 (N_10027,N_6922,N_8504);
or U10028 (N_10028,N_7378,N_7429);
xnor U10029 (N_10029,N_7457,N_8999);
or U10030 (N_10030,N_7606,N_7577);
nand U10031 (N_10031,N_7303,N_8594);
nand U10032 (N_10032,N_6438,N_8162);
or U10033 (N_10033,N_6829,N_7476);
nor U10034 (N_10034,N_7449,N_6780);
xor U10035 (N_10035,N_8956,N_8893);
nand U10036 (N_10036,N_6871,N_8256);
xor U10037 (N_10037,N_8447,N_7904);
or U10038 (N_10038,N_8359,N_6691);
nor U10039 (N_10039,N_6309,N_8719);
nor U10040 (N_10040,N_6117,N_7578);
xnor U10041 (N_10041,N_7741,N_8546);
nor U10042 (N_10042,N_8483,N_6156);
and U10043 (N_10043,N_8521,N_6666);
xor U10044 (N_10044,N_7743,N_7915);
nand U10045 (N_10045,N_6383,N_6824);
xnor U10046 (N_10046,N_8039,N_7071);
and U10047 (N_10047,N_8472,N_6681);
nand U10048 (N_10048,N_7832,N_7232);
nor U10049 (N_10049,N_6983,N_8090);
nand U10050 (N_10050,N_6869,N_6199);
xor U10051 (N_10051,N_6942,N_6344);
or U10052 (N_10052,N_6056,N_6924);
and U10053 (N_10053,N_7338,N_6984);
nand U10054 (N_10054,N_6788,N_7184);
or U10055 (N_10055,N_8815,N_8275);
nand U10056 (N_10056,N_8797,N_8880);
nand U10057 (N_10057,N_8759,N_8816);
nand U10058 (N_10058,N_8303,N_6202);
nand U10059 (N_10059,N_8909,N_6598);
and U10060 (N_10060,N_6140,N_7885);
nand U10061 (N_10061,N_6903,N_6484);
nand U10062 (N_10062,N_6741,N_7711);
nand U10063 (N_10063,N_8225,N_6021);
xnor U10064 (N_10064,N_7332,N_8181);
nand U10065 (N_10065,N_6152,N_6759);
and U10066 (N_10066,N_8608,N_7572);
or U10067 (N_10067,N_7715,N_7942);
nand U10068 (N_10068,N_6276,N_7047);
nand U10069 (N_10069,N_6842,N_7622);
and U10070 (N_10070,N_8245,N_6456);
nor U10071 (N_10071,N_8083,N_7197);
xor U10072 (N_10072,N_6135,N_8511);
nand U10073 (N_10073,N_6646,N_7358);
nor U10074 (N_10074,N_7975,N_8197);
nand U10075 (N_10075,N_6868,N_7751);
xor U10076 (N_10076,N_7542,N_8996);
and U10077 (N_10077,N_8294,N_7871);
nor U10078 (N_10078,N_6506,N_6350);
or U10079 (N_10079,N_8111,N_7080);
or U10080 (N_10080,N_6913,N_8189);
nand U10081 (N_10081,N_6011,N_8265);
nand U10082 (N_10082,N_8541,N_8124);
xor U10083 (N_10083,N_7483,N_8325);
or U10084 (N_10084,N_7628,N_7773);
nor U10085 (N_10085,N_7668,N_7160);
and U10086 (N_10086,N_8161,N_8471);
nor U10087 (N_10087,N_7818,N_8531);
xnor U10088 (N_10088,N_6266,N_6864);
xor U10089 (N_10089,N_7292,N_7973);
nor U10090 (N_10090,N_8579,N_7705);
nor U10091 (N_10091,N_6395,N_8620);
or U10092 (N_10092,N_6314,N_8886);
or U10093 (N_10093,N_7916,N_7591);
nand U10094 (N_10094,N_6196,N_7478);
and U10095 (N_10095,N_6294,N_7985);
xor U10096 (N_10096,N_7994,N_6817);
and U10097 (N_10097,N_7091,N_6126);
xnor U10098 (N_10098,N_7506,N_7589);
nor U10099 (N_10099,N_6045,N_7156);
nor U10100 (N_10100,N_7725,N_7772);
or U10101 (N_10101,N_6284,N_8102);
and U10102 (N_10102,N_6374,N_7198);
nor U10103 (N_10103,N_8012,N_8408);
nor U10104 (N_10104,N_8712,N_7514);
nor U10105 (N_10105,N_8600,N_6620);
xor U10106 (N_10106,N_8522,N_8751);
nor U10107 (N_10107,N_8392,N_8244);
and U10108 (N_10108,N_6060,N_8978);
nand U10109 (N_10109,N_6381,N_8057);
nand U10110 (N_10110,N_8872,N_7481);
nand U10111 (N_10111,N_8518,N_7049);
and U10112 (N_10112,N_8215,N_7012);
and U10113 (N_10113,N_6937,N_6685);
xnor U10114 (N_10114,N_8077,N_8803);
or U10115 (N_10115,N_8524,N_6485);
nand U10116 (N_10116,N_8078,N_8270);
xnor U10117 (N_10117,N_8574,N_6443);
nand U10118 (N_10118,N_7586,N_7403);
and U10119 (N_10119,N_8241,N_8141);
or U10120 (N_10120,N_7191,N_6064);
nor U10121 (N_10121,N_8459,N_6887);
xor U10122 (N_10122,N_6706,N_8505);
nand U10123 (N_10123,N_7943,N_8138);
or U10124 (N_10124,N_7311,N_7401);
nor U10125 (N_10125,N_8393,N_6536);
xor U10126 (N_10126,N_6244,N_7331);
nand U10127 (N_10127,N_8382,N_7634);
nor U10128 (N_10128,N_7322,N_7647);
nor U10129 (N_10129,N_8493,N_6148);
and U10130 (N_10130,N_8750,N_8038);
or U10131 (N_10131,N_7978,N_8375);
or U10132 (N_10132,N_8576,N_8771);
nor U10133 (N_10133,N_6962,N_8969);
or U10134 (N_10134,N_6027,N_7783);
nand U10135 (N_10135,N_8502,N_8687);
or U10136 (N_10136,N_8445,N_8995);
nand U10137 (N_10137,N_6481,N_8168);
nand U10138 (N_10138,N_7888,N_8126);
xnor U10139 (N_10139,N_8568,N_7557);
nor U10140 (N_10140,N_6985,N_6175);
xnor U10141 (N_10141,N_6479,N_6798);
nand U10142 (N_10142,N_7834,N_6193);
nor U10143 (N_10143,N_6404,N_7939);
xnor U10144 (N_10144,N_7284,N_7061);
and U10145 (N_10145,N_8718,N_8824);
or U10146 (N_10146,N_7726,N_6384);
and U10147 (N_10147,N_8677,N_7702);
and U10148 (N_10148,N_6500,N_6366);
nor U10149 (N_10149,N_8478,N_8884);
or U10150 (N_10150,N_7159,N_6546);
nand U10151 (N_10151,N_8963,N_8779);
nand U10152 (N_10152,N_6236,N_6859);
xor U10153 (N_10153,N_7039,N_8201);
and U10154 (N_10154,N_8795,N_6316);
xor U10155 (N_10155,N_6571,N_7494);
nand U10156 (N_10156,N_6877,N_6393);
or U10157 (N_10157,N_8179,N_7017);
xor U10158 (N_10158,N_8774,N_6278);
nor U10159 (N_10159,N_7013,N_7614);
nand U10160 (N_10160,N_8221,N_6154);
nor U10161 (N_10161,N_8679,N_8386);
nor U10162 (N_10162,N_8833,N_8388);
or U10163 (N_10163,N_8506,N_7050);
nand U10164 (N_10164,N_8367,N_8476);
nor U10165 (N_10165,N_7139,N_7937);
xnor U10166 (N_10166,N_7417,N_8312);
xor U10167 (N_10167,N_7593,N_6899);
nand U10168 (N_10168,N_6225,N_6349);
nor U10169 (N_10169,N_8144,N_8212);
and U10170 (N_10170,N_7551,N_6977);
and U10171 (N_10171,N_8965,N_6449);
nand U10172 (N_10172,N_7833,N_6626);
or U10173 (N_10173,N_8878,N_6570);
nor U10174 (N_10174,N_7443,N_8399);
and U10175 (N_10175,N_7554,N_8930);
nand U10176 (N_10176,N_6981,N_7658);
or U10177 (N_10177,N_7068,N_7736);
nand U10178 (N_10178,N_8347,N_7782);
nor U10179 (N_10179,N_8173,N_8879);
nor U10180 (N_10180,N_6169,N_8609);
nand U10181 (N_10181,N_6811,N_6062);
nand U10182 (N_10182,N_6143,N_8115);
nor U10183 (N_10183,N_8674,N_8233);
nor U10184 (N_10184,N_8414,N_8204);
nand U10185 (N_10185,N_6480,N_6168);
and U10186 (N_10186,N_7172,N_7125);
or U10187 (N_10187,N_6325,N_8501);
nor U10188 (N_10188,N_7812,N_8802);
and U10189 (N_10189,N_7587,N_8402);
or U10190 (N_10190,N_7682,N_8510);
xnor U10191 (N_10191,N_7574,N_8085);
or U10192 (N_10192,N_8164,N_7518);
and U10193 (N_10193,N_7629,N_8199);
and U10194 (N_10194,N_8783,N_7902);
and U10195 (N_10195,N_8851,N_8171);
and U10196 (N_10196,N_8671,N_7085);
or U10197 (N_10197,N_8811,N_6260);
and U10198 (N_10198,N_7177,N_8001);
xnor U10199 (N_10199,N_7490,N_8379);
nor U10200 (N_10200,N_6497,N_6566);
nor U10201 (N_10201,N_8129,N_6772);
or U10202 (N_10202,N_8611,N_6948);
nor U10203 (N_10203,N_6614,N_7794);
nand U10204 (N_10204,N_7361,N_7492);
xor U10205 (N_10205,N_8700,N_8946);
nand U10206 (N_10206,N_6704,N_6376);
nor U10207 (N_10207,N_6410,N_8185);
nand U10208 (N_10208,N_7810,N_6081);
nor U10209 (N_10209,N_7793,N_6302);
nand U10210 (N_10210,N_6991,N_6113);
xor U10211 (N_10211,N_8155,N_8661);
nand U10212 (N_10212,N_6789,N_8358);
or U10213 (N_10213,N_8152,N_8332);
and U10214 (N_10214,N_8693,N_6805);
or U10215 (N_10215,N_8362,N_8832);
nand U10216 (N_10216,N_7541,N_6882);
nand U10217 (N_10217,N_7503,N_6401);
nor U10218 (N_10218,N_6766,N_7785);
xor U10219 (N_10219,N_8876,N_8158);
or U10220 (N_10220,N_6758,N_8607);
nor U10221 (N_10221,N_7195,N_8662);
or U10222 (N_10222,N_7337,N_8433);
or U10223 (N_10223,N_7189,N_8907);
xor U10224 (N_10224,N_7059,N_6171);
or U10225 (N_10225,N_7105,N_7007);
xnor U10226 (N_10226,N_7757,N_8263);
and U10227 (N_10227,N_8527,N_6624);
and U10228 (N_10228,N_8926,N_7267);
nand U10229 (N_10229,N_6776,N_6514);
and U10230 (N_10230,N_8681,N_8578);
or U10231 (N_10231,N_8723,N_7157);
nor U10232 (N_10232,N_6441,N_7666);
nand U10233 (N_10233,N_8336,N_8737);
nor U10234 (N_10234,N_8651,N_8120);
or U10235 (N_10235,N_7580,N_6834);
and U10236 (N_10236,N_8495,N_8900);
nand U10237 (N_10237,N_7309,N_6952);
xnor U10238 (N_10238,N_7944,N_7134);
or U10239 (N_10239,N_7062,N_6568);
nand U10240 (N_10240,N_7598,N_6738);
or U10241 (N_10241,N_7251,N_6893);
or U10242 (N_10242,N_6253,N_8196);
xor U10243 (N_10243,N_8112,N_7671);
xnor U10244 (N_10244,N_6790,N_8320);
nor U10245 (N_10245,N_7294,N_6203);
nand U10246 (N_10246,N_6932,N_8791);
or U10247 (N_10247,N_7286,N_6635);
and U10248 (N_10248,N_7745,N_7323);
and U10249 (N_10249,N_7205,N_7095);
or U10250 (N_10250,N_8850,N_6525);
or U10251 (N_10251,N_7595,N_7719);
nand U10252 (N_10252,N_8400,N_6076);
or U10253 (N_10253,N_8354,N_7979);
nand U10254 (N_10254,N_7209,N_7867);
xor U10255 (N_10255,N_7399,N_7274);
or U10256 (N_10256,N_7803,N_7723);
and U10257 (N_10257,N_7742,N_7976);
nand U10258 (N_10258,N_7960,N_8821);
and U10259 (N_10259,N_7064,N_8855);
and U10260 (N_10260,N_6264,N_6682);
nand U10261 (N_10261,N_7811,N_7438);
or U10262 (N_10262,N_7765,N_6696);
nor U10263 (N_10263,N_7965,N_7369);
or U10264 (N_10264,N_7659,N_8149);
nor U10265 (N_10265,N_6775,N_6512);
nor U10266 (N_10266,N_7499,N_7655);
nor U10267 (N_10267,N_6222,N_7922);
or U10268 (N_10268,N_6086,N_7394);
xor U10269 (N_10269,N_7579,N_7544);
or U10270 (N_10270,N_7289,N_7056);
xnor U10271 (N_10271,N_6740,N_7218);
nand U10272 (N_10272,N_8329,N_6974);
nand U10273 (N_10273,N_6390,N_8055);
xor U10274 (N_10274,N_7566,N_6373);
nor U10275 (N_10275,N_6394,N_8058);
nand U10276 (N_10276,N_7997,N_7446);
nor U10277 (N_10277,N_8130,N_7607);
or U10278 (N_10278,N_8377,N_6944);
nor U10279 (N_10279,N_7669,N_7689);
xnor U10280 (N_10280,N_8764,N_7122);
nor U10281 (N_10281,N_6668,N_7282);
xor U10282 (N_10282,N_8103,N_7150);
and U10283 (N_10283,N_8732,N_7637);
nor U10284 (N_10284,N_8520,N_6970);
xnor U10285 (N_10285,N_7998,N_8614);
or U10286 (N_10286,N_8461,N_8819);
and U10287 (N_10287,N_6271,N_7569);
xnor U10288 (N_10288,N_7208,N_7597);
nand U10289 (N_10289,N_7545,N_7084);
nor U10290 (N_10290,N_8285,N_6157);
xor U10291 (N_10291,N_8939,N_7496);
or U10292 (N_10292,N_7549,N_7275);
nor U10293 (N_10293,N_7260,N_8983);
nor U10294 (N_10294,N_6760,N_6762);
nor U10295 (N_10295,N_6888,N_7424);
nand U10296 (N_10296,N_6852,N_8772);
and U10297 (N_10297,N_8566,N_7023);
and U10298 (N_10298,N_6433,N_6413);
nand U10299 (N_10299,N_6753,N_6097);
or U10300 (N_10300,N_6569,N_8137);
or U10301 (N_10301,N_7787,N_7307);
or U10302 (N_10302,N_6289,N_6651);
and U10303 (N_10303,N_6623,N_7747);
nor U10304 (N_10304,N_7487,N_8599);
or U10305 (N_10305,N_6402,N_8373);
and U10306 (N_10306,N_6414,N_7171);
or U10307 (N_10307,N_7474,N_6173);
xor U10308 (N_10308,N_7249,N_6936);
xor U10309 (N_10309,N_6856,N_8839);
nand U10310 (N_10310,N_6358,N_7152);
xnor U10311 (N_10311,N_8638,N_6661);
nor U10312 (N_10312,N_7701,N_8480);
xnor U10313 (N_10313,N_6177,N_7281);
and U10314 (N_10314,N_8966,N_7278);
xor U10315 (N_10315,N_8728,N_7759);
and U10316 (N_10316,N_8987,N_7838);
or U10317 (N_10317,N_6520,N_6605);
or U10318 (N_10318,N_7840,N_7900);
or U10319 (N_10319,N_6259,N_6929);
nor U10320 (N_10320,N_6655,N_6335);
and U10321 (N_10321,N_7860,N_8727);
xor U10322 (N_10322,N_8222,N_7505);
xor U10323 (N_10323,N_6557,N_8086);
or U10324 (N_10324,N_8148,N_7762);
nor U10325 (N_10325,N_6444,N_8826);
nand U10326 (N_10326,N_7739,N_7540);
and U10327 (N_10327,N_7206,N_8841);
xnor U10328 (N_10328,N_8380,N_6257);
and U10329 (N_10329,N_8153,N_6997);
xnor U10330 (N_10330,N_6355,N_7422);
nor U10331 (N_10331,N_8809,N_7670);
nand U10332 (N_10332,N_7957,N_8615);
xor U10333 (N_10333,N_6095,N_8762);
xnor U10334 (N_10334,N_6517,N_8545);
or U10335 (N_10335,N_8093,N_8022);
nand U10336 (N_10336,N_7592,N_8912);
or U10337 (N_10337,N_7089,N_8870);
nand U10338 (N_10338,N_7616,N_8387);
xor U10339 (N_10339,N_6494,N_7784);
and U10340 (N_10340,N_7252,N_8953);
nor U10341 (N_10341,N_6149,N_6987);
xnor U10342 (N_10342,N_8349,N_7226);
or U10343 (N_10343,N_6828,N_7250);
or U10344 (N_10344,N_7948,N_6367);
or U10345 (N_10345,N_7352,N_6840);
and U10346 (N_10346,N_6041,N_7786);
xor U10347 (N_10347,N_7502,N_8013);
nand U10348 (N_10348,N_7456,N_7565);
or U10349 (N_10349,N_7158,N_8788);
or U10350 (N_10350,N_6164,N_8268);
nand U10351 (N_10351,N_7717,N_7901);
or U10352 (N_10352,N_8964,N_6191);
nor U10353 (N_10353,N_8176,N_7555);
xnor U10354 (N_10354,N_8940,N_8888);
nand U10355 (N_10355,N_6782,N_6068);
nor U10356 (N_10356,N_6245,N_7695);
nor U10357 (N_10357,N_7259,N_8026);
and U10358 (N_10358,N_8626,N_6610);
xor U10359 (N_10359,N_7356,N_8259);
nand U10360 (N_10360,N_7248,N_8194);
and U10361 (N_10361,N_6417,N_6918);
and U10362 (N_10362,N_6310,N_8104);
nand U10363 (N_10363,N_8381,N_8655);
xor U10364 (N_10364,N_7185,N_7420);
nand U10365 (N_10365,N_6291,N_6839);
and U10366 (N_10366,N_6631,N_6555);
and U10367 (N_10367,N_8789,N_8738);
nand U10368 (N_10368,N_8572,N_8780);
or U10369 (N_10369,N_8767,N_8237);
nand U10370 (N_10370,N_6360,N_8147);
nand U10371 (N_10371,N_6251,N_7744);
xor U10372 (N_10372,N_6428,N_6061);
and U10373 (N_10373,N_8934,N_7065);
or U10374 (N_10374,N_6958,N_8786);
nor U10375 (N_10375,N_7202,N_7992);
nand U10376 (N_10376,N_6724,N_8432);
nor U10377 (N_10377,N_7970,N_7758);
nor U10378 (N_10378,N_7253,N_6369);
nor U10379 (N_10379,N_7377,N_7257);
nor U10380 (N_10380,N_8979,N_6382);
nand U10381 (N_10381,N_8613,N_6036);
or U10382 (N_10382,N_6996,N_7217);
or U10383 (N_10383,N_7660,N_6638);
and U10384 (N_10384,N_6416,N_7170);
nor U10385 (N_10385,N_8060,N_7909);
xnor U10386 (N_10386,N_7450,N_8896);
or U10387 (N_10387,N_8463,N_8056);
nand U10388 (N_10388,N_8955,N_6530);
xnor U10389 (N_10389,N_8849,N_6528);
nand U10390 (N_10390,N_6518,N_7008);
or U10391 (N_10391,N_6006,N_6055);
nand U10392 (N_10392,N_7321,N_8384);
nand U10393 (N_10393,N_7890,N_8061);
nand U10394 (N_10394,N_7835,N_7982);
or U10395 (N_10395,N_6346,N_6621);
nand U10396 (N_10396,N_8765,N_6455);
and U10397 (N_10397,N_7529,N_6628);
and U10398 (N_10398,N_6065,N_8557);
nand U10399 (N_10399,N_7790,N_6820);
and U10400 (N_10400,N_6471,N_7863);
xnor U10401 (N_10401,N_6226,N_6710);
or U10402 (N_10402,N_8406,N_6452);
nor U10403 (N_10403,N_7142,N_8667);
xnor U10404 (N_10404,N_8398,N_8894);
or U10405 (N_10405,N_8968,N_6184);
nand U10406 (N_10406,N_7415,N_7855);
xor U10407 (N_10407,N_6285,N_8794);
or U10408 (N_10408,N_8704,N_8547);
nor U10409 (N_10409,N_6941,N_6165);
nor U10410 (N_10410,N_6058,N_7364);
nor U10411 (N_10411,N_6796,N_6466);
and U10412 (N_10412,N_6023,N_7178);
nand U10413 (N_10413,N_6978,N_7004);
or U10414 (N_10414,N_6158,N_7100);
nand U10415 (N_10415,N_6756,N_7384);
or U10416 (N_10416,N_8159,N_8713);
nand U10417 (N_10417,N_6695,N_6522);
nor U10418 (N_10418,N_6545,N_7673);
xor U10419 (N_10419,N_6342,N_8869);
nand U10420 (N_10420,N_6907,N_8079);
nand U10421 (N_10421,N_6088,N_6396);
nor U10422 (N_10422,N_7135,N_6209);
and U10423 (N_10423,N_7339,N_8014);
nand U10424 (N_10424,N_8220,N_7903);
xnor U10425 (N_10425,N_8514,N_6034);
nand U10426 (N_10426,N_7844,N_8310);
or U10427 (N_10427,N_7406,N_7083);
xnor U10428 (N_10428,N_8217,N_7564);
nor U10429 (N_10429,N_7270,N_8997);
nand U10430 (N_10430,N_6079,N_7263);
and U10431 (N_10431,N_6070,N_6957);
nor U10432 (N_10432,N_6896,N_8749);
nor U10433 (N_10433,N_7663,N_8848);
nor U10434 (N_10434,N_8464,N_7410);
nor U10435 (N_10435,N_6085,N_6280);
nand U10436 (N_10436,N_6491,N_6939);
or U10437 (N_10437,N_6084,N_8954);
nand U10438 (N_10438,N_7611,N_6787);
nand U10439 (N_10439,N_6583,N_8734);
nand U10440 (N_10440,N_6641,N_7482);
or U10441 (N_10441,N_8720,N_6297);
nor U10442 (N_10442,N_6066,N_7907);
nand U10443 (N_10443,N_7029,N_7760);
or U10444 (N_10444,N_6779,N_7442);
xnor U10445 (N_10445,N_6223,N_6645);
xnor U10446 (N_10446,N_6938,N_6563);
xor U10447 (N_10447,N_8843,N_7193);
and U10448 (N_10448,N_6955,N_6694);
and U10449 (N_10449,N_6928,N_7454);
nor U10450 (N_10450,N_8218,N_6387);
nand U10451 (N_10451,N_7373,N_8895);
and U10452 (N_10452,N_7034,N_6311);
and U10453 (N_10453,N_8702,N_7826);
nand U10454 (N_10454,N_8282,N_7141);
or U10455 (N_10455,N_6732,N_7277);
xor U10456 (N_10456,N_6167,N_7908);
xor U10457 (N_10457,N_6044,N_7934);
nor U10458 (N_10458,N_6594,N_8296);
xor U10459 (N_10459,N_6577,N_7507);
nand U10460 (N_10460,N_8368,N_7878);
nor U10461 (N_10461,N_6912,N_6136);
and U10462 (N_10462,N_7489,N_7453);
xnor U10463 (N_10463,N_7063,N_7440);
and U10464 (N_10464,N_6835,N_6093);
nand U10465 (N_10465,N_6425,N_6560);
or U10466 (N_10466,N_7072,N_6132);
xor U10467 (N_10467,N_8434,N_6926);
nand U10468 (N_10468,N_7842,N_8807);
xor U10469 (N_10469,N_8228,N_7841);
nand U10470 (N_10470,N_8069,N_7187);
nand U10471 (N_10471,N_8335,N_7635);
xor U10472 (N_10472,N_6435,N_8395);
nand U10473 (N_10473,N_8597,N_8110);
nand U10474 (N_10474,N_8128,N_6590);
nor U10475 (N_10475,N_8891,N_7241);
or U10476 (N_10476,N_6336,N_7853);
nor U10477 (N_10477,N_7213,N_7060);
xnor U10478 (N_10478,N_6727,N_6138);
and U10479 (N_10479,N_7585,N_8761);
nand U10480 (N_10480,N_7353,N_6072);
xor U10481 (N_10481,N_8885,N_6786);
xnor U10482 (N_10482,N_7416,N_7687);
or U10483 (N_10483,N_6118,N_6905);
nand U10484 (N_10484,N_6470,N_7874);
nand U10485 (N_10485,N_6473,N_7696);
nor U10486 (N_10486,N_8363,N_7653);
nand U10487 (N_10487,N_8287,N_8513);
nor U10488 (N_10488,N_7313,N_7830);
nand U10489 (N_10489,N_8180,N_8512);
and U10490 (N_10490,N_7694,N_6647);
or U10491 (N_10491,N_6744,N_8177);
nand U10492 (N_10492,N_6800,N_7539);
and U10493 (N_10493,N_6865,N_7043);
nand U10494 (N_10494,N_8002,N_7276);
or U10495 (N_10495,N_8246,N_8680);
xnor U10496 (N_10496,N_7684,N_8284);
nor U10497 (N_10497,N_8458,N_6483);
or U10498 (N_10498,N_6534,N_8065);
nand U10499 (N_10499,N_7333,N_7109);
and U10500 (N_10500,N_7579,N_6331);
xnor U10501 (N_10501,N_8065,N_6201);
xnor U10502 (N_10502,N_7219,N_7198);
nand U10503 (N_10503,N_6394,N_6063);
nor U10504 (N_10504,N_6001,N_7649);
nor U10505 (N_10505,N_8809,N_8733);
or U10506 (N_10506,N_8493,N_8094);
or U10507 (N_10507,N_6147,N_6370);
nor U10508 (N_10508,N_7304,N_7141);
and U10509 (N_10509,N_8959,N_7549);
nand U10510 (N_10510,N_7668,N_6960);
or U10511 (N_10511,N_8487,N_8623);
nor U10512 (N_10512,N_8444,N_7621);
or U10513 (N_10513,N_8802,N_7250);
and U10514 (N_10514,N_7329,N_8737);
nand U10515 (N_10515,N_7117,N_6805);
and U10516 (N_10516,N_6487,N_6787);
or U10517 (N_10517,N_6579,N_6823);
nor U10518 (N_10518,N_7454,N_8843);
or U10519 (N_10519,N_8210,N_8071);
or U10520 (N_10520,N_8506,N_8841);
xnor U10521 (N_10521,N_8657,N_6089);
and U10522 (N_10522,N_7672,N_6900);
or U10523 (N_10523,N_7083,N_7989);
and U10524 (N_10524,N_8892,N_8003);
and U10525 (N_10525,N_7285,N_6307);
nand U10526 (N_10526,N_7353,N_6483);
and U10527 (N_10527,N_7303,N_7333);
or U10528 (N_10528,N_7054,N_6775);
or U10529 (N_10529,N_8098,N_6219);
and U10530 (N_10530,N_6581,N_8515);
or U10531 (N_10531,N_8003,N_6031);
or U10532 (N_10532,N_6984,N_6292);
nor U10533 (N_10533,N_7264,N_6316);
nor U10534 (N_10534,N_8285,N_8563);
xor U10535 (N_10535,N_7748,N_8200);
nor U10536 (N_10536,N_7883,N_8158);
xnor U10537 (N_10537,N_6343,N_6926);
xnor U10538 (N_10538,N_6443,N_6708);
nand U10539 (N_10539,N_8674,N_7866);
and U10540 (N_10540,N_7629,N_8293);
nand U10541 (N_10541,N_8348,N_7416);
or U10542 (N_10542,N_6542,N_7558);
nor U10543 (N_10543,N_6717,N_6170);
or U10544 (N_10544,N_6706,N_8296);
nor U10545 (N_10545,N_8176,N_6742);
nand U10546 (N_10546,N_7012,N_7225);
and U10547 (N_10547,N_6683,N_7523);
xnor U10548 (N_10548,N_7779,N_6314);
nor U10549 (N_10549,N_8675,N_6137);
nand U10550 (N_10550,N_7733,N_6567);
and U10551 (N_10551,N_6619,N_8632);
or U10552 (N_10552,N_8498,N_8397);
or U10553 (N_10553,N_6241,N_8426);
nor U10554 (N_10554,N_8368,N_7561);
nor U10555 (N_10555,N_6640,N_8519);
xor U10556 (N_10556,N_8651,N_7035);
and U10557 (N_10557,N_7855,N_7024);
or U10558 (N_10558,N_7277,N_7616);
nor U10559 (N_10559,N_6875,N_6144);
nor U10560 (N_10560,N_7907,N_8913);
or U10561 (N_10561,N_6543,N_6300);
xor U10562 (N_10562,N_6287,N_7247);
or U10563 (N_10563,N_7529,N_6100);
and U10564 (N_10564,N_6529,N_7080);
or U10565 (N_10565,N_8174,N_8058);
nand U10566 (N_10566,N_7001,N_8679);
nand U10567 (N_10567,N_8616,N_8266);
and U10568 (N_10568,N_7361,N_6223);
or U10569 (N_10569,N_6698,N_8794);
and U10570 (N_10570,N_7459,N_7447);
nor U10571 (N_10571,N_7733,N_7634);
xor U10572 (N_10572,N_6448,N_8033);
or U10573 (N_10573,N_6447,N_8058);
nand U10574 (N_10574,N_6436,N_8191);
nand U10575 (N_10575,N_6366,N_6982);
or U10576 (N_10576,N_6922,N_6328);
nand U10577 (N_10577,N_6901,N_7160);
nor U10578 (N_10578,N_7318,N_6871);
xor U10579 (N_10579,N_7449,N_8421);
and U10580 (N_10580,N_6228,N_6107);
nand U10581 (N_10581,N_6533,N_6817);
nor U10582 (N_10582,N_7177,N_7329);
or U10583 (N_10583,N_7293,N_8335);
xor U10584 (N_10584,N_7439,N_8264);
nor U10585 (N_10585,N_7961,N_7775);
or U10586 (N_10586,N_7884,N_8556);
nand U10587 (N_10587,N_7610,N_6374);
nand U10588 (N_10588,N_6420,N_7347);
or U10589 (N_10589,N_8650,N_8365);
or U10590 (N_10590,N_8856,N_7235);
or U10591 (N_10591,N_7068,N_6230);
nand U10592 (N_10592,N_6056,N_8631);
and U10593 (N_10593,N_7619,N_6258);
nand U10594 (N_10594,N_7985,N_6108);
nand U10595 (N_10595,N_7567,N_6776);
nand U10596 (N_10596,N_6453,N_7368);
nand U10597 (N_10597,N_6072,N_6384);
nand U10598 (N_10598,N_8527,N_7344);
and U10599 (N_10599,N_7116,N_6497);
nand U10600 (N_10600,N_8735,N_7865);
or U10601 (N_10601,N_7400,N_8269);
nor U10602 (N_10602,N_8007,N_8832);
nor U10603 (N_10603,N_8974,N_6959);
xnor U10604 (N_10604,N_7827,N_7090);
and U10605 (N_10605,N_8447,N_6096);
or U10606 (N_10606,N_6868,N_6545);
nor U10607 (N_10607,N_7613,N_8706);
nand U10608 (N_10608,N_6951,N_7026);
nor U10609 (N_10609,N_8256,N_7811);
nor U10610 (N_10610,N_6264,N_7558);
nor U10611 (N_10611,N_7365,N_7392);
and U10612 (N_10612,N_7320,N_8548);
or U10613 (N_10613,N_7535,N_7424);
and U10614 (N_10614,N_7874,N_6912);
and U10615 (N_10615,N_7940,N_8315);
nor U10616 (N_10616,N_6508,N_7917);
nor U10617 (N_10617,N_6541,N_7243);
nor U10618 (N_10618,N_8334,N_6209);
nor U10619 (N_10619,N_7659,N_7554);
nor U10620 (N_10620,N_8958,N_6367);
nand U10621 (N_10621,N_6932,N_6245);
or U10622 (N_10622,N_6784,N_6919);
nor U10623 (N_10623,N_8354,N_8953);
or U10624 (N_10624,N_6795,N_7332);
xnor U10625 (N_10625,N_8588,N_8247);
nor U10626 (N_10626,N_8514,N_8614);
nand U10627 (N_10627,N_8308,N_6259);
nor U10628 (N_10628,N_7589,N_7402);
or U10629 (N_10629,N_8287,N_6158);
or U10630 (N_10630,N_6646,N_7153);
nand U10631 (N_10631,N_8137,N_8705);
nor U10632 (N_10632,N_8702,N_8811);
nor U10633 (N_10633,N_7756,N_7229);
xnor U10634 (N_10634,N_8171,N_6039);
nand U10635 (N_10635,N_6687,N_7171);
or U10636 (N_10636,N_6916,N_6400);
nor U10637 (N_10637,N_6392,N_8467);
or U10638 (N_10638,N_8807,N_6810);
nand U10639 (N_10639,N_8845,N_6353);
xnor U10640 (N_10640,N_8284,N_8779);
and U10641 (N_10641,N_7264,N_7066);
nor U10642 (N_10642,N_6705,N_7116);
nor U10643 (N_10643,N_8626,N_7708);
nand U10644 (N_10644,N_7384,N_8198);
nor U10645 (N_10645,N_6564,N_7236);
and U10646 (N_10646,N_8261,N_7842);
nand U10647 (N_10647,N_8158,N_6011);
nand U10648 (N_10648,N_6299,N_7806);
or U10649 (N_10649,N_8944,N_8534);
nor U10650 (N_10650,N_8979,N_6997);
or U10651 (N_10651,N_8405,N_7535);
and U10652 (N_10652,N_8840,N_7295);
or U10653 (N_10653,N_8434,N_7302);
and U10654 (N_10654,N_8445,N_7580);
and U10655 (N_10655,N_7006,N_7196);
nor U10656 (N_10656,N_8033,N_8413);
or U10657 (N_10657,N_6368,N_6860);
nor U10658 (N_10658,N_8901,N_8153);
xnor U10659 (N_10659,N_7026,N_6335);
nand U10660 (N_10660,N_6495,N_6121);
xor U10661 (N_10661,N_8974,N_8634);
nand U10662 (N_10662,N_6603,N_7209);
xnor U10663 (N_10663,N_6477,N_8154);
or U10664 (N_10664,N_7842,N_6582);
xnor U10665 (N_10665,N_8972,N_8750);
and U10666 (N_10666,N_6794,N_8239);
and U10667 (N_10667,N_8791,N_7643);
and U10668 (N_10668,N_7654,N_8969);
xor U10669 (N_10669,N_8843,N_6978);
xor U10670 (N_10670,N_7762,N_7810);
xor U10671 (N_10671,N_6636,N_8684);
xnor U10672 (N_10672,N_7278,N_7125);
nand U10673 (N_10673,N_8829,N_6936);
nand U10674 (N_10674,N_7179,N_7400);
or U10675 (N_10675,N_8921,N_6413);
or U10676 (N_10676,N_8591,N_7467);
xnor U10677 (N_10677,N_8728,N_7218);
or U10678 (N_10678,N_8355,N_8128);
nor U10679 (N_10679,N_8698,N_8196);
nor U10680 (N_10680,N_7314,N_7654);
and U10681 (N_10681,N_8350,N_7353);
and U10682 (N_10682,N_8225,N_7299);
nand U10683 (N_10683,N_6845,N_8582);
or U10684 (N_10684,N_7897,N_7670);
nand U10685 (N_10685,N_6890,N_8015);
nor U10686 (N_10686,N_6924,N_6791);
xor U10687 (N_10687,N_6365,N_7818);
xor U10688 (N_10688,N_8459,N_6018);
xnor U10689 (N_10689,N_8458,N_6254);
or U10690 (N_10690,N_7635,N_6378);
nor U10691 (N_10691,N_8301,N_8124);
and U10692 (N_10692,N_8726,N_6279);
and U10693 (N_10693,N_7877,N_7679);
or U10694 (N_10694,N_6597,N_6189);
nor U10695 (N_10695,N_6486,N_7744);
nor U10696 (N_10696,N_8759,N_7533);
xnor U10697 (N_10697,N_6865,N_7624);
xor U10698 (N_10698,N_6642,N_8346);
nand U10699 (N_10699,N_8921,N_6614);
nor U10700 (N_10700,N_6730,N_8604);
nand U10701 (N_10701,N_8778,N_8893);
xnor U10702 (N_10702,N_8516,N_8931);
xnor U10703 (N_10703,N_7673,N_8488);
xor U10704 (N_10704,N_7617,N_6735);
xnor U10705 (N_10705,N_6493,N_6978);
xnor U10706 (N_10706,N_7369,N_6635);
or U10707 (N_10707,N_8608,N_7161);
and U10708 (N_10708,N_7122,N_8124);
nor U10709 (N_10709,N_8343,N_8039);
and U10710 (N_10710,N_8435,N_7062);
or U10711 (N_10711,N_8388,N_7171);
and U10712 (N_10712,N_8903,N_7400);
nand U10713 (N_10713,N_7920,N_8288);
and U10714 (N_10714,N_7310,N_7964);
nor U10715 (N_10715,N_6593,N_6800);
and U10716 (N_10716,N_8938,N_8200);
nor U10717 (N_10717,N_6369,N_6030);
nor U10718 (N_10718,N_8806,N_8295);
nor U10719 (N_10719,N_8816,N_8459);
xor U10720 (N_10720,N_6610,N_7365);
nand U10721 (N_10721,N_8952,N_8491);
nand U10722 (N_10722,N_6981,N_8750);
or U10723 (N_10723,N_8837,N_7638);
and U10724 (N_10724,N_8161,N_7247);
and U10725 (N_10725,N_7223,N_6604);
or U10726 (N_10726,N_7414,N_7870);
or U10727 (N_10727,N_7059,N_6848);
xnor U10728 (N_10728,N_7895,N_7650);
and U10729 (N_10729,N_8633,N_8866);
nand U10730 (N_10730,N_8052,N_7233);
nand U10731 (N_10731,N_7306,N_6786);
nor U10732 (N_10732,N_7974,N_8246);
xnor U10733 (N_10733,N_6320,N_8322);
nand U10734 (N_10734,N_6479,N_7289);
nor U10735 (N_10735,N_6081,N_8444);
and U10736 (N_10736,N_8672,N_8780);
nand U10737 (N_10737,N_8732,N_6792);
nor U10738 (N_10738,N_8981,N_7457);
xnor U10739 (N_10739,N_6473,N_8462);
and U10740 (N_10740,N_8624,N_7247);
or U10741 (N_10741,N_6624,N_6905);
nor U10742 (N_10742,N_6049,N_6399);
and U10743 (N_10743,N_6376,N_8566);
nand U10744 (N_10744,N_6090,N_8381);
xor U10745 (N_10745,N_8759,N_6774);
or U10746 (N_10746,N_6200,N_6923);
and U10747 (N_10747,N_7105,N_7844);
nor U10748 (N_10748,N_6840,N_7262);
nand U10749 (N_10749,N_7818,N_8199);
nor U10750 (N_10750,N_7867,N_8545);
xnor U10751 (N_10751,N_7278,N_7256);
xnor U10752 (N_10752,N_7548,N_6574);
xor U10753 (N_10753,N_8842,N_8887);
nor U10754 (N_10754,N_8131,N_8655);
or U10755 (N_10755,N_7999,N_7285);
xnor U10756 (N_10756,N_8566,N_7002);
nor U10757 (N_10757,N_6112,N_7734);
xnor U10758 (N_10758,N_8731,N_7421);
nor U10759 (N_10759,N_7206,N_8677);
or U10760 (N_10760,N_6969,N_6505);
and U10761 (N_10761,N_7637,N_6036);
xor U10762 (N_10762,N_7877,N_6436);
nand U10763 (N_10763,N_6703,N_7639);
and U10764 (N_10764,N_8280,N_7046);
xnor U10765 (N_10765,N_6886,N_6055);
and U10766 (N_10766,N_6929,N_7003);
xnor U10767 (N_10767,N_6324,N_8012);
and U10768 (N_10768,N_7141,N_6741);
nor U10769 (N_10769,N_6287,N_8386);
nand U10770 (N_10770,N_6632,N_6303);
and U10771 (N_10771,N_8010,N_8384);
or U10772 (N_10772,N_7179,N_7845);
or U10773 (N_10773,N_7348,N_7372);
nand U10774 (N_10774,N_6433,N_6867);
xnor U10775 (N_10775,N_7446,N_6463);
or U10776 (N_10776,N_6705,N_6260);
xnor U10777 (N_10777,N_7538,N_8566);
or U10778 (N_10778,N_7516,N_7175);
xnor U10779 (N_10779,N_7934,N_7403);
xor U10780 (N_10780,N_8399,N_8295);
or U10781 (N_10781,N_6528,N_8775);
nand U10782 (N_10782,N_6498,N_7049);
nand U10783 (N_10783,N_7313,N_6893);
xnor U10784 (N_10784,N_7768,N_6443);
nand U10785 (N_10785,N_6497,N_8831);
nand U10786 (N_10786,N_8931,N_8937);
xor U10787 (N_10787,N_7527,N_8206);
or U10788 (N_10788,N_8064,N_8758);
nor U10789 (N_10789,N_6655,N_6829);
nor U10790 (N_10790,N_8163,N_6834);
nor U10791 (N_10791,N_7731,N_6514);
or U10792 (N_10792,N_6553,N_7665);
nand U10793 (N_10793,N_6725,N_6372);
or U10794 (N_10794,N_6137,N_7748);
and U10795 (N_10795,N_6451,N_8858);
nand U10796 (N_10796,N_7039,N_7560);
nand U10797 (N_10797,N_8302,N_6131);
and U10798 (N_10798,N_6682,N_8794);
xnor U10799 (N_10799,N_8922,N_8082);
nor U10800 (N_10800,N_8002,N_8272);
or U10801 (N_10801,N_8754,N_7302);
nor U10802 (N_10802,N_6464,N_6495);
nand U10803 (N_10803,N_8080,N_6681);
nand U10804 (N_10804,N_8192,N_8813);
nor U10805 (N_10805,N_8574,N_6721);
nor U10806 (N_10806,N_6226,N_7672);
and U10807 (N_10807,N_7633,N_6631);
xor U10808 (N_10808,N_8348,N_8294);
nand U10809 (N_10809,N_7525,N_6334);
nor U10810 (N_10810,N_6872,N_6597);
nor U10811 (N_10811,N_8518,N_6988);
and U10812 (N_10812,N_7117,N_7429);
nor U10813 (N_10813,N_7408,N_7318);
nand U10814 (N_10814,N_7334,N_8505);
nor U10815 (N_10815,N_6411,N_8394);
xor U10816 (N_10816,N_7178,N_8398);
nand U10817 (N_10817,N_8751,N_6630);
and U10818 (N_10818,N_6074,N_7035);
or U10819 (N_10819,N_7467,N_6340);
nand U10820 (N_10820,N_7991,N_8687);
and U10821 (N_10821,N_8145,N_7831);
and U10822 (N_10822,N_8007,N_8889);
or U10823 (N_10823,N_6823,N_6376);
nand U10824 (N_10824,N_8513,N_7601);
or U10825 (N_10825,N_8301,N_8867);
nor U10826 (N_10826,N_6410,N_8132);
and U10827 (N_10827,N_8291,N_8866);
nor U10828 (N_10828,N_8740,N_7363);
xnor U10829 (N_10829,N_7590,N_8921);
or U10830 (N_10830,N_6829,N_7828);
xnor U10831 (N_10831,N_7350,N_6525);
and U10832 (N_10832,N_7104,N_6218);
xnor U10833 (N_10833,N_8150,N_6656);
nand U10834 (N_10834,N_6884,N_7556);
xnor U10835 (N_10835,N_8956,N_7324);
or U10836 (N_10836,N_8075,N_6306);
nand U10837 (N_10837,N_6426,N_7949);
or U10838 (N_10838,N_8487,N_7826);
nand U10839 (N_10839,N_8165,N_8692);
or U10840 (N_10840,N_7661,N_6445);
and U10841 (N_10841,N_7091,N_8221);
nand U10842 (N_10842,N_7815,N_6208);
xnor U10843 (N_10843,N_6225,N_7070);
or U10844 (N_10844,N_6767,N_8722);
nor U10845 (N_10845,N_8520,N_8099);
or U10846 (N_10846,N_8506,N_7266);
nand U10847 (N_10847,N_7997,N_8293);
nand U10848 (N_10848,N_7095,N_6932);
or U10849 (N_10849,N_8103,N_8775);
and U10850 (N_10850,N_6586,N_6880);
xnor U10851 (N_10851,N_6173,N_7166);
nor U10852 (N_10852,N_8300,N_6309);
nand U10853 (N_10853,N_6470,N_8548);
and U10854 (N_10854,N_8332,N_6328);
or U10855 (N_10855,N_6310,N_6839);
and U10856 (N_10856,N_8016,N_7567);
xor U10857 (N_10857,N_6584,N_8873);
or U10858 (N_10858,N_8840,N_8120);
or U10859 (N_10859,N_7387,N_8725);
and U10860 (N_10860,N_7444,N_7583);
nand U10861 (N_10861,N_6004,N_6956);
xnor U10862 (N_10862,N_6152,N_6101);
or U10863 (N_10863,N_6398,N_8047);
and U10864 (N_10864,N_6057,N_6834);
or U10865 (N_10865,N_8018,N_7932);
and U10866 (N_10866,N_6938,N_8031);
nor U10867 (N_10867,N_8877,N_7558);
nand U10868 (N_10868,N_6113,N_7550);
or U10869 (N_10869,N_8169,N_8235);
xnor U10870 (N_10870,N_8461,N_6937);
nand U10871 (N_10871,N_7216,N_6159);
or U10872 (N_10872,N_7162,N_6596);
and U10873 (N_10873,N_8832,N_6769);
nand U10874 (N_10874,N_7108,N_6407);
nor U10875 (N_10875,N_7456,N_8638);
or U10876 (N_10876,N_8009,N_7730);
nor U10877 (N_10877,N_7490,N_7063);
or U10878 (N_10878,N_8895,N_7484);
and U10879 (N_10879,N_6882,N_6205);
nand U10880 (N_10880,N_8925,N_8028);
or U10881 (N_10881,N_6378,N_8070);
or U10882 (N_10882,N_6284,N_7649);
or U10883 (N_10883,N_7669,N_7225);
nand U10884 (N_10884,N_8661,N_8562);
and U10885 (N_10885,N_7443,N_8386);
nand U10886 (N_10886,N_8052,N_8673);
nand U10887 (N_10887,N_7383,N_7155);
nor U10888 (N_10888,N_8342,N_6549);
or U10889 (N_10889,N_7464,N_8469);
or U10890 (N_10890,N_8515,N_8458);
nand U10891 (N_10891,N_8662,N_7624);
and U10892 (N_10892,N_6697,N_6086);
nand U10893 (N_10893,N_8051,N_8256);
and U10894 (N_10894,N_8902,N_8931);
and U10895 (N_10895,N_6114,N_8439);
and U10896 (N_10896,N_7124,N_8044);
nand U10897 (N_10897,N_6482,N_6695);
nand U10898 (N_10898,N_7578,N_6337);
nand U10899 (N_10899,N_8622,N_8796);
and U10900 (N_10900,N_8221,N_6183);
nand U10901 (N_10901,N_8116,N_8070);
or U10902 (N_10902,N_6343,N_8829);
nand U10903 (N_10903,N_6525,N_7565);
nor U10904 (N_10904,N_6965,N_6018);
nor U10905 (N_10905,N_7995,N_6468);
or U10906 (N_10906,N_7226,N_6462);
and U10907 (N_10907,N_8258,N_7586);
nand U10908 (N_10908,N_7530,N_7656);
or U10909 (N_10909,N_6899,N_6212);
nand U10910 (N_10910,N_6905,N_6882);
or U10911 (N_10911,N_8402,N_8870);
nor U10912 (N_10912,N_8400,N_8712);
xnor U10913 (N_10913,N_6305,N_7888);
or U10914 (N_10914,N_8616,N_7407);
xor U10915 (N_10915,N_7941,N_8544);
xor U10916 (N_10916,N_6920,N_7364);
xnor U10917 (N_10917,N_6016,N_6672);
nand U10918 (N_10918,N_6527,N_7144);
xor U10919 (N_10919,N_7828,N_7840);
nand U10920 (N_10920,N_7593,N_7296);
nor U10921 (N_10921,N_7437,N_6972);
nand U10922 (N_10922,N_8708,N_6519);
nand U10923 (N_10923,N_8362,N_6423);
and U10924 (N_10924,N_7417,N_8067);
and U10925 (N_10925,N_8199,N_7530);
nand U10926 (N_10926,N_8493,N_8866);
nand U10927 (N_10927,N_7835,N_7697);
and U10928 (N_10928,N_6401,N_8356);
or U10929 (N_10929,N_7692,N_7515);
nand U10930 (N_10930,N_6226,N_8249);
nor U10931 (N_10931,N_7515,N_8444);
nor U10932 (N_10932,N_8084,N_8440);
and U10933 (N_10933,N_7542,N_7999);
or U10934 (N_10934,N_8145,N_6671);
or U10935 (N_10935,N_6271,N_8533);
xnor U10936 (N_10936,N_8911,N_7301);
and U10937 (N_10937,N_7738,N_8862);
xnor U10938 (N_10938,N_6996,N_7213);
and U10939 (N_10939,N_8575,N_8947);
or U10940 (N_10940,N_7080,N_6995);
nor U10941 (N_10941,N_8614,N_7397);
nand U10942 (N_10942,N_7520,N_6267);
nor U10943 (N_10943,N_8341,N_8196);
nor U10944 (N_10944,N_7536,N_6532);
nor U10945 (N_10945,N_6378,N_7925);
or U10946 (N_10946,N_7699,N_7043);
or U10947 (N_10947,N_8952,N_8134);
nand U10948 (N_10948,N_8592,N_7490);
nor U10949 (N_10949,N_8388,N_7396);
and U10950 (N_10950,N_7661,N_6421);
nor U10951 (N_10951,N_7040,N_8879);
and U10952 (N_10952,N_8761,N_8647);
xnor U10953 (N_10953,N_6492,N_8806);
and U10954 (N_10954,N_8518,N_6948);
nand U10955 (N_10955,N_7780,N_6471);
or U10956 (N_10956,N_6161,N_6904);
nand U10957 (N_10957,N_7108,N_7031);
or U10958 (N_10958,N_7995,N_6711);
nand U10959 (N_10959,N_7605,N_7094);
and U10960 (N_10960,N_7610,N_6873);
or U10961 (N_10961,N_8221,N_6003);
and U10962 (N_10962,N_8186,N_7595);
nor U10963 (N_10963,N_7821,N_6723);
xnor U10964 (N_10964,N_7058,N_6769);
nor U10965 (N_10965,N_6569,N_6095);
nor U10966 (N_10966,N_7992,N_8730);
or U10967 (N_10967,N_8305,N_6084);
nand U10968 (N_10968,N_7828,N_8092);
xor U10969 (N_10969,N_7429,N_6330);
or U10970 (N_10970,N_6895,N_6893);
and U10971 (N_10971,N_8268,N_8333);
and U10972 (N_10972,N_7395,N_7267);
and U10973 (N_10973,N_8716,N_7906);
and U10974 (N_10974,N_7547,N_6169);
or U10975 (N_10975,N_6046,N_6620);
xor U10976 (N_10976,N_7966,N_6345);
xor U10977 (N_10977,N_7686,N_8484);
or U10978 (N_10978,N_7766,N_8539);
xor U10979 (N_10979,N_6329,N_8407);
nor U10980 (N_10980,N_8181,N_6141);
xor U10981 (N_10981,N_7577,N_7056);
or U10982 (N_10982,N_8677,N_7764);
nor U10983 (N_10983,N_8340,N_7856);
or U10984 (N_10984,N_8796,N_8970);
xor U10985 (N_10985,N_6003,N_6947);
or U10986 (N_10986,N_8055,N_8622);
or U10987 (N_10987,N_7706,N_8709);
and U10988 (N_10988,N_8849,N_7297);
xor U10989 (N_10989,N_7437,N_6940);
nand U10990 (N_10990,N_7148,N_8542);
and U10991 (N_10991,N_8479,N_8139);
or U10992 (N_10992,N_7227,N_8112);
nor U10993 (N_10993,N_8780,N_6745);
xor U10994 (N_10994,N_8071,N_8606);
and U10995 (N_10995,N_6553,N_8832);
nand U10996 (N_10996,N_6220,N_8900);
or U10997 (N_10997,N_8200,N_8532);
nand U10998 (N_10998,N_8266,N_8959);
xor U10999 (N_10999,N_8960,N_7511);
nand U11000 (N_11000,N_7034,N_6334);
and U11001 (N_11001,N_7080,N_6937);
nor U11002 (N_11002,N_7466,N_8685);
nor U11003 (N_11003,N_6487,N_7809);
and U11004 (N_11004,N_6125,N_8294);
nor U11005 (N_11005,N_8757,N_6172);
and U11006 (N_11006,N_6874,N_6479);
xor U11007 (N_11007,N_6342,N_7795);
and U11008 (N_11008,N_8976,N_7536);
xor U11009 (N_11009,N_8530,N_7604);
or U11010 (N_11010,N_7860,N_8499);
or U11011 (N_11011,N_7106,N_7989);
or U11012 (N_11012,N_7055,N_8687);
or U11013 (N_11013,N_6750,N_6973);
nand U11014 (N_11014,N_8881,N_7032);
or U11015 (N_11015,N_8611,N_8897);
nor U11016 (N_11016,N_7122,N_6207);
or U11017 (N_11017,N_7288,N_6303);
or U11018 (N_11018,N_7915,N_6605);
or U11019 (N_11019,N_6175,N_8212);
nand U11020 (N_11020,N_7865,N_7273);
nand U11021 (N_11021,N_8495,N_6723);
or U11022 (N_11022,N_6736,N_7908);
nor U11023 (N_11023,N_6623,N_7252);
or U11024 (N_11024,N_7835,N_7654);
or U11025 (N_11025,N_6107,N_7049);
xor U11026 (N_11026,N_8112,N_6771);
and U11027 (N_11027,N_8049,N_7365);
xor U11028 (N_11028,N_8949,N_7868);
nand U11029 (N_11029,N_8522,N_8845);
nor U11030 (N_11030,N_7792,N_7229);
xnor U11031 (N_11031,N_6015,N_7911);
or U11032 (N_11032,N_7226,N_7461);
or U11033 (N_11033,N_7804,N_8066);
nor U11034 (N_11034,N_6133,N_6003);
or U11035 (N_11035,N_6097,N_7124);
xor U11036 (N_11036,N_8292,N_8490);
nor U11037 (N_11037,N_8412,N_8466);
and U11038 (N_11038,N_6359,N_6346);
nand U11039 (N_11039,N_7896,N_8932);
and U11040 (N_11040,N_6727,N_7990);
xnor U11041 (N_11041,N_6652,N_6794);
xnor U11042 (N_11042,N_6673,N_8520);
nor U11043 (N_11043,N_8637,N_8793);
nor U11044 (N_11044,N_6823,N_8343);
nor U11045 (N_11045,N_6358,N_6269);
and U11046 (N_11046,N_7523,N_8435);
xnor U11047 (N_11047,N_6493,N_6691);
xor U11048 (N_11048,N_7314,N_7431);
and U11049 (N_11049,N_6403,N_6687);
and U11050 (N_11050,N_7568,N_7986);
nor U11051 (N_11051,N_6672,N_6423);
xor U11052 (N_11052,N_6939,N_8505);
nand U11053 (N_11053,N_8088,N_6252);
and U11054 (N_11054,N_7745,N_6702);
nand U11055 (N_11055,N_8605,N_7504);
nor U11056 (N_11056,N_8846,N_6985);
nor U11057 (N_11057,N_8658,N_6945);
or U11058 (N_11058,N_6094,N_7876);
or U11059 (N_11059,N_6645,N_6122);
and U11060 (N_11060,N_8065,N_7616);
nand U11061 (N_11061,N_7992,N_8430);
nor U11062 (N_11062,N_6752,N_6735);
nand U11063 (N_11063,N_7142,N_8008);
nand U11064 (N_11064,N_7259,N_7606);
xnor U11065 (N_11065,N_8144,N_8746);
and U11066 (N_11066,N_8809,N_7592);
or U11067 (N_11067,N_8149,N_7186);
nor U11068 (N_11068,N_7688,N_6761);
xnor U11069 (N_11069,N_7642,N_8994);
xor U11070 (N_11070,N_8746,N_6628);
nor U11071 (N_11071,N_8348,N_6728);
and U11072 (N_11072,N_6124,N_6747);
xnor U11073 (N_11073,N_6404,N_6102);
xnor U11074 (N_11074,N_7123,N_6059);
and U11075 (N_11075,N_7702,N_7722);
or U11076 (N_11076,N_7133,N_7117);
or U11077 (N_11077,N_6541,N_8552);
nand U11078 (N_11078,N_8801,N_8062);
nor U11079 (N_11079,N_7345,N_7728);
xor U11080 (N_11080,N_8745,N_7977);
or U11081 (N_11081,N_8692,N_8129);
nand U11082 (N_11082,N_8117,N_6535);
nand U11083 (N_11083,N_7770,N_6064);
nor U11084 (N_11084,N_6393,N_8114);
and U11085 (N_11085,N_7641,N_8458);
nor U11086 (N_11086,N_7781,N_7116);
xnor U11087 (N_11087,N_7895,N_7204);
nand U11088 (N_11088,N_8266,N_8352);
and U11089 (N_11089,N_8461,N_7810);
nor U11090 (N_11090,N_7949,N_8678);
or U11091 (N_11091,N_6512,N_7963);
or U11092 (N_11092,N_8099,N_6232);
or U11093 (N_11093,N_6313,N_6201);
or U11094 (N_11094,N_8974,N_8119);
xor U11095 (N_11095,N_6778,N_6790);
nand U11096 (N_11096,N_6682,N_7388);
xor U11097 (N_11097,N_8445,N_6484);
and U11098 (N_11098,N_8345,N_8532);
and U11099 (N_11099,N_7430,N_7752);
and U11100 (N_11100,N_8594,N_8620);
or U11101 (N_11101,N_6563,N_6430);
and U11102 (N_11102,N_7928,N_8844);
nand U11103 (N_11103,N_7981,N_8948);
and U11104 (N_11104,N_6400,N_8910);
and U11105 (N_11105,N_7234,N_7882);
nand U11106 (N_11106,N_8405,N_8743);
nor U11107 (N_11107,N_6403,N_8414);
and U11108 (N_11108,N_6717,N_6073);
or U11109 (N_11109,N_6064,N_8448);
and U11110 (N_11110,N_8517,N_7818);
nand U11111 (N_11111,N_6303,N_7847);
nand U11112 (N_11112,N_8227,N_6109);
nand U11113 (N_11113,N_7185,N_6634);
and U11114 (N_11114,N_6353,N_6754);
xor U11115 (N_11115,N_8408,N_7945);
nor U11116 (N_11116,N_6314,N_8712);
nor U11117 (N_11117,N_7355,N_7698);
nand U11118 (N_11118,N_8701,N_6544);
and U11119 (N_11119,N_6574,N_7874);
nand U11120 (N_11120,N_6591,N_6095);
nor U11121 (N_11121,N_6832,N_8357);
xnor U11122 (N_11122,N_8998,N_6042);
or U11123 (N_11123,N_8079,N_7125);
xor U11124 (N_11124,N_6552,N_6656);
or U11125 (N_11125,N_7469,N_7034);
xnor U11126 (N_11126,N_7848,N_6046);
xnor U11127 (N_11127,N_6863,N_6284);
nand U11128 (N_11128,N_8726,N_8277);
and U11129 (N_11129,N_7738,N_8376);
and U11130 (N_11130,N_7796,N_6986);
xor U11131 (N_11131,N_7294,N_8019);
xor U11132 (N_11132,N_7605,N_8891);
xnor U11133 (N_11133,N_7729,N_6803);
xor U11134 (N_11134,N_7501,N_8100);
and U11135 (N_11135,N_6342,N_7891);
xor U11136 (N_11136,N_7358,N_6932);
and U11137 (N_11137,N_7353,N_8930);
nand U11138 (N_11138,N_6965,N_6857);
nor U11139 (N_11139,N_6226,N_7370);
and U11140 (N_11140,N_8142,N_6810);
and U11141 (N_11141,N_6448,N_8962);
nand U11142 (N_11142,N_8367,N_6551);
nand U11143 (N_11143,N_8052,N_6195);
and U11144 (N_11144,N_8680,N_6168);
nor U11145 (N_11145,N_8100,N_7444);
nor U11146 (N_11146,N_8546,N_8894);
nand U11147 (N_11147,N_8511,N_8542);
and U11148 (N_11148,N_6660,N_8227);
nor U11149 (N_11149,N_6436,N_8945);
nor U11150 (N_11150,N_8352,N_8512);
and U11151 (N_11151,N_8667,N_6190);
nor U11152 (N_11152,N_8916,N_6008);
xor U11153 (N_11153,N_6513,N_8879);
nor U11154 (N_11154,N_8357,N_6370);
xnor U11155 (N_11155,N_7676,N_6972);
nand U11156 (N_11156,N_8969,N_7176);
xor U11157 (N_11157,N_6244,N_6974);
or U11158 (N_11158,N_6231,N_8603);
and U11159 (N_11159,N_6634,N_7346);
and U11160 (N_11160,N_7444,N_6638);
xnor U11161 (N_11161,N_7569,N_6492);
or U11162 (N_11162,N_8533,N_6722);
nor U11163 (N_11163,N_6665,N_8935);
xnor U11164 (N_11164,N_7459,N_7545);
xor U11165 (N_11165,N_6161,N_6752);
nand U11166 (N_11166,N_6538,N_7335);
and U11167 (N_11167,N_6596,N_6780);
nand U11168 (N_11168,N_6777,N_6314);
nand U11169 (N_11169,N_7432,N_7763);
nor U11170 (N_11170,N_6299,N_8031);
xnor U11171 (N_11171,N_7427,N_7635);
xor U11172 (N_11172,N_8146,N_7586);
or U11173 (N_11173,N_8281,N_6949);
or U11174 (N_11174,N_6248,N_7135);
and U11175 (N_11175,N_6460,N_6726);
or U11176 (N_11176,N_7626,N_7013);
or U11177 (N_11177,N_8865,N_7006);
or U11178 (N_11178,N_8970,N_6922);
nand U11179 (N_11179,N_7591,N_7477);
nor U11180 (N_11180,N_8735,N_7160);
or U11181 (N_11181,N_7879,N_6820);
and U11182 (N_11182,N_6155,N_6144);
nor U11183 (N_11183,N_8815,N_6811);
xnor U11184 (N_11184,N_6574,N_8236);
nor U11185 (N_11185,N_8314,N_8477);
or U11186 (N_11186,N_6011,N_8219);
or U11187 (N_11187,N_7468,N_8769);
xor U11188 (N_11188,N_6690,N_6947);
and U11189 (N_11189,N_6779,N_8288);
and U11190 (N_11190,N_6382,N_7628);
xnor U11191 (N_11191,N_7416,N_7542);
and U11192 (N_11192,N_7135,N_8883);
nor U11193 (N_11193,N_6327,N_6943);
or U11194 (N_11194,N_6847,N_6988);
or U11195 (N_11195,N_8692,N_8282);
nand U11196 (N_11196,N_6790,N_8476);
nand U11197 (N_11197,N_7523,N_8483);
or U11198 (N_11198,N_7046,N_8586);
xnor U11199 (N_11199,N_6360,N_7525);
or U11200 (N_11200,N_6665,N_6124);
or U11201 (N_11201,N_6046,N_6230);
or U11202 (N_11202,N_6363,N_8201);
or U11203 (N_11203,N_6156,N_6030);
and U11204 (N_11204,N_7156,N_6297);
or U11205 (N_11205,N_8339,N_7309);
or U11206 (N_11206,N_6629,N_8158);
nand U11207 (N_11207,N_7567,N_6223);
nor U11208 (N_11208,N_6287,N_8381);
nand U11209 (N_11209,N_8808,N_7517);
xnor U11210 (N_11210,N_7212,N_8233);
nand U11211 (N_11211,N_7716,N_7492);
nor U11212 (N_11212,N_6971,N_8490);
xnor U11213 (N_11213,N_8570,N_7398);
nor U11214 (N_11214,N_8917,N_8534);
or U11215 (N_11215,N_6952,N_8992);
or U11216 (N_11216,N_7681,N_8876);
and U11217 (N_11217,N_7383,N_6925);
xnor U11218 (N_11218,N_6767,N_6893);
nor U11219 (N_11219,N_6525,N_6322);
nand U11220 (N_11220,N_7663,N_7965);
or U11221 (N_11221,N_8973,N_8411);
xor U11222 (N_11222,N_8906,N_8257);
xor U11223 (N_11223,N_6508,N_8016);
or U11224 (N_11224,N_7477,N_7674);
and U11225 (N_11225,N_6786,N_6211);
and U11226 (N_11226,N_7867,N_8213);
or U11227 (N_11227,N_7840,N_6639);
or U11228 (N_11228,N_8087,N_8360);
or U11229 (N_11229,N_6701,N_6122);
nand U11230 (N_11230,N_6401,N_6643);
nor U11231 (N_11231,N_8112,N_8939);
nor U11232 (N_11232,N_6244,N_6071);
or U11233 (N_11233,N_8672,N_8665);
nor U11234 (N_11234,N_7056,N_8627);
or U11235 (N_11235,N_6842,N_6191);
nor U11236 (N_11236,N_8050,N_8801);
or U11237 (N_11237,N_7184,N_8099);
nor U11238 (N_11238,N_8570,N_6631);
nor U11239 (N_11239,N_7704,N_7547);
nor U11240 (N_11240,N_8679,N_7507);
nand U11241 (N_11241,N_8364,N_6398);
nand U11242 (N_11242,N_8866,N_7328);
or U11243 (N_11243,N_7444,N_7095);
and U11244 (N_11244,N_7315,N_7946);
nand U11245 (N_11245,N_7540,N_6705);
and U11246 (N_11246,N_6720,N_6203);
nand U11247 (N_11247,N_7254,N_7976);
nor U11248 (N_11248,N_6187,N_8634);
nor U11249 (N_11249,N_6440,N_6269);
and U11250 (N_11250,N_8528,N_7435);
or U11251 (N_11251,N_7431,N_8179);
nand U11252 (N_11252,N_8318,N_7400);
or U11253 (N_11253,N_6883,N_7842);
and U11254 (N_11254,N_6986,N_7503);
or U11255 (N_11255,N_7186,N_7415);
and U11256 (N_11256,N_7656,N_7624);
and U11257 (N_11257,N_8108,N_7840);
and U11258 (N_11258,N_7783,N_8127);
or U11259 (N_11259,N_6238,N_6347);
xor U11260 (N_11260,N_8240,N_6093);
nor U11261 (N_11261,N_6948,N_8060);
nor U11262 (N_11262,N_8932,N_8584);
nor U11263 (N_11263,N_6792,N_6635);
xor U11264 (N_11264,N_7508,N_8325);
and U11265 (N_11265,N_7712,N_6754);
or U11266 (N_11266,N_7252,N_8648);
nand U11267 (N_11267,N_7555,N_8669);
nand U11268 (N_11268,N_8159,N_8274);
nand U11269 (N_11269,N_8878,N_8336);
and U11270 (N_11270,N_6295,N_7463);
or U11271 (N_11271,N_7044,N_6019);
nand U11272 (N_11272,N_6511,N_8231);
nand U11273 (N_11273,N_6410,N_8856);
and U11274 (N_11274,N_8324,N_7540);
and U11275 (N_11275,N_6779,N_7702);
xor U11276 (N_11276,N_7341,N_6850);
nand U11277 (N_11277,N_8703,N_6224);
nor U11278 (N_11278,N_8741,N_8928);
nor U11279 (N_11279,N_6094,N_7802);
nand U11280 (N_11280,N_6700,N_8876);
nand U11281 (N_11281,N_7987,N_8093);
or U11282 (N_11282,N_7326,N_7756);
nand U11283 (N_11283,N_6539,N_8528);
nand U11284 (N_11284,N_6706,N_7920);
nor U11285 (N_11285,N_6542,N_6745);
and U11286 (N_11286,N_7750,N_8646);
nand U11287 (N_11287,N_7333,N_7482);
nand U11288 (N_11288,N_6302,N_8994);
nand U11289 (N_11289,N_8428,N_7664);
xnor U11290 (N_11290,N_6452,N_8499);
nand U11291 (N_11291,N_6002,N_7923);
nor U11292 (N_11292,N_7496,N_8339);
and U11293 (N_11293,N_6367,N_7993);
or U11294 (N_11294,N_7583,N_7743);
nand U11295 (N_11295,N_8229,N_8857);
nand U11296 (N_11296,N_8362,N_8723);
xnor U11297 (N_11297,N_6794,N_8367);
xor U11298 (N_11298,N_8420,N_7212);
nand U11299 (N_11299,N_6025,N_7387);
nand U11300 (N_11300,N_8186,N_6874);
and U11301 (N_11301,N_6113,N_8167);
nor U11302 (N_11302,N_6934,N_8761);
xnor U11303 (N_11303,N_7922,N_6155);
nand U11304 (N_11304,N_6934,N_7343);
nand U11305 (N_11305,N_7958,N_6839);
nor U11306 (N_11306,N_6119,N_8398);
and U11307 (N_11307,N_8853,N_6858);
xnor U11308 (N_11308,N_7020,N_7090);
nand U11309 (N_11309,N_8403,N_6139);
nand U11310 (N_11310,N_7084,N_6884);
nand U11311 (N_11311,N_6853,N_7470);
nand U11312 (N_11312,N_6938,N_6627);
nor U11313 (N_11313,N_8855,N_7705);
nand U11314 (N_11314,N_7096,N_8387);
and U11315 (N_11315,N_7031,N_7818);
nand U11316 (N_11316,N_7218,N_7934);
nor U11317 (N_11317,N_8295,N_6893);
xor U11318 (N_11318,N_6854,N_8737);
or U11319 (N_11319,N_6039,N_7373);
nor U11320 (N_11320,N_8207,N_6573);
nor U11321 (N_11321,N_8211,N_7875);
and U11322 (N_11322,N_7484,N_7112);
and U11323 (N_11323,N_6214,N_7869);
nand U11324 (N_11324,N_6574,N_8395);
or U11325 (N_11325,N_6565,N_8695);
xnor U11326 (N_11326,N_7917,N_8571);
nand U11327 (N_11327,N_7461,N_6274);
nand U11328 (N_11328,N_6094,N_8896);
nor U11329 (N_11329,N_8243,N_6161);
nor U11330 (N_11330,N_7432,N_7926);
nand U11331 (N_11331,N_8800,N_7657);
and U11332 (N_11332,N_6307,N_6160);
nor U11333 (N_11333,N_7850,N_8220);
and U11334 (N_11334,N_6040,N_7126);
xnor U11335 (N_11335,N_6238,N_8282);
and U11336 (N_11336,N_7177,N_6924);
and U11337 (N_11337,N_6648,N_7934);
and U11338 (N_11338,N_6018,N_6824);
nor U11339 (N_11339,N_7701,N_6414);
or U11340 (N_11340,N_8486,N_6878);
xor U11341 (N_11341,N_6703,N_7526);
xnor U11342 (N_11342,N_7512,N_8398);
or U11343 (N_11343,N_8776,N_8678);
and U11344 (N_11344,N_6984,N_7406);
xor U11345 (N_11345,N_7723,N_8314);
xor U11346 (N_11346,N_8354,N_6254);
and U11347 (N_11347,N_7119,N_7131);
nand U11348 (N_11348,N_8546,N_8404);
nand U11349 (N_11349,N_8593,N_6016);
or U11350 (N_11350,N_7376,N_7057);
and U11351 (N_11351,N_6805,N_6185);
xor U11352 (N_11352,N_6742,N_7508);
nand U11353 (N_11353,N_8015,N_6630);
and U11354 (N_11354,N_7718,N_6961);
nor U11355 (N_11355,N_7948,N_7850);
or U11356 (N_11356,N_6930,N_6566);
and U11357 (N_11357,N_7811,N_6431);
or U11358 (N_11358,N_8883,N_7440);
xor U11359 (N_11359,N_8009,N_8076);
nand U11360 (N_11360,N_6470,N_8654);
and U11361 (N_11361,N_6955,N_7982);
xnor U11362 (N_11362,N_8419,N_8834);
and U11363 (N_11363,N_8699,N_7800);
and U11364 (N_11364,N_8444,N_7893);
nand U11365 (N_11365,N_6957,N_8116);
nor U11366 (N_11366,N_6620,N_7438);
nor U11367 (N_11367,N_6606,N_8091);
or U11368 (N_11368,N_7579,N_6406);
nand U11369 (N_11369,N_6327,N_6388);
or U11370 (N_11370,N_8294,N_8352);
and U11371 (N_11371,N_7160,N_8577);
nand U11372 (N_11372,N_7052,N_7824);
nor U11373 (N_11373,N_6960,N_8701);
nor U11374 (N_11374,N_6697,N_7539);
or U11375 (N_11375,N_7934,N_6605);
xor U11376 (N_11376,N_6308,N_8338);
and U11377 (N_11377,N_8215,N_6474);
and U11378 (N_11378,N_6325,N_6754);
xnor U11379 (N_11379,N_7857,N_8326);
or U11380 (N_11380,N_8436,N_8010);
and U11381 (N_11381,N_8077,N_6225);
nand U11382 (N_11382,N_7950,N_8627);
nor U11383 (N_11383,N_6874,N_6248);
nand U11384 (N_11384,N_8395,N_6976);
nor U11385 (N_11385,N_7289,N_7988);
xor U11386 (N_11386,N_7879,N_6551);
or U11387 (N_11387,N_7533,N_8134);
or U11388 (N_11388,N_8804,N_8982);
xnor U11389 (N_11389,N_7996,N_8765);
nor U11390 (N_11390,N_7206,N_8899);
xnor U11391 (N_11391,N_8469,N_7344);
nand U11392 (N_11392,N_7642,N_7843);
and U11393 (N_11393,N_7684,N_6661);
or U11394 (N_11394,N_8075,N_7772);
or U11395 (N_11395,N_6971,N_8083);
xor U11396 (N_11396,N_7172,N_7124);
nand U11397 (N_11397,N_8454,N_7111);
and U11398 (N_11398,N_7953,N_8017);
nor U11399 (N_11399,N_8055,N_8775);
nand U11400 (N_11400,N_7364,N_6625);
nor U11401 (N_11401,N_7044,N_8780);
nand U11402 (N_11402,N_6837,N_7174);
xnor U11403 (N_11403,N_8551,N_7246);
nand U11404 (N_11404,N_8478,N_8939);
nor U11405 (N_11405,N_7588,N_8102);
or U11406 (N_11406,N_6458,N_6700);
nor U11407 (N_11407,N_6793,N_7793);
and U11408 (N_11408,N_8490,N_7077);
xnor U11409 (N_11409,N_8378,N_8499);
or U11410 (N_11410,N_6779,N_6469);
nor U11411 (N_11411,N_8100,N_7613);
or U11412 (N_11412,N_7621,N_6692);
nor U11413 (N_11413,N_6152,N_7321);
xor U11414 (N_11414,N_7670,N_7956);
or U11415 (N_11415,N_7124,N_6734);
nor U11416 (N_11416,N_7988,N_8964);
nand U11417 (N_11417,N_7978,N_6890);
and U11418 (N_11418,N_6934,N_6423);
nor U11419 (N_11419,N_8306,N_6396);
or U11420 (N_11420,N_8348,N_8026);
nand U11421 (N_11421,N_6558,N_6367);
nor U11422 (N_11422,N_8386,N_7116);
nand U11423 (N_11423,N_6606,N_8044);
xnor U11424 (N_11424,N_7226,N_8484);
xor U11425 (N_11425,N_6562,N_8847);
and U11426 (N_11426,N_7079,N_7445);
xor U11427 (N_11427,N_8275,N_8555);
or U11428 (N_11428,N_6317,N_8725);
or U11429 (N_11429,N_8294,N_8336);
and U11430 (N_11430,N_7233,N_6241);
nand U11431 (N_11431,N_7304,N_8002);
xnor U11432 (N_11432,N_8726,N_6385);
xnor U11433 (N_11433,N_7678,N_6629);
nand U11434 (N_11434,N_8211,N_8099);
xor U11435 (N_11435,N_6003,N_7144);
xnor U11436 (N_11436,N_7432,N_8396);
nor U11437 (N_11437,N_6816,N_7262);
nor U11438 (N_11438,N_7319,N_8918);
nand U11439 (N_11439,N_8118,N_7272);
xnor U11440 (N_11440,N_6127,N_7002);
nand U11441 (N_11441,N_7092,N_6858);
nor U11442 (N_11442,N_8311,N_7882);
nand U11443 (N_11443,N_6750,N_8875);
xnor U11444 (N_11444,N_8321,N_8284);
and U11445 (N_11445,N_7376,N_8604);
and U11446 (N_11446,N_6237,N_8501);
or U11447 (N_11447,N_6545,N_8038);
and U11448 (N_11448,N_7550,N_6633);
and U11449 (N_11449,N_6394,N_7361);
and U11450 (N_11450,N_6838,N_8484);
nor U11451 (N_11451,N_7824,N_8160);
nand U11452 (N_11452,N_7556,N_6079);
nand U11453 (N_11453,N_6764,N_6369);
nand U11454 (N_11454,N_6869,N_8994);
nor U11455 (N_11455,N_6484,N_6234);
nor U11456 (N_11456,N_7330,N_6673);
xor U11457 (N_11457,N_6806,N_7684);
and U11458 (N_11458,N_6273,N_7289);
nand U11459 (N_11459,N_7976,N_7236);
nand U11460 (N_11460,N_6405,N_6959);
and U11461 (N_11461,N_6142,N_8660);
nand U11462 (N_11462,N_7097,N_6826);
or U11463 (N_11463,N_6968,N_6156);
nor U11464 (N_11464,N_6084,N_6669);
nor U11465 (N_11465,N_6141,N_7258);
nand U11466 (N_11466,N_6923,N_8400);
nand U11467 (N_11467,N_6880,N_8542);
xor U11468 (N_11468,N_6421,N_6345);
xnor U11469 (N_11469,N_7026,N_6795);
or U11470 (N_11470,N_8995,N_8408);
or U11471 (N_11471,N_6471,N_6425);
or U11472 (N_11472,N_8819,N_6823);
or U11473 (N_11473,N_7096,N_8518);
and U11474 (N_11474,N_6023,N_8511);
nand U11475 (N_11475,N_8660,N_7191);
or U11476 (N_11476,N_8381,N_8044);
nand U11477 (N_11477,N_8432,N_6801);
and U11478 (N_11478,N_8221,N_8281);
and U11479 (N_11479,N_6128,N_7235);
xor U11480 (N_11480,N_8688,N_8874);
xnor U11481 (N_11481,N_8453,N_6162);
nor U11482 (N_11482,N_7350,N_7563);
or U11483 (N_11483,N_6920,N_6315);
and U11484 (N_11484,N_6535,N_7527);
xor U11485 (N_11485,N_7413,N_7608);
or U11486 (N_11486,N_6611,N_6198);
and U11487 (N_11487,N_8091,N_7432);
nand U11488 (N_11488,N_8026,N_6213);
nand U11489 (N_11489,N_8357,N_6953);
and U11490 (N_11490,N_6196,N_7299);
nor U11491 (N_11491,N_8324,N_7097);
nor U11492 (N_11492,N_6831,N_7968);
and U11493 (N_11493,N_6911,N_8742);
xor U11494 (N_11494,N_8840,N_7097);
and U11495 (N_11495,N_7020,N_8632);
or U11496 (N_11496,N_8217,N_7835);
nand U11497 (N_11497,N_6430,N_6585);
nand U11498 (N_11498,N_6637,N_6251);
and U11499 (N_11499,N_7917,N_8983);
xor U11500 (N_11500,N_6761,N_6373);
nor U11501 (N_11501,N_7762,N_8608);
xnor U11502 (N_11502,N_7107,N_7611);
or U11503 (N_11503,N_6557,N_6179);
nand U11504 (N_11504,N_8715,N_8646);
or U11505 (N_11505,N_6341,N_7284);
or U11506 (N_11506,N_7261,N_6638);
nand U11507 (N_11507,N_7646,N_8043);
nor U11508 (N_11508,N_8726,N_7730);
xor U11509 (N_11509,N_8058,N_7804);
nor U11510 (N_11510,N_8646,N_6729);
xor U11511 (N_11511,N_6246,N_7803);
and U11512 (N_11512,N_8338,N_6107);
or U11513 (N_11513,N_8180,N_6659);
nor U11514 (N_11514,N_7401,N_7722);
xnor U11515 (N_11515,N_7004,N_8493);
or U11516 (N_11516,N_7084,N_7758);
nand U11517 (N_11517,N_8151,N_7329);
and U11518 (N_11518,N_7908,N_7730);
xor U11519 (N_11519,N_8855,N_6368);
xnor U11520 (N_11520,N_8763,N_8275);
nand U11521 (N_11521,N_6940,N_7537);
xnor U11522 (N_11522,N_8581,N_8563);
nand U11523 (N_11523,N_7505,N_8086);
nand U11524 (N_11524,N_8669,N_7951);
and U11525 (N_11525,N_7425,N_7195);
nor U11526 (N_11526,N_7922,N_6792);
and U11527 (N_11527,N_7053,N_6081);
xnor U11528 (N_11528,N_7063,N_7116);
and U11529 (N_11529,N_8175,N_6564);
xnor U11530 (N_11530,N_6199,N_7709);
nand U11531 (N_11531,N_7187,N_6038);
nand U11532 (N_11532,N_6957,N_7033);
nand U11533 (N_11533,N_8038,N_8662);
nand U11534 (N_11534,N_8141,N_7063);
or U11535 (N_11535,N_6969,N_7153);
nand U11536 (N_11536,N_6464,N_6224);
nor U11537 (N_11537,N_6577,N_8857);
nor U11538 (N_11538,N_6769,N_8740);
xnor U11539 (N_11539,N_8487,N_8079);
and U11540 (N_11540,N_7910,N_8896);
and U11541 (N_11541,N_8252,N_6735);
and U11542 (N_11542,N_6933,N_7041);
or U11543 (N_11543,N_6834,N_7926);
or U11544 (N_11544,N_8361,N_8899);
nor U11545 (N_11545,N_6653,N_7862);
xor U11546 (N_11546,N_8195,N_6594);
nor U11547 (N_11547,N_7548,N_6886);
xor U11548 (N_11548,N_8572,N_6170);
xnor U11549 (N_11549,N_8341,N_8333);
nor U11550 (N_11550,N_6669,N_6489);
nor U11551 (N_11551,N_7612,N_8239);
and U11552 (N_11552,N_8327,N_8387);
nand U11553 (N_11553,N_8531,N_6154);
nor U11554 (N_11554,N_6513,N_6022);
xnor U11555 (N_11555,N_6946,N_8882);
nor U11556 (N_11556,N_6065,N_6486);
and U11557 (N_11557,N_8705,N_8454);
and U11558 (N_11558,N_6664,N_8364);
or U11559 (N_11559,N_6579,N_6134);
or U11560 (N_11560,N_8017,N_8114);
nand U11561 (N_11561,N_8929,N_7859);
or U11562 (N_11562,N_7367,N_6769);
and U11563 (N_11563,N_7018,N_7795);
or U11564 (N_11564,N_7518,N_6842);
xnor U11565 (N_11565,N_7304,N_8249);
or U11566 (N_11566,N_7786,N_8221);
nand U11567 (N_11567,N_7322,N_6616);
nand U11568 (N_11568,N_8545,N_6678);
nor U11569 (N_11569,N_8285,N_6675);
and U11570 (N_11570,N_6705,N_7472);
nand U11571 (N_11571,N_8524,N_7928);
xnor U11572 (N_11572,N_8587,N_7113);
and U11573 (N_11573,N_8514,N_6791);
or U11574 (N_11574,N_8975,N_7709);
xnor U11575 (N_11575,N_6607,N_6472);
and U11576 (N_11576,N_7988,N_8218);
and U11577 (N_11577,N_7294,N_6587);
nor U11578 (N_11578,N_8539,N_8543);
and U11579 (N_11579,N_8956,N_6246);
xor U11580 (N_11580,N_7582,N_7140);
xnor U11581 (N_11581,N_7883,N_8683);
nor U11582 (N_11582,N_6676,N_6048);
or U11583 (N_11583,N_6490,N_8795);
nand U11584 (N_11584,N_7843,N_7520);
nand U11585 (N_11585,N_7998,N_7109);
nor U11586 (N_11586,N_8644,N_8472);
and U11587 (N_11587,N_6582,N_8863);
nand U11588 (N_11588,N_6948,N_7761);
xor U11589 (N_11589,N_7961,N_8385);
nand U11590 (N_11590,N_8679,N_7689);
and U11591 (N_11591,N_6620,N_6239);
xnor U11592 (N_11592,N_6263,N_6744);
and U11593 (N_11593,N_6870,N_8226);
xor U11594 (N_11594,N_7909,N_8908);
or U11595 (N_11595,N_8004,N_6831);
nand U11596 (N_11596,N_7603,N_6091);
xor U11597 (N_11597,N_7648,N_8065);
nand U11598 (N_11598,N_7765,N_8503);
or U11599 (N_11599,N_8814,N_8031);
or U11600 (N_11600,N_8213,N_6576);
nor U11601 (N_11601,N_8497,N_7764);
nand U11602 (N_11602,N_7235,N_6379);
nor U11603 (N_11603,N_7991,N_7684);
nand U11604 (N_11604,N_8135,N_7770);
and U11605 (N_11605,N_8274,N_8464);
and U11606 (N_11606,N_6581,N_7988);
nand U11607 (N_11607,N_7350,N_6251);
xnor U11608 (N_11608,N_7388,N_6487);
xnor U11609 (N_11609,N_8791,N_8760);
xnor U11610 (N_11610,N_6052,N_6690);
and U11611 (N_11611,N_8916,N_8871);
and U11612 (N_11612,N_7716,N_7110);
nand U11613 (N_11613,N_7791,N_6399);
or U11614 (N_11614,N_8662,N_7841);
nand U11615 (N_11615,N_8385,N_8514);
and U11616 (N_11616,N_8223,N_6408);
or U11617 (N_11617,N_7862,N_6399);
nand U11618 (N_11618,N_8625,N_7946);
nand U11619 (N_11619,N_8127,N_8292);
or U11620 (N_11620,N_7286,N_8429);
nor U11621 (N_11621,N_7990,N_8727);
nor U11622 (N_11622,N_6137,N_8987);
or U11623 (N_11623,N_6067,N_7891);
nor U11624 (N_11624,N_8698,N_7444);
nand U11625 (N_11625,N_8315,N_8764);
xor U11626 (N_11626,N_7032,N_8380);
nand U11627 (N_11627,N_8370,N_7702);
xnor U11628 (N_11628,N_6653,N_8023);
nor U11629 (N_11629,N_6284,N_8722);
nand U11630 (N_11630,N_8006,N_7156);
and U11631 (N_11631,N_8922,N_7555);
and U11632 (N_11632,N_6027,N_7632);
nor U11633 (N_11633,N_7315,N_6258);
nand U11634 (N_11634,N_8722,N_7110);
nor U11635 (N_11635,N_8771,N_8987);
and U11636 (N_11636,N_7372,N_7090);
or U11637 (N_11637,N_6828,N_7829);
or U11638 (N_11638,N_7557,N_7507);
nor U11639 (N_11639,N_7887,N_6561);
nor U11640 (N_11640,N_7026,N_6661);
and U11641 (N_11641,N_7409,N_8930);
or U11642 (N_11642,N_7694,N_8359);
and U11643 (N_11643,N_6783,N_8648);
xnor U11644 (N_11644,N_7237,N_8332);
nor U11645 (N_11645,N_6080,N_7126);
or U11646 (N_11646,N_7990,N_8271);
nor U11647 (N_11647,N_6077,N_8782);
nand U11648 (N_11648,N_8693,N_6415);
and U11649 (N_11649,N_7916,N_7901);
or U11650 (N_11650,N_8199,N_8540);
xor U11651 (N_11651,N_6118,N_8312);
nor U11652 (N_11652,N_7667,N_6054);
nand U11653 (N_11653,N_6285,N_8993);
or U11654 (N_11654,N_8886,N_6205);
xnor U11655 (N_11655,N_7837,N_7267);
or U11656 (N_11656,N_6522,N_6342);
nor U11657 (N_11657,N_6571,N_8656);
nand U11658 (N_11658,N_8537,N_6819);
or U11659 (N_11659,N_7048,N_6272);
xnor U11660 (N_11660,N_7577,N_7453);
nor U11661 (N_11661,N_7736,N_6582);
or U11662 (N_11662,N_8516,N_7444);
nand U11663 (N_11663,N_6224,N_8517);
nor U11664 (N_11664,N_7973,N_8010);
or U11665 (N_11665,N_7371,N_6113);
and U11666 (N_11666,N_6070,N_8842);
and U11667 (N_11667,N_8124,N_6455);
xor U11668 (N_11668,N_6327,N_6624);
or U11669 (N_11669,N_8844,N_6810);
nand U11670 (N_11670,N_7164,N_7888);
or U11671 (N_11671,N_8481,N_6912);
or U11672 (N_11672,N_7156,N_6631);
and U11673 (N_11673,N_7047,N_8728);
nor U11674 (N_11674,N_8496,N_7134);
xnor U11675 (N_11675,N_7052,N_6099);
nand U11676 (N_11676,N_6288,N_8278);
xnor U11677 (N_11677,N_8238,N_8100);
nand U11678 (N_11678,N_6271,N_6504);
nor U11679 (N_11679,N_6865,N_6554);
or U11680 (N_11680,N_8989,N_6852);
or U11681 (N_11681,N_6036,N_7720);
and U11682 (N_11682,N_8536,N_6124);
xnor U11683 (N_11683,N_7856,N_7160);
or U11684 (N_11684,N_7043,N_7053);
nand U11685 (N_11685,N_7316,N_6339);
and U11686 (N_11686,N_6802,N_8526);
and U11687 (N_11687,N_6650,N_8787);
nand U11688 (N_11688,N_8934,N_7337);
nor U11689 (N_11689,N_8461,N_8339);
or U11690 (N_11690,N_6689,N_8210);
nand U11691 (N_11691,N_8781,N_6528);
nand U11692 (N_11692,N_6388,N_8456);
or U11693 (N_11693,N_7024,N_7717);
xnor U11694 (N_11694,N_6725,N_7398);
nand U11695 (N_11695,N_6555,N_6982);
or U11696 (N_11696,N_6403,N_6540);
and U11697 (N_11697,N_6943,N_6226);
or U11698 (N_11698,N_6845,N_7889);
or U11699 (N_11699,N_6209,N_8844);
nor U11700 (N_11700,N_8516,N_8021);
nand U11701 (N_11701,N_7482,N_6196);
xor U11702 (N_11702,N_8413,N_8102);
nand U11703 (N_11703,N_8651,N_8737);
nand U11704 (N_11704,N_6758,N_6279);
and U11705 (N_11705,N_7083,N_6422);
nand U11706 (N_11706,N_6815,N_6753);
or U11707 (N_11707,N_6375,N_7068);
nor U11708 (N_11708,N_7626,N_8664);
xnor U11709 (N_11709,N_8253,N_8346);
xor U11710 (N_11710,N_8943,N_6908);
and U11711 (N_11711,N_8159,N_8209);
nor U11712 (N_11712,N_6284,N_6111);
nor U11713 (N_11713,N_6636,N_7615);
nor U11714 (N_11714,N_8186,N_8315);
nor U11715 (N_11715,N_6800,N_6083);
and U11716 (N_11716,N_8409,N_6090);
xor U11717 (N_11717,N_8936,N_6405);
or U11718 (N_11718,N_7103,N_7616);
or U11719 (N_11719,N_8306,N_7313);
nor U11720 (N_11720,N_7919,N_8574);
nor U11721 (N_11721,N_6863,N_8242);
and U11722 (N_11722,N_6342,N_7495);
nand U11723 (N_11723,N_8026,N_7899);
nand U11724 (N_11724,N_7850,N_6174);
xnor U11725 (N_11725,N_8739,N_6430);
xor U11726 (N_11726,N_6508,N_6970);
nor U11727 (N_11727,N_6643,N_6691);
nor U11728 (N_11728,N_8650,N_8232);
nor U11729 (N_11729,N_8199,N_7758);
nor U11730 (N_11730,N_6288,N_6422);
and U11731 (N_11731,N_7839,N_8986);
nand U11732 (N_11732,N_8234,N_6600);
and U11733 (N_11733,N_6388,N_8039);
and U11734 (N_11734,N_8992,N_7070);
nand U11735 (N_11735,N_8669,N_6645);
or U11736 (N_11736,N_8263,N_7894);
nand U11737 (N_11737,N_7525,N_8833);
and U11738 (N_11738,N_8578,N_8480);
or U11739 (N_11739,N_8064,N_6793);
xor U11740 (N_11740,N_8322,N_6780);
or U11741 (N_11741,N_6441,N_6876);
or U11742 (N_11742,N_7230,N_7718);
and U11743 (N_11743,N_7939,N_7631);
or U11744 (N_11744,N_8119,N_8111);
xor U11745 (N_11745,N_6778,N_6160);
nand U11746 (N_11746,N_6294,N_7106);
nand U11747 (N_11747,N_6107,N_6094);
nor U11748 (N_11748,N_6279,N_8499);
nor U11749 (N_11749,N_6104,N_6920);
and U11750 (N_11750,N_7076,N_8013);
or U11751 (N_11751,N_6721,N_6847);
nor U11752 (N_11752,N_6865,N_6144);
or U11753 (N_11753,N_7179,N_8816);
nand U11754 (N_11754,N_6290,N_6801);
nor U11755 (N_11755,N_8525,N_7757);
xnor U11756 (N_11756,N_8647,N_8310);
or U11757 (N_11757,N_7512,N_8517);
nor U11758 (N_11758,N_7121,N_7040);
or U11759 (N_11759,N_7380,N_6395);
or U11760 (N_11760,N_6778,N_7433);
or U11761 (N_11761,N_7569,N_6713);
xnor U11762 (N_11762,N_7571,N_8872);
or U11763 (N_11763,N_7610,N_7763);
nor U11764 (N_11764,N_7874,N_8916);
nor U11765 (N_11765,N_8766,N_6932);
nor U11766 (N_11766,N_7446,N_7552);
nand U11767 (N_11767,N_8120,N_8652);
xnor U11768 (N_11768,N_7718,N_8682);
nor U11769 (N_11769,N_6971,N_8879);
or U11770 (N_11770,N_8450,N_7274);
nor U11771 (N_11771,N_8722,N_8701);
nand U11772 (N_11772,N_8047,N_8718);
nor U11773 (N_11773,N_6131,N_7315);
or U11774 (N_11774,N_8466,N_6732);
nand U11775 (N_11775,N_6249,N_8490);
nor U11776 (N_11776,N_6073,N_7409);
or U11777 (N_11777,N_7826,N_7500);
and U11778 (N_11778,N_7439,N_7726);
nand U11779 (N_11779,N_7539,N_6239);
nor U11780 (N_11780,N_7050,N_6186);
and U11781 (N_11781,N_7567,N_8031);
or U11782 (N_11782,N_8095,N_6958);
or U11783 (N_11783,N_7957,N_6812);
and U11784 (N_11784,N_6727,N_6495);
and U11785 (N_11785,N_6303,N_7634);
nor U11786 (N_11786,N_7087,N_7203);
xor U11787 (N_11787,N_7004,N_7891);
and U11788 (N_11788,N_8294,N_7626);
or U11789 (N_11789,N_8728,N_8943);
nor U11790 (N_11790,N_6963,N_7722);
nand U11791 (N_11791,N_6051,N_6551);
xnor U11792 (N_11792,N_7299,N_7684);
nand U11793 (N_11793,N_6888,N_8789);
nand U11794 (N_11794,N_8977,N_6326);
xnor U11795 (N_11795,N_6217,N_7220);
and U11796 (N_11796,N_7619,N_7397);
and U11797 (N_11797,N_8390,N_8987);
xnor U11798 (N_11798,N_6984,N_8977);
nand U11799 (N_11799,N_8798,N_6196);
nor U11800 (N_11800,N_6190,N_6025);
nand U11801 (N_11801,N_8594,N_8778);
xnor U11802 (N_11802,N_8545,N_6240);
or U11803 (N_11803,N_7704,N_6080);
or U11804 (N_11804,N_8619,N_6217);
nand U11805 (N_11805,N_6750,N_8396);
xor U11806 (N_11806,N_7297,N_6135);
and U11807 (N_11807,N_6223,N_8175);
nand U11808 (N_11808,N_7611,N_8631);
nand U11809 (N_11809,N_8405,N_6734);
xor U11810 (N_11810,N_8505,N_7993);
and U11811 (N_11811,N_8699,N_7015);
and U11812 (N_11812,N_6239,N_7213);
or U11813 (N_11813,N_8136,N_8942);
and U11814 (N_11814,N_6868,N_6235);
xnor U11815 (N_11815,N_8860,N_8666);
nor U11816 (N_11816,N_7337,N_7721);
or U11817 (N_11817,N_8218,N_8575);
and U11818 (N_11818,N_8821,N_7747);
and U11819 (N_11819,N_6641,N_7961);
or U11820 (N_11820,N_8872,N_6635);
and U11821 (N_11821,N_8941,N_7290);
or U11822 (N_11822,N_8410,N_7452);
and U11823 (N_11823,N_7122,N_7276);
xnor U11824 (N_11824,N_8730,N_7304);
and U11825 (N_11825,N_6696,N_6258);
or U11826 (N_11826,N_8589,N_6534);
or U11827 (N_11827,N_6909,N_6382);
and U11828 (N_11828,N_8316,N_8656);
and U11829 (N_11829,N_7651,N_7603);
xnor U11830 (N_11830,N_7629,N_8652);
or U11831 (N_11831,N_6492,N_7433);
and U11832 (N_11832,N_7235,N_7629);
nand U11833 (N_11833,N_8873,N_7417);
xor U11834 (N_11834,N_8608,N_8113);
nand U11835 (N_11835,N_7059,N_6036);
xor U11836 (N_11836,N_6644,N_6540);
xnor U11837 (N_11837,N_8718,N_8587);
nand U11838 (N_11838,N_7644,N_8307);
nand U11839 (N_11839,N_6797,N_6601);
nor U11840 (N_11840,N_8378,N_7162);
nor U11841 (N_11841,N_6444,N_6928);
or U11842 (N_11842,N_8736,N_8338);
or U11843 (N_11843,N_8274,N_6052);
nand U11844 (N_11844,N_7509,N_6317);
and U11845 (N_11845,N_6967,N_6315);
and U11846 (N_11846,N_8314,N_6255);
or U11847 (N_11847,N_8320,N_7845);
nand U11848 (N_11848,N_6913,N_8599);
or U11849 (N_11849,N_8735,N_7704);
and U11850 (N_11850,N_6160,N_7311);
nor U11851 (N_11851,N_7977,N_6566);
nand U11852 (N_11852,N_6822,N_8172);
or U11853 (N_11853,N_6780,N_8432);
nor U11854 (N_11854,N_6088,N_7931);
xor U11855 (N_11855,N_6444,N_7173);
or U11856 (N_11856,N_7752,N_6172);
or U11857 (N_11857,N_7475,N_8656);
nand U11858 (N_11858,N_6912,N_8877);
and U11859 (N_11859,N_6567,N_6059);
and U11860 (N_11860,N_8191,N_7093);
nand U11861 (N_11861,N_8650,N_6826);
xor U11862 (N_11862,N_7457,N_8966);
and U11863 (N_11863,N_8568,N_8877);
xor U11864 (N_11864,N_7437,N_7581);
or U11865 (N_11865,N_7232,N_8295);
nand U11866 (N_11866,N_6754,N_6104);
nand U11867 (N_11867,N_8092,N_7289);
and U11868 (N_11868,N_8997,N_7862);
nand U11869 (N_11869,N_7949,N_6284);
nor U11870 (N_11870,N_8732,N_6698);
nand U11871 (N_11871,N_7853,N_8657);
xnor U11872 (N_11872,N_6413,N_7784);
nor U11873 (N_11873,N_8827,N_6741);
nor U11874 (N_11874,N_6764,N_7208);
nor U11875 (N_11875,N_6545,N_8613);
xor U11876 (N_11876,N_6565,N_7982);
nand U11877 (N_11877,N_7516,N_7041);
nand U11878 (N_11878,N_7373,N_6614);
nand U11879 (N_11879,N_7939,N_7512);
or U11880 (N_11880,N_6928,N_7481);
xnor U11881 (N_11881,N_7233,N_6366);
nor U11882 (N_11882,N_7018,N_7986);
xnor U11883 (N_11883,N_7564,N_6735);
or U11884 (N_11884,N_6062,N_6464);
nand U11885 (N_11885,N_7710,N_8923);
nor U11886 (N_11886,N_6931,N_8555);
nand U11887 (N_11887,N_7989,N_6703);
and U11888 (N_11888,N_7238,N_6615);
xor U11889 (N_11889,N_8452,N_6857);
nor U11890 (N_11890,N_6441,N_8991);
nor U11891 (N_11891,N_7795,N_6979);
or U11892 (N_11892,N_6271,N_8435);
nand U11893 (N_11893,N_6401,N_7536);
or U11894 (N_11894,N_8670,N_7440);
nand U11895 (N_11895,N_8644,N_7031);
nor U11896 (N_11896,N_7769,N_8897);
nand U11897 (N_11897,N_7288,N_6478);
xnor U11898 (N_11898,N_8419,N_8518);
nor U11899 (N_11899,N_8703,N_6589);
nor U11900 (N_11900,N_6870,N_7220);
nor U11901 (N_11901,N_7433,N_6609);
or U11902 (N_11902,N_7521,N_6644);
nand U11903 (N_11903,N_7508,N_8668);
and U11904 (N_11904,N_7955,N_6092);
and U11905 (N_11905,N_8527,N_7473);
xnor U11906 (N_11906,N_7090,N_6300);
or U11907 (N_11907,N_8898,N_7111);
and U11908 (N_11908,N_6647,N_7678);
nor U11909 (N_11909,N_8620,N_8455);
nand U11910 (N_11910,N_6879,N_8873);
and U11911 (N_11911,N_6860,N_7855);
xnor U11912 (N_11912,N_6930,N_8714);
nand U11913 (N_11913,N_6174,N_7764);
nand U11914 (N_11914,N_8017,N_6085);
nand U11915 (N_11915,N_7390,N_8528);
and U11916 (N_11916,N_7970,N_7926);
nor U11917 (N_11917,N_6129,N_8024);
xnor U11918 (N_11918,N_7884,N_7989);
or U11919 (N_11919,N_7905,N_7107);
nand U11920 (N_11920,N_7043,N_8853);
nor U11921 (N_11921,N_8033,N_8784);
and U11922 (N_11922,N_6447,N_6935);
nand U11923 (N_11923,N_7182,N_8313);
xnor U11924 (N_11924,N_7714,N_8864);
nand U11925 (N_11925,N_6010,N_7830);
xnor U11926 (N_11926,N_7805,N_7354);
or U11927 (N_11927,N_8237,N_6211);
xor U11928 (N_11928,N_8416,N_8182);
and U11929 (N_11929,N_7723,N_8681);
nand U11930 (N_11930,N_8474,N_6505);
nor U11931 (N_11931,N_8830,N_6099);
nor U11932 (N_11932,N_7607,N_6930);
nand U11933 (N_11933,N_6779,N_6065);
nand U11934 (N_11934,N_7815,N_7471);
nand U11935 (N_11935,N_6764,N_8442);
nand U11936 (N_11936,N_8151,N_8341);
nand U11937 (N_11937,N_8865,N_6354);
and U11938 (N_11938,N_7439,N_6618);
or U11939 (N_11939,N_6520,N_6497);
xnor U11940 (N_11940,N_8227,N_7137);
and U11941 (N_11941,N_8296,N_7571);
nor U11942 (N_11942,N_7915,N_8325);
or U11943 (N_11943,N_7846,N_6253);
xnor U11944 (N_11944,N_6305,N_6361);
nand U11945 (N_11945,N_6449,N_6528);
nor U11946 (N_11946,N_6175,N_6916);
and U11947 (N_11947,N_7149,N_8386);
xnor U11948 (N_11948,N_7158,N_7501);
nand U11949 (N_11949,N_8507,N_8115);
or U11950 (N_11950,N_7357,N_6559);
and U11951 (N_11951,N_6171,N_7112);
xor U11952 (N_11952,N_8600,N_8857);
and U11953 (N_11953,N_7949,N_6324);
nor U11954 (N_11954,N_7756,N_8042);
and U11955 (N_11955,N_6269,N_7195);
nor U11956 (N_11956,N_7039,N_8402);
nand U11957 (N_11957,N_8983,N_7332);
nand U11958 (N_11958,N_7019,N_8850);
xnor U11959 (N_11959,N_6130,N_7653);
or U11960 (N_11960,N_8129,N_7772);
or U11961 (N_11961,N_6133,N_6250);
nor U11962 (N_11962,N_7865,N_6291);
xor U11963 (N_11963,N_6782,N_6959);
xor U11964 (N_11964,N_7934,N_8460);
xnor U11965 (N_11965,N_7172,N_8398);
or U11966 (N_11966,N_6966,N_6213);
nand U11967 (N_11967,N_8536,N_6556);
nand U11968 (N_11968,N_6828,N_8438);
or U11969 (N_11969,N_6234,N_6867);
xnor U11970 (N_11970,N_6854,N_6492);
xor U11971 (N_11971,N_7392,N_6163);
nor U11972 (N_11972,N_8718,N_8105);
nor U11973 (N_11973,N_6515,N_8699);
or U11974 (N_11974,N_7986,N_6783);
or U11975 (N_11975,N_6898,N_8810);
or U11976 (N_11976,N_6192,N_6813);
xnor U11977 (N_11977,N_6923,N_8188);
or U11978 (N_11978,N_7545,N_6868);
nor U11979 (N_11979,N_7933,N_7891);
xor U11980 (N_11980,N_7139,N_8175);
xor U11981 (N_11981,N_7345,N_6435);
and U11982 (N_11982,N_7111,N_6772);
xnor U11983 (N_11983,N_8520,N_6622);
and U11984 (N_11984,N_8389,N_8002);
nor U11985 (N_11985,N_7022,N_6531);
nand U11986 (N_11986,N_7905,N_8641);
and U11987 (N_11987,N_6009,N_8620);
and U11988 (N_11988,N_6128,N_8598);
nor U11989 (N_11989,N_7692,N_7680);
or U11990 (N_11990,N_7422,N_8202);
xor U11991 (N_11991,N_7185,N_6230);
xnor U11992 (N_11992,N_8797,N_7878);
xor U11993 (N_11993,N_8943,N_8555);
and U11994 (N_11994,N_6967,N_8240);
and U11995 (N_11995,N_6602,N_7068);
nand U11996 (N_11996,N_8232,N_8206);
and U11997 (N_11997,N_7953,N_8537);
and U11998 (N_11998,N_7163,N_6954);
nor U11999 (N_11999,N_7640,N_8093);
xnor U12000 (N_12000,N_11075,N_10013);
nor U12001 (N_12001,N_11101,N_11529);
nand U12002 (N_12002,N_11449,N_9887);
xnor U12003 (N_12003,N_10372,N_9730);
xor U12004 (N_12004,N_10364,N_9572);
and U12005 (N_12005,N_9033,N_9988);
or U12006 (N_12006,N_10869,N_9619);
xnor U12007 (N_12007,N_11240,N_11431);
and U12008 (N_12008,N_10440,N_10874);
and U12009 (N_12009,N_11480,N_9255);
and U12010 (N_12010,N_10395,N_9426);
nor U12011 (N_12011,N_9154,N_11589);
nor U12012 (N_12012,N_10268,N_10156);
xnor U12013 (N_12013,N_11619,N_11693);
xnor U12014 (N_12014,N_11256,N_10975);
and U12015 (N_12015,N_10474,N_10996);
or U12016 (N_12016,N_10266,N_9833);
and U12017 (N_12017,N_11024,N_11754);
and U12018 (N_12018,N_11765,N_10202);
or U12019 (N_12019,N_10931,N_11466);
nor U12020 (N_12020,N_10680,N_10167);
nand U12021 (N_12021,N_9280,N_9910);
xor U12022 (N_12022,N_10154,N_11519);
or U12023 (N_12023,N_10531,N_10522);
and U12024 (N_12024,N_9179,N_10646);
nand U12025 (N_12025,N_11530,N_10872);
xor U12026 (N_12026,N_10622,N_9026);
xnor U12027 (N_12027,N_9024,N_11143);
nand U12028 (N_12028,N_9173,N_10318);
nor U12029 (N_12029,N_9145,N_9886);
xnor U12030 (N_12030,N_11369,N_9251);
or U12031 (N_12031,N_9906,N_11363);
and U12032 (N_12032,N_9620,N_11925);
or U12033 (N_12033,N_10660,N_9881);
or U12034 (N_12034,N_11081,N_9905);
nor U12035 (N_12035,N_11474,N_9562);
and U12036 (N_12036,N_11883,N_9659);
nand U12037 (N_12037,N_11722,N_10687);
and U12038 (N_12038,N_9935,N_10348);
nand U12039 (N_12039,N_9837,N_9820);
or U12040 (N_12040,N_11669,N_11406);
or U12041 (N_12041,N_11318,N_9359);
xor U12042 (N_12042,N_9706,N_11473);
and U12043 (N_12043,N_11761,N_9057);
xor U12044 (N_12044,N_11877,N_9556);
xor U12045 (N_12045,N_9438,N_10175);
xor U12046 (N_12046,N_11346,N_9188);
nor U12047 (N_12047,N_11884,N_11961);
nor U12048 (N_12048,N_9648,N_11926);
nor U12049 (N_12049,N_11935,N_10773);
xnor U12050 (N_12050,N_9711,N_11167);
xnor U12051 (N_12051,N_9960,N_11223);
nand U12052 (N_12052,N_9455,N_10123);
nand U12053 (N_12053,N_10292,N_10473);
xor U12054 (N_12054,N_11061,N_10153);
nand U12055 (N_12055,N_10124,N_10562);
nor U12056 (N_12056,N_9044,N_10957);
or U12057 (N_12057,N_9680,N_10170);
nand U12058 (N_12058,N_11315,N_9846);
nor U12059 (N_12059,N_11510,N_10674);
nor U12060 (N_12060,N_11834,N_9600);
nor U12061 (N_12061,N_11556,N_9403);
nor U12062 (N_12062,N_11399,N_10418);
and U12063 (N_12063,N_9553,N_9640);
nand U12064 (N_12064,N_11854,N_10045);
xor U12065 (N_12065,N_9337,N_10788);
nor U12066 (N_12066,N_10520,N_10621);
nand U12067 (N_12067,N_11823,N_10691);
and U12068 (N_12068,N_9127,N_9571);
nor U12069 (N_12069,N_11413,N_10523);
nand U12070 (N_12070,N_10637,N_9235);
nand U12071 (N_12071,N_10300,N_9368);
and U12072 (N_12072,N_10050,N_10443);
or U12073 (N_12073,N_11420,N_9664);
xnor U12074 (N_12074,N_10686,N_9317);
and U12075 (N_12075,N_9966,N_10091);
xnor U12076 (N_12076,N_9329,N_10306);
or U12077 (N_12077,N_11724,N_11940);
or U12078 (N_12078,N_9654,N_9313);
nand U12079 (N_12079,N_9198,N_10378);
nand U12080 (N_12080,N_11165,N_9926);
nand U12081 (N_12081,N_10947,N_9101);
and U12082 (N_12082,N_10070,N_10939);
nand U12083 (N_12083,N_10628,N_10067);
xnor U12084 (N_12084,N_10386,N_9172);
nor U12085 (N_12085,N_10583,N_9183);
or U12086 (N_12086,N_11440,N_10461);
and U12087 (N_12087,N_10235,N_11389);
nor U12088 (N_12088,N_9615,N_9987);
or U12089 (N_12089,N_10671,N_11763);
or U12090 (N_12090,N_11591,N_11342);
nor U12091 (N_12091,N_10608,N_10712);
or U12092 (N_12092,N_10126,N_11164);
or U12093 (N_12093,N_10827,N_11978);
nor U12094 (N_12094,N_10875,N_11042);
nor U12095 (N_12095,N_10594,N_10243);
xnor U12096 (N_12096,N_9842,N_9717);
nor U12097 (N_12097,N_9272,N_11584);
xnor U12098 (N_12098,N_9034,N_10880);
and U12099 (N_12099,N_9611,N_9892);
xnor U12100 (N_12100,N_10639,N_10427);
or U12101 (N_12101,N_10792,N_10643);
nor U12102 (N_12102,N_10758,N_10718);
or U12103 (N_12103,N_10128,N_11445);
and U12104 (N_12104,N_11816,N_9772);
and U12105 (N_12105,N_11371,N_10388);
nor U12106 (N_12106,N_9757,N_10766);
and U12107 (N_12107,N_9082,N_10441);
and U12108 (N_12108,N_10840,N_11567);
nand U12109 (N_12109,N_9440,N_10759);
and U12110 (N_12110,N_11219,N_10798);
nand U12111 (N_12111,N_9570,N_9192);
and U12112 (N_12112,N_11997,N_10977);
nor U12113 (N_12113,N_10730,N_9027);
or U12114 (N_12114,N_10181,N_11234);
xnor U12115 (N_12115,N_9746,N_11019);
or U12116 (N_12116,N_10737,N_11860);
nor U12117 (N_12117,N_11666,N_11962);
and U12118 (N_12118,N_9267,N_9817);
nand U12119 (N_12119,N_10648,N_11411);
and U12120 (N_12120,N_10519,N_9702);
nor U12121 (N_12121,N_11870,N_9003);
and U12122 (N_12122,N_10214,N_9370);
nand U12123 (N_12123,N_10460,N_11683);
and U12124 (N_12124,N_9448,N_10141);
xor U12125 (N_12125,N_10896,N_10631);
or U12126 (N_12126,N_10336,N_11946);
nor U12127 (N_12127,N_9819,N_9930);
nand U12128 (N_12128,N_9918,N_9104);
and U12129 (N_12129,N_9340,N_9124);
nor U12130 (N_12130,N_9625,N_9231);
xnor U12131 (N_12131,N_10756,N_9610);
and U12132 (N_12132,N_11437,N_10638);
or U12133 (N_12133,N_9551,N_9719);
xor U12134 (N_12134,N_9561,N_11719);
nand U12135 (N_12135,N_9509,N_10787);
nand U12136 (N_12136,N_11829,N_10407);
xor U12137 (N_12137,N_10993,N_10494);
nand U12138 (N_12138,N_10165,N_11715);
nor U12139 (N_12139,N_9009,N_11840);
nor U12140 (N_12140,N_11203,N_10158);
and U12141 (N_12141,N_9445,N_9739);
or U12142 (N_12142,N_9281,N_11911);
nor U12143 (N_12143,N_11541,N_9090);
nand U12144 (N_12144,N_9681,N_11907);
or U12145 (N_12145,N_9979,N_10470);
nor U12146 (N_12146,N_9047,N_10271);
nand U12147 (N_12147,N_9688,N_9691);
and U12148 (N_12148,N_11792,N_10915);
or U12149 (N_12149,N_10887,N_9185);
nor U12150 (N_12150,N_10376,N_11456);
nand U12151 (N_12151,N_9635,N_11295);
nor U12152 (N_12152,N_10291,N_9547);
and U12153 (N_12153,N_10366,N_9229);
nand U12154 (N_12154,N_11932,N_10248);
nand U12155 (N_12155,N_9683,N_9297);
xor U12156 (N_12156,N_10065,N_9582);
nor U12157 (N_12157,N_11309,N_9588);
or U12158 (N_12158,N_10451,N_10424);
nor U12159 (N_12159,N_10961,N_9676);
and U12160 (N_12160,N_10920,N_9092);
xnor U12161 (N_12161,N_9394,N_9937);
xor U12162 (N_12162,N_10286,N_10908);
or U12163 (N_12163,N_9517,N_10510);
nor U12164 (N_12164,N_9642,N_9663);
or U12165 (N_12165,N_11964,N_11299);
xor U12166 (N_12166,N_9971,N_9279);
nand U12167 (N_12167,N_11463,N_9078);
xnor U12168 (N_12168,N_11634,N_9226);
nand U12169 (N_12169,N_10491,N_11447);
or U12170 (N_12170,N_10564,N_9375);
and U12171 (N_12171,N_11646,N_11422);
or U12172 (N_12172,N_9028,N_11172);
or U12173 (N_12173,N_9170,N_9500);
or U12174 (N_12174,N_11286,N_9039);
and U12175 (N_12175,N_9481,N_9446);
nor U12176 (N_12176,N_10782,N_9234);
and U12177 (N_12177,N_10959,N_11557);
xnor U12178 (N_12178,N_10179,N_11728);
nand U12179 (N_12179,N_9331,N_9768);
nand U12180 (N_12180,N_9669,N_10351);
and U12181 (N_12181,N_9404,N_11742);
nand U12182 (N_12182,N_11068,N_11138);
nor U12183 (N_12183,N_9502,N_11535);
and U12184 (N_12184,N_9737,N_10813);
nor U12185 (N_12185,N_9384,N_11434);
nand U12186 (N_12186,N_10554,N_11455);
or U12187 (N_12187,N_9933,N_9818);
nor U12188 (N_12188,N_9766,N_10437);
and U12189 (N_12189,N_10682,N_9849);
xor U12190 (N_12190,N_9984,N_10408);
nor U12191 (N_12191,N_10998,N_10539);
nor U12192 (N_12192,N_9697,N_9285);
nand U12193 (N_12193,N_11284,N_9113);
nor U12194 (N_12194,N_11914,N_9564);
and U12195 (N_12195,N_10725,N_10727);
xnor U12196 (N_12196,N_9965,N_10585);
nand U12197 (N_12197,N_10889,N_9335);
or U12198 (N_12198,N_9275,N_11822);
or U12199 (N_12199,N_10826,N_10810);
xor U12200 (N_12200,N_9157,N_10568);
and U12201 (N_12201,N_11603,N_9042);
or U12202 (N_12202,N_11890,N_10464);
nand U12203 (N_12203,N_10349,N_10755);
and U12204 (N_12204,N_11993,N_11242);
and U12205 (N_12205,N_10471,N_10354);
nand U12206 (N_12206,N_11468,N_10650);
xnor U12207 (N_12207,N_10342,N_9653);
or U12208 (N_12208,N_9148,N_9828);
nand U12209 (N_12209,N_10118,N_9233);
nor U12210 (N_12210,N_10774,N_10681);
and U12211 (N_12211,N_9529,N_9967);
and U12212 (N_12212,N_11528,N_9146);
or U12213 (N_12213,N_10652,N_11737);
and U12214 (N_12214,N_10350,N_9004);
xnor U12215 (N_12215,N_10086,N_11968);
or U12216 (N_12216,N_9815,N_10930);
and U12217 (N_12217,N_11245,N_11703);
nor U12218 (N_12218,N_11384,N_10733);
nand U12219 (N_12219,N_9838,N_10060);
and U12220 (N_12220,N_9542,N_10016);
and U12221 (N_12221,N_10757,N_11858);
xor U12222 (N_12222,N_10741,N_10558);
xor U12223 (N_12223,N_10341,N_10463);
nor U12224 (N_12224,N_11382,N_9451);
xor U12225 (N_12225,N_11502,N_11410);
nor U12226 (N_12226,N_10343,N_10188);
xor U12227 (N_12227,N_11671,N_9465);
or U12228 (N_12228,N_11806,N_9834);
nor U12229 (N_12229,N_11059,N_10784);
and U12230 (N_12230,N_9388,N_11210);
xor U12231 (N_12231,N_11253,N_10180);
xnor U12232 (N_12232,N_9323,N_11654);
nor U12233 (N_12233,N_9661,N_10593);
or U12234 (N_12234,N_10617,N_9633);
nor U12235 (N_12235,N_10358,N_9084);
xor U12236 (N_12236,N_11488,N_10056);
xnor U12237 (N_12237,N_9969,N_9406);
nor U12238 (N_12238,N_9922,N_9431);
nand U12239 (N_12239,N_10498,N_11327);
nor U12240 (N_12240,N_10340,N_11921);
xor U12241 (N_12241,N_11514,N_11049);
and U12242 (N_12242,N_11695,N_10532);
xnor U12243 (N_12243,N_10824,N_10096);
and U12244 (N_12244,N_11435,N_11667);
xor U12245 (N_12245,N_9373,N_9634);
nand U12246 (N_12246,N_10685,N_9512);
nand U12247 (N_12247,N_11425,N_9576);
xor U12248 (N_12248,N_10406,N_10397);
or U12249 (N_12249,N_11385,N_9774);
or U12250 (N_12250,N_9258,N_9327);
nand U12251 (N_12251,N_11617,N_11423);
nor U12252 (N_12252,N_10574,N_9803);
and U12253 (N_12253,N_11265,N_9025);
nand U12254 (N_12254,N_11720,N_9133);
nand U12255 (N_12255,N_10224,N_11361);
or U12256 (N_12256,N_9310,N_9708);
or U12257 (N_12257,N_11637,N_10347);
nand U12258 (N_12258,N_11982,N_11891);
nor U12259 (N_12259,N_9497,N_10048);
and U12260 (N_12260,N_9573,N_11032);
nor U12261 (N_12261,N_10428,N_9098);
xor U12262 (N_12262,N_9333,N_10855);
nor U12263 (N_12263,N_9686,N_11733);
or U12264 (N_12264,N_11461,N_10722);
or U12265 (N_12265,N_9868,N_11321);
xnor U12266 (N_12266,N_10137,N_11071);
nor U12267 (N_12267,N_11475,N_10111);
xor U12268 (N_12268,N_10719,N_9908);
nor U12269 (N_12269,N_11118,N_11937);
xnor U12270 (N_12270,N_9351,N_10864);
nor U12271 (N_12271,N_11663,N_10657);
nor U12272 (N_12272,N_9298,N_9941);
nor U12273 (N_12273,N_11756,N_11041);
and U12274 (N_12274,N_10616,N_10285);
nor U12275 (N_12275,N_11459,N_11696);
nor U12276 (N_12276,N_9832,N_10990);
nor U12277 (N_12277,N_10579,N_11835);
xnor U12278 (N_12278,N_11758,N_10983);
xnor U12279 (N_12279,N_10053,N_10216);
or U12280 (N_12280,N_9189,N_10177);
and U12281 (N_12281,N_11493,N_9952);
xnor U12282 (N_12282,N_11659,N_10288);
nand U12283 (N_12283,N_9475,N_9767);
or U12284 (N_12284,N_9736,N_11582);
xnor U12285 (N_12285,N_11119,N_10634);
nand U12286 (N_12286,N_11272,N_9603);
or U12287 (N_12287,N_9350,N_9424);
xor U12288 (N_12288,N_10548,N_10866);
nand U12289 (N_12289,N_9609,N_10120);
nand U12290 (N_12290,N_10515,N_10851);
nor U12291 (N_12291,N_11105,N_11904);
or U12292 (N_12292,N_10190,N_9714);
nand U12293 (N_12293,N_10417,N_11392);
nor U12294 (N_12294,N_9592,N_9346);
or U12295 (N_12295,N_9002,N_10570);
xnor U12296 (N_12296,N_10995,N_10117);
or U12297 (N_12297,N_10183,N_9811);
nand U12298 (N_12298,N_11853,N_11200);
or U12299 (N_12299,N_10466,N_11824);
nor U12300 (N_12300,N_10469,N_9548);
or U12301 (N_12301,N_11832,N_11970);
nand U12302 (N_12302,N_10449,N_11512);
or U12303 (N_12303,N_11375,N_10768);
or U12304 (N_12304,N_10385,N_10231);
xor U12305 (N_12305,N_9490,N_11175);
xor U12306 (N_12306,N_9765,N_9468);
nand U12307 (N_12307,N_10400,N_11707);
nand U12308 (N_12308,N_9690,N_11527);
nor U12309 (N_12309,N_11776,N_11882);
nand U12310 (N_12310,N_11114,N_11624);
xor U12311 (N_12311,N_10328,N_11625);
and U12312 (N_12312,N_11708,N_11706);
and U12313 (N_12313,N_9347,N_10485);
nand U12314 (N_12314,N_11430,N_10009);
xor U12315 (N_12315,N_10610,N_10832);
nor U12316 (N_12316,N_10816,N_10736);
and U12317 (N_12317,N_9797,N_10390);
and U12318 (N_12318,N_9479,N_10949);
nor U12319 (N_12319,N_10237,N_9223);
nor U12320 (N_12320,N_11034,N_9397);
or U12321 (N_12321,N_11380,N_11780);
nand U12322 (N_12322,N_9062,N_11319);
nand U12323 (N_12323,N_11745,N_9749);
nor U12324 (N_12324,N_9513,N_10511);
and U12325 (N_12325,N_9056,N_10796);
xnor U12326 (N_12326,N_10185,N_9802);
xor U12327 (N_12327,N_9063,N_11391);
nand U12328 (N_12328,N_11573,N_9020);
xnor U12329 (N_12329,N_9201,N_10015);
and U12330 (N_12330,N_9032,N_10546);
and U12331 (N_12331,N_9117,N_9771);
nand U12332 (N_12332,N_11665,N_9421);
or U12333 (N_12333,N_9726,N_11559);
or U12334 (N_12334,N_9873,N_9094);
nor U12335 (N_12335,N_9217,N_10109);
nand U12336 (N_12336,N_11918,N_11827);
and U12337 (N_12337,N_9147,N_11866);
nand U12338 (N_12338,N_10201,N_9067);
xnor U12339 (N_12339,N_9972,N_10134);
or U12340 (N_12340,N_9443,N_11629);
xor U12341 (N_12341,N_9862,N_9439);
xnor U12342 (N_12342,N_10979,N_9636);
xnor U12343 (N_12343,N_11097,N_11439);
or U12344 (N_12344,N_11896,N_9704);
nand U12345 (N_12345,N_10909,N_11846);
and U12346 (N_12346,N_11607,N_11536);
nor U12347 (N_12347,N_9083,N_11862);
and U12348 (N_12348,N_11815,N_9364);
nor U12349 (N_12349,N_11644,N_11465);
and U12350 (N_12350,N_10873,N_10913);
nand U12351 (N_12351,N_9460,N_11838);
and U12352 (N_12352,N_10173,N_9525);
nand U12353 (N_12353,N_9787,N_9806);
xnor U12354 (N_12354,N_11208,N_10371);
xnor U12355 (N_12355,N_10448,N_10678);
xor U12356 (N_12356,N_10778,N_9385);
and U12357 (N_12357,N_10061,N_11509);
nand U12358 (N_12358,N_9283,N_9429);
nand U12359 (N_12359,N_9103,N_11741);
xnor U12360 (N_12360,N_9072,N_9108);
and U12361 (N_12361,N_11429,N_11524);
or U12362 (N_12362,N_10104,N_9301);
or U12363 (N_12363,N_10458,N_10812);
xnor U12364 (N_12364,N_11955,N_10377);
or U12365 (N_12365,N_10982,N_11558);
nor U12366 (N_12366,N_10204,N_10694);
nand U12367 (N_12367,N_9510,N_9111);
nor U12368 (N_12368,N_9679,N_11367);
nand U12369 (N_12369,N_11421,N_9955);
and U12370 (N_12370,N_9864,N_9228);
nand U12371 (N_12371,N_9998,N_11161);
nand U12372 (N_12372,N_9891,N_11148);
or U12373 (N_12373,N_10063,N_10475);
nor U12374 (N_12374,N_10601,N_11368);
nand U12375 (N_12375,N_10431,N_9626);
nor U12376 (N_12376,N_9695,N_10541);
nand U12377 (N_12377,N_11004,N_10801);
or U12378 (N_12378,N_11350,N_10745);
xor U12379 (N_12379,N_10442,N_11923);
xor U12380 (N_12380,N_9874,N_9639);
nand U12381 (N_12381,N_11942,N_9422);
xor U12382 (N_12382,N_9357,N_9597);
nor U12383 (N_12383,N_10025,N_10199);
nor U12384 (N_12384,N_9902,N_10215);
nor U12385 (N_12385,N_9934,N_11296);
nand U12386 (N_12386,N_11581,N_9248);
or U12387 (N_12387,N_10409,N_10355);
or U12388 (N_12388,N_10743,N_11688);
nor U12389 (N_12389,N_10313,N_11267);
nand U12390 (N_12390,N_11176,N_10693);
xor U12391 (N_12391,N_9349,N_10273);
and U12392 (N_12392,N_10367,N_11215);
xnor U12393 (N_12393,N_11405,N_10289);
nand U12394 (N_12394,N_11147,N_11195);
and U12395 (N_12395,N_11444,N_10043);
xor U12396 (N_12396,N_11910,N_9013);
xnor U12397 (N_12397,N_9796,N_10375);
nand U12398 (N_12398,N_11781,N_9011);
or U12399 (N_12399,N_9921,N_10572);
nand U12400 (N_12400,N_9110,N_10919);
and U12401 (N_12401,N_9486,N_9053);
or U12402 (N_12402,N_11912,N_9474);
nand U12403 (N_12403,N_9543,N_11320);
nor U12404 (N_12404,N_11228,N_9861);
or U12405 (N_12405,N_9376,N_11214);
nand U12406 (N_12406,N_9036,N_11712);
and U12407 (N_12407,N_11141,N_10706);
and U12408 (N_12408,N_9177,N_10234);
and U12409 (N_12409,N_10699,N_10857);
nand U12410 (N_12410,N_11098,N_11479);
nand U12411 (N_12411,N_11575,N_9425);
nor U12412 (N_12412,N_9016,N_10595);
xnor U12413 (N_12413,N_9140,N_11915);
nand U12414 (N_12414,N_9214,N_9135);
xnor U12415 (N_12415,N_10482,N_9069);
or U12416 (N_12416,N_11000,N_10769);
nor U12417 (N_12417,N_10151,N_9498);
or U12418 (N_12418,N_10174,N_10459);
nand U12419 (N_12419,N_9759,N_11356);
xnor U12420 (N_12420,N_11158,N_11606);
and U12421 (N_12421,N_10781,N_11458);
or U12422 (N_12422,N_11630,N_9536);
or U12423 (N_12423,N_11684,N_10709);
nor U12424 (N_12424,N_10966,N_11264);
xnor U12425 (N_12425,N_11795,N_10439);
or U12426 (N_12426,N_10825,N_11571);
nand U12427 (N_12427,N_10837,N_9293);
nor U12428 (N_12428,N_10080,N_9048);
nor U12429 (N_12429,N_10105,N_11083);
and U12430 (N_12430,N_9306,N_10081);
or U12431 (N_12431,N_11574,N_10928);
xor U12432 (N_12432,N_11856,N_9637);
and U12433 (N_12433,N_9758,N_11274);
nand U12434 (N_12434,N_9417,N_10994);
or U12435 (N_12435,N_9700,N_9958);
and U12436 (N_12436,N_11187,N_9086);
and U12437 (N_12437,N_11258,N_11686);
xnor U12438 (N_12438,N_9537,N_11091);
and U12439 (N_12439,N_9945,N_11504);
and U12440 (N_12440,N_11553,N_10749);
or U12441 (N_12441,N_10814,N_10503);
and U12442 (N_12442,N_9444,N_10945);
nor U12443 (N_12443,N_9793,N_10000);
nor U12444 (N_12444,N_9869,N_10166);
nor U12445 (N_12445,N_10250,N_10894);
nand U12446 (N_12446,N_11349,N_11250);
nor U12447 (N_12447,N_11338,N_10748);
xor U12448 (N_12448,N_11332,N_9476);
xor U12449 (N_12449,N_11287,N_10036);
or U12450 (N_12450,N_10635,N_11954);
nand U12451 (N_12451,N_10890,N_10152);
nand U12452 (N_12452,N_11636,N_9792);
nor U12453 (N_12453,N_10144,N_9607);
nand U12454 (N_12454,N_9790,N_11304);
nand U12455 (N_12455,N_11023,N_9665);
nor U12456 (N_12456,N_10346,N_11700);
or U12457 (N_12457,N_9249,N_11401);
nand U12458 (N_12458,N_10430,N_10950);
xnor U12459 (N_12459,N_9341,N_11366);
xor U12460 (N_12460,N_11263,N_11828);
or U12461 (N_12461,N_11054,N_9856);
xor U12462 (N_12462,N_9540,N_10839);
or U12463 (N_12463,N_10582,N_10877);
and U12464 (N_12464,N_11969,N_10499);
nor U12465 (N_12465,N_9418,N_9079);
and U12466 (N_12466,N_9964,N_11612);
nand U12467 (N_12467,N_11549,N_10335);
nor U12468 (N_12468,N_11533,N_11221);
nor U12469 (N_12469,N_9363,N_10831);
and U12470 (N_12470,N_11008,N_10217);
nor U12471 (N_12471,N_11839,N_11916);
nand U12472 (N_12472,N_10416,N_9756);
nand U12473 (N_12473,N_10240,N_11777);
xor U12474 (N_12474,N_10083,N_10937);
nor U12475 (N_12475,N_11813,N_10393);
and U12476 (N_12476,N_9781,N_10436);
or U12477 (N_12477,N_9718,N_11550);
or U12478 (N_12478,N_9764,N_10037);
nand U12479 (N_12479,N_11279,N_9520);
or U12480 (N_12480,N_9579,N_10333);
xor U12481 (N_12481,N_9487,N_11796);
or U12482 (N_12482,N_11074,N_11036);
or U12483 (N_12483,N_11331,N_10135);
or U12484 (N_12484,N_9401,N_9358);
or U12485 (N_12485,N_9302,N_10549);
nor U12486 (N_12486,N_11400,N_10559);
and U12487 (N_12487,N_10804,N_9246);
or U12488 (N_12488,N_11852,N_11275);
and U12489 (N_12489,N_10462,N_11206);
or U12490 (N_12490,N_10819,N_10838);
nor U12491 (N_12491,N_11268,N_11308);
xnor U12492 (N_12492,N_9269,N_9995);
xnor U12493 (N_12493,N_9077,N_9212);
and U12494 (N_12494,N_9106,N_9541);
or U12495 (N_12495,N_11738,N_11494);
nand U12496 (N_12496,N_10321,N_10618);
xor U12497 (N_12497,N_10543,N_9105);
or U12498 (N_12498,N_11341,N_11058);
nand U12499 (N_12499,N_9216,N_10963);
and U12500 (N_12500,N_9420,N_10613);
nor U12501 (N_12501,N_10807,N_9343);
nand U12502 (N_12502,N_10262,N_9904);
or U12503 (N_12503,N_10171,N_11908);
xnor U12504 (N_12504,N_9581,N_9557);
nand U12505 (N_12505,N_11588,N_10968);
nor U12506 (N_12506,N_11826,N_9470);
or U12507 (N_12507,N_9088,N_10131);
or U12508 (N_12508,N_9872,N_9247);
xor U12509 (N_12509,N_11144,N_11808);
xor U12510 (N_12510,N_10164,N_10042);
nand U12511 (N_12511,N_11698,N_10938);
and U12512 (N_12512,N_10252,N_11554);
or U12513 (N_12513,N_10420,N_10127);
nor U12514 (N_12514,N_9956,N_11766);
nor U12515 (N_12515,N_9339,N_9342);
or U12516 (N_12516,N_9909,N_9996);
nor U12517 (N_12517,N_10238,N_11352);
nor U12518 (N_12518,N_10941,N_10978);
nor U12519 (N_12519,N_9225,N_10598);
or U12520 (N_12520,N_9155,N_11198);
xnor U12521 (N_12521,N_9136,N_11927);
or U12522 (N_12522,N_10192,N_10072);
or U12523 (N_12523,N_11329,N_9740);
nand U12524 (N_12524,N_11650,N_11022);
or U12525 (N_12525,N_9701,N_11772);
nand U12526 (N_12526,N_9860,N_9854);
or U12527 (N_12527,N_10242,N_9356);
or U12528 (N_12528,N_11889,N_9528);
and U12529 (N_12529,N_11163,N_9585);
nand U12530 (N_12530,N_10479,N_11355);
xor U12531 (N_12531,N_9578,N_9010);
and U12532 (N_12532,N_10544,N_10396);
nor U12533 (N_12533,N_9328,N_9489);
and U12534 (N_12534,N_11623,N_9866);
xor U12535 (N_12535,N_10948,N_11673);
xnor U12536 (N_12536,N_9107,N_9565);
xnor U12537 (N_12537,N_10509,N_10150);
nor U12538 (N_12538,N_10507,N_9959);
xnor U12539 (N_12539,N_11192,N_10952);
or U12540 (N_12540,N_11364,N_10155);
or U12541 (N_12541,N_9658,N_11378);
xor U12542 (N_12542,N_11564,N_9709);
nand U12543 (N_12543,N_11457,N_11516);
nand U12544 (N_12544,N_11974,N_11609);
or U12545 (N_12545,N_9857,N_10658);
or U12546 (N_12546,N_10607,N_9441);
and U12547 (N_12547,N_11060,N_9387);
and U12548 (N_12548,N_9863,N_11948);
xor U12549 (N_12549,N_10692,N_10434);
and U12550 (N_12550,N_10656,N_10912);
or U12551 (N_12551,N_9878,N_9112);
and U12552 (N_12552,N_9219,N_9184);
nor U12553 (N_12553,N_9716,N_10103);
and U12554 (N_12554,N_9250,N_10642);
nand U12555 (N_12555,N_10965,N_9974);
nor U12556 (N_12556,N_11376,N_10747);
or U12557 (N_12557,N_11987,N_10835);
and U12558 (N_12558,N_10933,N_9710);
nor U12559 (N_12559,N_11330,N_11930);
or U12560 (N_12560,N_11188,N_10581);
or U12561 (N_12561,N_11685,N_9186);
xnor U12562 (N_12562,N_10100,N_11812);
nand U12563 (N_12563,N_11095,N_9469);
or U12564 (N_12564,N_9591,N_9760);
and U12565 (N_12565,N_11934,N_9132);
nor U12566 (N_12566,N_11608,N_10708);
xor U12567 (N_12567,N_11334,N_11784);
nand U12568 (N_12568,N_11517,N_10304);
nand U12569 (N_12569,N_9182,N_11960);
nor U12570 (N_12570,N_10700,N_10881);
and U12571 (N_12571,N_11130,N_11779);
or U12572 (N_12572,N_9632,N_9893);
and U12573 (N_12573,N_9671,N_11682);
nor U12574 (N_12574,N_9081,N_11830);
nand U12575 (N_12575,N_10878,N_9006);
nor U12576 (N_12576,N_10811,N_9023);
xor U12577 (N_12577,N_10883,N_11515);
nor U12578 (N_12578,N_10654,N_9289);
and U12579 (N_12579,N_11774,N_11403);
xnor U12580 (N_12580,N_9361,N_11928);
or U12581 (N_12581,N_11180,N_11132);
and U12582 (N_12582,N_11136,N_10049);
xnor U12583 (N_12583,N_9606,N_9755);
nor U12584 (N_12584,N_10573,N_9175);
nor U12585 (N_12585,N_10951,N_9396);
and U12586 (N_12586,N_11289,N_10244);
xnor U12587 (N_12587,N_9442,N_9845);
xor U12588 (N_12588,N_9666,N_11864);
xor U12589 (N_12589,N_11335,N_10829);
and U12590 (N_12590,N_10034,N_11428);
or U12591 (N_12591,N_10611,N_11232);
and U12592 (N_12592,N_9144,N_10003);
nand U12593 (N_12593,N_9075,N_11931);
and U12594 (N_12594,N_11122,N_11441);
xor U12595 (N_12595,N_10954,N_10974);
nand U12596 (N_12596,N_10481,N_10704);
xor U12597 (N_12597,N_9943,N_10592);
xor U12598 (N_12598,N_10834,N_11088);
or U12599 (N_12599,N_9435,N_11953);
xnor U12600 (N_12600,N_11734,N_11526);
nor U12601 (N_12601,N_9731,N_9232);
and U12602 (N_12602,N_10666,N_11035);
xnor U12603 (N_12603,N_10972,N_10911);
nand U12604 (N_12604,N_9506,N_11988);
xor U12605 (N_12605,N_9574,N_9030);
or U12606 (N_12606,N_10808,N_10750);
xnor U12607 (N_12607,N_9816,N_9207);
and U12608 (N_12608,N_11995,N_10223);
nor U12609 (N_12609,N_9794,N_10815);
xnor U12610 (N_12610,N_10969,N_11252);
nor U12611 (N_12611,N_9651,N_9142);
or U12612 (N_12612,N_10859,N_10627);
nor U12613 (N_12613,N_9994,N_11277);
xnor U12614 (N_12614,N_9598,N_11370);
and U12615 (N_12615,N_9779,N_11181);
nand U12616 (N_12616,N_9012,N_11941);
or U12617 (N_12617,N_10645,N_9021);
nand U12618 (N_12618,N_11383,N_9348);
nor U12619 (N_12619,N_11751,N_11432);
or U12620 (N_12620,N_10504,N_11842);
xor U12621 (N_12621,N_11464,N_11260);
and U12622 (N_12622,N_10399,N_9305);
and U12623 (N_12623,N_10079,N_9526);
and U12624 (N_12624,N_9102,N_11753);
nor U12625 (N_12625,N_11409,N_9595);
and U12626 (N_12626,N_10455,N_10320);
or U12627 (N_12627,N_10496,N_9953);
xnor U12628 (N_12628,N_10090,N_11129);
nor U12629 (N_12629,N_9825,N_10698);
xor U12630 (N_12630,N_10888,N_9091);
nand U12631 (N_12631,N_9278,N_9130);
and U12632 (N_12632,N_10849,N_9052);
nor U12633 (N_12633,N_9321,N_10823);
or U12634 (N_12634,N_10257,N_11238);
or U12635 (N_12635,N_11174,N_9949);
xor U12636 (N_12636,N_11985,N_10944);
nand U12637 (N_12637,N_10102,N_9074);
nor U12638 (N_12638,N_11085,N_9577);
nor U12639 (N_12639,N_10551,N_11750);
nand U12640 (N_12640,N_11791,N_9245);
or U12641 (N_12641,N_11863,N_9371);
nor U12642 (N_12642,N_9523,N_10567);
or U12643 (N_12643,N_9282,N_10245);
xnor U12644 (N_12644,N_10379,N_11442);
xnor U12645 (N_12645,N_11507,N_9322);
nor U12646 (N_12646,N_10677,N_11140);
nor U12647 (N_12647,N_11600,N_10319);
and U12648 (N_12648,N_10999,N_9409);
and U12649 (N_12649,N_10476,N_9485);
xor U12650 (N_12650,N_11973,N_11506);
nand U12651 (N_12651,N_9824,N_10030);
and U12652 (N_12652,N_10361,N_10497);
nand U12653 (N_12653,N_11963,N_9554);
nand U12654 (N_12654,N_9823,N_11133);
nor U12655 (N_12655,N_11281,N_11137);
nand U12656 (N_12656,N_9419,N_11798);
nand U12657 (N_12657,N_9060,N_11077);
or U12658 (N_12658,N_11848,N_10344);
and U12659 (N_12659,N_11177,N_11297);
and U12660 (N_12660,N_9049,N_9689);
nand U12661 (N_12661,N_10765,N_9196);
and U12662 (N_12662,N_9213,N_11855);
and U12663 (N_12663,N_11501,N_11762);
and U12664 (N_12664,N_11407,N_9973);
and U12665 (N_12665,N_9058,N_10071);
or U12666 (N_12666,N_9288,N_9389);
xnor U12667 (N_12667,N_9655,N_9993);
or U12668 (N_12668,N_10850,N_9936);
nand U12669 (N_12669,N_10219,N_11374);
nand U12670 (N_12670,N_10716,N_10556);
and U12671 (N_12671,N_11160,N_9805);
and U12672 (N_12672,N_9195,N_10007);
and U12673 (N_12673,N_11967,N_11810);
or U12674 (N_12674,N_10014,N_10454);
or U12675 (N_12675,N_9035,N_9449);
xnor U12676 (N_12676,N_9149,N_11894);
or U12677 (N_12677,N_9705,N_10852);
nand U12678 (N_12678,N_10953,N_9978);
or U12679 (N_12679,N_9544,N_10900);
and U12680 (N_12680,N_11112,N_10445);
and U12681 (N_12681,N_9890,N_9261);
nand U12682 (N_12682,N_11892,N_11755);
nand U12683 (N_12683,N_11895,N_11620);
or U12684 (N_12684,N_9751,N_9378);
and U12685 (N_12685,N_11531,N_9882);
xnor U12686 (N_12686,N_9237,N_11545);
nor U12687 (N_12687,N_9986,N_9284);
nand U12688 (N_12688,N_9734,N_10917);
nand U12689 (N_12689,N_10054,N_11843);
xnor U12690 (N_12690,N_10345,N_11288);
or U12691 (N_12691,N_11802,N_11314);
xnor U12692 (N_12692,N_9181,N_9521);
or U12693 (N_12693,N_10672,N_11212);
or U12694 (N_12694,N_10892,N_11729);
xnor U12695 (N_12695,N_11540,N_10800);
nand U12696 (N_12696,N_11801,N_10066);
or U12697 (N_12697,N_10210,N_11090);
nor U12698 (N_12698,N_10263,N_10536);
xnor U12699 (N_12699,N_10898,N_11099);
nor U12700 (N_12700,N_11115,N_9462);
nand U12701 (N_12701,N_10147,N_10114);
and U12702 (N_12702,N_11631,N_11626);
nor U12703 (N_12703,N_10337,N_9118);
or U12704 (N_12704,N_9631,N_9798);
and U12705 (N_12705,N_10339,N_10278);
nor U12706 (N_12706,N_11546,N_9116);
nor U12707 (N_12707,N_10178,N_9068);
nor U12708 (N_12708,N_10830,N_11080);
nand U12709 (N_12709,N_10265,N_9000);
and U12710 (N_12710,N_9391,N_10516);
xor U12711 (N_12711,N_11599,N_9344);
xnor U12712 (N_12712,N_11084,N_10641);
nand U12713 (N_12713,N_9673,N_10665);
nor U12714 (N_12714,N_9732,N_11390);
or U12715 (N_12715,N_10258,N_10044);
nand U12716 (N_12716,N_11067,N_9123);
xnor U12717 (N_12717,N_11014,N_9051);
nand U12718 (N_12718,N_11065,N_9242);
and U12719 (N_12719,N_11873,N_10157);
xnor U12720 (N_12720,N_11408,N_9723);
and U12721 (N_12721,N_11876,N_11076);
and U12722 (N_12722,N_11952,N_10557);
and U12723 (N_12723,N_9386,N_9031);
nand U12724 (N_12724,N_9622,N_11675);
nand U12725 (N_12725,N_11222,N_10380);
and U12726 (N_12726,N_11759,N_11471);
or U12727 (N_12727,N_10024,N_11725);
or U12728 (N_12728,N_11543,N_9877);
nor U12729 (N_12729,N_10411,N_9095);
nor U12730 (N_12730,N_11011,N_9126);
nor U12731 (N_12731,N_9256,N_11202);
xnor U12732 (N_12732,N_9616,N_10149);
xor U12733 (N_12733,N_9464,N_10176);
xnor U12734 (N_12734,N_11446,N_10916);
nor U12735 (N_12735,N_11692,N_11622);
and U12736 (N_12736,N_10195,N_9727);
or U12737 (N_12737,N_9338,N_9780);
nor U12738 (N_12738,N_10055,N_11348);
or U12739 (N_12739,N_11735,N_11658);
or U12740 (N_12740,N_9159,N_10662);
or U12741 (N_12741,N_10226,N_10116);
xor U12742 (N_12742,N_10283,N_9813);
or U12743 (N_12743,N_11899,N_10793);
nand U12744 (N_12744,N_11482,N_9745);
nand U12745 (N_12745,N_10160,N_11495);
xnor U12746 (N_12746,N_10267,N_11207);
nand U12747 (N_12747,N_10629,N_10524);
and U12748 (N_12748,N_9366,N_9215);
and U12749 (N_12749,N_9589,N_11470);
xnor U12750 (N_12750,N_9814,N_10452);
xnor U12751 (N_12751,N_10895,N_11721);
and U12752 (N_12752,N_10317,N_9839);
and U12753 (N_12753,N_11628,N_11959);
or U12754 (N_12754,N_11045,N_11472);
nand U12755 (N_12755,N_9017,N_9494);
or U12756 (N_12756,N_9239,N_10738);
nand U12757 (N_12757,N_9931,N_9162);
xor U12758 (N_12758,N_10981,N_11668);
or U12759 (N_12759,N_10918,N_10547);
nand U12760 (N_12760,N_11108,N_11498);
or U12761 (N_12761,N_11324,N_9410);
xnor U12762 (N_12762,N_10227,N_11344);
or U12763 (N_12763,N_9352,N_11351);
and U12764 (N_12764,N_10534,N_9156);
and U12765 (N_12765,N_11009,N_10777);
or U12766 (N_12766,N_9575,N_11233);
nand U12767 (N_12767,N_10405,N_11026);
and U12768 (N_12768,N_9900,N_9241);
or U12769 (N_12769,N_10967,N_11278);
nand U12770 (N_12770,N_10382,N_10754);
nand U12771 (N_12771,N_9924,N_11094);
xnor U12772 (N_12772,N_10253,N_11057);
or U12773 (N_12773,N_11373,N_11053);
nand U12774 (N_12774,N_10853,N_11949);
or U12775 (N_12775,N_11113,N_9980);
nor U12776 (N_12776,N_10425,N_10683);
xnor U12777 (N_12777,N_10064,N_9096);
xnor U12778 (N_12778,N_10163,N_10297);
xnor U12779 (N_12779,N_9970,N_11128);
and U12780 (N_12780,N_10653,N_9427);
nor U12781 (N_12781,N_11534,N_10012);
or U12782 (N_12782,N_10389,N_11424);
xor U12783 (N_12783,N_11305,N_10605);
and U12784 (N_12784,N_11072,N_10576);
nor U12785 (N_12785,N_10457,N_10121);
or U12786 (N_12786,N_10886,N_11454);
nor U12787 (N_12787,N_10841,N_10241);
nand U12788 (N_12788,N_10212,N_11602);
xnor U12789 (N_12789,N_10290,N_10493);
nor U12790 (N_12790,N_10620,N_10752);
and U12791 (N_12791,N_9743,N_10676);
and U12792 (N_12792,N_10228,N_11986);
and U12793 (N_12793,N_11301,N_9163);
and U12794 (N_12794,N_10391,N_9687);
and U12795 (N_12795,N_11757,N_10589);
and U12796 (N_12796,N_10906,N_9066);
xnor U12797 (N_12797,N_11551,N_11394);
or U12798 (N_12798,N_9452,N_10914);
or U12799 (N_12799,N_9667,N_10538);
xnor U12800 (N_12800,N_9152,N_10776);
nand U12801 (N_12801,N_11497,N_9532);
and U12802 (N_12802,N_10272,N_9005);
nand U12803 (N_12803,N_11271,N_11580);
nor U12804 (N_12804,N_9461,N_9826);
and U12805 (N_12805,N_11958,N_9413);
and U12806 (N_12806,N_11525,N_10040);
xnor U12807 (N_12807,N_11875,N_10517);
and U12808 (N_12808,N_10186,N_11360);
xor U12809 (N_12809,N_11185,N_9405);
or U12810 (N_12810,N_9501,N_9202);
or U12811 (N_12811,N_9143,N_10035);
and U12812 (N_12812,N_11345,N_10028);
nand U12813 (N_12813,N_11585,N_10514);
xnor U12814 (N_12814,N_11655,N_11583);
nor U12815 (N_12815,N_11121,N_9855);
nor U12816 (N_12816,N_11100,N_10940);
nor U12817 (N_12817,N_9568,N_11577);
nand U12818 (N_12818,N_9947,N_10775);
or U12819 (N_12819,N_9355,N_11674);
nand U12820 (N_12820,N_11171,N_11888);
or U12821 (N_12821,N_9319,N_9549);
and U12822 (N_12822,N_10923,N_10429);
nand U12823 (N_12823,N_9236,N_11805);
and U12824 (N_12824,N_11552,N_9720);
xnor U12825 (N_12825,N_10095,N_10381);
and U12826 (N_12826,N_9645,N_9822);
nor U12827 (N_12827,N_10023,N_11157);
and U12828 (N_12828,N_10805,N_11306);
and U12829 (N_12829,N_9602,N_9957);
or U12830 (N_12830,N_10647,N_9722);
xor U12831 (N_12831,N_9046,N_11837);
or U12832 (N_12832,N_10904,N_9552);
xnor U12833 (N_12833,N_10450,N_11811);
nand U12834 (N_12834,N_9114,N_9061);
nand U12835 (N_12835,N_11249,N_10533);
nor U12836 (N_12836,N_11632,N_9160);
and U12837 (N_12837,N_9018,N_10701);
and U12838 (N_12838,N_9721,N_11209);
xor U12839 (N_12839,N_9038,N_10566);
xor U12840 (N_12840,N_10483,N_11872);
or U12841 (N_12841,N_11152,N_10312);
or U12842 (N_12842,N_10022,N_10062);
xnor U12843 (N_12843,N_9097,N_11593);
nor U12844 (N_12844,N_10767,N_10599);
nor U12845 (N_12845,N_9991,N_11066);
or U12846 (N_12846,N_10943,N_11283);
nand U12847 (N_12847,N_11193,N_10082);
nor U12848 (N_12848,N_10357,N_9374);
nor U12849 (N_12849,N_11491,N_9224);
nand U12850 (N_12850,N_11881,N_10619);
nand U12851 (N_12851,N_10352,N_10004);
or U12852 (N_12852,N_10932,N_10484);
xnor U12853 (N_12853,N_9345,N_9728);
nor U12854 (N_12854,N_9309,N_10305);
nand U12855 (N_12855,N_10760,N_10970);
nor U12856 (N_12856,N_9291,N_10203);
nand U12857 (N_12857,N_10962,N_11711);
or U12858 (N_12858,N_11189,N_11496);
and U12859 (N_12859,N_10115,N_11786);
nand U12860 (N_12860,N_9623,N_10910);
nand U12861 (N_12861,N_9961,N_9416);
nand U12862 (N_12862,N_9166,N_9210);
and U12863 (N_12863,N_11956,N_11006);
or U12864 (N_12864,N_9896,N_9871);
or U12865 (N_12865,N_9243,N_9534);
and U12866 (N_12866,N_9503,N_9300);
and U12867 (N_12867,N_9065,N_11878);
xor U12868 (N_12868,N_11365,N_11560);
or U12869 (N_12869,N_11672,N_10225);
xnor U12870 (N_12870,N_11687,N_11598);
or U12871 (N_12871,N_9332,N_9567);
or U12872 (N_12872,N_10922,N_11038);
xnor U12873 (N_12873,N_10848,N_10363);
and U12874 (N_12874,N_11051,N_11216);
nand U12875 (N_12875,N_9550,N_11205);
nand U12876 (N_12876,N_11484,N_9775);
xnor U12877 (N_12877,N_11183,N_10438);
or U12878 (N_12878,N_11310,N_9560);
nor U12879 (N_12879,N_9411,N_11184);
xor U12880 (N_12880,N_9360,N_9989);
and U12881 (N_12881,N_9608,N_10324);
xor U12882 (N_12882,N_9982,N_11867);
xnor U12883 (N_12883,N_11971,N_10088);
nand U12884 (N_12884,N_9408,N_11261);
xor U12885 (N_12885,N_9761,N_9100);
nor U12886 (N_12886,N_11485,N_11641);
or U12887 (N_12887,N_9428,N_11218);
nand U12888 (N_12888,N_11901,N_10031);
and U12889 (N_12889,N_9087,N_10084);
nor U12890 (N_12890,N_9584,N_10897);
and U12891 (N_12891,N_10833,N_10373);
and U12892 (N_12892,N_9412,N_10246);
xnor U12893 (N_12893,N_10707,N_11123);
xor U12894 (N_12894,N_10125,N_11586);
nor U12895 (N_12895,N_10563,N_11191);
nand U12896 (N_12896,N_11651,N_11270);
nor U12897 (N_12897,N_11965,N_11414);
nand U12898 (N_12898,N_10018,N_11800);
nor U12899 (N_12899,N_9827,N_11230);
nand U12900 (N_12900,N_9875,N_11723);
and U12901 (N_12901,N_11749,N_9276);
xor U12902 (N_12902,N_11592,N_11450);
nor U12903 (N_12903,N_10946,N_9007);
nor U12904 (N_12904,N_11012,N_9330);
and U12905 (N_12905,N_11887,N_9812);
xnor U12906 (N_12906,N_9271,N_11594);
nor U12907 (N_12907,N_9480,N_9482);
xor U12908 (N_12908,N_11259,N_10006);
xnor U12909 (N_12909,N_10038,N_9050);
nand U12910 (N_12910,N_11752,N_11033);
nand U12911 (N_12911,N_9913,N_10208);
xor U12912 (N_12912,N_10369,N_9851);
nor U12913 (N_12913,N_9206,N_10971);
xor U12914 (N_12914,N_9161,N_10087);
xor U12915 (N_12915,N_10960,N_11047);
nand U12916 (N_12916,N_10565,N_10846);
xnor U12917 (N_12917,N_11448,N_10771);
nand U12918 (N_12918,N_11417,N_9253);
and U12919 (N_12919,N_9685,N_11291);
and U12920 (N_12920,N_11050,N_10327);
nor U12921 (N_12921,N_9738,N_10161);
or U12922 (N_12922,N_10675,N_9171);
nand U12923 (N_12923,N_9128,N_9776);
or U12924 (N_12924,N_10663,N_10870);
xnor U12925 (N_12925,N_11992,N_10368);
nor U12926 (N_12926,N_11015,N_11555);
nand U12927 (N_12927,N_11726,N_11836);
or U12928 (N_12928,N_10426,N_10578);
nand U12929 (N_12929,N_11154,N_10218);
or U12930 (N_12930,N_9599,N_11618);
nor U12931 (N_12931,N_11566,N_10980);
nand U12932 (N_12932,N_10545,N_11262);
and U12933 (N_12933,N_9392,N_9450);
or U12934 (N_12934,N_10809,N_9054);
nor U12935 (N_12935,N_10734,N_10623);
xnor U12936 (N_12936,N_9477,N_10577);
nor U12937 (N_12937,N_9511,N_11247);
or U12938 (N_12938,N_10169,N_10688);
nor U12939 (N_12939,N_11505,N_10818);
or U12940 (N_12940,N_9992,N_10353);
and U12941 (N_12941,N_10891,N_10027);
and U12942 (N_12942,N_10085,N_10232);
nor U12943 (N_12943,N_9071,N_11469);
nand U12944 (N_12944,N_9294,N_11150);
nor U12945 (N_12945,N_9436,N_9912);
and U12946 (N_12946,N_10282,N_9590);
or U12947 (N_12947,N_11694,N_9844);
or U12948 (N_12948,N_10732,N_9883);
xor U12949 (N_12949,N_9125,N_11640);
xnor U12950 (N_12950,N_11257,N_11886);
nand U12951 (N_12951,N_9997,N_9657);
xor U12952 (N_12952,N_10307,N_9914);
nand U12953 (N_12953,N_11078,N_9514);
xor U12954 (N_12954,N_10446,N_9209);
nor U12955 (N_12955,N_10786,N_10206);
xnor U12956 (N_12956,N_9180,N_9120);
xor U12957 (N_12957,N_9178,N_11521);
nor U12958 (N_12958,N_11697,N_9456);
or U12959 (N_12959,N_11522,N_9299);
and U12960 (N_12960,N_10402,N_11031);
xor U12961 (N_12961,N_10059,N_10822);
or U12962 (N_12962,N_11357,N_10625);
or U12963 (N_12963,N_10394,N_10571);
nor U12964 (N_12964,N_10205,N_10537);
nor U12965 (N_12965,N_11290,N_11002);
or U12966 (N_12966,N_11817,N_11280);
xor U12967 (N_12967,N_10332,N_10590);
nor U12968 (N_12968,N_9968,N_10032);
or U12969 (N_12969,N_10842,N_9365);
nor U12970 (N_12970,N_10518,N_9252);
nand U12971 (N_12971,N_11021,N_11676);
or U12972 (N_12972,N_11542,N_10828);
and U12973 (N_12973,N_10626,N_10821);
xor U12974 (N_12974,N_10600,N_10991);
nor U12975 (N_12975,N_10478,N_10112);
xnor U12976 (N_12976,N_9677,N_9985);
or U12977 (N_12977,N_9211,N_10029);
xor U12978 (N_12978,N_9942,N_9747);
or U12979 (N_12979,N_11046,N_11922);
nand U12980 (N_12980,N_9773,N_10615);
nand U12981 (N_12981,N_9907,N_9218);
nor U12982 (N_12982,N_11920,N_9848);
xor U12983 (N_12983,N_10415,N_9203);
nand U12984 (N_12984,N_11229,N_11211);
and U12985 (N_12985,N_9990,N_9630);
nor U12986 (N_12986,N_10325,N_9646);
nand U12987 (N_12987,N_11699,N_9296);
nor U12988 (N_12988,N_10143,N_10453);
xnor U12989 (N_12989,N_11125,N_9897);
nand U12990 (N_12990,N_11398,N_11568);
nand U12991 (N_12991,N_11226,N_10097);
nand U12992 (N_12992,N_10640,N_10633);
or U12993 (N_12993,N_9307,N_10731);
nor U12994 (N_12994,N_11131,N_10296);
and U12995 (N_12995,N_9093,N_9865);
and U12996 (N_12996,N_10274,N_11972);
nor U12997 (N_12997,N_10404,N_10779);
nand U12998 (N_12998,N_11819,N_9522);
nor U12999 (N_12999,N_11005,N_11126);
nor U13000 (N_13000,N_11627,N_10715);
xor U13001 (N_13001,N_11999,N_9605);
and U13002 (N_13002,N_10761,N_9274);
or U13003 (N_13003,N_11303,N_11670);
and U13004 (N_13004,N_10322,N_9859);
nor U13005 (N_13005,N_11354,N_10284);
xor U13006 (N_13006,N_10433,N_10148);
nand U13007 (N_13007,N_11285,N_11186);
nor U13008 (N_13008,N_9495,N_9563);
nor U13009 (N_13009,N_11087,N_11718);
nand U13010 (N_13010,N_11266,N_9853);
xnor U13011 (N_13011,N_11572,N_11990);
nor U13012 (N_13012,N_10772,N_11576);
nand U13013 (N_13013,N_10521,N_10603);
xnor U13014 (N_13014,N_9729,N_10421);
and U13015 (N_13015,N_10744,N_9800);
or U13016 (N_13016,N_9407,N_11789);
and U13017 (N_13017,N_10492,N_10092);
xnor U13018 (N_13018,N_11379,N_10444);
nor U13019 (N_13019,N_10362,N_9131);
nand U13020 (N_13020,N_9220,N_11162);
or U13021 (N_13021,N_9594,N_10467);
or U13022 (N_13022,N_11269,N_11241);
nand U13023 (N_13023,N_11438,N_11426);
xor U13024 (N_13024,N_10746,N_9944);
or U13025 (N_13025,N_10222,N_9799);
xor U13026 (N_13026,N_10487,N_10057);
or U13027 (N_13027,N_10501,N_9587);
nor U13028 (N_13028,N_10992,N_10588);
and U13029 (N_13029,N_10281,N_9334);
nor U13030 (N_13030,N_9457,N_10142);
nor U13031 (N_13031,N_9040,N_9459);
xnor U13032 (N_13032,N_9672,N_9647);
or U13033 (N_13033,N_10955,N_11037);
and U13034 (N_13034,N_10360,N_11511);
or U13035 (N_13035,N_9259,N_11007);
nor U13036 (N_13036,N_11736,N_9884);
nor U13037 (N_13037,N_10495,N_11898);
and U13038 (N_13038,N_11642,N_10789);
nand U13039 (N_13039,N_10106,N_11547);
nand U13040 (N_13040,N_9624,N_9903);
nand U13041 (N_13041,N_9492,N_9888);
xor U13042 (N_13042,N_9744,N_11427);
nand U13043 (N_13043,N_11052,N_11778);
or U13044 (N_13044,N_9694,N_11282);
and U13045 (N_13045,N_11924,N_10542);
xnor U13046 (N_13046,N_9354,N_10026);
nor U13047 (N_13047,N_10884,N_10277);
or U13048 (N_13048,N_11251,N_9898);
xor U13049 (N_13049,N_11343,N_9119);
and U13050 (N_13050,N_9070,N_9569);
or U13051 (N_13051,N_11093,N_11857);
or U13052 (N_13052,N_9353,N_11166);
xnor U13053 (N_13053,N_11981,N_11859);
and U13054 (N_13054,N_10529,N_11539);
nand U13055 (N_13055,N_11604,N_10233);
nand U13056 (N_13056,N_11451,N_10119);
xor U13057 (N_13057,N_9762,N_9917);
xnor U13058 (N_13058,N_10287,N_11294);
nand U13059 (N_13059,N_10803,N_11197);
nand U13060 (N_13060,N_10302,N_11243);
nand U13061 (N_13061,N_11690,N_10655);
nor U13062 (N_13062,N_11767,N_11803);
and U13063 (N_13063,N_10107,N_9187);
nor U13064 (N_13064,N_10200,N_9019);
nand U13065 (N_13065,N_11747,N_10047);
or U13066 (N_13066,N_9894,N_10196);
nor U13067 (N_13067,N_9398,N_9273);
nor U13068 (N_13068,N_10089,N_9169);
or U13069 (N_13069,N_11977,N_11040);
nor U13070 (N_13070,N_9733,N_10033);
or U13071 (N_13071,N_10705,N_9383);
or U13072 (N_13072,N_11797,N_10078);
and U13073 (N_13073,N_11134,N_9693);
and U13074 (N_13074,N_11679,N_11149);
nor U13075 (N_13075,N_11064,N_11980);
or U13076 (N_13076,N_9041,N_10723);
nand U13077 (N_13077,N_9975,N_11486);
and U13078 (N_13078,N_10280,N_9434);
or U13079 (N_13079,N_9262,N_10553);
xnor U13080 (N_13080,N_9496,N_9786);
or U13081 (N_13081,N_10703,N_11994);
xor U13082 (N_13082,N_11467,N_11833);
xnor U13083 (N_13083,N_9692,N_9326);
nand U13084 (N_13084,N_9399,N_10770);
or U13085 (N_13085,N_9880,N_9015);
nor U13086 (N_13086,N_10477,N_10392);
and U13087 (N_13087,N_9644,N_11013);
nor U13088 (N_13088,N_9153,N_9530);
nor U13089 (N_13089,N_10198,N_10973);
and U13090 (N_13090,N_11807,N_9948);
and U13091 (N_13091,N_11387,N_11048);
nand U13092 (N_13092,N_11477,N_11874);
nand U13093 (N_13093,N_11939,N_10295);
nand U13094 (N_13094,N_11336,N_10717);
xor U13095 (N_13095,N_11102,N_11016);
and U13096 (N_13096,N_10410,N_11704);
and U13097 (N_13097,N_9566,N_11787);
xnor U13098 (N_13098,N_10956,N_11979);
nor U13099 (N_13099,N_11975,N_9555);
or U13100 (N_13100,N_9257,N_10294);
and U13101 (N_13101,N_9981,N_10398);
and U13102 (N_13102,N_11489,N_10591);
and U13103 (N_13103,N_10885,N_10301);
nor U13104 (N_13104,N_11681,N_9109);
nor U13105 (N_13105,N_10871,N_10468);
or U13106 (N_13106,N_9810,N_10907);
or U13107 (N_13107,N_10587,N_11317);
nor U13108 (N_13108,N_11142,N_9129);
nor U13109 (N_13109,N_10269,N_10882);
nor U13110 (N_13110,N_9821,N_9545);
xnor U13111 (N_13111,N_10270,N_10435);
nor U13112 (N_13112,N_9656,N_10984);
xnor U13113 (N_13113,N_9899,N_10136);
or U13114 (N_13114,N_9850,N_10138);
or U13115 (N_13115,N_10795,N_11851);
and U13116 (N_13116,N_9929,N_10329);
or U13117 (N_13117,N_9916,N_10860);
nor U13118 (N_13118,N_9999,N_11809);
or U13119 (N_13119,N_11481,N_10794);
or U13120 (N_13120,N_11818,N_11513);
nor U13121 (N_13121,N_10934,N_9777);
and U13122 (N_13122,N_11900,N_10365);
or U13123 (N_13123,N_11983,N_9254);
nand U13124 (N_13124,N_10093,N_11254);
and U13125 (N_13125,N_10569,N_10505);
and U13126 (N_13126,N_10713,N_10903);
nor U13127 (N_13127,N_11096,N_11322);
and U13128 (N_13128,N_10256,N_10580);
nand U13129 (N_13129,N_9954,N_11744);
xnor U13130 (N_13130,N_11453,N_9190);
nand U13131 (N_13131,N_11643,N_11043);
xnor U13132 (N_13132,N_11044,N_11649);
xor U13133 (N_13133,N_11082,N_9432);
nor U13134 (N_13134,N_9447,N_9911);
or U13135 (N_13135,N_10323,N_11326);
xnor U13136 (N_13136,N_10472,N_9939);
and U13137 (N_13137,N_11339,N_11705);
and U13138 (N_13138,N_11885,N_9454);
and U13139 (N_13139,N_10924,N_11678);
xor U13140 (N_13140,N_11677,N_10667);
xnor U13141 (N_13141,N_9199,N_11825);
nor U13142 (N_13142,N_10586,N_9580);
and U13143 (N_13143,N_11518,N_10069);
xor U13144 (N_13144,N_11785,N_11478);
and U13145 (N_13145,N_9089,N_11943);
nand U13146 (N_13146,N_9754,N_10858);
nand U13147 (N_13147,N_10001,N_10051);
or U13148 (N_13148,N_11849,N_10785);
nor U13149 (N_13149,N_11746,N_11030);
nor U13150 (N_13150,N_11701,N_10525);
nand U13151 (N_13151,N_10422,N_11788);
nor U13152 (N_13152,N_10936,N_10695);
nor U13153 (N_13153,N_10005,N_9533);
nor U13154 (N_13154,N_10099,N_9303);
or U13155 (N_13155,N_11388,N_9963);
xor U13156 (N_13156,N_9372,N_10338);
and U13157 (N_13157,N_11793,N_11028);
nand U13158 (N_13158,N_10735,N_11307);
nor U13159 (N_13159,N_9423,N_11661);
nor U13160 (N_13160,N_9194,N_10868);
or U13161 (N_13161,N_10751,N_9795);
xnor U13162 (N_13162,N_11146,N_11645);
and U13163 (N_13163,N_9029,N_10843);
xnor U13164 (N_13164,N_9286,N_11316);
and U13165 (N_13165,N_9643,N_9221);
xnor U13166 (N_13166,N_9504,N_9518);
nand U13167 (N_13167,N_11402,N_9650);
nand U13168 (N_13168,N_11127,N_11520);
and U13169 (N_13169,N_9527,N_10985);
nand U13170 (N_13170,N_10414,N_11944);
or U13171 (N_13171,N_10530,N_11079);
and U13172 (N_13172,N_9478,N_10989);
nor U13173 (N_13173,N_10865,N_9932);
or U13174 (N_13174,N_9287,N_11775);
or U13175 (N_13175,N_10528,N_11194);
nand U13176 (N_13176,N_9022,N_11201);
xor U13177 (N_13177,N_9508,N_10684);
or U13178 (N_13178,N_11933,N_11027);
nand U13179 (N_13179,N_11462,N_11227);
nor U13180 (N_13180,N_10275,N_10387);
nand U13181 (N_13181,N_10068,N_10575);
and U13182 (N_13182,N_9713,N_10926);
or U13183 (N_13183,N_9336,N_10710);
and U13184 (N_13184,N_11893,N_11156);
nor U13185 (N_13185,N_10726,N_11325);
xor U13186 (N_13186,N_11957,N_10728);
and U13187 (N_13187,N_10052,N_10260);
xor U13188 (N_13188,N_11713,N_9843);
and U13189 (N_13189,N_11561,N_9043);
and U13190 (N_13190,N_9763,N_11109);
or U13191 (N_13191,N_9785,N_9835);
nor U13192 (N_13192,N_9260,N_9670);
or U13193 (N_13193,N_9141,N_11595);
or U13194 (N_13194,N_10847,N_9263);
xor U13195 (N_13195,N_10612,N_9707);
or U13196 (N_13196,N_9099,N_10502);
nand U13197 (N_13197,N_9085,N_11664);
nor U13198 (N_13198,N_10632,N_11235);
and U13199 (N_13199,N_10753,N_11769);
nor U13200 (N_13200,N_11532,N_9467);
nor U13201 (N_13201,N_11865,N_9684);
nand U13202 (N_13202,N_10964,N_9191);
nand U13203 (N_13203,N_9059,N_9369);
xnor U13204 (N_13204,N_10929,N_11998);
xor U13205 (N_13205,N_9808,N_10011);
nand U13206 (N_13206,N_11110,N_11596);
or U13207 (N_13207,N_10456,N_9076);
and U13208 (N_13208,N_10721,N_11386);
xnor U13209 (N_13209,N_10584,N_10423);
and U13210 (N_13210,N_10927,N_11903);
xor U13211 (N_13211,N_11347,N_10298);
xnor U13212 (N_13212,N_11300,N_10845);
nor U13213 (N_13213,N_10259,N_10552);
nand U13214 (N_13214,N_9977,N_11337);
nand U13215 (N_13215,N_10383,N_9222);
nand U13216 (N_13216,N_9205,N_10401);
and U13217 (N_13217,N_10696,N_10740);
or U13218 (N_13218,N_9167,N_10374);
nand U13219 (N_13219,N_9507,N_9976);
nand U13220 (N_13220,N_11562,N_10021);
nor U13221 (N_13221,N_9473,N_10020);
or U13222 (N_13222,N_10739,N_9395);
or U13223 (N_13223,N_11302,N_10689);
nor U13224 (N_13224,N_11236,N_10879);
nand U13225 (N_13225,N_9791,N_10679);
nor U13226 (N_13226,N_9829,N_9867);
and U13227 (N_13227,N_11764,N_10314);
and U13228 (N_13228,N_10251,N_10550);
or U13229 (N_13229,N_9168,N_9390);
and U13230 (N_13230,N_11660,N_9001);
nor U13231 (N_13231,N_10636,N_9742);
nand U13232 (N_13232,N_10239,N_11841);
or U13233 (N_13233,N_11412,N_9983);
and U13234 (N_13234,N_11611,N_11880);
or U13235 (N_13235,N_9122,N_9788);
or U13236 (N_13236,N_9315,N_11393);
or U13237 (N_13237,N_9698,N_9200);
or U13238 (N_13238,N_11847,N_10649);
and U13239 (N_13239,N_9770,N_9703);
and U13240 (N_13240,N_10309,N_10844);
or U13241 (N_13241,N_11680,N_10867);
or U13242 (N_13242,N_11353,N_10076);
or U13243 (N_13243,N_9546,N_9879);
nor U13244 (N_13244,N_11821,N_9804);
nor U13245 (N_13245,N_9238,N_10315);
nor U13246 (N_13246,N_11062,N_9471);
or U13247 (N_13247,N_11714,N_11613);
or U13248 (N_13248,N_11716,N_9139);
nor U13249 (N_13249,N_11117,N_11107);
nor U13250 (N_13250,N_10229,N_10187);
nor U13251 (N_13251,N_11017,N_11204);
nand U13252 (N_13252,N_11139,N_10101);
nor U13253 (N_13253,N_10184,N_9367);
or U13254 (N_13254,N_10602,N_9836);
and U13255 (N_13255,N_11224,N_10403);
nor U13256 (N_13256,N_9270,N_10836);
nor U13257 (N_13257,N_11503,N_9925);
or U13258 (N_13258,N_11003,N_11092);
nor U13259 (N_13259,N_9753,N_9920);
or U13260 (N_13260,N_9660,N_9535);
nor U13261 (N_13261,N_10331,N_9801);
nor U13262 (N_13262,N_11689,N_11178);
or U13263 (N_13263,N_9682,N_11359);
xor U13264 (N_13264,N_10310,N_11947);
xor U13265 (N_13265,N_9415,N_11217);
nor U13266 (N_13266,N_11731,N_9265);
nand U13267 (N_13267,N_11653,N_11544);
or U13268 (N_13268,N_10506,N_9208);
or U13269 (N_13269,N_10094,N_11790);
or U13270 (N_13270,N_9268,N_11638);
xnor U13271 (N_13271,N_10191,N_10236);
or U13272 (N_13272,N_9045,N_11702);
xor U13273 (N_13273,N_9499,N_11597);
or U13274 (N_13274,N_9951,N_10697);
nand U13275 (N_13275,N_11089,N_9174);
or U13276 (N_13276,N_11029,N_10512);
nand U13277 (N_13277,N_9402,N_10604);
nand U13278 (N_13278,N_9741,N_11362);
nor U13279 (N_13279,N_9678,N_9483);
or U13280 (N_13280,N_11919,N_11662);
and U13281 (N_13281,N_10139,N_9324);
or U13282 (N_13282,N_11476,N_9014);
xnor U13283 (N_13283,N_9735,N_9641);
and U13284 (N_13284,N_11381,N_9629);
xor U13285 (N_13285,N_10921,N_10122);
nand U13286 (N_13286,N_10077,N_10899);
xnor U13287 (N_13287,N_10074,N_10986);
nand U13288 (N_13288,N_9151,N_10764);
xor U13289 (N_13289,N_11615,N_11635);
or U13290 (N_13290,N_11436,N_10661);
xnor U13291 (N_13291,N_11237,N_11292);
nand U13292 (N_13292,N_11902,N_11298);
nand U13293 (N_13293,N_11313,N_11814);
xnor U13294 (N_13294,N_9158,N_11748);
nand U13295 (N_13295,N_10714,N_10925);
nor U13296 (N_13296,N_9037,N_10797);
nand U13297 (N_13297,N_11358,N_11492);
nor U13298 (N_13298,N_11799,N_11182);
and U13299 (N_13299,N_10255,N_9769);
xnor U13300 (N_13300,N_11938,N_9008);
nor U13301 (N_13301,N_11104,N_9292);
nor U13302 (N_13302,N_10276,N_11276);
or U13303 (N_13303,N_9165,N_10893);
nor U13304 (N_13304,N_11086,N_11225);
nor U13305 (N_13305,N_11372,N_10720);
or U13306 (N_13306,N_10958,N_11159);
and U13307 (N_13307,N_9621,N_10976);
nand U13308 (N_13308,N_10668,N_9612);
xnor U13309 (N_13309,N_11273,N_11404);
and U13310 (N_13310,N_11850,N_9055);
and U13311 (N_13311,N_10041,N_9458);
or U13312 (N_13312,N_10447,N_9316);
nor U13313 (N_13313,N_11831,N_9807);
nor U13314 (N_13314,N_11116,N_10017);
xor U13315 (N_13315,N_11293,N_10370);
or U13316 (N_13316,N_9379,N_11020);
nor U13317 (N_13317,N_10762,N_11616);
nor U13318 (N_13318,N_9919,N_9073);
or U13319 (N_13319,N_10560,N_11587);
nand U13320 (N_13320,N_10690,N_10330);
nor U13321 (N_13321,N_11570,N_9750);
or U13322 (N_13322,N_9613,N_10670);
and U13323 (N_13323,N_11869,N_11782);
or U13324 (N_13324,N_10854,N_11169);
nor U13325 (N_13325,N_11563,N_10669);
and U13326 (N_13326,N_10820,N_10997);
xnor U13327 (N_13327,N_9586,N_9724);
and U13328 (N_13328,N_11897,N_11010);
xor U13329 (N_13329,N_10876,N_11460);
or U13330 (N_13330,N_11231,N_11913);
or U13331 (N_13331,N_10356,N_11648);
and U13332 (N_13332,N_9308,N_11246);
xor U13333 (N_13333,N_10133,N_9414);
and U13334 (N_13334,N_9712,N_10508);
or U13335 (N_13335,N_11418,N_11906);
nor U13336 (N_13336,N_9204,N_11120);
and U13337 (N_13337,N_11483,N_10465);
xnor U13338 (N_13338,N_9752,N_11905);
or U13339 (N_13339,N_9696,N_10596);
and U13340 (N_13340,N_10651,N_9138);
nand U13341 (N_13341,N_11732,N_10555);
and U13342 (N_13342,N_10664,N_11768);
nor U13343 (N_13343,N_9638,N_9493);
nand U13344 (N_13344,N_9725,N_10303);
and U13345 (N_13345,N_11656,N_10987);
nor U13346 (N_13346,N_9558,N_11173);
xnor U13347 (N_13347,N_11244,N_11220);
nor U13348 (N_13348,N_10326,N_10073);
nor U13349 (N_13349,N_9876,N_11499);
nor U13350 (N_13350,N_9176,N_11966);
and U13351 (N_13351,N_11168,N_9377);
and U13352 (N_13352,N_10742,N_11179);
and U13353 (N_13353,N_11073,N_10008);
or U13354 (N_13354,N_10098,N_9400);
and U13355 (N_13355,N_11621,N_11124);
and U13356 (N_13356,N_10527,N_11578);
and U13357 (N_13357,N_9519,N_11601);
xnor U13358 (N_13358,N_10901,N_9858);
nand U13359 (N_13359,N_10606,N_10230);
or U13360 (N_13360,N_9277,N_10488);
nand U13361 (N_13361,N_9115,N_9314);
nor U13362 (N_13362,N_9380,N_11996);
and U13363 (N_13363,N_9311,N_10146);
and U13364 (N_13364,N_10513,N_11647);
xor U13365 (N_13365,N_10207,N_11312);
nand U13366 (N_13366,N_11590,N_10384);
xnor U13367 (N_13367,N_11945,N_11909);
or U13368 (N_13368,N_9430,N_10182);
nor U13369 (N_13369,N_10075,N_11657);
xor U13370 (N_13370,N_9312,N_9784);
nor U13371 (N_13371,N_9453,N_10308);
nand U13372 (N_13372,N_11153,N_10168);
and U13373 (N_13373,N_9393,N_9831);
nand U13374 (N_13374,N_10802,N_10791);
or U13375 (N_13375,N_11717,N_9841);
nor U13376 (N_13376,N_11111,N_11508);
nor U13377 (N_13377,N_9382,N_10213);
or U13378 (N_13378,N_10614,N_10540);
nor U13379 (N_13379,N_11538,N_10526);
or U13380 (N_13380,N_9928,N_11614);
nor U13381 (N_13381,N_9895,N_10490);
and U13382 (N_13382,N_11579,N_9531);
and U13383 (N_13383,N_9668,N_10535);
nand U13384 (N_13384,N_9295,N_9064);
xor U13385 (N_13385,N_10159,N_10799);
and U13386 (N_13386,N_9962,N_9870);
xor U13387 (N_13387,N_10711,N_11871);
and U13388 (N_13388,N_10942,N_9778);
xnor U13389 (N_13389,N_9080,N_10486);
nor U13390 (N_13390,N_10220,N_10129);
nor U13391 (N_13391,N_11991,N_11770);
nor U13392 (N_13392,N_9782,N_10597);
and U13393 (N_13393,N_9230,N_9583);
nand U13394 (N_13394,N_9601,N_11610);
xnor U13395 (N_13395,N_11727,N_10247);
or U13396 (N_13396,N_10002,N_10010);
nor U13397 (N_13397,N_9627,N_9505);
xnor U13398 (N_13398,N_9266,N_11396);
nand U13399 (N_13399,N_10561,N_10046);
or U13400 (N_13400,N_10132,N_9304);
and U13401 (N_13401,N_11605,N_10113);
xor U13402 (N_13402,N_9433,N_9649);
xor U13403 (N_13403,N_9604,N_11773);
or U13404 (N_13404,N_11145,N_9614);
and U13405 (N_13405,N_10145,N_10480);
and U13406 (N_13406,N_11976,N_11135);
xnor U13407 (N_13407,N_11569,N_11740);
nand U13408 (N_13408,N_10110,N_10500);
nand U13409 (N_13409,N_10293,N_10905);
nor U13410 (N_13410,N_9783,N_9885);
nand U13411 (N_13411,N_9320,N_11844);
xnor U13412 (N_13412,N_11311,N_10162);
nor U13413 (N_13413,N_9538,N_10863);
nor U13414 (N_13414,N_9628,N_10817);
and U13415 (N_13415,N_9789,N_11103);
nand U13416 (N_13416,N_11443,N_10861);
and U13417 (N_13417,N_11055,N_10194);
and U13418 (N_13418,N_10644,N_10763);
nor U13419 (N_13419,N_11868,N_11377);
and U13420 (N_13420,N_10130,N_9938);
or U13421 (N_13421,N_11340,N_10299);
and U13422 (N_13422,N_10193,N_11950);
nand U13423 (N_13423,N_9923,N_11039);
nand U13424 (N_13424,N_9699,N_10862);
nand U13425 (N_13425,N_9652,N_11794);
nand U13426 (N_13426,N_10412,N_10254);
and U13427 (N_13427,N_11452,N_10729);
nor U13428 (N_13428,N_11652,N_9889);
nand U13429 (N_13429,N_11730,N_9950);
nand U13430 (N_13430,N_11415,N_10189);
xor U13431 (N_13431,N_10783,N_9362);
or U13432 (N_13432,N_9121,N_10197);
and U13433 (N_13433,N_11239,N_9466);
xor U13434 (N_13434,N_9437,N_10221);
nand U13435 (N_13435,N_11199,N_11917);
nand U13436 (N_13436,N_11397,N_9318);
and U13437 (N_13437,N_11328,N_10432);
nor U13438 (N_13438,N_10209,N_11929);
and U13439 (N_13439,N_11063,N_9381);
and U13440 (N_13440,N_11709,N_10261);
nand U13441 (N_13441,N_11639,N_9325);
or U13442 (N_13442,N_11951,N_11739);
xnor U13443 (N_13443,N_9539,N_9593);
and U13444 (N_13444,N_9927,N_11565);
and U13445 (N_13445,N_11001,N_9264);
and U13446 (N_13446,N_10673,N_11333);
and U13447 (N_13447,N_11196,N_9915);
nor U13448 (N_13448,N_11018,N_9516);
and U13449 (N_13449,N_9137,N_10140);
and U13450 (N_13450,N_10316,N_10790);
xor U13451 (N_13451,N_11419,N_11155);
nand U13452 (N_13452,N_11069,N_9240);
or U13453 (N_13453,N_9847,N_10108);
xnor U13454 (N_13454,N_11170,N_11537);
or U13455 (N_13455,N_10264,N_10935);
and U13456 (N_13456,N_11416,N_10019);
nor U13457 (N_13457,N_11820,N_11879);
or U13458 (N_13458,N_9193,N_11255);
or U13459 (N_13459,N_9227,N_10311);
and U13460 (N_13460,N_10988,N_9715);
or U13461 (N_13461,N_9524,N_9946);
and U13462 (N_13462,N_9662,N_11989);
or U13463 (N_13463,N_11523,N_10659);
and U13464 (N_13464,N_10413,N_9852);
nand U13465 (N_13465,N_9901,N_10856);
or U13466 (N_13466,N_10249,N_10624);
xnor U13467 (N_13467,N_9618,N_11213);
nand U13468 (N_13468,N_9809,N_9197);
and U13469 (N_13469,N_11323,N_9559);
nor U13470 (N_13470,N_9940,N_9164);
nor U13471 (N_13471,N_11743,N_11151);
nand U13472 (N_13472,N_11487,N_11804);
or U13473 (N_13473,N_9463,N_11845);
and U13474 (N_13474,N_11548,N_10489);
or U13475 (N_13475,N_11691,N_10902);
and U13476 (N_13476,N_11056,N_9244);
nand U13477 (N_13477,N_11936,N_9675);
or U13478 (N_13478,N_10334,N_11070);
and U13479 (N_13479,N_11025,N_11783);
nor U13480 (N_13480,N_10419,N_9830);
or U13481 (N_13481,N_11433,N_11710);
nand U13482 (N_13482,N_10039,N_10172);
nor U13483 (N_13483,N_9491,N_9748);
nor U13484 (N_13484,N_9134,N_9150);
and U13485 (N_13485,N_10058,N_11106);
or U13486 (N_13486,N_10609,N_10724);
xnor U13487 (N_13487,N_10806,N_10359);
nand U13488 (N_13488,N_11760,N_9472);
xnor U13489 (N_13489,N_9617,N_10211);
nand U13490 (N_13490,N_9484,N_9596);
or U13491 (N_13491,N_9290,N_10279);
and U13492 (N_13492,N_11771,N_11861);
or U13493 (N_13493,N_11984,N_10702);
xor U13494 (N_13494,N_9840,N_11248);
or U13495 (N_13495,N_11500,N_11633);
and U13496 (N_13496,N_11190,N_11395);
nand U13497 (N_13497,N_10630,N_9674);
and U13498 (N_13498,N_9488,N_9515);
xnor U13499 (N_13499,N_11490,N_10780);
xor U13500 (N_13500,N_10698,N_11644);
and U13501 (N_13501,N_11732,N_10408);
and U13502 (N_13502,N_10704,N_11024);
xor U13503 (N_13503,N_10928,N_9279);
nor U13504 (N_13504,N_11762,N_11000);
or U13505 (N_13505,N_11261,N_11018);
nor U13506 (N_13506,N_11215,N_11017);
and U13507 (N_13507,N_10990,N_10508);
nand U13508 (N_13508,N_10844,N_11473);
nand U13509 (N_13509,N_11814,N_10159);
xor U13510 (N_13510,N_9445,N_11906);
nand U13511 (N_13511,N_10866,N_10723);
and U13512 (N_13512,N_10994,N_9423);
xor U13513 (N_13513,N_9098,N_9593);
xnor U13514 (N_13514,N_10009,N_9696);
xor U13515 (N_13515,N_10122,N_10646);
xor U13516 (N_13516,N_9334,N_9037);
xor U13517 (N_13517,N_10307,N_9482);
or U13518 (N_13518,N_9471,N_9161);
nor U13519 (N_13519,N_10508,N_9411);
and U13520 (N_13520,N_9929,N_11016);
nor U13521 (N_13521,N_11801,N_11844);
xnor U13522 (N_13522,N_10598,N_9913);
or U13523 (N_13523,N_9096,N_10482);
xnor U13524 (N_13524,N_11137,N_10563);
nand U13525 (N_13525,N_10215,N_10226);
xor U13526 (N_13526,N_10040,N_11740);
and U13527 (N_13527,N_10994,N_11913);
or U13528 (N_13528,N_10432,N_11451);
or U13529 (N_13529,N_10323,N_11232);
and U13530 (N_13530,N_9852,N_10343);
xnor U13531 (N_13531,N_11341,N_11188);
xor U13532 (N_13532,N_9093,N_9028);
nand U13533 (N_13533,N_10603,N_10940);
xnor U13534 (N_13534,N_10369,N_9436);
or U13535 (N_13535,N_11666,N_11328);
and U13536 (N_13536,N_10882,N_9343);
nand U13537 (N_13537,N_10167,N_11355);
or U13538 (N_13538,N_11766,N_11395);
nand U13539 (N_13539,N_10219,N_10152);
and U13540 (N_13540,N_9046,N_11667);
or U13541 (N_13541,N_9797,N_11239);
or U13542 (N_13542,N_9761,N_10789);
xor U13543 (N_13543,N_10461,N_10841);
nor U13544 (N_13544,N_9508,N_11886);
and U13545 (N_13545,N_9490,N_9694);
nand U13546 (N_13546,N_9085,N_10575);
nor U13547 (N_13547,N_10066,N_10993);
xnor U13548 (N_13548,N_11911,N_10964);
or U13549 (N_13549,N_11065,N_9907);
nor U13550 (N_13550,N_10885,N_10942);
or U13551 (N_13551,N_10502,N_10238);
or U13552 (N_13552,N_10644,N_9876);
nor U13553 (N_13553,N_11016,N_11870);
xor U13554 (N_13554,N_9317,N_10094);
and U13555 (N_13555,N_11711,N_10913);
or U13556 (N_13556,N_9747,N_10596);
nand U13557 (N_13557,N_10448,N_11097);
or U13558 (N_13558,N_10476,N_10980);
or U13559 (N_13559,N_11368,N_10830);
and U13560 (N_13560,N_9334,N_9699);
or U13561 (N_13561,N_10133,N_9419);
xnor U13562 (N_13562,N_11894,N_10701);
nand U13563 (N_13563,N_10834,N_9794);
or U13564 (N_13564,N_9381,N_9218);
xor U13565 (N_13565,N_10153,N_9083);
or U13566 (N_13566,N_9324,N_10246);
or U13567 (N_13567,N_10466,N_11279);
xnor U13568 (N_13568,N_10944,N_10234);
nor U13569 (N_13569,N_11826,N_10119);
xor U13570 (N_13570,N_11059,N_11081);
nand U13571 (N_13571,N_11621,N_9419);
nand U13572 (N_13572,N_10501,N_11961);
xnor U13573 (N_13573,N_10675,N_10247);
or U13574 (N_13574,N_10386,N_10486);
and U13575 (N_13575,N_9788,N_10102);
or U13576 (N_13576,N_11464,N_10475);
xnor U13577 (N_13577,N_10840,N_11963);
or U13578 (N_13578,N_11302,N_9320);
or U13579 (N_13579,N_10491,N_11660);
nor U13580 (N_13580,N_10838,N_11013);
or U13581 (N_13581,N_11596,N_11824);
xnor U13582 (N_13582,N_10491,N_9558);
nor U13583 (N_13583,N_10106,N_9519);
nand U13584 (N_13584,N_9544,N_11484);
or U13585 (N_13585,N_9893,N_10565);
nor U13586 (N_13586,N_11361,N_10332);
nand U13587 (N_13587,N_11200,N_11408);
nor U13588 (N_13588,N_9676,N_10974);
or U13589 (N_13589,N_9456,N_9878);
xor U13590 (N_13590,N_9866,N_10763);
and U13591 (N_13591,N_11367,N_9501);
or U13592 (N_13592,N_10169,N_10916);
nand U13593 (N_13593,N_10337,N_11746);
nand U13594 (N_13594,N_9620,N_10588);
or U13595 (N_13595,N_11577,N_9501);
and U13596 (N_13596,N_10981,N_10166);
and U13597 (N_13597,N_10377,N_10003);
xor U13598 (N_13598,N_11963,N_10376);
nor U13599 (N_13599,N_10198,N_11071);
and U13600 (N_13600,N_9961,N_11187);
xnor U13601 (N_13601,N_11362,N_10174);
nand U13602 (N_13602,N_11377,N_9699);
nand U13603 (N_13603,N_10324,N_10142);
nand U13604 (N_13604,N_9893,N_10109);
nor U13605 (N_13605,N_11261,N_10806);
nor U13606 (N_13606,N_10323,N_11650);
xnor U13607 (N_13607,N_11881,N_11265);
nand U13608 (N_13608,N_11689,N_9259);
nor U13609 (N_13609,N_10729,N_9792);
and U13610 (N_13610,N_11649,N_11062);
nand U13611 (N_13611,N_11703,N_9294);
xnor U13612 (N_13612,N_10661,N_11267);
xnor U13613 (N_13613,N_10090,N_11726);
nand U13614 (N_13614,N_11497,N_10894);
xnor U13615 (N_13615,N_10193,N_10492);
and U13616 (N_13616,N_10820,N_9485);
or U13617 (N_13617,N_9643,N_10321);
or U13618 (N_13618,N_10297,N_11721);
xor U13619 (N_13619,N_11049,N_11638);
nor U13620 (N_13620,N_11197,N_11161);
or U13621 (N_13621,N_11227,N_11321);
nand U13622 (N_13622,N_9887,N_10271);
xor U13623 (N_13623,N_10323,N_11181);
xor U13624 (N_13624,N_11532,N_10862);
nor U13625 (N_13625,N_10754,N_11020);
xnor U13626 (N_13626,N_9997,N_10805);
nand U13627 (N_13627,N_9246,N_11963);
and U13628 (N_13628,N_9906,N_9398);
nand U13629 (N_13629,N_10567,N_9289);
nand U13630 (N_13630,N_9184,N_11303);
nand U13631 (N_13631,N_11319,N_9803);
nand U13632 (N_13632,N_10953,N_11321);
xor U13633 (N_13633,N_9879,N_11591);
xnor U13634 (N_13634,N_11129,N_11952);
nor U13635 (N_13635,N_11373,N_11761);
nand U13636 (N_13636,N_10250,N_9829);
nand U13637 (N_13637,N_11932,N_11204);
and U13638 (N_13638,N_10071,N_10217);
nand U13639 (N_13639,N_10249,N_9540);
or U13640 (N_13640,N_9588,N_10385);
nand U13641 (N_13641,N_9054,N_9929);
nor U13642 (N_13642,N_10901,N_10211);
or U13643 (N_13643,N_10517,N_11883);
xor U13644 (N_13644,N_10122,N_9573);
xor U13645 (N_13645,N_10360,N_9931);
nor U13646 (N_13646,N_9763,N_11341);
or U13647 (N_13647,N_9218,N_10035);
nor U13648 (N_13648,N_11087,N_9970);
xnor U13649 (N_13649,N_9329,N_9895);
and U13650 (N_13650,N_9005,N_9717);
or U13651 (N_13651,N_10195,N_10397);
nand U13652 (N_13652,N_9500,N_11263);
or U13653 (N_13653,N_9209,N_11923);
nor U13654 (N_13654,N_10337,N_11208);
and U13655 (N_13655,N_11106,N_11916);
xnor U13656 (N_13656,N_10617,N_9425);
and U13657 (N_13657,N_9209,N_10076);
and U13658 (N_13658,N_10528,N_10542);
and U13659 (N_13659,N_11531,N_10057);
xnor U13660 (N_13660,N_11049,N_9256);
xor U13661 (N_13661,N_10621,N_11820);
xor U13662 (N_13662,N_10957,N_11670);
nand U13663 (N_13663,N_10768,N_10947);
nor U13664 (N_13664,N_10048,N_9686);
xnor U13665 (N_13665,N_9662,N_9591);
nor U13666 (N_13666,N_11808,N_11464);
and U13667 (N_13667,N_11100,N_9504);
xnor U13668 (N_13668,N_9207,N_10746);
nand U13669 (N_13669,N_11987,N_9527);
and U13670 (N_13670,N_9758,N_10996);
nand U13671 (N_13671,N_10930,N_9114);
nand U13672 (N_13672,N_11987,N_10634);
xnor U13673 (N_13673,N_9427,N_10271);
nor U13674 (N_13674,N_11334,N_10093);
nand U13675 (N_13675,N_9887,N_10468);
or U13676 (N_13676,N_10575,N_11895);
xor U13677 (N_13677,N_9806,N_10628);
nand U13678 (N_13678,N_9102,N_9088);
nand U13679 (N_13679,N_11308,N_9967);
nor U13680 (N_13680,N_9587,N_11960);
nand U13681 (N_13681,N_11317,N_10724);
xnor U13682 (N_13682,N_9688,N_11662);
or U13683 (N_13683,N_11061,N_11342);
and U13684 (N_13684,N_10744,N_9631);
or U13685 (N_13685,N_10010,N_10761);
xor U13686 (N_13686,N_11733,N_11181);
nor U13687 (N_13687,N_10726,N_10956);
nand U13688 (N_13688,N_11673,N_11799);
nand U13689 (N_13689,N_10356,N_9032);
xor U13690 (N_13690,N_10288,N_9113);
nand U13691 (N_13691,N_10005,N_10333);
nor U13692 (N_13692,N_9168,N_10654);
nor U13693 (N_13693,N_9377,N_10775);
nand U13694 (N_13694,N_10853,N_11364);
nor U13695 (N_13695,N_9643,N_10921);
nand U13696 (N_13696,N_9970,N_10533);
and U13697 (N_13697,N_11974,N_9476);
xor U13698 (N_13698,N_9585,N_9210);
xor U13699 (N_13699,N_9866,N_11969);
nor U13700 (N_13700,N_11150,N_9542);
nor U13701 (N_13701,N_11078,N_10208);
nand U13702 (N_13702,N_10504,N_10057);
or U13703 (N_13703,N_11367,N_11360);
or U13704 (N_13704,N_10585,N_11239);
or U13705 (N_13705,N_11716,N_10438);
or U13706 (N_13706,N_10905,N_9774);
nor U13707 (N_13707,N_10182,N_9926);
or U13708 (N_13708,N_9180,N_9332);
and U13709 (N_13709,N_11636,N_11984);
and U13710 (N_13710,N_11462,N_11674);
and U13711 (N_13711,N_11457,N_9334);
nor U13712 (N_13712,N_9047,N_11272);
and U13713 (N_13713,N_9177,N_11390);
or U13714 (N_13714,N_11266,N_9065);
and U13715 (N_13715,N_11471,N_10356);
nand U13716 (N_13716,N_10867,N_11273);
nand U13717 (N_13717,N_11544,N_11446);
and U13718 (N_13718,N_9568,N_11886);
nor U13719 (N_13719,N_10055,N_10149);
xor U13720 (N_13720,N_9323,N_11320);
nand U13721 (N_13721,N_11104,N_10383);
or U13722 (N_13722,N_10690,N_10592);
nand U13723 (N_13723,N_9288,N_10472);
and U13724 (N_13724,N_11475,N_9963);
xnor U13725 (N_13725,N_9582,N_10375);
nand U13726 (N_13726,N_9928,N_9359);
nand U13727 (N_13727,N_11826,N_10313);
and U13728 (N_13728,N_11423,N_11801);
xor U13729 (N_13729,N_11442,N_11845);
nor U13730 (N_13730,N_9447,N_11307);
xnor U13731 (N_13731,N_9234,N_11078);
nand U13732 (N_13732,N_10731,N_9420);
or U13733 (N_13733,N_11621,N_9076);
xor U13734 (N_13734,N_11872,N_11539);
or U13735 (N_13735,N_10373,N_11843);
or U13736 (N_13736,N_9119,N_11409);
and U13737 (N_13737,N_10614,N_10728);
and U13738 (N_13738,N_10292,N_10938);
nand U13739 (N_13739,N_10227,N_9568);
and U13740 (N_13740,N_9965,N_9007);
nor U13741 (N_13741,N_11323,N_10750);
nor U13742 (N_13742,N_11369,N_11247);
and U13743 (N_13743,N_10298,N_11923);
and U13744 (N_13744,N_10477,N_10752);
nand U13745 (N_13745,N_9699,N_10133);
or U13746 (N_13746,N_11940,N_10174);
or U13747 (N_13747,N_10179,N_11332);
and U13748 (N_13748,N_11391,N_9444);
xor U13749 (N_13749,N_10181,N_10487);
or U13750 (N_13750,N_9534,N_10013);
or U13751 (N_13751,N_9850,N_11648);
xor U13752 (N_13752,N_11355,N_10390);
nand U13753 (N_13753,N_11948,N_10253);
nor U13754 (N_13754,N_9651,N_10834);
or U13755 (N_13755,N_9696,N_9752);
xnor U13756 (N_13756,N_9703,N_10251);
and U13757 (N_13757,N_11056,N_11176);
and U13758 (N_13758,N_10207,N_10447);
xor U13759 (N_13759,N_11611,N_9984);
nor U13760 (N_13760,N_11602,N_11547);
or U13761 (N_13761,N_9337,N_10288);
xnor U13762 (N_13762,N_10393,N_9965);
nand U13763 (N_13763,N_11073,N_10754);
nor U13764 (N_13764,N_9636,N_11617);
or U13765 (N_13765,N_11348,N_11155);
or U13766 (N_13766,N_11565,N_11230);
nor U13767 (N_13767,N_10342,N_9237);
nand U13768 (N_13768,N_9552,N_9513);
nand U13769 (N_13769,N_9304,N_11211);
nand U13770 (N_13770,N_10847,N_10874);
nor U13771 (N_13771,N_9283,N_11887);
nor U13772 (N_13772,N_10342,N_11188);
and U13773 (N_13773,N_11791,N_10691);
nand U13774 (N_13774,N_11587,N_10603);
or U13775 (N_13775,N_11307,N_9041);
or U13776 (N_13776,N_11392,N_10925);
nor U13777 (N_13777,N_10554,N_9225);
xor U13778 (N_13778,N_11407,N_11535);
and U13779 (N_13779,N_10454,N_11523);
or U13780 (N_13780,N_10831,N_10880);
or U13781 (N_13781,N_11226,N_11077);
or U13782 (N_13782,N_11949,N_9488);
xnor U13783 (N_13783,N_10862,N_11150);
and U13784 (N_13784,N_11084,N_9390);
nand U13785 (N_13785,N_10705,N_11426);
nor U13786 (N_13786,N_9076,N_10459);
or U13787 (N_13787,N_10586,N_9890);
or U13788 (N_13788,N_11940,N_9128);
or U13789 (N_13789,N_9658,N_9318);
and U13790 (N_13790,N_10901,N_11795);
nor U13791 (N_13791,N_10334,N_11689);
or U13792 (N_13792,N_11830,N_9126);
and U13793 (N_13793,N_11259,N_11408);
and U13794 (N_13794,N_10906,N_9280);
or U13795 (N_13795,N_10273,N_9824);
and U13796 (N_13796,N_10779,N_11996);
nor U13797 (N_13797,N_10558,N_10530);
nor U13798 (N_13798,N_10575,N_9444);
xor U13799 (N_13799,N_10666,N_9459);
nor U13800 (N_13800,N_11491,N_11251);
or U13801 (N_13801,N_10804,N_11507);
nor U13802 (N_13802,N_11603,N_11824);
or U13803 (N_13803,N_10326,N_9195);
and U13804 (N_13804,N_10127,N_9204);
and U13805 (N_13805,N_10564,N_11041);
and U13806 (N_13806,N_9427,N_11670);
and U13807 (N_13807,N_11330,N_10357);
or U13808 (N_13808,N_9434,N_9263);
and U13809 (N_13809,N_11183,N_10175);
nor U13810 (N_13810,N_9044,N_11030);
and U13811 (N_13811,N_11050,N_11438);
nor U13812 (N_13812,N_9288,N_11479);
and U13813 (N_13813,N_10768,N_9264);
and U13814 (N_13814,N_11092,N_11509);
xor U13815 (N_13815,N_9293,N_9665);
and U13816 (N_13816,N_10424,N_9966);
nor U13817 (N_13817,N_9575,N_11668);
xor U13818 (N_13818,N_10722,N_11443);
xor U13819 (N_13819,N_11797,N_9098);
xor U13820 (N_13820,N_11506,N_9527);
and U13821 (N_13821,N_11997,N_9046);
nand U13822 (N_13822,N_9056,N_10113);
xnor U13823 (N_13823,N_9568,N_10446);
nand U13824 (N_13824,N_10669,N_9165);
nand U13825 (N_13825,N_11060,N_9141);
nand U13826 (N_13826,N_11489,N_10298);
nand U13827 (N_13827,N_11027,N_11841);
nor U13828 (N_13828,N_9850,N_9243);
nand U13829 (N_13829,N_10986,N_9400);
and U13830 (N_13830,N_10379,N_10049);
xor U13831 (N_13831,N_9447,N_11162);
xor U13832 (N_13832,N_10602,N_10169);
and U13833 (N_13833,N_10000,N_9088);
and U13834 (N_13834,N_9421,N_11700);
xor U13835 (N_13835,N_11434,N_11531);
nor U13836 (N_13836,N_9580,N_10774);
nand U13837 (N_13837,N_11057,N_10657);
and U13838 (N_13838,N_9778,N_9506);
nor U13839 (N_13839,N_9738,N_10406);
xor U13840 (N_13840,N_10644,N_9602);
nand U13841 (N_13841,N_10112,N_9840);
nor U13842 (N_13842,N_10670,N_9246);
nor U13843 (N_13843,N_10748,N_11912);
nor U13844 (N_13844,N_11900,N_11325);
or U13845 (N_13845,N_9901,N_11845);
and U13846 (N_13846,N_10294,N_9948);
nor U13847 (N_13847,N_10195,N_11165);
nand U13848 (N_13848,N_9424,N_11066);
nand U13849 (N_13849,N_11984,N_11532);
and U13850 (N_13850,N_10546,N_10580);
xor U13851 (N_13851,N_10484,N_10823);
and U13852 (N_13852,N_10757,N_10851);
nand U13853 (N_13853,N_9590,N_9847);
or U13854 (N_13854,N_10244,N_11433);
xnor U13855 (N_13855,N_11203,N_11285);
nor U13856 (N_13856,N_9425,N_10146);
nor U13857 (N_13857,N_11494,N_11981);
and U13858 (N_13858,N_11679,N_11180);
nand U13859 (N_13859,N_10968,N_11092);
xor U13860 (N_13860,N_9308,N_10109);
nand U13861 (N_13861,N_11456,N_10754);
nor U13862 (N_13862,N_11702,N_11842);
xor U13863 (N_13863,N_11150,N_10866);
and U13864 (N_13864,N_9776,N_11576);
nor U13865 (N_13865,N_11793,N_9184);
and U13866 (N_13866,N_11418,N_10012);
and U13867 (N_13867,N_10301,N_11086);
nand U13868 (N_13868,N_11324,N_9984);
and U13869 (N_13869,N_11182,N_10819);
or U13870 (N_13870,N_11677,N_11752);
nor U13871 (N_13871,N_11314,N_11102);
xor U13872 (N_13872,N_10370,N_11335);
or U13873 (N_13873,N_9617,N_10511);
xnor U13874 (N_13874,N_9810,N_9222);
or U13875 (N_13875,N_10259,N_11800);
or U13876 (N_13876,N_11974,N_9407);
or U13877 (N_13877,N_10025,N_11306);
nand U13878 (N_13878,N_9570,N_11964);
xor U13879 (N_13879,N_11924,N_10985);
xnor U13880 (N_13880,N_9333,N_10020);
nor U13881 (N_13881,N_11872,N_9615);
xnor U13882 (N_13882,N_10209,N_10145);
or U13883 (N_13883,N_11342,N_10453);
nor U13884 (N_13884,N_10600,N_10137);
or U13885 (N_13885,N_10995,N_9432);
and U13886 (N_13886,N_9494,N_9074);
and U13887 (N_13887,N_9418,N_9078);
nand U13888 (N_13888,N_10608,N_9769);
nor U13889 (N_13889,N_10763,N_11101);
or U13890 (N_13890,N_9296,N_10844);
xor U13891 (N_13891,N_11203,N_10016);
nor U13892 (N_13892,N_10741,N_10450);
nor U13893 (N_13893,N_9772,N_10061);
and U13894 (N_13894,N_11272,N_9700);
or U13895 (N_13895,N_9075,N_9924);
nand U13896 (N_13896,N_10367,N_11380);
and U13897 (N_13897,N_10656,N_10170);
xor U13898 (N_13898,N_11217,N_10601);
nor U13899 (N_13899,N_11155,N_10077);
xor U13900 (N_13900,N_10203,N_11683);
nor U13901 (N_13901,N_9157,N_10970);
nor U13902 (N_13902,N_10006,N_9846);
nor U13903 (N_13903,N_9580,N_9548);
or U13904 (N_13904,N_9234,N_11025);
or U13905 (N_13905,N_10552,N_10048);
or U13906 (N_13906,N_9766,N_10848);
nor U13907 (N_13907,N_10062,N_9479);
nand U13908 (N_13908,N_10903,N_9916);
nand U13909 (N_13909,N_10619,N_11072);
nor U13910 (N_13910,N_9015,N_9856);
or U13911 (N_13911,N_10436,N_11122);
and U13912 (N_13912,N_11261,N_9266);
or U13913 (N_13913,N_11856,N_9361);
nand U13914 (N_13914,N_10476,N_9112);
nand U13915 (N_13915,N_9507,N_10024);
nor U13916 (N_13916,N_9865,N_9586);
nor U13917 (N_13917,N_10308,N_9654);
xnor U13918 (N_13918,N_9845,N_11513);
nor U13919 (N_13919,N_9513,N_11889);
and U13920 (N_13920,N_11245,N_10834);
nand U13921 (N_13921,N_11270,N_10922);
or U13922 (N_13922,N_11265,N_11343);
and U13923 (N_13923,N_9104,N_10341);
and U13924 (N_13924,N_11194,N_9874);
or U13925 (N_13925,N_10417,N_10051);
and U13926 (N_13926,N_9066,N_10485);
and U13927 (N_13927,N_10051,N_9781);
nand U13928 (N_13928,N_9547,N_11923);
or U13929 (N_13929,N_10476,N_9051);
nor U13930 (N_13930,N_11608,N_9441);
nor U13931 (N_13931,N_9171,N_9058);
and U13932 (N_13932,N_11092,N_10469);
nor U13933 (N_13933,N_9269,N_11320);
or U13934 (N_13934,N_11819,N_11118);
nand U13935 (N_13935,N_11365,N_9304);
nand U13936 (N_13936,N_10160,N_10848);
or U13937 (N_13937,N_10404,N_10745);
xor U13938 (N_13938,N_11191,N_9664);
xor U13939 (N_13939,N_9153,N_11109);
xor U13940 (N_13940,N_10094,N_11633);
nor U13941 (N_13941,N_10075,N_10549);
xnor U13942 (N_13942,N_11098,N_11265);
nor U13943 (N_13943,N_11302,N_11510);
or U13944 (N_13944,N_11426,N_10047);
and U13945 (N_13945,N_10936,N_11260);
nand U13946 (N_13946,N_10976,N_10534);
xor U13947 (N_13947,N_11451,N_9116);
xnor U13948 (N_13948,N_9468,N_9728);
nor U13949 (N_13949,N_9467,N_11060);
nand U13950 (N_13950,N_9426,N_10026);
nand U13951 (N_13951,N_10274,N_9315);
or U13952 (N_13952,N_11145,N_11931);
nor U13953 (N_13953,N_11869,N_10215);
and U13954 (N_13954,N_9948,N_10072);
nand U13955 (N_13955,N_9371,N_11337);
and U13956 (N_13956,N_11278,N_9425);
and U13957 (N_13957,N_11842,N_10433);
nand U13958 (N_13958,N_11381,N_11862);
and U13959 (N_13959,N_10781,N_10187);
nor U13960 (N_13960,N_11091,N_10639);
or U13961 (N_13961,N_9448,N_11446);
or U13962 (N_13962,N_9323,N_11337);
xnor U13963 (N_13963,N_9136,N_9075);
nor U13964 (N_13964,N_9694,N_9144);
nor U13965 (N_13965,N_10395,N_11989);
or U13966 (N_13966,N_9197,N_11281);
or U13967 (N_13967,N_9076,N_10421);
nor U13968 (N_13968,N_11319,N_11593);
xor U13969 (N_13969,N_11527,N_10579);
and U13970 (N_13970,N_10843,N_9958);
or U13971 (N_13971,N_10411,N_11246);
xnor U13972 (N_13972,N_9589,N_9422);
xnor U13973 (N_13973,N_11166,N_9884);
and U13974 (N_13974,N_9381,N_9741);
xnor U13975 (N_13975,N_9200,N_9330);
nor U13976 (N_13976,N_9280,N_9102);
xor U13977 (N_13977,N_9775,N_10306);
or U13978 (N_13978,N_10866,N_10683);
nor U13979 (N_13979,N_9307,N_10205);
nor U13980 (N_13980,N_10996,N_9641);
and U13981 (N_13981,N_10202,N_10184);
nor U13982 (N_13982,N_10236,N_11351);
or U13983 (N_13983,N_10940,N_9122);
or U13984 (N_13984,N_10916,N_11010);
or U13985 (N_13985,N_9406,N_10342);
nand U13986 (N_13986,N_11313,N_9832);
nor U13987 (N_13987,N_9556,N_9987);
xor U13988 (N_13988,N_11878,N_9667);
xnor U13989 (N_13989,N_10583,N_11584);
nor U13990 (N_13990,N_9790,N_9588);
or U13991 (N_13991,N_11172,N_10891);
or U13992 (N_13992,N_10918,N_11985);
nor U13993 (N_13993,N_9343,N_10561);
or U13994 (N_13994,N_10541,N_11705);
or U13995 (N_13995,N_10722,N_11533);
and U13996 (N_13996,N_9912,N_10195);
nor U13997 (N_13997,N_11674,N_9917);
nand U13998 (N_13998,N_11320,N_11584);
or U13999 (N_13999,N_9360,N_9964);
or U14000 (N_14000,N_11963,N_10025);
and U14001 (N_14001,N_9590,N_11135);
and U14002 (N_14002,N_9176,N_9737);
and U14003 (N_14003,N_10176,N_10039);
xor U14004 (N_14004,N_9881,N_11167);
nand U14005 (N_14005,N_9940,N_10123);
nor U14006 (N_14006,N_10400,N_10595);
and U14007 (N_14007,N_10780,N_11015);
or U14008 (N_14008,N_10884,N_9838);
xor U14009 (N_14009,N_10392,N_10813);
nand U14010 (N_14010,N_11263,N_11151);
and U14011 (N_14011,N_11338,N_11660);
and U14012 (N_14012,N_9375,N_9961);
or U14013 (N_14013,N_9699,N_11679);
nor U14014 (N_14014,N_10246,N_9795);
xnor U14015 (N_14015,N_11582,N_9274);
xnor U14016 (N_14016,N_9697,N_9979);
or U14017 (N_14017,N_10040,N_9941);
xnor U14018 (N_14018,N_11097,N_10532);
and U14019 (N_14019,N_9084,N_11018);
and U14020 (N_14020,N_11888,N_10914);
nand U14021 (N_14021,N_9163,N_11600);
nand U14022 (N_14022,N_10737,N_9382);
xor U14023 (N_14023,N_9317,N_9761);
xor U14024 (N_14024,N_10705,N_10121);
nand U14025 (N_14025,N_11132,N_11434);
or U14026 (N_14026,N_10151,N_11883);
xor U14027 (N_14027,N_11228,N_9503);
nor U14028 (N_14028,N_10184,N_11263);
nand U14029 (N_14029,N_10767,N_10055);
and U14030 (N_14030,N_11214,N_11916);
or U14031 (N_14031,N_11668,N_11317);
nor U14032 (N_14032,N_11678,N_11436);
and U14033 (N_14033,N_10378,N_10535);
and U14034 (N_14034,N_9904,N_10923);
nand U14035 (N_14035,N_9315,N_10678);
or U14036 (N_14036,N_11454,N_11013);
nand U14037 (N_14037,N_9386,N_11579);
or U14038 (N_14038,N_10349,N_11702);
or U14039 (N_14039,N_11465,N_11095);
or U14040 (N_14040,N_9131,N_10793);
nor U14041 (N_14041,N_11633,N_11654);
xnor U14042 (N_14042,N_9360,N_10483);
xor U14043 (N_14043,N_10401,N_9495);
nand U14044 (N_14044,N_9885,N_10804);
and U14045 (N_14045,N_11855,N_11754);
and U14046 (N_14046,N_11640,N_10611);
nor U14047 (N_14047,N_11341,N_11403);
nor U14048 (N_14048,N_11269,N_11821);
or U14049 (N_14049,N_10238,N_9252);
and U14050 (N_14050,N_9017,N_10795);
xnor U14051 (N_14051,N_11052,N_10806);
or U14052 (N_14052,N_9611,N_10840);
xor U14053 (N_14053,N_10050,N_9157);
nor U14054 (N_14054,N_10584,N_9899);
and U14055 (N_14055,N_11961,N_11957);
nor U14056 (N_14056,N_10268,N_10648);
and U14057 (N_14057,N_9124,N_10429);
xor U14058 (N_14058,N_10063,N_10860);
and U14059 (N_14059,N_11491,N_10585);
nand U14060 (N_14060,N_10029,N_11877);
xor U14061 (N_14061,N_11083,N_9695);
xor U14062 (N_14062,N_11476,N_9113);
or U14063 (N_14063,N_10245,N_9321);
nor U14064 (N_14064,N_11954,N_9883);
nand U14065 (N_14065,N_11275,N_11519);
or U14066 (N_14066,N_10616,N_11772);
nor U14067 (N_14067,N_11161,N_11569);
nor U14068 (N_14068,N_11430,N_9174);
nand U14069 (N_14069,N_10480,N_9711);
nand U14070 (N_14070,N_10332,N_11918);
and U14071 (N_14071,N_9866,N_10558);
or U14072 (N_14072,N_10521,N_11544);
or U14073 (N_14073,N_9383,N_9999);
nand U14074 (N_14074,N_9315,N_11345);
nand U14075 (N_14075,N_9354,N_9159);
or U14076 (N_14076,N_10466,N_11805);
and U14077 (N_14077,N_9031,N_11362);
or U14078 (N_14078,N_9611,N_9313);
nand U14079 (N_14079,N_11596,N_10968);
nor U14080 (N_14080,N_11881,N_11638);
and U14081 (N_14081,N_9221,N_10899);
and U14082 (N_14082,N_9456,N_10331);
xnor U14083 (N_14083,N_9436,N_11420);
nand U14084 (N_14084,N_9942,N_9102);
xor U14085 (N_14085,N_10897,N_11754);
nor U14086 (N_14086,N_9133,N_11566);
nor U14087 (N_14087,N_10022,N_10749);
nand U14088 (N_14088,N_11874,N_9616);
or U14089 (N_14089,N_9756,N_10995);
or U14090 (N_14090,N_9179,N_10128);
or U14091 (N_14091,N_10899,N_10145);
nand U14092 (N_14092,N_11473,N_9795);
or U14093 (N_14093,N_11982,N_9954);
nor U14094 (N_14094,N_11818,N_11426);
xor U14095 (N_14095,N_9234,N_11833);
nand U14096 (N_14096,N_9754,N_10799);
nand U14097 (N_14097,N_9303,N_9952);
nand U14098 (N_14098,N_9850,N_9631);
and U14099 (N_14099,N_9917,N_10525);
and U14100 (N_14100,N_9558,N_10399);
nand U14101 (N_14101,N_10651,N_11001);
or U14102 (N_14102,N_10660,N_11712);
nor U14103 (N_14103,N_10712,N_10287);
or U14104 (N_14104,N_9757,N_11457);
xnor U14105 (N_14105,N_9073,N_10065);
or U14106 (N_14106,N_11061,N_11170);
nand U14107 (N_14107,N_9918,N_10231);
nor U14108 (N_14108,N_11959,N_9663);
or U14109 (N_14109,N_11696,N_10373);
and U14110 (N_14110,N_10219,N_10979);
or U14111 (N_14111,N_9203,N_10407);
nand U14112 (N_14112,N_9075,N_11280);
or U14113 (N_14113,N_11184,N_9944);
and U14114 (N_14114,N_9916,N_11100);
xor U14115 (N_14115,N_10115,N_11036);
nor U14116 (N_14116,N_9921,N_11498);
and U14117 (N_14117,N_10075,N_11713);
and U14118 (N_14118,N_10917,N_11965);
or U14119 (N_14119,N_11432,N_10212);
nand U14120 (N_14120,N_10241,N_10578);
nand U14121 (N_14121,N_9285,N_10339);
or U14122 (N_14122,N_11190,N_11496);
and U14123 (N_14123,N_11226,N_9945);
xor U14124 (N_14124,N_9489,N_9402);
nor U14125 (N_14125,N_11837,N_11920);
nand U14126 (N_14126,N_10301,N_11355);
nand U14127 (N_14127,N_10376,N_11606);
nor U14128 (N_14128,N_11492,N_11942);
nand U14129 (N_14129,N_11825,N_9551);
nor U14130 (N_14130,N_9940,N_9527);
nand U14131 (N_14131,N_11254,N_9485);
and U14132 (N_14132,N_9305,N_9333);
or U14133 (N_14133,N_11913,N_9071);
nand U14134 (N_14134,N_9419,N_10181);
nand U14135 (N_14135,N_9758,N_10722);
xnor U14136 (N_14136,N_9971,N_10084);
nand U14137 (N_14137,N_9549,N_9628);
nor U14138 (N_14138,N_10546,N_9047);
nand U14139 (N_14139,N_9089,N_9137);
nand U14140 (N_14140,N_11691,N_10543);
nand U14141 (N_14141,N_9587,N_11936);
xnor U14142 (N_14142,N_11285,N_10053);
and U14143 (N_14143,N_9890,N_10226);
and U14144 (N_14144,N_9017,N_11981);
or U14145 (N_14145,N_10261,N_11003);
or U14146 (N_14146,N_10079,N_10817);
and U14147 (N_14147,N_11299,N_10136);
and U14148 (N_14148,N_10864,N_10487);
nand U14149 (N_14149,N_11660,N_10065);
and U14150 (N_14150,N_10998,N_10008);
or U14151 (N_14151,N_10347,N_10227);
nor U14152 (N_14152,N_11857,N_9639);
xor U14153 (N_14153,N_10108,N_10724);
nand U14154 (N_14154,N_11463,N_11457);
nor U14155 (N_14155,N_11935,N_9622);
or U14156 (N_14156,N_9467,N_9929);
nor U14157 (N_14157,N_9499,N_9427);
xor U14158 (N_14158,N_10899,N_10322);
xor U14159 (N_14159,N_9030,N_10699);
and U14160 (N_14160,N_9601,N_10292);
and U14161 (N_14161,N_10384,N_9362);
xnor U14162 (N_14162,N_10342,N_11310);
nor U14163 (N_14163,N_11407,N_9802);
nor U14164 (N_14164,N_10724,N_9085);
nand U14165 (N_14165,N_9770,N_9166);
xor U14166 (N_14166,N_10844,N_10498);
nand U14167 (N_14167,N_10747,N_9090);
nor U14168 (N_14168,N_10305,N_9536);
nor U14169 (N_14169,N_11171,N_9653);
nor U14170 (N_14170,N_11831,N_10161);
or U14171 (N_14171,N_10368,N_9110);
nand U14172 (N_14172,N_9031,N_11471);
nand U14173 (N_14173,N_10246,N_11074);
xor U14174 (N_14174,N_11699,N_11929);
nand U14175 (N_14175,N_11327,N_9915);
and U14176 (N_14176,N_9556,N_9109);
xor U14177 (N_14177,N_9167,N_9233);
or U14178 (N_14178,N_10950,N_11343);
xor U14179 (N_14179,N_11750,N_10169);
nand U14180 (N_14180,N_10981,N_11914);
or U14181 (N_14181,N_9958,N_9333);
and U14182 (N_14182,N_10993,N_11207);
nor U14183 (N_14183,N_11439,N_11502);
nand U14184 (N_14184,N_10127,N_9422);
and U14185 (N_14185,N_11895,N_10107);
nand U14186 (N_14186,N_9568,N_11720);
nor U14187 (N_14187,N_9873,N_11988);
and U14188 (N_14188,N_9759,N_11155);
nor U14189 (N_14189,N_10281,N_9850);
nand U14190 (N_14190,N_10516,N_10252);
xor U14191 (N_14191,N_11836,N_11363);
nor U14192 (N_14192,N_9978,N_10773);
nand U14193 (N_14193,N_11096,N_10913);
or U14194 (N_14194,N_9741,N_10319);
nor U14195 (N_14195,N_9953,N_9053);
and U14196 (N_14196,N_11389,N_9039);
nor U14197 (N_14197,N_11599,N_10828);
nor U14198 (N_14198,N_10345,N_9123);
nand U14199 (N_14199,N_9058,N_10121);
nand U14200 (N_14200,N_10989,N_10103);
and U14201 (N_14201,N_11473,N_11416);
or U14202 (N_14202,N_11541,N_10822);
xnor U14203 (N_14203,N_11801,N_10353);
nor U14204 (N_14204,N_9500,N_11273);
or U14205 (N_14205,N_9226,N_10106);
and U14206 (N_14206,N_9752,N_11835);
xnor U14207 (N_14207,N_10585,N_10843);
nor U14208 (N_14208,N_9210,N_10278);
nor U14209 (N_14209,N_9366,N_11238);
nor U14210 (N_14210,N_9312,N_9358);
xor U14211 (N_14211,N_11703,N_11050);
nand U14212 (N_14212,N_11933,N_9759);
nand U14213 (N_14213,N_9112,N_9330);
nor U14214 (N_14214,N_10948,N_11415);
and U14215 (N_14215,N_9069,N_9954);
or U14216 (N_14216,N_9294,N_10409);
nor U14217 (N_14217,N_10822,N_9694);
nor U14218 (N_14218,N_9672,N_10191);
nor U14219 (N_14219,N_10208,N_11436);
or U14220 (N_14220,N_11459,N_11650);
or U14221 (N_14221,N_11094,N_9979);
or U14222 (N_14222,N_11106,N_11682);
and U14223 (N_14223,N_9949,N_11423);
xor U14224 (N_14224,N_10118,N_10031);
nand U14225 (N_14225,N_10745,N_9205);
or U14226 (N_14226,N_9843,N_10525);
or U14227 (N_14227,N_9400,N_10443);
nand U14228 (N_14228,N_9607,N_10154);
nor U14229 (N_14229,N_11230,N_10290);
or U14230 (N_14230,N_10768,N_11130);
or U14231 (N_14231,N_11053,N_11567);
or U14232 (N_14232,N_10813,N_10792);
nand U14233 (N_14233,N_9716,N_10383);
and U14234 (N_14234,N_10905,N_10443);
or U14235 (N_14235,N_11749,N_10248);
nor U14236 (N_14236,N_10766,N_11169);
or U14237 (N_14237,N_9664,N_11409);
nand U14238 (N_14238,N_9027,N_10781);
xor U14239 (N_14239,N_9332,N_11693);
or U14240 (N_14240,N_10847,N_11092);
nand U14241 (N_14241,N_10419,N_10902);
or U14242 (N_14242,N_9346,N_11786);
nand U14243 (N_14243,N_11352,N_10689);
and U14244 (N_14244,N_10301,N_9611);
nand U14245 (N_14245,N_10068,N_10867);
nand U14246 (N_14246,N_11483,N_11778);
nor U14247 (N_14247,N_10197,N_11739);
nor U14248 (N_14248,N_11421,N_9784);
and U14249 (N_14249,N_11101,N_10532);
nand U14250 (N_14250,N_9798,N_11463);
nor U14251 (N_14251,N_9387,N_10215);
nand U14252 (N_14252,N_9369,N_9862);
nand U14253 (N_14253,N_11600,N_10029);
nor U14254 (N_14254,N_9394,N_9547);
or U14255 (N_14255,N_10211,N_11261);
and U14256 (N_14256,N_9098,N_10980);
xor U14257 (N_14257,N_9180,N_9598);
nor U14258 (N_14258,N_11917,N_10892);
nor U14259 (N_14259,N_11853,N_11193);
xnor U14260 (N_14260,N_9772,N_10892);
and U14261 (N_14261,N_10320,N_10766);
nand U14262 (N_14262,N_11311,N_10053);
nand U14263 (N_14263,N_9917,N_9849);
xnor U14264 (N_14264,N_11084,N_9515);
and U14265 (N_14265,N_11257,N_11158);
nand U14266 (N_14266,N_9050,N_10367);
nor U14267 (N_14267,N_10560,N_9968);
nor U14268 (N_14268,N_9398,N_9831);
and U14269 (N_14269,N_9083,N_9562);
and U14270 (N_14270,N_11098,N_11116);
xnor U14271 (N_14271,N_10577,N_9445);
nor U14272 (N_14272,N_10496,N_9670);
nor U14273 (N_14273,N_9778,N_11887);
xor U14274 (N_14274,N_9595,N_9487);
nand U14275 (N_14275,N_11515,N_11755);
and U14276 (N_14276,N_11384,N_9949);
and U14277 (N_14277,N_10817,N_11578);
or U14278 (N_14278,N_9785,N_11142);
xnor U14279 (N_14279,N_10565,N_10048);
or U14280 (N_14280,N_9643,N_9249);
and U14281 (N_14281,N_11128,N_11597);
xor U14282 (N_14282,N_9961,N_10401);
xor U14283 (N_14283,N_9500,N_10814);
nand U14284 (N_14284,N_9461,N_10766);
nand U14285 (N_14285,N_10468,N_10092);
and U14286 (N_14286,N_10879,N_11869);
nand U14287 (N_14287,N_10405,N_11997);
nor U14288 (N_14288,N_10867,N_11253);
nand U14289 (N_14289,N_11937,N_9571);
xor U14290 (N_14290,N_9292,N_10363);
nor U14291 (N_14291,N_11144,N_10582);
and U14292 (N_14292,N_10029,N_11634);
and U14293 (N_14293,N_11363,N_11755);
and U14294 (N_14294,N_9839,N_9190);
or U14295 (N_14295,N_9187,N_9925);
or U14296 (N_14296,N_10667,N_11314);
nand U14297 (N_14297,N_9102,N_10045);
nand U14298 (N_14298,N_11954,N_10563);
and U14299 (N_14299,N_11784,N_11242);
and U14300 (N_14300,N_10493,N_11791);
nor U14301 (N_14301,N_11613,N_10170);
and U14302 (N_14302,N_10902,N_11987);
and U14303 (N_14303,N_10320,N_9173);
nor U14304 (N_14304,N_10752,N_11921);
or U14305 (N_14305,N_11011,N_11288);
or U14306 (N_14306,N_10851,N_9381);
nand U14307 (N_14307,N_9755,N_10277);
xor U14308 (N_14308,N_9273,N_10182);
or U14309 (N_14309,N_10819,N_9861);
xnor U14310 (N_14310,N_10531,N_9063);
xor U14311 (N_14311,N_10395,N_9748);
nor U14312 (N_14312,N_11864,N_10189);
or U14313 (N_14313,N_11049,N_10520);
xnor U14314 (N_14314,N_11711,N_10413);
or U14315 (N_14315,N_10326,N_10604);
nand U14316 (N_14316,N_9169,N_11008);
xnor U14317 (N_14317,N_10856,N_9659);
nand U14318 (N_14318,N_11446,N_11315);
or U14319 (N_14319,N_11983,N_11080);
and U14320 (N_14320,N_11777,N_9866);
xnor U14321 (N_14321,N_11046,N_10218);
xor U14322 (N_14322,N_11997,N_9422);
nor U14323 (N_14323,N_9336,N_9537);
or U14324 (N_14324,N_11186,N_10973);
and U14325 (N_14325,N_10974,N_9580);
nand U14326 (N_14326,N_9819,N_9301);
nand U14327 (N_14327,N_9699,N_11899);
nand U14328 (N_14328,N_10156,N_11217);
or U14329 (N_14329,N_11169,N_10620);
nand U14330 (N_14330,N_10285,N_9178);
or U14331 (N_14331,N_10509,N_10618);
and U14332 (N_14332,N_10708,N_11219);
xnor U14333 (N_14333,N_9541,N_10019);
nand U14334 (N_14334,N_10159,N_10991);
xnor U14335 (N_14335,N_10084,N_11596);
xor U14336 (N_14336,N_10114,N_11958);
xor U14337 (N_14337,N_9259,N_9993);
nor U14338 (N_14338,N_9936,N_9981);
nand U14339 (N_14339,N_10627,N_10140);
nor U14340 (N_14340,N_10192,N_10824);
and U14341 (N_14341,N_9821,N_9047);
nor U14342 (N_14342,N_10653,N_11082);
nand U14343 (N_14343,N_10927,N_10372);
or U14344 (N_14344,N_11213,N_10044);
and U14345 (N_14345,N_9230,N_10989);
or U14346 (N_14346,N_10270,N_11164);
or U14347 (N_14347,N_11110,N_9412);
xor U14348 (N_14348,N_9029,N_10211);
and U14349 (N_14349,N_10948,N_11071);
xor U14350 (N_14350,N_10039,N_10961);
or U14351 (N_14351,N_10896,N_11522);
or U14352 (N_14352,N_9250,N_9682);
and U14353 (N_14353,N_11289,N_10451);
and U14354 (N_14354,N_11603,N_11795);
nand U14355 (N_14355,N_11722,N_10665);
and U14356 (N_14356,N_9036,N_11510);
nand U14357 (N_14357,N_11149,N_9135);
nor U14358 (N_14358,N_10113,N_10643);
nand U14359 (N_14359,N_11451,N_9505);
or U14360 (N_14360,N_10372,N_10558);
nand U14361 (N_14361,N_10029,N_11976);
nand U14362 (N_14362,N_9906,N_10544);
and U14363 (N_14363,N_11860,N_9210);
or U14364 (N_14364,N_10124,N_9768);
or U14365 (N_14365,N_11305,N_11446);
nand U14366 (N_14366,N_11326,N_10244);
nand U14367 (N_14367,N_9717,N_9589);
nand U14368 (N_14368,N_9396,N_9310);
and U14369 (N_14369,N_9902,N_9480);
xnor U14370 (N_14370,N_11742,N_9324);
and U14371 (N_14371,N_11422,N_11977);
and U14372 (N_14372,N_10998,N_9296);
xor U14373 (N_14373,N_9165,N_10094);
and U14374 (N_14374,N_10890,N_9275);
nand U14375 (N_14375,N_9024,N_11282);
and U14376 (N_14376,N_10962,N_9092);
xor U14377 (N_14377,N_9326,N_10616);
and U14378 (N_14378,N_9543,N_11210);
nand U14379 (N_14379,N_9304,N_10035);
nand U14380 (N_14380,N_10660,N_11293);
or U14381 (N_14381,N_10425,N_9449);
xnor U14382 (N_14382,N_9080,N_11612);
xnor U14383 (N_14383,N_11659,N_11852);
nand U14384 (N_14384,N_11158,N_9164);
nor U14385 (N_14385,N_9351,N_9690);
nand U14386 (N_14386,N_10896,N_11820);
nand U14387 (N_14387,N_10484,N_10473);
nor U14388 (N_14388,N_10816,N_9546);
nand U14389 (N_14389,N_11564,N_9722);
nand U14390 (N_14390,N_10970,N_9667);
and U14391 (N_14391,N_11462,N_9321);
or U14392 (N_14392,N_11573,N_11827);
nor U14393 (N_14393,N_9428,N_11148);
or U14394 (N_14394,N_10295,N_9478);
nand U14395 (N_14395,N_10302,N_10765);
nor U14396 (N_14396,N_11473,N_11345);
and U14397 (N_14397,N_10791,N_9536);
nor U14398 (N_14398,N_9678,N_11620);
nor U14399 (N_14399,N_11457,N_11378);
xor U14400 (N_14400,N_10409,N_10673);
xor U14401 (N_14401,N_11064,N_10716);
and U14402 (N_14402,N_11082,N_9150);
nand U14403 (N_14403,N_9040,N_11232);
xnor U14404 (N_14404,N_11860,N_9466);
or U14405 (N_14405,N_11260,N_10880);
nor U14406 (N_14406,N_9743,N_10967);
nand U14407 (N_14407,N_11100,N_11474);
and U14408 (N_14408,N_11550,N_9050);
xnor U14409 (N_14409,N_10904,N_11319);
or U14410 (N_14410,N_11936,N_9732);
or U14411 (N_14411,N_11539,N_9236);
nand U14412 (N_14412,N_10529,N_10070);
nand U14413 (N_14413,N_11895,N_9296);
xnor U14414 (N_14414,N_9140,N_10226);
and U14415 (N_14415,N_10612,N_11810);
and U14416 (N_14416,N_10611,N_10673);
nor U14417 (N_14417,N_11743,N_11909);
nand U14418 (N_14418,N_11391,N_9918);
nor U14419 (N_14419,N_11358,N_10950);
or U14420 (N_14420,N_9633,N_9915);
or U14421 (N_14421,N_9935,N_10705);
or U14422 (N_14422,N_11050,N_9264);
and U14423 (N_14423,N_11031,N_11408);
or U14424 (N_14424,N_9046,N_11953);
or U14425 (N_14425,N_10653,N_10665);
nand U14426 (N_14426,N_9669,N_9309);
nor U14427 (N_14427,N_10805,N_9179);
or U14428 (N_14428,N_11226,N_9720);
and U14429 (N_14429,N_9252,N_10618);
xor U14430 (N_14430,N_9695,N_10341);
nand U14431 (N_14431,N_10529,N_10438);
and U14432 (N_14432,N_11458,N_10468);
nand U14433 (N_14433,N_10001,N_10389);
nand U14434 (N_14434,N_9226,N_9064);
xor U14435 (N_14435,N_10562,N_11341);
xor U14436 (N_14436,N_11743,N_9145);
nor U14437 (N_14437,N_9586,N_10655);
or U14438 (N_14438,N_11197,N_9443);
nand U14439 (N_14439,N_11305,N_9239);
and U14440 (N_14440,N_10835,N_11295);
xnor U14441 (N_14441,N_10671,N_9395);
nor U14442 (N_14442,N_10302,N_10291);
and U14443 (N_14443,N_10150,N_10775);
nor U14444 (N_14444,N_9164,N_11997);
and U14445 (N_14445,N_9578,N_9766);
and U14446 (N_14446,N_9729,N_9772);
xor U14447 (N_14447,N_9620,N_11953);
xnor U14448 (N_14448,N_10891,N_9499);
nand U14449 (N_14449,N_9821,N_9964);
nor U14450 (N_14450,N_9194,N_9462);
or U14451 (N_14451,N_9130,N_11527);
nor U14452 (N_14452,N_9008,N_11664);
or U14453 (N_14453,N_10758,N_9813);
or U14454 (N_14454,N_11688,N_11542);
xor U14455 (N_14455,N_11085,N_11026);
nand U14456 (N_14456,N_9044,N_11310);
nor U14457 (N_14457,N_9575,N_9576);
nand U14458 (N_14458,N_10614,N_10134);
or U14459 (N_14459,N_9453,N_11033);
or U14460 (N_14460,N_10554,N_9307);
nor U14461 (N_14461,N_11582,N_9040);
xnor U14462 (N_14462,N_9355,N_9631);
nand U14463 (N_14463,N_9260,N_9737);
xnor U14464 (N_14464,N_10794,N_9067);
or U14465 (N_14465,N_11082,N_9357);
nor U14466 (N_14466,N_9609,N_9177);
and U14467 (N_14467,N_11716,N_11502);
nand U14468 (N_14468,N_11078,N_11711);
or U14469 (N_14469,N_9891,N_10109);
xor U14470 (N_14470,N_11340,N_9266);
or U14471 (N_14471,N_10905,N_9742);
nor U14472 (N_14472,N_9530,N_10135);
xor U14473 (N_14473,N_11660,N_11727);
or U14474 (N_14474,N_10057,N_9465);
nor U14475 (N_14475,N_11290,N_10247);
nor U14476 (N_14476,N_9387,N_9308);
nor U14477 (N_14477,N_10464,N_9546);
or U14478 (N_14478,N_11950,N_9061);
nand U14479 (N_14479,N_10351,N_10692);
nor U14480 (N_14480,N_10010,N_11739);
nand U14481 (N_14481,N_11495,N_11182);
and U14482 (N_14482,N_10308,N_9352);
xnor U14483 (N_14483,N_11574,N_9792);
nor U14484 (N_14484,N_9838,N_11068);
and U14485 (N_14485,N_10346,N_10059);
nand U14486 (N_14486,N_9603,N_10778);
and U14487 (N_14487,N_10893,N_11827);
xnor U14488 (N_14488,N_9707,N_11489);
xnor U14489 (N_14489,N_10009,N_10215);
and U14490 (N_14490,N_9133,N_11097);
nor U14491 (N_14491,N_11695,N_10086);
and U14492 (N_14492,N_9185,N_10895);
nand U14493 (N_14493,N_10669,N_9204);
xor U14494 (N_14494,N_11603,N_11421);
nand U14495 (N_14495,N_10571,N_10669);
and U14496 (N_14496,N_9235,N_9708);
or U14497 (N_14497,N_9006,N_10943);
and U14498 (N_14498,N_9310,N_10192);
nand U14499 (N_14499,N_9556,N_10640);
and U14500 (N_14500,N_11912,N_9586);
and U14501 (N_14501,N_11569,N_11441);
nand U14502 (N_14502,N_9317,N_11030);
nand U14503 (N_14503,N_9781,N_11844);
or U14504 (N_14504,N_9058,N_9456);
xnor U14505 (N_14505,N_9895,N_10821);
and U14506 (N_14506,N_9341,N_11984);
and U14507 (N_14507,N_11811,N_9123);
nor U14508 (N_14508,N_10147,N_9502);
and U14509 (N_14509,N_11875,N_9090);
xor U14510 (N_14510,N_11950,N_11987);
nor U14511 (N_14511,N_9263,N_9833);
xnor U14512 (N_14512,N_10782,N_10851);
nand U14513 (N_14513,N_9895,N_9607);
or U14514 (N_14514,N_11205,N_9402);
or U14515 (N_14515,N_9573,N_11993);
or U14516 (N_14516,N_10352,N_10732);
nor U14517 (N_14517,N_10557,N_10046);
xnor U14518 (N_14518,N_11390,N_9154);
or U14519 (N_14519,N_9598,N_11598);
nor U14520 (N_14520,N_9071,N_10753);
and U14521 (N_14521,N_11670,N_11146);
nand U14522 (N_14522,N_11163,N_11758);
nor U14523 (N_14523,N_9937,N_11913);
and U14524 (N_14524,N_10220,N_10989);
and U14525 (N_14525,N_10537,N_9709);
xor U14526 (N_14526,N_10842,N_10354);
and U14527 (N_14527,N_9466,N_11210);
nor U14528 (N_14528,N_10867,N_11662);
nand U14529 (N_14529,N_11108,N_9246);
nor U14530 (N_14530,N_10822,N_10804);
nand U14531 (N_14531,N_11013,N_11173);
nand U14532 (N_14532,N_11474,N_9838);
or U14533 (N_14533,N_9963,N_9306);
and U14534 (N_14534,N_11057,N_9685);
or U14535 (N_14535,N_10950,N_11979);
xnor U14536 (N_14536,N_11082,N_10656);
nand U14537 (N_14537,N_9024,N_9694);
nor U14538 (N_14538,N_10741,N_11745);
nand U14539 (N_14539,N_11911,N_11424);
xnor U14540 (N_14540,N_10075,N_10921);
or U14541 (N_14541,N_9907,N_10737);
or U14542 (N_14542,N_11802,N_11684);
nand U14543 (N_14543,N_10370,N_11155);
xnor U14544 (N_14544,N_9041,N_9100);
xnor U14545 (N_14545,N_11967,N_9566);
nor U14546 (N_14546,N_10806,N_9060);
and U14547 (N_14547,N_9438,N_10072);
and U14548 (N_14548,N_11732,N_9804);
and U14549 (N_14549,N_11444,N_11438);
or U14550 (N_14550,N_9325,N_9043);
and U14551 (N_14551,N_10762,N_10542);
or U14552 (N_14552,N_9064,N_9445);
and U14553 (N_14553,N_10916,N_9153);
xor U14554 (N_14554,N_10504,N_9668);
xnor U14555 (N_14555,N_10171,N_9982);
and U14556 (N_14556,N_11808,N_11047);
or U14557 (N_14557,N_10863,N_9517);
or U14558 (N_14558,N_10285,N_9312);
nand U14559 (N_14559,N_11414,N_10888);
nand U14560 (N_14560,N_11227,N_11291);
or U14561 (N_14561,N_9260,N_11935);
nor U14562 (N_14562,N_9231,N_10198);
or U14563 (N_14563,N_11276,N_11504);
or U14564 (N_14564,N_11188,N_11967);
or U14565 (N_14565,N_11939,N_9781);
and U14566 (N_14566,N_11020,N_9277);
nor U14567 (N_14567,N_9151,N_10156);
and U14568 (N_14568,N_10211,N_11432);
or U14569 (N_14569,N_11193,N_10851);
and U14570 (N_14570,N_10878,N_11306);
nand U14571 (N_14571,N_11798,N_9670);
and U14572 (N_14572,N_11181,N_11247);
xnor U14573 (N_14573,N_11458,N_10866);
and U14574 (N_14574,N_9224,N_11169);
nand U14575 (N_14575,N_9993,N_9175);
xnor U14576 (N_14576,N_10627,N_11187);
nor U14577 (N_14577,N_10330,N_10998);
and U14578 (N_14578,N_11508,N_11520);
and U14579 (N_14579,N_11426,N_11374);
or U14580 (N_14580,N_9149,N_10453);
nand U14581 (N_14581,N_11426,N_9484);
and U14582 (N_14582,N_9158,N_10102);
nand U14583 (N_14583,N_9215,N_10621);
nor U14584 (N_14584,N_11650,N_10227);
and U14585 (N_14585,N_9244,N_10703);
nand U14586 (N_14586,N_11881,N_10287);
nand U14587 (N_14587,N_11698,N_10057);
and U14588 (N_14588,N_11194,N_9697);
xnor U14589 (N_14589,N_11469,N_9952);
nand U14590 (N_14590,N_10647,N_9716);
and U14591 (N_14591,N_9340,N_9353);
xnor U14592 (N_14592,N_10803,N_9364);
and U14593 (N_14593,N_11042,N_10637);
and U14594 (N_14594,N_9707,N_11490);
or U14595 (N_14595,N_10210,N_10566);
and U14596 (N_14596,N_11663,N_11825);
xor U14597 (N_14597,N_9359,N_9216);
and U14598 (N_14598,N_9668,N_11783);
and U14599 (N_14599,N_10309,N_10337);
xnor U14600 (N_14600,N_11701,N_11067);
and U14601 (N_14601,N_10444,N_10186);
xor U14602 (N_14602,N_11940,N_11249);
or U14603 (N_14603,N_11484,N_11442);
xnor U14604 (N_14604,N_9079,N_9967);
nor U14605 (N_14605,N_9520,N_10340);
nor U14606 (N_14606,N_11836,N_9099);
nand U14607 (N_14607,N_11587,N_9726);
xnor U14608 (N_14608,N_9414,N_10860);
or U14609 (N_14609,N_9654,N_11632);
nor U14610 (N_14610,N_11585,N_11360);
xor U14611 (N_14611,N_9768,N_11439);
nand U14612 (N_14612,N_9542,N_9325);
and U14613 (N_14613,N_9533,N_11926);
nor U14614 (N_14614,N_11408,N_11459);
xnor U14615 (N_14615,N_11228,N_9111);
nand U14616 (N_14616,N_9816,N_10358);
or U14617 (N_14617,N_10069,N_11659);
nor U14618 (N_14618,N_10267,N_10318);
and U14619 (N_14619,N_10436,N_10933);
and U14620 (N_14620,N_10718,N_11166);
nand U14621 (N_14621,N_10830,N_9885);
nand U14622 (N_14622,N_9956,N_10802);
nor U14623 (N_14623,N_10185,N_9664);
nor U14624 (N_14624,N_9254,N_9660);
or U14625 (N_14625,N_11047,N_10731);
and U14626 (N_14626,N_11446,N_11948);
nor U14627 (N_14627,N_9758,N_10071);
nor U14628 (N_14628,N_10579,N_10536);
nor U14629 (N_14629,N_11412,N_9642);
nor U14630 (N_14630,N_10227,N_9096);
nand U14631 (N_14631,N_10285,N_9254);
nor U14632 (N_14632,N_10674,N_11669);
nand U14633 (N_14633,N_10450,N_10478);
and U14634 (N_14634,N_9872,N_11526);
xnor U14635 (N_14635,N_11231,N_10103);
xnor U14636 (N_14636,N_9151,N_10081);
and U14637 (N_14637,N_9682,N_10078);
nor U14638 (N_14638,N_9558,N_11602);
and U14639 (N_14639,N_10703,N_11850);
xor U14640 (N_14640,N_11297,N_10314);
and U14641 (N_14641,N_9144,N_11191);
nand U14642 (N_14642,N_11977,N_11660);
nand U14643 (N_14643,N_11533,N_11910);
nor U14644 (N_14644,N_11135,N_9548);
or U14645 (N_14645,N_11624,N_10447);
and U14646 (N_14646,N_10830,N_10456);
and U14647 (N_14647,N_9196,N_9945);
xnor U14648 (N_14648,N_10863,N_11721);
nor U14649 (N_14649,N_9323,N_10567);
and U14650 (N_14650,N_11461,N_9219);
nand U14651 (N_14651,N_9174,N_10422);
nor U14652 (N_14652,N_11045,N_9409);
or U14653 (N_14653,N_11052,N_9866);
nand U14654 (N_14654,N_9106,N_9441);
and U14655 (N_14655,N_9665,N_10668);
nor U14656 (N_14656,N_11913,N_9798);
and U14657 (N_14657,N_10854,N_10622);
and U14658 (N_14658,N_11781,N_9882);
nor U14659 (N_14659,N_10761,N_11345);
nand U14660 (N_14660,N_11754,N_9271);
or U14661 (N_14661,N_11306,N_11102);
nor U14662 (N_14662,N_11914,N_11466);
xnor U14663 (N_14663,N_11357,N_10007);
nand U14664 (N_14664,N_10109,N_9565);
nand U14665 (N_14665,N_9779,N_9621);
xor U14666 (N_14666,N_10963,N_9302);
nor U14667 (N_14667,N_10954,N_11811);
and U14668 (N_14668,N_11373,N_11968);
and U14669 (N_14669,N_11245,N_10649);
nand U14670 (N_14670,N_9208,N_10363);
or U14671 (N_14671,N_10098,N_9010);
or U14672 (N_14672,N_11763,N_10197);
xor U14673 (N_14673,N_9249,N_11532);
xnor U14674 (N_14674,N_10751,N_10768);
nor U14675 (N_14675,N_9180,N_9744);
nand U14676 (N_14676,N_10663,N_10087);
nand U14677 (N_14677,N_9901,N_9012);
or U14678 (N_14678,N_10879,N_9970);
nand U14679 (N_14679,N_11803,N_11595);
nor U14680 (N_14680,N_9078,N_9528);
nor U14681 (N_14681,N_9464,N_9485);
nor U14682 (N_14682,N_11069,N_10996);
nand U14683 (N_14683,N_10246,N_10575);
nand U14684 (N_14684,N_11228,N_9668);
xnor U14685 (N_14685,N_11510,N_10572);
nand U14686 (N_14686,N_9102,N_11712);
xnor U14687 (N_14687,N_11314,N_10347);
or U14688 (N_14688,N_11004,N_10760);
xor U14689 (N_14689,N_10539,N_11385);
xor U14690 (N_14690,N_9105,N_10682);
xor U14691 (N_14691,N_9434,N_10077);
xnor U14692 (N_14692,N_11414,N_11439);
xnor U14693 (N_14693,N_11772,N_9213);
and U14694 (N_14694,N_9028,N_10838);
xor U14695 (N_14695,N_9870,N_11684);
or U14696 (N_14696,N_9862,N_9267);
or U14697 (N_14697,N_10208,N_9053);
nand U14698 (N_14698,N_10093,N_11794);
nand U14699 (N_14699,N_9327,N_11291);
or U14700 (N_14700,N_9606,N_10913);
xnor U14701 (N_14701,N_9682,N_9443);
nor U14702 (N_14702,N_11788,N_11643);
nor U14703 (N_14703,N_11694,N_11202);
nand U14704 (N_14704,N_11330,N_11215);
nor U14705 (N_14705,N_10836,N_9398);
nand U14706 (N_14706,N_10505,N_9544);
nand U14707 (N_14707,N_9270,N_11443);
nand U14708 (N_14708,N_11487,N_10946);
xnor U14709 (N_14709,N_10269,N_10773);
and U14710 (N_14710,N_9266,N_10127);
xnor U14711 (N_14711,N_11358,N_9840);
or U14712 (N_14712,N_9419,N_10112);
xor U14713 (N_14713,N_10190,N_10614);
and U14714 (N_14714,N_10632,N_11464);
xor U14715 (N_14715,N_9780,N_10973);
and U14716 (N_14716,N_10317,N_9760);
and U14717 (N_14717,N_10326,N_11458);
or U14718 (N_14718,N_9568,N_9804);
and U14719 (N_14719,N_10499,N_9317);
nand U14720 (N_14720,N_9365,N_10891);
nor U14721 (N_14721,N_10225,N_10175);
nand U14722 (N_14722,N_9872,N_10807);
nand U14723 (N_14723,N_9618,N_10094);
nand U14724 (N_14724,N_11798,N_9550);
xnor U14725 (N_14725,N_10392,N_11001);
or U14726 (N_14726,N_9159,N_9990);
nor U14727 (N_14727,N_10212,N_9049);
and U14728 (N_14728,N_9647,N_10713);
or U14729 (N_14729,N_11941,N_11389);
nand U14730 (N_14730,N_10163,N_9857);
and U14731 (N_14731,N_11592,N_10493);
and U14732 (N_14732,N_11327,N_9544);
and U14733 (N_14733,N_9965,N_10891);
xnor U14734 (N_14734,N_11493,N_11849);
nor U14735 (N_14735,N_10786,N_9836);
and U14736 (N_14736,N_9595,N_10478);
nand U14737 (N_14737,N_10390,N_9240);
xnor U14738 (N_14738,N_10341,N_9528);
and U14739 (N_14739,N_11622,N_9382);
xnor U14740 (N_14740,N_9192,N_11489);
nand U14741 (N_14741,N_9519,N_10935);
xor U14742 (N_14742,N_9688,N_11627);
or U14743 (N_14743,N_11775,N_10236);
and U14744 (N_14744,N_11840,N_11279);
nand U14745 (N_14745,N_9388,N_10635);
and U14746 (N_14746,N_10292,N_9580);
or U14747 (N_14747,N_10657,N_11705);
xnor U14748 (N_14748,N_9158,N_11179);
nand U14749 (N_14749,N_11391,N_10300);
or U14750 (N_14750,N_9553,N_10203);
nor U14751 (N_14751,N_9680,N_10962);
xor U14752 (N_14752,N_9660,N_11679);
or U14753 (N_14753,N_10913,N_10410);
nand U14754 (N_14754,N_9652,N_9118);
xor U14755 (N_14755,N_11308,N_9384);
or U14756 (N_14756,N_11135,N_9940);
nor U14757 (N_14757,N_11059,N_9141);
and U14758 (N_14758,N_10602,N_11117);
nand U14759 (N_14759,N_9099,N_9523);
nand U14760 (N_14760,N_10869,N_10067);
nor U14761 (N_14761,N_10825,N_10449);
nand U14762 (N_14762,N_11812,N_10474);
and U14763 (N_14763,N_10113,N_10641);
nand U14764 (N_14764,N_9573,N_11659);
or U14765 (N_14765,N_11114,N_11709);
nor U14766 (N_14766,N_10703,N_9615);
nand U14767 (N_14767,N_10084,N_10142);
xor U14768 (N_14768,N_11152,N_9349);
nor U14769 (N_14769,N_10735,N_10148);
or U14770 (N_14770,N_9027,N_10922);
nor U14771 (N_14771,N_10286,N_11440);
or U14772 (N_14772,N_11230,N_11324);
nand U14773 (N_14773,N_9863,N_9191);
nand U14774 (N_14774,N_10773,N_10616);
and U14775 (N_14775,N_9659,N_10248);
xnor U14776 (N_14776,N_10577,N_9300);
nor U14777 (N_14777,N_9566,N_10889);
and U14778 (N_14778,N_11200,N_9229);
or U14779 (N_14779,N_10317,N_10470);
nand U14780 (N_14780,N_10074,N_11650);
or U14781 (N_14781,N_9121,N_10995);
or U14782 (N_14782,N_10644,N_11374);
or U14783 (N_14783,N_9843,N_10712);
or U14784 (N_14784,N_10487,N_10960);
and U14785 (N_14785,N_10407,N_11404);
xnor U14786 (N_14786,N_11701,N_11048);
or U14787 (N_14787,N_10964,N_9762);
or U14788 (N_14788,N_10064,N_10272);
or U14789 (N_14789,N_11663,N_9153);
or U14790 (N_14790,N_9669,N_11161);
or U14791 (N_14791,N_9949,N_9399);
or U14792 (N_14792,N_11065,N_11764);
or U14793 (N_14793,N_11522,N_10250);
and U14794 (N_14794,N_10701,N_9102);
nand U14795 (N_14795,N_10491,N_11963);
and U14796 (N_14796,N_10827,N_10222);
nor U14797 (N_14797,N_11402,N_9916);
nor U14798 (N_14798,N_10478,N_10728);
xor U14799 (N_14799,N_9970,N_9061);
or U14800 (N_14800,N_10236,N_11154);
nand U14801 (N_14801,N_10258,N_9501);
nor U14802 (N_14802,N_10420,N_9962);
xor U14803 (N_14803,N_9444,N_11154);
or U14804 (N_14804,N_9279,N_11784);
nor U14805 (N_14805,N_11907,N_10460);
xnor U14806 (N_14806,N_9686,N_11013);
xor U14807 (N_14807,N_11131,N_11471);
and U14808 (N_14808,N_9632,N_9706);
and U14809 (N_14809,N_11707,N_9761);
and U14810 (N_14810,N_9973,N_11488);
nand U14811 (N_14811,N_9765,N_10331);
xor U14812 (N_14812,N_11794,N_11575);
nand U14813 (N_14813,N_10945,N_10323);
xnor U14814 (N_14814,N_9953,N_11120);
or U14815 (N_14815,N_9267,N_11471);
and U14816 (N_14816,N_10562,N_11220);
nand U14817 (N_14817,N_9054,N_11660);
and U14818 (N_14818,N_11943,N_10078);
or U14819 (N_14819,N_11485,N_11201);
and U14820 (N_14820,N_9513,N_11403);
and U14821 (N_14821,N_11140,N_10472);
nor U14822 (N_14822,N_11858,N_11486);
xor U14823 (N_14823,N_10438,N_10969);
nand U14824 (N_14824,N_9355,N_9632);
or U14825 (N_14825,N_11716,N_11801);
xnor U14826 (N_14826,N_10953,N_11015);
and U14827 (N_14827,N_9400,N_10862);
or U14828 (N_14828,N_10117,N_10853);
xnor U14829 (N_14829,N_10774,N_9630);
nor U14830 (N_14830,N_11434,N_11711);
xor U14831 (N_14831,N_10283,N_10799);
nand U14832 (N_14832,N_9580,N_9101);
and U14833 (N_14833,N_11436,N_10872);
xor U14834 (N_14834,N_9048,N_11719);
nand U14835 (N_14835,N_10170,N_11864);
nor U14836 (N_14836,N_9873,N_10881);
xnor U14837 (N_14837,N_9942,N_9639);
and U14838 (N_14838,N_11605,N_10397);
and U14839 (N_14839,N_10300,N_11603);
nor U14840 (N_14840,N_11486,N_11289);
nand U14841 (N_14841,N_10757,N_11680);
nor U14842 (N_14842,N_10035,N_11811);
nand U14843 (N_14843,N_9568,N_10006);
nor U14844 (N_14844,N_9601,N_10357);
nor U14845 (N_14845,N_11924,N_11200);
nand U14846 (N_14846,N_11642,N_10185);
nor U14847 (N_14847,N_9840,N_10910);
nand U14848 (N_14848,N_11603,N_9793);
nor U14849 (N_14849,N_9064,N_10080);
nor U14850 (N_14850,N_9311,N_10626);
nor U14851 (N_14851,N_10047,N_10080);
or U14852 (N_14852,N_11972,N_10533);
nand U14853 (N_14853,N_10273,N_10778);
or U14854 (N_14854,N_9261,N_10399);
nor U14855 (N_14855,N_9754,N_10780);
nor U14856 (N_14856,N_9179,N_10870);
xnor U14857 (N_14857,N_11788,N_9181);
nor U14858 (N_14858,N_11220,N_10554);
xor U14859 (N_14859,N_9874,N_10670);
and U14860 (N_14860,N_10431,N_11145);
xor U14861 (N_14861,N_9199,N_11818);
and U14862 (N_14862,N_10849,N_10540);
and U14863 (N_14863,N_10551,N_9003);
and U14864 (N_14864,N_11596,N_11028);
and U14865 (N_14865,N_9064,N_11779);
or U14866 (N_14866,N_10850,N_11858);
or U14867 (N_14867,N_11295,N_11573);
or U14868 (N_14868,N_11719,N_10030);
or U14869 (N_14869,N_10860,N_10464);
nand U14870 (N_14870,N_11457,N_10869);
nand U14871 (N_14871,N_9452,N_11244);
nand U14872 (N_14872,N_10415,N_10457);
nor U14873 (N_14873,N_10843,N_10488);
xor U14874 (N_14874,N_11816,N_9566);
xnor U14875 (N_14875,N_9575,N_10058);
or U14876 (N_14876,N_9244,N_11170);
nor U14877 (N_14877,N_10189,N_10918);
nor U14878 (N_14878,N_11466,N_9125);
and U14879 (N_14879,N_10822,N_9601);
or U14880 (N_14880,N_11463,N_11114);
nor U14881 (N_14881,N_9125,N_11666);
nand U14882 (N_14882,N_10294,N_11100);
or U14883 (N_14883,N_11159,N_10913);
and U14884 (N_14884,N_10299,N_11775);
or U14885 (N_14885,N_10828,N_9236);
and U14886 (N_14886,N_11697,N_9546);
xor U14887 (N_14887,N_9377,N_9281);
or U14888 (N_14888,N_11829,N_10990);
nor U14889 (N_14889,N_9986,N_10968);
or U14890 (N_14890,N_11307,N_11903);
and U14891 (N_14891,N_10273,N_10327);
nand U14892 (N_14892,N_9722,N_9413);
and U14893 (N_14893,N_9351,N_9759);
xor U14894 (N_14894,N_9372,N_10228);
or U14895 (N_14895,N_9025,N_11850);
or U14896 (N_14896,N_9836,N_11854);
nor U14897 (N_14897,N_9712,N_11485);
and U14898 (N_14898,N_9701,N_10117);
xor U14899 (N_14899,N_11705,N_9468);
and U14900 (N_14900,N_11247,N_9898);
nor U14901 (N_14901,N_9004,N_10179);
or U14902 (N_14902,N_11238,N_10349);
or U14903 (N_14903,N_9244,N_9425);
xor U14904 (N_14904,N_9740,N_11276);
xnor U14905 (N_14905,N_11735,N_10568);
xor U14906 (N_14906,N_9142,N_9395);
or U14907 (N_14907,N_10356,N_10385);
nor U14908 (N_14908,N_11488,N_9931);
or U14909 (N_14909,N_10116,N_9263);
xnor U14910 (N_14910,N_11738,N_9260);
xnor U14911 (N_14911,N_10902,N_11173);
and U14912 (N_14912,N_11164,N_11195);
and U14913 (N_14913,N_9459,N_10928);
nand U14914 (N_14914,N_11999,N_9587);
nand U14915 (N_14915,N_11478,N_11084);
or U14916 (N_14916,N_10250,N_9089);
nand U14917 (N_14917,N_9942,N_11309);
nor U14918 (N_14918,N_11586,N_9136);
nand U14919 (N_14919,N_11910,N_9720);
xnor U14920 (N_14920,N_10771,N_10340);
or U14921 (N_14921,N_10550,N_11829);
nor U14922 (N_14922,N_11248,N_9422);
xor U14923 (N_14923,N_10032,N_9960);
and U14924 (N_14924,N_9478,N_10309);
nor U14925 (N_14925,N_10981,N_9995);
xnor U14926 (N_14926,N_9873,N_11385);
and U14927 (N_14927,N_10736,N_11218);
and U14928 (N_14928,N_11283,N_10863);
or U14929 (N_14929,N_11205,N_10546);
and U14930 (N_14930,N_9066,N_10233);
and U14931 (N_14931,N_9775,N_9465);
nand U14932 (N_14932,N_11239,N_11060);
xor U14933 (N_14933,N_11236,N_11625);
nor U14934 (N_14934,N_10325,N_9536);
nor U14935 (N_14935,N_10254,N_10929);
and U14936 (N_14936,N_9261,N_11884);
nand U14937 (N_14937,N_11057,N_9654);
nand U14938 (N_14938,N_10149,N_10884);
or U14939 (N_14939,N_9647,N_9799);
or U14940 (N_14940,N_11915,N_10757);
and U14941 (N_14941,N_10285,N_10178);
nand U14942 (N_14942,N_10854,N_11319);
and U14943 (N_14943,N_10902,N_9916);
xnor U14944 (N_14944,N_9099,N_11591);
xnor U14945 (N_14945,N_11966,N_11969);
xnor U14946 (N_14946,N_9857,N_10719);
nand U14947 (N_14947,N_10736,N_10668);
nor U14948 (N_14948,N_10712,N_11153);
and U14949 (N_14949,N_10587,N_9932);
nor U14950 (N_14950,N_9935,N_11504);
and U14951 (N_14951,N_10508,N_9452);
and U14952 (N_14952,N_11402,N_11529);
nand U14953 (N_14953,N_11037,N_10569);
nor U14954 (N_14954,N_9039,N_9369);
nor U14955 (N_14955,N_9974,N_11485);
nand U14956 (N_14956,N_9743,N_9590);
nor U14957 (N_14957,N_10707,N_11501);
xor U14958 (N_14958,N_9331,N_9709);
xor U14959 (N_14959,N_9360,N_10399);
and U14960 (N_14960,N_11975,N_11958);
or U14961 (N_14961,N_11517,N_11338);
and U14962 (N_14962,N_11904,N_11196);
nor U14963 (N_14963,N_11889,N_11015);
and U14964 (N_14964,N_9712,N_11448);
nand U14965 (N_14965,N_11971,N_11746);
xnor U14966 (N_14966,N_11973,N_11828);
or U14967 (N_14967,N_11006,N_10077);
and U14968 (N_14968,N_9443,N_10221);
xor U14969 (N_14969,N_11292,N_11707);
nand U14970 (N_14970,N_10818,N_11667);
xor U14971 (N_14971,N_11226,N_10026);
nor U14972 (N_14972,N_11043,N_9661);
and U14973 (N_14973,N_10021,N_11443);
xnor U14974 (N_14974,N_10681,N_10451);
nor U14975 (N_14975,N_10759,N_11216);
xnor U14976 (N_14976,N_11454,N_10482);
and U14977 (N_14977,N_10129,N_9764);
nand U14978 (N_14978,N_9503,N_10843);
or U14979 (N_14979,N_11206,N_11549);
nand U14980 (N_14980,N_11781,N_9633);
nand U14981 (N_14981,N_10810,N_11563);
nand U14982 (N_14982,N_10687,N_9545);
and U14983 (N_14983,N_10746,N_11393);
xnor U14984 (N_14984,N_9049,N_10617);
nand U14985 (N_14985,N_9288,N_10394);
and U14986 (N_14986,N_9391,N_11755);
nand U14987 (N_14987,N_9594,N_10286);
nand U14988 (N_14988,N_11798,N_10582);
nor U14989 (N_14989,N_10542,N_11685);
and U14990 (N_14990,N_11183,N_10583);
nand U14991 (N_14991,N_10750,N_9155);
xor U14992 (N_14992,N_11694,N_11936);
xnor U14993 (N_14993,N_11384,N_10794);
xor U14994 (N_14994,N_10073,N_11271);
or U14995 (N_14995,N_10406,N_9763);
xnor U14996 (N_14996,N_9653,N_10144);
or U14997 (N_14997,N_11934,N_11860);
nand U14998 (N_14998,N_11754,N_11636);
nor U14999 (N_14999,N_9295,N_9635);
nor U15000 (N_15000,N_12173,N_12542);
xnor U15001 (N_15001,N_13990,N_12258);
xor U15002 (N_15002,N_13820,N_13120);
or U15003 (N_15003,N_13171,N_13720);
and U15004 (N_15004,N_12005,N_13375);
and U15005 (N_15005,N_12041,N_12358);
and U15006 (N_15006,N_14360,N_13695);
or U15007 (N_15007,N_14902,N_13381);
and U15008 (N_15008,N_13573,N_13559);
nand U15009 (N_15009,N_14586,N_13692);
and U15010 (N_15010,N_13275,N_14112);
and U15011 (N_15011,N_14654,N_12737);
and U15012 (N_15012,N_13551,N_12325);
nor U15013 (N_15013,N_14831,N_14688);
nand U15014 (N_15014,N_13116,N_13723);
and U15015 (N_15015,N_13525,N_14712);
nor U15016 (N_15016,N_12130,N_13217);
or U15017 (N_15017,N_13958,N_12416);
xor U15018 (N_15018,N_12611,N_12863);
nor U15019 (N_15019,N_12397,N_13192);
nand U15020 (N_15020,N_14630,N_14009);
or U15021 (N_15021,N_14834,N_14737);
or U15022 (N_15022,N_13486,N_14619);
or U15023 (N_15023,N_14919,N_14217);
and U15024 (N_15024,N_14943,N_12393);
and U15025 (N_15025,N_14136,N_14304);
or U15026 (N_15026,N_12370,N_13665);
or U15027 (N_15027,N_12981,N_12197);
nor U15028 (N_15028,N_12294,N_12208);
nand U15029 (N_15029,N_14507,N_13207);
xor U15030 (N_15030,N_13930,N_12374);
nand U15031 (N_15031,N_13554,N_12302);
xor U15032 (N_15032,N_12944,N_12570);
and U15033 (N_15033,N_13014,N_12025);
xor U15034 (N_15034,N_14195,N_13762);
nand U15035 (N_15035,N_14940,N_14730);
nand U15036 (N_15036,N_12257,N_13511);
nor U15037 (N_15037,N_13356,N_13556);
or U15038 (N_15038,N_14419,N_12424);
xor U15039 (N_15039,N_13267,N_12878);
nand U15040 (N_15040,N_12379,N_12743);
nand U15041 (N_15041,N_13727,N_14692);
and U15042 (N_15042,N_12028,N_13080);
or U15043 (N_15043,N_12266,N_12506);
xnor U15044 (N_15044,N_12313,N_14910);
nand U15045 (N_15045,N_12118,N_12603);
nor U15046 (N_15046,N_12514,N_14584);
and U15047 (N_15047,N_12732,N_12591);
nor U15048 (N_15048,N_14708,N_12515);
nor U15049 (N_15049,N_14656,N_12177);
and U15050 (N_15050,N_13834,N_14955);
or U15051 (N_15051,N_12823,N_13542);
nor U15052 (N_15052,N_13659,N_13054);
or U15053 (N_15053,N_14732,N_13589);
nand U15054 (N_15054,N_13307,N_13165);
xor U15055 (N_15055,N_14398,N_14331);
nor U15056 (N_15056,N_14048,N_14828);
and U15057 (N_15057,N_12955,N_12982);
xnor U15058 (N_15058,N_12085,N_13445);
nor U15059 (N_15059,N_12960,N_12421);
nor U15060 (N_15060,N_13785,N_13143);
or U15061 (N_15061,N_14721,N_13774);
or U15062 (N_15062,N_12939,N_14521);
or U15063 (N_15063,N_13633,N_14582);
nor U15064 (N_15064,N_12324,N_13948);
nor U15065 (N_15065,N_12436,N_14290);
nand U15066 (N_15066,N_12880,N_12655);
xnor U15067 (N_15067,N_12711,N_12274);
and U15068 (N_15068,N_12022,N_14556);
and U15069 (N_15069,N_14853,N_14799);
xnor U15070 (N_15070,N_14237,N_14030);
xnor U15071 (N_15071,N_13044,N_12661);
nand U15072 (N_15072,N_13691,N_14034);
nor U15073 (N_15073,N_14565,N_12652);
or U15074 (N_15074,N_14364,N_13297);
nor U15075 (N_15075,N_13992,N_12073);
and U15076 (N_15076,N_12705,N_13470);
nand U15077 (N_15077,N_13840,N_14043);
nand U15078 (N_15078,N_12192,N_13138);
nand U15079 (N_15079,N_14776,N_12327);
and U15080 (N_15080,N_12024,N_13400);
xor U15081 (N_15081,N_14281,N_12253);
xor U15082 (N_15082,N_12228,N_14618);
or U15083 (N_15083,N_14527,N_12355);
xnor U15084 (N_15084,N_12605,N_14923);
nor U15085 (N_15085,N_12282,N_13802);
nor U15086 (N_15086,N_12383,N_13056);
and U15087 (N_15087,N_14413,N_14514);
nand U15088 (N_15088,N_13202,N_13117);
xor U15089 (N_15089,N_12268,N_14566);
xor U15090 (N_15090,N_12456,N_12080);
or U15091 (N_15091,N_14523,N_14942);
and U15092 (N_15092,N_13332,N_14354);
nand U15093 (N_15093,N_13372,N_14323);
xnor U15094 (N_15094,N_14675,N_13137);
xnor U15095 (N_15095,N_12101,N_12149);
or U15096 (N_15096,N_13708,N_13450);
or U15097 (N_15097,N_12914,N_12773);
nand U15098 (N_15098,N_13805,N_12599);
xor U15099 (N_15099,N_12278,N_12115);
xnor U15100 (N_15100,N_13623,N_12622);
or U15101 (N_15101,N_14664,N_14599);
nand U15102 (N_15102,N_14286,N_13485);
and U15103 (N_15103,N_13367,N_12754);
and U15104 (N_15104,N_14744,N_14472);
nand U15105 (N_15105,N_14231,N_14138);
or U15106 (N_15106,N_12047,N_12909);
or U15107 (N_15107,N_14023,N_12059);
or U15108 (N_15108,N_12812,N_14669);
and U15109 (N_15109,N_12550,N_14441);
or U15110 (N_15110,N_12986,N_13684);
xnor U15111 (N_15111,N_12789,N_14626);
xor U15112 (N_15112,N_12116,N_14309);
nor U15113 (N_15113,N_14199,N_13399);
nor U15114 (N_15114,N_12160,N_12869);
nand U15115 (N_15115,N_12065,N_14438);
nand U15116 (N_15116,N_13827,N_13033);
and U15117 (N_15117,N_12345,N_13235);
nand U15118 (N_15118,N_12633,N_14247);
or U15119 (N_15119,N_14899,N_14386);
or U15120 (N_15120,N_12592,N_14738);
and U15121 (N_15121,N_12326,N_12105);
and U15122 (N_15122,N_14307,N_12348);
and U15123 (N_15123,N_13568,N_12169);
xnor U15124 (N_15124,N_13850,N_14239);
and U15125 (N_15125,N_14118,N_12290);
or U15126 (N_15126,N_12568,N_13678);
or U15127 (N_15127,N_12261,N_14020);
nand U15128 (N_15128,N_12061,N_14857);
and U15129 (N_15129,N_12497,N_12488);
or U15130 (N_15130,N_13985,N_14187);
nor U15131 (N_15131,N_12910,N_13815);
and U15132 (N_15132,N_13787,N_13913);
nor U15133 (N_15133,N_13466,N_13318);
nand U15134 (N_15134,N_13639,N_13861);
or U15135 (N_15135,N_14442,N_12104);
nor U15136 (N_15136,N_13422,N_14612);
and U15137 (N_15137,N_13680,N_14215);
nand U15138 (N_15138,N_12207,N_14068);
or U15139 (N_15139,N_12484,N_13614);
nor U15140 (N_15140,N_13387,N_13225);
xnor U15141 (N_15141,N_14934,N_12174);
or U15142 (N_15142,N_13984,N_14851);
xor U15143 (N_15143,N_12749,N_14054);
xor U15144 (N_15144,N_12153,N_14314);
xnor U15145 (N_15145,N_12018,N_12466);
nor U15146 (N_15146,N_12913,N_14969);
xnor U15147 (N_15147,N_12224,N_14303);
xnor U15148 (N_15148,N_14985,N_13208);
or U15149 (N_15149,N_14097,N_14752);
and U15150 (N_15150,N_12434,N_14840);
and U15151 (N_15151,N_12539,N_12412);
xor U15152 (N_15152,N_12482,N_12013);
nand U15153 (N_15153,N_13089,N_13915);
nor U15154 (N_15154,N_14078,N_13880);
xor U15155 (N_15155,N_12481,N_13465);
or U15156 (N_15156,N_12492,N_13978);
and U15157 (N_15157,N_13546,N_12810);
and U15158 (N_15158,N_13900,N_14476);
and U15159 (N_15159,N_12446,N_14515);
xnor U15160 (N_15160,N_14850,N_14003);
xor U15161 (N_15161,N_14720,N_13376);
xor U15162 (N_15162,N_12091,N_13083);
nand U15163 (N_15163,N_12043,N_14803);
nor U15164 (N_15164,N_14461,N_13418);
or U15165 (N_15165,N_12631,N_13016);
and U15166 (N_15166,N_13847,N_13241);
nor U15167 (N_15167,N_13273,N_14494);
and U15168 (N_15168,N_12010,N_14298);
nand U15169 (N_15169,N_12624,N_14065);
or U15170 (N_15170,N_12175,N_14497);
or U15171 (N_15171,N_12537,N_13547);
nor U15172 (N_15172,N_13876,N_12185);
nor U15173 (N_15173,N_12796,N_13715);
or U15174 (N_15174,N_12447,N_12276);
xnor U15175 (N_15175,N_14946,N_13963);
xnor U15176 (N_15176,N_14904,N_12628);
or U15177 (N_15177,N_12577,N_12837);
or U15178 (N_15178,N_14271,N_13378);
nor U15179 (N_15179,N_14905,N_12021);
or U15180 (N_15180,N_13611,N_13074);
nand U15181 (N_15181,N_12865,N_14150);
xor U15182 (N_15182,N_13062,N_14255);
nor U15183 (N_15183,N_13673,N_13187);
and U15184 (N_15184,N_14777,N_14953);
xnor U15185 (N_15185,N_13177,N_14723);
and U15186 (N_15186,N_13725,N_13687);
nand U15187 (N_15187,N_12833,N_14643);
nand U15188 (N_15188,N_13446,N_14986);
or U15189 (N_15189,N_14207,N_14872);
nand U15190 (N_15190,N_13879,N_13620);
nand U15191 (N_15191,N_12825,N_12522);
xnor U15192 (N_15192,N_14225,N_13726);
nand U15193 (N_15193,N_12180,N_12891);
nand U15194 (N_15194,N_13778,N_14547);
or U15195 (N_15195,N_14633,N_12656);
xor U15196 (N_15196,N_14498,N_14211);
and U15197 (N_15197,N_13451,N_14074);
and U15198 (N_15198,N_14987,N_12887);
and U15199 (N_15199,N_13025,N_12181);
nand U15200 (N_15200,N_13150,N_12708);
xnor U15201 (N_15201,N_12214,N_14775);
and U15202 (N_15202,N_12694,N_13262);
and U15203 (N_15203,N_13058,N_14763);
nand U15204 (N_15204,N_12395,N_13944);
and U15205 (N_15205,N_13188,N_14410);
nand U15206 (N_15206,N_13951,N_13925);
or U15207 (N_15207,N_12988,N_14022);
and U15208 (N_15208,N_12161,N_13388);
and U15209 (N_15209,N_13218,N_14597);
and U15210 (N_15210,N_12513,N_12961);
or U15211 (N_15211,N_14448,N_13411);
xor U15212 (N_15212,N_12541,N_14321);
or U15213 (N_15213,N_12834,N_13652);
or U15214 (N_15214,N_13705,N_14809);
xnor U15215 (N_15215,N_12643,N_12042);
nor U15216 (N_15216,N_13108,N_14100);
xnor U15217 (N_15217,N_14079,N_13352);
or U15218 (N_15218,N_13416,N_13917);
and U15219 (N_15219,N_13906,N_12333);
nand U15220 (N_15220,N_12686,N_13882);
or U15221 (N_15221,N_13460,N_13185);
xor U15222 (N_15222,N_13902,N_13309);
and U15223 (N_15223,N_13027,N_13512);
xnor U15224 (N_15224,N_13069,N_13361);
or U15225 (N_15225,N_13085,N_13059);
or U15226 (N_15226,N_13467,N_13480);
nor U15227 (N_15227,N_12963,N_13205);
or U15228 (N_15228,N_12965,N_13908);
nor U15229 (N_15229,N_13515,N_13812);
nand U15230 (N_15230,N_14788,N_12584);
or U15231 (N_15231,N_12574,N_12525);
nand U15232 (N_15232,N_13934,N_12895);
xnor U15233 (N_15233,N_12793,N_12874);
and U15234 (N_15234,N_14812,N_14791);
xor U15235 (N_15235,N_12365,N_12163);
nand U15236 (N_15236,N_12002,N_12848);
xor U15237 (N_15237,N_12719,N_12741);
or U15238 (N_15238,N_12517,N_14362);
nor U15239 (N_15239,N_13417,N_13575);
nor U15240 (N_15240,N_14361,N_14474);
or U15241 (N_15241,N_12875,N_13532);
or U15242 (N_15242,N_13312,N_12146);
xnor U15243 (N_15243,N_12461,N_13959);
nor U15244 (N_15244,N_14184,N_14610);
and U15245 (N_15245,N_13191,N_14844);
nand U15246 (N_15246,N_13580,N_12016);
nor U15247 (N_15247,N_13008,N_14085);
nor U15248 (N_15248,N_14722,N_12150);
nor U15249 (N_15249,N_12236,N_13162);
nor U15250 (N_15250,N_12120,N_14911);
xor U15251 (N_15251,N_12337,N_14459);
nor U15252 (N_15252,N_13326,N_13330);
nor U15253 (N_15253,N_13023,N_14188);
xnor U15254 (N_15254,N_13569,N_12563);
nor U15255 (N_15255,N_12629,N_13055);
or U15256 (N_15256,N_13997,N_12778);
xnor U15257 (N_15257,N_12809,N_14778);
nand U15258 (N_15258,N_13746,N_13303);
nor U15259 (N_15259,N_14593,N_14734);
nand U15260 (N_15260,N_14363,N_14223);
or U15261 (N_15261,N_13872,N_14843);
nor U15262 (N_15262,N_14384,N_14014);
and U15263 (N_15263,N_14457,N_12193);
or U15264 (N_15264,N_13000,N_14089);
and U15265 (N_15265,N_13282,N_13338);
nor U15266 (N_15266,N_14701,N_13604);
and U15267 (N_15267,N_13586,N_12870);
xor U15268 (N_15268,N_12435,N_13178);
nand U15269 (N_15269,N_14815,N_14502);
xnor U15270 (N_15270,N_14168,N_12382);
and U15271 (N_15271,N_14756,N_12746);
nor U15272 (N_15272,N_13764,N_14257);
nor U15273 (N_15273,N_14587,N_12400);
or U15274 (N_15274,N_13777,N_12219);
nand U15275 (N_15275,N_13219,N_13548);
nor U15276 (N_15276,N_14149,N_13989);
nor U15277 (N_15277,N_12221,N_12677);
nand U15278 (N_15278,N_12508,N_13365);
nor U15279 (N_15279,N_13160,N_12191);
nand U15280 (N_15280,N_14259,N_14278);
nand U15281 (N_15281,N_12331,N_13829);
or U15282 (N_15282,N_13881,N_14050);
and U15283 (N_15283,N_13118,N_12996);
or U15284 (N_15284,N_14007,N_13730);
nand U15285 (N_15285,N_12103,N_12269);
or U15286 (N_15286,N_13447,N_12272);
and U15287 (N_15287,N_14277,N_13223);
nor U15288 (N_15288,N_14931,N_12453);
nand U15289 (N_15289,N_12849,N_13813);
nor U15290 (N_15290,N_14491,N_12134);
xor U15291 (N_15291,N_14092,N_12084);
xnor U15292 (N_15292,N_14885,N_14864);
nor U15293 (N_15293,N_13866,N_12625);
or U15294 (N_15294,N_13701,N_13270);
nand U15295 (N_15295,N_14997,N_14948);
xnor U15296 (N_15296,N_12317,N_13030);
or U15297 (N_15297,N_12441,N_13032);
xor U15298 (N_15298,N_12738,N_13851);
xnor U15299 (N_15299,N_13714,N_14390);
nand U15300 (N_15300,N_13170,N_14169);
or U15301 (N_15301,N_13587,N_13344);
nor U15302 (N_15302,N_12557,N_13197);
nor U15303 (N_15303,N_12926,N_13919);
nand U15304 (N_15304,N_14867,N_14596);
or U15305 (N_15305,N_12143,N_12703);
or U15306 (N_15306,N_12035,N_12666);
or U15307 (N_15307,N_13671,N_14280);
or U15308 (N_15308,N_12538,N_12889);
nor U15309 (N_15309,N_14095,N_13891);
or U15310 (N_15310,N_13250,N_13644);
and U15311 (N_15311,N_13981,N_14288);
xor U15312 (N_15312,N_14016,N_14403);
and U15313 (N_15313,N_14486,N_13564);
or U15314 (N_15314,N_12170,N_12945);
nand U15315 (N_15315,N_12255,N_13078);
and U15316 (N_15316,N_13412,N_14975);
or U15317 (N_15317,N_12725,N_12690);
nor U15318 (N_15318,N_13535,N_12921);
nor U15319 (N_15319,N_14427,N_14965);
nand U15320 (N_15320,N_14519,N_12606);
xnor U15321 (N_15321,N_14120,N_14141);
xor U15322 (N_15322,N_14534,N_14518);
xor U15323 (N_15323,N_12136,N_14532);
xnor U15324 (N_15324,N_14665,N_13859);
xnor U15325 (N_15325,N_14289,N_14103);
and U15326 (N_15326,N_12798,N_13885);
xor U15327 (N_15327,N_12263,N_13093);
nand U15328 (N_15328,N_14718,N_14276);
nor U15329 (N_15329,N_12868,N_14914);
nand U15330 (N_15330,N_13733,N_13144);
or U15331 (N_15331,N_13822,N_14176);
nand U15332 (N_15332,N_12908,N_13592);
nor U15333 (N_15333,N_14130,N_12227);
xnor U15334 (N_15334,N_14185,N_14949);
or U15335 (N_15335,N_13193,N_12756);
and U15336 (N_15336,N_13686,N_12051);
xnor U15337 (N_15337,N_13227,N_12604);
nand U15338 (N_15338,N_12375,N_12581);
and U15339 (N_15339,N_13619,N_14595);
nor U15340 (N_15340,N_14039,N_13555);
or U15341 (N_15341,N_13499,N_13938);
or U15342 (N_15342,N_12768,N_12060);
nor U15343 (N_15343,N_12437,N_13111);
nand U15344 (N_15344,N_14898,N_13816);
and U15345 (N_15345,N_12415,N_13622);
nor U15346 (N_15346,N_14495,N_14637);
or U15347 (N_15347,N_12423,N_14880);
or U15348 (N_15348,N_14273,N_14310);
nand U15349 (N_15349,N_12480,N_13797);
nor U15350 (N_15350,N_13368,N_12784);
nor U15351 (N_15351,N_12128,N_14159);
nand U15352 (N_15352,N_12767,N_14699);
xor U15353 (N_15353,N_14069,N_12439);
or U15354 (N_15354,N_12905,N_12695);
and U15355 (N_15355,N_12171,N_13645);
nand U15356 (N_15356,N_14397,N_13302);
and U15357 (N_15357,N_12413,N_12699);
or U15358 (N_15358,N_12806,N_12818);
nor U15359 (N_15359,N_14837,N_14516);
nor U15360 (N_15360,N_12552,N_12354);
nand U15361 (N_15361,N_14040,N_14585);
xnor U15362 (N_15362,N_14797,N_14155);
nor U15363 (N_15363,N_13489,N_14966);
nor U15364 (N_15364,N_12546,N_13563);
nand U15365 (N_15365,N_13122,N_12826);
nand U15366 (N_15366,N_14719,N_12598);
xor U15367 (N_15367,N_14200,N_12927);
nor U15368 (N_15368,N_14261,N_14663);
nand U15369 (N_15369,N_13583,N_13732);
nand U15370 (N_15370,N_12138,N_12619);
nor U15371 (N_15371,N_13947,N_13301);
or U15372 (N_15372,N_13638,N_14465);
or U15373 (N_15373,N_14394,N_12600);
or U15374 (N_15374,N_13869,N_14370);
xnor U15375 (N_15375,N_13221,N_12094);
or U15376 (N_15376,N_13230,N_12954);
nor U15377 (N_15377,N_13998,N_13432);
xnor U15378 (N_15378,N_13413,N_12831);
xor U15379 (N_15379,N_13967,N_13738);
nand U15380 (N_15380,N_14579,N_12839);
nand U15381 (N_15381,N_13286,N_13293);
xor U15382 (N_15382,N_12657,N_13401);
xnor U15383 (N_15383,N_13006,N_14460);
or U15384 (N_15384,N_13779,N_14806);
nor U15385 (N_15385,N_13590,N_13156);
nor U15386 (N_15386,N_13928,N_14174);
and U15387 (N_15387,N_12271,N_14983);
nor U15388 (N_15388,N_14808,N_12275);
nor U15389 (N_15389,N_14606,N_14392);
nor U15390 (N_15390,N_12941,N_12009);
and U15391 (N_15391,N_14423,N_14380);
or U15392 (N_15392,N_13019,N_14711);
and U15393 (N_15393,N_12820,N_14396);
or U15394 (N_15394,N_14232,N_13814);
or U15395 (N_15395,N_13518,N_13359);
or U15396 (N_15396,N_13035,N_13536);
xnor U15397 (N_15397,N_13776,N_14052);
nor U15398 (N_15398,N_14716,N_13077);
nand U15399 (N_15399,N_13456,N_14031);
and U15400 (N_15400,N_13427,N_12338);
xnor U15401 (N_15401,N_14127,N_13741);
nand U15402 (N_15402,N_13040,N_14385);
nor U15403 (N_15403,N_13767,N_12242);
nor U15404 (N_15404,N_13824,N_12045);
nand U15405 (N_15405,N_14096,N_13272);
nand U15406 (N_15406,N_12001,N_13449);
nor U15407 (N_15407,N_12007,N_14084);
nand U15408 (N_15408,N_14066,N_13434);
xor U15409 (N_15409,N_13943,N_14449);
or U15410 (N_15410,N_13544,N_14639);
and U15411 (N_15411,N_13801,N_12332);
nand U15412 (N_15412,N_14861,N_14725);
nand U15413 (N_15413,N_12168,N_14567);
or U15414 (N_15414,N_14877,N_12378);
nand U15415 (N_15415,N_13625,N_14827);
xor U15416 (N_15416,N_12772,N_14359);
and U15417 (N_15417,N_14773,N_13174);
and U15418 (N_15418,N_12478,N_14035);
and U15419 (N_15419,N_14166,N_13895);
or U15420 (N_15420,N_12621,N_12178);
nor U15421 (N_15421,N_13189,N_12698);
or U15422 (N_15422,N_12373,N_12167);
and U15423 (N_15423,N_12534,N_13596);
nand U15424 (N_15424,N_13740,N_12298);
and U15425 (N_15425,N_14779,N_13960);
nor U15426 (N_15426,N_13119,N_12917);
nand U15427 (N_15427,N_13103,N_14935);
nor U15428 (N_15428,N_12885,N_14027);
and U15429 (N_15429,N_12477,N_14430);
and U15430 (N_15430,N_12308,N_14830);
xnor U15431 (N_15431,N_12310,N_13971);
or U15432 (N_15432,N_13903,N_14334);
and U15433 (N_15433,N_14726,N_13579);
or U15434 (N_15434,N_12556,N_12819);
or U15435 (N_15435,N_13941,N_14535);
nor U15436 (N_15436,N_13212,N_12206);
nor U15437 (N_15437,N_13045,N_14865);
nand U15438 (N_15438,N_14499,N_14767);
or U15439 (N_15439,N_14018,N_14302);
nor U15440 (N_15440,N_13752,N_13707);
and U15441 (N_15441,N_13127,N_13249);
and U15442 (N_15442,N_14644,N_13458);
and U15443 (N_15443,N_12750,N_14691);
nor U15444 (N_15444,N_14750,N_13567);
nor U15445 (N_15445,N_13711,N_12545);
xor U15446 (N_15446,N_13134,N_12349);
nand U15447 (N_15447,N_14616,N_14871);
or U15448 (N_15448,N_14748,N_13609);
xor U15449 (N_15449,N_14440,N_14444);
nor U15450 (N_15450,N_13371,N_13244);
nor U15451 (N_15451,N_13237,N_14818);
and U15452 (N_15452,N_13521,N_13694);
nor U15453 (N_15453,N_12840,N_14512);
and U15454 (N_15454,N_13786,N_13584);
xnor U15455 (N_15455,N_12736,N_13558);
xor U15456 (N_15456,N_13440,N_12390);
nor U15457 (N_15457,N_12691,N_13268);
or U15458 (N_15458,N_13630,N_12978);
and U15459 (N_15459,N_14724,N_14993);
nand U15460 (N_15460,N_12925,N_14537);
and U15461 (N_15461,N_13139,N_14551);
nand U15462 (N_15462,N_14424,N_13113);
nand U15463 (N_15463,N_13246,N_13722);
nand U15464 (N_15464,N_13163,N_13522);
or U15465 (N_15465,N_12056,N_14319);
xor U15466 (N_15466,N_12089,N_14399);
nor U15467 (N_15467,N_12493,N_13345);
and U15468 (N_15468,N_13939,N_12547);
nand U15469 (N_15469,N_14742,N_14208);
or U15470 (N_15470,N_12209,N_12392);
or U15471 (N_15471,N_12335,N_14869);
xor U15472 (N_15472,N_12046,N_12553);
or U15473 (N_15473,N_12100,N_13041);
xor U15474 (N_15474,N_14958,N_12700);
xnor U15475 (N_15475,N_14580,N_14123);
nor U15476 (N_15476,N_14794,N_12472);
nand U15477 (N_15477,N_13735,N_12845);
and U15478 (N_15478,N_14624,N_14558);
or U15479 (N_15479,N_14336,N_14995);
and U15480 (N_15480,N_14160,N_12249);
nand U15481 (N_15481,N_13168,N_14685);
nand U15482 (N_15482,N_13390,N_12496);
or U15483 (N_15483,N_14901,N_14501);
or U15484 (N_15484,N_14504,N_12816);
xnor U15485 (N_15485,N_12821,N_14526);
nand U15486 (N_15486,N_12585,N_14408);
nand U15487 (N_15487,N_12503,N_13593);
xor U15488 (N_15488,N_12246,N_12295);
and U15489 (N_15489,N_14574,N_14407);
or U15490 (N_15490,N_12890,N_13130);
and U15491 (N_15491,N_12616,N_14836);
nor U15492 (N_15492,N_12199,N_14759);
nand U15493 (N_15493,N_13600,N_12764);
or U15494 (N_15494,N_13763,N_13676);
nor U15495 (N_15495,N_12906,N_12494);
xor U15496 (N_15496,N_12951,N_14793);
or U15497 (N_15497,N_13457,N_13995);
nand U15498 (N_15498,N_12303,N_13104);
xnor U15499 (N_15499,N_12918,N_12576);
nor U15500 (N_15500,N_12283,N_14792);
or U15501 (N_15501,N_14436,N_12237);
or U15502 (N_15502,N_14908,N_13601);
or U15503 (N_15503,N_13647,N_12184);
and U15504 (N_15504,N_12836,N_12144);
and U15505 (N_15505,N_14761,N_13184);
nor U15506 (N_15506,N_14932,N_13835);
nand U15507 (N_15507,N_14377,N_14876);
and U15508 (N_15508,N_14470,N_12562);
nor U15509 (N_15509,N_12030,N_14513);
nor U15510 (N_15510,N_14249,N_13396);
nand U15511 (N_15511,N_13655,N_13806);
or U15512 (N_15512,N_14689,N_14332);
and U15513 (N_15513,N_13677,N_13255);
nand U15514 (N_15514,N_12452,N_12969);
or U15515 (N_15515,N_12429,N_13905);
xor U15516 (N_15516,N_12858,N_12922);
xnor U15517 (N_15517,N_13724,N_12543);
nor U15518 (N_15518,N_14121,N_12882);
and U15519 (N_15519,N_12759,N_12187);
nand U15520 (N_15520,N_13355,N_12057);
nand U15521 (N_15521,N_13716,N_12614);
nor U15522 (N_15522,N_14219,N_13317);
or U15523 (N_15523,N_14250,N_13051);
and U15524 (N_15524,N_12312,N_13749);
nor U15525 (N_15525,N_13509,N_13240);
and U15526 (N_15526,N_13321,N_14735);
and U15527 (N_15527,N_14038,N_13602);
nand U15528 (N_15528,N_13911,N_14171);
or U15529 (N_15529,N_13242,N_12223);
and U15530 (N_15530,N_13453,N_14417);
and U15531 (N_15531,N_14197,N_13610);
nand U15532 (N_15532,N_13328,N_12139);
nor U15533 (N_15533,N_13053,N_13322);
or U15534 (N_15534,N_12709,N_14086);
or U15535 (N_15535,N_14265,N_12530);
nand U15536 (N_15536,N_14835,N_13860);
nand U15537 (N_15537,N_13845,N_14433);
nand U15538 (N_15538,N_12993,N_12911);
nand U15539 (N_15539,N_12339,N_12899);
or U15540 (N_15540,N_14144,N_14676);
xor U15541 (N_15541,N_12975,N_14894);
or U15542 (N_15542,N_14157,N_14651);
xnor U15543 (N_15543,N_13914,N_13410);
or U15544 (N_15544,N_14146,N_12641);
and U15545 (N_15545,N_14667,N_14952);
or U15546 (N_15546,N_12037,N_14431);
nor U15547 (N_15547,N_12897,N_12505);
xor U15548 (N_15548,N_14642,N_14177);
nand U15549 (N_15549,N_13565,N_12790);
and U15550 (N_15550,N_13169,N_13795);
xor U15551 (N_15551,N_13742,N_14071);
or U15552 (N_15552,N_14072,N_12549);
and U15553 (N_15553,N_14937,N_13442);
nand U15554 (N_15554,N_13825,N_13574);
xnor U15555 (N_15555,N_14391,N_14740);
xnor U15556 (N_15556,N_14496,N_14640);
or U15557 (N_15557,N_12259,N_14925);
nand U15558 (N_15558,N_12110,N_13199);
nor U15559 (N_15559,N_12182,N_13682);
nor U15560 (N_15560,N_12659,N_14520);
nand U15561 (N_15561,N_12256,N_13662);
and U15562 (N_15562,N_12667,N_12995);
nand U15563 (N_15563,N_14341,N_14786);
xnor U15564 (N_15564,N_12938,N_14170);
nor U15565 (N_15565,N_12524,N_14056);
or U15566 (N_15566,N_13818,N_13910);
and U15567 (N_15567,N_12824,N_14019);
xnor U15568 (N_15568,N_14137,N_12937);
and U15569 (N_15569,N_12835,N_13865);
nand U15570 (N_15570,N_13700,N_13887);
xnor U15571 (N_15571,N_14992,N_13498);
or U15572 (N_15572,N_14475,N_14409);
nor U15573 (N_15573,N_14075,N_14156);
nor U15574 (N_15574,N_13634,N_14154);
and U15575 (N_15575,N_14511,N_14820);
xnor U15576 (N_15576,N_13490,N_14706);
or U15577 (N_15577,N_12164,N_13699);
or U15578 (N_15578,N_12114,N_12487);
nor U15579 (N_15579,N_13871,N_14469);
nand U15580 (N_15580,N_13497,N_12127);
xnor U15581 (N_15581,N_12521,N_13531);
and U15582 (N_15582,N_14178,N_12610);
and U15583 (N_15583,N_14493,N_12797);
xnor U15584 (N_15584,N_14214,N_14324);
nor U15585 (N_15585,N_14209,N_12476);
and U15586 (N_15586,N_12471,N_12417);
xnor U15587 (N_15587,N_13670,N_12758);
xnor U15588 (N_15588,N_14213,N_12284);
xor U15589 (N_15589,N_13794,N_13266);
or U15590 (N_15590,N_14680,N_14057);
xnor U15591 (N_15591,N_12036,N_12498);
or U15592 (N_15592,N_14655,N_14351);
xnor U15593 (N_15593,N_13216,N_14968);
and U15594 (N_15594,N_13379,N_14848);
or U15595 (N_15595,N_14634,N_13916);
and U15596 (N_15596,N_12967,N_13897);
nor U15597 (N_15597,N_12142,N_13591);
and U15598 (N_15598,N_13131,N_12004);
nand U15599 (N_15599,N_12222,N_12763);
xor U15600 (N_15600,N_14743,N_14372);
nor U15601 (N_15601,N_14152,N_12314);
nor U15602 (N_15602,N_13493,N_13760);
or U15603 (N_15603,N_12742,N_14927);
and U15604 (N_15604,N_13263,N_14450);
nand U15605 (N_15605,N_12287,N_12664);
nor U15606 (N_15606,N_12702,N_14173);
or U15607 (N_15607,N_12919,N_13276);
nand U15608 (N_15608,N_13494,N_14856);
or U15609 (N_15609,N_12722,N_14106);
nor U15610 (N_15610,N_14813,N_12082);
nand U15611 (N_15611,N_13836,N_14690);
and U15612 (N_15612,N_12343,N_13210);
nand U15613 (N_15613,N_13049,N_13505);
xnor U15614 (N_15614,N_14037,N_13823);
nand U15615 (N_15615,N_12915,N_14886);
nor U15616 (N_15616,N_12930,N_12410);
nor U15617 (N_15617,N_12893,N_13979);
xor U15618 (N_15618,N_14013,N_12300);
or U15619 (N_15619,N_12724,N_14868);
and U15620 (N_15620,N_12583,N_13628);
or U15621 (N_15621,N_12328,N_12853);
nor U15622 (N_15622,N_12306,N_12490);
xor U15623 (N_15623,N_14789,N_13966);
xor U15624 (N_15624,N_13478,N_13471);
or U15625 (N_15625,N_12152,N_13406);
nor U15626 (N_15626,N_12788,N_13855);
nor U15627 (N_15627,N_13452,N_13920);
nand U15628 (N_15628,N_14487,N_12843);
xor U15629 (N_15629,N_12155,N_14531);
or U15630 (N_15630,N_14024,N_12638);
and U15631 (N_15631,N_14122,N_14212);
or U15632 (N_15632,N_14234,N_14939);
nand U15633 (N_15633,N_12623,N_13022);
xor U15634 (N_15634,N_14055,N_12385);
and U15635 (N_15635,N_13793,N_12215);
or U15636 (N_15636,N_13037,N_12544);
nor U15637 (N_15637,N_13172,N_14621);
and U15638 (N_15638,N_12589,N_13152);
nor U15639 (N_15639,N_13061,N_14984);
and U15640 (N_15640,N_14432,N_14422);
nand U15641 (N_15641,N_12247,N_12445);
nand U15642 (N_15642,N_14822,N_12860);
or U15643 (N_15643,N_12267,N_13179);
nor U15644 (N_15644,N_12959,N_14682);
and U15645 (N_15645,N_14674,N_14389);
or U15646 (N_15646,N_13146,N_13927);
and U15647 (N_15647,N_12704,N_14179);
xnor U15648 (N_15648,N_12696,N_12066);
nor U15649 (N_15649,N_12609,N_12109);
xor U15650 (N_15650,N_14903,N_13063);
or U15651 (N_15651,N_14172,N_12250);
nand U15652 (N_15652,N_12877,N_12923);
xnor U15653 (N_15653,N_12712,N_14479);
nor U15654 (N_15654,N_13310,N_14653);
xor U15655 (N_15655,N_13788,N_13649);
nand U15656 (N_15656,N_12186,N_12693);
or U15657 (N_15657,N_12122,N_14731);
xnor U15658 (N_15658,N_14804,N_12730);
and U15659 (N_15659,N_14393,N_12239);
or U15660 (N_15660,N_13624,N_14814);
nor U15661 (N_15661,N_13429,N_14196);
nor U15662 (N_15662,N_12289,N_12262);
nor U15663 (N_15663,N_14306,N_13042);
or U15664 (N_15664,N_14238,N_13578);
xnor U15665 (N_15665,N_14453,N_12176);
nor U15666 (N_15666,N_12361,N_13397);
and U15667 (N_15667,N_13688,N_12039);
xnor U15668 (N_15668,N_13472,N_14972);
or U15669 (N_15669,N_12855,N_12594);
nor U15670 (N_15670,N_12140,N_14042);
xnor U15671 (N_15671,N_12968,N_12117);
nand U15672 (N_15672,N_12952,N_13560);
and U15673 (N_15673,N_13392,N_12369);
and U15674 (N_15674,N_14349,N_14705);
and U15675 (N_15675,N_14026,N_12755);
xor U15676 (N_15676,N_13693,N_13968);
xnor U15677 (N_15677,N_12658,N_12033);
and U15678 (N_15678,N_12019,N_12912);
and U15679 (N_15679,N_13181,N_12901);
or U15680 (N_15680,N_14204,N_14117);
and U15681 (N_15681,N_12462,N_13068);
or U15682 (N_15682,N_13349,N_14322);
nand U15683 (N_15683,N_14641,N_14978);
nand U15684 (N_15684,N_14796,N_14227);
xor U15685 (N_15685,N_14229,N_14605);
nor U15686 (N_15686,N_13804,N_12540);
nor U15687 (N_15687,N_14546,N_13926);
nor U15688 (N_15688,N_12612,N_14044);
and U15689 (N_15689,N_13519,N_14330);
nand U15690 (N_15690,N_14525,N_13753);
nor U15691 (N_15691,N_14583,N_13768);
xnor U15692 (N_15692,N_14458,N_13849);
or U15693 (N_15693,N_13380,N_14147);
nand U15694 (N_15694,N_14490,N_13710);
nor U15695 (N_15695,N_12814,N_14863);
nand U15696 (N_15696,N_12636,N_12774);
xor U15697 (N_15697,N_13363,N_13718);
xnor U15698 (N_15698,N_12285,N_12273);
xnor U15699 (N_15699,N_13870,N_12292);
or U15700 (N_15700,N_14961,N_14126);
or U15701 (N_15701,N_12277,N_13781);
nand U15702 (N_15702,N_12958,N_13510);
nand U15703 (N_15703,N_14981,N_13353);
nand U15704 (N_15704,N_14198,N_13100);
or U15705 (N_15705,N_13907,N_13358);
xnor U15706 (N_15706,N_13956,N_14573);
and U15707 (N_15707,N_12086,N_12555);
nand U15708 (N_15708,N_14571,N_13306);
or U15709 (N_15709,N_14190,N_13347);
nor U15710 (N_15710,N_14694,N_14887);
nand U15711 (N_15711,N_13102,N_12980);
nor U15712 (N_15712,N_12404,N_12096);
or U15713 (N_15713,N_12745,N_12678);
nor U15714 (N_15714,N_14262,N_12427);
nor U15715 (N_15715,N_12977,N_14819);
and U15716 (N_15716,N_12723,N_13502);
xnor U15717 (N_15717,N_13260,N_14845);
nor U15718 (N_15718,N_13454,N_14870);
xnor U15719 (N_15719,N_13479,N_12304);
and U15720 (N_15720,N_12832,N_12217);
xor U15721 (N_15721,N_14548,N_13878);
nor U15722 (N_15722,N_12972,N_12166);
and U15723 (N_15723,N_14781,N_12634);
nor U15724 (N_15724,N_12561,N_12838);
xor U15725 (N_15725,N_14661,N_14000);
xnor U15726 (N_15726,N_14455,N_14283);
nor U15727 (N_15727,N_14326,N_12714);
or U15728 (N_15728,N_13946,N_12675);
xnor U15729 (N_15729,N_13996,N_13274);
and U15730 (N_15730,N_13043,N_14464);
and U15731 (N_15731,N_14638,N_12602);
or U15732 (N_15732,N_14437,N_13704);
nand U15733 (N_15733,N_12684,N_13972);
nor U15734 (N_15734,N_13615,N_14866);
nor U15735 (N_15735,N_13316,N_14405);
xor U15736 (N_15736,N_13252,N_12098);
nand U15737 (N_15737,N_13790,N_14660);
xor U15738 (N_15738,N_12856,N_13807);
and U15739 (N_15739,N_13389,N_14603);
nor U15740 (N_15740,N_13046,N_13962);
nand U15741 (N_15741,N_14798,N_12740);
nor U15742 (N_15742,N_13298,N_12203);
xnor U15743 (N_15743,N_13517,N_12428);
and U15744 (N_15744,N_14308,N_13538);
nor U15745 (N_15745,N_12113,N_14555);
or U15746 (N_15746,N_12999,N_12034);
nor U15747 (N_15747,N_14505,N_14693);
nand U15748 (N_15748,N_12252,N_13304);
or U15749 (N_15749,N_14560,N_14936);
and U15750 (N_15750,N_14045,N_13313);
nand U15751 (N_15751,N_12637,N_14246);
nor U15752 (N_15752,N_14061,N_13712);
xor U15753 (N_15753,N_14539,N_12147);
nand U15754 (N_15754,N_14540,N_14082);
nand U15755 (N_15755,N_14649,N_13585);
nor U15756 (N_15756,N_12640,N_13036);
xnor U15757 (N_15757,N_13702,N_14924);
and U15758 (N_15758,N_14787,N_12372);
or U15759 (N_15759,N_13889,N_14017);
nand U15760 (N_15760,N_12055,N_14379);
nor U15761 (N_15761,N_14451,N_12847);
xnor U15762 (N_15762,N_14167,N_12067);
and U15763 (N_15763,N_12558,N_14594);
or U15764 (N_15764,N_14622,N_14272);
nor U15765 (N_15765,N_14950,N_12351);
or U15766 (N_15766,N_13898,N_12425);
xor U15767 (N_15767,N_14976,N_14559);
xor U15768 (N_15768,N_14878,N_14447);
nand U15769 (N_15769,N_12111,N_13674);
nand U15770 (N_15770,N_12731,N_12575);
nor U15771 (N_15771,N_14011,N_14148);
or U15772 (N_15772,N_13299,N_14080);
nand U15773 (N_15773,N_12299,N_14698);
and U15774 (N_15774,N_13430,N_13799);
or U15775 (N_15775,N_12531,N_12936);
or U15776 (N_15776,N_14506,N_12419);
or U15777 (N_15777,N_12017,N_13561);
xor U15778 (N_15778,N_14918,N_13492);
nand U15779 (N_15779,N_13384,N_12817);
nand U15780 (N_15780,N_14647,N_12133);
nand U15781 (N_15781,N_14268,N_14221);
nor U15782 (N_15782,N_14373,N_14254);
nor U15783 (N_15783,N_12883,N_13888);
or U15784 (N_15784,N_13843,N_14313);
and U15785 (N_15785,N_13029,N_13350);
xor U15786 (N_15786,N_14260,N_13106);
and U15787 (N_15787,N_13476,N_14826);
nor U15788 (N_15788,N_13775,N_12050);
nor U15789 (N_15789,N_12907,N_12929);
xor U15790 (N_15790,N_12669,N_12560);
nand U15791 (N_15791,N_13437,N_14615);
or U15792 (N_15792,N_14001,N_14846);
nand U15793 (N_15793,N_14847,N_12830);
nor U15794 (N_15794,N_14824,N_12770);
xnor U15795 (N_15795,N_14832,N_14628);
or U15796 (N_15796,N_14376,N_12673);
nand U15797 (N_15797,N_13066,N_12364);
nor U15798 (N_15798,N_14180,N_12000);
nand U15799 (N_15799,N_14059,N_12420);
xor U15800 (N_15800,N_13524,N_13342);
xor U15801 (N_15801,N_13483,N_14305);
nand U15802 (N_15802,N_14107,N_14356);
and U15803 (N_15803,N_14400,N_12587);
xor U15804 (N_15804,N_14226,N_12596);
nor U15805 (N_15805,N_12291,N_14087);
and U15806 (N_15806,N_13566,N_13653);
or U15807 (N_15807,N_14347,N_12235);
nor U15808 (N_15808,N_12336,N_14996);
or U15809 (N_15809,N_13936,N_12728);
or U15810 (N_15810,N_13839,N_12353);
nand U15811 (N_15811,N_14098,N_12608);
and U15812 (N_15812,N_13713,N_13279);
and U15813 (N_15813,N_14012,N_14713);
or U15814 (N_15814,N_13076,N_13195);
and U15815 (N_15815,N_14350,N_12992);
nor U15816 (N_15816,N_13506,N_13238);
or U15817 (N_15817,N_12486,N_13394);
nand U15818 (N_15818,N_14600,N_12473);
xor U15819 (N_15819,N_13114,N_12099);
nand U15820 (N_15820,N_14695,N_13696);
and U15821 (N_15821,N_14348,N_14550);
nor U15822 (N_15822,N_13198,N_12251);
or U15823 (N_15823,N_14707,N_12108);
or U15824 (N_15824,N_14029,N_14175);
xnor U15825 (N_15825,N_14849,N_13886);
xnor U15826 (N_15826,N_13128,N_14947);
xnor U15827 (N_15827,N_14093,N_14129);
or U15828 (N_15828,N_13772,N_14083);
nand U15829 (N_15829,N_13523,N_12802);
xnor U15830 (N_15830,N_14471,N_12465);
nor U15831 (N_15831,N_12485,N_14563);
nor U15832 (N_15832,N_13346,N_12551);
and U15833 (N_15833,N_12953,N_12573);
nor U15834 (N_15834,N_14771,N_13351);
xor U15835 (N_15835,N_14589,N_12976);
xnor U15836 (N_15836,N_13415,N_13842);
or U15837 (N_15837,N_12406,N_13110);
xor U15838 (N_15838,N_12460,N_13901);
and U15839 (N_15839,N_12861,N_13269);
nand U15840 (N_15840,N_14327,N_12935);
xor U15841 (N_15841,N_12044,N_13026);
or U15842 (N_15842,N_13157,N_13287);
nand U15843 (N_15843,N_12595,N_13013);
nand U15844 (N_15844,N_12020,N_14090);
or U15845 (N_15845,N_14388,N_14552);
nor U15846 (N_15846,N_14269,N_14545);
and U15847 (N_15847,N_12985,N_13455);
or U15848 (N_15848,N_13099,N_13402);
or U15849 (N_15849,N_14151,N_12630);
or U15850 (N_15850,N_12571,N_13892);
xnor U15851 (N_15851,N_14970,N_14374);
or U15852 (N_15852,N_14554,N_12776);
or U15853 (N_15853,N_14769,N_14933);
nor U15854 (N_15854,N_12450,N_12618);
xnor U15855 (N_15855,N_14163,N_13894);
and U15856 (N_15856,N_13426,N_12381);
nor U15857 (N_15857,N_14623,N_14625);
nand U15858 (N_15858,N_12356,N_12757);
nor U15859 (N_15859,N_13308,N_13209);
nor U15860 (N_15860,N_13239,N_13819);
nor U15861 (N_15861,N_13658,N_12689);
xnor U15862 (N_15862,N_14979,N_14194);
and U15863 (N_15863,N_14244,N_12068);
or U15864 (N_15864,N_14687,N_12132);
xnor U15865 (N_15865,N_14785,N_14192);
nand U15866 (N_15866,N_12987,N_13656);
xor U15867 (N_15867,N_13448,N_14755);
nand U15868 (N_15868,N_13654,N_13867);
or U15869 (N_15869,N_14412,N_13213);
nor U15870 (N_15870,N_13441,N_13679);
xnor U15871 (N_15871,N_12871,N_13320);
xor U15872 (N_15872,N_13838,N_12377);
or U15873 (N_15873,N_14790,N_14646);
and U15874 (N_15874,N_14954,N_13101);
xnor U15875 (N_15875,N_13617,N_13540);
and U15876 (N_15876,N_12970,N_12933);
and U15877 (N_15877,N_13248,N_14369);
xnor U15878 (N_15878,N_13142,N_14570);
xor U15879 (N_15879,N_13520,N_14366);
nand U15880 (N_15880,N_12479,N_12307);
or U15881 (N_15881,N_14414,N_13292);
nand U15882 (N_15882,N_12038,N_14746);
and U15883 (N_15883,N_12032,N_13754);
nor U15884 (N_15884,N_13190,N_12844);
nand U15885 (N_15885,N_14406,N_13832);
or U15886 (N_15886,N_13873,N_14216);
or U15887 (N_15887,N_12829,N_12363);
or U15888 (N_15888,N_12867,N_14772);
or U15889 (N_15889,N_12957,N_14115);
xor U15890 (N_15890,N_14760,N_12718);
or U15891 (N_15891,N_12994,N_13974);
nand U15892 (N_15892,N_13616,N_14951);
xnor U15893 (N_15893,N_12394,N_12566);
nand U15894 (N_15894,N_14517,N_12644);
nor U15895 (N_15895,N_12683,N_13765);
nor U15896 (N_15896,N_12559,N_14757);
nand U15897 (N_15897,N_12455,N_13047);
and U15898 (N_15898,N_13828,N_13253);
and U15899 (N_15899,N_13009,N_14710);
nand U15900 (N_15900,N_14404,N_12451);
and U15901 (N_15901,N_14657,N_14312);
xnor U15902 (N_15902,N_14562,N_13329);
nand U15903 (N_15903,N_13087,N_13862);
nand U15904 (N_15904,N_14242,N_13123);
nor U15905 (N_15905,N_13729,N_13291);
xnor U15906 (N_15906,N_14342,N_12727);
xnor U15907 (N_15907,N_13988,N_13612);
nor U15908 (N_15908,N_14425,N_12532);
and U15909 (N_15909,N_14145,N_13539);
and U15910 (N_15910,N_13672,N_12131);
nor U15911 (N_15911,N_13952,N_13599);
xnor U15912 (N_15912,N_14131,N_12200);
or U15913 (N_15913,N_14881,N_12864);
nor U15914 (N_15914,N_12454,N_12665);
xor U15915 (N_15915,N_13425,N_14920);
nor U15916 (N_15916,N_12129,N_13495);
nor U15917 (N_15917,N_14135,N_13534);
nand U15918 (N_15918,N_13983,N_12701);
nand U15919 (N_15919,N_12270,N_14909);
xnor U15920 (N_15920,N_12866,N_13245);
nand U15921 (N_15921,N_12391,N_12685);
or U15922 (N_15922,N_14294,N_14049);
xor U15923 (N_15923,N_12238,N_12063);
nand U15924 (N_15924,N_12811,N_14318);
or U15925 (N_15925,N_14295,N_12650);
xnor U15926 (N_15926,N_12660,N_13553);
nor U15927 (N_15927,N_12516,N_14588);
nor U15928 (N_15928,N_14611,N_14235);
or U15929 (N_15929,N_12225,N_13993);
xor U15930 (N_15930,N_13261,N_12286);
and U15931 (N_15931,N_12426,N_12510);
and U15932 (N_15932,N_14709,N_13844);
and U15933 (N_15933,N_14977,N_13052);
nor U15934 (N_15934,N_14275,N_12859);
and U15935 (N_15935,N_12956,N_12949);
xor U15936 (N_15936,N_13607,N_14784);
nor U15937 (N_15937,N_13005,N_12813);
nand U15938 (N_15938,N_13929,N_12613);
or U15939 (N_15939,N_14124,N_12646);
or U15940 (N_15940,N_13003,N_12964);
and U15941 (N_15941,N_14142,N_14480);
and U15942 (N_15942,N_13629,N_13909);
nor U15943 (N_15943,N_12779,N_12398);
xnor U15944 (N_15944,N_13613,N_14852);
nor U15945 (N_15945,N_12464,N_13296);
nor U15946 (N_15946,N_14182,N_14411);
nor U15947 (N_15947,N_13133,N_14672);
nand U15948 (N_15948,N_13800,N_14053);
or U15949 (N_15949,N_14454,N_13529);
nor U15950 (N_15950,N_14897,N_14959);
xor U15951 (N_15951,N_14811,N_14883);
and U15952 (N_15952,N_13528,N_12075);
nand U15953 (N_15953,N_13734,N_13154);
and U15954 (N_15954,N_13354,N_12799);
nand U15955 (N_15955,N_12565,N_14002);
xor U15956 (N_15956,N_12218,N_13148);
nor U15957 (N_15957,N_13211,N_14764);
or U15958 (N_15958,N_14921,N_13516);
nand U15959 (N_15959,N_12396,N_13572);
nand U15960 (N_15960,N_13004,N_12924);
nor U15961 (N_15961,N_12990,N_13404);
and U15962 (N_15962,N_13258,N_13141);
and U15963 (N_15963,N_14782,N_14073);
or U15964 (N_15964,N_13079,N_14875);
and U15965 (N_15965,N_14980,N_12124);
xnor U15966 (N_15966,N_12795,N_13194);
or U15967 (N_15967,N_13771,N_12896);
nand U15968 (N_15968,N_14557,N_13098);
nor U15969 (N_15969,N_13094,N_13391);
nand U15970 (N_15970,N_14749,N_13868);
nand U15971 (N_15971,N_12097,N_14236);
nor U15972 (N_15972,N_12204,N_14291);
xor U15973 (N_15973,N_14102,N_13474);
and U15974 (N_15974,N_14252,N_12344);
and U15975 (N_15975,N_12680,N_13743);
xnor U15976 (N_15976,N_14770,N_14700);
nand U15977 (N_15977,N_14697,N_14645);
or U15978 (N_15978,N_12210,N_13748);
nand U15979 (N_15979,N_12651,N_14285);
or U15980 (N_15980,N_13020,N_14111);
nor U15981 (N_15981,N_14344,N_12023);
and U15982 (N_15982,N_13065,N_14279);
and U15983 (N_15983,N_13791,N_12288);
nand U15984 (N_15984,N_13745,N_14067);
or U15985 (N_15985,N_12264,N_14415);
and U15986 (N_15986,N_14094,N_13105);
nand U15987 (N_15987,N_13167,N_12668);
or U15988 (N_15988,N_13935,N_12422);
xnor U15989 (N_15989,N_13236,N_14228);
or U15990 (N_15990,N_13594,N_14762);
nand U15991 (N_15991,N_12647,N_14337);
xor U15992 (N_15992,N_12777,N_13964);
nor U15993 (N_15993,N_12783,N_12894);
nand U15994 (N_15994,N_13487,N_13731);
nand U15995 (N_15995,N_12162,N_14032);
nor U15996 (N_15996,N_12322,N_12070);
nand U15997 (N_15997,N_13933,N_12318);
xnor U15998 (N_15998,N_12852,N_14378);
and U15999 (N_15999,N_12330,N_14823);
nor U16000 (N_16000,N_12360,N_13182);
and U16001 (N_16001,N_14833,N_14816);
nand U16002 (N_16002,N_12165,N_14938);
nor U16003 (N_16003,N_13526,N_14008);
nand U16004 (N_16004,N_13340,N_14335);
or U16005 (N_16005,N_14592,N_14728);
nand U16006 (N_16006,N_13300,N_13782);
nand U16007 (N_16007,N_13527,N_14482);
xor U16008 (N_16008,N_13537,N_12402);
xnor U16009 (N_16009,N_14896,N_14485);
xor U16010 (N_16010,N_13550,N_13136);
xnor U16011 (N_16011,N_12841,N_12407);
nor U16012 (N_16012,N_13232,N_12463);
nor U16013 (N_16013,N_13697,N_14481);
and U16014 (N_16014,N_13436,N_14768);
nand U16015 (N_16015,N_12386,N_14210);
or U16016 (N_16016,N_13259,N_12158);
or U16017 (N_16017,N_14890,N_12205);
nand U16018 (N_16018,N_14357,N_14945);
nor U16019 (N_16019,N_13689,N_14099);
nor U16020 (N_16020,N_12123,N_14668);
xor U16021 (N_16021,N_12920,N_14401);
and U16022 (N_16022,N_14028,N_12948);
xnor U16023 (N_16023,N_12430,N_12528);
nand U16024 (N_16024,N_13398,N_14101);
nor U16025 (N_16025,N_13348,N_14266);
and U16026 (N_16026,N_14917,N_12090);
nor U16027 (N_16027,N_12662,N_14696);
and U16028 (N_16028,N_14446,N_13706);
xor U16029 (N_16029,N_14503,N_14429);
nand U16030 (N_16030,N_13153,N_12347);
nor U16031 (N_16031,N_14006,N_13635);
xor U16032 (N_16032,N_13940,N_12940);
xnor U16033 (N_16033,N_12232,N_13024);
nor U16034 (N_16034,N_12265,N_14274);
or U16035 (N_16035,N_13038,N_12787);
or U16036 (N_16036,N_13370,N_14608);
and U16037 (N_16037,N_14258,N_13883);
xnor U16038 (N_16038,N_12495,N_12188);
xor U16039 (N_16039,N_12707,N_14134);
or U16040 (N_16040,N_14577,N_12766);
nand U16041 (N_16041,N_14005,N_14765);
xor U16042 (N_16042,N_14021,N_12697);
xor U16043 (N_16043,N_14325,N_14119);
nand U16044 (N_16044,N_13780,N_12077);
xor U16045 (N_16045,N_14684,N_14333);
and U16046 (N_16046,N_13783,N_14681);
and U16047 (N_16047,N_13675,N_12726);
or U16048 (N_16048,N_12380,N_13874);
nand U16049 (N_16049,N_14010,N_14445);
or U16050 (N_16050,N_14944,N_13508);
and U16051 (N_16051,N_12141,N_14753);
nand U16052 (N_16052,N_14928,N_14114);
nor U16053 (N_16053,N_13661,N_14105);
nor U16054 (N_16054,N_12692,N_14683);
nor U16055 (N_16055,N_13923,N_14542);
nand U16056 (N_16056,N_13481,N_14109);
nand U16057 (N_16057,N_12567,N_12499);
nor U16058 (N_16058,N_12183,N_13459);
and U16059 (N_16059,N_13975,N_13496);
nand U16060 (N_16060,N_12058,N_14508);
nand U16061 (N_16061,N_12230,N_14733);
nand U16062 (N_16062,N_14662,N_13164);
and U16063 (N_16063,N_14287,N_13222);
or U16064 (N_16064,N_12973,N_14879);
and U16065 (N_16065,N_13552,N_12997);
nand U16066 (N_16066,N_13294,N_13737);
or U16067 (N_16067,N_13284,N_12775);
nor U16068 (N_16068,N_14854,N_12311);
xnor U16069 (N_16069,N_12340,N_12822);
nor U16070 (N_16070,N_14161,N_14590);
nor U16071 (N_16071,N_12904,N_12172);
xnor U16072 (N_16072,N_13973,N_13374);
or U16073 (N_16073,N_12942,N_13031);
nor U16074 (N_16074,N_13149,N_13271);
xnor U16075 (N_16075,N_13204,N_13646);
xnor U16076 (N_16076,N_13631,N_13627);
xor U16077 (N_16077,N_14678,N_13140);
xnor U16078 (N_16078,N_13853,N_14889);
xnor U16079 (N_16079,N_14810,N_13683);
and U16080 (N_16080,N_12095,N_12554);
or U16081 (N_16081,N_12512,N_13290);
nor U16082 (N_16082,N_13931,N_12881);
nor U16083 (N_16083,N_14635,N_12069);
nor U16084 (N_16084,N_13385,N_12119);
and U16085 (N_16085,N_14509,N_13097);
nand U16086 (N_16086,N_13201,N_13681);
or U16087 (N_16087,N_12501,N_13176);
nand U16088 (N_16088,N_14686,N_13991);
nand U16089 (N_16089,N_14329,N_13709);
xor U16090 (N_16090,N_14193,N_14860);
xor U16091 (N_16091,N_12418,N_12828);
nor U16092 (N_16092,N_12320,N_14841);
nor U16093 (N_16093,N_12888,N_13409);
nand U16094 (N_16094,N_13405,N_14108);
xnor U16095 (N_16095,N_12761,N_12946);
and U16096 (N_16096,N_13407,N_14463);
nand U16097 (N_16097,N_13667,N_14533);
nand U16098 (N_16098,N_14544,N_12389);
xnor U16099 (N_16099,N_12635,N_13357);
nor U16100 (N_16100,N_14140,N_14780);
nand U16101 (N_16101,N_14340,N_14128);
nand U16102 (N_16102,N_12245,N_12234);
xor U16103 (N_16103,N_14352,N_13018);
and U16104 (N_16104,N_12523,N_14181);
nor U16105 (N_16105,N_12157,N_13543);
xnor U16106 (N_16106,N_12189,N_13175);
or U16107 (N_16107,N_13751,N_14375);
or U16108 (N_16108,N_14991,N_13932);
nand U16109 (N_16109,N_12281,N_13491);
xor U16110 (N_16110,N_12076,N_14164);
or U16111 (N_16111,N_12366,N_12241);
and U16112 (N_16112,N_14165,N_14536);
nand U16113 (N_16113,N_14158,N_13382);
nand U16114 (N_16114,N_14990,N_13719);
nor U16115 (N_16115,N_13650,N_14328);
or U16116 (N_16116,N_14842,N_14466);
nand U16117 (N_16117,N_12533,N_14477);
and U16118 (N_16118,N_13295,N_13419);
and U16119 (N_16119,N_13588,N_13424);
nand U16120 (N_16120,N_12713,N_13755);
xor U16121 (N_16121,N_13809,N_12491);
and U16122 (N_16122,N_12201,N_12753);
xor U16123 (N_16123,N_12156,N_13057);
or U16124 (N_16124,N_12519,N_14297);
or U16125 (N_16125,N_13473,N_12807);
nand U16126 (N_16126,N_14572,N_14613);
and U16127 (N_16127,N_13852,N_13817);
nand U16128 (N_16128,N_12803,N_13854);
and U16129 (N_16129,N_12916,N_12649);
xor U16130 (N_16130,N_13075,N_13107);
nand U16131 (N_16131,N_12642,N_12350);
and U16132 (N_16132,N_12088,N_13257);
nand U16133 (N_16133,N_14483,N_13319);
or U16134 (N_16134,N_13183,N_13125);
nor U16135 (N_16135,N_12072,N_13810);
nand U16136 (N_16136,N_12226,N_12442);
nand U16137 (N_16137,N_12459,N_14568);
nor U16138 (N_16138,N_14888,N_14817);
xnor U16139 (N_16139,N_12087,N_12903);
xor U16140 (N_16140,N_12049,N_13826);
or U16141 (N_16141,N_14365,N_13469);
or U16142 (N_16142,N_13792,N_14679);
nand U16143 (N_16143,N_13403,N_12054);
nor U16144 (N_16144,N_12760,N_12971);
xor U16145 (N_16145,N_13922,N_13017);
or U16146 (N_16146,N_14478,N_12898);
and U16147 (N_16147,N_14839,N_13421);
xor U16148 (N_16148,N_13050,N_12432);
and U16149 (N_16149,N_12107,N_14741);
or U16150 (N_16150,N_13987,N_14859);
nand U16151 (N_16151,N_12805,N_12672);
and U16152 (N_16152,N_12433,N_14320);
and U16153 (N_16153,N_13980,N_12765);
and U16154 (N_16154,N_13690,N_12342);
nand U16155 (N_16155,N_14727,N_14263);
and U16156 (N_16156,N_12006,N_14434);
nor U16157 (N_16157,N_12507,N_12511);
and U16158 (N_16158,N_12509,N_13265);
and U16159 (N_16159,N_12145,N_13504);
xor U16160 (N_16160,N_12305,N_12468);
nor U16161 (N_16161,N_14617,N_14468);
nand U16162 (N_16162,N_13081,N_14882);
and U16163 (N_16163,N_13067,N_14143);
or U16164 (N_16164,N_12902,N_12751);
xnor U16165 (N_16165,N_12074,N_13603);
or U16166 (N_16166,N_14941,N_12012);
or U16167 (N_16167,N_13285,N_12458);
or U16168 (N_16168,N_14220,N_14926);
nor U16169 (N_16169,N_12027,N_12934);
or U16170 (N_16170,N_14462,N_14704);
nand U16171 (N_16171,N_13135,N_14632);
nand U16172 (N_16172,N_13435,N_13698);
or U16173 (N_16173,N_13937,N_13444);
nor U16174 (N_16174,N_14994,N_14522);
xnor U16175 (N_16175,N_12617,N_13581);
or U16176 (N_16176,N_12564,N_12083);
or U16177 (N_16177,N_12791,N_13088);
or U16178 (N_16178,N_12842,N_14296);
or U16179 (N_16179,N_14104,N_12244);
xor U16180 (N_16180,N_14795,N_13821);
nand U16181 (N_16181,N_14292,N_12639);
and U16182 (N_16182,N_12125,N_12931);
and U16183 (N_16183,N_12579,N_12804);
and U16184 (N_16184,N_14648,N_14598);
and U16185 (N_16185,N_13803,N_14650);
nand U16186 (N_16186,N_12529,N_14677);
and U16187 (N_16187,N_14435,N_14652);
nor U16188 (N_16188,N_12093,N_12003);
nor U16189 (N_16189,N_13048,N_14230);
and U16190 (N_16190,N_14576,N_12815);
nand U16191 (N_16191,N_13945,N_12932);
xnor U16192 (N_16192,N_14402,N_12748);
nand U16193 (N_16193,N_13577,N_14971);
and U16194 (N_16194,N_14081,N_14293);
or U16195 (N_16195,N_13893,N_13145);
nor U16196 (N_16196,N_13500,N_12747);
and U16197 (N_16197,N_13766,N_12862);
and U16198 (N_16198,N_13950,N_14829);
nor U16199 (N_16199,N_12808,N_13648);
and U16200 (N_16200,N_12928,N_12653);
nand U16201 (N_16201,N_14241,N_14088);
nand U16202 (N_16202,N_12213,N_12008);
nand U16203 (N_16203,N_14601,N_13717);
or U16204 (N_16204,N_13595,N_13034);
or U16205 (N_16205,N_12752,N_13461);
or U16206 (N_16206,N_14802,N_13863);
and U16207 (N_16207,N_14183,N_13021);
nand U16208 (N_16208,N_13721,N_12785);
xnor U16209 (N_16209,N_12319,N_12720);
xor U16210 (N_16210,N_13597,N_13090);
xor U16211 (N_16211,N_12071,N_13637);
or U16212 (N_16212,N_12357,N_14381);
nor U16213 (N_16213,N_14666,N_12632);
or U16214 (N_16214,N_12443,N_14076);
or U16215 (N_16215,N_12670,N_12475);
nand U16216 (N_16216,N_13501,N_13173);
nor U16217 (N_16217,N_13229,N_13341);
or U16218 (N_16218,N_14549,N_14077);
or U16219 (N_16219,N_12857,N_12367);
and U16220 (N_16220,N_12873,N_13362);
and U16221 (N_16221,N_13438,N_12801);
nor U16222 (N_16222,N_12989,N_14702);
or U16223 (N_16223,N_12663,N_14530);
nand U16224 (N_16224,N_12102,N_14064);
xor U16225 (N_16225,N_13533,N_14284);
nand U16226 (N_16226,N_12593,N_13278);
xnor U16227 (N_16227,N_12280,N_13598);
or U16228 (N_16228,N_13875,N_14873);
or U16229 (N_16229,N_14133,N_12352);
nand U16230 (N_16230,N_13147,N_14930);
nand U16231 (N_16231,N_12800,N_13884);
and U16232 (N_16232,N_12687,N_12048);
xor U16233 (N_16233,N_12078,N_13002);
nand U16234 (N_16234,N_12615,N_14999);
or U16235 (N_16235,N_14729,N_12233);
nor U16236 (N_16236,N_12588,N_13576);
and U16237 (N_16237,N_12947,N_13012);
or U16238 (N_16238,N_13383,N_14627);
xor U16239 (N_16239,N_14368,N_13750);
or U16240 (N_16240,N_13770,N_13728);
nand U16241 (N_16241,N_14956,N_14395);
xor U16242 (N_16242,N_14253,N_14528);
or U16243 (N_16243,N_14607,N_13640);
or U16244 (N_16244,N_13666,N_14338);
and U16245 (N_16245,N_14614,N_14439);
or U16246 (N_16246,N_14739,N_13606);
nor U16247 (N_16247,N_12026,N_14343);
and U16248 (N_16248,N_13283,N_14636);
or U16249 (N_16249,N_13507,N_13256);
or U16250 (N_16250,N_12900,N_12316);
or U16251 (N_16251,N_14421,N_13247);
nand U16252 (N_16252,N_13335,N_14256);
xnor U16253 (N_16253,N_12601,N_14311);
nand U16254 (N_16254,N_12648,N_13251);
and U16255 (N_16255,N_14240,N_14051);
nand U16256 (N_16256,N_14543,N_12502);
or U16257 (N_16257,N_13921,N_12744);
or U16258 (N_16258,N_13769,N_14063);
and U16259 (N_16259,N_12984,N_13369);
or U16260 (N_16260,N_14428,N_12739);
or U16261 (N_16261,N_12212,N_12582);
nand U16262 (N_16262,N_13010,N_14113);
nor U16263 (N_16263,N_13331,N_12444);
and U16264 (N_16264,N_12368,N_14218);
and U16265 (N_16265,N_13339,N_13336);
nor U16266 (N_16266,N_12717,N_12966);
or U16267 (N_16267,N_12679,N_12781);
and U16268 (N_16268,N_14671,N_12449);
nand U16269 (N_16269,N_14251,N_12202);
nor U16270 (N_16270,N_13513,N_12710);
nand U16271 (N_16271,N_13428,N_14299);
nor U16272 (N_16272,N_13660,N_12309);
or U16273 (N_16273,N_12240,N_14058);
and U16274 (N_16274,N_13621,N_12771);
nor U16275 (N_16275,N_13095,N_13669);
nor U16276 (N_16276,N_14153,N_12578);
nand U16277 (N_16277,N_12607,N_13082);
nor U16278 (N_16278,N_12196,N_14629);
or U16279 (N_16279,N_12062,N_14047);
xnor U16280 (N_16280,N_13642,N_12674);
nand U16281 (N_16281,N_13789,N_13747);
nand U16282 (N_16282,N_13626,N_13126);
nand U16283 (N_16283,N_14510,N_12408);
and U16284 (N_16284,N_12879,N_12297);
and U16285 (N_16285,N_13541,N_12254);
and U16286 (N_16286,N_14205,N_14243);
xnor U16287 (N_16287,N_13758,N_14673);
xor U16288 (N_16288,N_13073,N_12220);
nor U16289 (N_16289,N_14033,N_14456);
and U16290 (N_16290,N_14916,N_12346);
and U16291 (N_16291,N_12892,N_13408);
nand U16292 (N_16292,N_14418,N_13756);
and U16293 (N_16293,N_13977,N_13280);
and U16294 (N_16294,N_12376,N_14245);
or U16295 (N_16295,N_12011,N_12323);
xor U16296 (N_16296,N_13757,N_13311);
xor U16297 (N_16297,N_13323,N_13364);
nor U16298 (N_16298,N_12359,N_13224);
and U16299 (N_16299,N_13833,N_12734);
and U16300 (N_16300,N_14015,N_12671);
nor U16301 (N_16301,N_12448,N_14825);
nor U16302 (N_16302,N_14703,N_12092);
nand U16303 (N_16303,N_12527,N_13982);
and U16304 (N_16304,N_14162,N_12401);
nand U16305 (N_16305,N_14963,N_13327);
nor U16306 (N_16306,N_14631,N_14346);
nor U16307 (N_16307,N_14659,N_14025);
nor U16308 (N_16308,N_12040,N_12535);
nand U16309 (N_16309,N_12489,N_13664);
nand U16310 (N_16310,N_13129,N_13464);
or U16311 (N_16311,N_13484,N_13186);
xnor U16312 (N_16312,N_13064,N_13226);
nand U16313 (N_16313,N_13856,N_13158);
or U16314 (N_16314,N_12121,N_14805);
nor U16315 (N_16315,N_13857,N_12064);
nand U16316 (N_16316,N_13288,N_14747);
and U16317 (N_16317,N_13393,N_13657);
nor U16318 (N_16318,N_13955,N_13924);
or U16319 (N_16319,N_13663,N_13957);
nand U16320 (N_16320,N_14758,N_13203);
or U16321 (N_16321,N_12597,N_12216);
or U16322 (N_16322,N_13605,N_12676);
xnor U16323 (N_16323,N_14892,N_13488);
nor U16324 (N_16324,N_12409,N_13007);
nand U16325 (N_16325,N_13858,N_14998);
xnor U16326 (N_16326,N_14467,N_14915);
nand U16327 (N_16327,N_13360,N_14139);
nand U16328 (N_16328,N_14046,N_14929);
and U16329 (N_16329,N_12148,N_12279);
and U16330 (N_16330,N_14670,N_13414);
nor U16331 (N_16331,N_14922,N_13324);
nor U16332 (N_16332,N_12682,N_13468);
xnor U16333 (N_16333,N_14561,N_14907);
xor U16334 (N_16334,N_13096,N_13773);
and U16335 (N_16335,N_14383,N_14591);
and U16336 (N_16336,N_12846,N_12411);
nor U16337 (N_16337,N_13264,N_12979);
nor U16338 (N_16338,N_12794,N_14264);
xor U16339 (N_16339,N_14489,N_13651);
and U16340 (N_16340,N_13373,N_13477);
xnor U16341 (N_16341,N_14186,N_14282);
xor U16342 (N_16342,N_14957,N_12315);
or U16343 (N_16343,N_14201,N_13530);
nand U16344 (N_16344,N_14541,N_12151);
nor U16345 (N_16345,N_13070,N_14222);
xor U16346 (N_16346,N_12371,N_12190);
or U16347 (N_16347,N_14270,N_12580);
or U16348 (N_16348,N_14960,N_12500);
xnor U16349 (N_16349,N_12229,N_12154);
nor U16350 (N_16350,N_12329,N_12399);
nor U16351 (N_16351,N_12293,N_12526);
nand U16352 (N_16352,N_13200,N_12504);
xnor U16353 (N_16353,N_12572,N_12780);
or U16354 (N_16354,N_14316,N_13325);
and U16355 (N_16355,N_13736,N_14125);
or U16356 (N_16356,N_12194,N_13433);
nor U16357 (N_16357,N_13831,N_12469);
xor U16358 (N_16358,N_13462,N_12301);
nor U16359 (N_16359,N_12198,N_14783);
nor U16360 (N_16360,N_12735,N_12645);
or U16361 (N_16361,N_12341,N_12872);
or U16362 (N_16362,N_12548,N_14484);
nor U16363 (N_16363,N_14962,N_12231);
nor U16364 (N_16364,N_13562,N_14973);
xnor U16365 (N_16365,N_14964,N_14766);
xnor U16366 (N_16366,N_14736,N_13431);
xnor U16367 (N_16367,N_13234,N_14745);
xor U16368 (N_16368,N_13166,N_14191);
nor U16369 (N_16369,N_12792,N_13899);
xnor U16370 (N_16370,N_14578,N_12769);
or U16371 (N_16371,N_14248,N_12854);
xnor U16372 (N_16372,N_13439,N_12943);
or U16373 (N_16373,N_13668,N_13503);
nor U16374 (N_16374,N_14443,N_13243);
nor U16375 (N_16375,N_13334,N_13641);
nand U16376 (N_16376,N_14473,N_13115);
or U16377 (N_16377,N_14553,N_13608);
xor U16378 (N_16378,N_14110,N_13395);
and U16379 (N_16379,N_14906,N_12457);
or U16380 (N_16380,N_13015,N_14420);
or U16381 (N_16381,N_12106,N_14300);
nand U16382 (N_16382,N_14524,N_12884);
nand U16383 (N_16383,N_14345,N_12179);
and U16384 (N_16384,N_13846,N_13796);
and U16385 (N_16385,N_12876,N_12135);
xor U16386 (N_16386,N_14569,N_12081);
or U16387 (N_16387,N_12159,N_12586);
and U16388 (N_16388,N_13028,N_13949);
or U16389 (N_16389,N_14658,N_14751);
nor U16390 (N_16390,N_12243,N_12851);
or U16391 (N_16391,N_12014,N_13039);
nor U16392 (N_16392,N_14893,N_13830);
and U16393 (N_16393,N_14060,N_13132);
xor U16394 (N_16394,N_12721,N_14581);
nand U16395 (N_16395,N_13196,N_14895);
xnor U16396 (N_16396,N_13808,N_14912);
or U16397 (N_16397,N_12296,N_12474);
nor U16398 (N_16398,N_14800,N_13942);
and U16399 (N_16399,N_14855,N_13954);
or U16400 (N_16400,N_13965,N_14604);
nand U16401 (N_16401,N_13912,N_13784);
or U16402 (N_16402,N_12195,N_13918);
and U16403 (N_16403,N_14036,N_13060);
nor U16404 (N_16404,N_12827,N_14206);
xnor U16405 (N_16405,N_13798,N_13386);
nand U16406 (N_16406,N_13155,N_13315);
or U16407 (N_16407,N_14967,N_13685);
xor U16408 (N_16408,N_14989,N_13423);
or U16409 (N_16409,N_14900,N_13180);
xor U16410 (N_16410,N_13759,N_14062);
or U16411 (N_16411,N_14070,N_12729);
nor U16412 (N_16412,N_13206,N_14620);
xor U16413 (N_16413,N_13091,N_13739);
nor U16414 (N_16414,N_13848,N_13072);
nor U16415 (N_16415,N_12211,N_13337);
or U16416 (N_16416,N_13071,N_14452);
nor U16417 (N_16417,N_13999,N_12998);
nor U16418 (N_16418,N_13314,N_12620);
nand U16419 (N_16419,N_12260,N_14862);
nand U16420 (N_16420,N_12052,N_14575);
or U16421 (N_16421,N_13557,N_12626);
or U16422 (N_16422,N_13151,N_14884);
nand U16423 (N_16423,N_13744,N_13231);
nand U16424 (N_16424,N_12590,N_12569);
and U16425 (N_16425,N_14339,N_12974);
or U16426 (N_16426,N_12688,N_12950);
and U16427 (N_16427,N_13289,N_14358);
xor U16428 (N_16428,N_14132,N_14529);
or U16429 (N_16429,N_12886,N_14492);
or U16430 (N_16430,N_12053,N_14387);
nand U16431 (N_16431,N_12715,N_12112);
nor U16432 (N_16432,N_12733,N_13969);
nand U16433 (N_16433,N_12762,N_12031);
nor U16434 (N_16434,N_12029,N_14838);
nor U16435 (N_16435,N_14301,N_13214);
or U16436 (N_16436,N_12470,N_13761);
xnor U16437 (N_16437,N_13514,N_14382);
and U16438 (N_16438,N_13254,N_12991);
xor U16439 (N_16439,N_12137,N_14602);
or U16440 (N_16440,N_13994,N_12431);
or U16441 (N_16441,N_13953,N_14224);
or U16442 (N_16442,N_13976,N_12015);
and U16443 (N_16443,N_13864,N_14116);
nand U16444 (N_16444,N_14538,N_13549);
nand U16445 (N_16445,N_14189,N_12248);
and U16446 (N_16446,N_12414,N_12782);
or U16447 (N_16447,N_14355,N_13121);
or U16448 (N_16448,N_12403,N_12536);
nand U16449 (N_16449,N_13001,N_12706);
xnor U16450 (N_16450,N_13092,N_14774);
and U16451 (N_16451,N_12716,N_14202);
and U16452 (N_16452,N_14315,N_14609);
nor U16453 (N_16453,N_14041,N_14091);
and U16454 (N_16454,N_13475,N_14891);
nand U16455 (N_16455,N_14974,N_14988);
nand U16456 (N_16456,N_13124,N_14317);
and U16457 (N_16457,N_13636,N_13896);
or U16458 (N_16458,N_12388,N_12362);
nand U16459 (N_16459,N_14717,N_13571);
xor U16460 (N_16460,N_13084,N_13011);
xor U16461 (N_16461,N_12518,N_13618);
xor U16462 (N_16462,N_14801,N_13904);
or U16463 (N_16463,N_12384,N_12126);
nand U16464 (N_16464,N_12387,N_13159);
and U16465 (N_16465,N_13890,N_13086);
and U16466 (N_16466,N_13986,N_14982);
and U16467 (N_16467,N_14353,N_13482);
and U16468 (N_16468,N_13811,N_13961);
or U16469 (N_16469,N_13582,N_14426);
and U16470 (N_16470,N_14564,N_13109);
and U16471 (N_16471,N_14488,N_14714);
or U16472 (N_16472,N_12786,N_13420);
xnor U16473 (N_16473,N_13343,N_13841);
nor U16474 (N_16474,N_13443,N_13161);
or U16475 (N_16475,N_12321,N_12654);
nand U16476 (N_16476,N_13377,N_13545);
nor U16477 (N_16477,N_13281,N_13632);
or U16478 (N_16478,N_12962,N_13570);
nand U16479 (N_16479,N_12438,N_12681);
xnor U16480 (N_16480,N_13703,N_13305);
or U16481 (N_16481,N_14233,N_13220);
or U16482 (N_16482,N_14416,N_12405);
or U16483 (N_16483,N_12079,N_12440);
nor U16484 (N_16484,N_14371,N_13333);
and U16485 (N_16485,N_13970,N_12483);
and U16486 (N_16486,N_14267,N_12627);
nand U16487 (N_16487,N_13215,N_14715);
nand U16488 (N_16488,N_14821,N_14004);
and U16489 (N_16489,N_14367,N_13366);
or U16490 (N_16490,N_12983,N_14913);
and U16491 (N_16491,N_14807,N_14754);
xor U16492 (N_16492,N_14203,N_13463);
and U16493 (N_16493,N_12467,N_12520);
nor U16494 (N_16494,N_13277,N_13643);
or U16495 (N_16495,N_12334,N_13877);
xnor U16496 (N_16496,N_14500,N_13112);
or U16497 (N_16497,N_13228,N_13233);
xnor U16498 (N_16498,N_13837,N_14858);
or U16499 (N_16499,N_14874,N_12850);
xnor U16500 (N_16500,N_12890,N_13510);
nand U16501 (N_16501,N_14093,N_12250);
and U16502 (N_16502,N_13684,N_12050);
or U16503 (N_16503,N_14519,N_14784);
nand U16504 (N_16504,N_14551,N_12398);
nor U16505 (N_16505,N_13920,N_12617);
or U16506 (N_16506,N_12413,N_12349);
nor U16507 (N_16507,N_13117,N_14558);
and U16508 (N_16508,N_13431,N_13587);
nor U16509 (N_16509,N_13590,N_13161);
and U16510 (N_16510,N_12890,N_13402);
and U16511 (N_16511,N_12416,N_14756);
xor U16512 (N_16512,N_12574,N_12554);
and U16513 (N_16513,N_12965,N_13339);
nand U16514 (N_16514,N_14254,N_13368);
and U16515 (N_16515,N_13471,N_13663);
xor U16516 (N_16516,N_12786,N_14867);
xor U16517 (N_16517,N_14410,N_12633);
xnor U16518 (N_16518,N_12471,N_14374);
xnor U16519 (N_16519,N_12518,N_13242);
nor U16520 (N_16520,N_14167,N_14577);
nor U16521 (N_16521,N_14905,N_12142);
and U16522 (N_16522,N_13787,N_14929);
or U16523 (N_16523,N_13463,N_12192);
or U16524 (N_16524,N_13803,N_14973);
and U16525 (N_16525,N_12623,N_12246);
xor U16526 (N_16526,N_12167,N_13109);
and U16527 (N_16527,N_14631,N_14697);
nor U16528 (N_16528,N_13638,N_12453);
nor U16529 (N_16529,N_12838,N_14668);
nor U16530 (N_16530,N_14318,N_13847);
nand U16531 (N_16531,N_14153,N_13500);
and U16532 (N_16532,N_13949,N_14574);
nand U16533 (N_16533,N_14936,N_12498);
or U16534 (N_16534,N_12288,N_13687);
or U16535 (N_16535,N_12317,N_14507);
and U16536 (N_16536,N_12733,N_14838);
or U16537 (N_16537,N_14119,N_14697);
xor U16538 (N_16538,N_12860,N_14784);
and U16539 (N_16539,N_13837,N_12997);
and U16540 (N_16540,N_13489,N_13707);
and U16541 (N_16541,N_12357,N_12080);
and U16542 (N_16542,N_12625,N_13660);
and U16543 (N_16543,N_12990,N_12384);
nand U16544 (N_16544,N_13474,N_12313);
or U16545 (N_16545,N_13757,N_13859);
and U16546 (N_16546,N_13148,N_12409);
nand U16547 (N_16547,N_13811,N_14517);
and U16548 (N_16548,N_14709,N_13286);
and U16549 (N_16549,N_12356,N_14861);
and U16550 (N_16550,N_14633,N_12669);
or U16551 (N_16551,N_12733,N_14961);
nor U16552 (N_16552,N_12735,N_13878);
nor U16553 (N_16553,N_13327,N_12482);
xor U16554 (N_16554,N_14555,N_14991);
nor U16555 (N_16555,N_12146,N_12528);
xnor U16556 (N_16556,N_14908,N_14285);
xnor U16557 (N_16557,N_13201,N_13809);
nand U16558 (N_16558,N_12999,N_12228);
nand U16559 (N_16559,N_12847,N_12655);
xor U16560 (N_16560,N_13843,N_12554);
xor U16561 (N_16561,N_13070,N_12213);
nand U16562 (N_16562,N_12295,N_12875);
nand U16563 (N_16563,N_13216,N_13841);
nor U16564 (N_16564,N_14450,N_12197);
or U16565 (N_16565,N_12187,N_13387);
xor U16566 (N_16566,N_13338,N_14942);
or U16567 (N_16567,N_13110,N_14907);
nor U16568 (N_16568,N_12482,N_14085);
nor U16569 (N_16569,N_14592,N_14023);
nor U16570 (N_16570,N_13329,N_12875);
nand U16571 (N_16571,N_12577,N_12802);
or U16572 (N_16572,N_14429,N_12810);
or U16573 (N_16573,N_13454,N_13194);
xor U16574 (N_16574,N_12197,N_14613);
xor U16575 (N_16575,N_14048,N_13171);
and U16576 (N_16576,N_12221,N_14606);
nor U16577 (N_16577,N_12426,N_12638);
xnor U16578 (N_16578,N_13772,N_12437);
nand U16579 (N_16579,N_13572,N_14300);
xor U16580 (N_16580,N_12457,N_12141);
and U16581 (N_16581,N_13718,N_12467);
nor U16582 (N_16582,N_12673,N_12181);
and U16583 (N_16583,N_14063,N_12191);
nor U16584 (N_16584,N_14135,N_12580);
nor U16585 (N_16585,N_14794,N_12503);
and U16586 (N_16586,N_12461,N_13277);
nor U16587 (N_16587,N_13890,N_13678);
nand U16588 (N_16588,N_12259,N_12463);
nor U16589 (N_16589,N_12666,N_14877);
and U16590 (N_16590,N_12149,N_13210);
and U16591 (N_16591,N_14290,N_12299);
or U16592 (N_16592,N_13087,N_12530);
nor U16593 (N_16593,N_12703,N_14426);
and U16594 (N_16594,N_14511,N_13063);
or U16595 (N_16595,N_13622,N_12070);
and U16596 (N_16596,N_13196,N_14071);
nor U16597 (N_16597,N_12657,N_12253);
nor U16598 (N_16598,N_12546,N_12794);
xor U16599 (N_16599,N_14647,N_13153);
nor U16600 (N_16600,N_14356,N_12200);
or U16601 (N_16601,N_14609,N_14715);
nand U16602 (N_16602,N_14028,N_13973);
nand U16603 (N_16603,N_14750,N_13479);
or U16604 (N_16604,N_12015,N_14788);
xor U16605 (N_16605,N_14734,N_13072);
xnor U16606 (N_16606,N_13460,N_12667);
nand U16607 (N_16607,N_12336,N_13380);
or U16608 (N_16608,N_12708,N_13563);
nand U16609 (N_16609,N_12734,N_14131);
nand U16610 (N_16610,N_13791,N_14419);
nand U16611 (N_16611,N_14664,N_13826);
xor U16612 (N_16612,N_12639,N_12328);
and U16613 (N_16613,N_13207,N_13961);
and U16614 (N_16614,N_13399,N_12030);
nor U16615 (N_16615,N_14500,N_12740);
xnor U16616 (N_16616,N_14182,N_13901);
nor U16617 (N_16617,N_13705,N_14440);
or U16618 (N_16618,N_14105,N_12667);
and U16619 (N_16619,N_14215,N_14674);
xor U16620 (N_16620,N_12596,N_13812);
xnor U16621 (N_16621,N_14582,N_12094);
or U16622 (N_16622,N_13756,N_13982);
or U16623 (N_16623,N_13122,N_13852);
nand U16624 (N_16624,N_14986,N_14224);
or U16625 (N_16625,N_12148,N_12997);
and U16626 (N_16626,N_12265,N_14233);
xnor U16627 (N_16627,N_13767,N_14960);
and U16628 (N_16628,N_14367,N_14133);
or U16629 (N_16629,N_14829,N_12692);
nand U16630 (N_16630,N_12016,N_12752);
or U16631 (N_16631,N_13743,N_13878);
nand U16632 (N_16632,N_14980,N_13418);
nand U16633 (N_16633,N_14407,N_13452);
nand U16634 (N_16634,N_12802,N_12220);
nor U16635 (N_16635,N_14411,N_14258);
or U16636 (N_16636,N_12154,N_14924);
nor U16637 (N_16637,N_14185,N_14721);
nand U16638 (N_16638,N_14837,N_13462);
or U16639 (N_16639,N_13103,N_12784);
nand U16640 (N_16640,N_12238,N_14596);
or U16641 (N_16641,N_12252,N_14482);
nor U16642 (N_16642,N_12725,N_13704);
xor U16643 (N_16643,N_14230,N_13846);
nand U16644 (N_16644,N_12235,N_13575);
or U16645 (N_16645,N_12339,N_14021);
nor U16646 (N_16646,N_14002,N_14772);
or U16647 (N_16647,N_12098,N_12334);
and U16648 (N_16648,N_14817,N_14100);
xor U16649 (N_16649,N_14422,N_13126);
xor U16650 (N_16650,N_12131,N_12002);
nor U16651 (N_16651,N_12480,N_12223);
nand U16652 (N_16652,N_13912,N_14694);
xnor U16653 (N_16653,N_13833,N_14907);
nor U16654 (N_16654,N_12114,N_13853);
xnor U16655 (N_16655,N_14295,N_14161);
and U16656 (N_16656,N_13665,N_14736);
and U16657 (N_16657,N_14517,N_14144);
or U16658 (N_16658,N_12415,N_12216);
or U16659 (N_16659,N_12398,N_14160);
and U16660 (N_16660,N_13778,N_12948);
nor U16661 (N_16661,N_13280,N_14355);
or U16662 (N_16662,N_13565,N_12148);
xnor U16663 (N_16663,N_12647,N_13669);
and U16664 (N_16664,N_14419,N_12146);
xor U16665 (N_16665,N_13886,N_13689);
nand U16666 (N_16666,N_14672,N_13246);
nand U16667 (N_16667,N_12081,N_14266);
xnor U16668 (N_16668,N_14917,N_13934);
nand U16669 (N_16669,N_13746,N_14571);
nand U16670 (N_16670,N_12014,N_13622);
and U16671 (N_16671,N_12340,N_12660);
nor U16672 (N_16672,N_13381,N_14343);
nor U16673 (N_16673,N_13390,N_12835);
or U16674 (N_16674,N_14037,N_12637);
or U16675 (N_16675,N_13140,N_12880);
xnor U16676 (N_16676,N_14033,N_14633);
and U16677 (N_16677,N_14294,N_12379);
xnor U16678 (N_16678,N_12181,N_13820);
and U16679 (N_16679,N_13048,N_14455);
or U16680 (N_16680,N_12855,N_13018);
and U16681 (N_16681,N_13989,N_14871);
nand U16682 (N_16682,N_14622,N_13424);
and U16683 (N_16683,N_13057,N_14621);
and U16684 (N_16684,N_12597,N_14756);
and U16685 (N_16685,N_14361,N_13208);
xor U16686 (N_16686,N_13285,N_12632);
xnor U16687 (N_16687,N_12784,N_12008);
nand U16688 (N_16688,N_14341,N_13428);
nor U16689 (N_16689,N_12832,N_14418);
or U16690 (N_16690,N_12600,N_14059);
nor U16691 (N_16691,N_14005,N_12449);
or U16692 (N_16692,N_12456,N_13247);
xor U16693 (N_16693,N_14626,N_14516);
xnor U16694 (N_16694,N_12166,N_13995);
nor U16695 (N_16695,N_12292,N_14498);
or U16696 (N_16696,N_13218,N_14224);
xnor U16697 (N_16697,N_13479,N_14780);
xor U16698 (N_16698,N_13999,N_14949);
and U16699 (N_16699,N_14628,N_14305);
xor U16700 (N_16700,N_13824,N_13514);
nor U16701 (N_16701,N_14377,N_13472);
nand U16702 (N_16702,N_12875,N_12692);
xor U16703 (N_16703,N_13244,N_13528);
xor U16704 (N_16704,N_13701,N_12297);
and U16705 (N_16705,N_12090,N_13564);
xnor U16706 (N_16706,N_14718,N_13815);
xor U16707 (N_16707,N_12738,N_14563);
xor U16708 (N_16708,N_14444,N_14456);
nand U16709 (N_16709,N_13585,N_13091);
nor U16710 (N_16710,N_12368,N_12920);
xor U16711 (N_16711,N_14101,N_14477);
and U16712 (N_16712,N_13875,N_12794);
or U16713 (N_16713,N_12827,N_14506);
nor U16714 (N_16714,N_13195,N_13437);
xor U16715 (N_16715,N_12985,N_14864);
nor U16716 (N_16716,N_13073,N_13181);
and U16717 (N_16717,N_13965,N_12736);
nor U16718 (N_16718,N_14830,N_14155);
nor U16719 (N_16719,N_12682,N_12032);
or U16720 (N_16720,N_14811,N_14242);
and U16721 (N_16721,N_13056,N_13185);
nand U16722 (N_16722,N_13639,N_13608);
and U16723 (N_16723,N_14387,N_12634);
nor U16724 (N_16724,N_13684,N_14733);
nand U16725 (N_16725,N_14476,N_12987);
and U16726 (N_16726,N_13223,N_12306);
nand U16727 (N_16727,N_14742,N_12539);
xor U16728 (N_16728,N_12317,N_12515);
or U16729 (N_16729,N_14274,N_13706);
or U16730 (N_16730,N_12561,N_14816);
xor U16731 (N_16731,N_13152,N_12235);
nand U16732 (N_16732,N_12399,N_12520);
nand U16733 (N_16733,N_13391,N_13679);
nand U16734 (N_16734,N_12720,N_12668);
and U16735 (N_16735,N_13967,N_12046);
nand U16736 (N_16736,N_13673,N_12569);
nor U16737 (N_16737,N_14748,N_12900);
or U16738 (N_16738,N_12351,N_14294);
nand U16739 (N_16739,N_13304,N_12584);
nor U16740 (N_16740,N_12008,N_13821);
nand U16741 (N_16741,N_12191,N_12536);
xor U16742 (N_16742,N_12086,N_14989);
nor U16743 (N_16743,N_14579,N_13665);
xor U16744 (N_16744,N_12537,N_13596);
or U16745 (N_16745,N_13003,N_13582);
or U16746 (N_16746,N_13023,N_12744);
xor U16747 (N_16747,N_14809,N_12761);
xnor U16748 (N_16748,N_12518,N_14678);
nand U16749 (N_16749,N_13422,N_12642);
nor U16750 (N_16750,N_12821,N_13449);
xor U16751 (N_16751,N_12329,N_14030);
and U16752 (N_16752,N_12663,N_14761);
xor U16753 (N_16753,N_12981,N_13669);
nor U16754 (N_16754,N_14455,N_14763);
and U16755 (N_16755,N_13783,N_14843);
or U16756 (N_16756,N_13221,N_12163);
and U16757 (N_16757,N_13934,N_14241);
nand U16758 (N_16758,N_12477,N_13494);
and U16759 (N_16759,N_14126,N_12034);
and U16760 (N_16760,N_14969,N_12662);
and U16761 (N_16761,N_13543,N_13694);
and U16762 (N_16762,N_14223,N_14097);
xnor U16763 (N_16763,N_14135,N_13823);
nor U16764 (N_16764,N_13620,N_14516);
and U16765 (N_16765,N_14892,N_13584);
or U16766 (N_16766,N_12586,N_13567);
and U16767 (N_16767,N_12023,N_13934);
or U16768 (N_16768,N_12265,N_14801);
and U16769 (N_16769,N_13302,N_14847);
nand U16770 (N_16770,N_12520,N_14954);
or U16771 (N_16771,N_14015,N_14707);
and U16772 (N_16772,N_14426,N_14535);
nor U16773 (N_16773,N_13540,N_14300);
nand U16774 (N_16774,N_12357,N_14567);
or U16775 (N_16775,N_14558,N_13378);
and U16776 (N_16776,N_12920,N_14856);
and U16777 (N_16777,N_13793,N_12346);
or U16778 (N_16778,N_14012,N_13072);
nand U16779 (N_16779,N_14597,N_14170);
nor U16780 (N_16780,N_14699,N_14318);
nor U16781 (N_16781,N_14372,N_13293);
or U16782 (N_16782,N_12524,N_13116);
and U16783 (N_16783,N_12666,N_14992);
and U16784 (N_16784,N_12731,N_14445);
xor U16785 (N_16785,N_12343,N_14909);
nand U16786 (N_16786,N_12096,N_14282);
or U16787 (N_16787,N_12565,N_14213);
xnor U16788 (N_16788,N_13383,N_13656);
xor U16789 (N_16789,N_12884,N_13660);
nand U16790 (N_16790,N_13786,N_14428);
xor U16791 (N_16791,N_12960,N_14481);
nor U16792 (N_16792,N_12056,N_14149);
and U16793 (N_16793,N_13410,N_13296);
and U16794 (N_16794,N_12729,N_12779);
nand U16795 (N_16795,N_13715,N_14429);
nor U16796 (N_16796,N_14014,N_14473);
nor U16797 (N_16797,N_14537,N_13796);
xnor U16798 (N_16798,N_14032,N_14551);
and U16799 (N_16799,N_13612,N_12286);
nand U16800 (N_16800,N_12658,N_13050);
nor U16801 (N_16801,N_14146,N_13908);
or U16802 (N_16802,N_13724,N_12053);
xor U16803 (N_16803,N_12815,N_12666);
nor U16804 (N_16804,N_12943,N_13485);
nand U16805 (N_16805,N_13265,N_14050);
or U16806 (N_16806,N_14722,N_13782);
nor U16807 (N_16807,N_12109,N_12954);
or U16808 (N_16808,N_14207,N_12484);
nor U16809 (N_16809,N_12617,N_12735);
xnor U16810 (N_16810,N_12490,N_13317);
nor U16811 (N_16811,N_12575,N_12754);
and U16812 (N_16812,N_13153,N_12248);
nor U16813 (N_16813,N_12115,N_12142);
or U16814 (N_16814,N_14929,N_14048);
or U16815 (N_16815,N_13317,N_13604);
xor U16816 (N_16816,N_14171,N_14861);
and U16817 (N_16817,N_13187,N_14971);
xnor U16818 (N_16818,N_13168,N_12870);
and U16819 (N_16819,N_14310,N_13783);
nand U16820 (N_16820,N_13369,N_12360);
nor U16821 (N_16821,N_12795,N_12415);
xor U16822 (N_16822,N_14521,N_14054);
nand U16823 (N_16823,N_13048,N_14795);
xnor U16824 (N_16824,N_12829,N_14164);
or U16825 (N_16825,N_12664,N_14927);
and U16826 (N_16826,N_13705,N_14069);
nand U16827 (N_16827,N_12864,N_14890);
or U16828 (N_16828,N_12674,N_14032);
and U16829 (N_16829,N_14241,N_13861);
or U16830 (N_16830,N_12873,N_12319);
xor U16831 (N_16831,N_12731,N_14032);
xor U16832 (N_16832,N_12576,N_12865);
nand U16833 (N_16833,N_13019,N_14688);
and U16834 (N_16834,N_12329,N_12070);
nor U16835 (N_16835,N_13526,N_13270);
or U16836 (N_16836,N_12320,N_14119);
and U16837 (N_16837,N_12561,N_14209);
nand U16838 (N_16838,N_14569,N_13554);
or U16839 (N_16839,N_14830,N_13520);
nor U16840 (N_16840,N_12433,N_12705);
and U16841 (N_16841,N_12202,N_14083);
nor U16842 (N_16842,N_12801,N_14285);
and U16843 (N_16843,N_14124,N_13508);
nand U16844 (N_16844,N_14857,N_13618);
and U16845 (N_16845,N_14868,N_14246);
xnor U16846 (N_16846,N_14871,N_12334);
and U16847 (N_16847,N_13724,N_14067);
nand U16848 (N_16848,N_14794,N_12179);
or U16849 (N_16849,N_12336,N_12703);
or U16850 (N_16850,N_13272,N_12602);
and U16851 (N_16851,N_12913,N_14890);
nand U16852 (N_16852,N_13428,N_13414);
nor U16853 (N_16853,N_13869,N_12069);
nor U16854 (N_16854,N_14778,N_13439);
nor U16855 (N_16855,N_13486,N_12833);
nand U16856 (N_16856,N_12006,N_12919);
nand U16857 (N_16857,N_14289,N_13831);
nand U16858 (N_16858,N_14673,N_12320);
nand U16859 (N_16859,N_13719,N_14437);
xnor U16860 (N_16860,N_12658,N_12303);
nor U16861 (N_16861,N_13836,N_12835);
and U16862 (N_16862,N_14853,N_12301);
nand U16863 (N_16863,N_13811,N_14509);
nand U16864 (N_16864,N_12105,N_14418);
nand U16865 (N_16865,N_12840,N_12196);
xnor U16866 (N_16866,N_13010,N_14395);
and U16867 (N_16867,N_13117,N_13389);
nand U16868 (N_16868,N_13838,N_13908);
nor U16869 (N_16869,N_12052,N_14421);
nand U16870 (N_16870,N_14539,N_14905);
nand U16871 (N_16871,N_13076,N_13570);
nand U16872 (N_16872,N_13459,N_14754);
nand U16873 (N_16873,N_12625,N_14271);
and U16874 (N_16874,N_14875,N_12251);
nand U16875 (N_16875,N_14104,N_13361);
xor U16876 (N_16876,N_13765,N_13486);
and U16877 (N_16877,N_14327,N_13108);
nor U16878 (N_16878,N_13704,N_14120);
or U16879 (N_16879,N_12484,N_12706);
xor U16880 (N_16880,N_13262,N_13354);
and U16881 (N_16881,N_13455,N_12526);
and U16882 (N_16882,N_14983,N_14899);
or U16883 (N_16883,N_14164,N_14046);
xnor U16884 (N_16884,N_12456,N_12760);
and U16885 (N_16885,N_13188,N_14086);
and U16886 (N_16886,N_13283,N_14417);
and U16887 (N_16887,N_12560,N_13941);
nand U16888 (N_16888,N_14870,N_13371);
and U16889 (N_16889,N_14969,N_14376);
or U16890 (N_16890,N_12288,N_14693);
or U16891 (N_16891,N_13700,N_12079);
and U16892 (N_16892,N_12136,N_13211);
xor U16893 (N_16893,N_14807,N_12991);
or U16894 (N_16894,N_13559,N_12091);
or U16895 (N_16895,N_12181,N_13339);
nand U16896 (N_16896,N_14628,N_13000);
nor U16897 (N_16897,N_12684,N_14055);
nand U16898 (N_16898,N_12235,N_13490);
or U16899 (N_16899,N_12382,N_12169);
or U16900 (N_16900,N_13537,N_12286);
xnor U16901 (N_16901,N_12068,N_12141);
nor U16902 (N_16902,N_13089,N_12138);
nand U16903 (N_16903,N_14311,N_12010);
or U16904 (N_16904,N_12841,N_13708);
nand U16905 (N_16905,N_14239,N_13624);
nand U16906 (N_16906,N_13404,N_12798);
nand U16907 (N_16907,N_13109,N_12299);
or U16908 (N_16908,N_14375,N_14470);
xor U16909 (N_16909,N_14725,N_13012);
nand U16910 (N_16910,N_13605,N_13270);
nand U16911 (N_16911,N_13000,N_13291);
and U16912 (N_16912,N_14381,N_12465);
xor U16913 (N_16913,N_13549,N_13338);
nor U16914 (N_16914,N_14502,N_12425);
nor U16915 (N_16915,N_14480,N_13986);
and U16916 (N_16916,N_13268,N_12486);
nor U16917 (N_16917,N_12245,N_14790);
nand U16918 (N_16918,N_14895,N_12794);
or U16919 (N_16919,N_13923,N_14953);
nand U16920 (N_16920,N_13320,N_12155);
nor U16921 (N_16921,N_12321,N_13427);
and U16922 (N_16922,N_13485,N_12605);
xnor U16923 (N_16923,N_12615,N_14243);
xnor U16924 (N_16924,N_12776,N_13496);
nand U16925 (N_16925,N_13619,N_13539);
and U16926 (N_16926,N_14975,N_14723);
nor U16927 (N_16927,N_13758,N_12617);
or U16928 (N_16928,N_14930,N_12499);
nor U16929 (N_16929,N_14295,N_14381);
and U16930 (N_16930,N_14570,N_12365);
xor U16931 (N_16931,N_12898,N_12939);
nor U16932 (N_16932,N_12045,N_14365);
or U16933 (N_16933,N_13588,N_13764);
nor U16934 (N_16934,N_14547,N_14471);
or U16935 (N_16935,N_13166,N_12346);
nor U16936 (N_16936,N_13432,N_14975);
xor U16937 (N_16937,N_13587,N_14907);
or U16938 (N_16938,N_13894,N_12759);
or U16939 (N_16939,N_13638,N_12521);
and U16940 (N_16940,N_12139,N_12222);
xnor U16941 (N_16941,N_14018,N_14917);
and U16942 (N_16942,N_14491,N_14589);
nand U16943 (N_16943,N_12410,N_12750);
and U16944 (N_16944,N_14288,N_14829);
nor U16945 (N_16945,N_12811,N_14385);
and U16946 (N_16946,N_13379,N_13880);
nand U16947 (N_16947,N_13833,N_12222);
or U16948 (N_16948,N_12927,N_13032);
xor U16949 (N_16949,N_14940,N_14274);
xnor U16950 (N_16950,N_12437,N_12741);
xnor U16951 (N_16951,N_14318,N_12412);
nand U16952 (N_16952,N_13794,N_13703);
nor U16953 (N_16953,N_12122,N_14755);
xor U16954 (N_16954,N_13926,N_12875);
nand U16955 (N_16955,N_14584,N_13956);
and U16956 (N_16956,N_12545,N_13270);
or U16957 (N_16957,N_12184,N_13332);
nand U16958 (N_16958,N_13583,N_14608);
nand U16959 (N_16959,N_14838,N_12343);
nand U16960 (N_16960,N_14215,N_13252);
and U16961 (N_16961,N_14049,N_13334);
and U16962 (N_16962,N_12937,N_13121);
xor U16963 (N_16963,N_14268,N_13920);
nor U16964 (N_16964,N_12993,N_12055);
xor U16965 (N_16965,N_14864,N_14760);
and U16966 (N_16966,N_14529,N_12862);
or U16967 (N_16967,N_12176,N_13923);
nor U16968 (N_16968,N_12088,N_12502);
nor U16969 (N_16969,N_14093,N_14813);
and U16970 (N_16970,N_12280,N_12512);
or U16971 (N_16971,N_14585,N_12574);
and U16972 (N_16972,N_12359,N_14197);
nor U16973 (N_16973,N_13178,N_13957);
xor U16974 (N_16974,N_12393,N_14660);
nor U16975 (N_16975,N_14146,N_14935);
nor U16976 (N_16976,N_14790,N_12800);
and U16977 (N_16977,N_12145,N_13754);
nand U16978 (N_16978,N_12270,N_12090);
nand U16979 (N_16979,N_12200,N_13967);
nor U16980 (N_16980,N_13717,N_12682);
xnor U16981 (N_16981,N_13314,N_14284);
nor U16982 (N_16982,N_12735,N_14538);
nor U16983 (N_16983,N_14513,N_14687);
nor U16984 (N_16984,N_14115,N_12083);
or U16985 (N_16985,N_13528,N_13795);
or U16986 (N_16986,N_12385,N_13559);
nand U16987 (N_16987,N_14379,N_12872);
nor U16988 (N_16988,N_13200,N_14934);
and U16989 (N_16989,N_14010,N_13065);
nor U16990 (N_16990,N_13614,N_13556);
nand U16991 (N_16991,N_12402,N_14593);
nand U16992 (N_16992,N_12037,N_13433);
xnor U16993 (N_16993,N_14633,N_13767);
xor U16994 (N_16994,N_13006,N_13261);
xor U16995 (N_16995,N_12955,N_12827);
nor U16996 (N_16996,N_13621,N_14549);
xnor U16997 (N_16997,N_14295,N_13955);
nor U16998 (N_16998,N_13257,N_13772);
or U16999 (N_16999,N_13899,N_14611);
nor U17000 (N_17000,N_14584,N_13095);
nand U17001 (N_17001,N_13104,N_13479);
and U17002 (N_17002,N_12440,N_14262);
nor U17003 (N_17003,N_14468,N_14922);
nand U17004 (N_17004,N_14674,N_14850);
xor U17005 (N_17005,N_13141,N_14649);
nand U17006 (N_17006,N_14559,N_14140);
and U17007 (N_17007,N_12107,N_14622);
or U17008 (N_17008,N_12768,N_14133);
nand U17009 (N_17009,N_12413,N_14136);
nor U17010 (N_17010,N_14578,N_13448);
nor U17011 (N_17011,N_13933,N_12270);
xnor U17012 (N_17012,N_12418,N_14337);
or U17013 (N_17013,N_12593,N_12940);
or U17014 (N_17014,N_13726,N_13187);
or U17015 (N_17015,N_12000,N_14316);
xor U17016 (N_17016,N_12981,N_14763);
nor U17017 (N_17017,N_13820,N_14793);
or U17018 (N_17018,N_13905,N_13020);
nand U17019 (N_17019,N_13229,N_13685);
and U17020 (N_17020,N_13964,N_12617);
nand U17021 (N_17021,N_12827,N_14726);
nor U17022 (N_17022,N_12697,N_12594);
or U17023 (N_17023,N_13605,N_13565);
and U17024 (N_17024,N_14558,N_13434);
and U17025 (N_17025,N_13749,N_14857);
nand U17026 (N_17026,N_12683,N_12354);
nand U17027 (N_17027,N_13494,N_13708);
xnor U17028 (N_17028,N_13749,N_14062);
or U17029 (N_17029,N_12281,N_12381);
nand U17030 (N_17030,N_14696,N_13832);
nand U17031 (N_17031,N_12172,N_12178);
xnor U17032 (N_17032,N_14499,N_14047);
xor U17033 (N_17033,N_14451,N_14979);
and U17034 (N_17034,N_14692,N_13943);
nor U17035 (N_17035,N_12907,N_13839);
or U17036 (N_17036,N_12566,N_14798);
or U17037 (N_17037,N_14204,N_13618);
or U17038 (N_17038,N_14397,N_12607);
xor U17039 (N_17039,N_12591,N_12418);
nand U17040 (N_17040,N_14899,N_12630);
and U17041 (N_17041,N_12885,N_14198);
xnor U17042 (N_17042,N_13701,N_13654);
nand U17043 (N_17043,N_13152,N_12639);
and U17044 (N_17044,N_14529,N_12719);
and U17045 (N_17045,N_12330,N_12126);
nand U17046 (N_17046,N_14812,N_12661);
nand U17047 (N_17047,N_14512,N_12892);
nor U17048 (N_17048,N_13974,N_14633);
and U17049 (N_17049,N_13784,N_13119);
and U17050 (N_17050,N_13654,N_12659);
xnor U17051 (N_17051,N_12810,N_13895);
nand U17052 (N_17052,N_14765,N_12914);
nand U17053 (N_17053,N_12526,N_13244);
xor U17054 (N_17054,N_13709,N_13774);
or U17055 (N_17055,N_13814,N_14514);
and U17056 (N_17056,N_13461,N_13924);
and U17057 (N_17057,N_13557,N_13192);
nand U17058 (N_17058,N_14041,N_12542);
or U17059 (N_17059,N_14483,N_12039);
nor U17060 (N_17060,N_12075,N_14696);
and U17061 (N_17061,N_14099,N_12073);
nor U17062 (N_17062,N_12858,N_13948);
xor U17063 (N_17063,N_14254,N_14450);
nor U17064 (N_17064,N_14633,N_14423);
nand U17065 (N_17065,N_13926,N_12301);
or U17066 (N_17066,N_13362,N_12327);
or U17067 (N_17067,N_14633,N_13264);
nand U17068 (N_17068,N_13912,N_14784);
nor U17069 (N_17069,N_12662,N_13345);
nand U17070 (N_17070,N_13963,N_14629);
and U17071 (N_17071,N_14808,N_14310);
and U17072 (N_17072,N_12551,N_12206);
nand U17073 (N_17073,N_13851,N_14941);
nor U17074 (N_17074,N_14737,N_13533);
xnor U17075 (N_17075,N_13889,N_13651);
and U17076 (N_17076,N_14757,N_14467);
xnor U17077 (N_17077,N_14938,N_13692);
xor U17078 (N_17078,N_13642,N_12960);
and U17079 (N_17079,N_12544,N_13272);
nand U17080 (N_17080,N_13043,N_13873);
xnor U17081 (N_17081,N_12373,N_12427);
and U17082 (N_17082,N_13525,N_12695);
xnor U17083 (N_17083,N_14422,N_14369);
nor U17084 (N_17084,N_12700,N_13083);
or U17085 (N_17085,N_13671,N_12471);
and U17086 (N_17086,N_13713,N_12251);
or U17087 (N_17087,N_12974,N_13442);
nor U17088 (N_17088,N_13368,N_13474);
and U17089 (N_17089,N_13954,N_13353);
and U17090 (N_17090,N_12458,N_14470);
xor U17091 (N_17091,N_14195,N_12484);
nand U17092 (N_17092,N_14405,N_13340);
and U17093 (N_17093,N_12431,N_13702);
or U17094 (N_17094,N_12789,N_12905);
or U17095 (N_17095,N_13603,N_14222);
or U17096 (N_17096,N_14706,N_14139);
nor U17097 (N_17097,N_14583,N_14471);
xnor U17098 (N_17098,N_14677,N_13773);
nand U17099 (N_17099,N_12942,N_12196);
nand U17100 (N_17100,N_12740,N_13872);
nand U17101 (N_17101,N_13633,N_14132);
and U17102 (N_17102,N_12351,N_12091);
or U17103 (N_17103,N_12779,N_12653);
or U17104 (N_17104,N_12572,N_12182);
nand U17105 (N_17105,N_12754,N_14274);
nor U17106 (N_17106,N_14968,N_13101);
nor U17107 (N_17107,N_14966,N_13904);
nand U17108 (N_17108,N_13460,N_12512);
xor U17109 (N_17109,N_14426,N_13831);
and U17110 (N_17110,N_12073,N_13646);
xnor U17111 (N_17111,N_13496,N_13062);
xor U17112 (N_17112,N_12263,N_12193);
xnor U17113 (N_17113,N_12753,N_12411);
and U17114 (N_17114,N_13236,N_14937);
xnor U17115 (N_17115,N_13446,N_12118);
and U17116 (N_17116,N_14344,N_12282);
nand U17117 (N_17117,N_14971,N_12184);
xnor U17118 (N_17118,N_14362,N_12739);
nor U17119 (N_17119,N_13352,N_13454);
xnor U17120 (N_17120,N_14897,N_13448);
xor U17121 (N_17121,N_14494,N_13748);
xnor U17122 (N_17122,N_12387,N_13243);
xor U17123 (N_17123,N_14963,N_14298);
xor U17124 (N_17124,N_14969,N_13894);
and U17125 (N_17125,N_13485,N_13861);
nand U17126 (N_17126,N_14777,N_12603);
xnor U17127 (N_17127,N_12066,N_14944);
nor U17128 (N_17128,N_14259,N_12842);
nor U17129 (N_17129,N_14266,N_12190);
xnor U17130 (N_17130,N_13156,N_14344);
nand U17131 (N_17131,N_12389,N_13905);
nand U17132 (N_17132,N_13420,N_13820);
and U17133 (N_17133,N_12918,N_14286);
and U17134 (N_17134,N_14278,N_12868);
nor U17135 (N_17135,N_13426,N_14527);
xnor U17136 (N_17136,N_13340,N_13962);
and U17137 (N_17137,N_12666,N_12818);
or U17138 (N_17138,N_12347,N_14397);
and U17139 (N_17139,N_14881,N_14597);
and U17140 (N_17140,N_12554,N_12299);
or U17141 (N_17141,N_12221,N_12104);
and U17142 (N_17142,N_14321,N_12324);
xnor U17143 (N_17143,N_12033,N_13223);
xnor U17144 (N_17144,N_12783,N_12714);
xnor U17145 (N_17145,N_14923,N_12081);
xnor U17146 (N_17146,N_13584,N_12745);
and U17147 (N_17147,N_12568,N_12553);
xnor U17148 (N_17148,N_12276,N_14148);
and U17149 (N_17149,N_13334,N_14411);
nor U17150 (N_17150,N_12786,N_14313);
nand U17151 (N_17151,N_14327,N_13050);
and U17152 (N_17152,N_12690,N_13007);
nor U17153 (N_17153,N_14925,N_14519);
and U17154 (N_17154,N_14816,N_12572);
or U17155 (N_17155,N_13828,N_13942);
xnor U17156 (N_17156,N_12633,N_12361);
nor U17157 (N_17157,N_14887,N_13822);
nor U17158 (N_17158,N_12199,N_14685);
xor U17159 (N_17159,N_12962,N_13759);
nor U17160 (N_17160,N_14295,N_12610);
nand U17161 (N_17161,N_12465,N_13461);
or U17162 (N_17162,N_13080,N_14266);
and U17163 (N_17163,N_14205,N_12164);
or U17164 (N_17164,N_14055,N_13927);
xnor U17165 (N_17165,N_14924,N_13644);
nor U17166 (N_17166,N_12639,N_12522);
or U17167 (N_17167,N_14701,N_14816);
xor U17168 (N_17168,N_13620,N_13791);
xor U17169 (N_17169,N_12874,N_14080);
nor U17170 (N_17170,N_12164,N_12878);
and U17171 (N_17171,N_12316,N_13808);
and U17172 (N_17172,N_14239,N_13007);
or U17173 (N_17173,N_12840,N_14630);
and U17174 (N_17174,N_12444,N_13655);
and U17175 (N_17175,N_12202,N_12861);
xnor U17176 (N_17176,N_14651,N_12916);
nand U17177 (N_17177,N_14831,N_13831);
nand U17178 (N_17178,N_14028,N_12307);
nor U17179 (N_17179,N_12428,N_13639);
or U17180 (N_17180,N_13914,N_12771);
or U17181 (N_17181,N_12381,N_14444);
nand U17182 (N_17182,N_12177,N_12839);
or U17183 (N_17183,N_13238,N_14955);
nand U17184 (N_17184,N_13159,N_13556);
nand U17185 (N_17185,N_14817,N_14983);
xor U17186 (N_17186,N_14533,N_14285);
nand U17187 (N_17187,N_13755,N_12430);
or U17188 (N_17188,N_14149,N_13000);
nand U17189 (N_17189,N_13663,N_13429);
or U17190 (N_17190,N_12270,N_12131);
nand U17191 (N_17191,N_14421,N_12087);
xnor U17192 (N_17192,N_13644,N_13045);
or U17193 (N_17193,N_13174,N_12426);
xor U17194 (N_17194,N_12517,N_12459);
nand U17195 (N_17195,N_12316,N_14605);
and U17196 (N_17196,N_14408,N_12349);
nor U17197 (N_17197,N_13907,N_12225);
nor U17198 (N_17198,N_13149,N_13300);
nor U17199 (N_17199,N_12741,N_12021);
or U17200 (N_17200,N_14145,N_13460);
nand U17201 (N_17201,N_12259,N_12058);
and U17202 (N_17202,N_13503,N_13667);
nand U17203 (N_17203,N_13965,N_12041);
xor U17204 (N_17204,N_13366,N_13946);
xor U17205 (N_17205,N_13362,N_12792);
xnor U17206 (N_17206,N_14384,N_14487);
and U17207 (N_17207,N_13831,N_12901);
or U17208 (N_17208,N_14063,N_12694);
nor U17209 (N_17209,N_12295,N_14753);
nand U17210 (N_17210,N_14606,N_13163);
or U17211 (N_17211,N_13203,N_12238);
xor U17212 (N_17212,N_14317,N_13203);
nor U17213 (N_17213,N_14398,N_13149);
nor U17214 (N_17214,N_13023,N_12476);
nand U17215 (N_17215,N_14555,N_13638);
nand U17216 (N_17216,N_14863,N_13235);
nand U17217 (N_17217,N_14642,N_14324);
and U17218 (N_17218,N_12916,N_12505);
nor U17219 (N_17219,N_12797,N_14490);
and U17220 (N_17220,N_13145,N_13841);
and U17221 (N_17221,N_14210,N_12046);
xor U17222 (N_17222,N_14889,N_12960);
or U17223 (N_17223,N_13089,N_13848);
or U17224 (N_17224,N_12830,N_14963);
and U17225 (N_17225,N_12921,N_12161);
nand U17226 (N_17226,N_14644,N_12215);
nor U17227 (N_17227,N_12628,N_14104);
nand U17228 (N_17228,N_12064,N_13856);
nor U17229 (N_17229,N_12860,N_14744);
nand U17230 (N_17230,N_12275,N_12682);
xor U17231 (N_17231,N_14256,N_13554);
nand U17232 (N_17232,N_13814,N_13684);
nor U17233 (N_17233,N_13516,N_14588);
and U17234 (N_17234,N_13042,N_13435);
nor U17235 (N_17235,N_13430,N_12970);
xor U17236 (N_17236,N_14512,N_12855);
nand U17237 (N_17237,N_14322,N_14391);
and U17238 (N_17238,N_14407,N_12306);
and U17239 (N_17239,N_14899,N_12043);
nor U17240 (N_17240,N_13229,N_12657);
nand U17241 (N_17241,N_13419,N_13787);
nand U17242 (N_17242,N_13583,N_14253);
and U17243 (N_17243,N_14270,N_12196);
or U17244 (N_17244,N_14351,N_14542);
or U17245 (N_17245,N_12176,N_13718);
xor U17246 (N_17246,N_13648,N_12990);
nand U17247 (N_17247,N_13600,N_13701);
xnor U17248 (N_17248,N_12534,N_12985);
xnor U17249 (N_17249,N_12180,N_14192);
xnor U17250 (N_17250,N_13631,N_14258);
nand U17251 (N_17251,N_12474,N_12229);
xor U17252 (N_17252,N_12070,N_14418);
or U17253 (N_17253,N_14341,N_12001);
xor U17254 (N_17254,N_12764,N_12592);
and U17255 (N_17255,N_13326,N_13065);
nand U17256 (N_17256,N_12786,N_14516);
or U17257 (N_17257,N_13079,N_12663);
or U17258 (N_17258,N_13716,N_14407);
nand U17259 (N_17259,N_14738,N_14807);
or U17260 (N_17260,N_12298,N_12263);
nor U17261 (N_17261,N_12951,N_13413);
and U17262 (N_17262,N_12191,N_12587);
nor U17263 (N_17263,N_14758,N_14388);
or U17264 (N_17264,N_13349,N_14885);
nand U17265 (N_17265,N_12838,N_12559);
nand U17266 (N_17266,N_12021,N_14869);
nor U17267 (N_17267,N_13534,N_13423);
nand U17268 (N_17268,N_14918,N_12638);
and U17269 (N_17269,N_12064,N_12013);
nand U17270 (N_17270,N_14404,N_13629);
or U17271 (N_17271,N_14211,N_12578);
or U17272 (N_17272,N_12151,N_14770);
nand U17273 (N_17273,N_14315,N_12597);
nor U17274 (N_17274,N_13925,N_14561);
or U17275 (N_17275,N_13323,N_14566);
nor U17276 (N_17276,N_13269,N_13912);
and U17277 (N_17277,N_13469,N_13270);
nor U17278 (N_17278,N_12596,N_12210);
and U17279 (N_17279,N_13224,N_14307);
or U17280 (N_17280,N_13801,N_14789);
or U17281 (N_17281,N_14330,N_14443);
or U17282 (N_17282,N_12861,N_12903);
and U17283 (N_17283,N_14032,N_12435);
and U17284 (N_17284,N_12302,N_14222);
or U17285 (N_17285,N_13596,N_14103);
nor U17286 (N_17286,N_14945,N_12201);
nand U17287 (N_17287,N_12094,N_14524);
xnor U17288 (N_17288,N_13036,N_12345);
or U17289 (N_17289,N_12302,N_14714);
or U17290 (N_17290,N_12519,N_12293);
nand U17291 (N_17291,N_14893,N_13712);
nor U17292 (N_17292,N_13777,N_14455);
nor U17293 (N_17293,N_13668,N_12750);
and U17294 (N_17294,N_12638,N_14974);
nor U17295 (N_17295,N_13978,N_13293);
or U17296 (N_17296,N_12155,N_13171);
nor U17297 (N_17297,N_13075,N_12369);
and U17298 (N_17298,N_14254,N_13454);
or U17299 (N_17299,N_14362,N_12966);
xor U17300 (N_17300,N_12361,N_12122);
nor U17301 (N_17301,N_12233,N_13489);
nand U17302 (N_17302,N_13271,N_13890);
or U17303 (N_17303,N_12160,N_13863);
xor U17304 (N_17304,N_12831,N_12628);
nor U17305 (N_17305,N_13988,N_14855);
nand U17306 (N_17306,N_14255,N_13813);
nor U17307 (N_17307,N_12374,N_14886);
or U17308 (N_17308,N_12395,N_13677);
and U17309 (N_17309,N_13222,N_14129);
xnor U17310 (N_17310,N_12144,N_12211);
xnor U17311 (N_17311,N_13605,N_13201);
nor U17312 (N_17312,N_12214,N_12477);
and U17313 (N_17313,N_13157,N_14801);
or U17314 (N_17314,N_12919,N_12430);
nor U17315 (N_17315,N_14154,N_12413);
and U17316 (N_17316,N_13199,N_12264);
or U17317 (N_17317,N_12366,N_14388);
xor U17318 (N_17318,N_13080,N_14524);
nand U17319 (N_17319,N_12069,N_14101);
xnor U17320 (N_17320,N_13302,N_13892);
xnor U17321 (N_17321,N_13706,N_14053);
xor U17322 (N_17322,N_13262,N_13611);
nor U17323 (N_17323,N_12349,N_13215);
and U17324 (N_17324,N_12677,N_12168);
nor U17325 (N_17325,N_14389,N_13977);
and U17326 (N_17326,N_14386,N_14583);
nor U17327 (N_17327,N_12587,N_14368);
xnor U17328 (N_17328,N_13816,N_12589);
xnor U17329 (N_17329,N_12727,N_13504);
or U17330 (N_17330,N_13103,N_13858);
xnor U17331 (N_17331,N_12771,N_14963);
and U17332 (N_17332,N_12555,N_14301);
xnor U17333 (N_17333,N_12985,N_13649);
nand U17334 (N_17334,N_14989,N_14617);
nand U17335 (N_17335,N_13209,N_14681);
nand U17336 (N_17336,N_13495,N_13842);
nand U17337 (N_17337,N_14490,N_14227);
xnor U17338 (N_17338,N_12022,N_12875);
and U17339 (N_17339,N_12576,N_14109);
xnor U17340 (N_17340,N_12386,N_14220);
nand U17341 (N_17341,N_12729,N_13706);
nor U17342 (N_17342,N_13337,N_13229);
and U17343 (N_17343,N_12819,N_12361);
and U17344 (N_17344,N_14560,N_12471);
xor U17345 (N_17345,N_14069,N_13537);
and U17346 (N_17346,N_13853,N_14621);
xnor U17347 (N_17347,N_13431,N_13624);
and U17348 (N_17348,N_14812,N_14575);
or U17349 (N_17349,N_12718,N_13539);
nand U17350 (N_17350,N_14638,N_13882);
nand U17351 (N_17351,N_12722,N_12867);
or U17352 (N_17352,N_14367,N_14218);
nor U17353 (N_17353,N_13698,N_12921);
nor U17354 (N_17354,N_13571,N_12516);
nor U17355 (N_17355,N_14377,N_13492);
nor U17356 (N_17356,N_14169,N_13927);
xor U17357 (N_17357,N_12628,N_12090);
nor U17358 (N_17358,N_12129,N_14690);
or U17359 (N_17359,N_12963,N_14455);
and U17360 (N_17360,N_12073,N_14186);
or U17361 (N_17361,N_12708,N_12817);
nand U17362 (N_17362,N_12387,N_12855);
xor U17363 (N_17363,N_14514,N_14890);
or U17364 (N_17364,N_12268,N_12698);
nand U17365 (N_17365,N_13057,N_14390);
and U17366 (N_17366,N_13155,N_12675);
or U17367 (N_17367,N_14474,N_13707);
and U17368 (N_17368,N_13131,N_13692);
nor U17369 (N_17369,N_13611,N_14417);
nor U17370 (N_17370,N_13792,N_14451);
and U17371 (N_17371,N_13190,N_13601);
or U17372 (N_17372,N_12716,N_13498);
or U17373 (N_17373,N_12234,N_12826);
nand U17374 (N_17374,N_12777,N_12759);
nor U17375 (N_17375,N_14972,N_13537);
nor U17376 (N_17376,N_12479,N_14506);
or U17377 (N_17377,N_12079,N_12431);
and U17378 (N_17378,N_14620,N_13404);
and U17379 (N_17379,N_13633,N_14371);
or U17380 (N_17380,N_12946,N_13721);
or U17381 (N_17381,N_14500,N_12971);
nand U17382 (N_17382,N_14920,N_12685);
and U17383 (N_17383,N_13002,N_12636);
nand U17384 (N_17384,N_13539,N_14084);
nand U17385 (N_17385,N_13169,N_12570);
xor U17386 (N_17386,N_13404,N_12404);
nor U17387 (N_17387,N_14577,N_13260);
and U17388 (N_17388,N_13949,N_12037);
xnor U17389 (N_17389,N_14871,N_13330);
or U17390 (N_17390,N_12490,N_12596);
nand U17391 (N_17391,N_14626,N_12716);
nor U17392 (N_17392,N_13332,N_13050);
nor U17393 (N_17393,N_13588,N_13700);
nor U17394 (N_17394,N_12157,N_12155);
nor U17395 (N_17395,N_14865,N_14735);
nand U17396 (N_17396,N_12602,N_12819);
and U17397 (N_17397,N_13199,N_13657);
and U17398 (N_17398,N_13749,N_14146);
nand U17399 (N_17399,N_13149,N_13018);
or U17400 (N_17400,N_14063,N_12285);
or U17401 (N_17401,N_12465,N_14194);
nand U17402 (N_17402,N_12886,N_14652);
nand U17403 (N_17403,N_14720,N_12020);
nand U17404 (N_17404,N_13687,N_12942);
or U17405 (N_17405,N_12791,N_13260);
nand U17406 (N_17406,N_13904,N_13892);
and U17407 (N_17407,N_14723,N_12752);
xor U17408 (N_17408,N_14742,N_13548);
nor U17409 (N_17409,N_12402,N_12812);
or U17410 (N_17410,N_13093,N_14376);
nand U17411 (N_17411,N_14871,N_14194);
nor U17412 (N_17412,N_14614,N_14298);
or U17413 (N_17413,N_14732,N_12977);
or U17414 (N_17414,N_14441,N_12930);
nand U17415 (N_17415,N_14837,N_13646);
nand U17416 (N_17416,N_14010,N_14646);
and U17417 (N_17417,N_13987,N_13129);
xor U17418 (N_17418,N_12487,N_14597);
and U17419 (N_17419,N_12022,N_14931);
nor U17420 (N_17420,N_12178,N_12581);
and U17421 (N_17421,N_12732,N_14645);
nand U17422 (N_17422,N_13638,N_14869);
or U17423 (N_17423,N_14140,N_13999);
or U17424 (N_17424,N_12693,N_12783);
or U17425 (N_17425,N_14029,N_12658);
nand U17426 (N_17426,N_13028,N_12604);
or U17427 (N_17427,N_12031,N_14687);
nand U17428 (N_17428,N_14974,N_12491);
xor U17429 (N_17429,N_12502,N_12915);
xor U17430 (N_17430,N_12187,N_13749);
and U17431 (N_17431,N_13766,N_14049);
nor U17432 (N_17432,N_14339,N_12415);
nand U17433 (N_17433,N_13184,N_12249);
xnor U17434 (N_17434,N_13824,N_14190);
and U17435 (N_17435,N_13608,N_12347);
xnor U17436 (N_17436,N_14996,N_14373);
or U17437 (N_17437,N_14073,N_12995);
and U17438 (N_17438,N_13303,N_12866);
and U17439 (N_17439,N_14242,N_12199);
nand U17440 (N_17440,N_13077,N_12472);
or U17441 (N_17441,N_13132,N_14530);
nand U17442 (N_17442,N_14963,N_13928);
and U17443 (N_17443,N_14466,N_12323);
nand U17444 (N_17444,N_13821,N_13500);
nand U17445 (N_17445,N_13208,N_13613);
or U17446 (N_17446,N_12577,N_13903);
and U17447 (N_17447,N_12572,N_14950);
nand U17448 (N_17448,N_13570,N_13928);
nor U17449 (N_17449,N_12573,N_13548);
nand U17450 (N_17450,N_12063,N_13146);
nor U17451 (N_17451,N_12834,N_14785);
or U17452 (N_17452,N_12543,N_12083);
xnor U17453 (N_17453,N_13086,N_14059);
xor U17454 (N_17454,N_14205,N_13143);
nand U17455 (N_17455,N_13622,N_13951);
nor U17456 (N_17456,N_14933,N_14577);
xor U17457 (N_17457,N_12853,N_12317);
and U17458 (N_17458,N_13062,N_14827);
nor U17459 (N_17459,N_14289,N_13416);
or U17460 (N_17460,N_12838,N_13539);
or U17461 (N_17461,N_14677,N_13882);
nor U17462 (N_17462,N_12019,N_12414);
and U17463 (N_17463,N_13957,N_13602);
nor U17464 (N_17464,N_14370,N_12887);
or U17465 (N_17465,N_14853,N_13448);
nor U17466 (N_17466,N_12697,N_14618);
xnor U17467 (N_17467,N_14291,N_13883);
and U17468 (N_17468,N_14121,N_12130);
xor U17469 (N_17469,N_14878,N_14641);
nand U17470 (N_17470,N_13486,N_14594);
xor U17471 (N_17471,N_14478,N_14791);
xnor U17472 (N_17472,N_14249,N_14167);
or U17473 (N_17473,N_14331,N_13725);
nand U17474 (N_17474,N_12547,N_14138);
and U17475 (N_17475,N_13901,N_12851);
or U17476 (N_17476,N_13401,N_12108);
and U17477 (N_17477,N_12907,N_14559);
and U17478 (N_17478,N_13344,N_13050);
nand U17479 (N_17479,N_13721,N_12998);
or U17480 (N_17480,N_14585,N_12057);
and U17481 (N_17481,N_14255,N_14920);
xor U17482 (N_17482,N_14800,N_13189);
nand U17483 (N_17483,N_14534,N_14700);
and U17484 (N_17484,N_12168,N_14024);
nand U17485 (N_17485,N_14008,N_13191);
xnor U17486 (N_17486,N_12877,N_12455);
or U17487 (N_17487,N_12503,N_12289);
or U17488 (N_17488,N_13981,N_13728);
or U17489 (N_17489,N_13131,N_12044);
nor U17490 (N_17490,N_12693,N_14755);
xnor U17491 (N_17491,N_12613,N_13611);
nand U17492 (N_17492,N_14136,N_13950);
and U17493 (N_17493,N_13499,N_12710);
and U17494 (N_17494,N_14308,N_14946);
and U17495 (N_17495,N_13066,N_13623);
nand U17496 (N_17496,N_12249,N_14235);
nand U17497 (N_17497,N_14799,N_13915);
nor U17498 (N_17498,N_13309,N_12922);
xor U17499 (N_17499,N_12720,N_12214);
and U17500 (N_17500,N_12518,N_13001);
xor U17501 (N_17501,N_13385,N_14620);
and U17502 (N_17502,N_13431,N_13312);
nor U17503 (N_17503,N_12838,N_12020);
nor U17504 (N_17504,N_14546,N_12536);
and U17505 (N_17505,N_13518,N_13054);
and U17506 (N_17506,N_12362,N_13030);
nor U17507 (N_17507,N_14164,N_13361);
nor U17508 (N_17508,N_13510,N_12188);
nor U17509 (N_17509,N_12080,N_13480);
nand U17510 (N_17510,N_12051,N_12405);
nor U17511 (N_17511,N_13611,N_14725);
and U17512 (N_17512,N_14965,N_13177);
and U17513 (N_17513,N_13709,N_13218);
nor U17514 (N_17514,N_12956,N_14108);
nand U17515 (N_17515,N_14699,N_12093);
and U17516 (N_17516,N_13429,N_14289);
and U17517 (N_17517,N_13555,N_13250);
xor U17518 (N_17518,N_12568,N_13513);
or U17519 (N_17519,N_12446,N_14985);
and U17520 (N_17520,N_13910,N_12471);
nand U17521 (N_17521,N_14443,N_12668);
or U17522 (N_17522,N_12805,N_14453);
nor U17523 (N_17523,N_13295,N_12277);
nor U17524 (N_17524,N_12929,N_13109);
and U17525 (N_17525,N_14395,N_13452);
nor U17526 (N_17526,N_12139,N_12461);
nor U17527 (N_17527,N_12884,N_13217);
xor U17528 (N_17528,N_14026,N_12797);
nor U17529 (N_17529,N_14456,N_13376);
nor U17530 (N_17530,N_13865,N_14638);
and U17531 (N_17531,N_14803,N_13632);
nor U17532 (N_17532,N_12124,N_13412);
xnor U17533 (N_17533,N_12548,N_12365);
or U17534 (N_17534,N_14242,N_14167);
xor U17535 (N_17535,N_13598,N_14216);
xnor U17536 (N_17536,N_12122,N_12724);
nor U17537 (N_17537,N_14711,N_14358);
nor U17538 (N_17538,N_14176,N_14831);
and U17539 (N_17539,N_12564,N_14694);
or U17540 (N_17540,N_12354,N_14946);
or U17541 (N_17541,N_12456,N_13968);
xor U17542 (N_17542,N_12931,N_12031);
and U17543 (N_17543,N_14119,N_13217);
or U17544 (N_17544,N_12374,N_12546);
xnor U17545 (N_17545,N_12118,N_13029);
nor U17546 (N_17546,N_12358,N_12412);
or U17547 (N_17547,N_12788,N_12619);
or U17548 (N_17548,N_14748,N_14693);
or U17549 (N_17549,N_13189,N_14897);
xnor U17550 (N_17550,N_12130,N_14970);
xnor U17551 (N_17551,N_14258,N_13451);
nor U17552 (N_17552,N_12829,N_12935);
xor U17553 (N_17553,N_13246,N_14887);
nand U17554 (N_17554,N_12388,N_12300);
or U17555 (N_17555,N_14613,N_12721);
xor U17556 (N_17556,N_13603,N_14412);
xnor U17557 (N_17557,N_14406,N_14214);
xnor U17558 (N_17558,N_13090,N_12376);
nand U17559 (N_17559,N_13832,N_13478);
or U17560 (N_17560,N_13836,N_13817);
nor U17561 (N_17561,N_14652,N_14564);
nor U17562 (N_17562,N_14192,N_14649);
and U17563 (N_17563,N_12115,N_13919);
nor U17564 (N_17564,N_12905,N_14365);
xnor U17565 (N_17565,N_14534,N_14717);
nand U17566 (N_17566,N_12760,N_13330);
or U17567 (N_17567,N_12659,N_12224);
nand U17568 (N_17568,N_13582,N_13129);
nor U17569 (N_17569,N_13784,N_13288);
xor U17570 (N_17570,N_12058,N_14274);
and U17571 (N_17571,N_13278,N_12147);
xor U17572 (N_17572,N_13436,N_13485);
nor U17573 (N_17573,N_13406,N_12255);
nand U17574 (N_17574,N_13808,N_14623);
or U17575 (N_17575,N_13588,N_12952);
nand U17576 (N_17576,N_14550,N_13516);
or U17577 (N_17577,N_13654,N_12227);
nor U17578 (N_17578,N_14228,N_14039);
nand U17579 (N_17579,N_13599,N_14973);
or U17580 (N_17580,N_12110,N_14012);
xor U17581 (N_17581,N_14658,N_13129);
xor U17582 (N_17582,N_13920,N_13114);
xnor U17583 (N_17583,N_12061,N_13312);
nor U17584 (N_17584,N_13945,N_14028);
and U17585 (N_17585,N_13628,N_13110);
nand U17586 (N_17586,N_13589,N_14297);
nor U17587 (N_17587,N_14093,N_14460);
nand U17588 (N_17588,N_12438,N_13092);
xor U17589 (N_17589,N_14840,N_12405);
and U17590 (N_17590,N_14567,N_12030);
nor U17591 (N_17591,N_12886,N_13031);
or U17592 (N_17592,N_12529,N_12622);
and U17593 (N_17593,N_13482,N_13973);
nor U17594 (N_17594,N_14717,N_12922);
or U17595 (N_17595,N_14355,N_12963);
nand U17596 (N_17596,N_12714,N_13077);
or U17597 (N_17597,N_14684,N_14306);
xor U17598 (N_17598,N_12692,N_14951);
and U17599 (N_17599,N_13814,N_13742);
nand U17600 (N_17600,N_13311,N_12150);
xor U17601 (N_17601,N_14345,N_12977);
xnor U17602 (N_17602,N_13316,N_13449);
xnor U17603 (N_17603,N_13312,N_12774);
or U17604 (N_17604,N_13813,N_14087);
xor U17605 (N_17605,N_13842,N_12810);
nand U17606 (N_17606,N_13257,N_14920);
nor U17607 (N_17607,N_14135,N_14314);
nand U17608 (N_17608,N_12574,N_14925);
and U17609 (N_17609,N_12174,N_13827);
or U17610 (N_17610,N_13367,N_14216);
nor U17611 (N_17611,N_14224,N_13429);
nor U17612 (N_17612,N_13649,N_13635);
nor U17613 (N_17613,N_13469,N_12238);
nand U17614 (N_17614,N_12344,N_12447);
or U17615 (N_17615,N_13924,N_12000);
or U17616 (N_17616,N_12169,N_14069);
or U17617 (N_17617,N_12212,N_13748);
nor U17618 (N_17618,N_14559,N_12002);
and U17619 (N_17619,N_14916,N_14073);
or U17620 (N_17620,N_12243,N_14816);
xnor U17621 (N_17621,N_14668,N_13587);
nand U17622 (N_17622,N_13864,N_12828);
xnor U17623 (N_17623,N_13541,N_14217);
and U17624 (N_17624,N_13717,N_14880);
xor U17625 (N_17625,N_13710,N_14205);
or U17626 (N_17626,N_13010,N_14426);
nor U17627 (N_17627,N_13564,N_12976);
nor U17628 (N_17628,N_12270,N_14705);
nand U17629 (N_17629,N_12600,N_14478);
xnor U17630 (N_17630,N_14059,N_14672);
or U17631 (N_17631,N_13296,N_14549);
or U17632 (N_17632,N_12421,N_12263);
or U17633 (N_17633,N_12955,N_13258);
nand U17634 (N_17634,N_12331,N_13826);
nand U17635 (N_17635,N_12534,N_13904);
and U17636 (N_17636,N_13375,N_12235);
and U17637 (N_17637,N_12064,N_13697);
or U17638 (N_17638,N_12822,N_12618);
nand U17639 (N_17639,N_14609,N_13060);
xnor U17640 (N_17640,N_13680,N_14737);
xnor U17641 (N_17641,N_14967,N_13566);
or U17642 (N_17642,N_13901,N_12940);
or U17643 (N_17643,N_13440,N_13194);
or U17644 (N_17644,N_14878,N_12587);
nand U17645 (N_17645,N_14015,N_13081);
and U17646 (N_17646,N_14486,N_14852);
or U17647 (N_17647,N_13666,N_13197);
xnor U17648 (N_17648,N_12229,N_12742);
nand U17649 (N_17649,N_13427,N_13843);
nor U17650 (N_17650,N_14992,N_12756);
or U17651 (N_17651,N_12717,N_13466);
xnor U17652 (N_17652,N_13143,N_12539);
and U17653 (N_17653,N_12805,N_12990);
xnor U17654 (N_17654,N_12086,N_12396);
xnor U17655 (N_17655,N_12956,N_14604);
and U17656 (N_17656,N_12954,N_13093);
or U17657 (N_17657,N_14374,N_12761);
and U17658 (N_17658,N_14890,N_13900);
xnor U17659 (N_17659,N_12207,N_14139);
and U17660 (N_17660,N_12811,N_12588);
nand U17661 (N_17661,N_12285,N_12849);
and U17662 (N_17662,N_12581,N_12004);
or U17663 (N_17663,N_13410,N_14832);
or U17664 (N_17664,N_12137,N_13899);
nor U17665 (N_17665,N_12483,N_12919);
nand U17666 (N_17666,N_14852,N_13007);
xnor U17667 (N_17667,N_12061,N_12742);
nand U17668 (N_17668,N_12991,N_13607);
nor U17669 (N_17669,N_12163,N_13541);
or U17670 (N_17670,N_14140,N_13730);
xnor U17671 (N_17671,N_13965,N_14155);
nand U17672 (N_17672,N_14938,N_14057);
nand U17673 (N_17673,N_13430,N_12362);
nor U17674 (N_17674,N_13151,N_14961);
and U17675 (N_17675,N_14720,N_12360);
or U17676 (N_17676,N_12200,N_14044);
and U17677 (N_17677,N_13588,N_12756);
xor U17678 (N_17678,N_13287,N_13373);
or U17679 (N_17679,N_13385,N_13174);
xnor U17680 (N_17680,N_13527,N_14840);
nor U17681 (N_17681,N_12788,N_13631);
xnor U17682 (N_17682,N_14809,N_13277);
and U17683 (N_17683,N_12009,N_13545);
nor U17684 (N_17684,N_13539,N_13987);
nor U17685 (N_17685,N_14907,N_13294);
xor U17686 (N_17686,N_12701,N_13687);
or U17687 (N_17687,N_12261,N_14916);
nor U17688 (N_17688,N_13767,N_12827);
and U17689 (N_17689,N_12959,N_12669);
nand U17690 (N_17690,N_12783,N_12087);
nand U17691 (N_17691,N_14933,N_14203);
nor U17692 (N_17692,N_13807,N_14460);
xnor U17693 (N_17693,N_13860,N_13260);
or U17694 (N_17694,N_13337,N_12573);
nor U17695 (N_17695,N_12067,N_12142);
nand U17696 (N_17696,N_14110,N_12197);
nor U17697 (N_17697,N_14092,N_12350);
xnor U17698 (N_17698,N_12283,N_14806);
nand U17699 (N_17699,N_12953,N_12704);
xor U17700 (N_17700,N_14674,N_13718);
or U17701 (N_17701,N_14511,N_13780);
and U17702 (N_17702,N_12080,N_14991);
nor U17703 (N_17703,N_12509,N_14165);
and U17704 (N_17704,N_12244,N_14023);
nor U17705 (N_17705,N_12400,N_14528);
or U17706 (N_17706,N_12026,N_14367);
or U17707 (N_17707,N_14331,N_12811);
nand U17708 (N_17708,N_13113,N_14618);
nor U17709 (N_17709,N_12399,N_13843);
nor U17710 (N_17710,N_12322,N_14663);
and U17711 (N_17711,N_13051,N_13249);
xor U17712 (N_17712,N_14608,N_13524);
xnor U17713 (N_17713,N_14940,N_13734);
nand U17714 (N_17714,N_14014,N_14032);
or U17715 (N_17715,N_13628,N_13051);
nor U17716 (N_17716,N_12753,N_13541);
nor U17717 (N_17717,N_13149,N_12852);
xnor U17718 (N_17718,N_14763,N_13075);
and U17719 (N_17719,N_13530,N_13587);
or U17720 (N_17720,N_13395,N_12964);
nor U17721 (N_17721,N_12398,N_12852);
nand U17722 (N_17722,N_12940,N_14964);
and U17723 (N_17723,N_14303,N_14936);
and U17724 (N_17724,N_13999,N_12679);
nand U17725 (N_17725,N_12614,N_14243);
xnor U17726 (N_17726,N_13786,N_14352);
nor U17727 (N_17727,N_12739,N_13570);
xnor U17728 (N_17728,N_14077,N_13230);
and U17729 (N_17729,N_14138,N_13590);
and U17730 (N_17730,N_13620,N_14406);
xor U17731 (N_17731,N_13424,N_12783);
nor U17732 (N_17732,N_14466,N_13368);
xor U17733 (N_17733,N_13997,N_13721);
xnor U17734 (N_17734,N_14365,N_13348);
nand U17735 (N_17735,N_14381,N_14984);
and U17736 (N_17736,N_12898,N_12656);
nor U17737 (N_17737,N_13730,N_12984);
and U17738 (N_17738,N_13242,N_13029);
nor U17739 (N_17739,N_13766,N_13787);
xnor U17740 (N_17740,N_14622,N_13101);
nor U17741 (N_17741,N_13453,N_13328);
xor U17742 (N_17742,N_14773,N_12925);
or U17743 (N_17743,N_13006,N_12703);
or U17744 (N_17744,N_12177,N_12686);
nand U17745 (N_17745,N_12959,N_14892);
nor U17746 (N_17746,N_14211,N_13929);
xnor U17747 (N_17747,N_13153,N_14191);
and U17748 (N_17748,N_13800,N_12654);
or U17749 (N_17749,N_12716,N_14070);
or U17750 (N_17750,N_14244,N_12102);
xor U17751 (N_17751,N_14946,N_13571);
nor U17752 (N_17752,N_14415,N_13014);
nand U17753 (N_17753,N_14858,N_13479);
and U17754 (N_17754,N_12938,N_14495);
and U17755 (N_17755,N_12544,N_12121);
or U17756 (N_17756,N_12643,N_13609);
nor U17757 (N_17757,N_14124,N_14318);
nor U17758 (N_17758,N_13754,N_13702);
nand U17759 (N_17759,N_14586,N_14537);
xnor U17760 (N_17760,N_12994,N_13008);
xor U17761 (N_17761,N_12684,N_13101);
xnor U17762 (N_17762,N_12289,N_13125);
nand U17763 (N_17763,N_13138,N_13130);
xor U17764 (N_17764,N_14256,N_13650);
xor U17765 (N_17765,N_12957,N_13258);
nand U17766 (N_17766,N_12943,N_12551);
nand U17767 (N_17767,N_14529,N_14867);
or U17768 (N_17768,N_13661,N_12597);
nor U17769 (N_17769,N_13424,N_14176);
nor U17770 (N_17770,N_12440,N_12562);
nor U17771 (N_17771,N_13866,N_13926);
nand U17772 (N_17772,N_12877,N_14240);
nand U17773 (N_17773,N_14273,N_13859);
and U17774 (N_17774,N_14044,N_13950);
xnor U17775 (N_17775,N_14222,N_12314);
nor U17776 (N_17776,N_14701,N_13912);
and U17777 (N_17777,N_12354,N_13023);
nor U17778 (N_17778,N_14613,N_12837);
nor U17779 (N_17779,N_13761,N_12707);
and U17780 (N_17780,N_14473,N_14271);
nand U17781 (N_17781,N_14851,N_12572);
and U17782 (N_17782,N_12997,N_12291);
nor U17783 (N_17783,N_14209,N_14694);
or U17784 (N_17784,N_12248,N_14949);
xnor U17785 (N_17785,N_13914,N_14719);
nand U17786 (N_17786,N_13510,N_12603);
xor U17787 (N_17787,N_12607,N_12077);
nand U17788 (N_17788,N_13293,N_13620);
nor U17789 (N_17789,N_13101,N_12811);
nand U17790 (N_17790,N_12022,N_14625);
nor U17791 (N_17791,N_12187,N_13954);
nand U17792 (N_17792,N_12844,N_13452);
or U17793 (N_17793,N_12103,N_12282);
xor U17794 (N_17794,N_14176,N_12570);
nor U17795 (N_17795,N_14048,N_14750);
nor U17796 (N_17796,N_13927,N_12874);
or U17797 (N_17797,N_12092,N_12125);
xnor U17798 (N_17798,N_14393,N_12931);
nand U17799 (N_17799,N_13465,N_12800);
xnor U17800 (N_17800,N_14924,N_13447);
nand U17801 (N_17801,N_12071,N_12444);
nor U17802 (N_17802,N_13366,N_14304);
or U17803 (N_17803,N_12768,N_14450);
xor U17804 (N_17804,N_14020,N_12235);
nand U17805 (N_17805,N_12568,N_14409);
and U17806 (N_17806,N_12196,N_13810);
xor U17807 (N_17807,N_12160,N_14386);
nor U17808 (N_17808,N_14031,N_13874);
nand U17809 (N_17809,N_13813,N_12523);
or U17810 (N_17810,N_13354,N_13211);
xnor U17811 (N_17811,N_13533,N_14487);
nor U17812 (N_17812,N_12834,N_13180);
xor U17813 (N_17813,N_14579,N_12067);
nand U17814 (N_17814,N_13039,N_13073);
or U17815 (N_17815,N_13912,N_13846);
or U17816 (N_17816,N_13132,N_14372);
xnor U17817 (N_17817,N_12855,N_13611);
or U17818 (N_17818,N_14819,N_14502);
nor U17819 (N_17819,N_13594,N_13157);
or U17820 (N_17820,N_14017,N_13598);
and U17821 (N_17821,N_13543,N_12707);
and U17822 (N_17822,N_13358,N_13019);
and U17823 (N_17823,N_13114,N_13014);
nor U17824 (N_17824,N_12046,N_13343);
xnor U17825 (N_17825,N_12730,N_13133);
nand U17826 (N_17826,N_13811,N_14215);
nand U17827 (N_17827,N_14330,N_13241);
nor U17828 (N_17828,N_14069,N_14267);
nor U17829 (N_17829,N_13066,N_14786);
nor U17830 (N_17830,N_14924,N_12300);
xor U17831 (N_17831,N_13812,N_13116);
and U17832 (N_17832,N_12188,N_12545);
xor U17833 (N_17833,N_14952,N_13119);
or U17834 (N_17834,N_13124,N_14566);
and U17835 (N_17835,N_13060,N_12694);
nor U17836 (N_17836,N_14204,N_13376);
or U17837 (N_17837,N_13654,N_12395);
and U17838 (N_17838,N_13305,N_14502);
xnor U17839 (N_17839,N_12261,N_13350);
and U17840 (N_17840,N_12510,N_14777);
and U17841 (N_17841,N_14683,N_14794);
nand U17842 (N_17842,N_14383,N_12968);
xnor U17843 (N_17843,N_14551,N_12840);
nand U17844 (N_17844,N_12403,N_12887);
xnor U17845 (N_17845,N_13990,N_14090);
nand U17846 (N_17846,N_12752,N_12390);
and U17847 (N_17847,N_12313,N_13370);
and U17848 (N_17848,N_13289,N_12495);
nand U17849 (N_17849,N_13128,N_14162);
xnor U17850 (N_17850,N_13579,N_12585);
xor U17851 (N_17851,N_14595,N_13006);
nor U17852 (N_17852,N_12732,N_13090);
nand U17853 (N_17853,N_12078,N_14721);
nand U17854 (N_17854,N_13562,N_14799);
or U17855 (N_17855,N_12488,N_14089);
nand U17856 (N_17856,N_14570,N_12128);
and U17857 (N_17857,N_14810,N_12573);
and U17858 (N_17858,N_12331,N_12384);
nor U17859 (N_17859,N_13863,N_12690);
xor U17860 (N_17860,N_12879,N_13692);
xor U17861 (N_17861,N_14142,N_12372);
nand U17862 (N_17862,N_13768,N_13587);
or U17863 (N_17863,N_13510,N_14088);
nor U17864 (N_17864,N_13669,N_14200);
xor U17865 (N_17865,N_12667,N_12254);
or U17866 (N_17866,N_12166,N_13954);
nand U17867 (N_17867,N_13707,N_13617);
nor U17868 (N_17868,N_14812,N_12781);
and U17869 (N_17869,N_12975,N_13617);
nand U17870 (N_17870,N_14907,N_12136);
xnor U17871 (N_17871,N_12883,N_14969);
and U17872 (N_17872,N_12580,N_13260);
and U17873 (N_17873,N_13454,N_12731);
xnor U17874 (N_17874,N_12200,N_12274);
xnor U17875 (N_17875,N_13558,N_13807);
and U17876 (N_17876,N_14264,N_12221);
and U17877 (N_17877,N_13588,N_12904);
and U17878 (N_17878,N_12223,N_12297);
and U17879 (N_17879,N_14599,N_14065);
xnor U17880 (N_17880,N_13876,N_14057);
nor U17881 (N_17881,N_13825,N_13498);
or U17882 (N_17882,N_12985,N_13942);
and U17883 (N_17883,N_13867,N_12311);
nand U17884 (N_17884,N_12501,N_14459);
xor U17885 (N_17885,N_13021,N_12741);
nand U17886 (N_17886,N_13387,N_13782);
xnor U17887 (N_17887,N_12118,N_12549);
or U17888 (N_17888,N_12781,N_13363);
and U17889 (N_17889,N_12267,N_12653);
nand U17890 (N_17890,N_12149,N_12145);
nor U17891 (N_17891,N_12886,N_14889);
and U17892 (N_17892,N_12566,N_14026);
xnor U17893 (N_17893,N_12709,N_13483);
and U17894 (N_17894,N_14551,N_13718);
and U17895 (N_17895,N_13120,N_13048);
and U17896 (N_17896,N_12806,N_12440);
and U17897 (N_17897,N_14314,N_12524);
xor U17898 (N_17898,N_13709,N_13461);
nand U17899 (N_17899,N_14777,N_12268);
and U17900 (N_17900,N_14284,N_13386);
and U17901 (N_17901,N_12850,N_12205);
nor U17902 (N_17902,N_12499,N_12782);
nand U17903 (N_17903,N_14319,N_13531);
nand U17904 (N_17904,N_14789,N_12281);
nor U17905 (N_17905,N_13320,N_12949);
nand U17906 (N_17906,N_14605,N_12001);
nand U17907 (N_17907,N_14243,N_12067);
xor U17908 (N_17908,N_13621,N_14281);
and U17909 (N_17909,N_13374,N_13864);
nand U17910 (N_17910,N_14051,N_14736);
xor U17911 (N_17911,N_13225,N_14517);
nand U17912 (N_17912,N_12637,N_14650);
xor U17913 (N_17913,N_12466,N_14694);
nand U17914 (N_17914,N_14552,N_13430);
nand U17915 (N_17915,N_12109,N_13960);
nand U17916 (N_17916,N_12484,N_13754);
xnor U17917 (N_17917,N_12638,N_13161);
or U17918 (N_17918,N_12735,N_13780);
and U17919 (N_17919,N_12969,N_12532);
nand U17920 (N_17920,N_14646,N_13983);
xnor U17921 (N_17921,N_12522,N_13612);
and U17922 (N_17922,N_12856,N_12146);
nand U17923 (N_17923,N_12846,N_14904);
nor U17924 (N_17924,N_13000,N_13461);
xnor U17925 (N_17925,N_13703,N_13663);
and U17926 (N_17926,N_14504,N_13841);
nand U17927 (N_17927,N_13405,N_13871);
nand U17928 (N_17928,N_12129,N_14472);
nor U17929 (N_17929,N_14116,N_12239);
nor U17930 (N_17930,N_13748,N_12312);
nand U17931 (N_17931,N_13191,N_12208);
nor U17932 (N_17932,N_14829,N_13235);
nand U17933 (N_17933,N_12707,N_13996);
nor U17934 (N_17934,N_14223,N_14140);
xor U17935 (N_17935,N_12220,N_12316);
nor U17936 (N_17936,N_13232,N_12007);
nand U17937 (N_17937,N_14286,N_12565);
nor U17938 (N_17938,N_12270,N_14418);
nand U17939 (N_17939,N_13938,N_12976);
nor U17940 (N_17940,N_12372,N_14599);
or U17941 (N_17941,N_12437,N_12607);
xor U17942 (N_17942,N_14266,N_14804);
nor U17943 (N_17943,N_12277,N_13437);
nor U17944 (N_17944,N_13860,N_14115);
and U17945 (N_17945,N_14509,N_14820);
xor U17946 (N_17946,N_14614,N_12172);
and U17947 (N_17947,N_12162,N_12951);
nand U17948 (N_17948,N_14095,N_12278);
nand U17949 (N_17949,N_12667,N_12851);
or U17950 (N_17950,N_13108,N_14971);
and U17951 (N_17951,N_12505,N_12281);
nor U17952 (N_17952,N_14739,N_12139);
or U17953 (N_17953,N_14050,N_12389);
or U17954 (N_17954,N_14550,N_13130);
nand U17955 (N_17955,N_14337,N_12577);
nand U17956 (N_17956,N_14537,N_12893);
xor U17957 (N_17957,N_14835,N_14042);
or U17958 (N_17958,N_13693,N_14894);
or U17959 (N_17959,N_12170,N_12446);
or U17960 (N_17960,N_13705,N_13090);
xnor U17961 (N_17961,N_12585,N_12009);
and U17962 (N_17962,N_13813,N_13330);
xor U17963 (N_17963,N_12567,N_12697);
nand U17964 (N_17964,N_13139,N_13431);
or U17965 (N_17965,N_13968,N_13508);
nand U17966 (N_17966,N_13046,N_14793);
and U17967 (N_17967,N_14803,N_13974);
and U17968 (N_17968,N_14437,N_12370);
xnor U17969 (N_17969,N_14148,N_12238);
xnor U17970 (N_17970,N_12387,N_13190);
and U17971 (N_17971,N_13410,N_13078);
nor U17972 (N_17972,N_14259,N_13680);
xor U17973 (N_17973,N_14183,N_12444);
or U17974 (N_17974,N_12263,N_12406);
nor U17975 (N_17975,N_12531,N_14517);
or U17976 (N_17976,N_13847,N_13937);
nand U17977 (N_17977,N_13057,N_14423);
nor U17978 (N_17978,N_12976,N_14177);
and U17979 (N_17979,N_14869,N_14905);
and U17980 (N_17980,N_13375,N_14852);
or U17981 (N_17981,N_13067,N_14008);
nor U17982 (N_17982,N_14955,N_14977);
and U17983 (N_17983,N_14668,N_12921);
and U17984 (N_17984,N_13679,N_13965);
or U17985 (N_17985,N_12712,N_12404);
nand U17986 (N_17986,N_13778,N_13075);
xor U17987 (N_17987,N_14554,N_12399);
nor U17988 (N_17988,N_13256,N_12695);
nand U17989 (N_17989,N_12522,N_14007);
or U17990 (N_17990,N_14890,N_14832);
or U17991 (N_17991,N_14632,N_13595);
and U17992 (N_17992,N_12228,N_14773);
xor U17993 (N_17993,N_14369,N_14939);
and U17994 (N_17994,N_14965,N_12186);
xor U17995 (N_17995,N_12303,N_13409);
and U17996 (N_17996,N_12074,N_13014);
xnor U17997 (N_17997,N_12728,N_13594);
xnor U17998 (N_17998,N_14919,N_13581);
or U17999 (N_17999,N_13300,N_14012);
nand U18000 (N_18000,N_16701,N_16245);
and U18001 (N_18001,N_16135,N_15677);
and U18002 (N_18002,N_15055,N_16306);
or U18003 (N_18003,N_16722,N_15756);
or U18004 (N_18004,N_15169,N_15872);
xnor U18005 (N_18005,N_15237,N_17337);
nor U18006 (N_18006,N_17861,N_15998);
nor U18007 (N_18007,N_15278,N_16630);
nand U18008 (N_18008,N_17726,N_17524);
nor U18009 (N_18009,N_16996,N_15087);
nor U18010 (N_18010,N_16379,N_16700);
or U18011 (N_18011,N_15528,N_16443);
nand U18012 (N_18012,N_17187,N_17910);
and U18013 (N_18013,N_16965,N_17918);
nand U18014 (N_18014,N_15880,N_16896);
and U18015 (N_18015,N_16961,N_16102);
nor U18016 (N_18016,N_16865,N_15916);
nand U18017 (N_18017,N_15956,N_16403);
nor U18018 (N_18018,N_17755,N_15754);
or U18019 (N_18019,N_15355,N_17076);
or U18020 (N_18020,N_16442,N_16811);
nor U18021 (N_18021,N_17090,N_15639);
xor U18022 (N_18022,N_16252,N_15137);
and U18023 (N_18023,N_15127,N_16385);
xor U18024 (N_18024,N_15682,N_16480);
nand U18025 (N_18025,N_17807,N_15808);
or U18026 (N_18026,N_16613,N_17385);
and U18027 (N_18027,N_17749,N_17701);
and U18028 (N_18028,N_17848,N_15707);
nor U18029 (N_18029,N_17556,N_15630);
or U18030 (N_18030,N_17388,N_15969);
and U18031 (N_18031,N_15233,N_16827);
nor U18032 (N_18032,N_15035,N_15256);
nor U18033 (N_18033,N_15176,N_17546);
and U18034 (N_18034,N_15503,N_17885);
xnor U18035 (N_18035,N_17793,N_15687);
or U18036 (N_18036,N_17395,N_16161);
or U18037 (N_18037,N_17014,N_16649);
xnor U18038 (N_18038,N_15920,N_17510);
nand U18039 (N_18039,N_15668,N_16163);
xor U18040 (N_18040,N_15941,N_15504);
xnor U18041 (N_18041,N_16978,N_17302);
nand U18042 (N_18042,N_15519,N_15710);
or U18043 (N_18043,N_15244,N_16511);
and U18044 (N_18044,N_17597,N_17651);
xnor U18045 (N_18045,N_16348,N_17340);
nor U18046 (N_18046,N_17485,N_16046);
nor U18047 (N_18047,N_17901,N_17877);
nand U18048 (N_18048,N_17012,N_15307);
nor U18049 (N_18049,N_16971,N_17784);
xor U18050 (N_18050,N_17528,N_17938);
or U18051 (N_18051,N_17627,N_15840);
or U18052 (N_18052,N_17205,N_15304);
xor U18053 (N_18053,N_17874,N_17600);
nand U18054 (N_18054,N_16880,N_17121);
and U18055 (N_18055,N_15726,N_16512);
and U18056 (N_18056,N_15581,N_15767);
xor U18057 (N_18057,N_17212,N_15182);
and U18058 (N_18058,N_15994,N_17046);
or U18059 (N_18059,N_17206,N_16429);
and U18060 (N_18060,N_17890,N_17278);
or U18061 (N_18061,N_15225,N_15138);
and U18062 (N_18062,N_16851,N_16713);
xnor U18063 (N_18063,N_16593,N_17330);
xnor U18064 (N_18064,N_17441,N_15220);
nor U18065 (N_18065,N_16980,N_16795);
and U18066 (N_18066,N_15255,N_17378);
nor U18067 (N_18067,N_16693,N_17465);
or U18068 (N_18068,N_17355,N_17350);
or U18069 (N_18069,N_17345,N_15522);
and U18070 (N_18070,N_17326,N_16242);
or U18071 (N_18071,N_16424,N_16397);
nand U18072 (N_18072,N_16190,N_16502);
and U18073 (N_18073,N_16782,N_15796);
or U18074 (N_18074,N_16938,N_16372);
and U18075 (N_18075,N_16300,N_16453);
or U18076 (N_18076,N_16285,N_16193);
nor U18077 (N_18077,N_16121,N_15243);
and U18078 (N_18078,N_17899,N_16903);
nand U18079 (N_18079,N_17349,N_16665);
nor U18080 (N_18080,N_15624,N_15399);
nor U18081 (N_18081,N_15569,N_16493);
or U18082 (N_18082,N_17935,N_16947);
xor U18083 (N_18083,N_15080,N_16714);
or U18084 (N_18084,N_16181,N_17564);
xor U18085 (N_18085,N_15972,N_16092);
nand U18086 (N_18086,N_17751,N_15029);
nand U18087 (N_18087,N_17280,N_16157);
and U18088 (N_18088,N_16038,N_15172);
nor U18089 (N_18089,N_17599,N_15531);
nor U18090 (N_18090,N_16617,N_16755);
nor U18091 (N_18091,N_16094,N_15798);
or U18092 (N_18092,N_17480,N_15868);
or U18093 (N_18093,N_16670,N_17027);
and U18094 (N_18094,N_15006,N_15902);
or U18095 (N_18095,N_17748,N_17773);
nand U18096 (N_18096,N_15621,N_16262);
and U18097 (N_18097,N_17715,N_17710);
and U18098 (N_18098,N_15913,N_17975);
xnor U18099 (N_18099,N_15812,N_15986);
nand U18100 (N_18100,N_16384,N_15893);
or U18101 (N_18101,N_15724,N_17450);
xor U18102 (N_18102,N_16249,N_16779);
nor U18103 (N_18103,N_17131,N_15146);
xor U18104 (N_18104,N_17942,N_15303);
nor U18105 (N_18105,N_17057,N_16439);
or U18106 (N_18106,N_17342,N_15082);
nor U18107 (N_18107,N_16077,N_17661);
nor U18108 (N_18108,N_16095,N_16072);
or U18109 (N_18109,N_17903,N_16726);
nand U18110 (N_18110,N_17936,N_15934);
xnor U18111 (N_18111,N_17018,N_15075);
and U18112 (N_18112,N_17353,N_15269);
xnor U18113 (N_18113,N_16552,N_16998);
or U18114 (N_18114,N_16118,N_16205);
and U18115 (N_18115,N_16934,N_17718);
xor U18116 (N_18116,N_16198,N_15249);
nand U18117 (N_18117,N_15235,N_15928);
nand U18118 (N_18118,N_16796,N_16414);
or U18119 (N_18119,N_16745,N_15856);
nor U18120 (N_18120,N_16603,N_16197);
or U18121 (N_18121,N_16660,N_15715);
nand U18122 (N_18122,N_16476,N_16967);
and U18123 (N_18123,N_16818,N_17507);
or U18124 (N_18124,N_16555,N_17282);
or U18125 (N_18125,N_16800,N_16567);
nor U18126 (N_18126,N_15215,N_17292);
nand U18127 (N_18127,N_16224,N_17503);
and U18128 (N_18128,N_16661,N_17428);
and U18129 (N_18129,N_16082,N_16776);
xnor U18130 (N_18130,N_15081,N_16330);
xnor U18131 (N_18131,N_16981,N_15953);
nand U18132 (N_18132,N_15449,N_17976);
nand U18133 (N_18133,N_16091,N_17258);
or U18134 (N_18134,N_15454,N_16199);
nor U18135 (N_18135,N_16211,N_17109);
xor U18136 (N_18136,N_17436,N_16069);
nand U18137 (N_18137,N_17454,N_17126);
xnor U18138 (N_18138,N_15136,N_17334);
and U18139 (N_18139,N_16410,N_15529);
xor U18140 (N_18140,N_17967,N_17895);
or U18141 (N_18141,N_17314,N_15592);
xor U18142 (N_18142,N_15482,N_15790);
and U18143 (N_18143,N_15362,N_15310);
or U18144 (N_18144,N_15978,N_16768);
or U18145 (N_18145,N_17338,N_15989);
xnor U18146 (N_18146,N_17692,N_16437);
xor U18147 (N_18147,N_15755,N_16604);
nand U18148 (N_18148,N_16635,N_17192);
or U18149 (N_18149,N_17409,N_16136);
nand U18150 (N_18150,N_15054,N_17298);
or U18151 (N_18151,N_16979,N_15466);
nor U18152 (N_18152,N_16957,N_17537);
nor U18153 (N_18153,N_17943,N_15842);
or U18154 (N_18154,N_16358,N_16332);
or U18155 (N_18155,N_17045,N_17218);
xnor U18156 (N_18156,N_16029,N_15234);
nor U18157 (N_18157,N_17137,N_16120);
or U18158 (N_18158,N_15188,N_15619);
xor U18159 (N_18159,N_17179,N_17794);
nand U18160 (N_18160,N_17888,N_17493);
xor U18161 (N_18161,N_16837,N_17707);
nor U18162 (N_18162,N_17495,N_15699);
xor U18163 (N_18163,N_17202,N_15321);
nor U18164 (N_18164,N_16498,N_17308);
xor U18165 (N_18165,N_16111,N_15031);
or U18166 (N_18166,N_17083,N_17028);
nor U18167 (N_18167,N_16844,N_15759);
xnor U18168 (N_18168,N_17889,N_15280);
nor U18169 (N_18169,N_17632,N_16342);
and U18170 (N_18170,N_16158,N_17226);
or U18171 (N_18171,N_17633,N_15047);
nor U18172 (N_18172,N_15486,N_15462);
nand U18173 (N_18173,N_17584,N_16001);
xor U18174 (N_18174,N_17184,N_16122);
nand U18175 (N_18175,N_15572,N_17115);
xor U18176 (N_18176,N_17367,N_16454);
xor U18177 (N_18177,N_16590,N_15882);
nand U18178 (N_18178,N_16011,N_17359);
and U18179 (N_18179,N_16902,N_16508);
nor U18180 (N_18180,N_17371,N_15252);
and U18181 (N_18181,N_16487,N_15871);
nand U18182 (N_18182,N_15982,N_16805);
and U18183 (N_18183,N_15465,N_15515);
nand U18184 (N_18184,N_15284,N_17419);
xor U18185 (N_18185,N_16033,N_15794);
nand U18186 (N_18186,N_16615,N_15210);
or U18187 (N_18187,N_16325,N_15479);
nand U18188 (N_18188,N_16803,N_16166);
or U18189 (N_18189,N_16043,N_16114);
or U18190 (N_18190,N_15923,N_15156);
xnor U18191 (N_18191,N_15720,N_16056);
nand U18192 (N_18192,N_16950,N_16201);
and U18193 (N_18193,N_16405,N_17044);
nand U18194 (N_18194,N_16337,N_15505);
or U18195 (N_18195,N_17864,N_15145);
xor U18196 (N_18196,N_16041,N_17674);
or U18197 (N_18197,N_15187,N_17102);
or U18198 (N_18198,N_17968,N_16380);
and U18199 (N_18199,N_15723,N_17132);
or U18200 (N_18200,N_15262,N_16290);
or U18201 (N_18201,N_15483,N_17081);
and U18202 (N_18202,N_17971,N_15866);
nand U18203 (N_18203,N_17396,N_17164);
nand U18204 (N_18204,N_16734,N_15890);
and U18205 (N_18205,N_17527,N_16129);
or U18206 (N_18206,N_17919,N_16840);
and U18207 (N_18207,N_16176,N_15068);
nand U18208 (N_18208,N_16892,N_15422);
and U18209 (N_18209,N_17303,N_17636);
and U18210 (N_18210,N_15020,N_17032);
xnor U18211 (N_18211,N_16537,N_16286);
nor U18212 (N_18212,N_17455,N_17365);
and U18213 (N_18213,N_17145,N_15478);
nor U18214 (N_18214,N_15057,N_15704);
or U18215 (N_18215,N_16601,N_16983);
nor U18216 (N_18216,N_17199,N_17249);
nand U18217 (N_18217,N_17035,N_16561);
nand U18218 (N_18218,N_17460,N_17194);
xnor U18219 (N_18219,N_15356,N_17228);
or U18220 (N_18220,N_16723,N_16448);
nand U18221 (N_18221,N_15543,N_16566);
nand U18222 (N_18222,N_17851,N_16756);
and U18223 (N_18223,N_17185,N_17065);
or U18224 (N_18224,N_15128,N_16172);
and U18225 (N_18225,N_15032,N_15556);
nand U18226 (N_18226,N_16107,N_16349);
xnor U18227 (N_18227,N_15589,N_15123);
nand U18228 (N_18228,N_15769,N_17621);
or U18229 (N_18229,N_16717,N_17769);
nand U18230 (N_18230,N_15011,N_17357);
xnor U18231 (N_18231,N_17135,N_15761);
nand U18232 (N_18232,N_15175,N_17497);
nand U18233 (N_18233,N_17117,N_16952);
nor U18234 (N_18234,N_17243,N_17312);
and U18235 (N_18235,N_17103,N_17050);
xnor U18236 (N_18236,N_16515,N_17760);
nor U18237 (N_18237,N_16625,N_17582);
xnor U18238 (N_18238,N_16110,N_16817);
or U18239 (N_18239,N_16706,N_15700);
nor U18240 (N_18240,N_16667,N_17991);
nor U18241 (N_18241,N_16562,N_17608);
and U18242 (N_18242,N_17849,N_17005);
xnor U18243 (N_18243,N_15410,N_17483);
nand U18244 (N_18244,N_16543,N_17703);
and U18245 (N_18245,N_15095,N_16912);
nand U18246 (N_18246,N_15268,N_17870);
xor U18247 (N_18247,N_17148,N_17125);
xnor U18248 (N_18248,N_16406,N_17729);
nand U18249 (N_18249,N_16207,N_15846);
nor U18250 (N_18250,N_16449,N_17149);
and U18251 (N_18251,N_16855,N_16654);
nand U18252 (N_18252,N_17411,N_16253);
nor U18253 (N_18253,N_15010,N_17679);
and U18254 (N_18254,N_17602,N_16452);
or U18255 (N_18255,N_17095,N_15990);
or U18256 (N_18256,N_16074,N_15258);
and U18257 (N_18257,N_17262,N_15048);
xnor U18258 (N_18258,N_17417,N_16113);
xnor U18259 (N_18259,N_17000,N_15766);
and U18260 (N_18260,N_17924,N_16145);
nand U18261 (N_18261,N_17315,N_17666);
nor U18262 (N_18262,N_17542,N_17697);
xor U18263 (N_18263,N_17172,N_17642);
and U18264 (N_18264,N_16875,N_15740);
xnor U18265 (N_18265,N_17623,N_15506);
xnor U18266 (N_18266,N_17295,N_16943);
nor U18267 (N_18267,N_17787,N_16382);
and U18268 (N_18268,N_17680,N_17138);
xor U18269 (N_18269,N_16391,N_17607);
xnor U18270 (N_18270,N_17394,N_15874);
xnor U18271 (N_18271,N_16160,N_17144);
xnor U18272 (N_18272,N_17306,N_17116);
and U18273 (N_18273,N_15167,N_17629);
and U18274 (N_18274,N_16749,N_15375);
nand U18275 (N_18275,N_15357,N_15413);
and U18276 (N_18276,N_15965,N_16637);
nand U18277 (N_18277,N_16150,N_16895);
and U18278 (N_18278,N_15491,N_16153);
xnor U18279 (N_18279,N_17423,N_17213);
and U18280 (N_18280,N_15932,N_17380);
or U18281 (N_18281,N_15312,N_17979);
and U18282 (N_18282,N_16521,N_17063);
and U18283 (N_18283,N_17550,N_15066);
xnor U18284 (N_18284,N_15405,N_15614);
or U18285 (N_18285,N_15885,N_15800);
nand U18286 (N_18286,N_16246,N_17802);
or U18287 (N_18287,N_15663,N_17959);
or U18288 (N_18288,N_17242,N_15587);
nand U18289 (N_18289,N_17384,N_16016);
xor U18290 (N_18290,N_17472,N_15636);
nor U18291 (N_18291,N_15660,N_15579);
and U18292 (N_18292,N_17168,N_16616);
nor U18293 (N_18293,N_15785,N_16576);
and U18294 (N_18294,N_17836,N_17830);
nor U18295 (N_18295,N_15634,N_16289);
and U18296 (N_18296,N_16142,N_15649);
nor U18297 (N_18297,N_15298,N_15226);
xnor U18298 (N_18298,N_17712,N_17796);
and U18299 (N_18299,N_17640,N_16856);
or U18300 (N_18300,N_15602,N_16341);
nand U18301 (N_18301,N_15148,N_17806);
xor U18302 (N_18302,N_16538,N_16640);
xnor U18303 (N_18303,N_17174,N_17171);
nand U18304 (N_18304,N_17084,N_17110);
and U18305 (N_18305,N_16731,N_15365);
or U18306 (N_18306,N_15900,N_16940);
nor U18307 (N_18307,N_16915,N_15052);
and U18308 (N_18308,N_16859,N_17934);
or U18309 (N_18309,N_17487,N_15461);
nor U18310 (N_18310,N_16139,N_15096);
and U18311 (N_18311,N_17853,N_15658);
xnor U18312 (N_18312,N_15381,N_17061);
or U18313 (N_18313,N_17949,N_15870);
nand U18314 (N_18314,N_15678,N_15977);
nand U18315 (N_18315,N_16832,N_16119);
xnor U18316 (N_18316,N_17316,N_17002);
and U18317 (N_18317,N_16293,N_16220);
nor U18318 (N_18318,N_17944,N_15536);
and U18319 (N_18319,N_16729,N_15196);
xnor U18320 (N_18320,N_15521,N_17559);
and U18321 (N_18321,N_17933,N_15714);
and U18322 (N_18322,N_17271,N_16581);
xnor U18323 (N_18323,N_15099,N_16557);
nor U18324 (N_18324,N_17620,N_17476);
nand U18325 (N_18325,N_15437,N_17800);
nor U18326 (N_18326,N_17927,N_17561);
nor U18327 (N_18327,N_15575,N_15523);
nand U18328 (N_18328,N_17047,N_15058);
nor U18329 (N_18329,N_16219,N_15626);
and U18330 (N_18330,N_17668,N_17469);
nor U18331 (N_18331,N_17157,N_17766);
nand U18332 (N_18332,N_16522,N_15014);
nand U18333 (N_18333,N_15946,N_17809);
and U18334 (N_18334,N_16079,N_15784);
nor U18335 (N_18335,N_15083,N_16564);
or U18336 (N_18336,N_17286,N_15816);
or U18337 (N_18337,N_16497,N_16783);
nand U18338 (N_18338,N_17225,N_16999);
and U18339 (N_18339,N_15013,N_17301);
nand U18340 (N_18340,N_17087,N_15933);
and U18341 (N_18341,N_17754,N_15371);
nor U18342 (N_18342,N_16707,N_17891);
or U18343 (N_18343,N_16222,N_17276);
and U18344 (N_18344,N_16824,N_15173);
and U18345 (N_18345,N_17630,N_17348);
xnor U18346 (N_18346,N_17190,N_16563);
xor U18347 (N_18347,N_17804,N_15878);
nand U18348 (N_18348,N_15727,N_17643);
nand U18349 (N_18349,N_15787,N_15997);
xor U18350 (N_18350,N_16462,N_15938);
nand U18351 (N_18351,N_17215,N_16802);
and U18352 (N_18352,N_15591,N_16968);
and U18353 (N_18353,N_17778,N_15595);
xnor U18354 (N_18354,N_15441,N_15993);
or U18355 (N_18355,N_16000,N_15867);
and U18356 (N_18356,N_16280,N_17579);
nor U18357 (N_18357,N_16048,N_17279);
nor U18358 (N_18358,N_15331,N_15161);
nor U18359 (N_18359,N_16156,N_17878);
xor U18360 (N_18360,N_17565,N_15108);
xnor U18361 (N_18361,N_17008,N_15984);
nand U18362 (N_18362,N_15180,N_16377);
xnor U18363 (N_18363,N_15223,N_15495);
nor U18364 (N_18364,N_15459,N_15251);
xor U18365 (N_18365,N_16678,N_16032);
nor U18366 (N_18366,N_17761,N_17129);
or U18367 (N_18367,N_15738,N_17641);
or U18368 (N_18368,N_17369,N_15493);
nor U18369 (N_18369,N_15670,N_15958);
and U18370 (N_18370,N_16314,N_16946);
nand U18371 (N_18371,N_17563,N_16598);
nand U18372 (N_18372,N_17331,N_17305);
or U18373 (N_18373,N_15527,N_15511);
nand U18374 (N_18374,N_17058,N_17739);
nand U18375 (N_18375,N_16993,N_15897);
nand U18376 (N_18376,N_15332,N_15174);
nand U18377 (N_18377,N_17745,N_16834);
and U18378 (N_18378,N_15545,N_15260);
and U18379 (N_18379,N_15289,N_15033);
nand U18380 (N_18380,N_16829,N_16657);
nand U18381 (N_18381,N_16434,N_16319);
nand U18382 (N_18382,N_16843,N_17956);
and U18383 (N_18383,N_17026,N_17850);
and U18384 (N_18384,N_17744,N_16527);
nand U18385 (N_18385,N_15910,N_17554);
nor U18386 (N_18386,N_15686,N_16230);
or U18387 (N_18387,N_17591,N_15203);
nor U18388 (N_18388,N_15214,N_16162);
nand U18389 (N_18389,N_15570,N_17248);
and U18390 (N_18390,N_17268,N_17275);
xor U18391 (N_18391,N_16404,N_15648);
nand U18392 (N_18392,N_17293,N_17624);
or U18393 (N_18393,N_15324,N_17819);
or U18394 (N_18394,N_15807,N_16910);
nor U18395 (N_18395,N_16928,N_16884);
and U18396 (N_18396,N_15447,N_17752);
nor U18397 (N_18397,N_17932,N_15899);
or U18398 (N_18398,N_17973,N_15016);
xor U18399 (N_18399,N_16730,N_17585);
and U18400 (N_18400,N_17731,N_16194);
or U18401 (N_18401,N_16422,N_16570);
xor U18402 (N_18402,N_16737,N_16954);
nor U18403 (N_18403,N_15396,N_17327);
xor U18404 (N_18404,N_16949,N_15949);
nand U18405 (N_18405,N_15774,N_15450);
nor U18406 (N_18406,N_15265,N_15320);
nand U18407 (N_18407,N_17952,N_16112);
nand U18408 (N_18408,N_17708,N_16408);
nor U18409 (N_18409,N_16184,N_15597);
nor U18410 (N_18410,N_15633,N_15186);
nor U18411 (N_18411,N_16468,N_15209);
and U18412 (N_18412,N_17558,N_15696);
and U18413 (N_18413,N_17658,N_15326);
xnor U18414 (N_18414,N_17031,N_16312);
or U18415 (N_18415,N_15440,N_17165);
nand U18416 (N_18416,N_16992,N_15758);
nand U18417 (N_18417,N_15420,N_16645);
nor U18418 (N_18418,N_16897,N_16235);
xnor U18419 (N_18419,N_16006,N_16815);
nand U18420 (N_18420,N_17788,N_15818);
or U18421 (N_18421,N_16945,N_16313);
and U18422 (N_18422,N_16492,N_15285);
nand U18423 (N_18423,N_15825,N_16258);
and U18424 (N_18424,N_17862,N_17015);
or U18425 (N_18425,N_17908,N_15344);
xor U18426 (N_18426,N_16247,N_17108);
and U18427 (N_18427,N_17209,N_17798);
xnor U18428 (N_18428,N_16504,N_17598);
nand U18429 (N_18429,N_17458,N_15526);
xor U18430 (N_18430,N_15829,N_16867);
or U18431 (N_18431,N_17984,N_15403);
nand U18432 (N_18432,N_16901,N_15361);
xor U18433 (N_18433,N_15603,N_15005);
and U18434 (N_18434,N_16232,N_15976);
nand U18435 (N_18435,N_15485,N_16799);
nor U18436 (N_18436,N_15004,N_16766);
or U18437 (N_18437,N_16316,N_17987);
xor U18438 (N_18438,N_17659,N_17053);
nor U18439 (N_18439,N_15747,N_16417);
nand U18440 (N_18440,N_17531,N_16676);
nand U18441 (N_18441,N_17650,N_15272);
or U18442 (N_18442,N_15151,N_15703);
nor U18443 (N_18443,N_16760,N_17586);
xnor U18444 (N_18444,N_16421,N_15929);
or U18445 (N_18445,N_15142,N_16320);
nor U18446 (N_18446,N_17930,N_15065);
or U18447 (N_18447,N_15921,N_15257);
or U18448 (N_18448,N_15101,N_16906);
nand U18449 (N_18449,N_15653,N_16012);
nor U18450 (N_18450,N_15317,N_16569);
nand U18451 (N_18451,N_17427,N_16970);
nand U18452 (N_18452,N_15364,N_17471);
nor U18453 (N_18453,N_17175,N_16283);
nor U18454 (N_18454,N_17776,N_16109);
xnor U18455 (N_18455,N_15426,N_16309);
nor U18456 (N_18456,N_16647,N_16689);
nor U18457 (N_18457,N_17551,N_15637);
nand U18458 (N_18458,N_17266,N_16845);
nand U18459 (N_18459,N_15078,N_17954);
nor U18460 (N_18460,N_16619,N_17368);
and U18461 (N_18461,N_16123,N_16057);
and U18462 (N_18462,N_16582,N_17432);
nand U18463 (N_18463,N_17593,N_15041);
nand U18464 (N_18464,N_16956,N_15673);
xnor U18465 (N_18465,N_17881,N_17287);
and U18466 (N_18466,N_15538,N_15091);
nand U18467 (N_18467,N_16592,N_17204);
nor U18468 (N_18468,N_16479,N_16644);
nor U18469 (N_18469,N_16386,N_15448);
nand U18470 (N_18470,N_15644,N_17086);
nor U18471 (N_18471,N_16683,N_17917);
nand U18472 (N_18472,N_16392,N_16777);
nand U18473 (N_18473,N_17705,N_16638);
nor U18474 (N_18474,N_15301,N_15692);
and U18475 (N_18475,N_16663,N_17902);
nor U18476 (N_18476,N_16271,N_15793);
or U18477 (N_18477,N_17894,N_15408);
xor U18478 (N_18478,N_16228,N_16535);
nor U18479 (N_18479,N_17897,N_16212);
xnor U18480 (N_18480,N_17310,N_17098);
xor U18481 (N_18481,N_16841,N_17962);
or U18482 (N_18482,N_17351,N_17082);
nor U18483 (N_18483,N_17505,N_17589);
xnor U18484 (N_18484,N_15132,N_17133);
nor U18485 (N_18485,N_16878,N_16752);
and U18486 (N_18486,N_17615,N_16798);
or U18487 (N_18487,N_17957,N_16624);
xnor U18488 (N_18488,N_17541,N_15778);
or U18489 (N_18489,N_17492,N_17609);
and U18490 (N_18490,N_17033,N_15042);
nor U18491 (N_18491,N_15951,N_16831);
xnor U18492 (N_18492,N_17547,N_16887);
or U18493 (N_18493,N_15473,N_15883);
and U18494 (N_18494,N_16296,N_16360);
nand U18495 (N_18495,N_15917,N_17681);
nand U18496 (N_18496,N_16060,N_16725);
nor U18497 (N_18497,N_16931,N_15114);
nand U18498 (N_18498,N_17412,N_17601);
and U18499 (N_18499,N_17964,N_17690);
or U18500 (N_18500,N_16338,N_17229);
nand U18501 (N_18501,N_16823,N_16869);
nor U18502 (N_18502,N_15814,N_16499);
nand U18503 (N_18503,N_15254,N_15959);
nand U18504 (N_18504,N_15957,N_17363);
and U18505 (N_18505,N_17222,N_16067);
and U18506 (N_18506,N_15021,N_17509);
or U18507 (N_18507,N_15906,N_15728);
xor U18508 (N_18508,N_17420,N_16456);
xor U18509 (N_18509,N_17970,N_17224);
nand U18510 (N_18510,N_15768,N_17843);
xnor U18511 (N_18511,N_16556,N_15788);
or U18512 (N_18512,N_15152,N_16472);
nand U18513 (N_18513,N_17685,N_15841);
or U18514 (N_18514,N_15105,N_15826);
xnor U18515 (N_18515,N_17141,N_16073);
nor U18516 (N_18516,N_17914,N_16668);
nand U18517 (N_18517,N_17223,N_15499);
and U18518 (N_18518,N_17288,N_15125);
nor U18519 (N_18519,N_16863,N_15157);
nand U18520 (N_18520,N_15566,N_16986);
or U18521 (N_18521,N_16727,N_17486);
nand U18522 (N_18522,N_16131,N_17038);
xnor U18523 (N_18523,N_15657,N_16496);
nor U18524 (N_18524,N_17594,N_17533);
and U18525 (N_18525,N_17844,N_17498);
nand U18526 (N_18526,N_16302,N_16955);
or U18527 (N_18527,N_17572,N_15467);
xor U18528 (N_18528,N_17198,N_15323);
or U18529 (N_18529,N_16475,N_16853);
xnor U18530 (N_18530,N_16732,N_16974);
or U18531 (N_18531,N_15501,N_15739);
and U18532 (N_18532,N_15039,N_16720);
or U18533 (N_18533,N_15084,N_16093);
and U18534 (N_18534,N_15373,N_16051);
nand U18535 (N_18535,N_17402,N_17415);
nand U18536 (N_18536,N_16491,N_15742);
nor U18537 (N_18537,N_17343,N_16927);
or U18538 (N_18538,N_16839,N_17191);
and U18539 (N_18539,N_17376,N_15776);
or U18540 (N_18540,N_16399,N_15974);
or U18541 (N_18541,N_16539,N_16010);
or U18542 (N_18542,N_16780,N_16771);
and U18543 (N_18543,N_17167,N_15008);
xnor U18544 (N_18544,N_17625,N_17734);
or U18545 (N_18545,N_17704,N_16500);
nand U18546 (N_18546,N_16825,N_16335);
nand U18547 (N_18547,N_16297,N_17473);
or U18548 (N_18548,N_16389,N_17667);
nand U18549 (N_18549,N_15551,N_16191);
xor U18550 (N_18550,N_17158,N_15424);
nand U18551 (N_18551,N_16466,N_15183);
xnor U18552 (N_18552,N_17398,N_15576);
nor U18553 (N_18553,N_17617,N_15019);
or U18554 (N_18554,N_16054,N_16872);
or U18555 (N_18555,N_16688,N_16044);
nor U18556 (N_18556,N_15983,N_16478);
and U18557 (N_18557,N_15073,N_15985);
and U18558 (N_18558,N_17182,N_15248);
xnor U18559 (N_18559,N_15185,N_15097);
nor U18560 (N_18560,N_17635,N_17255);
nor U18561 (N_18561,N_15313,N_17512);
or U18562 (N_18562,N_16239,N_16641);
nand U18563 (N_18563,N_15855,N_15227);
or U18564 (N_18564,N_17237,N_17173);
nand U18565 (N_18565,N_17457,N_15417);
nor U18566 (N_18566,N_16599,N_17577);
nor U18567 (N_18567,N_16510,N_16987);
nor U18568 (N_18568,N_17177,N_17618);
nor U18569 (N_18569,N_15760,N_15221);
nand U18570 (N_18570,N_16007,N_15571);
nor U18571 (N_18571,N_16550,N_17162);
nor U18572 (N_18572,N_15074,N_15231);
and U18573 (N_18573,N_17691,N_15126);
and U18574 (N_18574,N_16594,N_17783);
nand U18575 (N_18575,N_15701,N_15034);
xnor U18576 (N_18576,N_17817,N_15216);
nand U18577 (N_18577,N_15197,N_17818);
nor U18578 (N_18578,N_16708,N_15698);
nor U18579 (N_18579,N_15745,N_17246);
and U18580 (N_18580,N_17724,N_15198);
nand U18581 (N_18581,N_15530,N_16982);
xnor U18582 (N_18582,N_16886,N_17399);
xnor U18583 (N_18583,N_15232,N_16214);
or U18584 (N_18584,N_16618,N_17515);
nand U18585 (N_18585,N_15694,N_16365);
nor U18586 (N_18586,N_15201,N_16307);
nor U18587 (N_18587,N_16866,N_17040);
or U18588 (N_18588,N_16053,N_17810);
or U18589 (N_18589,N_17181,N_17325);
or U18590 (N_18590,N_17779,N_17662);
xnor U18591 (N_18591,N_17725,N_17088);
nand U18592 (N_18592,N_16764,N_15372);
xnor U18593 (N_18593,N_17346,N_15891);
or U18594 (N_18594,N_17328,N_17019);
or U18595 (N_18595,N_17834,N_16327);
nor U18596 (N_18596,N_16709,N_16165);
nand U18597 (N_18597,N_17863,N_16694);
xor U18598 (N_18598,N_17143,N_15553);
or U18599 (N_18599,N_15040,N_16573);
nand U18600 (N_18600,N_17277,N_16941);
and U18601 (N_18601,N_16607,N_16005);
nand U18602 (N_18602,N_16821,N_17759);
nand U18603 (N_18603,N_16888,N_15713);
xnor U18604 (N_18604,N_17433,N_15887);
or U18605 (N_18605,N_16259,N_15743);
xnor U18606 (N_18606,N_16423,N_17247);
and U18607 (N_18607,N_16097,N_17323);
nand U18608 (N_18608,N_16108,N_15432);
or U18609 (N_18609,N_16770,N_16216);
nand U18610 (N_18610,N_17926,N_15120);
nor U18611 (N_18611,N_17612,N_15554);
or U18612 (N_18612,N_15346,N_16256);
and U18613 (N_18613,N_15541,N_17413);
nand U18614 (N_18614,N_17152,N_16596);
xnor U18615 (N_18615,N_17387,N_15253);
nor U18616 (N_18616,N_17422,N_16105);
and U18617 (N_18617,N_15282,N_17682);
xor U18618 (N_18618,N_17079,N_17906);
and U18619 (N_18619,N_15434,N_17566);
or U18620 (N_18620,N_15291,N_16958);
xnor U18621 (N_18621,N_17146,N_15212);
nor U18622 (N_18622,N_15514,N_17442);
and U18623 (N_18623,N_16329,N_16907);
nand U18624 (N_18624,N_16809,N_15489);
nor U18625 (N_18625,N_15088,N_15160);
and U18626 (N_18626,N_15822,N_16140);
and U18627 (N_18627,N_15433,N_17921);
or U18628 (N_18628,N_15337,N_16292);
and U18629 (N_18629,N_15705,N_16045);
nand U18630 (N_18630,N_17525,N_16767);
nor U18631 (N_18631,N_17931,N_15349);
or U18632 (N_18632,N_16820,N_16432);
nand U18633 (N_18633,N_17136,N_16301);
nor U18634 (N_18634,N_15049,N_16769);
nand U18635 (N_18635,N_17405,N_16850);
and U18636 (N_18636,N_17735,N_16227);
nor U18637 (N_18637,N_15352,N_16765);
and U18638 (N_18638,N_16458,N_15245);
nor U18639 (N_18639,N_17475,N_16233);
nor U18640 (N_18640,N_15815,N_15667);
and U18641 (N_18641,N_15149,N_15286);
xnor U18642 (N_18642,N_15604,N_15401);
and U18643 (N_18643,N_16063,N_17321);
and U18644 (N_18644,N_16147,N_15409);
nand U18645 (N_18645,N_15999,N_15963);
xor U18646 (N_18646,N_15294,N_15488);
xor U18647 (N_18647,N_17085,N_15849);
nand U18648 (N_18648,N_16375,N_15343);
and U18649 (N_18649,N_16346,N_15416);
or U18650 (N_18650,N_15817,N_15338);
and U18651 (N_18651,N_16972,N_16168);
and U18652 (N_18652,N_17898,N_15139);
xor U18653 (N_18653,N_17464,N_16786);
nand U18654 (N_18654,N_15930,N_15051);
or U18655 (N_18655,N_16318,N_17251);
nor U18656 (N_18656,N_17039,N_17260);
xor U18657 (N_18657,N_16750,N_17812);
nand U18658 (N_18658,N_17997,N_17884);
and U18659 (N_18659,N_16620,N_16146);
or U18660 (N_18660,N_16642,N_17421);
or U18661 (N_18661,N_17813,N_16547);
nor U18662 (N_18662,N_16355,N_15070);
or U18663 (N_18663,N_17879,N_15753);
and U18664 (N_18664,N_15712,N_16368);
xnor U18665 (N_18665,N_15549,N_15943);
nand U18666 (N_18666,N_15915,N_15805);
and U18667 (N_18667,N_16482,N_16255);
nor U18668 (N_18668,N_15567,N_16340);
xnor U18669 (N_18669,N_15564,N_16751);
xor U18670 (N_18670,N_16807,N_17696);
or U18671 (N_18671,N_15555,N_15762);
nor U18672 (N_18672,N_16484,N_15446);
and U18673 (N_18673,N_17453,N_17900);
xor U18674 (N_18674,N_17447,N_15498);
and U18675 (N_18675,N_16464,N_15456);
nand U18676 (N_18676,N_16103,N_17780);
nand U18677 (N_18677,N_17448,N_16935);
nor U18678 (N_18678,N_16559,N_17837);
nor U18679 (N_18679,N_17443,N_15520);
nand U18680 (N_18680,N_16816,N_15045);
nand U18681 (N_18681,N_17827,N_16431);
xnor U18682 (N_18682,N_16261,N_17689);
and U18683 (N_18683,N_16636,N_17669);
xnor U18684 (N_18684,N_16533,N_16847);
nand U18685 (N_18685,N_17123,N_15927);
nor U18686 (N_18686,N_15009,N_15270);
nor U18687 (N_18687,N_15746,N_16913);
and U18688 (N_18688,N_16321,N_17245);
xor U18689 (N_18689,N_15907,N_15512);
xor U18690 (N_18690,N_15802,N_15423);
nor U18691 (N_18691,N_16412,N_16882);
or U18692 (N_18692,N_17151,N_16411);
xnor U18693 (N_18693,N_15539,N_17426);
or U18694 (N_18694,N_16849,N_15979);
or U18695 (N_18695,N_16876,N_16891);
nor U18696 (N_18696,N_17573,N_17553);
or U18697 (N_18697,N_15804,N_15862);
or U18698 (N_18698,N_16387,N_15327);
or U18699 (N_18699,N_17540,N_16898);
nand U18700 (N_18700,N_15370,N_17939);
or U18701 (N_18701,N_17216,N_16517);
or U18702 (N_18702,N_16206,N_16237);
nor U18703 (N_18703,N_17313,N_15610);
xnor U18704 (N_18704,N_16842,N_17758);
or U18705 (N_18705,N_16746,N_17297);
or U18706 (N_18706,N_16975,N_17880);
or U18707 (N_18707,N_17484,N_15366);
nor U18708 (N_18708,N_16461,N_17502);
nand U18709 (N_18709,N_17001,N_17960);
xor U18710 (N_18710,N_16583,N_15578);
or U18711 (N_18711,N_16273,N_17534);
and U18712 (N_18712,N_15908,N_16899);
xnor U18713 (N_18713,N_17341,N_16627);
or U18714 (N_18714,N_17922,N_16704);
and U18715 (N_18715,N_16506,N_16427);
xnor U18716 (N_18716,N_16666,N_16126);
or U18717 (N_18717,N_17709,N_16648);
xor U18718 (N_18718,N_17211,N_17883);
nor U18719 (N_18719,N_15017,N_16215);
nand U18720 (N_18720,N_17250,N_17781);
nand U18721 (N_18721,N_17264,N_16331);
or U18722 (N_18722,N_15411,N_15288);
nand U18723 (N_18723,N_16848,N_16277);
nor U18724 (N_18724,N_15721,N_15240);
nor U18725 (N_18725,N_17911,N_16804);
nand U18726 (N_18726,N_16083,N_15001);
nand U18727 (N_18727,N_16858,N_15067);
nor U18728 (N_18728,N_16361,N_15407);
or U18729 (N_18729,N_17360,N_16819);
nand U18730 (N_18730,N_16529,N_16835);
nor U18731 (N_18731,N_17071,N_16836);
nand U18732 (N_18732,N_17434,N_17474);
nor U18733 (N_18733,N_17815,N_17060);
xnor U18734 (N_18734,N_17730,N_17743);
and U18735 (N_18735,N_17339,N_16234);
xor U18736 (N_18736,N_16294,N_15922);
xnor U18737 (N_18737,N_15706,N_15189);
and U18738 (N_18738,N_16914,N_17056);
nor U18739 (N_18739,N_15468,N_17309);
nand U18740 (N_18740,N_15722,N_16806);
nor U18741 (N_18741,N_16366,N_17096);
nand U18742 (N_18742,N_17459,N_17267);
nor U18743 (N_18743,N_15025,N_16023);
nor U18744 (N_18744,N_15560,N_16513);
xnor U18745 (N_18745,N_17916,N_15732);
or U18746 (N_18746,N_17831,N_15190);
xnor U18747 (N_18747,N_15781,N_15909);
xor U18748 (N_18748,N_15302,N_17491);
or U18749 (N_18749,N_17406,N_17532);
xnor U18750 (N_18750,N_17768,N_17285);
nor U18751 (N_18751,N_16893,N_16420);
and U18752 (N_18752,N_16200,N_16463);
nand U18753 (N_18753,N_15605,N_15388);
and U18754 (N_18754,N_16838,N_15018);
xnor U18755 (N_18755,N_17361,N_15811);
or U18756 (N_18756,N_16930,N_16035);
nor U18757 (N_18757,N_15429,N_17720);
xnor U18758 (N_18758,N_15616,N_16602);
or U18759 (N_18759,N_17721,N_15588);
nand U18760 (N_18760,N_16268,N_15476);
or U18761 (N_18761,N_17477,N_15594);
and U18762 (N_18762,N_17066,N_17771);
nor U18763 (N_18763,N_17119,N_16339);
nand U18764 (N_18764,N_16225,N_17284);
or U18765 (N_18765,N_16177,N_17571);
or U18766 (N_18766,N_15651,N_16584);
nand U18767 (N_18767,N_17283,N_16440);
xor U18768 (N_18768,N_15618,N_16021);
nand U18769 (N_18769,N_17740,N_16632);
nor U18770 (N_18770,N_17166,N_16685);
and U18771 (N_18771,N_17741,N_16580);
nand U18772 (N_18772,N_17407,N_17189);
or U18773 (N_18773,N_15079,N_17011);
and U18774 (N_18774,N_16305,N_15502);
or U18775 (N_18775,N_15850,N_15904);
or U18776 (N_18776,N_16334,N_17451);
nand U18777 (N_18777,N_15532,N_15847);
or U18778 (N_18778,N_16474,N_15524);
nand U18779 (N_18779,N_16343,N_15022);
nor U18780 (N_18780,N_17538,N_17868);
xor U18781 (N_18781,N_15492,N_17677);
nor U18782 (N_18782,N_16020,N_17481);
nand U18783 (N_18783,N_16303,N_17947);
nand U18784 (N_18784,N_16002,N_15071);
nand U18785 (N_18785,N_16679,N_15333);
nand U18786 (N_18786,N_16352,N_17048);
nand U18787 (N_18787,N_15064,N_17857);
and U18788 (N_18788,N_16269,N_17291);
and U18789 (N_18789,N_17430,N_15107);
nor U18790 (N_18790,N_15803,N_16587);
nor U18791 (N_18791,N_16393,N_15632);
nand U18792 (N_18792,N_17240,N_16141);
nor U18793 (N_18793,N_17560,N_15470);
xnor U18794 (N_18794,N_17404,N_16773);
or U18795 (N_18795,N_16578,N_15876);
or U18796 (N_18796,N_16115,N_15056);
nand U18797 (N_18797,N_16467,N_16672);
nand U18798 (N_18798,N_15513,N_15683);
nor U18799 (N_18799,N_15497,N_17296);
xor U18800 (N_18800,N_15898,N_15295);
nor U18801 (N_18801,N_17606,N_16354);
xor U18802 (N_18802,N_17763,N_15736);
or U18803 (N_18803,N_15612,N_15092);
and U18804 (N_18804,N_16433,N_15463);
nand U18805 (N_18805,N_16278,N_15093);
nand U18806 (N_18806,N_15439,N_17329);
nor U18807 (N_18807,N_17713,N_17501);
and U18808 (N_18808,N_16985,N_15110);
xor U18809 (N_18809,N_15104,N_16551);
xor U18810 (N_18810,N_16742,N_17557);
nor U18811 (N_18811,N_16918,N_16098);
xor U18812 (N_18812,N_17847,N_15709);
or U18813 (N_18813,N_16167,N_16988);
nand U18814 (N_18814,N_15267,N_15222);
nand U18815 (N_18815,N_15119,N_17858);
and U18816 (N_18816,N_16741,N_17822);
xnor U18817 (N_18817,N_16681,N_16792);
nor U18818 (N_18818,N_16323,N_15770);
or U18819 (N_18819,N_17969,N_16812);
or U18820 (N_18820,N_16871,N_16116);
nor U18821 (N_18821,N_15028,N_15681);
xnor U18822 (N_18822,N_17333,N_15200);
nand U18823 (N_18823,N_17100,N_17153);
nor U18824 (N_18824,N_15389,N_16287);
nand U18825 (N_18825,N_17535,N_15444);
nor U18826 (N_18826,N_15402,N_16548);
nand U18827 (N_18827,N_15573,N_17139);
and U18828 (N_18828,N_16728,N_15266);
and U18829 (N_18829,N_15342,N_15708);
xnor U18830 (N_18830,N_17737,N_15797);
nor U18831 (N_18831,N_15378,N_15296);
xor U18832 (N_18832,N_15319,N_16132);
and U18833 (N_18833,N_16740,N_16560);
xor U18834 (N_18834,N_15995,N_17688);
nand U18835 (N_18835,N_16367,N_17238);
xnor U18836 (N_18836,N_15451,N_16003);
and U18837 (N_18837,N_15130,N_17099);
xor U18838 (N_18838,N_17403,N_17429);
or U18839 (N_18839,N_15398,N_16398);
and U18840 (N_18840,N_17281,N_15980);
nand U18841 (N_18841,N_15261,N_15274);
nor U18842 (N_18842,N_16034,N_17985);
or U18843 (N_18843,N_17826,N_16787);
nor U18844 (N_18844,N_16868,N_15044);
xor U18845 (N_18845,N_16061,N_16260);
xnor U18846 (N_18846,N_15397,N_15050);
xor U18847 (N_18847,N_15427,N_17114);
nand U18848 (N_18848,N_17049,N_16014);
nand U18849 (N_18849,N_17016,N_17294);
and U18850 (N_18850,N_16170,N_16407);
nor U18851 (N_18851,N_16675,N_16419);
nor U18852 (N_18852,N_16264,N_15775);
nand U18853 (N_18853,N_17257,N_16173);
and U18854 (N_18854,N_15455,N_16995);
or U18855 (N_18855,N_15368,N_16396);
nand U18856 (N_18856,N_16364,N_15643);
nand U18857 (N_18857,N_15336,N_16486);
xnor U18858 (N_18858,N_17992,N_15219);
nor U18859 (N_18859,N_16690,N_15379);
nor U18860 (N_18860,N_15211,N_16953);
xor U18861 (N_18861,N_15435,N_17774);
xor U18862 (N_18862,N_15955,N_15935);
nand U18863 (N_18863,N_16733,N_15043);
nand U18864 (N_18864,N_16267,N_15112);
or U18865 (N_18865,N_15358,N_15386);
and U18866 (N_18866,N_17996,N_17410);
xor U18867 (N_18867,N_15428,N_16217);
or U18868 (N_18868,N_15164,N_16789);
and U18869 (N_18869,N_16018,N_15425);
and U18870 (N_18870,N_16659,N_16413);
nand U18871 (N_18871,N_16171,N_16315);
and U18872 (N_18872,N_15936,N_15584);
nor U18873 (N_18873,N_15059,N_16295);
xor U18874 (N_18874,N_16646,N_16127);
or U18875 (N_18875,N_15918,N_16049);
and U18876 (N_18876,N_15675,N_15779);
nand U18877 (N_18877,N_16159,N_15359);
or U18878 (N_18878,N_15544,N_16549);
xor U18879 (N_18879,N_16310,N_15652);
and U18880 (N_18880,N_16076,N_15702);
xnor U18881 (N_18881,N_15496,N_16814);
nor U18882 (N_18882,N_17479,N_15559);
or U18883 (N_18883,N_16695,N_15911);
nor U18884 (N_18884,N_15077,N_15629);
xnor U18885 (N_18885,N_15574,N_17539);
nand U18886 (N_18886,N_17431,N_16944);
nor U18887 (N_18887,N_17445,N_17370);
xnor U18888 (N_18888,N_15580,N_15442);
and U18889 (N_18889,N_16775,N_16395);
or U18890 (N_18890,N_16208,N_15299);
xor U18891 (N_18891,N_15460,N_16736);
xor U18892 (N_18892,N_17366,N_15208);
nor U18893 (N_18893,N_15300,N_15824);
nor U18894 (N_18894,N_15195,N_16251);
nand U18895 (N_18895,N_16240,N_16025);
or U18896 (N_18896,N_16757,N_16748);
nor U18897 (N_18897,N_15679,N_16932);
and U18898 (N_18898,N_15480,N_16774);
nand U18899 (N_18899,N_16523,N_15283);
nand U18900 (N_18900,N_17080,N_17603);
nand U18901 (N_18901,N_17336,N_17183);
and U18902 (N_18902,N_17068,N_16009);
nor U18903 (N_18903,N_16236,N_17335);
nand U18904 (N_18904,N_15487,N_17318);
xor U18905 (N_18905,N_16179,N_15414);
nor U18906 (N_18906,N_16908,N_15383);
or U18907 (N_18907,N_16629,N_15737);
nand U18908 (N_18908,N_17094,N_17508);
or U18909 (N_18909,N_17698,N_17511);
or U18910 (N_18910,N_17188,N_15163);
nor U18911 (N_18911,N_16698,N_16650);
or U18912 (N_18912,N_17263,N_16705);
xor U18913 (N_18913,N_15641,N_16920);
xnor U18914 (N_18914,N_16794,N_16495);
nand U18915 (N_18915,N_16540,N_17762);
and U18916 (N_18916,N_17808,N_16436);
xor U18917 (N_18917,N_15672,N_16024);
or U18918 (N_18918,N_15948,N_16359);
or U18919 (N_18919,N_16042,N_17037);
xor U18920 (N_18920,N_16390,N_15582);
and U18921 (N_18921,N_17549,N_16860);
and U18922 (N_18922,N_16106,N_15242);
nand U18923 (N_18923,N_15436,N_17852);
or U18924 (N_18924,N_17521,N_16554);
and U18925 (N_18925,N_16401,N_17972);
nor U18926 (N_18926,N_16703,N_17180);
nand U18927 (N_18927,N_16244,N_17373);
nor U18928 (N_18928,N_16658,N_16611);
nor U18929 (N_18929,N_16070,N_15194);
or U18930 (N_18930,N_17953,N_16879);
xor U18931 (N_18931,N_17186,N_16558);
xor U18932 (N_18932,N_15015,N_15475);
nand U18933 (N_18933,N_17456,N_17785);
or U18934 (N_18934,N_17197,N_15400);
nor U18935 (N_18935,N_16738,N_15611);
xnor U18936 (N_18936,N_17062,N_15973);
nand U18937 (N_18937,N_17227,N_17489);
and U18938 (N_18938,N_17648,N_17974);
xnor U18939 (N_18939,N_15628,N_17886);
nor U18940 (N_18940,N_16862,N_15693);
nor U18941 (N_18941,N_15229,N_15676);
nand U18942 (N_18942,N_15664,N_15061);
or U18943 (N_18943,N_15140,N_17253);
or U18944 (N_18944,N_16164,N_15179);
and U18945 (N_18945,N_15162,N_15996);
or U18946 (N_18946,N_17522,N_16036);
nor U18947 (N_18947,N_17958,N_17169);
nand U18948 (N_18948,N_15952,N_15944);
xor U18949 (N_18949,N_16143,N_15865);
nand U18950 (N_18950,N_17887,N_15622);
xor U18951 (N_18951,N_17004,N_16013);
nand U18952 (N_18952,N_16977,N_15159);
or U18953 (N_18953,N_16857,N_16577);
nand U18954 (N_18954,N_16696,N_17723);
xnor U18955 (N_18955,N_16960,N_17506);
xnor U18956 (N_18956,N_15165,N_17256);
xor U18957 (N_18957,N_17665,N_15642);
nand U18958 (N_18958,N_16441,N_16631);
or U18959 (N_18959,N_17687,N_15860);
or U18960 (N_18960,N_15674,N_16605);
nor U18961 (N_18961,N_16250,N_17070);
xor U18962 (N_18962,N_15430,N_15599);
nor U18963 (N_18963,N_17803,N_17414);
nand U18964 (N_18964,N_15827,N_15277);
xnor U18965 (N_18965,N_17678,N_17319);
and U18966 (N_18966,N_15831,N_17221);
nand U18967 (N_18967,N_16526,N_15086);
or U18968 (N_18968,N_15150,N_15118);
xnor U18969 (N_18969,N_16963,N_15561);
and U18970 (N_18970,N_17344,N_15646);
nand U18971 (N_18971,N_15771,N_15819);
xor U18972 (N_18972,N_16925,N_16808);
xnor U18973 (N_18973,N_16545,N_15206);
xor U18974 (N_18974,N_17611,N_17234);
and U18975 (N_18975,N_16861,N_16791);
xnor U18976 (N_18976,N_16298,N_16050);
nand U18977 (N_18977,N_16909,N_17978);
xnor U18978 (N_18978,N_16671,N_17074);
and U18979 (N_18979,N_16883,N_15550);
nor U18980 (N_18980,N_17576,N_15547);
or U18981 (N_18981,N_17876,N_16152);
and U18982 (N_18982,N_16175,N_16553);
and U18983 (N_18983,N_16916,N_16459);
nand U18984 (N_18984,N_17244,N_15335);
nand U18985 (N_18985,N_16213,N_16402);
or U18986 (N_18986,N_16939,N_17647);
xnor U18987 (N_18987,N_16483,N_16394);
nand U18988 (N_18988,N_17986,N_15275);
nor U18989 (N_18989,N_16125,N_17220);
xor U18990 (N_18990,N_15443,N_16532);
or U18991 (N_18991,N_16444,N_16793);
nand U18992 (N_18992,N_17437,N_17239);
nand U18993 (N_18993,N_15689,N_15748);
nand U18994 (N_18994,N_17913,N_17882);
and U18995 (N_18995,N_15115,N_17529);
xnor U18996 (N_18996,N_17418,N_16536);
xnor U18997 (N_18997,N_17105,N_15931);
and U18998 (N_18998,N_17631,N_17989);
nor U18999 (N_18999,N_16192,N_17393);
xnor U19000 (N_19000,N_16080,N_16852);
nand U19001 (N_19001,N_16218,N_15586);
nor U19002 (N_19002,N_17628,N_16503);
or U19003 (N_19003,N_17616,N_15224);
or U19004 (N_19004,N_15508,N_15293);
xnor U19005 (N_19005,N_15109,N_15276);
and U19006 (N_19006,N_16133,N_16308);
xnor U19007 (N_19007,N_15510,N_17795);
xor U19008 (N_19008,N_17728,N_16610);
nand U19009 (N_19009,N_16052,N_16430);
nor U19010 (N_19010,N_17756,N_17995);
xnor U19011 (N_19011,N_16772,N_15177);
nand U19012 (N_19012,N_15102,N_15894);
nand U19013 (N_19013,N_17893,N_16317);
or U19014 (N_19014,N_16284,N_16008);
nor U19015 (N_19015,N_16609,N_16081);
nand U19016 (N_19016,N_16951,N_15828);
nor U19017 (N_19017,N_17570,N_17854);
xnor U19018 (N_19018,N_16881,N_17128);
or U19019 (N_19019,N_17929,N_17024);
nand U19020 (N_19020,N_17790,N_15236);
xnor U19021 (N_19021,N_15609,N_15650);
xnor U19022 (N_19022,N_15003,N_17961);
nor U19023 (N_19023,N_16047,N_17770);
and U19024 (N_19024,N_16275,N_15144);
or U19025 (N_19025,N_17867,N_16311);
nor U19026 (N_19026,N_16221,N_16677);
and U19027 (N_19027,N_17254,N_15950);
xnor U19028 (N_19028,N_15795,N_17928);
nor U19029 (N_19029,N_17828,N_17424);
or U19030 (N_19030,N_17866,N_15354);
nor U19031 (N_19031,N_15845,N_16575);
and U19032 (N_19032,N_15458,N_15391);
and U19033 (N_19033,N_16154,N_15729);
and U19034 (N_19034,N_16797,N_16196);
and U19035 (N_19035,N_16997,N_17439);
nor U19036 (N_19036,N_15863,N_17022);
nand U19037 (N_19037,N_15098,N_17552);
and U19038 (N_19038,N_15438,N_15085);
or U19039 (N_19039,N_17452,N_17657);
nor U19040 (N_19040,N_17289,N_17694);
xnor U19041 (N_19041,N_16291,N_17772);
nand U19042 (N_19042,N_15348,N_17777);
or U19043 (N_19043,N_17134,N_15171);
xor U19044 (N_19044,N_17990,N_16272);
xor U19045 (N_19045,N_15178,N_15117);
and U19046 (N_19046,N_16418,N_16662);
xnor U19047 (N_19047,N_17732,N_15690);
xnor U19048 (N_19048,N_17569,N_17236);
nor U19049 (N_19049,N_15864,N_17655);
xnor U19050 (N_19050,N_17782,N_16017);
nor U19051 (N_19051,N_17488,N_16064);
nor U19052 (N_19052,N_17377,N_17208);
xor U19053 (N_19053,N_17998,N_15002);
xnor U19054 (N_19054,N_15090,N_15246);
and U19055 (N_19055,N_17178,N_17307);
nand U19056 (N_19056,N_16055,N_15469);
nand U19057 (N_19057,N_15153,N_16565);
nor U19058 (N_19058,N_17142,N_16469);
xor U19059 (N_19059,N_15193,N_15471);
and U19060 (N_19060,N_17873,N_17683);
nor U19061 (N_19061,N_15263,N_16004);
nor U19062 (N_19062,N_15960,N_17416);
nand U19063 (N_19063,N_15548,N_16336);
and U19064 (N_19064,N_16905,N_15247);
nor U19065 (N_19065,N_17494,N_15158);
xnor U19066 (N_19066,N_17590,N_17383);
nor U19067 (N_19067,N_15757,N_15615);
nand U19068 (N_19068,N_15945,N_16989);
nand U19069 (N_19069,N_15852,N_15988);
nor U19070 (N_19070,N_17013,N_17671);
xor U19071 (N_19071,N_16270,N_16813);
and U19072 (N_19072,N_15837,N_17029);
xnor U19073 (N_19073,N_15947,N_15192);
nor U19074 (N_19074,N_16282,N_17120);
or U19075 (N_19075,N_16697,N_15385);
or U19076 (N_19076,N_17892,N_17093);
xor U19077 (N_19077,N_17043,N_15106);
and U19078 (N_19078,N_15879,N_17219);
nand U19079 (N_19079,N_16353,N_16299);
and U19080 (N_19080,N_15241,N_16969);
or U19081 (N_19081,N_16546,N_15851);
xnor U19082 (N_19082,N_15281,N_17104);
xnor U19083 (N_19083,N_16169,N_16924);
and U19084 (N_19084,N_16784,N_15669);
or U19085 (N_19085,N_17176,N_16623);
and U19086 (N_19086,N_17261,N_17462);
and U19087 (N_19087,N_16874,N_15991);
nand U19088 (N_19088,N_15228,N_15330);
or U19089 (N_19089,N_17400,N_17444);
nor U19090 (N_19090,N_15415,N_17767);
or U19091 (N_19091,N_15027,N_16761);
xor U19092 (N_19092,N_15568,N_16682);
and U19093 (N_19093,N_15046,N_16716);
or U19094 (N_19094,N_17676,N_17449);
or U19095 (N_19095,N_17738,N_17575);
xor U19096 (N_19096,N_16833,N_17364);
nand U19097 (N_19097,N_16451,N_15662);
xnor U19098 (N_19098,N_15751,N_17006);
and U19099 (N_19099,N_16885,N_16691);
nor U19100 (N_19100,N_17408,N_17389);
and U19101 (N_19101,N_16415,N_16137);
or U19102 (N_19102,N_15661,N_17200);
xnor U19103 (N_19103,N_15036,N_15390);
nand U19104 (N_19104,N_17699,N_16188);
or U19105 (N_19105,N_16078,N_16488);
nand U19106 (N_19106,N_15924,N_16134);
nand U19107 (N_19107,N_16626,N_17829);
nand U19108 (N_19108,N_15334,N_15558);
and U19109 (N_19109,N_17646,N_16066);
nor U19110 (N_19110,N_16333,N_17805);
and U19111 (N_19111,N_16229,N_17580);
or U19112 (N_19112,N_15838,N_17846);
xnor U19113 (N_19113,N_17955,N_17127);
and U19114 (N_19114,N_17381,N_16990);
or U19115 (N_19115,N_15881,N_16099);
xnor U19116 (N_19116,N_15431,N_15671);
xnor U19117 (N_19117,N_16877,N_16656);
xnor U19118 (N_19118,N_15975,N_17865);
xor U19119 (N_19119,N_15477,N_17036);
or U19120 (N_19120,N_15154,N_17375);
and U19121 (N_19121,N_15404,N_16085);
xor U19122 (N_19122,N_15308,N_17915);
nor U19123 (N_19123,N_15230,N_17374);
or U19124 (N_19124,N_17078,N_15369);
and U19125 (N_19125,N_17764,N_17548);
nor U19126 (N_19126,N_16680,N_15525);
nor U19127 (N_19127,N_15895,N_15367);
xor U19128 (N_19128,N_15412,N_16586);
nor U19129 (N_19129,N_16639,N_16274);
xor U19130 (N_19130,N_17382,N_16595);
nor U19131 (N_19131,N_16288,N_17235);
nor U19132 (N_19132,N_15380,N_17478);
or U19133 (N_19133,N_16324,N_15799);
or U19134 (N_19134,N_15848,N_16481);
nor U19135 (N_19135,N_15971,N_17702);
or U19136 (N_19136,N_16151,N_16759);
or U19137 (N_19137,N_16180,N_15481);
or U19138 (N_19138,N_17925,N_15691);
nor U19139 (N_19139,N_15940,N_16948);
or U19140 (N_19140,N_17193,N_16976);
and U19141 (N_19141,N_17792,N_16438);
nand U19142 (N_19142,N_17097,N_15925);
or U19143 (N_19143,N_15452,N_16686);
nand U19144 (N_19144,N_17514,N_17672);
and U19145 (N_19145,N_16059,N_16037);
nor U19146 (N_19146,N_16416,N_17232);
or U19147 (N_19147,N_16031,N_15987);
and U19148 (N_19148,N_15509,N_16186);
nand U19149 (N_19149,N_15786,N_16019);
nand U19150 (N_19150,N_15484,N_17530);
and U19151 (N_19151,N_16494,N_15184);
nor U19152 (N_19152,N_16096,N_17347);
nand U19153 (N_19153,N_17161,N_16223);
xnor U19154 (N_19154,N_17994,N_17020);
nor U19155 (N_19155,N_16758,N_15875);
nor U19156 (N_19156,N_15133,N_16263);
nand U19157 (N_19157,N_17118,N_15314);
and U19158 (N_19158,N_15861,N_16281);
nand U19159 (N_19159,N_16790,N_16518);
or U19160 (N_19160,N_15563,N_15733);
xnor U19161 (N_19161,N_17499,N_17711);
or U19162 (N_19162,N_16501,N_15557);
or U19163 (N_19163,N_16376,N_17963);
nand U19164 (N_19164,N_15577,N_15062);
nor U19165 (N_19165,N_15122,N_17467);
or U19166 (N_19166,N_17567,N_16450);
and U19167 (N_19167,N_15585,N_16347);
nor U19168 (N_19168,N_16753,N_16425);
nand U19169 (N_19169,N_16187,N_15060);
nand U19170 (N_19170,N_15834,N_15617);
or U19171 (N_19171,N_15857,N_15858);
nand U19172 (N_19172,N_17811,N_15623);
xnor U19173 (N_19173,N_17203,N_15717);
and U19174 (N_19174,N_16345,N_15445);
and U19175 (N_19175,N_17536,N_17269);
and U19176 (N_19176,N_15565,N_15535);
nor U19177 (N_19177,N_15654,N_16572);
xor U19178 (N_19178,N_15290,N_15518);
nand U19179 (N_19179,N_17791,N_15328);
xnor U19180 (N_19180,N_17645,N_16890);
and U19181 (N_19181,N_15684,N_16606);
xnor U19182 (N_19182,N_16062,N_17273);
and U19183 (N_19183,N_17075,N_15204);
and U19184 (N_19184,N_15782,N_16388);
xnor U19185 (N_19185,N_17466,N_17170);
nand U19186 (N_19186,N_17010,N_16762);
nor U19187 (N_19187,N_17059,N_16266);
and U19188 (N_19188,N_16994,N_15309);
or U19189 (N_19189,N_15772,N_15939);
xnor U19190 (N_19190,N_16090,N_15873);
and U19191 (N_19191,N_17670,N_17733);
nand U19192 (N_19192,N_17797,N_16030);
nand U19193 (N_19193,N_17230,N_15457);
and U19194 (N_19194,N_15406,N_15250);
or U19195 (N_19195,N_17578,N_15666);
or U19196 (N_19196,N_17113,N_15552);
nand U19197 (N_19197,N_16455,N_16754);
xor U19198 (N_19198,N_16477,N_17077);
nor U19199 (N_19199,N_17290,N_15374);
xnor U19200 (N_19200,N_15353,N_16248);
and U19201 (N_19201,N_15124,N_17069);
and U19202 (N_19202,N_15823,N_15069);
and U19203 (N_19203,N_15533,N_15744);
xor U19204 (N_19204,N_17425,N_17030);
nand U19205 (N_19205,N_17825,N_15718);
nor U19206 (N_19206,N_16516,N_16138);
xor U19207 (N_19207,N_16673,N_16195);
and U19208 (N_19208,N_16643,N_16900);
or U19209 (N_19209,N_15832,N_16534);
or U19210 (N_19210,N_17072,N_16086);
nor U19211 (N_19211,N_17981,N_16071);
or U19212 (N_19212,N_15490,N_15821);
nor U19213 (N_19213,N_17154,N_16241);
or U19214 (N_19214,N_15377,N_17461);
nor U19215 (N_19215,N_16959,N_16520);
and U19216 (N_19216,N_17317,N_17604);
nor U19217 (N_19217,N_15601,N_15593);
or U19218 (N_19218,N_15562,N_16718);
and U19219 (N_19219,N_16371,N_15645);
xnor U19220 (N_19220,N_17905,N_16702);
xor U19221 (N_19221,N_17092,N_15264);
or U19222 (N_19222,N_15968,N_15311);
nand U19223 (N_19223,N_15877,N_17869);
or U19224 (N_19224,N_15350,N_15135);
xnor U19225 (N_19225,N_16039,N_16471);
or U19226 (N_19226,N_17614,N_17799);
and U19227 (N_19227,N_17210,N_15854);
xnor U19228 (N_19228,N_16470,N_16243);
or U19229 (N_19229,N_17299,N_17824);
nor U19230 (N_19230,N_16279,N_17017);
and U19231 (N_19231,N_17838,N_15801);
xnor U19232 (N_19232,N_17089,N_17025);
nand U19233 (N_19233,N_17379,N_17840);
xor U19234 (N_19234,N_17021,N_17945);
and U19235 (N_19235,N_15472,N_17820);
or U19236 (N_19236,N_17588,N_15305);
xnor U19237 (N_19237,N_15780,N_15322);
nand U19238 (N_19238,N_15394,N_15912);
nand U19239 (N_19239,N_15859,N_15103);
nor U19240 (N_19240,N_16828,N_15647);
nand U19241 (N_19241,N_17051,N_15271);
and U19242 (N_19242,N_17842,N_15809);
xnor U19243 (N_19243,N_17832,N_16363);
xnor U19244 (N_19244,N_16489,N_16447);
nor U19245 (N_19245,N_15749,N_17605);
or U19246 (N_19246,N_16356,N_16568);
or U19247 (N_19247,N_17106,N_15111);
and U19248 (N_19248,N_17101,N_15964);
xor U19249 (N_19249,N_15213,N_16600);
or U19250 (N_19250,N_16185,N_15688);
nor U19251 (N_19251,N_17073,N_15792);
xnor U19252 (N_19252,N_15590,N_15608);
and U19253 (N_19253,N_16628,N_15037);
nand U19254 (N_19254,N_17446,N_15239);
nand U19255 (N_19255,N_17356,N_17052);
nand U19256 (N_19256,N_16622,N_17111);
nand U19257 (N_19257,N_15600,N_17587);
and U19258 (N_19258,N_17856,N_16591);
or U19259 (N_19259,N_15170,N_16065);
or U19260 (N_19260,N_15141,N_15730);
nand U19261 (N_19261,N_16028,N_16743);
xnor U19262 (N_19262,N_15962,N_17217);
nand U19263 (N_19263,N_15884,N_15735);
or U19264 (N_19264,N_16088,N_15835);
and U19265 (N_19265,N_16585,N_15896);
xor U19266 (N_19266,N_15038,N_16846);
nor U19267 (N_19267,N_16801,N_15053);
and U19268 (N_19268,N_15607,N_15942);
and U19269 (N_19269,N_15339,N_16328);
or U19270 (N_19270,N_15464,N_16633);
nand U19271 (N_19271,N_15542,N_17150);
xnor U19272 (N_19272,N_17595,N_15199);
nor U19273 (N_19273,N_17272,N_17091);
nor U19274 (N_19274,N_16710,N_16984);
nand U19275 (N_19275,N_15716,N_15836);
or U19276 (N_19276,N_15325,N_17241);
nand U19277 (N_19277,N_16507,N_17274);
or U19278 (N_19278,N_15741,N_15534);
and U19279 (N_19279,N_17727,N_16873);
xnor U19280 (N_19280,N_16763,N_17311);
and U19281 (N_19281,N_15731,N_16026);
nor U19282 (N_19282,N_15685,N_15719);
or U19283 (N_19283,N_17653,N_17845);
nor U19284 (N_19284,N_15833,N_16426);
and U19285 (N_19285,N_16350,N_15129);
nor U19286 (N_19286,N_17518,N_15094);
xor U19287 (N_19287,N_17265,N_15474);
nand U19288 (N_19288,N_15297,N_16712);
xnor U19289 (N_19289,N_17839,N_15888);
and U19290 (N_19290,N_17948,N_15116);
and U19291 (N_19291,N_16149,N_16724);
nor U19292 (N_19292,N_17007,N_16226);
or U19293 (N_19293,N_16189,N_15516);
xnor U19294 (N_19294,N_16778,N_16922);
or U19295 (N_19295,N_16155,N_15121);
xnor U19296 (N_19296,N_16964,N_16962);
xor U19297 (N_19297,N_15810,N_15007);
and U19298 (N_19298,N_17581,N_17652);
or U19299 (N_19299,N_16530,N_16075);
nand U19300 (N_19300,N_17814,N_16747);
nor U19301 (N_19301,N_15659,N_16921);
nand U19302 (N_19302,N_17520,N_16326);
xnor U19303 (N_19303,N_15387,N_17965);
xnor U19304 (N_19304,N_17392,N_15537);
nor U19305 (N_19305,N_16597,N_16652);
xnor U19306 (N_19306,N_17654,N_17362);
or U19307 (N_19307,N_17872,N_17664);
nor U19308 (N_19308,N_16973,N_15351);
or U19309 (N_19309,N_17300,N_15347);
and U19310 (N_19310,N_16936,N_17871);
nor U19311 (N_19311,N_17993,N_17358);
xor U19312 (N_19312,N_16485,N_16473);
xor U19313 (N_19313,N_17390,N_16711);
and U19314 (N_19314,N_15012,N_15205);
xnor U19315 (N_19315,N_16100,N_17747);
and U19316 (N_19316,N_17523,N_17041);
or U19317 (N_19317,N_15620,N_16178);
nor U19318 (N_19318,N_15292,N_15830);
nand U19319 (N_19319,N_15627,N_17988);
or U19320 (N_19320,N_15418,N_17816);
or U19321 (N_19321,N_16209,N_15217);
xnor U19322 (N_19322,N_17496,N_16519);
nand U19323 (N_19323,N_17722,N_17440);
or U19324 (N_19324,N_17504,N_17982);
and U19325 (N_19325,N_17626,N_17644);
nand U19326 (N_19326,N_16589,N_17122);
and U19327 (N_19327,N_15419,N_17753);
nor U19328 (N_19328,N_15089,N_17999);
and U19329 (N_19329,N_16374,N_15926);
or U19330 (N_19330,N_16937,N_16699);
xor U19331 (N_19331,N_15546,N_17324);
or U19332 (N_19332,N_15000,N_16692);
xnor U19333 (N_19333,N_17966,N_17855);
nand U19334 (N_19334,N_15202,N_16739);
and U19335 (N_19335,N_15024,N_16117);
nand U19336 (N_19336,N_16933,N_17649);
nand U19337 (N_19337,N_15903,N_17950);
nand U19338 (N_19338,N_17042,N_17613);
and U19339 (N_19339,N_17663,N_16344);
or U19340 (N_19340,N_17977,N_17067);
nor U19341 (N_19341,N_15421,N_15919);
or U19342 (N_19342,N_17517,N_17941);
xnor U19343 (N_19343,N_17574,N_15279);
nand U19344 (N_19344,N_15844,N_15752);
nor U19345 (N_19345,N_17583,N_17320);
or U19346 (N_19346,N_17545,N_17619);
and U19347 (N_19347,N_17259,N_15583);
nand U19348 (N_19348,N_16810,N_15966);
nand U19349 (N_19349,N_17923,N_17775);
nor U19350 (N_19350,N_15382,N_15967);
and U19351 (N_19351,N_16022,N_16505);
nand U19352 (N_19352,N_15393,N_17639);
nand U19353 (N_19353,N_17860,N_16445);
nor U19354 (N_19354,N_17656,N_16894);
and U19355 (N_19355,N_15507,N_17252);
and U19356 (N_19356,N_16942,N_17875);
or U19357 (N_19357,N_16101,N_17637);
xnor U19358 (N_19358,N_16669,N_16144);
nor U19359 (N_19359,N_17951,N_15886);
nand U19360 (N_19360,N_15695,N_17555);
nand U19361 (N_19361,N_17909,N_16904);
or U19362 (N_19362,N_15030,N_17835);
xor U19363 (N_19363,N_17841,N_17719);
and U19364 (N_19364,N_15839,N_17196);
nor U19365 (N_19365,N_15655,N_17904);
xor U19366 (N_19366,N_17003,N_16183);
nand U19367 (N_19367,N_15725,N_17786);
nand U19368 (N_19368,N_17516,N_17746);
xnor U19369 (N_19369,N_15791,N_17750);
xor U19370 (N_19370,N_16409,N_15076);
nor U19371 (N_19371,N_17064,N_17159);
nor U19372 (N_19372,N_15750,N_15777);
xor U19373 (N_19373,N_17214,N_17155);
xor U19374 (N_19374,N_17231,N_17596);
nor U19375 (N_19375,N_15806,N_15764);
nor U19376 (N_19376,N_16991,N_15680);
or U19377 (N_19377,N_16104,N_17757);
and U19378 (N_19378,N_16911,N_17821);
and U19379 (N_19379,N_17401,N_16381);
or U19380 (N_19380,N_17391,N_15981);
nand U19381 (N_19381,N_17352,N_17500);
xor U19382 (N_19382,N_17543,N_17907);
nor U19383 (N_19383,N_16203,N_15914);
or U19384 (N_19384,N_15656,N_16087);
or U19385 (N_19385,N_16322,N_16588);
nor U19386 (N_19386,N_15763,N_17372);
or U19387 (N_19387,N_17695,N_15063);
and U19388 (N_19388,N_15166,N_16490);
xor U19389 (N_19389,N_15143,N_15340);
nor U19390 (N_19390,N_16231,N_15500);
nor U19391 (N_19391,N_15889,N_17201);
xnor U19392 (N_19392,N_17693,N_17438);
nand U19393 (N_19393,N_16542,N_17714);
nand U19394 (N_19394,N_16435,N_16015);
or U19395 (N_19395,N_17638,N_16919);
xnor U19396 (N_19396,N_16089,N_17163);
nand U19397 (N_19397,N_16854,N_17519);
or U19398 (N_19398,N_16514,N_17946);
nor U19399 (N_19399,N_16400,N_16446);
xnor U19400 (N_19400,N_17716,N_15869);
xnor U19401 (N_19401,N_15954,N_16027);
and U19402 (N_19402,N_17684,N_16579);
or U19403 (N_19403,N_17526,N_16254);
nand U19404 (N_19404,N_15306,N_15905);
and U19405 (N_19405,N_17610,N_17034);
nand U19406 (N_19406,N_16687,N_16889);
or U19407 (N_19407,N_17568,N_16362);
xor U19408 (N_19408,N_15892,N_17195);
nor U19409 (N_19409,N_15961,N_15023);
xnor U19410 (N_19410,N_15181,N_15218);
nand U19411 (N_19411,N_15789,N_17160);
and U19412 (N_19412,N_16058,N_15665);
or U19413 (N_19413,N_16210,N_16148);
xor U19414 (N_19414,N_17112,N_16174);
or U19415 (N_19415,N_16653,N_17686);
nand U19416 (N_19416,N_16674,N_16917);
xnor U19417 (N_19417,N_16531,N_17634);
or U19418 (N_19418,N_17937,N_16864);
and U19419 (N_19419,N_17544,N_15345);
nand U19420 (N_19420,N_16608,N_17107);
and U19421 (N_19421,N_17482,N_16614);
xor U19422 (N_19422,N_15316,N_16822);
xor U19423 (N_19423,N_15606,N_16238);
or U19424 (N_19424,N_17124,N_16460);
xnor U19425 (N_19425,N_17700,N_15517);
xor U19426 (N_19426,N_17660,N_15853);
and U19427 (N_19427,N_17736,N_17055);
or U19428 (N_19428,N_15134,N_15697);
and U19429 (N_19429,N_15259,N_17801);
xor U19430 (N_19430,N_16351,N_17470);
nor U19431 (N_19431,N_16040,N_17156);
xnor U19432 (N_19432,N_15901,N_15072);
nor U19433 (N_19433,N_15992,N_16428);
nor U19434 (N_19434,N_16655,N_15970);
or U19435 (N_19435,N_17140,N_15392);
or U19436 (N_19436,N_15329,N_17980);
xnor U19437 (N_19437,N_17940,N_16509);
and U19438 (N_19438,N_15147,N_17468);
nand U19439 (N_19439,N_15191,N_16525);
nand U19440 (N_19440,N_15596,N_15494);
nor U19441 (N_19441,N_16721,N_16202);
nand U19442 (N_19442,N_16830,N_17983);
and U19443 (N_19443,N_15773,N_16684);
and U19444 (N_19444,N_15155,N_16571);
and U19445 (N_19445,N_16923,N_15238);
nor U19446 (N_19446,N_15384,N_15843);
xor U19447 (N_19447,N_16744,N_16378);
and U19448 (N_19448,N_16124,N_16926);
xor U19449 (N_19449,N_16544,N_16719);
or U19450 (N_19450,N_15813,N_16574);
and U19451 (N_19451,N_17789,N_16370);
nand U19452 (N_19452,N_15341,N_17896);
xnor U19453 (N_19453,N_15937,N_16715);
nand U19454 (N_19454,N_16373,N_16788);
or U19455 (N_19455,N_17675,N_17322);
xor U19456 (N_19456,N_16084,N_15635);
xor U19457 (N_19457,N_15315,N_17717);
nor U19458 (N_19458,N_15453,N_17765);
or U19459 (N_19459,N_15638,N_16130);
nor U19460 (N_19460,N_17622,N_16651);
nand U19461 (N_19461,N_15540,N_17920);
nand U19462 (N_19462,N_16528,N_16204);
or U19463 (N_19463,N_17742,N_16276);
nand U19464 (N_19464,N_15734,N_17354);
xor U19465 (N_19465,N_16524,N_15395);
nand U19466 (N_19466,N_15765,N_17859);
and U19467 (N_19467,N_16265,N_15613);
nor U19468 (N_19468,N_16465,N_16128);
nor U19469 (N_19469,N_17833,N_16357);
nor U19470 (N_19470,N_15168,N_16781);
nand U19471 (N_19471,N_15711,N_17332);
xor U19472 (N_19472,N_17912,N_15100);
nand U19473 (N_19473,N_17009,N_15820);
xor U19474 (N_19474,N_16257,N_16785);
nor U19475 (N_19475,N_16929,N_17463);
nand U19476 (N_19476,N_16621,N_17304);
xor U19477 (N_19477,N_17706,N_15131);
nor U19478 (N_19478,N_16383,N_17233);
nand U19479 (N_19479,N_16182,N_15360);
xor U19480 (N_19480,N_17386,N_17397);
and U19481 (N_19481,N_16541,N_15625);
nand U19482 (N_19482,N_17490,N_15640);
nor U19483 (N_19483,N_16612,N_15598);
nor U19484 (N_19484,N_15026,N_15287);
nand U19485 (N_19485,N_17054,N_16966);
and U19486 (N_19486,N_17513,N_16369);
nand U19487 (N_19487,N_17823,N_16068);
or U19488 (N_19488,N_16826,N_16634);
and U19489 (N_19489,N_15273,N_17207);
nand U19490 (N_19490,N_17023,N_15363);
xor U19491 (N_19491,N_15113,N_17147);
and U19492 (N_19492,N_16457,N_17562);
nand U19493 (N_19493,N_15207,N_15783);
or U19494 (N_19494,N_17435,N_17673);
nand U19495 (N_19495,N_15318,N_17130);
and U19496 (N_19496,N_16304,N_15376);
xnor U19497 (N_19497,N_16735,N_17270);
and U19498 (N_19498,N_15631,N_17592);
or U19499 (N_19499,N_16870,N_16664);
xnor U19500 (N_19500,N_16800,N_15658);
and U19501 (N_19501,N_16307,N_17647);
xnor U19502 (N_19502,N_17667,N_16965);
nor U19503 (N_19503,N_15617,N_15796);
or U19504 (N_19504,N_16515,N_17754);
and U19505 (N_19505,N_17528,N_16752);
or U19506 (N_19506,N_16691,N_16500);
nand U19507 (N_19507,N_15206,N_17453);
xor U19508 (N_19508,N_15202,N_15083);
nand U19509 (N_19509,N_16988,N_15550);
nand U19510 (N_19510,N_15567,N_17263);
xnor U19511 (N_19511,N_15495,N_17242);
nor U19512 (N_19512,N_16666,N_16378);
nor U19513 (N_19513,N_15771,N_16716);
and U19514 (N_19514,N_15014,N_16870);
or U19515 (N_19515,N_17087,N_16601);
and U19516 (N_19516,N_16940,N_16021);
or U19517 (N_19517,N_17727,N_17346);
nor U19518 (N_19518,N_16818,N_17783);
nor U19519 (N_19519,N_16285,N_15221);
xor U19520 (N_19520,N_15296,N_17353);
nor U19521 (N_19521,N_16501,N_17446);
or U19522 (N_19522,N_15750,N_16325);
nand U19523 (N_19523,N_15396,N_16397);
xor U19524 (N_19524,N_15666,N_15659);
xnor U19525 (N_19525,N_15932,N_16716);
or U19526 (N_19526,N_17333,N_16461);
nor U19527 (N_19527,N_15230,N_16014);
nor U19528 (N_19528,N_17261,N_17339);
nand U19529 (N_19529,N_16899,N_16517);
and U19530 (N_19530,N_15819,N_16761);
nand U19531 (N_19531,N_16875,N_15852);
or U19532 (N_19532,N_17457,N_17068);
nand U19533 (N_19533,N_16335,N_15679);
nor U19534 (N_19534,N_15871,N_15201);
nand U19535 (N_19535,N_17879,N_15381);
and U19536 (N_19536,N_16537,N_15931);
nor U19537 (N_19537,N_17199,N_17027);
and U19538 (N_19538,N_17575,N_16843);
xnor U19539 (N_19539,N_15264,N_15377);
or U19540 (N_19540,N_17276,N_15099);
xnor U19541 (N_19541,N_15407,N_15435);
nand U19542 (N_19542,N_17139,N_16259);
or U19543 (N_19543,N_16297,N_16461);
nand U19544 (N_19544,N_15165,N_17742);
nor U19545 (N_19545,N_15254,N_16740);
nor U19546 (N_19546,N_15594,N_17599);
or U19547 (N_19547,N_16146,N_15715);
and U19548 (N_19548,N_15604,N_15485);
or U19549 (N_19549,N_15072,N_15991);
and U19550 (N_19550,N_15094,N_17178);
nor U19551 (N_19551,N_17654,N_16389);
nand U19552 (N_19552,N_17823,N_15575);
and U19553 (N_19553,N_15801,N_16014);
nand U19554 (N_19554,N_17379,N_16976);
xor U19555 (N_19555,N_16602,N_15820);
or U19556 (N_19556,N_16265,N_17703);
and U19557 (N_19557,N_16795,N_17512);
nand U19558 (N_19558,N_15983,N_17590);
xor U19559 (N_19559,N_15964,N_16785);
xor U19560 (N_19560,N_16049,N_17455);
and U19561 (N_19561,N_16961,N_16035);
or U19562 (N_19562,N_15059,N_17043);
nor U19563 (N_19563,N_16218,N_17587);
xnor U19564 (N_19564,N_17032,N_15354);
nor U19565 (N_19565,N_16893,N_17909);
xor U19566 (N_19566,N_15169,N_17121);
and U19567 (N_19567,N_15538,N_16544);
nand U19568 (N_19568,N_15634,N_15840);
nand U19569 (N_19569,N_15700,N_16181);
xnor U19570 (N_19570,N_16105,N_15620);
and U19571 (N_19571,N_17140,N_17204);
xnor U19572 (N_19572,N_17139,N_15120);
and U19573 (N_19573,N_17172,N_16277);
nand U19574 (N_19574,N_17677,N_16764);
and U19575 (N_19575,N_16199,N_15735);
xor U19576 (N_19576,N_15680,N_16130);
or U19577 (N_19577,N_15970,N_16048);
xor U19578 (N_19578,N_15114,N_16822);
or U19579 (N_19579,N_16769,N_16549);
nand U19580 (N_19580,N_16470,N_17068);
nor U19581 (N_19581,N_15850,N_17502);
nor U19582 (N_19582,N_17701,N_15417);
nand U19583 (N_19583,N_16015,N_16299);
nor U19584 (N_19584,N_17197,N_16423);
xnor U19585 (N_19585,N_15087,N_15997);
nand U19586 (N_19586,N_16191,N_15558);
nor U19587 (N_19587,N_17500,N_15586);
or U19588 (N_19588,N_17947,N_15742);
xor U19589 (N_19589,N_16979,N_16879);
and U19590 (N_19590,N_16308,N_15641);
or U19591 (N_19591,N_15900,N_16187);
and U19592 (N_19592,N_17156,N_15784);
or U19593 (N_19593,N_16236,N_16845);
nor U19594 (N_19594,N_16176,N_15353);
xor U19595 (N_19595,N_16740,N_15938);
nand U19596 (N_19596,N_15053,N_17229);
nand U19597 (N_19597,N_17894,N_16007);
nor U19598 (N_19598,N_16122,N_15520);
nand U19599 (N_19599,N_16042,N_17208);
xnor U19600 (N_19600,N_15451,N_17426);
or U19601 (N_19601,N_15583,N_15563);
nand U19602 (N_19602,N_16541,N_15355);
xor U19603 (N_19603,N_16065,N_17599);
and U19604 (N_19604,N_17517,N_17903);
or U19605 (N_19605,N_16467,N_16533);
or U19606 (N_19606,N_15079,N_16282);
or U19607 (N_19607,N_17424,N_16042);
nand U19608 (N_19608,N_15384,N_15794);
nand U19609 (N_19609,N_15692,N_15026);
xnor U19610 (N_19610,N_17716,N_15976);
or U19611 (N_19611,N_15626,N_15550);
xnor U19612 (N_19612,N_15005,N_16013);
nand U19613 (N_19613,N_16689,N_16073);
nand U19614 (N_19614,N_16895,N_16049);
or U19615 (N_19615,N_15578,N_17408);
xnor U19616 (N_19616,N_17954,N_15886);
nand U19617 (N_19617,N_16851,N_16649);
and U19618 (N_19618,N_17217,N_17179);
nand U19619 (N_19619,N_17635,N_16652);
nor U19620 (N_19620,N_15991,N_16464);
nand U19621 (N_19621,N_16606,N_15116);
nor U19622 (N_19622,N_16548,N_15242);
or U19623 (N_19623,N_17068,N_15250);
or U19624 (N_19624,N_15005,N_16289);
xnor U19625 (N_19625,N_17592,N_16862);
nor U19626 (N_19626,N_17274,N_15286);
nor U19627 (N_19627,N_15617,N_15613);
xnor U19628 (N_19628,N_17958,N_15754);
or U19629 (N_19629,N_17176,N_17564);
nor U19630 (N_19630,N_15484,N_15953);
and U19631 (N_19631,N_16159,N_15119);
nand U19632 (N_19632,N_16420,N_17884);
xnor U19633 (N_19633,N_15612,N_16727);
or U19634 (N_19634,N_17060,N_16779);
or U19635 (N_19635,N_17558,N_17731);
nand U19636 (N_19636,N_16393,N_17956);
nor U19637 (N_19637,N_16269,N_16512);
or U19638 (N_19638,N_16028,N_16475);
and U19639 (N_19639,N_15653,N_17178);
nand U19640 (N_19640,N_15103,N_16879);
and U19641 (N_19641,N_16400,N_17568);
or U19642 (N_19642,N_16361,N_15372);
nand U19643 (N_19643,N_15257,N_16453);
and U19644 (N_19644,N_17408,N_15830);
nand U19645 (N_19645,N_16229,N_17528);
and U19646 (N_19646,N_17258,N_17168);
and U19647 (N_19647,N_16392,N_16041);
nand U19648 (N_19648,N_16318,N_16777);
nand U19649 (N_19649,N_17241,N_16775);
nor U19650 (N_19650,N_16199,N_17226);
nand U19651 (N_19651,N_17650,N_15038);
and U19652 (N_19652,N_17920,N_17552);
and U19653 (N_19653,N_17952,N_15727);
nand U19654 (N_19654,N_16888,N_15987);
or U19655 (N_19655,N_16390,N_17979);
and U19656 (N_19656,N_16198,N_17213);
xor U19657 (N_19657,N_15837,N_15955);
nor U19658 (N_19658,N_17922,N_17730);
nand U19659 (N_19659,N_16346,N_15706);
or U19660 (N_19660,N_17924,N_15252);
nand U19661 (N_19661,N_16382,N_16134);
or U19662 (N_19662,N_17327,N_17423);
nor U19663 (N_19663,N_15010,N_16304);
nand U19664 (N_19664,N_17289,N_15610);
and U19665 (N_19665,N_17530,N_15986);
or U19666 (N_19666,N_17092,N_17207);
nor U19667 (N_19667,N_16547,N_16689);
xor U19668 (N_19668,N_15651,N_16369);
nand U19669 (N_19669,N_15228,N_16296);
and U19670 (N_19670,N_17901,N_16009);
xnor U19671 (N_19671,N_17633,N_17151);
nor U19672 (N_19672,N_16943,N_15564);
nor U19673 (N_19673,N_16735,N_17696);
nor U19674 (N_19674,N_15363,N_15186);
xor U19675 (N_19675,N_16910,N_16710);
or U19676 (N_19676,N_16188,N_17065);
nand U19677 (N_19677,N_15658,N_17682);
xor U19678 (N_19678,N_16461,N_15384);
nand U19679 (N_19679,N_15800,N_16936);
xor U19680 (N_19680,N_17079,N_16833);
xnor U19681 (N_19681,N_16512,N_15638);
nor U19682 (N_19682,N_15230,N_16518);
and U19683 (N_19683,N_16279,N_15743);
nand U19684 (N_19684,N_15036,N_17581);
and U19685 (N_19685,N_16906,N_15352);
xnor U19686 (N_19686,N_17500,N_16000);
or U19687 (N_19687,N_16368,N_15511);
xor U19688 (N_19688,N_15697,N_16751);
nand U19689 (N_19689,N_15946,N_15646);
and U19690 (N_19690,N_17834,N_15241);
and U19691 (N_19691,N_16627,N_17438);
nor U19692 (N_19692,N_16633,N_17210);
nor U19693 (N_19693,N_16774,N_17503);
nand U19694 (N_19694,N_17865,N_17937);
nand U19695 (N_19695,N_15476,N_15575);
nor U19696 (N_19696,N_15376,N_16635);
or U19697 (N_19697,N_17480,N_15080);
and U19698 (N_19698,N_17271,N_16607);
or U19699 (N_19699,N_16997,N_17207);
and U19700 (N_19700,N_16877,N_16054);
nand U19701 (N_19701,N_16203,N_15933);
xor U19702 (N_19702,N_17479,N_15759);
nor U19703 (N_19703,N_16641,N_15390);
xnor U19704 (N_19704,N_16823,N_16356);
or U19705 (N_19705,N_17409,N_16978);
nand U19706 (N_19706,N_17629,N_15307);
xnor U19707 (N_19707,N_16538,N_16165);
xor U19708 (N_19708,N_17180,N_15146);
xor U19709 (N_19709,N_16318,N_17991);
xnor U19710 (N_19710,N_15821,N_17511);
and U19711 (N_19711,N_17694,N_15403);
xor U19712 (N_19712,N_16976,N_17315);
nand U19713 (N_19713,N_15660,N_17646);
or U19714 (N_19714,N_15601,N_16284);
or U19715 (N_19715,N_16639,N_15887);
or U19716 (N_19716,N_16682,N_15988);
nor U19717 (N_19717,N_16486,N_17073);
and U19718 (N_19718,N_16192,N_15420);
nor U19719 (N_19719,N_16507,N_16184);
nand U19720 (N_19720,N_15549,N_15158);
or U19721 (N_19721,N_17924,N_15900);
nand U19722 (N_19722,N_16652,N_16623);
nand U19723 (N_19723,N_16934,N_17434);
nor U19724 (N_19724,N_15560,N_17266);
nand U19725 (N_19725,N_16337,N_17268);
xor U19726 (N_19726,N_17933,N_16992);
nand U19727 (N_19727,N_15894,N_15044);
or U19728 (N_19728,N_17574,N_16417);
or U19729 (N_19729,N_17107,N_16231);
or U19730 (N_19730,N_17341,N_15609);
nand U19731 (N_19731,N_16062,N_17819);
or U19732 (N_19732,N_16618,N_16253);
nand U19733 (N_19733,N_16982,N_17981);
nand U19734 (N_19734,N_16243,N_15638);
xnor U19735 (N_19735,N_15613,N_16488);
and U19736 (N_19736,N_16839,N_17438);
nor U19737 (N_19737,N_16373,N_16142);
nor U19738 (N_19738,N_17376,N_15855);
nand U19739 (N_19739,N_15955,N_16302);
xor U19740 (N_19740,N_16450,N_17041);
nand U19741 (N_19741,N_15824,N_16565);
nand U19742 (N_19742,N_15277,N_15244);
xor U19743 (N_19743,N_17095,N_17583);
nand U19744 (N_19744,N_15345,N_16525);
and U19745 (N_19745,N_15930,N_16756);
xnor U19746 (N_19746,N_15442,N_15280);
xnor U19747 (N_19747,N_16155,N_16765);
xnor U19748 (N_19748,N_16980,N_17193);
and U19749 (N_19749,N_17740,N_17100);
and U19750 (N_19750,N_17580,N_16964);
xor U19751 (N_19751,N_16283,N_17046);
nor U19752 (N_19752,N_17977,N_16315);
or U19753 (N_19753,N_16639,N_17822);
nor U19754 (N_19754,N_15243,N_16475);
and U19755 (N_19755,N_15792,N_17991);
and U19756 (N_19756,N_17803,N_17180);
or U19757 (N_19757,N_15319,N_16526);
or U19758 (N_19758,N_16317,N_16114);
nand U19759 (N_19759,N_17140,N_15169);
xnor U19760 (N_19760,N_15655,N_17255);
or U19761 (N_19761,N_15211,N_16124);
nand U19762 (N_19762,N_17393,N_16250);
xor U19763 (N_19763,N_17814,N_16503);
or U19764 (N_19764,N_15035,N_16627);
nor U19765 (N_19765,N_16953,N_17480);
nand U19766 (N_19766,N_16613,N_17314);
or U19767 (N_19767,N_15648,N_17262);
xnor U19768 (N_19768,N_15292,N_16433);
or U19769 (N_19769,N_16043,N_17641);
xor U19770 (N_19770,N_15756,N_16041);
nor U19771 (N_19771,N_15304,N_16869);
nor U19772 (N_19772,N_17741,N_17436);
and U19773 (N_19773,N_17990,N_15290);
nand U19774 (N_19774,N_16586,N_15404);
xor U19775 (N_19775,N_17887,N_16446);
or U19776 (N_19776,N_17066,N_15375);
xnor U19777 (N_19777,N_15496,N_17692);
or U19778 (N_19778,N_15466,N_17372);
nor U19779 (N_19779,N_16210,N_17904);
nor U19780 (N_19780,N_16540,N_15405);
xnor U19781 (N_19781,N_16224,N_15052);
nand U19782 (N_19782,N_15513,N_16916);
xnor U19783 (N_19783,N_17921,N_17162);
nand U19784 (N_19784,N_15030,N_17622);
nand U19785 (N_19785,N_16886,N_16526);
or U19786 (N_19786,N_15975,N_17802);
xnor U19787 (N_19787,N_16148,N_15022);
nand U19788 (N_19788,N_15368,N_17734);
nand U19789 (N_19789,N_15041,N_15821);
or U19790 (N_19790,N_15225,N_16718);
and U19791 (N_19791,N_17801,N_16703);
nor U19792 (N_19792,N_17800,N_16363);
xor U19793 (N_19793,N_15189,N_17546);
and U19794 (N_19794,N_17263,N_17789);
nor U19795 (N_19795,N_17998,N_15037);
nand U19796 (N_19796,N_17102,N_15139);
xor U19797 (N_19797,N_16837,N_17550);
nand U19798 (N_19798,N_17493,N_15409);
xor U19799 (N_19799,N_16210,N_15185);
xnor U19800 (N_19800,N_17610,N_17467);
nor U19801 (N_19801,N_17556,N_16494);
nand U19802 (N_19802,N_15259,N_17706);
nand U19803 (N_19803,N_17353,N_16558);
nor U19804 (N_19804,N_15106,N_15029);
nor U19805 (N_19805,N_17432,N_15232);
and U19806 (N_19806,N_15444,N_17369);
nand U19807 (N_19807,N_17629,N_16277);
nand U19808 (N_19808,N_15243,N_17234);
and U19809 (N_19809,N_17939,N_15939);
nand U19810 (N_19810,N_15202,N_17814);
xnor U19811 (N_19811,N_16930,N_16031);
nor U19812 (N_19812,N_17996,N_15783);
and U19813 (N_19813,N_15236,N_16693);
nand U19814 (N_19814,N_15477,N_15317);
nor U19815 (N_19815,N_16388,N_15737);
nand U19816 (N_19816,N_16426,N_15288);
or U19817 (N_19817,N_16491,N_17380);
nand U19818 (N_19818,N_17622,N_17913);
and U19819 (N_19819,N_17347,N_17716);
or U19820 (N_19820,N_15923,N_17117);
nand U19821 (N_19821,N_17302,N_17142);
and U19822 (N_19822,N_17058,N_16493);
nand U19823 (N_19823,N_17065,N_15626);
xnor U19824 (N_19824,N_15001,N_15914);
or U19825 (N_19825,N_15794,N_17318);
and U19826 (N_19826,N_15417,N_15122);
or U19827 (N_19827,N_16989,N_15739);
and U19828 (N_19828,N_16720,N_16551);
xor U19829 (N_19829,N_17827,N_16615);
and U19830 (N_19830,N_17503,N_15388);
and U19831 (N_19831,N_15350,N_17355);
and U19832 (N_19832,N_17713,N_16025);
nand U19833 (N_19833,N_17216,N_15840);
xor U19834 (N_19834,N_15854,N_17620);
nand U19835 (N_19835,N_15010,N_15240);
nand U19836 (N_19836,N_17829,N_16387);
and U19837 (N_19837,N_15934,N_15643);
xor U19838 (N_19838,N_17941,N_16782);
or U19839 (N_19839,N_16761,N_17994);
xnor U19840 (N_19840,N_15295,N_16968);
nand U19841 (N_19841,N_17306,N_15611);
or U19842 (N_19842,N_16169,N_16217);
or U19843 (N_19843,N_16386,N_15902);
or U19844 (N_19844,N_17834,N_15195);
or U19845 (N_19845,N_17303,N_17242);
nand U19846 (N_19846,N_16735,N_15102);
xor U19847 (N_19847,N_15307,N_15538);
and U19848 (N_19848,N_15101,N_17005);
and U19849 (N_19849,N_15554,N_15878);
and U19850 (N_19850,N_17075,N_17157);
nand U19851 (N_19851,N_17857,N_15726);
and U19852 (N_19852,N_17031,N_15701);
or U19853 (N_19853,N_17495,N_16005);
nor U19854 (N_19854,N_17154,N_16943);
and U19855 (N_19855,N_17418,N_15289);
nand U19856 (N_19856,N_15165,N_16114);
or U19857 (N_19857,N_15920,N_15895);
or U19858 (N_19858,N_15485,N_15891);
xnor U19859 (N_19859,N_17421,N_16835);
nor U19860 (N_19860,N_16063,N_16604);
or U19861 (N_19861,N_16429,N_17560);
nor U19862 (N_19862,N_15467,N_17563);
nor U19863 (N_19863,N_15793,N_15988);
and U19864 (N_19864,N_16955,N_16909);
nor U19865 (N_19865,N_17151,N_16689);
xnor U19866 (N_19866,N_17040,N_16497);
nor U19867 (N_19867,N_17209,N_15783);
and U19868 (N_19868,N_17347,N_17480);
nor U19869 (N_19869,N_15875,N_17631);
nor U19870 (N_19870,N_16812,N_17167);
nor U19871 (N_19871,N_17372,N_15604);
and U19872 (N_19872,N_15128,N_15637);
xnor U19873 (N_19873,N_15378,N_15321);
nand U19874 (N_19874,N_15215,N_16986);
and U19875 (N_19875,N_16120,N_16881);
and U19876 (N_19876,N_17864,N_16004);
xnor U19877 (N_19877,N_15973,N_17110);
and U19878 (N_19878,N_17305,N_17383);
and U19879 (N_19879,N_16523,N_16747);
and U19880 (N_19880,N_15893,N_16000);
nand U19881 (N_19881,N_15022,N_15156);
and U19882 (N_19882,N_16071,N_15664);
nand U19883 (N_19883,N_16531,N_15184);
xor U19884 (N_19884,N_16550,N_16729);
and U19885 (N_19885,N_15968,N_17967);
and U19886 (N_19886,N_15678,N_16398);
or U19887 (N_19887,N_16321,N_15394);
and U19888 (N_19888,N_15585,N_16696);
and U19889 (N_19889,N_17241,N_15216);
nand U19890 (N_19890,N_17632,N_16323);
nor U19891 (N_19891,N_15848,N_17477);
nor U19892 (N_19892,N_16227,N_17933);
and U19893 (N_19893,N_17935,N_15831);
or U19894 (N_19894,N_17611,N_15189);
nor U19895 (N_19895,N_15114,N_15672);
nand U19896 (N_19896,N_16842,N_15388);
nand U19897 (N_19897,N_15849,N_17898);
nand U19898 (N_19898,N_15797,N_15204);
xor U19899 (N_19899,N_15269,N_15624);
and U19900 (N_19900,N_15205,N_15347);
or U19901 (N_19901,N_15741,N_17377);
xor U19902 (N_19902,N_16346,N_15268);
nor U19903 (N_19903,N_17557,N_17793);
nor U19904 (N_19904,N_16448,N_15167);
or U19905 (N_19905,N_16687,N_15241);
nand U19906 (N_19906,N_16238,N_16506);
nand U19907 (N_19907,N_16732,N_16774);
xnor U19908 (N_19908,N_15412,N_17261);
xor U19909 (N_19909,N_16838,N_16576);
xnor U19910 (N_19910,N_17796,N_16343);
or U19911 (N_19911,N_16088,N_17098);
nor U19912 (N_19912,N_17751,N_17585);
nor U19913 (N_19913,N_16914,N_17797);
nand U19914 (N_19914,N_15676,N_16014);
nor U19915 (N_19915,N_16943,N_15510);
xnor U19916 (N_19916,N_15522,N_16754);
xnor U19917 (N_19917,N_15216,N_16216);
and U19918 (N_19918,N_16368,N_17247);
xor U19919 (N_19919,N_15287,N_17300);
xnor U19920 (N_19920,N_15564,N_16912);
and U19921 (N_19921,N_15109,N_17768);
and U19922 (N_19922,N_15020,N_16387);
and U19923 (N_19923,N_16771,N_15626);
or U19924 (N_19924,N_16153,N_16687);
or U19925 (N_19925,N_16708,N_17783);
nand U19926 (N_19926,N_17928,N_15681);
nand U19927 (N_19927,N_16303,N_17688);
nand U19928 (N_19928,N_16607,N_15896);
nor U19929 (N_19929,N_15159,N_17042);
xor U19930 (N_19930,N_17899,N_17495);
xor U19931 (N_19931,N_16870,N_17184);
nor U19932 (N_19932,N_17742,N_16663);
nor U19933 (N_19933,N_17365,N_16375);
and U19934 (N_19934,N_15564,N_16783);
and U19935 (N_19935,N_17229,N_17803);
and U19936 (N_19936,N_17982,N_17790);
nor U19937 (N_19937,N_15085,N_15446);
xnor U19938 (N_19938,N_16363,N_15074);
nand U19939 (N_19939,N_17147,N_17527);
nand U19940 (N_19940,N_17531,N_16588);
xnor U19941 (N_19941,N_16981,N_17402);
and U19942 (N_19942,N_16657,N_17110);
or U19943 (N_19943,N_17692,N_16524);
nand U19944 (N_19944,N_15334,N_16638);
nor U19945 (N_19945,N_15160,N_16537);
or U19946 (N_19946,N_17859,N_17763);
nand U19947 (N_19947,N_15897,N_15164);
xnor U19948 (N_19948,N_15922,N_16483);
or U19949 (N_19949,N_15301,N_17523);
nor U19950 (N_19950,N_16033,N_16342);
nand U19951 (N_19951,N_17740,N_16724);
or U19952 (N_19952,N_16749,N_15176);
nand U19953 (N_19953,N_16468,N_15556);
nand U19954 (N_19954,N_16050,N_16085);
nor U19955 (N_19955,N_17710,N_15443);
and U19956 (N_19956,N_16817,N_17318);
nand U19957 (N_19957,N_16500,N_15246);
or U19958 (N_19958,N_17264,N_17152);
and U19959 (N_19959,N_15970,N_17076);
or U19960 (N_19960,N_16412,N_16287);
or U19961 (N_19961,N_15422,N_16186);
and U19962 (N_19962,N_15018,N_15900);
and U19963 (N_19963,N_15814,N_16996);
and U19964 (N_19964,N_17531,N_17431);
or U19965 (N_19965,N_15082,N_17755);
and U19966 (N_19966,N_15197,N_17352);
nor U19967 (N_19967,N_17057,N_16193);
nor U19968 (N_19968,N_15189,N_15272);
nand U19969 (N_19969,N_15882,N_16850);
or U19970 (N_19970,N_15191,N_17929);
nand U19971 (N_19971,N_15672,N_16134);
nor U19972 (N_19972,N_17973,N_17981);
or U19973 (N_19973,N_17478,N_17784);
or U19974 (N_19974,N_17427,N_15878);
nor U19975 (N_19975,N_15464,N_15454);
xnor U19976 (N_19976,N_17833,N_15695);
nor U19977 (N_19977,N_16413,N_16361);
or U19978 (N_19978,N_17654,N_17005);
nand U19979 (N_19979,N_15822,N_17106);
xnor U19980 (N_19980,N_16939,N_17498);
xnor U19981 (N_19981,N_15871,N_15889);
nor U19982 (N_19982,N_16964,N_15012);
xor U19983 (N_19983,N_17942,N_17496);
xnor U19984 (N_19984,N_15769,N_17945);
nand U19985 (N_19985,N_15813,N_16724);
and U19986 (N_19986,N_15923,N_16713);
xor U19987 (N_19987,N_16359,N_16587);
or U19988 (N_19988,N_15989,N_15898);
and U19989 (N_19989,N_16812,N_15527);
and U19990 (N_19990,N_15370,N_17334);
nor U19991 (N_19991,N_16028,N_17850);
or U19992 (N_19992,N_16370,N_17208);
nor U19993 (N_19993,N_17429,N_17782);
xor U19994 (N_19994,N_16851,N_15205);
nor U19995 (N_19995,N_17879,N_17356);
and U19996 (N_19996,N_16529,N_17765);
nor U19997 (N_19997,N_16813,N_15389);
and U19998 (N_19998,N_17082,N_17818);
nand U19999 (N_19999,N_16318,N_17018);
nand U20000 (N_20000,N_17844,N_17978);
xnor U20001 (N_20001,N_15211,N_16935);
xnor U20002 (N_20002,N_16327,N_15682);
nand U20003 (N_20003,N_17376,N_17273);
nand U20004 (N_20004,N_17906,N_15675);
nand U20005 (N_20005,N_17244,N_17657);
or U20006 (N_20006,N_17181,N_15532);
nor U20007 (N_20007,N_16571,N_16469);
nor U20008 (N_20008,N_16945,N_17177);
nand U20009 (N_20009,N_15103,N_17132);
xnor U20010 (N_20010,N_15363,N_15147);
and U20011 (N_20011,N_17606,N_15448);
nand U20012 (N_20012,N_17318,N_15062);
and U20013 (N_20013,N_15773,N_15915);
nor U20014 (N_20014,N_16807,N_16694);
or U20015 (N_20015,N_15180,N_16431);
and U20016 (N_20016,N_16585,N_15917);
and U20017 (N_20017,N_15975,N_17382);
xnor U20018 (N_20018,N_15029,N_15873);
nand U20019 (N_20019,N_15192,N_17647);
and U20020 (N_20020,N_16339,N_15291);
or U20021 (N_20021,N_17162,N_17792);
xor U20022 (N_20022,N_17646,N_15816);
nor U20023 (N_20023,N_16952,N_17871);
and U20024 (N_20024,N_17181,N_16710);
or U20025 (N_20025,N_17694,N_17192);
nor U20026 (N_20026,N_17486,N_15713);
xor U20027 (N_20027,N_15916,N_16653);
xor U20028 (N_20028,N_17615,N_15828);
or U20029 (N_20029,N_15104,N_15873);
xor U20030 (N_20030,N_17892,N_17338);
xnor U20031 (N_20031,N_15270,N_17147);
nand U20032 (N_20032,N_16918,N_15202);
or U20033 (N_20033,N_16507,N_17369);
and U20034 (N_20034,N_15280,N_15794);
or U20035 (N_20035,N_17757,N_15779);
or U20036 (N_20036,N_15008,N_17439);
and U20037 (N_20037,N_15920,N_16036);
and U20038 (N_20038,N_15829,N_16142);
or U20039 (N_20039,N_17318,N_15732);
xor U20040 (N_20040,N_15524,N_16776);
or U20041 (N_20041,N_15579,N_17612);
nand U20042 (N_20042,N_15330,N_15473);
nand U20043 (N_20043,N_15740,N_15148);
nor U20044 (N_20044,N_15837,N_16011);
nor U20045 (N_20045,N_16959,N_17260);
and U20046 (N_20046,N_16192,N_16959);
nor U20047 (N_20047,N_15872,N_16431);
nor U20048 (N_20048,N_17234,N_15840);
or U20049 (N_20049,N_17102,N_16817);
nand U20050 (N_20050,N_15333,N_17284);
xor U20051 (N_20051,N_17798,N_17777);
xnor U20052 (N_20052,N_16375,N_15509);
nor U20053 (N_20053,N_15302,N_16620);
and U20054 (N_20054,N_15738,N_16574);
xnor U20055 (N_20055,N_17859,N_16393);
nor U20056 (N_20056,N_17985,N_17692);
nor U20057 (N_20057,N_15668,N_15031);
nand U20058 (N_20058,N_15350,N_17258);
or U20059 (N_20059,N_15405,N_15736);
xor U20060 (N_20060,N_16774,N_17674);
nor U20061 (N_20061,N_16468,N_15977);
nor U20062 (N_20062,N_15807,N_16732);
xnor U20063 (N_20063,N_16603,N_17974);
nand U20064 (N_20064,N_16224,N_15249);
and U20065 (N_20065,N_15477,N_16552);
xor U20066 (N_20066,N_17792,N_15967);
nor U20067 (N_20067,N_15388,N_16437);
xor U20068 (N_20068,N_16038,N_15431);
xnor U20069 (N_20069,N_17981,N_16045);
nand U20070 (N_20070,N_17184,N_17024);
nand U20071 (N_20071,N_16963,N_16564);
xor U20072 (N_20072,N_16935,N_16729);
or U20073 (N_20073,N_16978,N_15089);
and U20074 (N_20074,N_17785,N_15880);
or U20075 (N_20075,N_16439,N_16028);
xor U20076 (N_20076,N_15031,N_15433);
or U20077 (N_20077,N_16125,N_15557);
nor U20078 (N_20078,N_16019,N_15638);
nand U20079 (N_20079,N_15142,N_15688);
and U20080 (N_20080,N_16432,N_17177);
or U20081 (N_20081,N_16914,N_16919);
xor U20082 (N_20082,N_15629,N_15415);
nor U20083 (N_20083,N_16085,N_16411);
xnor U20084 (N_20084,N_17216,N_17339);
nor U20085 (N_20085,N_15650,N_17353);
or U20086 (N_20086,N_16784,N_17254);
xor U20087 (N_20087,N_17269,N_16984);
xnor U20088 (N_20088,N_16805,N_16907);
nand U20089 (N_20089,N_16256,N_15434);
and U20090 (N_20090,N_15790,N_16965);
or U20091 (N_20091,N_15802,N_17426);
or U20092 (N_20092,N_15289,N_16793);
nor U20093 (N_20093,N_17651,N_17124);
nand U20094 (N_20094,N_16018,N_17591);
and U20095 (N_20095,N_15999,N_17344);
xor U20096 (N_20096,N_15454,N_16542);
xnor U20097 (N_20097,N_17414,N_15972);
xor U20098 (N_20098,N_16902,N_17015);
nor U20099 (N_20099,N_15349,N_16224);
or U20100 (N_20100,N_15499,N_16619);
nor U20101 (N_20101,N_15561,N_15721);
or U20102 (N_20102,N_15439,N_16738);
xnor U20103 (N_20103,N_16332,N_16779);
nor U20104 (N_20104,N_16262,N_15092);
and U20105 (N_20105,N_15428,N_17199);
nand U20106 (N_20106,N_15895,N_15588);
nand U20107 (N_20107,N_17493,N_16904);
and U20108 (N_20108,N_17022,N_17565);
and U20109 (N_20109,N_17139,N_17236);
and U20110 (N_20110,N_17882,N_16180);
xor U20111 (N_20111,N_15738,N_17925);
xor U20112 (N_20112,N_16975,N_15125);
nor U20113 (N_20113,N_15136,N_17506);
nor U20114 (N_20114,N_15111,N_16000);
or U20115 (N_20115,N_17858,N_17263);
or U20116 (N_20116,N_16298,N_16236);
nor U20117 (N_20117,N_16899,N_15071);
and U20118 (N_20118,N_15184,N_15411);
xor U20119 (N_20119,N_17587,N_15923);
and U20120 (N_20120,N_15676,N_16426);
xnor U20121 (N_20121,N_15929,N_15039);
nor U20122 (N_20122,N_15343,N_17947);
nor U20123 (N_20123,N_15602,N_17966);
nor U20124 (N_20124,N_16023,N_16473);
nor U20125 (N_20125,N_15273,N_16489);
or U20126 (N_20126,N_16156,N_16902);
or U20127 (N_20127,N_17945,N_17358);
xnor U20128 (N_20128,N_16741,N_17022);
or U20129 (N_20129,N_15932,N_16992);
xnor U20130 (N_20130,N_17379,N_17143);
xnor U20131 (N_20131,N_15784,N_16762);
or U20132 (N_20132,N_17355,N_16038);
nor U20133 (N_20133,N_15449,N_16186);
nor U20134 (N_20134,N_16540,N_16206);
nand U20135 (N_20135,N_15551,N_17406);
xor U20136 (N_20136,N_16231,N_15411);
or U20137 (N_20137,N_17352,N_15457);
nand U20138 (N_20138,N_17363,N_16819);
xnor U20139 (N_20139,N_16322,N_17250);
xor U20140 (N_20140,N_16023,N_17353);
and U20141 (N_20141,N_16134,N_17024);
nor U20142 (N_20142,N_17749,N_17359);
and U20143 (N_20143,N_17216,N_17156);
and U20144 (N_20144,N_17168,N_15017);
nor U20145 (N_20145,N_17688,N_15911);
and U20146 (N_20146,N_15831,N_17055);
xor U20147 (N_20147,N_15980,N_16107);
or U20148 (N_20148,N_17542,N_15489);
nand U20149 (N_20149,N_17920,N_17622);
nor U20150 (N_20150,N_16636,N_15145);
nand U20151 (N_20151,N_17234,N_16091);
nand U20152 (N_20152,N_16184,N_15755);
nand U20153 (N_20153,N_17798,N_15438);
and U20154 (N_20154,N_15731,N_16367);
nor U20155 (N_20155,N_15141,N_17196);
xnor U20156 (N_20156,N_17434,N_15987);
or U20157 (N_20157,N_15488,N_16919);
nor U20158 (N_20158,N_16574,N_15611);
nand U20159 (N_20159,N_15975,N_16285);
nand U20160 (N_20160,N_16433,N_16794);
xnor U20161 (N_20161,N_16168,N_17536);
nor U20162 (N_20162,N_17380,N_15448);
or U20163 (N_20163,N_17343,N_15757);
nor U20164 (N_20164,N_16780,N_16890);
and U20165 (N_20165,N_15568,N_17620);
xor U20166 (N_20166,N_17631,N_17035);
xnor U20167 (N_20167,N_15745,N_17443);
or U20168 (N_20168,N_16906,N_16037);
and U20169 (N_20169,N_16686,N_16597);
xor U20170 (N_20170,N_16391,N_17094);
or U20171 (N_20171,N_17311,N_17208);
nand U20172 (N_20172,N_16724,N_17313);
nand U20173 (N_20173,N_16959,N_15035);
and U20174 (N_20174,N_16391,N_15329);
and U20175 (N_20175,N_16340,N_17803);
or U20176 (N_20176,N_16320,N_16840);
nor U20177 (N_20177,N_15151,N_16157);
or U20178 (N_20178,N_15497,N_16679);
and U20179 (N_20179,N_16140,N_16429);
and U20180 (N_20180,N_16083,N_15672);
nor U20181 (N_20181,N_15834,N_17801);
nor U20182 (N_20182,N_16080,N_16349);
and U20183 (N_20183,N_17650,N_17455);
nand U20184 (N_20184,N_15757,N_16494);
nor U20185 (N_20185,N_17380,N_16998);
and U20186 (N_20186,N_15129,N_17914);
or U20187 (N_20187,N_16870,N_15779);
and U20188 (N_20188,N_16909,N_16339);
and U20189 (N_20189,N_15764,N_15626);
or U20190 (N_20190,N_15504,N_15881);
nand U20191 (N_20191,N_15309,N_17051);
nor U20192 (N_20192,N_16763,N_17208);
xnor U20193 (N_20193,N_15604,N_17750);
nor U20194 (N_20194,N_16311,N_16941);
xnor U20195 (N_20195,N_16002,N_15617);
or U20196 (N_20196,N_17550,N_15046);
or U20197 (N_20197,N_17127,N_15189);
nand U20198 (N_20198,N_16521,N_17787);
nand U20199 (N_20199,N_17705,N_16534);
nand U20200 (N_20200,N_17457,N_17557);
xor U20201 (N_20201,N_17141,N_16429);
xnor U20202 (N_20202,N_17386,N_17686);
xnor U20203 (N_20203,N_16883,N_17664);
nand U20204 (N_20204,N_17143,N_15008);
and U20205 (N_20205,N_15249,N_17269);
nor U20206 (N_20206,N_15543,N_15189);
and U20207 (N_20207,N_16600,N_15991);
or U20208 (N_20208,N_17274,N_17721);
and U20209 (N_20209,N_17607,N_17737);
nor U20210 (N_20210,N_15131,N_17082);
or U20211 (N_20211,N_17294,N_17710);
or U20212 (N_20212,N_15239,N_17021);
or U20213 (N_20213,N_17598,N_17513);
nand U20214 (N_20214,N_16474,N_15905);
nor U20215 (N_20215,N_15353,N_16189);
nand U20216 (N_20216,N_17291,N_15946);
and U20217 (N_20217,N_15956,N_16997);
and U20218 (N_20218,N_17747,N_17068);
nor U20219 (N_20219,N_17726,N_16076);
or U20220 (N_20220,N_16487,N_16794);
and U20221 (N_20221,N_17905,N_15184);
or U20222 (N_20222,N_17868,N_15930);
and U20223 (N_20223,N_17315,N_16519);
and U20224 (N_20224,N_16408,N_17609);
nor U20225 (N_20225,N_16223,N_16720);
nor U20226 (N_20226,N_17602,N_17395);
xnor U20227 (N_20227,N_16278,N_16019);
or U20228 (N_20228,N_15299,N_15498);
xnor U20229 (N_20229,N_16682,N_15321);
nand U20230 (N_20230,N_16260,N_15108);
xnor U20231 (N_20231,N_17428,N_16226);
and U20232 (N_20232,N_16520,N_17986);
xor U20233 (N_20233,N_15026,N_16427);
and U20234 (N_20234,N_17427,N_17197);
or U20235 (N_20235,N_16728,N_16365);
nand U20236 (N_20236,N_16453,N_17573);
xor U20237 (N_20237,N_17752,N_16513);
or U20238 (N_20238,N_15657,N_17746);
and U20239 (N_20239,N_15525,N_16725);
nand U20240 (N_20240,N_15165,N_17149);
nand U20241 (N_20241,N_16529,N_15022);
nor U20242 (N_20242,N_16974,N_15720);
nor U20243 (N_20243,N_15569,N_17504);
nand U20244 (N_20244,N_17131,N_16641);
nor U20245 (N_20245,N_15272,N_15421);
xnor U20246 (N_20246,N_16456,N_17387);
or U20247 (N_20247,N_15462,N_15972);
xor U20248 (N_20248,N_15392,N_16768);
nand U20249 (N_20249,N_15652,N_15150);
nand U20250 (N_20250,N_17819,N_17426);
and U20251 (N_20251,N_17003,N_16079);
and U20252 (N_20252,N_15466,N_17260);
and U20253 (N_20253,N_16294,N_16898);
xnor U20254 (N_20254,N_17519,N_15107);
and U20255 (N_20255,N_15715,N_17077);
nand U20256 (N_20256,N_15493,N_17139);
nor U20257 (N_20257,N_15009,N_16961);
nor U20258 (N_20258,N_16654,N_16703);
nand U20259 (N_20259,N_17569,N_16158);
nand U20260 (N_20260,N_16254,N_15265);
and U20261 (N_20261,N_17180,N_16250);
and U20262 (N_20262,N_16520,N_16592);
xnor U20263 (N_20263,N_16840,N_17225);
nand U20264 (N_20264,N_16017,N_15605);
xor U20265 (N_20265,N_17198,N_17926);
nand U20266 (N_20266,N_15906,N_17235);
nor U20267 (N_20267,N_15459,N_16929);
nand U20268 (N_20268,N_16315,N_16060);
and U20269 (N_20269,N_16036,N_15083);
or U20270 (N_20270,N_17575,N_17001);
nand U20271 (N_20271,N_15030,N_16178);
nand U20272 (N_20272,N_16120,N_15702);
and U20273 (N_20273,N_17783,N_16782);
nand U20274 (N_20274,N_16971,N_16991);
and U20275 (N_20275,N_17785,N_16579);
or U20276 (N_20276,N_16404,N_16296);
or U20277 (N_20277,N_16073,N_17310);
or U20278 (N_20278,N_15227,N_16782);
nor U20279 (N_20279,N_16326,N_15661);
and U20280 (N_20280,N_16747,N_17858);
xor U20281 (N_20281,N_17192,N_16631);
or U20282 (N_20282,N_15880,N_16069);
xor U20283 (N_20283,N_15172,N_16100);
and U20284 (N_20284,N_17343,N_15562);
nor U20285 (N_20285,N_17279,N_17553);
and U20286 (N_20286,N_16800,N_15128);
and U20287 (N_20287,N_17186,N_17213);
xnor U20288 (N_20288,N_15494,N_15713);
or U20289 (N_20289,N_16944,N_16033);
nor U20290 (N_20290,N_16719,N_17011);
and U20291 (N_20291,N_17215,N_17987);
and U20292 (N_20292,N_16924,N_15396);
xor U20293 (N_20293,N_17472,N_16607);
and U20294 (N_20294,N_17313,N_16835);
xor U20295 (N_20295,N_16543,N_17623);
nand U20296 (N_20296,N_15520,N_16650);
nand U20297 (N_20297,N_15204,N_17035);
xnor U20298 (N_20298,N_16444,N_16628);
nor U20299 (N_20299,N_16527,N_17958);
nor U20300 (N_20300,N_16086,N_17627);
and U20301 (N_20301,N_16307,N_15193);
or U20302 (N_20302,N_17750,N_17439);
xnor U20303 (N_20303,N_16302,N_17544);
nand U20304 (N_20304,N_15591,N_17547);
nand U20305 (N_20305,N_17972,N_17398);
nand U20306 (N_20306,N_17782,N_17287);
nand U20307 (N_20307,N_17463,N_16306);
nand U20308 (N_20308,N_16729,N_15984);
nor U20309 (N_20309,N_17727,N_16848);
and U20310 (N_20310,N_15401,N_17412);
and U20311 (N_20311,N_17556,N_15752);
or U20312 (N_20312,N_15105,N_16110);
or U20313 (N_20313,N_17686,N_17339);
nand U20314 (N_20314,N_17443,N_16713);
nand U20315 (N_20315,N_17750,N_15171);
nand U20316 (N_20316,N_15526,N_16534);
nor U20317 (N_20317,N_15201,N_15286);
xnor U20318 (N_20318,N_16732,N_15823);
and U20319 (N_20319,N_16174,N_16746);
xor U20320 (N_20320,N_15155,N_17455);
xnor U20321 (N_20321,N_16538,N_17415);
nand U20322 (N_20322,N_15294,N_15810);
or U20323 (N_20323,N_15752,N_17374);
or U20324 (N_20324,N_16175,N_15827);
nor U20325 (N_20325,N_16918,N_16214);
nor U20326 (N_20326,N_17287,N_15592);
nand U20327 (N_20327,N_17077,N_15348);
nor U20328 (N_20328,N_16018,N_16917);
nand U20329 (N_20329,N_17356,N_15623);
and U20330 (N_20330,N_16366,N_17959);
and U20331 (N_20331,N_16256,N_17216);
and U20332 (N_20332,N_16772,N_15817);
xnor U20333 (N_20333,N_15829,N_17200);
nor U20334 (N_20334,N_16518,N_17690);
nor U20335 (N_20335,N_15950,N_15758);
nand U20336 (N_20336,N_16689,N_17631);
and U20337 (N_20337,N_15107,N_17660);
or U20338 (N_20338,N_16381,N_16553);
or U20339 (N_20339,N_17108,N_16896);
and U20340 (N_20340,N_15781,N_17984);
and U20341 (N_20341,N_15819,N_15979);
or U20342 (N_20342,N_16017,N_15064);
or U20343 (N_20343,N_16897,N_17695);
and U20344 (N_20344,N_16168,N_15557);
nand U20345 (N_20345,N_17383,N_16654);
nand U20346 (N_20346,N_15929,N_16784);
nand U20347 (N_20347,N_15447,N_16664);
nor U20348 (N_20348,N_17478,N_15276);
nand U20349 (N_20349,N_16071,N_16426);
or U20350 (N_20350,N_17475,N_15758);
and U20351 (N_20351,N_16910,N_16362);
nand U20352 (N_20352,N_15895,N_15798);
xor U20353 (N_20353,N_15679,N_17800);
nor U20354 (N_20354,N_15338,N_15632);
xor U20355 (N_20355,N_17751,N_16818);
xor U20356 (N_20356,N_17384,N_16387);
xnor U20357 (N_20357,N_15642,N_16559);
and U20358 (N_20358,N_17123,N_16940);
xor U20359 (N_20359,N_15220,N_15208);
nand U20360 (N_20360,N_15782,N_15633);
nor U20361 (N_20361,N_15910,N_15204);
xnor U20362 (N_20362,N_15136,N_17512);
xor U20363 (N_20363,N_15099,N_15336);
xnor U20364 (N_20364,N_17215,N_17915);
nand U20365 (N_20365,N_17844,N_16019);
xnor U20366 (N_20366,N_15184,N_17081);
or U20367 (N_20367,N_16292,N_17027);
and U20368 (N_20368,N_16957,N_17978);
or U20369 (N_20369,N_16611,N_15278);
nand U20370 (N_20370,N_17095,N_17625);
nor U20371 (N_20371,N_15083,N_15717);
nand U20372 (N_20372,N_16829,N_16376);
and U20373 (N_20373,N_15934,N_16422);
and U20374 (N_20374,N_15498,N_15037);
nor U20375 (N_20375,N_17345,N_16453);
nand U20376 (N_20376,N_15050,N_16099);
nand U20377 (N_20377,N_17195,N_17167);
nor U20378 (N_20378,N_16770,N_16914);
nor U20379 (N_20379,N_17634,N_15432);
or U20380 (N_20380,N_15182,N_17242);
xnor U20381 (N_20381,N_17588,N_17098);
xnor U20382 (N_20382,N_17627,N_16319);
nor U20383 (N_20383,N_17182,N_16205);
xor U20384 (N_20384,N_17678,N_17425);
nor U20385 (N_20385,N_17913,N_15825);
nand U20386 (N_20386,N_15661,N_16072);
or U20387 (N_20387,N_17923,N_17832);
nand U20388 (N_20388,N_17729,N_16350);
xor U20389 (N_20389,N_16134,N_17946);
or U20390 (N_20390,N_16735,N_16908);
nor U20391 (N_20391,N_17604,N_15872);
nor U20392 (N_20392,N_15034,N_15074);
and U20393 (N_20393,N_15971,N_17725);
and U20394 (N_20394,N_15210,N_16591);
nor U20395 (N_20395,N_17677,N_17827);
nand U20396 (N_20396,N_16084,N_15906);
and U20397 (N_20397,N_15792,N_15708);
nor U20398 (N_20398,N_16809,N_15288);
xnor U20399 (N_20399,N_17868,N_16351);
xor U20400 (N_20400,N_16046,N_16476);
and U20401 (N_20401,N_17222,N_17376);
nand U20402 (N_20402,N_15996,N_17168);
nand U20403 (N_20403,N_15743,N_16408);
or U20404 (N_20404,N_17690,N_16201);
nand U20405 (N_20405,N_15255,N_17774);
or U20406 (N_20406,N_16269,N_15150);
or U20407 (N_20407,N_16892,N_15215);
and U20408 (N_20408,N_15429,N_17182);
nand U20409 (N_20409,N_16275,N_15291);
nor U20410 (N_20410,N_16024,N_17609);
nor U20411 (N_20411,N_17735,N_15893);
xnor U20412 (N_20412,N_15538,N_15116);
and U20413 (N_20413,N_15991,N_17897);
xnor U20414 (N_20414,N_16923,N_15857);
or U20415 (N_20415,N_16359,N_17149);
or U20416 (N_20416,N_17799,N_16732);
or U20417 (N_20417,N_16010,N_16638);
xnor U20418 (N_20418,N_15734,N_17917);
xor U20419 (N_20419,N_16336,N_17082);
or U20420 (N_20420,N_15407,N_17102);
and U20421 (N_20421,N_15101,N_16082);
and U20422 (N_20422,N_15634,N_17438);
and U20423 (N_20423,N_16643,N_16435);
nand U20424 (N_20424,N_16383,N_15039);
nand U20425 (N_20425,N_15982,N_17600);
or U20426 (N_20426,N_15455,N_15137);
and U20427 (N_20427,N_17210,N_15902);
and U20428 (N_20428,N_17713,N_16007);
xor U20429 (N_20429,N_17253,N_15397);
and U20430 (N_20430,N_15989,N_16768);
nand U20431 (N_20431,N_15771,N_17640);
or U20432 (N_20432,N_17846,N_16872);
and U20433 (N_20433,N_16726,N_17024);
nor U20434 (N_20434,N_16469,N_15483);
and U20435 (N_20435,N_15016,N_16491);
or U20436 (N_20436,N_15151,N_15958);
and U20437 (N_20437,N_17086,N_16552);
nor U20438 (N_20438,N_17973,N_15709);
or U20439 (N_20439,N_17803,N_16105);
or U20440 (N_20440,N_15217,N_15128);
nand U20441 (N_20441,N_16420,N_17980);
xor U20442 (N_20442,N_17748,N_17828);
nand U20443 (N_20443,N_15754,N_15811);
nor U20444 (N_20444,N_17671,N_16021);
nand U20445 (N_20445,N_16167,N_16618);
xnor U20446 (N_20446,N_16495,N_15193);
and U20447 (N_20447,N_15103,N_17724);
nor U20448 (N_20448,N_17069,N_16701);
nor U20449 (N_20449,N_15846,N_17981);
nor U20450 (N_20450,N_16298,N_15731);
and U20451 (N_20451,N_16265,N_17740);
nor U20452 (N_20452,N_17308,N_17132);
nand U20453 (N_20453,N_17355,N_15892);
and U20454 (N_20454,N_17325,N_16767);
xnor U20455 (N_20455,N_15552,N_15680);
xor U20456 (N_20456,N_15281,N_17456);
and U20457 (N_20457,N_16912,N_15623);
nand U20458 (N_20458,N_16083,N_16866);
or U20459 (N_20459,N_16394,N_16670);
nand U20460 (N_20460,N_15894,N_17395);
xor U20461 (N_20461,N_15018,N_16605);
and U20462 (N_20462,N_16979,N_16356);
nand U20463 (N_20463,N_15403,N_15778);
nand U20464 (N_20464,N_17886,N_17318);
nor U20465 (N_20465,N_17520,N_15731);
and U20466 (N_20466,N_16615,N_15562);
nor U20467 (N_20467,N_16430,N_15199);
nand U20468 (N_20468,N_17830,N_16073);
or U20469 (N_20469,N_17530,N_17393);
or U20470 (N_20470,N_15754,N_17038);
and U20471 (N_20471,N_17683,N_17792);
or U20472 (N_20472,N_17063,N_15469);
nand U20473 (N_20473,N_15453,N_15729);
or U20474 (N_20474,N_16961,N_15377);
nor U20475 (N_20475,N_15620,N_15222);
or U20476 (N_20476,N_15399,N_16550);
or U20477 (N_20477,N_16756,N_15504);
nor U20478 (N_20478,N_15716,N_16707);
nor U20479 (N_20479,N_15770,N_15397);
or U20480 (N_20480,N_17082,N_15475);
or U20481 (N_20481,N_17281,N_15727);
or U20482 (N_20482,N_15939,N_16927);
nand U20483 (N_20483,N_17202,N_16103);
or U20484 (N_20484,N_15876,N_16371);
nand U20485 (N_20485,N_17774,N_15848);
xnor U20486 (N_20486,N_16002,N_16493);
nand U20487 (N_20487,N_15612,N_16112);
nor U20488 (N_20488,N_15896,N_15930);
xnor U20489 (N_20489,N_17231,N_16769);
xnor U20490 (N_20490,N_15782,N_16362);
or U20491 (N_20491,N_17899,N_15247);
or U20492 (N_20492,N_15165,N_15883);
nand U20493 (N_20493,N_17314,N_15895);
nor U20494 (N_20494,N_17758,N_15325);
nand U20495 (N_20495,N_16740,N_15177);
xor U20496 (N_20496,N_16748,N_16610);
nor U20497 (N_20497,N_15893,N_16609);
and U20498 (N_20498,N_16236,N_17546);
nor U20499 (N_20499,N_16622,N_16294);
nand U20500 (N_20500,N_16332,N_15223);
nand U20501 (N_20501,N_16046,N_17607);
xor U20502 (N_20502,N_15184,N_15193);
and U20503 (N_20503,N_17331,N_16699);
or U20504 (N_20504,N_15867,N_15206);
and U20505 (N_20505,N_17748,N_16702);
and U20506 (N_20506,N_17384,N_15456);
xnor U20507 (N_20507,N_15667,N_17682);
xor U20508 (N_20508,N_16116,N_15520);
nor U20509 (N_20509,N_16946,N_17579);
and U20510 (N_20510,N_15077,N_15090);
and U20511 (N_20511,N_17696,N_17278);
nor U20512 (N_20512,N_17890,N_16473);
or U20513 (N_20513,N_17397,N_17724);
nor U20514 (N_20514,N_16696,N_15422);
and U20515 (N_20515,N_17586,N_16568);
and U20516 (N_20516,N_16568,N_15820);
xor U20517 (N_20517,N_16131,N_15141);
nor U20518 (N_20518,N_16620,N_17757);
nand U20519 (N_20519,N_16210,N_16631);
nand U20520 (N_20520,N_15192,N_17240);
and U20521 (N_20521,N_15651,N_17564);
xnor U20522 (N_20522,N_15718,N_15440);
and U20523 (N_20523,N_16262,N_16938);
nor U20524 (N_20524,N_15484,N_17790);
or U20525 (N_20525,N_17149,N_16533);
xor U20526 (N_20526,N_15878,N_17908);
or U20527 (N_20527,N_16232,N_15938);
or U20528 (N_20528,N_17850,N_17460);
and U20529 (N_20529,N_16007,N_16603);
or U20530 (N_20530,N_16167,N_17732);
nand U20531 (N_20531,N_17934,N_15257);
nand U20532 (N_20532,N_15973,N_16422);
nand U20533 (N_20533,N_17260,N_17387);
xor U20534 (N_20534,N_15349,N_16396);
or U20535 (N_20535,N_16949,N_17512);
xnor U20536 (N_20536,N_15031,N_16804);
or U20537 (N_20537,N_15910,N_17380);
or U20538 (N_20538,N_17657,N_16450);
nor U20539 (N_20539,N_17702,N_17292);
xnor U20540 (N_20540,N_17047,N_15579);
xnor U20541 (N_20541,N_17795,N_16985);
nor U20542 (N_20542,N_17268,N_15265);
nand U20543 (N_20543,N_17370,N_15775);
nor U20544 (N_20544,N_15208,N_16949);
nand U20545 (N_20545,N_15340,N_16937);
nand U20546 (N_20546,N_16411,N_16876);
xor U20547 (N_20547,N_15166,N_17204);
xnor U20548 (N_20548,N_16230,N_16840);
xor U20549 (N_20549,N_15767,N_17544);
xor U20550 (N_20550,N_17240,N_15808);
and U20551 (N_20551,N_15191,N_16056);
nand U20552 (N_20552,N_16226,N_17005);
or U20553 (N_20553,N_16346,N_16799);
xor U20554 (N_20554,N_17077,N_16390);
and U20555 (N_20555,N_15869,N_16618);
and U20556 (N_20556,N_15501,N_17496);
xnor U20557 (N_20557,N_16389,N_16588);
nor U20558 (N_20558,N_17206,N_17453);
nand U20559 (N_20559,N_15200,N_17635);
and U20560 (N_20560,N_17107,N_15617);
xor U20561 (N_20561,N_17934,N_16749);
nand U20562 (N_20562,N_17189,N_16707);
and U20563 (N_20563,N_15845,N_17116);
nor U20564 (N_20564,N_16917,N_16900);
or U20565 (N_20565,N_15626,N_17821);
nor U20566 (N_20566,N_15667,N_15771);
or U20567 (N_20567,N_17732,N_17325);
nand U20568 (N_20568,N_17157,N_16120);
nand U20569 (N_20569,N_17353,N_16732);
or U20570 (N_20570,N_16539,N_15779);
nand U20571 (N_20571,N_15969,N_16657);
or U20572 (N_20572,N_17031,N_15642);
and U20573 (N_20573,N_16135,N_15671);
xnor U20574 (N_20574,N_17288,N_17872);
nor U20575 (N_20575,N_17504,N_16616);
xnor U20576 (N_20576,N_16623,N_16485);
xor U20577 (N_20577,N_17621,N_17213);
xnor U20578 (N_20578,N_15768,N_17962);
nor U20579 (N_20579,N_15163,N_15423);
and U20580 (N_20580,N_15562,N_16327);
xnor U20581 (N_20581,N_16287,N_16693);
nand U20582 (N_20582,N_17492,N_16564);
or U20583 (N_20583,N_17584,N_15021);
and U20584 (N_20584,N_17466,N_16376);
or U20585 (N_20585,N_16335,N_17270);
xnor U20586 (N_20586,N_15292,N_16145);
nand U20587 (N_20587,N_16558,N_15236);
xor U20588 (N_20588,N_16982,N_15362);
or U20589 (N_20589,N_16335,N_16953);
nor U20590 (N_20590,N_16733,N_17718);
and U20591 (N_20591,N_15375,N_16523);
nand U20592 (N_20592,N_15673,N_15625);
or U20593 (N_20593,N_17166,N_16481);
nand U20594 (N_20594,N_17618,N_17718);
nor U20595 (N_20595,N_15790,N_16980);
or U20596 (N_20596,N_16187,N_17547);
or U20597 (N_20597,N_17866,N_17233);
nor U20598 (N_20598,N_17795,N_15809);
nand U20599 (N_20599,N_16746,N_15951);
or U20600 (N_20600,N_16216,N_17119);
nand U20601 (N_20601,N_16318,N_15123);
or U20602 (N_20602,N_17542,N_15335);
nand U20603 (N_20603,N_15953,N_16076);
nand U20604 (N_20604,N_15025,N_16427);
or U20605 (N_20605,N_16738,N_16613);
nand U20606 (N_20606,N_15256,N_15245);
nand U20607 (N_20607,N_17634,N_17382);
nor U20608 (N_20608,N_17757,N_15149);
xnor U20609 (N_20609,N_16277,N_15169);
and U20610 (N_20610,N_17999,N_16480);
nand U20611 (N_20611,N_17457,N_17463);
and U20612 (N_20612,N_15666,N_16118);
nand U20613 (N_20613,N_15060,N_16654);
or U20614 (N_20614,N_16218,N_17858);
xor U20615 (N_20615,N_15160,N_17883);
xor U20616 (N_20616,N_16846,N_17127);
xnor U20617 (N_20617,N_17713,N_15444);
or U20618 (N_20618,N_15853,N_15708);
nor U20619 (N_20619,N_16093,N_17176);
nand U20620 (N_20620,N_16191,N_15030);
and U20621 (N_20621,N_16130,N_15858);
xnor U20622 (N_20622,N_16833,N_16812);
or U20623 (N_20623,N_15132,N_17540);
and U20624 (N_20624,N_16566,N_17468);
or U20625 (N_20625,N_15626,N_17148);
and U20626 (N_20626,N_16609,N_17644);
nand U20627 (N_20627,N_15340,N_17850);
nor U20628 (N_20628,N_15290,N_16141);
nor U20629 (N_20629,N_15202,N_15496);
nand U20630 (N_20630,N_17336,N_16445);
or U20631 (N_20631,N_16817,N_15790);
nand U20632 (N_20632,N_16895,N_15968);
nor U20633 (N_20633,N_15713,N_17543);
or U20634 (N_20634,N_17490,N_15559);
or U20635 (N_20635,N_17446,N_16798);
or U20636 (N_20636,N_15877,N_15534);
nand U20637 (N_20637,N_17394,N_15972);
or U20638 (N_20638,N_17699,N_16632);
and U20639 (N_20639,N_17202,N_16997);
and U20640 (N_20640,N_16751,N_17547);
nand U20641 (N_20641,N_16811,N_15834);
xnor U20642 (N_20642,N_16733,N_16826);
or U20643 (N_20643,N_17160,N_16581);
or U20644 (N_20644,N_17021,N_15686);
and U20645 (N_20645,N_15214,N_15641);
nor U20646 (N_20646,N_17561,N_15287);
xor U20647 (N_20647,N_17890,N_16073);
xnor U20648 (N_20648,N_17860,N_16280);
or U20649 (N_20649,N_16294,N_16117);
xor U20650 (N_20650,N_16923,N_17531);
nand U20651 (N_20651,N_16036,N_15552);
or U20652 (N_20652,N_17760,N_17750);
nand U20653 (N_20653,N_16900,N_15762);
nand U20654 (N_20654,N_16830,N_15821);
xnor U20655 (N_20655,N_16477,N_16891);
or U20656 (N_20656,N_15647,N_17522);
xnor U20657 (N_20657,N_15522,N_17920);
and U20658 (N_20658,N_15671,N_17106);
xor U20659 (N_20659,N_17878,N_16778);
and U20660 (N_20660,N_16921,N_17198);
and U20661 (N_20661,N_17486,N_15657);
or U20662 (N_20662,N_15437,N_15142);
nor U20663 (N_20663,N_17268,N_15134);
or U20664 (N_20664,N_17543,N_15723);
and U20665 (N_20665,N_15623,N_16901);
and U20666 (N_20666,N_17386,N_15967);
nor U20667 (N_20667,N_15404,N_15810);
or U20668 (N_20668,N_17987,N_15700);
or U20669 (N_20669,N_16879,N_16334);
nand U20670 (N_20670,N_16646,N_16716);
or U20671 (N_20671,N_15935,N_15669);
xor U20672 (N_20672,N_16921,N_17260);
xnor U20673 (N_20673,N_15855,N_16047);
nor U20674 (N_20674,N_15534,N_15744);
xor U20675 (N_20675,N_17914,N_16457);
xnor U20676 (N_20676,N_17609,N_15915);
and U20677 (N_20677,N_15823,N_16849);
xor U20678 (N_20678,N_17724,N_17363);
and U20679 (N_20679,N_17083,N_16757);
or U20680 (N_20680,N_16536,N_17374);
nor U20681 (N_20681,N_15362,N_17485);
nor U20682 (N_20682,N_16311,N_17000);
nor U20683 (N_20683,N_17768,N_16666);
and U20684 (N_20684,N_16504,N_15650);
nand U20685 (N_20685,N_15780,N_15454);
xnor U20686 (N_20686,N_15718,N_16902);
or U20687 (N_20687,N_16370,N_17792);
or U20688 (N_20688,N_17296,N_15427);
xor U20689 (N_20689,N_17586,N_17961);
xnor U20690 (N_20690,N_16578,N_15612);
xor U20691 (N_20691,N_15426,N_15389);
xnor U20692 (N_20692,N_17117,N_17296);
and U20693 (N_20693,N_16447,N_17655);
xnor U20694 (N_20694,N_17684,N_16277);
xor U20695 (N_20695,N_17419,N_15491);
xnor U20696 (N_20696,N_15126,N_16191);
nor U20697 (N_20697,N_16514,N_16116);
nor U20698 (N_20698,N_17059,N_17381);
nor U20699 (N_20699,N_17344,N_16759);
nand U20700 (N_20700,N_17652,N_17545);
nand U20701 (N_20701,N_16239,N_16861);
or U20702 (N_20702,N_15881,N_17981);
nor U20703 (N_20703,N_17686,N_15038);
nand U20704 (N_20704,N_16760,N_17819);
xor U20705 (N_20705,N_15645,N_16453);
and U20706 (N_20706,N_17337,N_17770);
nor U20707 (N_20707,N_15723,N_17674);
nor U20708 (N_20708,N_15808,N_15422);
or U20709 (N_20709,N_17951,N_16740);
and U20710 (N_20710,N_15339,N_17950);
nor U20711 (N_20711,N_17972,N_16337);
nand U20712 (N_20712,N_17826,N_16316);
and U20713 (N_20713,N_17463,N_15289);
or U20714 (N_20714,N_17791,N_17827);
xor U20715 (N_20715,N_15071,N_16135);
xor U20716 (N_20716,N_16971,N_17534);
xnor U20717 (N_20717,N_17421,N_15896);
and U20718 (N_20718,N_16773,N_15115);
xnor U20719 (N_20719,N_17772,N_16416);
xnor U20720 (N_20720,N_15350,N_15807);
xor U20721 (N_20721,N_17087,N_16877);
nor U20722 (N_20722,N_15428,N_15495);
xnor U20723 (N_20723,N_15045,N_15389);
or U20724 (N_20724,N_17994,N_17252);
nor U20725 (N_20725,N_15951,N_16011);
xnor U20726 (N_20726,N_16090,N_15960);
xnor U20727 (N_20727,N_16564,N_17420);
nor U20728 (N_20728,N_15938,N_17460);
or U20729 (N_20729,N_15360,N_17963);
nand U20730 (N_20730,N_17780,N_16796);
or U20731 (N_20731,N_15946,N_16979);
and U20732 (N_20732,N_15288,N_17649);
xnor U20733 (N_20733,N_16080,N_16784);
nor U20734 (N_20734,N_15216,N_17525);
or U20735 (N_20735,N_15575,N_15258);
xor U20736 (N_20736,N_15171,N_15402);
xor U20737 (N_20737,N_17469,N_16552);
and U20738 (N_20738,N_17472,N_16023);
and U20739 (N_20739,N_16430,N_17661);
or U20740 (N_20740,N_17891,N_15739);
xnor U20741 (N_20741,N_15875,N_17242);
and U20742 (N_20742,N_17573,N_17818);
nand U20743 (N_20743,N_16137,N_17167);
nor U20744 (N_20744,N_16568,N_15584);
and U20745 (N_20745,N_16480,N_17433);
nand U20746 (N_20746,N_17058,N_15429);
and U20747 (N_20747,N_16157,N_16814);
and U20748 (N_20748,N_17292,N_17588);
or U20749 (N_20749,N_17463,N_16103);
xor U20750 (N_20750,N_16451,N_16606);
and U20751 (N_20751,N_16017,N_15267);
nand U20752 (N_20752,N_16357,N_17550);
xnor U20753 (N_20753,N_15347,N_16762);
xor U20754 (N_20754,N_17105,N_16325);
nand U20755 (N_20755,N_15725,N_15710);
xor U20756 (N_20756,N_16280,N_17620);
xor U20757 (N_20757,N_17412,N_17838);
or U20758 (N_20758,N_17677,N_16913);
nor U20759 (N_20759,N_16488,N_16849);
nand U20760 (N_20760,N_15793,N_17109);
nor U20761 (N_20761,N_17873,N_15704);
or U20762 (N_20762,N_15026,N_17778);
xor U20763 (N_20763,N_17219,N_16693);
xnor U20764 (N_20764,N_16441,N_16208);
nor U20765 (N_20765,N_17402,N_16607);
nand U20766 (N_20766,N_15392,N_16264);
nor U20767 (N_20767,N_16103,N_15038);
and U20768 (N_20768,N_15563,N_15920);
xor U20769 (N_20769,N_15767,N_15776);
nand U20770 (N_20770,N_15505,N_15570);
nor U20771 (N_20771,N_17029,N_16557);
or U20772 (N_20772,N_17771,N_15430);
and U20773 (N_20773,N_16711,N_15353);
nor U20774 (N_20774,N_17776,N_16480);
or U20775 (N_20775,N_15766,N_15054);
nor U20776 (N_20776,N_17541,N_16577);
or U20777 (N_20777,N_15715,N_17583);
xnor U20778 (N_20778,N_17856,N_16271);
nand U20779 (N_20779,N_16927,N_15279);
and U20780 (N_20780,N_16859,N_16064);
nor U20781 (N_20781,N_15512,N_15529);
and U20782 (N_20782,N_16863,N_17636);
and U20783 (N_20783,N_15557,N_15610);
nand U20784 (N_20784,N_15897,N_17232);
or U20785 (N_20785,N_16175,N_15876);
xnor U20786 (N_20786,N_16801,N_15143);
nor U20787 (N_20787,N_15052,N_16852);
xor U20788 (N_20788,N_15501,N_17128);
and U20789 (N_20789,N_17534,N_16617);
or U20790 (N_20790,N_15468,N_16176);
and U20791 (N_20791,N_15293,N_15419);
nand U20792 (N_20792,N_16248,N_16951);
nand U20793 (N_20793,N_15794,N_16244);
nand U20794 (N_20794,N_16169,N_15906);
nand U20795 (N_20795,N_16376,N_17235);
nor U20796 (N_20796,N_16674,N_15222);
nand U20797 (N_20797,N_15058,N_16543);
or U20798 (N_20798,N_15288,N_17545);
and U20799 (N_20799,N_16348,N_17259);
nor U20800 (N_20800,N_15212,N_16044);
and U20801 (N_20801,N_16919,N_17862);
or U20802 (N_20802,N_16545,N_15827);
or U20803 (N_20803,N_17906,N_15690);
nor U20804 (N_20804,N_15707,N_16411);
nand U20805 (N_20805,N_15925,N_15805);
xnor U20806 (N_20806,N_16146,N_17973);
and U20807 (N_20807,N_15158,N_17094);
and U20808 (N_20808,N_15777,N_15950);
xnor U20809 (N_20809,N_17512,N_17169);
or U20810 (N_20810,N_15608,N_15377);
xor U20811 (N_20811,N_15251,N_16900);
and U20812 (N_20812,N_15797,N_15097);
xnor U20813 (N_20813,N_17534,N_17491);
and U20814 (N_20814,N_15017,N_16580);
nand U20815 (N_20815,N_15341,N_15357);
or U20816 (N_20816,N_15367,N_16139);
and U20817 (N_20817,N_15023,N_17273);
xor U20818 (N_20818,N_17407,N_15615);
or U20819 (N_20819,N_15845,N_16784);
nor U20820 (N_20820,N_15419,N_16242);
or U20821 (N_20821,N_15133,N_16277);
and U20822 (N_20822,N_15166,N_15076);
nand U20823 (N_20823,N_16798,N_17828);
or U20824 (N_20824,N_17761,N_17842);
nor U20825 (N_20825,N_17746,N_17535);
xnor U20826 (N_20826,N_17477,N_17815);
or U20827 (N_20827,N_15425,N_16339);
xnor U20828 (N_20828,N_15056,N_15959);
xnor U20829 (N_20829,N_16246,N_16917);
xor U20830 (N_20830,N_17641,N_16877);
and U20831 (N_20831,N_17496,N_16420);
xnor U20832 (N_20832,N_15844,N_15766);
and U20833 (N_20833,N_17715,N_16293);
xnor U20834 (N_20834,N_17577,N_16905);
xnor U20835 (N_20835,N_16745,N_17738);
nor U20836 (N_20836,N_17665,N_15752);
and U20837 (N_20837,N_16915,N_16822);
nand U20838 (N_20838,N_17379,N_16832);
xnor U20839 (N_20839,N_15795,N_16077);
xnor U20840 (N_20840,N_17082,N_16772);
nand U20841 (N_20841,N_16564,N_17179);
nand U20842 (N_20842,N_17300,N_17262);
and U20843 (N_20843,N_16367,N_16227);
nor U20844 (N_20844,N_15842,N_17199);
and U20845 (N_20845,N_15375,N_16613);
or U20846 (N_20846,N_17079,N_15559);
xor U20847 (N_20847,N_17767,N_17344);
nor U20848 (N_20848,N_16801,N_16140);
xor U20849 (N_20849,N_15902,N_17672);
nor U20850 (N_20850,N_16161,N_17458);
nor U20851 (N_20851,N_16493,N_15990);
and U20852 (N_20852,N_17674,N_17702);
nand U20853 (N_20853,N_17176,N_17412);
nor U20854 (N_20854,N_16175,N_16834);
nor U20855 (N_20855,N_16654,N_17603);
xor U20856 (N_20856,N_17734,N_15405);
nand U20857 (N_20857,N_17727,N_17131);
or U20858 (N_20858,N_17469,N_16500);
xor U20859 (N_20859,N_17905,N_16291);
or U20860 (N_20860,N_16596,N_16015);
nand U20861 (N_20861,N_16015,N_15857);
or U20862 (N_20862,N_16723,N_16384);
nand U20863 (N_20863,N_16622,N_15933);
and U20864 (N_20864,N_16944,N_16932);
nor U20865 (N_20865,N_15918,N_15601);
nand U20866 (N_20866,N_17098,N_16718);
nor U20867 (N_20867,N_16349,N_16545);
and U20868 (N_20868,N_17517,N_17990);
nand U20869 (N_20869,N_16753,N_15935);
xnor U20870 (N_20870,N_17218,N_17539);
nor U20871 (N_20871,N_15210,N_16776);
xnor U20872 (N_20872,N_15297,N_15089);
or U20873 (N_20873,N_16883,N_17192);
and U20874 (N_20874,N_17321,N_15080);
or U20875 (N_20875,N_17829,N_15030);
nor U20876 (N_20876,N_17357,N_17913);
and U20877 (N_20877,N_17765,N_17438);
nand U20878 (N_20878,N_16500,N_15100);
nor U20879 (N_20879,N_16067,N_16068);
and U20880 (N_20880,N_15571,N_16150);
xor U20881 (N_20881,N_17471,N_16756);
nand U20882 (N_20882,N_16036,N_15793);
nand U20883 (N_20883,N_15868,N_17326);
or U20884 (N_20884,N_17226,N_16483);
nand U20885 (N_20885,N_16235,N_15135);
nand U20886 (N_20886,N_15008,N_16472);
and U20887 (N_20887,N_15917,N_15783);
nor U20888 (N_20888,N_15125,N_16410);
and U20889 (N_20889,N_16731,N_15824);
xor U20890 (N_20890,N_16346,N_15373);
nor U20891 (N_20891,N_16146,N_15536);
or U20892 (N_20892,N_16564,N_17601);
xor U20893 (N_20893,N_17074,N_16788);
or U20894 (N_20894,N_15593,N_15101);
xor U20895 (N_20895,N_15189,N_16813);
or U20896 (N_20896,N_15743,N_15552);
and U20897 (N_20897,N_16425,N_17904);
nand U20898 (N_20898,N_17462,N_15740);
xnor U20899 (N_20899,N_15273,N_15511);
nor U20900 (N_20900,N_17842,N_17926);
nand U20901 (N_20901,N_15192,N_17724);
nor U20902 (N_20902,N_15904,N_15143);
nor U20903 (N_20903,N_15864,N_15060);
nor U20904 (N_20904,N_15630,N_16631);
nor U20905 (N_20905,N_16732,N_17492);
and U20906 (N_20906,N_15154,N_15057);
and U20907 (N_20907,N_16542,N_16449);
nand U20908 (N_20908,N_15470,N_17179);
nor U20909 (N_20909,N_15395,N_15864);
nor U20910 (N_20910,N_15384,N_16443);
or U20911 (N_20911,N_15219,N_17498);
nor U20912 (N_20912,N_16455,N_15047);
and U20913 (N_20913,N_15435,N_16026);
nand U20914 (N_20914,N_16824,N_15384);
xnor U20915 (N_20915,N_16326,N_16587);
or U20916 (N_20916,N_16084,N_15081);
xor U20917 (N_20917,N_15792,N_16468);
nor U20918 (N_20918,N_16129,N_15425);
or U20919 (N_20919,N_15846,N_15913);
and U20920 (N_20920,N_15698,N_15252);
or U20921 (N_20921,N_16296,N_16893);
nor U20922 (N_20922,N_15364,N_15340);
nor U20923 (N_20923,N_15790,N_17410);
or U20924 (N_20924,N_16993,N_15630);
or U20925 (N_20925,N_16629,N_16920);
and U20926 (N_20926,N_17952,N_15467);
nand U20927 (N_20927,N_17223,N_15423);
nand U20928 (N_20928,N_15541,N_16910);
and U20929 (N_20929,N_16793,N_15435);
nor U20930 (N_20930,N_17520,N_16490);
and U20931 (N_20931,N_17612,N_16016);
or U20932 (N_20932,N_17705,N_16171);
xor U20933 (N_20933,N_17018,N_17002);
xnor U20934 (N_20934,N_16767,N_17514);
xor U20935 (N_20935,N_17421,N_17166);
xnor U20936 (N_20936,N_16924,N_16114);
or U20937 (N_20937,N_17945,N_15907);
and U20938 (N_20938,N_15901,N_15320);
or U20939 (N_20939,N_16821,N_16692);
or U20940 (N_20940,N_15974,N_15076);
or U20941 (N_20941,N_16862,N_17071);
or U20942 (N_20942,N_15315,N_17600);
nor U20943 (N_20943,N_16030,N_15790);
nor U20944 (N_20944,N_16814,N_17375);
nor U20945 (N_20945,N_16730,N_17854);
or U20946 (N_20946,N_17164,N_15681);
nand U20947 (N_20947,N_16370,N_16751);
xnor U20948 (N_20948,N_17768,N_16925);
and U20949 (N_20949,N_17327,N_17050);
nor U20950 (N_20950,N_17839,N_17147);
and U20951 (N_20951,N_17751,N_17481);
nand U20952 (N_20952,N_15914,N_17501);
nand U20953 (N_20953,N_17006,N_17050);
nor U20954 (N_20954,N_15316,N_16608);
nand U20955 (N_20955,N_15292,N_15736);
or U20956 (N_20956,N_15964,N_16608);
or U20957 (N_20957,N_17643,N_17471);
xnor U20958 (N_20958,N_16093,N_17986);
xor U20959 (N_20959,N_17177,N_15828);
or U20960 (N_20960,N_15605,N_15637);
nor U20961 (N_20961,N_17849,N_16270);
nor U20962 (N_20962,N_16654,N_15130);
or U20963 (N_20963,N_16113,N_15048);
xnor U20964 (N_20964,N_16456,N_15878);
nand U20965 (N_20965,N_16168,N_16549);
xnor U20966 (N_20966,N_15113,N_16607);
xnor U20967 (N_20967,N_15190,N_16840);
or U20968 (N_20968,N_15916,N_15240);
xor U20969 (N_20969,N_16030,N_16676);
and U20970 (N_20970,N_16146,N_16762);
xor U20971 (N_20971,N_15595,N_15552);
xor U20972 (N_20972,N_16663,N_15483);
or U20973 (N_20973,N_15239,N_15455);
or U20974 (N_20974,N_17509,N_17477);
xnor U20975 (N_20975,N_15912,N_15572);
or U20976 (N_20976,N_15054,N_15719);
and U20977 (N_20977,N_16582,N_15359);
nor U20978 (N_20978,N_17576,N_17328);
nand U20979 (N_20979,N_17130,N_16478);
nand U20980 (N_20980,N_15329,N_15107);
nand U20981 (N_20981,N_17590,N_17018);
nor U20982 (N_20982,N_16772,N_15517);
and U20983 (N_20983,N_15446,N_16874);
and U20984 (N_20984,N_16565,N_15075);
xnor U20985 (N_20985,N_16211,N_15786);
nand U20986 (N_20986,N_17377,N_17526);
xnor U20987 (N_20987,N_16338,N_15316);
and U20988 (N_20988,N_15027,N_16898);
nor U20989 (N_20989,N_15264,N_16003);
nor U20990 (N_20990,N_15105,N_17221);
or U20991 (N_20991,N_16763,N_17915);
nor U20992 (N_20992,N_17845,N_15422);
xnor U20993 (N_20993,N_15681,N_17389);
and U20994 (N_20994,N_17428,N_16912);
xor U20995 (N_20995,N_15370,N_15267);
nand U20996 (N_20996,N_16843,N_17836);
and U20997 (N_20997,N_17932,N_16241);
or U20998 (N_20998,N_17905,N_17734);
nand U20999 (N_20999,N_15703,N_17648);
xnor U21000 (N_21000,N_19252,N_20537);
nor U21001 (N_21001,N_18609,N_20457);
nor U21002 (N_21002,N_19707,N_18746);
and U21003 (N_21003,N_19161,N_18629);
and U21004 (N_21004,N_18909,N_19761);
nor U21005 (N_21005,N_19820,N_19106);
nand U21006 (N_21006,N_19262,N_19705);
nor U21007 (N_21007,N_20939,N_18017);
nand U21008 (N_21008,N_18992,N_18387);
and U21009 (N_21009,N_19101,N_19921);
xor U21010 (N_21010,N_18286,N_19347);
and U21011 (N_21011,N_18434,N_20616);
or U21012 (N_21012,N_18213,N_19778);
xor U21013 (N_21013,N_20302,N_19170);
or U21014 (N_21014,N_18329,N_20137);
nand U21015 (N_21015,N_18567,N_19397);
nor U21016 (N_21016,N_19677,N_18123);
or U21017 (N_21017,N_18845,N_20999);
and U21018 (N_21018,N_19418,N_18230);
or U21019 (N_21019,N_19165,N_19871);
nand U21020 (N_21020,N_18969,N_18541);
and U21021 (N_21021,N_20242,N_19643);
or U21022 (N_21022,N_19539,N_18924);
nand U21023 (N_21023,N_19672,N_19540);
nor U21024 (N_21024,N_18842,N_18703);
nor U21025 (N_21025,N_19934,N_18474);
and U21026 (N_21026,N_20210,N_19683);
xnor U21027 (N_21027,N_20186,N_18104);
xor U21028 (N_21028,N_20034,N_19512);
nor U21029 (N_21029,N_18343,N_20036);
xor U21030 (N_21030,N_20107,N_19107);
xnor U21031 (N_21031,N_19838,N_20161);
nand U21032 (N_21032,N_20546,N_20866);
or U21033 (N_21033,N_19823,N_19686);
and U21034 (N_21034,N_20521,N_20344);
nor U21035 (N_21035,N_18871,N_18222);
or U21036 (N_21036,N_20333,N_19119);
nand U21037 (N_21037,N_19728,N_19836);
nand U21038 (N_21038,N_20117,N_18624);
nand U21039 (N_21039,N_18143,N_18302);
xor U21040 (N_21040,N_19018,N_19324);
xnor U21041 (N_21041,N_19405,N_20744);
and U21042 (N_21042,N_20519,N_18594);
and U21043 (N_21043,N_18868,N_20135);
xor U21044 (N_21044,N_20269,N_18215);
and U21045 (N_21045,N_19981,N_20054);
xor U21046 (N_21046,N_19742,N_18423);
and U21047 (N_21047,N_20570,N_18178);
nor U21048 (N_21048,N_19373,N_19691);
or U21049 (N_21049,N_20730,N_19372);
and U21050 (N_21050,N_20804,N_18713);
nand U21051 (N_21051,N_19906,N_19759);
nand U21052 (N_21052,N_19822,N_20291);
or U21053 (N_21053,N_20737,N_18360);
nor U21054 (N_21054,N_19924,N_20162);
and U21055 (N_21055,N_19053,N_18031);
nand U21056 (N_21056,N_19003,N_19867);
nand U21057 (N_21057,N_19675,N_18151);
xor U21058 (N_21058,N_20230,N_20055);
nand U21059 (N_21059,N_19804,N_19491);
nor U21060 (N_21060,N_20900,N_20411);
nor U21061 (N_21061,N_20418,N_19073);
nor U21062 (N_21062,N_19434,N_20922);
or U21063 (N_21063,N_20000,N_20752);
or U21064 (N_21064,N_20402,N_18934);
xor U21065 (N_21065,N_19045,N_19942);
xnor U21066 (N_21066,N_18582,N_20528);
and U21067 (N_21067,N_19678,N_20393);
nand U21068 (N_21068,N_19134,N_18422);
and U21069 (N_21069,N_20791,N_18428);
or U21070 (N_21070,N_18849,N_18297);
nand U21071 (N_21071,N_18250,N_18931);
or U21072 (N_21072,N_20788,N_19515);
and U21073 (N_21073,N_18291,N_18783);
xor U21074 (N_21074,N_20822,N_20719);
or U21075 (N_21075,N_19574,N_18691);
or U21076 (N_21076,N_19627,N_18105);
nor U21077 (N_21077,N_18675,N_20207);
and U21078 (N_21078,N_20780,N_20139);
nor U21079 (N_21079,N_18885,N_18179);
or U21080 (N_21080,N_19327,N_19355);
and U21081 (N_21081,N_19211,N_18109);
nand U21082 (N_21082,N_19990,N_20094);
nand U21083 (N_21083,N_18115,N_20061);
and U21084 (N_21084,N_18470,N_20462);
nand U21085 (N_21085,N_19187,N_18910);
or U21086 (N_21086,N_20104,N_20324);
xnor U21087 (N_21087,N_18869,N_20090);
and U21088 (N_21088,N_18127,N_20338);
nor U21089 (N_21089,N_20968,N_19350);
and U21090 (N_21090,N_20314,N_20496);
nand U21091 (N_21091,N_19644,N_19098);
and U21092 (N_21092,N_19994,N_20184);
nand U21093 (N_21093,N_18636,N_19647);
and U21094 (N_21094,N_19464,N_18000);
nor U21095 (N_21095,N_20174,N_20516);
or U21096 (N_21096,N_20348,N_20657);
nand U21097 (N_21097,N_20643,N_20278);
nand U21098 (N_21098,N_19800,N_18976);
nor U21099 (N_21099,N_19341,N_19448);
or U21100 (N_21100,N_20726,N_19480);
nand U21101 (N_21101,N_20335,N_18039);
nand U21102 (N_21102,N_20739,N_18432);
or U21103 (N_21103,N_19966,N_19899);
nand U21104 (N_21104,N_20961,N_19105);
nand U21105 (N_21105,N_18158,N_19684);
nand U21106 (N_21106,N_18634,N_19305);
xnor U21107 (N_21107,N_19699,N_19783);
or U21108 (N_21108,N_18079,N_18526);
and U21109 (N_21109,N_18935,N_19905);
nor U21110 (N_21110,N_18518,N_20792);
nor U21111 (N_21111,N_20856,N_19494);
nor U21112 (N_21112,N_18872,N_18153);
and U21113 (N_21113,N_19930,N_19049);
and U21114 (N_21114,N_20538,N_19502);
or U21115 (N_21115,N_19633,N_18790);
nand U21116 (N_21116,N_18013,N_19976);
and U21117 (N_21117,N_18999,N_18183);
nor U21118 (N_21118,N_19493,N_19841);
xor U21119 (N_21119,N_19316,N_19922);
xnor U21120 (N_21120,N_18888,N_19888);
or U21121 (N_21121,N_18616,N_18765);
and U21122 (N_21122,N_19524,N_18604);
or U21123 (N_21123,N_20006,N_20023);
xnor U21124 (N_21124,N_19718,N_19342);
and U21125 (N_21125,N_19466,N_19791);
nand U21126 (N_21126,N_19777,N_20478);
and U21127 (N_21127,N_18515,N_20685);
and U21128 (N_21128,N_19664,N_18018);
nor U21129 (N_21129,N_18708,N_20800);
xor U21130 (N_21130,N_20937,N_18922);
or U21131 (N_21131,N_19848,N_20590);
nand U21132 (N_21132,N_20147,N_19220);
xor U21133 (N_21133,N_20136,N_18320);
nand U21134 (N_21134,N_18987,N_19167);
nand U21135 (N_21135,N_20965,N_18967);
xnor U21136 (N_21136,N_18226,N_18628);
or U21137 (N_21137,N_19587,N_18762);
xor U21138 (N_21138,N_18174,N_18099);
nor U21139 (N_21139,N_18895,N_18403);
xnor U21140 (N_21140,N_18417,N_18478);
and U21141 (N_21141,N_19645,N_20450);
nor U21142 (N_21142,N_20168,N_20951);
nand U21143 (N_21143,N_18346,N_20681);
or U21144 (N_21144,N_18224,N_18269);
or U21145 (N_21145,N_20383,N_19266);
xnor U21146 (N_21146,N_19843,N_19468);
or U21147 (N_21147,N_18107,N_19139);
nand U21148 (N_21148,N_20897,N_20138);
or U21149 (N_21149,N_19182,N_19757);
nand U21150 (N_21150,N_18473,N_18932);
xnor U21151 (N_21151,N_20913,N_20473);
and U21152 (N_21152,N_18248,N_20812);
and U21153 (N_21153,N_18315,N_19209);
nand U21154 (N_21154,N_19056,N_19268);
nor U21155 (N_21155,N_19065,N_18561);
and U21156 (N_21156,N_20366,N_18098);
or U21157 (N_21157,N_19965,N_20218);
nand U21158 (N_21158,N_20043,N_20245);
or U21159 (N_21159,N_18100,N_20647);
nand U21160 (N_21160,N_19485,N_18625);
or U21161 (N_21161,N_18770,N_18087);
nand U21162 (N_21162,N_18135,N_19242);
and U21163 (N_21163,N_19312,N_19743);
nand U21164 (N_21164,N_18789,N_18781);
xnor U21165 (N_21165,N_18456,N_18852);
or U21166 (N_21166,N_20573,N_18246);
and U21167 (N_21167,N_18943,N_18058);
and U21168 (N_21168,N_18394,N_19157);
nand U21169 (N_21169,N_18112,N_19668);
nand U21170 (N_21170,N_20018,N_20589);
nor U21171 (N_21171,N_19531,N_20330);
xnor U21172 (N_21172,N_18635,N_18085);
nand U21173 (N_21173,N_18319,N_19891);
xnor U21174 (N_21174,N_18968,N_19721);
xor U21175 (N_21175,N_20404,N_19293);
and U21176 (N_21176,N_19273,N_18768);
xor U21177 (N_21177,N_20003,N_19534);
xor U21178 (N_21178,N_20255,N_18181);
nand U21179 (N_21179,N_18575,N_20300);
or U21180 (N_21180,N_20196,N_18775);
xnor U21181 (N_21181,N_18114,N_18759);
or U21182 (N_21182,N_20838,N_20041);
xnor U21183 (N_21183,N_20171,N_19948);
and U21184 (N_21184,N_20631,N_18766);
or U21185 (N_21185,N_19789,N_20567);
or U21186 (N_21186,N_19185,N_19901);
and U21187 (N_21187,N_19102,N_18280);
and U21188 (N_21188,N_18535,N_18137);
nand U21189 (N_21189,N_19031,N_19690);
nor U21190 (N_21190,N_19022,N_20035);
or U21191 (N_21191,N_20881,N_20423);
xor U21192 (N_21192,N_18128,N_19160);
and U21193 (N_21193,N_18860,N_20665);
and U21194 (N_21194,N_19421,N_18384);
xnor U21195 (N_21195,N_19764,N_20518);
nand U21196 (N_21196,N_18238,N_18295);
and U21197 (N_21197,N_20994,N_20422);
nand U21198 (N_21198,N_20395,N_19663);
and U21199 (N_21199,N_20608,N_19681);
xor U21200 (N_21200,N_19436,N_19714);
and U21201 (N_21201,N_18756,N_18825);
and U21202 (N_21202,N_20845,N_18659);
xor U21203 (N_21203,N_18374,N_20776);
or U21204 (N_21204,N_19793,N_18929);
or U21205 (N_21205,N_20677,N_18711);
and U21206 (N_21206,N_18540,N_20307);
nor U21207 (N_21207,N_20007,N_19612);
nor U21208 (N_21208,N_19150,N_19632);
nor U21209 (N_21209,N_20784,N_20204);
and U21210 (N_21210,N_20306,N_18829);
nand U21211 (N_21211,N_20060,N_18672);
nand U21212 (N_21212,N_19857,N_20532);
and U21213 (N_21213,N_18267,N_19915);
and U21214 (N_21214,N_20783,N_19870);
nand U21215 (N_21215,N_19863,N_19114);
and U21216 (N_21216,N_19472,N_19925);
nand U21217 (N_21217,N_19566,N_20219);
nor U21218 (N_21218,N_20351,N_20603);
or U21219 (N_21219,N_20813,N_18828);
xnor U21220 (N_21220,N_18513,N_19259);
and U21221 (N_21221,N_20332,N_20111);
or U21222 (N_21222,N_19878,N_20952);
nor U21223 (N_21223,N_20653,N_18305);
and U21224 (N_21224,N_20001,N_20953);
xor U21225 (N_21225,N_20511,N_19460);
and U21226 (N_21226,N_20038,N_20028);
or U21227 (N_21227,N_18661,N_18089);
nor U21228 (N_21228,N_19950,N_18527);
or U21229 (N_21229,N_18771,N_18028);
and U21230 (N_21230,N_18406,N_20237);
and U21231 (N_21231,N_19855,N_20724);
or U21232 (N_21232,N_19175,N_19099);
nor U21233 (N_21233,N_20808,N_18965);
and U21234 (N_21234,N_20392,N_18680);
nor U21235 (N_21235,N_18330,N_19154);
nor U21236 (N_21236,N_18785,N_20096);
nand U21237 (N_21237,N_19991,N_19559);
nor U21238 (N_21238,N_18833,N_19737);
nor U21239 (N_21239,N_19058,N_20256);
nand U21240 (N_21240,N_18113,N_19709);
nand U21241 (N_21241,N_20806,N_18097);
nor U21242 (N_21242,N_18560,N_18637);
nor U21243 (N_21243,N_20942,N_19328);
nand U21244 (N_21244,N_19044,N_19335);
xor U21245 (N_21245,N_20249,N_19636);
or U21246 (N_21246,N_18276,N_18709);
nor U21247 (N_21247,N_19059,N_18091);
nor U21248 (N_21248,N_20901,N_18663);
xnor U21249 (N_21249,N_18697,N_20254);
nand U21250 (N_21250,N_20903,N_19600);
and U21251 (N_21251,N_20740,N_18858);
and U21252 (N_21252,N_19444,N_19348);
or U21253 (N_21253,N_18009,N_18342);
xor U21254 (N_21254,N_20440,N_18486);
or U21255 (N_21255,N_18409,N_20981);
nand U21256 (N_21256,N_19081,N_18900);
nor U21257 (N_21257,N_20695,N_20713);
and U21258 (N_21258,N_20557,N_19995);
nor U21259 (N_21259,N_18612,N_18024);
or U21260 (N_21260,N_19661,N_18679);
nor U21261 (N_21261,N_19951,N_19322);
nor U21262 (N_21262,N_20535,N_20520);
nand U21263 (N_21263,N_19523,N_20396);
or U21264 (N_21264,N_19492,N_19658);
nor U21265 (N_21265,N_18945,N_19489);
nand U21266 (N_21266,N_18283,N_20290);
nor U21267 (N_21267,N_19417,N_20830);
or U21268 (N_21268,N_18331,N_18814);
xor U21269 (N_21269,N_18500,N_20932);
and U21270 (N_21270,N_20274,N_19532);
or U21271 (N_21271,N_19998,N_20539);
and U21272 (N_21272,N_20331,N_19054);
and U21273 (N_21273,N_20293,N_18642);
nor U21274 (N_21274,N_20578,N_19295);
xnor U21275 (N_21275,N_18727,N_19459);
or U21276 (N_21276,N_20084,N_18553);
or U21277 (N_21277,N_19227,N_20257);
xnor U21278 (N_21278,N_18906,N_20052);
nand U21279 (N_21279,N_18277,N_20574);
xor U21280 (N_21280,N_18667,N_20233);
xnor U21281 (N_21281,N_20382,N_20931);
and U21282 (N_21282,N_20284,N_19551);
nand U21283 (N_21283,N_19155,N_18020);
or U21284 (N_21284,N_19307,N_20401);
xnor U21285 (N_21285,N_19475,N_18139);
and U21286 (N_21286,N_19301,N_20180);
nor U21287 (N_21287,N_18034,N_20352);
and U21288 (N_21288,N_19006,N_18673);
nor U21289 (N_21289,N_18410,N_20507);
or U21290 (N_21290,N_20599,N_20127);
nand U21291 (N_21291,N_19564,N_19428);
xnor U21292 (N_21292,N_18232,N_20093);
and U21293 (N_21293,N_20033,N_20214);
xnor U21294 (N_21294,N_18338,N_20735);
nand U21295 (N_21295,N_18348,N_18152);
nand U21296 (N_21296,N_19481,N_19488);
nand U21297 (N_21297,N_18517,N_20947);
nor U21298 (N_21298,N_20627,N_18207);
or U21299 (N_21299,N_18964,N_19581);
xor U21300 (N_21300,N_18457,N_20376);
nor U21301 (N_21301,N_18481,N_19954);
xnor U21302 (N_21302,N_19473,N_19203);
xnor U21303 (N_21303,N_19343,N_20834);
nor U21304 (N_21304,N_19550,N_19198);
and U21305 (N_21305,N_18106,N_18933);
nand U21306 (N_21306,N_18846,N_18510);
and U21307 (N_21307,N_19886,N_20849);
nor U21308 (N_21308,N_18893,N_19357);
or U21309 (N_21309,N_19774,N_18817);
xor U21310 (N_21310,N_18057,N_19613);
or U21311 (N_21311,N_20131,N_18260);
nand U21312 (N_21312,N_19110,N_18312);
or U21313 (N_21313,N_18471,N_20836);
xnor U21314 (N_21314,N_18068,N_19565);
xor U21315 (N_21315,N_19169,N_20372);
xnor U21316 (N_21316,N_19592,N_18204);
nand U21317 (N_21317,N_19898,N_18937);
nor U21318 (N_21318,N_18760,N_18608);
nor U21319 (N_21319,N_18095,N_20742);
or U21320 (N_21320,N_18040,N_19230);
or U21321 (N_21321,N_20588,N_20743);
and U21322 (N_21322,N_20621,N_18460);
nor U21323 (N_21323,N_18840,N_18060);
xnor U21324 (N_21324,N_18717,N_19958);
nand U21325 (N_21325,N_20159,N_20640);
nand U21326 (N_21326,N_20102,N_20201);
nor U21327 (N_21327,N_20341,N_19801);
nand U21328 (N_21328,N_18654,N_20078);
and U21329 (N_21329,N_20956,N_20683);
nor U21330 (N_21330,N_20424,N_19311);
and U21331 (N_21331,N_19497,N_20946);
nand U21332 (N_21332,N_19671,N_18764);
nand U21333 (N_21333,N_20945,N_18850);
nand U21334 (N_21334,N_18578,N_20364);
xor U21335 (N_21335,N_19547,N_20206);
and U21336 (N_21336,N_20173,N_18416);
nand U21337 (N_21337,N_18623,N_19255);
and U21338 (N_21338,N_19121,N_19693);
nand U21339 (N_21339,N_19153,N_18927);
and U21340 (N_21340,N_20040,N_18803);
nor U21341 (N_21341,N_18063,N_20654);
or U21342 (N_21342,N_19239,N_18281);
nand U21343 (N_21343,N_19713,N_19364);
xor U21344 (N_21344,N_20215,N_19947);
xor U21345 (N_21345,N_19556,N_18499);
xnor U21346 (N_21346,N_20438,N_20980);
or U21347 (N_21347,N_19651,N_18960);
or U21348 (N_21348,N_19496,N_20982);
nor U21349 (N_21349,N_20318,N_19811);
or U21350 (N_21350,N_18971,N_20056);
nor U21351 (N_21351,N_20772,N_19000);
or U21352 (N_21352,N_20696,N_18610);
nor U21353 (N_21353,N_18237,N_19505);
or U21354 (N_21354,N_19294,N_20809);
or U21355 (N_21355,N_18614,N_18993);
and U21356 (N_21356,N_20347,N_20187);
nand U21357 (N_21357,N_20633,N_20053);
xor U21358 (N_21358,N_20497,N_18395);
nand U21359 (N_21359,N_18630,N_20490);
xnor U21360 (N_21360,N_20228,N_20189);
nor U21361 (N_21361,N_18026,N_18718);
nor U21362 (N_21362,N_18714,N_19662);
nor U21363 (N_21363,N_20213,N_20864);
or U21364 (N_21364,N_18705,N_19750);
nand U21365 (N_21365,N_19095,N_20919);
xor U21366 (N_21366,N_18881,N_20110);
xor U21367 (N_21367,N_18073,N_20764);
or U21368 (N_21368,N_19984,N_18903);
nor U21369 (N_21369,N_19654,N_20100);
xnor U21370 (N_21370,N_19249,N_20313);
nor U21371 (N_21371,N_19563,N_19814);
and U21372 (N_21372,N_20671,N_20283);
nor U21373 (N_21373,N_18914,N_18355);
xor U21374 (N_21374,N_20465,N_18218);
and U21375 (N_21375,N_20157,N_18545);
nand U21376 (N_21376,N_18341,N_18660);
or U21377 (N_21377,N_19344,N_20770);
xnor U21378 (N_21378,N_19621,N_19927);
or U21379 (N_21379,N_18583,N_19456);
and U21380 (N_21380,N_18700,N_18195);
nor U21381 (N_21381,N_19089,N_19879);
xnor U21382 (N_21382,N_19111,N_20600);
and U21383 (N_21383,N_19264,N_20814);
or U21384 (N_21384,N_20042,N_19670);
xor U21385 (N_21385,N_20449,N_18876);
or U21386 (N_21386,N_20459,N_20680);
nor U21387 (N_21387,N_19270,N_18369);
and U21388 (N_21388,N_19725,N_18314);
nor U21389 (N_21389,N_18156,N_19688);
nand U21390 (N_21390,N_19463,N_18794);
and U21391 (N_21391,N_20560,N_18427);
nand U21392 (N_21392,N_18796,N_18658);
xor U21393 (N_21393,N_20577,N_20909);
and U21394 (N_21394,N_20581,N_19216);
xnor U21395 (N_21395,N_18581,N_19692);
or U21396 (N_21396,N_19385,N_18815);
nand U21397 (N_21397,N_20991,N_20753);
nand U21398 (N_21398,N_20381,N_18136);
nand U21399 (N_21399,N_19253,N_19964);
or U21400 (N_21400,N_20004,N_20145);
or U21401 (N_21401,N_19205,N_20360);
nor U21402 (N_21402,N_20399,N_20238);
xor U21403 (N_21403,N_19156,N_20533);
xor U21404 (N_21404,N_19201,N_20010);
xnor U21405 (N_21405,N_19116,N_18367);
xnor U21406 (N_21406,N_18150,N_18776);
nand U21407 (N_21407,N_19314,N_18546);
nand U21408 (N_21408,N_18777,N_18336);
and U21409 (N_21409,N_19824,N_20386);
xor U21410 (N_21410,N_19940,N_20527);
and U21411 (N_21411,N_18458,N_19642);
nor U21412 (N_21412,N_19383,N_18044);
xnor U21413 (N_21413,N_18002,N_19112);
xnor U21414 (N_21414,N_19507,N_18974);
nor U21415 (N_21415,N_18399,N_18755);
or U21416 (N_21416,N_20554,N_19807);
nor U21417 (N_21417,N_19286,N_19218);
nor U21418 (N_21418,N_19839,N_18884);
xnor U21419 (N_21419,N_20563,N_19263);
and U21420 (N_21420,N_18730,N_20309);
nor U21421 (N_21421,N_20350,N_19233);
or U21422 (N_21422,N_18901,N_20580);
nand U21423 (N_21423,N_18784,N_20950);
nand U21424 (N_21424,N_18596,N_18033);
and U21425 (N_21425,N_20299,N_20745);
nor U21426 (N_21426,N_18162,N_19517);
and U21427 (N_21427,N_20958,N_19889);
and U21428 (N_21428,N_18539,N_19362);
xnor U21429 (N_21429,N_20176,N_18589);
xnor U21430 (N_21430,N_18752,N_20750);
and U21431 (N_21431,N_18704,N_19988);
nand U21432 (N_21432,N_19299,N_18650);
and U21433 (N_21433,N_20941,N_19674);
xnor U21434 (N_21434,N_18602,N_19799);
nor U21435 (N_21435,N_18693,N_19103);
xnor U21436 (N_21436,N_19501,N_20893);
xnor U21437 (N_21437,N_18787,N_19461);
xor U21438 (N_21438,N_18576,N_19057);
nand U21439 (N_21439,N_20320,N_19403);
nand U21440 (N_21440,N_18306,N_18186);
nor U21441 (N_21441,N_18388,N_20166);
and U21442 (N_21442,N_20820,N_18468);
nor U21443 (N_21443,N_18140,N_20365);
or U21444 (N_21444,N_20669,N_19520);
xnor U21445 (N_21445,N_19180,N_18373);
xor U21446 (N_21446,N_18236,N_20618);
nand U21447 (N_21447,N_19197,N_20605);
or U21448 (N_21448,N_20771,N_20273);
or U21449 (N_21449,N_20039,N_19518);
xor U21450 (N_21450,N_18577,N_18822);
and U21451 (N_21451,N_18707,N_19552);
or U21452 (N_21452,N_20321,N_20667);
nand U21453 (N_21453,N_18984,N_18838);
nor U21454 (N_21454,N_18052,N_19479);
nor U21455 (N_21455,N_19407,N_18710);
nor U21456 (N_21456,N_20252,N_18287);
or U21457 (N_21457,N_18883,N_19186);
and U21458 (N_21458,N_20673,N_20623);
and U21459 (N_21459,N_19382,N_18688);
nand U21460 (N_21460,N_18078,N_19076);
and U21461 (N_21461,N_20378,N_19265);
nor U21462 (N_21462,N_20345,N_18864);
or U21463 (N_21463,N_20425,N_20996);
and U21464 (N_21464,N_18366,N_19993);
nand U21465 (N_21465,N_18598,N_18475);
nand U21466 (N_21466,N_20445,N_18379);
xnor U21467 (N_21467,N_19100,N_18414);
nor U21468 (N_21468,N_20543,N_18742);
nand U21469 (N_21469,N_20888,N_19238);
nor U21470 (N_21470,N_19177,N_18657);
nand U21471 (N_21471,N_19477,N_18670);
nand U21472 (N_21472,N_18251,N_20134);
and U21473 (N_21473,N_20629,N_18827);
and U21474 (N_21474,N_18668,N_18227);
xnor U21475 (N_21475,N_19500,N_18681);
or U21476 (N_21476,N_20485,N_19553);
or U21477 (N_21477,N_20502,N_19726);
and U21478 (N_21478,N_18368,N_18455);
and U21479 (N_21479,N_20568,N_19332);
nand U21480 (N_21480,N_20391,N_18193);
nor U21481 (N_21481,N_19088,N_18975);
xnor U21482 (N_21482,N_19237,N_19781);
and U21483 (N_21483,N_19094,N_18566);
and U21484 (N_21484,N_20799,N_18041);
xor U21485 (N_21485,N_20962,N_18122);
or U21486 (N_21486,N_18411,N_18646);
xor U21487 (N_21487,N_18365,N_18264);
nand U21488 (N_21488,N_20217,N_18599);
nand U21489 (N_21489,N_20524,N_19554);
or U21490 (N_21490,N_19427,N_19504);
nor U21491 (N_21491,N_20193,N_18726);
nand U21492 (N_21492,N_20451,N_19406);
or U21493 (N_21493,N_18439,N_19061);
nand U21494 (N_21494,N_19831,N_20178);
nand U21495 (N_21495,N_20601,N_19440);
xnor U21496 (N_21496,N_18733,N_19873);
and U21497 (N_21497,N_19845,N_18211);
nor U21498 (N_21498,N_20857,N_18645);
nor U21499 (N_21499,N_20286,N_19339);
nor U21500 (N_21500,N_20606,N_20689);
or U21501 (N_21501,N_18802,N_18160);
or U21502 (N_21502,N_19223,N_18254);
xnor U21503 (N_21503,N_20005,N_18351);
nand U21504 (N_21504,N_20656,N_20155);
and U21505 (N_21505,N_18443,N_20072);
xnor U21506 (N_21506,N_19248,N_19803);
nand U21507 (N_21507,N_19245,N_19923);
xnor U21508 (N_21508,N_20177,N_19351);
or U21509 (N_21509,N_19812,N_19439);
nor U21510 (N_21510,N_18197,N_20619);
or U21511 (N_21511,N_19377,N_20412);
and U21512 (N_21512,N_18531,N_18271);
nor U21513 (N_21513,N_19142,N_18737);
and U21514 (N_21514,N_20678,N_20182);
nand U21515 (N_21515,N_19019,N_19048);
xnor U21516 (N_21516,N_20712,N_18548);
and U21517 (N_21517,N_19835,N_18745);
nor U21518 (N_21518,N_18357,N_18205);
or U21519 (N_21519,N_18378,N_18464);
nand U21520 (N_21520,N_18669,N_18245);
and U21521 (N_21521,N_18958,N_19620);
and U21522 (N_21522,N_19345,N_20641);
nand U21523 (N_21523,N_18208,N_19068);
xor U21524 (N_21524,N_18132,N_20045);
or U21525 (N_21525,N_18461,N_20779);
nand U21526 (N_21526,N_20514,N_18744);
or U21527 (N_21527,N_20123,N_18376);
or U21528 (N_21528,N_18307,N_20662);
nor U21529 (N_21529,N_18380,N_18683);
xor U21530 (N_21530,N_20203,N_18308);
and U21531 (N_21531,N_19118,N_20759);
or U21532 (N_21532,N_18699,N_19676);
nand U21533 (N_21533,N_20684,N_18549);
nor U21534 (N_21534,N_19949,N_20655);
or U21535 (N_21535,N_18743,N_18223);
nor U21536 (N_21536,N_20595,N_20954);
nand U21537 (N_21537,N_19008,N_20966);
nor U21538 (N_21538,N_19618,N_18413);
nor U21539 (N_21539,N_18167,N_19132);
nor U21540 (N_21540,N_20421,N_19956);
or U21541 (N_21541,N_20855,N_20216);
or U21542 (N_21542,N_20013,N_20510);
or U21543 (N_21543,N_18234,N_20691);
or U21544 (N_21544,N_18096,N_18495);
and U21545 (N_21545,N_18956,N_20637);
and U21546 (N_21546,N_20796,N_18133);
or U21547 (N_21547,N_20085,N_20340);
xnor U21548 (N_21548,N_20463,N_20879);
nor U21549 (N_21549,N_19128,N_18029);
nand U21550 (N_21550,N_18911,N_20969);
and U21551 (N_21551,N_19166,N_18559);
xor U21552 (N_21552,N_19404,N_19413);
and U21553 (N_21553,N_20815,N_19247);
nand U21554 (N_21554,N_18289,N_18279);
xnor U21555 (N_21555,N_18217,N_20871);
xnor U21556 (N_21556,N_19340,N_20342);
nor U21557 (N_21557,N_18448,N_18278);
nor U21558 (N_21558,N_20470,N_19787);
nand U21559 (N_21559,N_19711,N_18919);
and U21560 (N_21560,N_19583,N_19920);
xor U21561 (N_21561,N_18192,N_20569);
or U21562 (N_21562,N_19623,N_19611);
xnor U21563 (N_21563,N_19082,N_20661);
or U21564 (N_21564,N_18061,N_18607);
xnor U21565 (N_21565,N_19744,N_19267);
or U21566 (N_21566,N_20160,N_18619);
xnor U21567 (N_21567,N_20068,N_19738);
and U21568 (N_21568,N_18339,N_20868);
or U21569 (N_21569,N_18818,N_20995);
and U21570 (N_21570,N_19776,N_18905);
nor U21571 (N_21571,N_18022,N_18731);
nand U21572 (N_21572,N_20363,N_19359);
nor U21573 (N_21573,N_20530,N_20448);
xnor U21574 (N_21574,N_18467,N_19893);
nor U21575 (N_21575,N_19970,N_18989);
nor U21576 (N_21576,N_18169,N_19607);
nand U21577 (N_21577,N_20862,N_18902);
nand U21578 (N_21578,N_20754,N_20622);
xnor U21579 (N_21579,N_20870,N_19578);
xor U21580 (N_21580,N_20592,N_18580);
nand U21581 (N_21581,N_18426,N_18450);
nor U21582 (N_21582,N_18212,N_19084);
nor U21583 (N_21583,N_20016,N_20547);
and U21584 (N_21584,N_19590,N_20628);
nand U21585 (N_21585,N_18520,N_18484);
nand U21586 (N_21586,N_19458,N_19816);
xnor U21587 (N_21587,N_20361,N_20063);
or U21588 (N_21588,N_18980,N_19689);
xnor U21589 (N_21589,N_19615,N_18750);
nand U21590 (N_21590,N_18389,N_20636);
nand U21591 (N_21591,N_19036,N_20062);
xnor U21592 (N_21592,N_20234,N_18149);
xnor U21593 (N_21593,N_19561,N_20679);
nor U21594 (N_21594,N_19859,N_18142);
and U21595 (N_21595,N_18506,N_18102);
or U21596 (N_21596,N_18532,N_19589);
xor U21597 (N_21597,N_18472,N_18719);
nor U21598 (N_21598,N_20634,N_20832);
nand U21599 (N_21599,N_18265,N_18735);
xor U21600 (N_21600,N_19025,N_18209);
nand U21601 (N_21601,N_20190,N_20587);
nor U21602 (N_21602,N_18154,N_19637);
xor U21603 (N_21603,N_20140,N_19055);
nor U21604 (N_21604,N_20874,N_20339);
xor U21605 (N_21605,N_18509,N_18228);
and U21606 (N_21606,N_20048,N_20329);
nand U21607 (N_21607,N_20141,N_19224);
or U21608 (N_21608,N_18401,N_18335);
nand U21609 (N_21609,N_18266,N_18333);
nand U21610 (N_21610,N_18042,N_19030);
nand U21611 (N_21611,N_19462,N_18702);
nand U21612 (N_21612,N_19775,N_20706);
xor U21613 (N_21613,N_18497,N_20370);
xor U21614 (N_21614,N_19960,N_19624);
nor U21615 (N_21615,N_20070,N_20786);
nand U21616 (N_21616,N_18847,N_20872);
and U21617 (N_21617,N_18844,N_18004);
or U21618 (N_21618,N_20967,N_18072);
xnor U21619 (N_21619,N_19544,N_19309);
xnor U21620 (N_21620,N_20688,N_19109);
nand U21621 (N_21621,N_19967,N_18168);
nor U21622 (N_21622,N_18334,N_18763);
nor U21623 (N_21623,N_20073,N_20829);
or U21624 (N_21624,N_19963,N_20513);
or U21625 (N_21625,N_19199,N_18898);
xor U21626 (N_21626,N_20846,N_18452);
or U21627 (N_21627,N_20151,N_20727);
and U21628 (N_21628,N_20443,N_18948);
nand U21629 (N_21629,N_19447,N_19570);
nand U21630 (N_21630,N_19290,N_20263);
nand U21631 (N_21631,N_20091,N_20992);
nor U21632 (N_21632,N_19035,N_19526);
and U21633 (N_21633,N_20807,N_19833);
nor U21634 (N_21634,N_18979,N_18897);
xor U21635 (N_21635,N_19370,N_18715);
xnor U21636 (N_21636,N_19120,N_20852);
or U21637 (N_21637,N_19399,N_19616);
xor U21638 (N_21638,N_18084,N_19549);
nor U21639 (N_21639,N_20672,N_19817);
or U21640 (N_21640,N_19179,N_19827);
or U21641 (N_21641,N_20801,N_20660);
nand U21642 (N_21642,N_18120,N_18587);
nand U21643 (N_21643,N_20191,N_20700);
nor U21644 (N_21644,N_18134,N_18954);
and U21645 (N_21645,N_19715,N_20185);
and U21646 (N_21646,N_18615,N_20202);
xor U21647 (N_21647,N_20358,N_19028);
nor U21648 (N_21648,N_18214,N_19173);
xor U21649 (N_21649,N_20997,N_19007);
or U21650 (N_21650,N_20398,N_20781);
nand U21651 (N_21651,N_18332,N_20506);
nand U21652 (N_21652,N_20928,N_18550);
nor U21653 (N_21653,N_18773,N_18723);
or U21654 (N_21654,N_19024,N_20489);
or U21655 (N_21655,N_18356,N_19498);
nor U21656 (N_21656,N_20782,N_20955);
or U21657 (N_21657,N_19584,N_20480);
nand U21658 (N_21658,N_19897,N_20702);
nor U21659 (N_21659,N_18397,N_19412);
xnor U21660 (N_21660,N_19535,N_20725);
xnor U21661 (N_21661,N_18621,N_19779);
or U21662 (N_21662,N_20927,N_20988);
nor U21663 (N_21663,N_19108,N_20295);
and U21664 (N_21664,N_19703,N_18555);
xor U21665 (N_21665,N_19246,N_19435);
or U21666 (N_21666,N_20549,N_20156);
and U21667 (N_21667,N_19337,N_20406);
nor U21668 (N_21668,N_20632,N_19389);
xor U21669 (N_21669,N_20272,N_18469);
nand U21670 (N_21670,N_18075,N_18164);
or U21671 (N_21671,N_18065,N_20987);
nand U21672 (N_21672,N_18070,N_19281);
nand U21673 (N_21673,N_18597,N_20328);
xnor U21674 (N_21674,N_18125,N_18400);
nor U21675 (N_21675,N_19652,N_18483);
xor U21676 (N_21676,N_20802,N_19411);
nor U21677 (N_21677,N_20359,N_18476);
and U21678 (N_21678,N_19918,N_19017);
nor U21679 (N_21679,N_20940,N_19336);
xnor U21680 (N_21680,N_19176,N_19484);
nand U21681 (N_21681,N_20758,N_20790);
nand U21682 (N_21682,N_18552,N_20163);
nor U21683 (N_21683,N_19241,N_19381);
or U21684 (N_21684,N_18285,N_19908);
and U21685 (N_21685,N_20747,N_19288);
or U21686 (N_21686,N_19868,N_18255);
nor U21687 (N_21687,N_19768,N_20024);
xnor U21688 (N_21688,N_20389,N_19020);
or U21689 (N_21689,N_19731,N_18558);
xor U21690 (N_21690,N_18835,N_19409);
xnor U21691 (N_21691,N_19014,N_18130);
nor U21692 (N_21692,N_19269,N_19666);
or U21693 (N_21693,N_18244,N_18522);
nor U21694 (N_21694,N_20316,N_18465);
xor U21695 (N_21695,N_20097,N_20429);
or U21696 (N_21696,N_19215,N_20251);
or U21697 (N_21697,N_19935,N_18321);
or U21698 (N_21698,N_20116,N_18877);
or U21699 (N_21699,N_20394,N_18706);
or U21700 (N_21700,N_18119,N_20736);
nand U21701 (N_21701,N_20793,N_18508);
and U21702 (N_21702,N_18118,N_19834);
or U21703 (N_21703,N_20477,N_19852);
nand U21704 (N_21704,N_18912,N_20923);
or U21705 (N_21705,N_19883,N_19712);
xnor U21706 (N_21706,N_19946,N_20491);
nor U21707 (N_21707,N_18916,N_18865);
and U21708 (N_21708,N_20275,N_20686);
nor U21709 (N_21709,N_19810,N_19358);
or U21710 (N_21710,N_18605,N_18689);
and U21711 (N_21711,N_20128,N_19384);
nand U21712 (N_21712,N_20575,N_20974);
nor U21713 (N_21713,N_18219,N_18011);
nand U21714 (N_21714,N_19503,N_20211);
or U21715 (N_21715,N_20624,N_20762);
and U21716 (N_21716,N_19773,N_20529);
nand U21717 (N_21717,N_20310,N_20277);
nand U21718 (N_21718,N_19387,N_18891);
nor U21719 (N_21719,N_18323,N_19786);
nand U21720 (N_21720,N_18565,N_18653);
or U21721 (N_21721,N_19232,N_20419);
xnor U21722 (N_21722,N_20247,N_19568);
xnor U21723 (N_21723,N_19980,N_20058);
or U21724 (N_21724,N_20933,N_18622);
xnor U21725 (N_21725,N_18839,N_19979);
nand U21726 (N_21726,N_19455,N_20646);
and U21727 (N_21727,N_18631,N_18145);
and U21728 (N_21728,N_19329,N_18564);
nand U21729 (N_21729,N_19213,N_18603);
and U21730 (N_21730,N_20690,N_20617);
nor U21731 (N_21731,N_20756,N_18344);
and U21732 (N_21732,N_20902,N_20734);
and U21733 (N_21733,N_18233,N_20875);
or U21734 (N_21734,N_18110,N_19722);
nor U21735 (N_21735,N_18595,N_20551);
nor U21736 (N_21736,N_18649,N_20960);
nand U21737 (N_21737,N_20586,N_19697);
or U21738 (N_21738,N_20464,N_18257);
xnor U21739 (N_21739,N_20224,N_19530);
nor U21740 (N_21740,N_18562,N_20397);
or U21741 (N_21741,N_20512,N_19441);
nand U21742 (N_21742,N_19365,N_20281);
nand U21743 (N_21743,N_18874,N_20541);
nand U21744 (N_21744,N_19609,N_20271);
xnor U21745 (N_21745,N_20778,N_19890);
nand U21746 (N_21746,N_19298,N_18198);
xnor U21747 (N_21747,N_20417,N_20635);
nor U21748 (N_21748,N_18200,N_20741);
nor U21749 (N_21749,N_18925,N_18479);
nor U21750 (N_21750,N_19667,N_19476);
nor U21751 (N_21751,N_18957,N_18358);
xor U21752 (N_21752,N_19346,N_20287);
or U21753 (N_21753,N_18729,N_18003);
and U21754 (N_21754,N_19283,N_18652);
nor U21755 (N_21755,N_20508,N_20357);
xnor U21756 (N_21756,N_20086,N_19596);
xor U21757 (N_21757,N_18438,N_18161);
and U21758 (N_21758,N_18951,N_19442);
xor U21759 (N_21759,N_19593,N_18570);
or U21760 (N_21760,N_20118,N_18686);
and U21761 (N_21761,N_18116,N_18025);
or U21762 (N_21762,N_20659,N_19303);
nor U21763 (N_21763,N_18793,N_20325);
nand U21764 (N_21764,N_20892,N_20031);
nor U21765 (N_21765,N_18080,N_18243);
xor U21766 (N_21766,N_20387,N_19158);
and U21767 (N_21767,N_18048,N_19657);
nand U21768 (N_21768,N_18391,N_19041);
nand U21769 (N_21769,N_19582,N_20917);
and U21770 (N_21770,N_20326,N_18676);
nand U21771 (N_21771,N_20971,N_20356);
nand U21772 (N_21772,N_18801,N_19957);
nand U21773 (N_21773,N_20693,N_20707);
xnor U21774 (N_21774,N_20373,N_18482);
or U21775 (N_21775,N_19914,N_18985);
and U21776 (N_21776,N_19577,N_18890);
or U21777 (N_21777,N_19136,N_19163);
or U21778 (N_21778,N_20323,N_20797);
nand U21779 (N_21779,N_20795,N_19354);
and U21780 (N_21780,N_20092,N_19528);
or U21781 (N_21781,N_20522,N_18894);
nand U21782 (N_21782,N_20146,N_18936);
xor U21783 (N_21783,N_19453,N_20584);
and U21784 (N_21784,N_19653,N_18682);
and U21785 (N_21785,N_20721,N_19603);
or U21786 (N_21786,N_18447,N_19083);
xor U21787 (N_21787,N_19770,N_19751);
and U21788 (N_21788,N_19471,N_20501);
nor U21789 (N_21789,N_19221,N_18007);
xor U21790 (N_21790,N_19602,N_19510);
nor U21791 (N_21791,N_18284,N_19302);
nand U21792 (N_21792,N_20843,N_20863);
or U21793 (N_21793,N_20983,N_18496);
and U21794 (N_21794,N_20929,N_19009);
and U21795 (N_21795,N_20239,N_19291);
and U21796 (N_21796,N_20261,N_20167);
and U21797 (N_21797,N_20088,N_18641);
xnor U21798 (N_21798,N_18311,N_19797);
or U21799 (N_21799,N_19277,N_20349);
and U21800 (N_21800,N_19075,N_19431);
nor U21801 (N_21801,N_20354,N_19195);
and U21802 (N_21802,N_19425,N_20265);
xor U21803 (N_21803,N_18083,N_19723);
xnor U21804 (N_21804,N_20500,N_18804);
nand U21805 (N_21805,N_18326,N_19569);
nand U21806 (N_21806,N_20427,N_19646);
nor U21807 (N_21807,N_18309,N_20414);
and U21808 (N_21808,N_20761,N_20375);
and U21809 (N_21809,N_20037,N_20833);
nand U21810 (N_21810,N_20243,N_20704);
or U21811 (N_21811,N_19474,N_20095);
or U21812 (N_21812,N_19204,N_18375);
nor U21813 (N_21813,N_18767,N_19380);
nand U21814 (N_21814,N_18449,N_19499);
nand U21815 (N_21815,N_18878,N_18677);
and U21816 (N_21816,N_20851,N_19509);
xor U21817 (N_21817,N_19070,N_18889);
nand U21818 (N_21818,N_20415,N_19698);
nand U21819 (N_21819,N_18998,N_18887);
or U21820 (N_21820,N_20842,N_19467);
and U21821 (N_21821,N_18203,N_19334);
and U21822 (N_21822,N_19219,N_18296);
xor U21823 (N_21823,N_20405,N_19240);
or U21824 (N_21824,N_18830,N_19933);
xor U21825 (N_21825,N_19426,N_19402);
nand U21826 (N_21826,N_19125,N_18728);
nand U21827 (N_21827,N_20602,N_20755);
or U21828 (N_21828,N_20630,N_20509);
xor U21829 (N_21829,N_20183,N_18908);
nand U21830 (N_21830,N_18944,N_19673);
nor U21831 (N_21831,N_20936,N_18834);
nand U21832 (N_21832,N_19911,N_20400);
xor U21833 (N_21833,N_19588,N_18997);
xnor U21834 (N_21834,N_19973,N_19060);
nand U21835 (N_21835,N_18175,N_19808);
xor U21836 (N_21836,N_19063,N_20195);
or U21837 (N_21837,N_19282,N_19830);
nor U21838 (N_21838,N_19236,N_18524);
nand U21839 (N_21839,N_19753,N_19541);
xnor U21840 (N_21840,N_18947,N_18533);
and U21841 (N_21841,N_19696,N_19256);
and U21842 (N_21842,N_19597,N_18592);
or U21843 (N_21843,N_19091,N_19244);
xnor U21844 (N_21844,N_19622,N_18940);
or U21845 (N_21845,N_18480,N_20390);
nor U21846 (N_21846,N_18970,N_20545);
xnor U21847 (N_21847,N_20749,N_18798);
or U21848 (N_21848,N_20260,N_19630);
or U21849 (N_21849,N_18288,N_20886);
or U21850 (N_21850,N_18514,N_19206);
or U21851 (N_21851,N_20819,N_18955);
nor U21852 (N_21852,N_18074,N_18370);
and U21853 (N_21853,N_19716,N_19913);
and U21854 (N_21854,N_20768,N_18441);
xor U21855 (N_21855,N_20235,N_20479);
nor U21856 (N_21856,N_19739,N_18551);
and U21857 (N_21857,N_18340,N_19416);
nor U21858 (N_21858,N_20082,N_19130);
or U21859 (N_21859,N_19276,N_19319);
and U21860 (N_21860,N_19331,N_19975);
and U21861 (N_21861,N_20825,N_19727);
nor U21862 (N_21862,N_19780,N_19961);
nand U21863 (N_21863,N_19939,N_18364);
nor U21864 (N_21864,N_19164,N_20668);
and U21865 (N_21865,N_20371,N_20517);
nand U21866 (N_21866,N_20246,N_19992);
xor U21867 (N_21867,N_19010,N_19420);
nor U21868 (N_21868,N_19608,N_18994);
or U21869 (N_21869,N_19884,N_19047);
and U21870 (N_21870,N_20841,N_19746);
xor U21871 (N_21871,N_19250,N_20908);
or U21872 (N_21872,N_20259,N_19971);
nand U21873 (N_21873,N_20663,N_20098);
xor U21874 (N_21874,N_19379,N_20250);
and U21875 (N_21875,N_19430,N_20847);
nand U21876 (N_21876,N_20978,N_19135);
or U21877 (N_21877,N_19141,N_19656);
nor U21878 (N_21878,N_19605,N_20074);
xnor U21879 (N_21879,N_19598,N_18725);
xnor U21880 (N_21880,N_19837,N_20883);
or U21881 (N_21881,N_20565,N_20080);
nor U21882 (N_21882,N_19601,N_20626);
nor U21883 (N_21883,N_18310,N_20150);
nand U21884 (N_21884,N_20555,N_18059);
nand U21885 (N_21885,N_19483,N_20152);
xnor U21886 (N_21886,N_20709,N_20108);
or U21887 (N_21887,N_20081,N_19599);
nand U21888 (N_21888,N_19080,N_18904);
xnor U21889 (N_21889,N_20826,N_19854);
nor U21890 (N_21890,N_20047,N_20562);
nand U21891 (N_21891,N_19944,N_19853);
or U21892 (N_21892,N_19685,N_20698);
nor U21893 (N_21893,N_19959,N_19926);
and U21894 (N_21894,N_19796,N_20194);
nor U21895 (N_21895,N_20317,N_19555);
and U21896 (N_21896,N_19638,N_19395);
or U21897 (N_21897,N_19192,N_19178);
nand U21898 (N_21898,N_19451,N_19758);
xor U21899 (N_21899,N_20311,N_19129);
xnor U21900 (N_21900,N_18644,N_18511);
nor U21901 (N_21901,N_20803,N_19506);
nand U21902 (N_21902,N_20612,N_18050);
nand U21903 (N_21903,N_18090,N_20484);
and U21904 (N_21904,N_20276,N_18820);
and U21905 (N_21905,N_20935,N_18431);
or U21906 (N_21906,N_20089,N_19754);
nor U21907 (N_21907,N_19184,N_18453);
xnor U21908 (N_21908,N_19034,N_20885);
nor U21909 (N_21909,N_19378,N_19752);
or U21910 (N_21910,N_19490,N_18189);
or U21911 (N_21911,N_18574,N_20926);
nand U21912 (N_21912,N_18617,N_19604);
nor U21913 (N_21913,N_20650,N_18579);
nand U21914 (N_21914,N_19985,N_19191);
or U21915 (N_21915,N_20760,N_19631);
xor U21916 (N_21916,N_20452,N_18361);
xor U21917 (N_21917,N_19026,N_19027);
nor U21918 (N_21918,N_20718,N_18507);
xor U21919 (N_21919,N_18247,N_19272);
nor U21920 (N_21920,N_19542,N_20288);
xor U21921 (N_21921,N_20487,N_19806);
nor U21922 (N_21922,N_19122,N_18299);
nand U21923 (N_21923,N_18505,N_20482);
or U21924 (N_21924,N_18377,N_20610);
and U21925 (N_21925,N_20876,N_19519);
nand U21926 (N_21926,N_19194,N_19228);
or U21927 (N_21927,N_19996,N_19320);
or U21928 (N_21928,N_19469,N_20687);
nand U21929 (N_21929,N_20441,N_19306);
and U21930 (N_21930,N_18585,N_19736);
or U21931 (N_21931,N_19614,N_20583);
or U21932 (N_21932,N_18444,N_18371);
and U21933 (N_21933,N_20993,N_18381);
or U21934 (N_21934,N_19977,N_19625);
or U21935 (N_21935,N_19819,N_18241);
nor U21936 (N_21936,N_18690,N_18722);
or U21937 (N_21937,N_18108,N_18536);
or U21938 (N_21938,N_19410,N_19900);
nand U21939 (N_21939,N_20944,N_20165);
nand U21940 (N_21940,N_18952,N_18235);
xnor U21941 (N_21941,N_19077,N_19087);
and U21942 (N_21942,N_20645,N_18035);
xnor U21943 (N_21943,N_18808,N_18030);
and U21944 (N_21944,N_18253,N_18813);
xnor U21945 (N_21945,N_20294,N_20212);
and U21946 (N_21946,N_19321,N_20231);
nand U21947 (N_21947,N_18404,N_18632);
xnor U21948 (N_21948,N_19821,N_18301);
or U21949 (N_21949,N_18220,N_19210);
and U21950 (N_21950,N_18316,N_18913);
or U21951 (N_21951,N_20920,N_18907);
nor U21952 (N_21952,N_18662,N_20817);
and U21953 (N_21953,N_20867,N_18221);
and U21954 (N_21954,N_20552,N_20337);
or U21955 (N_21955,N_18494,N_19315);
nor U21956 (N_21956,N_18942,N_18950);
or U21957 (N_21957,N_19529,N_20262);
and U21958 (N_21958,N_19585,N_18807);
nor U21959 (N_21959,N_19482,N_20732);
xnor U21960 (N_21960,N_18797,N_19892);
nor U21961 (N_21961,N_19756,N_19846);
or U21962 (N_21962,N_19200,N_18067);
and U21963 (N_21963,N_19767,N_20322);
nand U21964 (N_21964,N_20850,N_18268);
and U21965 (N_21965,N_18799,N_18487);
xnor U21966 (N_21966,N_19700,N_19766);
nand U21967 (N_21967,N_18103,N_18946);
or U21968 (N_21968,N_20553,N_18586);
and U21969 (N_21969,N_20525,N_19702);
nor U21970 (N_21970,N_18651,N_18436);
and U21971 (N_21971,N_19361,N_20604);
or U21972 (N_21972,N_18148,N_19818);
and U21973 (N_21973,N_19470,N_19978);
nand U21974 (N_21974,N_20523,N_18385);
nor U21975 (N_21975,N_20766,N_20505);
nor U21976 (N_21976,N_19669,N_19424);
and U21977 (N_21977,N_18537,N_20019);
or U21978 (N_21978,N_19987,N_18678);
xor U21979 (N_21979,N_20658,N_18538);
nand U21980 (N_21980,N_20544,N_19038);
and U21981 (N_21981,N_20699,N_19749);
nand U21982 (N_21982,N_18210,N_20670);
nand U21983 (N_21983,N_19659,N_19513);
or U21984 (N_21984,N_20142,N_18173);
xor U21985 (N_21985,N_20076,N_19349);
xor U21986 (N_21986,N_20458,N_18837);
or U21987 (N_21987,N_19353,N_19895);
and U21988 (N_21988,N_20763,N_20986);
xor U21989 (N_21989,N_20158,N_19310);
or U21990 (N_21990,N_20308,N_19423);
or U21991 (N_21991,N_19308,N_18015);
or U21992 (N_21992,N_18854,N_20369);
or U21993 (N_21993,N_19015,N_19050);
and U21994 (N_21994,N_19536,N_20327);
or U21995 (N_21995,N_19318,N_20079);
nor U21996 (N_21996,N_20436,N_18938);
nor U21997 (N_21997,N_18758,N_19708);
and U21998 (N_21998,N_20964,N_18081);
or U21999 (N_21999,N_19401,N_18037);
nor U22000 (N_22000,N_19606,N_19573);
or U22001 (N_22001,N_20409,N_18800);
and U22002 (N_22002,N_18146,N_20453);
xor U22003 (N_22003,N_18258,N_18093);
nand U22004 (N_22004,N_20241,N_18462);
nand U22005 (N_22005,N_18180,N_20651);
and U22006 (N_22006,N_20434,N_20949);
xor U22007 (N_22007,N_18856,N_18463);
or U22008 (N_22008,N_19649,N_19188);
or U22009 (N_22009,N_18692,N_19937);
and U22010 (N_22010,N_20859,N_18412);
xnor U22011 (N_22011,N_18440,N_18433);
xor U22012 (N_22012,N_20426,N_19792);
and U22013 (N_22013,N_18643,N_19078);
nor U22014 (N_22014,N_20708,N_19907);
nor U22015 (N_22015,N_18392,N_18202);
nor U22016 (N_22016,N_19557,N_20542);
xnor U22017 (N_22017,N_19366,N_19280);
xor U22018 (N_22018,N_20765,N_18256);
or U22019 (N_22019,N_19478,N_18736);
and U22020 (N_22020,N_19013,N_20248);
nand U22021 (N_22021,N_20703,N_20336);
and U22022 (N_22022,N_20591,N_19815);
xor U22023 (N_22023,N_19079,N_19085);
or U22024 (N_22024,N_18014,N_20878);
xnor U22025 (N_22025,N_18272,N_20420);
nand U22026 (N_22026,N_18982,N_18655);
nand U22027 (N_22027,N_20891,N_19682);
nor U22028 (N_22028,N_19287,N_20540);
or U22029 (N_22029,N_18270,N_19858);
xnor U22030 (N_22030,N_19147,N_20015);
nand U22031 (N_22031,N_20374,N_18191);
xnor U22032 (N_22032,N_19989,N_20298);
and U22033 (N_22033,N_18345,N_20697);
or U22034 (N_22034,N_18086,N_18290);
or U22035 (N_22035,N_20648,N_19955);
and U22036 (N_22036,N_18263,N_18973);
and U22037 (N_22037,N_19680,N_19046);
nand U22038 (N_22038,N_18861,N_18806);
nor U22039 (N_22039,N_19002,N_18196);
and U22040 (N_22040,N_18261,N_20112);
xnor U22041 (N_22041,N_19813,N_20748);
nand U22042 (N_22042,N_20877,N_18991);
nand U22043 (N_22043,N_19847,N_18390);
and U22044 (N_22044,N_19861,N_19798);
nand U22045 (N_22045,N_18961,N_20977);
or U22046 (N_22046,N_18821,N_18523);
nor U22047 (N_22047,N_19919,N_19093);
nor U22048 (N_22048,N_20083,N_19760);
nand U22049 (N_22049,N_20714,N_20410);
nor U22050 (N_22050,N_19445,N_18292);
and U22051 (N_22051,N_19398,N_19325);
or U22052 (N_22052,N_20620,N_19183);
and U22053 (N_22053,N_20664,N_19145);
or U22054 (N_22054,N_18337,N_18918);
xnor U22055 (N_22055,N_18780,N_20355);
xnor U22056 (N_22056,N_18021,N_19149);
nand U22057 (N_22057,N_20611,N_19575);
xnor U22058 (N_22058,N_20021,N_19734);
and U22059 (N_22059,N_18190,N_19012);
nand U22060 (N_22060,N_18049,N_20934);
or U22061 (N_22061,N_19665,N_18749);
and U22062 (N_22062,N_20811,N_18322);
xor U22063 (N_22063,N_20566,N_18584);
or U22064 (N_22064,N_19866,N_20865);
xor U22065 (N_22065,N_20649,N_18056);
and U22066 (N_22066,N_20075,N_20733);
nor U22067 (N_22067,N_20188,N_20973);
xor U22068 (N_22068,N_18571,N_20431);
and U22069 (N_22069,N_18353,N_19785);
nor U22070 (N_22070,N_20773,N_19152);
and U22071 (N_22071,N_20895,N_18147);
xor U22072 (N_22072,N_18853,N_19548);
nor U22073 (N_22073,N_20615,N_20492);
xor U22074 (N_22074,N_20362,N_20236);
nor U22075 (N_22075,N_20564,N_20114);
nor U22076 (N_22076,N_18327,N_20467);
xnor U22077 (N_22077,N_18405,N_18684);
nand U22078 (N_22078,N_18859,N_19104);
or U22079 (N_22079,N_18324,N_20924);
or U22080 (N_22080,N_18064,N_19521);
nand U22081 (N_22081,N_19454,N_19243);
or U22082 (N_22082,N_20896,N_18826);
or U22083 (N_22083,N_19001,N_18501);
or U22084 (N_22084,N_19229,N_19772);
or U22085 (N_22085,N_20515,N_20717);
nand U22086 (N_22086,N_19394,N_19097);
nor U22087 (N_22087,N_20585,N_19560);
and U22088 (N_22088,N_18023,N_20738);
and U22089 (N_22089,N_18359,N_19096);
and U22090 (N_22090,N_20794,N_18701);
nand U22091 (N_22091,N_18836,N_20258);
nor U22092 (N_22092,N_20122,N_19452);
or U22093 (N_22093,N_18131,N_19375);
nor U22094 (N_22094,N_19525,N_19591);
nand U22095 (N_22095,N_20379,N_20244);
xnor U22096 (N_22096,N_18300,N_20077);
and U22097 (N_22097,N_20025,N_18556);
xnor U22098 (N_22098,N_18362,N_18396);
and U22099 (N_22099,N_18926,N_19062);
or U22100 (N_22100,N_18863,N_18712);
nand U22101 (N_22101,N_19909,N_20169);
xor U22102 (N_22102,N_19885,N_18382);
or U22103 (N_22103,N_18185,N_18638);
nor U22104 (N_22104,N_19449,N_20915);
nor U22105 (N_22105,N_18117,N_20268);
nor U22106 (N_22106,N_19391,N_19217);
and U22107 (N_22107,N_19131,N_20172);
or U22108 (N_22108,N_19032,N_20472);
xnor U22109 (N_22109,N_19856,N_18988);
or U22110 (N_22110,N_20906,N_19392);
and U22111 (N_22111,N_20343,N_20179);
nor U22112 (N_22112,N_19172,N_20613);
and U22113 (N_22113,N_20488,N_20388);
nand U22114 (N_22114,N_20011,N_19896);
nand U22115 (N_22115,N_18995,N_19072);
nand U22116 (N_22116,N_19881,N_19457);
nor U22117 (N_22117,N_19733,N_18274);
nor U22118 (N_22118,N_20002,N_18788);
xor U22119 (N_22119,N_18303,N_18779);
xnor U22120 (N_22120,N_20442,N_20976);
nand U22121 (N_22121,N_18038,N_18990);
nand U22122 (N_22122,N_19313,N_18054);
nor U22123 (N_22123,N_18996,N_20990);
nor U22124 (N_22124,N_18062,N_20380);
nand U22125 (N_22125,N_19408,N_20894);
or U22126 (N_22126,N_19586,N_19275);
nor U22127 (N_22127,N_19437,N_19865);
nand U22128 (N_22128,N_20124,N_19212);
nand U22129 (N_22129,N_20625,N_19261);
xor U22130 (N_22130,N_18855,N_18528);
and U22131 (N_22131,N_19300,N_19052);
and U22132 (N_22132,N_20192,N_18963);
and U22133 (N_22133,N_20346,N_20066);
xor U22134 (N_22134,N_18188,N_20598);
nand U22135 (N_22135,N_18786,N_19805);
xor U22136 (N_22136,N_18187,N_18812);
xnor U22137 (N_22137,N_19655,N_18347);
xnor U22138 (N_22138,N_18857,N_20582);
or U22139 (N_22139,N_19903,N_20884);
nand U22140 (N_22140,N_20493,N_20805);
nand U22141 (N_22141,N_20270,N_19360);
nand U22142 (N_22142,N_18421,N_19634);
and U22143 (N_22143,N_18870,N_18239);
xor U22144 (N_22144,N_19226,N_19487);
or U22145 (N_22145,N_18170,N_18986);
nand U22146 (N_22146,N_19872,N_20130);
or U22147 (N_22147,N_20609,N_20898);
xnor U22148 (N_22148,N_19214,N_18298);
xor U22149 (N_22149,N_19067,N_19710);
xor U22150 (N_22150,N_18393,N_19572);
nand U22151 (N_22151,N_19438,N_19887);
or U22152 (N_22152,N_20844,N_19626);
and U22153 (N_22153,N_20115,N_20989);
nand U22154 (N_22154,N_20821,N_18121);
nor U22155 (N_22155,N_18489,N_18354);
or U22156 (N_22156,N_20057,N_20312);
and U22157 (N_22157,N_18408,N_20715);
nor U22158 (N_22158,N_18696,N_20860);
xnor U22159 (N_22159,N_18892,N_20106);
xnor U22160 (N_22160,N_19033,N_20938);
xor U22161 (N_22161,N_19231,N_18418);
nand U22162 (N_22162,N_19021,N_20787);
xor U22163 (N_22163,N_18734,N_18866);
and U22164 (N_22164,N_20014,N_20692);
nand U22165 (N_22165,N_19415,N_18809);
and U22166 (N_22166,N_18547,N_18155);
nor U22167 (N_22167,N_19687,N_18092);
and U22168 (N_22168,N_20416,N_20385);
and U22169 (N_22169,N_19579,N_20682);
nand U22170 (N_22170,N_19326,N_20918);
and U22171 (N_22171,N_19745,N_19124);
nor U22172 (N_22172,N_18590,N_20593);
nand U22173 (N_22173,N_19862,N_18446);
nor U22174 (N_22174,N_18512,N_20432);
nand U22175 (N_22175,N_20644,N_19842);
and U22176 (N_22176,N_18262,N_18259);
and U22177 (N_22177,N_20460,N_20858);
nor U22178 (N_22178,N_18053,N_18611);
xnor U22179 (N_22179,N_19388,N_19755);
xor U22180 (N_22180,N_20899,N_20720);
and U22181 (N_22181,N_18101,N_18782);
xor U22182 (N_22182,N_19279,N_18754);
and U22183 (N_22183,N_18516,N_20889);
or U22184 (N_22184,N_19802,N_20304);
or U22185 (N_22185,N_20132,N_18313);
nor U22186 (N_22186,N_20597,N_20407);
nand U22187 (N_22187,N_20498,N_19297);
nor U22188 (N_22188,N_19514,N_18419);
nor U22189 (N_22189,N_20044,N_19763);
nand U22190 (N_22190,N_20225,N_18732);
nor U22191 (N_22191,N_19706,N_19829);
nand U22192 (N_22192,N_19352,N_20531);
nor U22193 (N_22193,N_18240,N_20154);
xor U22194 (N_22194,N_20837,N_18747);
and U22195 (N_22195,N_20433,N_19051);
or U22196 (N_22196,N_20905,N_18563);
and U22197 (N_22197,N_19880,N_19869);
nand U22198 (N_22198,N_18492,N_18046);
and U22199 (N_22199,N_18032,N_20065);
xnor U22200 (N_22200,N_20957,N_18751);
nand U22201 (N_22201,N_20818,N_19064);
or U22202 (N_22202,N_20823,N_20315);
and U22203 (N_22203,N_18242,N_20666);
nand U22204 (N_22204,N_20912,N_18529);
or U22205 (N_22205,N_20471,N_19982);
nand U22206 (N_22206,N_19730,N_18129);
nor U22207 (N_22207,N_19151,N_19042);
or U22208 (N_22208,N_20854,N_19333);
or U22209 (N_22209,N_20880,N_20403);
nand U22210 (N_22210,N_19784,N_18383);
nor U22211 (N_22211,N_20728,N_19928);
xnor U22212 (N_22212,N_19446,N_19916);
and U22213 (N_22213,N_20716,N_18959);
nand U22214 (N_22214,N_20022,N_18618);
or U22215 (N_22215,N_20596,N_18816);
or U22216 (N_22216,N_19066,N_20675);
and U22217 (N_22217,N_20676,N_18880);
nor U22218 (N_22218,N_20861,N_20428);
xnor U22219 (N_22219,N_18685,N_20572);
xor U22220 (N_22220,N_20113,N_19117);
and U22221 (N_22221,N_18141,N_19004);
nor U22222 (N_22222,N_19558,N_20556);
and U22223 (N_22223,N_20998,N_18949);
or U22224 (N_22224,N_19069,N_18811);
or U22225 (N_22225,N_20297,N_19826);
or U22226 (N_22226,N_19527,N_20816);
and U22227 (N_22227,N_20143,N_19562);
nand U22228 (N_22228,N_20099,N_18843);
and U22229 (N_22229,N_18875,N_19113);
nand U22230 (N_22230,N_19171,N_18415);
or U22231 (N_22231,N_19849,N_19832);
nand U22232 (N_22232,N_19704,N_20170);
nand U22233 (N_22233,N_18138,N_20561);
or U22234 (N_22234,N_20280,N_18325);
and U22235 (N_22235,N_18216,N_19788);
and U22236 (N_22236,N_19193,N_20839);
nor U22237 (N_22237,N_19809,N_19146);
or U22238 (N_22238,N_19904,N_19356);
nand U22239 (N_22239,N_18656,N_19769);
and U22240 (N_22240,N_18012,N_20757);
nand U22241 (N_22241,N_20777,N_19043);
nand U22242 (N_22242,N_20914,N_18398);
nand U22243 (N_22243,N_20221,N_20384);
or U22244 (N_22244,N_18740,N_18005);
xor U22245 (N_22245,N_19986,N_18978);
xor U22246 (N_22246,N_20101,N_20970);
and U22247 (N_22247,N_18530,N_18966);
and U22248 (N_22248,N_18953,N_19594);
nand U22249 (N_22249,N_20175,N_18695);
or U22250 (N_22250,N_18019,N_20103);
nand U22251 (N_22251,N_18304,N_19371);
and U22252 (N_22252,N_20032,N_19617);
nand U22253 (N_22253,N_18036,N_18282);
nor U22254 (N_22254,N_19876,N_20848);
or U22255 (N_22255,N_19140,N_20455);
xor U22256 (N_22256,N_20289,N_18867);
and U22257 (N_22257,N_18199,N_19545);
and U22258 (N_22258,N_20959,N_18613);
nand U22259 (N_22259,N_19260,N_19400);
xor U22260 (N_22260,N_20208,N_18724);
nand U22261 (N_22261,N_20475,N_19189);
nand U22262 (N_22262,N_19877,N_19144);
nand U22263 (N_22263,N_18716,N_18055);
or U22264 (N_22264,N_19864,N_19011);
nand U22265 (N_22265,N_18176,N_18350);
or U22266 (N_22266,N_19720,N_20305);
nand U22267 (N_22267,N_19576,N_20008);
xnor U22268 (N_22268,N_19278,N_20199);
nor U22269 (N_22269,N_18488,N_19660);
nand U22270 (N_22270,N_19029,N_20353);
and U22271 (N_22271,N_20984,N_20222);
nor U22272 (N_22272,N_19292,N_19330);
or U22273 (N_22273,N_20887,N_19679);
and U22274 (N_22274,N_19695,N_20483);
or U22275 (N_22275,N_18748,N_19533);
nand U22276 (N_22276,N_20282,N_19932);
nor U22277 (N_22277,N_18459,N_19208);
nor U22278 (N_22278,N_19376,N_20105);
nand U22279 (N_22279,N_18088,N_19850);
or U22280 (N_22280,N_19580,N_19181);
and U22281 (N_22281,N_18082,N_18753);
nand U22282 (N_22282,N_19137,N_19148);
nand U22283 (N_22283,N_19732,N_19567);
nor U22284 (N_22284,N_18425,N_20705);
xnor U22285 (N_22285,N_19969,N_19369);
xor U22286 (N_22286,N_18620,N_18879);
nand U22287 (N_22287,N_18273,N_20232);
nand U22288 (N_22288,N_20468,N_19422);
nor U22289 (N_22289,N_18741,N_19762);
and U22290 (N_22290,N_20985,N_20026);
or U22291 (N_22291,N_20240,N_19844);
nand U22292 (N_22292,N_18294,N_18490);
nor U22293 (N_22293,N_18791,N_18206);
and U22294 (N_22294,N_20907,N_18534);
and U22295 (N_22295,N_18972,N_18166);
and U22296 (N_22296,N_19443,N_18066);
xor U22297 (N_22297,N_19390,N_18593);
nand U22298 (N_22298,N_20279,N_19953);
nand U22299 (N_22299,N_18069,N_20444);
nor U22300 (N_22300,N_18172,N_19433);
or U22301 (N_22301,N_20723,N_19571);
or U22302 (N_22302,N_20149,N_20064);
or U22303 (N_22303,N_20824,N_19610);
xnor U22304 (N_22304,N_20439,N_19701);
or U22305 (N_22305,N_20205,N_20253);
or U22306 (N_22306,N_19639,N_18721);
xnor U22307 (N_22307,N_18544,N_20469);
and U22308 (N_22308,N_20266,N_18823);
or U22309 (N_22309,N_19794,N_20367);
xnor U22310 (N_22310,N_20767,N_18601);
or U22311 (N_22311,N_20285,N_18674);
or U22312 (N_22312,N_19289,N_19968);
and U22313 (N_22313,N_20694,N_20890);
nand U22314 (N_22314,N_19735,N_19367);
nor U22315 (N_22315,N_20223,N_18633);
and U22316 (N_22316,N_18928,N_18430);
and U22317 (N_22317,N_18016,N_20810);
or U22318 (N_22318,N_18094,N_19486);
and U22319 (N_22319,N_20835,N_18451);
nor U22320 (N_22320,N_18006,N_18163);
nand U22321 (N_22321,N_20027,N_20446);
and U22322 (N_22322,N_18591,N_18899);
and U22323 (N_22323,N_20503,N_18442);
nand U22324 (N_22324,N_20227,N_19729);
xor U22325 (N_22325,N_19629,N_18051);
nor U22326 (N_22326,N_20200,N_19363);
and U22327 (N_22327,N_18896,N_18639);
and U22328 (N_22328,N_19717,N_20486);
or U22329 (N_22329,N_18810,N_19719);
and U22330 (N_22330,N_20267,N_18886);
or U22331 (N_22331,N_20109,N_19074);
or U22332 (N_22332,N_18437,N_19368);
nand U22333 (N_22333,N_20911,N_20499);
nand U22334 (N_22334,N_18739,N_18317);
and U22335 (N_22335,N_20576,N_19771);
xor U22336 (N_22336,N_20226,N_20009);
xor U22337 (N_22337,N_19546,N_19902);
or U22338 (N_22338,N_18962,N_18485);
xor U22339 (N_22339,N_20536,N_20121);
nand U22340 (N_22340,N_18491,N_20943);
xor U22341 (N_22341,N_18738,N_19207);
and U22342 (N_22342,N_18915,N_18352);
nor U22343 (N_22343,N_18832,N_18521);
nand U22344 (N_22344,N_18111,N_18349);
nor U22345 (N_22345,N_18194,N_18819);
and U22346 (N_22346,N_18977,N_18694);
xor U22347 (N_22347,N_20963,N_20447);
nor U22348 (N_22348,N_20051,N_18665);
and U22349 (N_22349,N_20930,N_18318);
and U22350 (N_22350,N_18554,N_19168);
or U22351 (N_22351,N_20910,N_19222);
xnor U22352 (N_22352,N_19495,N_18008);
xor U22353 (N_22353,N_18043,N_18525);
and U22354 (N_22354,N_20642,N_20229);
or U22355 (N_22355,N_20466,N_18851);
xor U22356 (N_22356,N_18795,N_18627);
xnor U22357 (N_22357,N_18648,N_19016);
nand U22358 (N_22358,N_19635,N_19543);
or U22359 (N_22359,N_19874,N_19127);
or U22360 (N_22360,N_20710,N_19943);
nand U22361 (N_22361,N_19825,N_18229);
xnor U22362 (N_22362,N_19393,N_20067);
or U22363 (N_22363,N_18184,N_18076);
nor U22364 (N_22364,N_18923,N_18454);
nand U22365 (N_22365,N_19694,N_20030);
and U22366 (N_22366,N_19619,N_20558);
or U22367 (N_22367,N_19159,N_18761);
or U22368 (N_22368,N_20087,N_20292);
nand U22369 (N_22369,N_18671,N_19023);
and U22370 (N_22370,N_19765,N_18435);
or U22371 (N_22371,N_18920,N_19782);
nand U22372 (N_22372,N_19271,N_18569);
nand U22373 (N_22373,N_19875,N_20869);
or U22374 (N_22374,N_18275,N_20853);
nor U22375 (N_22375,N_19296,N_19040);
and U22376 (N_22376,N_20769,N_18498);
nand U22377 (N_22377,N_19628,N_19747);
nand U22378 (N_22378,N_20550,N_20430);
nand U22379 (N_22379,N_18047,N_20559);
nand U22380 (N_22380,N_20789,N_19071);
nand U22381 (N_22381,N_19374,N_20798);
nor U22382 (N_22382,N_19595,N_18600);
nor U22383 (N_22383,N_18792,N_20882);
xor U22384 (N_22384,N_18588,N_19537);
nor U22385 (N_22385,N_20873,N_19917);
or U22386 (N_22386,N_18445,N_19511);
and U22387 (N_22387,N_19741,N_18939);
xnor U22388 (N_22388,N_18420,N_19929);
and U22389 (N_22389,N_18077,N_20746);
xnor U22390 (N_22390,N_19254,N_20144);
or U22391 (N_22391,N_18831,N_20481);
nand U22392 (N_22392,N_19338,N_20334);
and U22393 (N_22393,N_18171,N_19912);
and U22394 (N_22394,N_18010,N_18231);
and U22395 (N_22395,N_20775,N_18862);
nand U22396 (N_22396,N_19465,N_18687);
nor U22397 (N_22397,N_20831,N_19851);
nor U22398 (N_22398,N_20296,N_18477);
or U22399 (N_22399,N_20614,N_19450);
xnor U22400 (N_22400,N_20301,N_20638);
xnor U22401 (N_22401,N_20711,N_19882);
nor U22402 (N_22402,N_18805,N_18504);
or U22403 (N_22403,N_19945,N_19143);
and U22404 (N_22404,N_20198,N_20579);
and U22405 (N_22405,N_20377,N_18493);
xnor U22406 (N_22406,N_18386,N_19005);
xnor U22407 (N_22407,N_18543,N_19323);
or U22408 (N_22408,N_18225,N_18249);
or U22409 (N_22409,N_19999,N_19974);
nand U22410 (N_22410,N_19285,N_19414);
nand U22411 (N_22411,N_19952,N_18424);
xnor U22412 (N_22412,N_18572,N_18930);
nand U22413 (N_22413,N_20607,N_18293);
and U22414 (N_22414,N_19115,N_20701);
nor U22415 (N_22415,N_18045,N_19133);
nand U22416 (N_22416,N_19748,N_18769);
nor U22417 (N_22417,N_20071,N_20534);
and U22418 (N_22418,N_18407,N_20461);
nand U22419 (N_22419,N_20729,N_19162);
nand U22420 (N_22420,N_18640,N_20153);
nand U22421 (N_22421,N_20303,N_20029);
and U22422 (N_22422,N_19284,N_20476);
nand U22423 (N_22423,N_18201,N_18981);
or U22424 (N_22424,N_20059,N_19516);
or U22425 (N_22425,N_18027,N_19795);
and U22426 (N_22426,N_20722,N_18757);
xnor U22427 (N_22427,N_19941,N_18626);
nand U22428 (N_22428,N_19225,N_18126);
or U22429 (N_22429,N_20494,N_20119);
xnor U22430 (N_22430,N_19508,N_19538);
or U22431 (N_22431,N_20548,N_18568);
or U22432 (N_22432,N_20012,N_20774);
nand U22433 (N_22433,N_20904,N_20731);
xor U22434 (N_22434,N_20526,N_18328);
nor U22435 (N_22435,N_20413,N_18778);
nand U22436 (N_22436,N_18252,N_18698);
nand U22437 (N_22437,N_20975,N_18557);
nor U22438 (N_22438,N_18941,N_20828);
or U22439 (N_22439,N_20148,N_19648);
nor U22440 (N_22440,N_20674,N_19972);
or U22441 (N_22441,N_20751,N_20017);
or U22442 (N_22442,N_19910,N_18429);
nand U22443 (N_22443,N_20785,N_18503);
and U22444 (N_22444,N_20120,N_19640);
xnor U22445 (N_22445,N_18372,N_19317);
nor U22446 (N_22446,N_19828,N_19938);
nand U22447 (N_22447,N_19274,N_18502);
nor U22448 (N_22448,N_20133,N_18848);
nand U22449 (N_22449,N_19386,N_18144);
xnor U22450 (N_22450,N_18841,N_18666);
and U22451 (N_22451,N_19258,N_19304);
nor U22452 (N_22452,N_20049,N_19740);
xor U22453 (N_22453,N_20979,N_19138);
or U22454 (N_22454,N_19522,N_19962);
xnor U22455 (N_22455,N_20020,N_18824);
nor U22456 (N_22456,N_18519,N_20129);
xnor U22457 (N_22457,N_20050,N_19724);
nor U22458 (N_22458,N_19123,N_20594);
nand U22459 (N_22459,N_20827,N_18157);
xnor U22460 (N_22460,N_20125,N_18647);
xor U22461 (N_22461,N_20840,N_20921);
nor U22462 (N_22462,N_20435,N_19997);
nand U22463 (N_22463,N_19257,N_18402);
xor U22464 (N_22464,N_18921,N_18071);
nand U22465 (N_22465,N_20209,N_18917);
or U22466 (N_22466,N_18873,N_19196);
or U22467 (N_22467,N_18606,N_19090);
nand U22468 (N_22468,N_18124,N_20652);
and U22469 (N_22469,N_19432,N_18177);
xor U22470 (N_22470,N_19641,N_20126);
xnor U22471 (N_22471,N_18159,N_18664);
nor U22472 (N_22472,N_19419,N_20264);
and U22473 (N_22473,N_20368,N_19174);
nor U22474 (N_22474,N_20437,N_19894);
and U22475 (N_22475,N_20495,N_20639);
or U22476 (N_22476,N_20164,N_18466);
nor U22477 (N_22477,N_18573,N_18772);
xor U22478 (N_22478,N_18363,N_19650);
xor U22479 (N_22479,N_18182,N_20571);
nand U22480 (N_22480,N_20069,N_18542);
xor U22481 (N_22481,N_18774,N_20972);
nor U22482 (N_22482,N_19983,N_20197);
nand U22483 (N_22483,N_19190,N_19126);
or U22484 (N_22484,N_19429,N_20925);
nand U22485 (N_22485,N_18720,N_20319);
nor U22486 (N_22486,N_19936,N_19202);
or U22487 (N_22487,N_18882,N_20916);
nand U22488 (N_22488,N_18165,N_18001);
or U22489 (N_22489,N_19931,N_19251);
nand U22490 (N_22490,N_19037,N_19234);
nand U22491 (N_22491,N_20181,N_20948);
or U22492 (N_22492,N_20046,N_19396);
nand U22493 (N_22493,N_19092,N_19790);
nor U22494 (N_22494,N_20454,N_20504);
nand U22495 (N_22495,N_20220,N_18983);
or U22496 (N_22496,N_19840,N_19086);
nand U22497 (N_22497,N_20408,N_19235);
nand U22498 (N_22498,N_19860,N_20474);
or U22499 (N_22499,N_19039,N_20456);
nor U22500 (N_22500,N_20945,N_19537);
and U22501 (N_22501,N_20554,N_20565);
xnor U22502 (N_22502,N_19462,N_19832);
xor U22503 (N_22503,N_20303,N_18992);
or U22504 (N_22504,N_20617,N_19467);
xnor U22505 (N_22505,N_18416,N_18192);
xor U22506 (N_22506,N_20657,N_18761);
or U22507 (N_22507,N_19255,N_18624);
and U22508 (N_22508,N_20796,N_18482);
nand U22509 (N_22509,N_19514,N_18053);
or U22510 (N_22510,N_20870,N_19317);
or U22511 (N_22511,N_20832,N_18664);
or U22512 (N_22512,N_20411,N_20810);
and U22513 (N_22513,N_18051,N_19146);
or U22514 (N_22514,N_19668,N_19156);
or U22515 (N_22515,N_18240,N_20483);
nand U22516 (N_22516,N_18994,N_18627);
nand U22517 (N_22517,N_18871,N_20247);
nor U22518 (N_22518,N_18305,N_20804);
nand U22519 (N_22519,N_20397,N_18302);
nand U22520 (N_22520,N_19053,N_20146);
or U22521 (N_22521,N_20804,N_18447);
or U22522 (N_22522,N_19133,N_19291);
xnor U22523 (N_22523,N_18354,N_19216);
xnor U22524 (N_22524,N_20540,N_18278);
or U22525 (N_22525,N_20539,N_19271);
and U22526 (N_22526,N_19378,N_18846);
or U22527 (N_22527,N_19181,N_20167);
xor U22528 (N_22528,N_18653,N_18836);
nand U22529 (N_22529,N_20136,N_19715);
nor U22530 (N_22530,N_18257,N_19276);
or U22531 (N_22531,N_19515,N_20382);
nor U22532 (N_22532,N_19369,N_18342);
or U22533 (N_22533,N_19716,N_20867);
or U22534 (N_22534,N_19479,N_19913);
xor U22535 (N_22535,N_18662,N_18082);
nand U22536 (N_22536,N_18087,N_20717);
xnor U22537 (N_22537,N_18742,N_19550);
or U22538 (N_22538,N_18736,N_20154);
xor U22539 (N_22539,N_19430,N_20416);
and U22540 (N_22540,N_19447,N_18699);
or U22541 (N_22541,N_20018,N_19117);
nand U22542 (N_22542,N_19964,N_19644);
xor U22543 (N_22543,N_20836,N_19296);
and U22544 (N_22544,N_19335,N_18951);
nand U22545 (N_22545,N_18831,N_20763);
nor U22546 (N_22546,N_19010,N_19785);
or U22547 (N_22547,N_19218,N_20639);
nand U22548 (N_22548,N_20820,N_18434);
nor U22549 (N_22549,N_20308,N_19340);
or U22550 (N_22550,N_19919,N_20365);
nor U22551 (N_22551,N_20248,N_18516);
nand U22552 (N_22552,N_19030,N_20524);
nor U22553 (N_22553,N_18287,N_18938);
xor U22554 (N_22554,N_19457,N_20182);
or U22555 (N_22555,N_20573,N_18063);
nand U22556 (N_22556,N_18695,N_20674);
or U22557 (N_22557,N_20991,N_18942);
or U22558 (N_22558,N_20775,N_19884);
nor U22559 (N_22559,N_20758,N_20271);
xnor U22560 (N_22560,N_19154,N_18388);
xor U22561 (N_22561,N_18894,N_18161);
or U22562 (N_22562,N_18514,N_20642);
and U22563 (N_22563,N_18019,N_19583);
or U22564 (N_22564,N_18568,N_19950);
and U22565 (N_22565,N_18177,N_20088);
and U22566 (N_22566,N_19030,N_20709);
nor U22567 (N_22567,N_18982,N_19173);
and U22568 (N_22568,N_20066,N_19349);
and U22569 (N_22569,N_18452,N_20113);
or U22570 (N_22570,N_19160,N_19398);
nor U22571 (N_22571,N_18791,N_20052);
or U22572 (N_22572,N_18142,N_20071);
or U22573 (N_22573,N_19861,N_18158);
nand U22574 (N_22574,N_20975,N_20586);
nand U22575 (N_22575,N_18776,N_20070);
or U22576 (N_22576,N_20616,N_18878);
xnor U22577 (N_22577,N_19941,N_19838);
nor U22578 (N_22578,N_19537,N_19296);
or U22579 (N_22579,N_20782,N_18070);
or U22580 (N_22580,N_19445,N_18412);
xor U22581 (N_22581,N_19407,N_19480);
or U22582 (N_22582,N_20446,N_20331);
or U22583 (N_22583,N_20416,N_20474);
nor U22584 (N_22584,N_18720,N_18388);
xor U22585 (N_22585,N_19930,N_20613);
nor U22586 (N_22586,N_20997,N_19703);
or U22587 (N_22587,N_18912,N_20200);
nor U22588 (N_22588,N_18043,N_20447);
xor U22589 (N_22589,N_18821,N_18737);
nor U22590 (N_22590,N_18013,N_20284);
nor U22591 (N_22591,N_19357,N_20810);
xnor U22592 (N_22592,N_18613,N_20669);
nor U22593 (N_22593,N_20597,N_19811);
nor U22594 (N_22594,N_20645,N_18758);
nand U22595 (N_22595,N_18927,N_20008);
nand U22596 (N_22596,N_18027,N_19682);
nor U22597 (N_22597,N_18968,N_20388);
xor U22598 (N_22598,N_19986,N_18252);
and U22599 (N_22599,N_20362,N_19695);
xor U22600 (N_22600,N_18879,N_18661);
nor U22601 (N_22601,N_20799,N_20844);
nand U22602 (N_22602,N_18301,N_20778);
xor U22603 (N_22603,N_18969,N_20214);
and U22604 (N_22604,N_19043,N_18957);
xor U22605 (N_22605,N_18280,N_20250);
nor U22606 (N_22606,N_18073,N_18174);
xor U22607 (N_22607,N_20570,N_19740);
and U22608 (N_22608,N_19712,N_18462);
nor U22609 (N_22609,N_19678,N_18706);
nand U22610 (N_22610,N_20562,N_19968);
and U22611 (N_22611,N_20405,N_18305);
nor U22612 (N_22612,N_18160,N_20933);
or U22613 (N_22613,N_19862,N_18140);
and U22614 (N_22614,N_19118,N_19487);
nand U22615 (N_22615,N_18351,N_18173);
nor U22616 (N_22616,N_19904,N_20431);
nor U22617 (N_22617,N_20228,N_18115);
and U22618 (N_22618,N_19992,N_19851);
nand U22619 (N_22619,N_20918,N_19186);
xnor U22620 (N_22620,N_18630,N_18169);
nor U22621 (N_22621,N_19718,N_20529);
nor U22622 (N_22622,N_18663,N_20105);
nand U22623 (N_22623,N_18804,N_20635);
xnor U22624 (N_22624,N_20940,N_18955);
xnor U22625 (N_22625,N_19642,N_20920);
and U22626 (N_22626,N_18431,N_19984);
nor U22627 (N_22627,N_20399,N_20400);
and U22628 (N_22628,N_20193,N_18044);
xnor U22629 (N_22629,N_19893,N_18608);
and U22630 (N_22630,N_20818,N_19337);
and U22631 (N_22631,N_19473,N_18281);
or U22632 (N_22632,N_18808,N_18738);
nor U22633 (N_22633,N_20652,N_20648);
or U22634 (N_22634,N_19996,N_18541);
nor U22635 (N_22635,N_18689,N_20080);
nand U22636 (N_22636,N_20873,N_18099);
and U22637 (N_22637,N_20237,N_18694);
xnor U22638 (N_22638,N_18368,N_18976);
xor U22639 (N_22639,N_20559,N_19228);
xnor U22640 (N_22640,N_20160,N_18517);
nand U22641 (N_22641,N_20140,N_19299);
nand U22642 (N_22642,N_20447,N_20083);
and U22643 (N_22643,N_20958,N_20758);
xnor U22644 (N_22644,N_20671,N_19232);
nor U22645 (N_22645,N_18258,N_20134);
and U22646 (N_22646,N_18552,N_18979);
xnor U22647 (N_22647,N_18975,N_19392);
nor U22648 (N_22648,N_18266,N_20903);
or U22649 (N_22649,N_18187,N_18544);
nor U22650 (N_22650,N_19803,N_18346);
or U22651 (N_22651,N_20046,N_20365);
or U22652 (N_22652,N_18949,N_20418);
nand U22653 (N_22653,N_18950,N_18449);
xnor U22654 (N_22654,N_19942,N_19540);
or U22655 (N_22655,N_19724,N_18561);
nand U22656 (N_22656,N_18524,N_18368);
or U22657 (N_22657,N_18225,N_20980);
xnor U22658 (N_22658,N_20955,N_19425);
and U22659 (N_22659,N_20745,N_18147);
and U22660 (N_22660,N_20817,N_19535);
and U22661 (N_22661,N_20789,N_19810);
xnor U22662 (N_22662,N_18173,N_20024);
nor U22663 (N_22663,N_19601,N_19260);
or U22664 (N_22664,N_18975,N_19552);
nand U22665 (N_22665,N_20656,N_20535);
xnor U22666 (N_22666,N_19821,N_20522);
nand U22667 (N_22667,N_20779,N_19021);
xnor U22668 (N_22668,N_20091,N_18905);
xor U22669 (N_22669,N_18672,N_19345);
nor U22670 (N_22670,N_19513,N_19409);
nor U22671 (N_22671,N_20419,N_19463);
nor U22672 (N_22672,N_20473,N_20464);
or U22673 (N_22673,N_18635,N_20111);
or U22674 (N_22674,N_20665,N_19727);
xor U22675 (N_22675,N_20251,N_18147);
xnor U22676 (N_22676,N_20880,N_19453);
or U22677 (N_22677,N_18999,N_18203);
or U22678 (N_22678,N_20373,N_19075);
nand U22679 (N_22679,N_20340,N_20467);
nor U22680 (N_22680,N_19669,N_20598);
and U22681 (N_22681,N_20615,N_18287);
or U22682 (N_22682,N_20366,N_18588);
nand U22683 (N_22683,N_20797,N_19819);
xnor U22684 (N_22684,N_18482,N_19337);
nor U22685 (N_22685,N_20572,N_19840);
nor U22686 (N_22686,N_18690,N_19605);
xor U22687 (N_22687,N_20049,N_18329);
xnor U22688 (N_22688,N_19511,N_20184);
nor U22689 (N_22689,N_20585,N_20856);
nor U22690 (N_22690,N_20999,N_19948);
xnor U22691 (N_22691,N_18569,N_18903);
nand U22692 (N_22692,N_19032,N_18276);
nand U22693 (N_22693,N_19532,N_19743);
nand U22694 (N_22694,N_19434,N_18844);
xor U22695 (N_22695,N_18825,N_18850);
or U22696 (N_22696,N_18970,N_19559);
nor U22697 (N_22697,N_19131,N_20500);
and U22698 (N_22698,N_20683,N_19108);
or U22699 (N_22699,N_19357,N_20509);
or U22700 (N_22700,N_18008,N_18767);
or U22701 (N_22701,N_18652,N_20984);
nor U22702 (N_22702,N_20350,N_19160);
nor U22703 (N_22703,N_19266,N_20760);
and U22704 (N_22704,N_19098,N_20767);
nand U22705 (N_22705,N_18300,N_18541);
nor U22706 (N_22706,N_19130,N_19691);
nor U22707 (N_22707,N_20789,N_18252);
xor U22708 (N_22708,N_19905,N_19793);
and U22709 (N_22709,N_20849,N_19040);
nand U22710 (N_22710,N_19759,N_18019);
or U22711 (N_22711,N_18226,N_19144);
or U22712 (N_22712,N_19688,N_20055);
nor U22713 (N_22713,N_19394,N_20037);
nor U22714 (N_22714,N_18082,N_18615);
nor U22715 (N_22715,N_19172,N_20890);
nor U22716 (N_22716,N_20131,N_20939);
or U22717 (N_22717,N_20668,N_20181);
and U22718 (N_22718,N_20014,N_18765);
or U22719 (N_22719,N_19799,N_20579);
nand U22720 (N_22720,N_20879,N_20917);
nand U22721 (N_22721,N_20471,N_20973);
or U22722 (N_22722,N_18641,N_19558);
xor U22723 (N_22723,N_19497,N_19660);
nand U22724 (N_22724,N_19891,N_20343);
nor U22725 (N_22725,N_18258,N_19566);
nand U22726 (N_22726,N_19889,N_18042);
or U22727 (N_22727,N_19845,N_18745);
nor U22728 (N_22728,N_19907,N_18387);
xor U22729 (N_22729,N_19971,N_18739);
nor U22730 (N_22730,N_18325,N_18575);
xnor U22731 (N_22731,N_18850,N_20154);
and U22732 (N_22732,N_18914,N_19906);
nor U22733 (N_22733,N_18421,N_18452);
nand U22734 (N_22734,N_18586,N_19378);
xnor U22735 (N_22735,N_19186,N_20028);
nor U22736 (N_22736,N_18609,N_19486);
and U22737 (N_22737,N_19690,N_19714);
and U22738 (N_22738,N_18624,N_20043);
nor U22739 (N_22739,N_20444,N_19260);
nor U22740 (N_22740,N_18935,N_19183);
nand U22741 (N_22741,N_20420,N_18826);
or U22742 (N_22742,N_20835,N_18949);
nor U22743 (N_22743,N_20645,N_20351);
xor U22744 (N_22744,N_20930,N_20913);
xor U22745 (N_22745,N_19216,N_20276);
nand U22746 (N_22746,N_19928,N_18938);
xor U22747 (N_22747,N_20480,N_18099);
and U22748 (N_22748,N_18993,N_19373);
nor U22749 (N_22749,N_18545,N_19595);
and U22750 (N_22750,N_18607,N_18911);
and U22751 (N_22751,N_19853,N_20978);
nor U22752 (N_22752,N_20853,N_19726);
xnor U22753 (N_22753,N_18323,N_18142);
or U22754 (N_22754,N_20721,N_20697);
xor U22755 (N_22755,N_20318,N_18998);
or U22756 (N_22756,N_18741,N_20508);
nand U22757 (N_22757,N_20385,N_19028);
nand U22758 (N_22758,N_19045,N_19224);
nand U22759 (N_22759,N_18542,N_18295);
or U22760 (N_22760,N_20387,N_19142);
and U22761 (N_22761,N_20048,N_20692);
and U22762 (N_22762,N_19813,N_20623);
and U22763 (N_22763,N_20884,N_19252);
nor U22764 (N_22764,N_19925,N_18510);
nand U22765 (N_22765,N_19924,N_19402);
and U22766 (N_22766,N_20186,N_19228);
nor U22767 (N_22767,N_18400,N_19967);
xor U22768 (N_22768,N_19993,N_19712);
or U22769 (N_22769,N_19949,N_20945);
or U22770 (N_22770,N_19539,N_18501);
nor U22771 (N_22771,N_18057,N_18465);
and U22772 (N_22772,N_20854,N_18777);
and U22773 (N_22773,N_18212,N_20060);
or U22774 (N_22774,N_19301,N_20290);
nor U22775 (N_22775,N_20272,N_20300);
nor U22776 (N_22776,N_18846,N_18935);
nor U22777 (N_22777,N_20837,N_19262);
and U22778 (N_22778,N_19044,N_20799);
nor U22779 (N_22779,N_19504,N_20933);
xnor U22780 (N_22780,N_18478,N_19603);
xnor U22781 (N_22781,N_18092,N_20873);
xor U22782 (N_22782,N_19782,N_18816);
or U22783 (N_22783,N_18589,N_18498);
xor U22784 (N_22784,N_18282,N_18073);
and U22785 (N_22785,N_20573,N_19748);
nor U22786 (N_22786,N_19488,N_19399);
nor U22787 (N_22787,N_20370,N_18210);
nor U22788 (N_22788,N_20768,N_19506);
nor U22789 (N_22789,N_18371,N_20389);
xor U22790 (N_22790,N_20811,N_19265);
nand U22791 (N_22791,N_20618,N_19194);
xor U22792 (N_22792,N_19730,N_18626);
and U22793 (N_22793,N_20349,N_18641);
nor U22794 (N_22794,N_19513,N_20331);
nor U22795 (N_22795,N_19345,N_18342);
xnor U22796 (N_22796,N_18619,N_20740);
nor U22797 (N_22797,N_18097,N_19108);
or U22798 (N_22798,N_19726,N_20950);
xnor U22799 (N_22799,N_18682,N_19025);
or U22800 (N_22800,N_20391,N_19865);
nand U22801 (N_22801,N_19792,N_20953);
or U22802 (N_22802,N_18621,N_18487);
xnor U22803 (N_22803,N_18566,N_19345);
or U22804 (N_22804,N_18566,N_20673);
or U22805 (N_22805,N_20451,N_18433);
nor U22806 (N_22806,N_20058,N_19489);
xnor U22807 (N_22807,N_18285,N_19645);
nor U22808 (N_22808,N_19060,N_18236);
nand U22809 (N_22809,N_18608,N_18735);
or U22810 (N_22810,N_18898,N_18802);
or U22811 (N_22811,N_20042,N_18986);
and U22812 (N_22812,N_18288,N_18442);
nor U22813 (N_22813,N_20782,N_19647);
nor U22814 (N_22814,N_20896,N_20928);
nand U22815 (N_22815,N_20478,N_20633);
nor U22816 (N_22816,N_18343,N_18838);
nor U22817 (N_22817,N_20489,N_18072);
and U22818 (N_22818,N_19324,N_19381);
and U22819 (N_22819,N_20532,N_18319);
and U22820 (N_22820,N_20668,N_19427);
nand U22821 (N_22821,N_19417,N_20965);
and U22822 (N_22822,N_19424,N_19792);
nor U22823 (N_22823,N_20221,N_20719);
or U22824 (N_22824,N_20225,N_19118);
xnor U22825 (N_22825,N_18587,N_19334);
and U22826 (N_22826,N_19560,N_20886);
and U22827 (N_22827,N_20638,N_19611);
xor U22828 (N_22828,N_20216,N_18287);
nand U22829 (N_22829,N_19796,N_20090);
nor U22830 (N_22830,N_18374,N_19055);
nand U22831 (N_22831,N_18783,N_20872);
or U22832 (N_22832,N_18583,N_19954);
or U22833 (N_22833,N_20168,N_20032);
or U22834 (N_22834,N_19599,N_19380);
xor U22835 (N_22835,N_20020,N_18895);
xnor U22836 (N_22836,N_20970,N_18266);
nor U22837 (N_22837,N_20966,N_20554);
nand U22838 (N_22838,N_20091,N_18203);
or U22839 (N_22839,N_18374,N_19937);
nand U22840 (N_22840,N_18877,N_19462);
nand U22841 (N_22841,N_19925,N_18225);
nand U22842 (N_22842,N_18428,N_18594);
nor U22843 (N_22843,N_18926,N_18058);
nor U22844 (N_22844,N_18752,N_19451);
nor U22845 (N_22845,N_20885,N_20112);
and U22846 (N_22846,N_19675,N_20783);
nor U22847 (N_22847,N_19736,N_20892);
and U22848 (N_22848,N_18283,N_18929);
or U22849 (N_22849,N_19064,N_18346);
and U22850 (N_22850,N_20726,N_18776);
xnor U22851 (N_22851,N_20943,N_18233);
and U22852 (N_22852,N_18558,N_19908);
xnor U22853 (N_22853,N_18878,N_20797);
or U22854 (N_22854,N_20630,N_20675);
nor U22855 (N_22855,N_20452,N_19050);
nand U22856 (N_22856,N_19517,N_19589);
xnor U22857 (N_22857,N_19734,N_19762);
or U22858 (N_22858,N_19710,N_19163);
or U22859 (N_22859,N_19367,N_19914);
xnor U22860 (N_22860,N_18939,N_20198);
xor U22861 (N_22861,N_18392,N_20275);
xor U22862 (N_22862,N_18252,N_19410);
or U22863 (N_22863,N_19919,N_19390);
and U22864 (N_22864,N_19510,N_19643);
and U22865 (N_22865,N_18345,N_18475);
xor U22866 (N_22866,N_18525,N_18615);
nand U22867 (N_22867,N_20436,N_20009);
nor U22868 (N_22868,N_19092,N_18341);
xnor U22869 (N_22869,N_20136,N_18177);
nor U22870 (N_22870,N_20925,N_20389);
and U22871 (N_22871,N_18349,N_20978);
nand U22872 (N_22872,N_19250,N_20312);
xor U22873 (N_22873,N_19224,N_18412);
xor U22874 (N_22874,N_19544,N_20294);
or U22875 (N_22875,N_18150,N_18062);
or U22876 (N_22876,N_18064,N_20772);
nor U22877 (N_22877,N_20135,N_18346);
and U22878 (N_22878,N_20687,N_19043);
nand U22879 (N_22879,N_20687,N_18998);
nand U22880 (N_22880,N_18430,N_20762);
or U22881 (N_22881,N_18735,N_18035);
nor U22882 (N_22882,N_19673,N_18177);
xnor U22883 (N_22883,N_18269,N_18875);
xor U22884 (N_22884,N_20385,N_20717);
or U22885 (N_22885,N_20284,N_19363);
and U22886 (N_22886,N_19869,N_18480);
xnor U22887 (N_22887,N_20733,N_18787);
xor U22888 (N_22888,N_18962,N_19175);
nor U22889 (N_22889,N_20444,N_20151);
nand U22890 (N_22890,N_20009,N_18579);
nand U22891 (N_22891,N_19248,N_19182);
nand U22892 (N_22892,N_19550,N_20658);
nand U22893 (N_22893,N_20611,N_18699);
or U22894 (N_22894,N_18868,N_18765);
nor U22895 (N_22895,N_18134,N_18725);
nor U22896 (N_22896,N_19272,N_20927);
or U22897 (N_22897,N_18937,N_20012);
nor U22898 (N_22898,N_19070,N_18426);
xnor U22899 (N_22899,N_18383,N_18528);
nand U22900 (N_22900,N_20415,N_20609);
or U22901 (N_22901,N_19895,N_18148);
nor U22902 (N_22902,N_20944,N_18202);
nand U22903 (N_22903,N_18106,N_19947);
nor U22904 (N_22904,N_18707,N_18327);
or U22905 (N_22905,N_20123,N_20258);
or U22906 (N_22906,N_20778,N_19956);
nand U22907 (N_22907,N_20704,N_18809);
and U22908 (N_22908,N_19190,N_19134);
and U22909 (N_22909,N_18397,N_20667);
nor U22910 (N_22910,N_18988,N_19277);
nor U22911 (N_22911,N_20403,N_18978);
nor U22912 (N_22912,N_18067,N_20215);
nand U22913 (N_22913,N_18288,N_20273);
and U22914 (N_22914,N_18969,N_19152);
xnor U22915 (N_22915,N_20704,N_19414);
nor U22916 (N_22916,N_20136,N_19744);
nor U22917 (N_22917,N_19581,N_18845);
or U22918 (N_22918,N_19772,N_19463);
or U22919 (N_22919,N_19536,N_20079);
nor U22920 (N_22920,N_19998,N_19988);
and U22921 (N_22921,N_18994,N_19899);
or U22922 (N_22922,N_20621,N_20715);
nand U22923 (N_22923,N_18598,N_18718);
and U22924 (N_22924,N_19984,N_19873);
or U22925 (N_22925,N_20974,N_19444);
and U22926 (N_22926,N_19739,N_19113);
xnor U22927 (N_22927,N_18370,N_20695);
nand U22928 (N_22928,N_20410,N_19937);
nand U22929 (N_22929,N_20452,N_19295);
and U22930 (N_22930,N_18405,N_19922);
and U22931 (N_22931,N_20353,N_19475);
and U22932 (N_22932,N_19875,N_18401);
xnor U22933 (N_22933,N_20568,N_19040);
nor U22934 (N_22934,N_18375,N_18720);
xnor U22935 (N_22935,N_19369,N_18355);
xor U22936 (N_22936,N_19478,N_20199);
and U22937 (N_22937,N_20562,N_18625);
nand U22938 (N_22938,N_19922,N_19570);
xor U22939 (N_22939,N_18350,N_20878);
nand U22940 (N_22940,N_19759,N_19707);
nor U22941 (N_22941,N_20892,N_19172);
or U22942 (N_22942,N_19353,N_18451);
and U22943 (N_22943,N_19542,N_19104);
nor U22944 (N_22944,N_20105,N_19308);
xor U22945 (N_22945,N_20604,N_19604);
xnor U22946 (N_22946,N_20562,N_19958);
nor U22947 (N_22947,N_18839,N_19949);
nand U22948 (N_22948,N_18048,N_18912);
nand U22949 (N_22949,N_18853,N_18699);
and U22950 (N_22950,N_18432,N_18639);
or U22951 (N_22951,N_20237,N_20291);
and U22952 (N_22952,N_18499,N_19288);
xor U22953 (N_22953,N_19368,N_20944);
nor U22954 (N_22954,N_19641,N_20391);
and U22955 (N_22955,N_20490,N_19750);
xor U22956 (N_22956,N_19829,N_19024);
and U22957 (N_22957,N_18569,N_20365);
or U22958 (N_22958,N_20653,N_19556);
or U22959 (N_22959,N_18564,N_18782);
or U22960 (N_22960,N_18365,N_19005);
or U22961 (N_22961,N_20472,N_19720);
nand U22962 (N_22962,N_18763,N_19235);
nand U22963 (N_22963,N_18860,N_19630);
nand U22964 (N_22964,N_19209,N_20418);
or U22965 (N_22965,N_19721,N_20572);
or U22966 (N_22966,N_18914,N_18929);
and U22967 (N_22967,N_19806,N_20470);
nand U22968 (N_22968,N_19402,N_18441);
xnor U22969 (N_22969,N_19202,N_18855);
nand U22970 (N_22970,N_19418,N_19789);
nand U22971 (N_22971,N_18279,N_20430);
nor U22972 (N_22972,N_19551,N_18458);
nor U22973 (N_22973,N_18753,N_18178);
nand U22974 (N_22974,N_20100,N_18936);
nor U22975 (N_22975,N_18705,N_20251);
or U22976 (N_22976,N_18708,N_20862);
and U22977 (N_22977,N_19350,N_19203);
and U22978 (N_22978,N_20487,N_20736);
nor U22979 (N_22979,N_20648,N_18582);
nor U22980 (N_22980,N_18064,N_18026);
nand U22981 (N_22981,N_20427,N_18756);
nand U22982 (N_22982,N_18724,N_19354);
nor U22983 (N_22983,N_20712,N_20729);
nor U22984 (N_22984,N_19088,N_20043);
nand U22985 (N_22985,N_19213,N_19412);
or U22986 (N_22986,N_20875,N_20903);
or U22987 (N_22987,N_18087,N_20196);
xor U22988 (N_22988,N_19808,N_20958);
nor U22989 (N_22989,N_19360,N_19144);
or U22990 (N_22990,N_19641,N_20816);
nor U22991 (N_22991,N_19940,N_19997);
and U22992 (N_22992,N_19876,N_19444);
and U22993 (N_22993,N_20922,N_20249);
or U22994 (N_22994,N_18765,N_19005);
nand U22995 (N_22995,N_20577,N_18351);
nor U22996 (N_22996,N_20264,N_20775);
xor U22997 (N_22997,N_19078,N_20191);
and U22998 (N_22998,N_19764,N_20848);
nand U22999 (N_22999,N_20221,N_19360);
or U23000 (N_23000,N_19817,N_19777);
xnor U23001 (N_23001,N_19125,N_18980);
nor U23002 (N_23002,N_18578,N_20989);
xor U23003 (N_23003,N_18354,N_20473);
nand U23004 (N_23004,N_18420,N_18816);
xnor U23005 (N_23005,N_18523,N_20333);
xor U23006 (N_23006,N_18362,N_20931);
xnor U23007 (N_23007,N_20039,N_19928);
or U23008 (N_23008,N_20339,N_18137);
nand U23009 (N_23009,N_18926,N_20762);
and U23010 (N_23010,N_20828,N_20819);
and U23011 (N_23011,N_19872,N_18403);
xor U23012 (N_23012,N_20634,N_18142);
and U23013 (N_23013,N_20367,N_18787);
nand U23014 (N_23014,N_19287,N_19731);
and U23015 (N_23015,N_20133,N_18280);
xor U23016 (N_23016,N_18004,N_18631);
or U23017 (N_23017,N_18397,N_18550);
nand U23018 (N_23018,N_18349,N_18960);
nor U23019 (N_23019,N_19180,N_19622);
nand U23020 (N_23020,N_19146,N_20543);
xor U23021 (N_23021,N_19520,N_20671);
nor U23022 (N_23022,N_18726,N_20419);
xnor U23023 (N_23023,N_19650,N_18492);
xor U23024 (N_23024,N_19030,N_18338);
nand U23025 (N_23025,N_19689,N_19577);
nor U23026 (N_23026,N_19888,N_20640);
or U23027 (N_23027,N_18386,N_20777);
xnor U23028 (N_23028,N_19104,N_19505);
nand U23029 (N_23029,N_19888,N_19827);
and U23030 (N_23030,N_20133,N_20871);
xnor U23031 (N_23031,N_20447,N_18796);
xnor U23032 (N_23032,N_19762,N_19497);
nor U23033 (N_23033,N_19339,N_19556);
xnor U23034 (N_23034,N_20478,N_20868);
xor U23035 (N_23035,N_18154,N_19246);
xnor U23036 (N_23036,N_18871,N_18843);
xnor U23037 (N_23037,N_20163,N_20375);
nand U23038 (N_23038,N_19624,N_20303);
nand U23039 (N_23039,N_18784,N_18607);
nand U23040 (N_23040,N_19825,N_18620);
or U23041 (N_23041,N_19772,N_20474);
or U23042 (N_23042,N_19308,N_20485);
and U23043 (N_23043,N_19355,N_20490);
and U23044 (N_23044,N_20386,N_19754);
and U23045 (N_23045,N_18589,N_20328);
or U23046 (N_23046,N_20793,N_19048);
xnor U23047 (N_23047,N_19125,N_19319);
and U23048 (N_23048,N_20159,N_19113);
nand U23049 (N_23049,N_18899,N_20898);
or U23050 (N_23050,N_19994,N_19810);
or U23051 (N_23051,N_19453,N_20945);
and U23052 (N_23052,N_20872,N_20863);
nand U23053 (N_23053,N_18709,N_19924);
nand U23054 (N_23054,N_19773,N_20073);
xnor U23055 (N_23055,N_19910,N_18840);
and U23056 (N_23056,N_19133,N_18727);
and U23057 (N_23057,N_18420,N_18239);
nor U23058 (N_23058,N_20056,N_19489);
or U23059 (N_23059,N_19442,N_18038);
xnor U23060 (N_23060,N_18962,N_20765);
nand U23061 (N_23061,N_20686,N_20357);
xnor U23062 (N_23062,N_20378,N_18673);
nor U23063 (N_23063,N_19900,N_18381);
nor U23064 (N_23064,N_18504,N_19010);
nor U23065 (N_23065,N_19657,N_20607);
nand U23066 (N_23066,N_18671,N_19937);
nor U23067 (N_23067,N_19423,N_20453);
nand U23068 (N_23068,N_20172,N_19895);
and U23069 (N_23069,N_20979,N_20954);
or U23070 (N_23070,N_19430,N_18488);
xor U23071 (N_23071,N_18661,N_18822);
and U23072 (N_23072,N_19261,N_20872);
nand U23073 (N_23073,N_19820,N_18939);
or U23074 (N_23074,N_20911,N_18289);
and U23075 (N_23075,N_18656,N_18418);
nor U23076 (N_23076,N_19638,N_18014);
xor U23077 (N_23077,N_18767,N_20513);
xnor U23078 (N_23078,N_20240,N_20170);
xnor U23079 (N_23079,N_19292,N_20515);
nand U23080 (N_23080,N_18111,N_19460);
nand U23081 (N_23081,N_18011,N_20153);
xor U23082 (N_23082,N_19355,N_20288);
or U23083 (N_23083,N_19709,N_18136);
xnor U23084 (N_23084,N_19124,N_19972);
nor U23085 (N_23085,N_20814,N_18340);
nand U23086 (N_23086,N_20273,N_18480);
xor U23087 (N_23087,N_19018,N_20023);
xnor U23088 (N_23088,N_18533,N_19738);
nand U23089 (N_23089,N_20247,N_19567);
and U23090 (N_23090,N_19635,N_20345);
nand U23091 (N_23091,N_19038,N_18715);
nor U23092 (N_23092,N_19922,N_19407);
nand U23093 (N_23093,N_18712,N_19506);
xnor U23094 (N_23094,N_18351,N_20427);
and U23095 (N_23095,N_19573,N_20565);
and U23096 (N_23096,N_20751,N_19481);
nor U23097 (N_23097,N_19880,N_18515);
nor U23098 (N_23098,N_20404,N_20563);
and U23099 (N_23099,N_19669,N_18321);
xor U23100 (N_23100,N_19973,N_19239);
and U23101 (N_23101,N_20484,N_19579);
xor U23102 (N_23102,N_18178,N_19349);
or U23103 (N_23103,N_19882,N_18013);
nand U23104 (N_23104,N_20084,N_18210);
nand U23105 (N_23105,N_20768,N_18958);
nand U23106 (N_23106,N_19451,N_18202);
and U23107 (N_23107,N_18415,N_20506);
nand U23108 (N_23108,N_20319,N_20439);
or U23109 (N_23109,N_18586,N_19573);
nand U23110 (N_23110,N_18459,N_18345);
xor U23111 (N_23111,N_19215,N_18743);
nand U23112 (N_23112,N_20754,N_18855);
and U23113 (N_23113,N_20504,N_20183);
xnor U23114 (N_23114,N_20966,N_19049);
xor U23115 (N_23115,N_20389,N_20074);
xor U23116 (N_23116,N_18861,N_19610);
xnor U23117 (N_23117,N_20688,N_18792);
nor U23118 (N_23118,N_19439,N_20746);
or U23119 (N_23119,N_20498,N_20360);
nand U23120 (N_23120,N_19815,N_18332);
and U23121 (N_23121,N_20287,N_20727);
and U23122 (N_23122,N_19456,N_18022);
nor U23123 (N_23123,N_18333,N_20128);
or U23124 (N_23124,N_18867,N_20231);
xor U23125 (N_23125,N_19243,N_20053);
xnor U23126 (N_23126,N_18843,N_18399);
nand U23127 (N_23127,N_20798,N_19385);
and U23128 (N_23128,N_20571,N_19894);
or U23129 (N_23129,N_18794,N_20028);
and U23130 (N_23130,N_20921,N_20510);
xnor U23131 (N_23131,N_18838,N_18225);
nor U23132 (N_23132,N_20395,N_18433);
xnor U23133 (N_23133,N_18800,N_18420);
nor U23134 (N_23134,N_20768,N_19688);
nand U23135 (N_23135,N_19674,N_19409);
or U23136 (N_23136,N_18178,N_20714);
or U23137 (N_23137,N_18089,N_19184);
and U23138 (N_23138,N_20392,N_19074);
nand U23139 (N_23139,N_18230,N_18842);
nand U23140 (N_23140,N_20470,N_20056);
or U23141 (N_23141,N_18240,N_19579);
nor U23142 (N_23142,N_18231,N_20490);
or U23143 (N_23143,N_20681,N_20564);
xnor U23144 (N_23144,N_18255,N_18434);
xnor U23145 (N_23145,N_20778,N_19137);
nor U23146 (N_23146,N_19394,N_20527);
nor U23147 (N_23147,N_20474,N_19739);
xnor U23148 (N_23148,N_18734,N_18837);
nand U23149 (N_23149,N_20284,N_19431);
and U23150 (N_23150,N_20621,N_18388);
xor U23151 (N_23151,N_20443,N_20931);
or U23152 (N_23152,N_19087,N_18433);
and U23153 (N_23153,N_18042,N_19382);
and U23154 (N_23154,N_18211,N_18193);
and U23155 (N_23155,N_19878,N_19036);
nor U23156 (N_23156,N_18980,N_20079);
and U23157 (N_23157,N_18387,N_20227);
or U23158 (N_23158,N_18048,N_20085);
or U23159 (N_23159,N_19631,N_19785);
and U23160 (N_23160,N_20559,N_20280);
xnor U23161 (N_23161,N_18613,N_18013);
and U23162 (N_23162,N_19686,N_20107);
or U23163 (N_23163,N_20754,N_20955);
xnor U23164 (N_23164,N_20850,N_19513);
nor U23165 (N_23165,N_19451,N_19754);
xor U23166 (N_23166,N_20943,N_18917);
nor U23167 (N_23167,N_19248,N_19402);
or U23168 (N_23168,N_20633,N_20245);
xnor U23169 (N_23169,N_19099,N_20276);
nand U23170 (N_23170,N_19091,N_20781);
xnor U23171 (N_23171,N_20311,N_20898);
xor U23172 (N_23172,N_19098,N_19030);
and U23173 (N_23173,N_20159,N_18614);
nand U23174 (N_23174,N_19206,N_19795);
or U23175 (N_23175,N_18484,N_18879);
nand U23176 (N_23176,N_18070,N_19978);
xor U23177 (N_23177,N_19045,N_19513);
xor U23178 (N_23178,N_19550,N_18097);
nor U23179 (N_23179,N_20426,N_20618);
xor U23180 (N_23180,N_18413,N_18376);
or U23181 (N_23181,N_18690,N_20349);
nand U23182 (N_23182,N_20366,N_19247);
nor U23183 (N_23183,N_18694,N_18945);
nor U23184 (N_23184,N_20670,N_19889);
or U23185 (N_23185,N_20526,N_19210);
and U23186 (N_23186,N_19609,N_19637);
nor U23187 (N_23187,N_19450,N_18714);
xnor U23188 (N_23188,N_20471,N_18990);
and U23189 (N_23189,N_19402,N_18663);
nor U23190 (N_23190,N_18235,N_20743);
and U23191 (N_23191,N_18030,N_19446);
or U23192 (N_23192,N_20543,N_20635);
nand U23193 (N_23193,N_19541,N_18576);
xor U23194 (N_23194,N_20856,N_19683);
and U23195 (N_23195,N_19301,N_18723);
or U23196 (N_23196,N_20707,N_20947);
and U23197 (N_23197,N_20826,N_19101);
and U23198 (N_23198,N_18148,N_20599);
or U23199 (N_23199,N_20182,N_18578);
nor U23200 (N_23200,N_19892,N_18351);
xnor U23201 (N_23201,N_18217,N_18880);
xor U23202 (N_23202,N_18028,N_20243);
nor U23203 (N_23203,N_19997,N_20335);
or U23204 (N_23204,N_20950,N_19639);
and U23205 (N_23205,N_19073,N_19972);
nand U23206 (N_23206,N_20924,N_20695);
nor U23207 (N_23207,N_18242,N_19896);
nor U23208 (N_23208,N_19812,N_18785);
nand U23209 (N_23209,N_18408,N_20705);
nor U23210 (N_23210,N_20706,N_19154);
nand U23211 (N_23211,N_18374,N_20218);
and U23212 (N_23212,N_18683,N_20155);
nand U23213 (N_23213,N_20990,N_19277);
and U23214 (N_23214,N_18675,N_18674);
nor U23215 (N_23215,N_19006,N_20179);
nand U23216 (N_23216,N_18680,N_20322);
nor U23217 (N_23217,N_19543,N_18837);
or U23218 (N_23218,N_20153,N_20517);
or U23219 (N_23219,N_20216,N_19754);
nor U23220 (N_23220,N_19096,N_18957);
xnor U23221 (N_23221,N_20642,N_20187);
nand U23222 (N_23222,N_20915,N_20853);
nor U23223 (N_23223,N_20845,N_18008);
or U23224 (N_23224,N_19646,N_18150);
or U23225 (N_23225,N_19129,N_20292);
xor U23226 (N_23226,N_20163,N_19718);
xor U23227 (N_23227,N_18547,N_19593);
and U23228 (N_23228,N_20721,N_20792);
nand U23229 (N_23229,N_18141,N_18546);
nand U23230 (N_23230,N_19679,N_19051);
xor U23231 (N_23231,N_20540,N_18546);
xor U23232 (N_23232,N_19629,N_18539);
xnor U23233 (N_23233,N_19487,N_20498);
xor U23234 (N_23234,N_20760,N_18883);
or U23235 (N_23235,N_19135,N_19527);
xor U23236 (N_23236,N_18282,N_19071);
nor U23237 (N_23237,N_19308,N_20085);
or U23238 (N_23238,N_19592,N_18903);
and U23239 (N_23239,N_20387,N_19372);
xnor U23240 (N_23240,N_20483,N_20631);
and U23241 (N_23241,N_18509,N_19255);
xor U23242 (N_23242,N_19015,N_19548);
or U23243 (N_23243,N_20613,N_20473);
and U23244 (N_23244,N_18207,N_19504);
and U23245 (N_23245,N_18266,N_18877);
xor U23246 (N_23246,N_20383,N_20098);
nor U23247 (N_23247,N_19144,N_20694);
or U23248 (N_23248,N_20251,N_20752);
xor U23249 (N_23249,N_20167,N_18329);
nand U23250 (N_23250,N_19893,N_19707);
or U23251 (N_23251,N_20671,N_20294);
xnor U23252 (N_23252,N_19936,N_18149);
xnor U23253 (N_23253,N_19679,N_20905);
nor U23254 (N_23254,N_20415,N_20775);
nand U23255 (N_23255,N_18745,N_19721);
and U23256 (N_23256,N_19738,N_19327);
nand U23257 (N_23257,N_20749,N_20381);
or U23258 (N_23258,N_18767,N_19946);
xnor U23259 (N_23259,N_18495,N_20731);
or U23260 (N_23260,N_20777,N_19749);
xor U23261 (N_23261,N_20942,N_18946);
or U23262 (N_23262,N_19913,N_20396);
and U23263 (N_23263,N_19627,N_20339);
or U23264 (N_23264,N_19745,N_19635);
and U23265 (N_23265,N_19564,N_18165);
nand U23266 (N_23266,N_19481,N_20728);
nor U23267 (N_23267,N_18104,N_20798);
nand U23268 (N_23268,N_18894,N_19212);
nand U23269 (N_23269,N_20679,N_19062);
xnor U23270 (N_23270,N_18553,N_18741);
or U23271 (N_23271,N_18065,N_19227);
xnor U23272 (N_23272,N_20099,N_18169);
xnor U23273 (N_23273,N_18967,N_19903);
or U23274 (N_23274,N_19544,N_19929);
or U23275 (N_23275,N_18376,N_20776);
or U23276 (N_23276,N_20615,N_19547);
xor U23277 (N_23277,N_20798,N_20305);
nand U23278 (N_23278,N_18473,N_18642);
and U23279 (N_23279,N_18485,N_18594);
xnor U23280 (N_23280,N_20683,N_18990);
or U23281 (N_23281,N_18810,N_20687);
or U23282 (N_23282,N_18742,N_19943);
and U23283 (N_23283,N_19787,N_18564);
or U23284 (N_23284,N_18468,N_18852);
and U23285 (N_23285,N_19952,N_19701);
nand U23286 (N_23286,N_20766,N_19676);
nand U23287 (N_23287,N_19574,N_19750);
xor U23288 (N_23288,N_20248,N_18853);
nor U23289 (N_23289,N_18824,N_20178);
nand U23290 (N_23290,N_20670,N_20743);
or U23291 (N_23291,N_18811,N_20836);
nand U23292 (N_23292,N_19418,N_18503);
and U23293 (N_23293,N_18367,N_18382);
nor U23294 (N_23294,N_18514,N_20672);
xor U23295 (N_23295,N_19139,N_18064);
nor U23296 (N_23296,N_19133,N_19279);
or U23297 (N_23297,N_19437,N_18425);
and U23298 (N_23298,N_19697,N_19168);
nand U23299 (N_23299,N_20381,N_18140);
or U23300 (N_23300,N_19641,N_19017);
and U23301 (N_23301,N_18810,N_19160);
or U23302 (N_23302,N_18371,N_18893);
or U23303 (N_23303,N_20393,N_18584);
nand U23304 (N_23304,N_19341,N_19909);
nand U23305 (N_23305,N_20491,N_19642);
and U23306 (N_23306,N_18323,N_20675);
and U23307 (N_23307,N_19911,N_18625);
nor U23308 (N_23308,N_19780,N_18829);
and U23309 (N_23309,N_20357,N_18960);
xnor U23310 (N_23310,N_20149,N_20421);
and U23311 (N_23311,N_19240,N_18354);
xnor U23312 (N_23312,N_20794,N_19143);
or U23313 (N_23313,N_19682,N_18385);
nor U23314 (N_23314,N_20733,N_18165);
xor U23315 (N_23315,N_20257,N_19381);
xnor U23316 (N_23316,N_18412,N_19609);
nor U23317 (N_23317,N_20580,N_19707);
nor U23318 (N_23318,N_18610,N_20385);
nor U23319 (N_23319,N_19671,N_20310);
nor U23320 (N_23320,N_19960,N_18011);
nand U23321 (N_23321,N_18409,N_19786);
nand U23322 (N_23322,N_19136,N_19941);
and U23323 (N_23323,N_18085,N_19094);
xor U23324 (N_23324,N_19526,N_20016);
and U23325 (N_23325,N_19955,N_18490);
nor U23326 (N_23326,N_20154,N_19409);
or U23327 (N_23327,N_19908,N_19406);
and U23328 (N_23328,N_19799,N_20598);
nor U23329 (N_23329,N_19686,N_18786);
or U23330 (N_23330,N_20561,N_18331);
xnor U23331 (N_23331,N_18725,N_18909);
nor U23332 (N_23332,N_19024,N_19438);
nand U23333 (N_23333,N_20201,N_20465);
nand U23334 (N_23334,N_20624,N_20031);
xor U23335 (N_23335,N_19339,N_20544);
and U23336 (N_23336,N_19686,N_19635);
xnor U23337 (N_23337,N_19257,N_20419);
nand U23338 (N_23338,N_19233,N_20902);
nand U23339 (N_23339,N_18064,N_19264);
and U23340 (N_23340,N_18055,N_18424);
and U23341 (N_23341,N_18341,N_18047);
or U23342 (N_23342,N_20884,N_18046);
nor U23343 (N_23343,N_18178,N_18049);
xnor U23344 (N_23344,N_19174,N_19217);
xor U23345 (N_23345,N_19476,N_20618);
or U23346 (N_23346,N_20700,N_20203);
nand U23347 (N_23347,N_18975,N_18782);
xnor U23348 (N_23348,N_19015,N_18172);
nand U23349 (N_23349,N_18551,N_19993);
nand U23350 (N_23350,N_20520,N_19406);
nand U23351 (N_23351,N_18074,N_19007);
xor U23352 (N_23352,N_20683,N_19523);
and U23353 (N_23353,N_18020,N_19094);
or U23354 (N_23354,N_18757,N_18064);
nor U23355 (N_23355,N_19001,N_19816);
nand U23356 (N_23356,N_19920,N_20498);
nand U23357 (N_23357,N_18595,N_20218);
or U23358 (N_23358,N_20189,N_18691);
xor U23359 (N_23359,N_18009,N_18214);
or U23360 (N_23360,N_20128,N_18809);
nor U23361 (N_23361,N_20105,N_18066);
nor U23362 (N_23362,N_18680,N_20298);
and U23363 (N_23363,N_19151,N_19733);
xnor U23364 (N_23364,N_19682,N_19690);
nor U23365 (N_23365,N_20684,N_19661);
xor U23366 (N_23366,N_20767,N_18737);
nor U23367 (N_23367,N_19236,N_19580);
and U23368 (N_23368,N_19208,N_19156);
nor U23369 (N_23369,N_18137,N_18994);
nor U23370 (N_23370,N_19814,N_19562);
or U23371 (N_23371,N_18169,N_19497);
nor U23372 (N_23372,N_19641,N_20157);
nand U23373 (N_23373,N_20593,N_19475);
nor U23374 (N_23374,N_18625,N_20021);
nor U23375 (N_23375,N_20608,N_20270);
or U23376 (N_23376,N_18515,N_18572);
and U23377 (N_23377,N_20258,N_18542);
and U23378 (N_23378,N_20038,N_18966);
xor U23379 (N_23379,N_19704,N_18804);
nand U23380 (N_23380,N_19894,N_19529);
nand U23381 (N_23381,N_19089,N_18982);
and U23382 (N_23382,N_18747,N_19630);
nand U23383 (N_23383,N_20123,N_19542);
xor U23384 (N_23384,N_19356,N_18322);
nand U23385 (N_23385,N_20496,N_19985);
nor U23386 (N_23386,N_19076,N_18176);
or U23387 (N_23387,N_20846,N_19761);
and U23388 (N_23388,N_19528,N_18892);
and U23389 (N_23389,N_19390,N_19053);
and U23390 (N_23390,N_19327,N_20048);
xor U23391 (N_23391,N_19282,N_20822);
nand U23392 (N_23392,N_18521,N_18305);
xnor U23393 (N_23393,N_20034,N_19420);
xor U23394 (N_23394,N_18562,N_19309);
nor U23395 (N_23395,N_20290,N_18754);
xnor U23396 (N_23396,N_18749,N_18028);
nand U23397 (N_23397,N_19949,N_20744);
and U23398 (N_23398,N_19496,N_18376);
nand U23399 (N_23399,N_20329,N_20453);
xnor U23400 (N_23400,N_20639,N_18230);
and U23401 (N_23401,N_18847,N_20333);
or U23402 (N_23402,N_19505,N_18383);
or U23403 (N_23403,N_18830,N_20182);
and U23404 (N_23404,N_20541,N_19681);
xor U23405 (N_23405,N_19944,N_18324);
nand U23406 (N_23406,N_20508,N_18853);
nand U23407 (N_23407,N_19827,N_20977);
nor U23408 (N_23408,N_19819,N_18915);
nand U23409 (N_23409,N_19771,N_19522);
or U23410 (N_23410,N_18475,N_20104);
nor U23411 (N_23411,N_19019,N_18930);
or U23412 (N_23412,N_19458,N_20261);
nand U23413 (N_23413,N_20505,N_18841);
xnor U23414 (N_23414,N_19824,N_20064);
nand U23415 (N_23415,N_18480,N_18406);
nor U23416 (N_23416,N_19794,N_18015);
xnor U23417 (N_23417,N_19808,N_19844);
or U23418 (N_23418,N_20301,N_18617);
nand U23419 (N_23419,N_19209,N_18269);
or U23420 (N_23420,N_19942,N_18228);
and U23421 (N_23421,N_20519,N_18507);
and U23422 (N_23422,N_18408,N_19934);
nor U23423 (N_23423,N_18866,N_20575);
nor U23424 (N_23424,N_19593,N_20086);
or U23425 (N_23425,N_18393,N_19582);
nor U23426 (N_23426,N_20884,N_18870);
or U23427 (N_23427,N_19062,N_20215);
and U23428 (N_23428,N_18367,N_18926);
and U23429 (N_23429,N_19810,N_19741);
or U23430 (N_23430,N_19488,N_18311);
and U23431 (N_23431,N_20985,N_20143);
or U23432 (N_23432,N_20796,N_18312);
xor U23433 (N_23433,N_19701,N_18303);
xor U23434 (N_23434,N_19315,N_20338);
and U23435 (N_23435,N_19331,N_20015);
nor U23436 (N_23436,N_18704,N_20094);
nand U23437 (N_23437,N_20847,N_18888);
nand U23438 (N_23438,N_19204,N_18706);
and U23439 (N_23439,N_18704,N_19563);
nor U23440 (N_23440,N_20700,N_20136);
and U23441 (N_23441,N_19237,N_18893);
nand U23442 (N_23442,N_19777,N_18270);
nand U23443 (N_23443,N_19543,N_18932);
nand U23444 (N_23444,N_18144,N_19955);
nand U23445 (N_23445,N_19991,N_18614);
xor U23446 (N_23446,N_20784,N_19689);
xor U23447 (N_23447,N_18318,N_20866);
nor U23448 (N_23448,N_18166,N_19556);
or U23449 (N_23449,N_20375,N_19814);
or U23450 (N_23450,N_18481,N_18626);
xor U23451 (N_23451,N_19444,N_20096);
and U23452 (N_23452,N_18750,N_18911);
or U23453 (N_23453,N_18335,N_18255);
nand U23454 (N_23454,N_20117,N_18998);
nand U23455 (N_23455,N_19364,N_19893);
and U23456 (N_23456,N_20547,N_18785);
nand U23457 (N_23457,N_18936,N_18342);
or U23458 (N_23458,N_19573,N_19059);
nor U23459 (N_23459,N_20581,N_20827);
nor U23460 (N_23460,N_18157,N_20953);
nand U23461 (N_23461,N_18659,N_18673);
nor U23462 (N_23462,N_19470,N_19236);
and U23463 (N_23463,N_19605,N_20584);
xnor U23464 (N_23464,N_19055,N_19029);
nand U23465 (N_23465,N_18582,N_18816);
or U23466 (N_23466,N_18962,N_19087);
nor U23467 (N_23467,N_18986,N_18676);
nor U23468 (N_23468,N_20017,N_18083);
xor U23469 (N_23469,N_18759,N_18810);
or U23470 (N_23470,N_20386,N_18681);
or U23471 (N_23471,N_19589,N_19080);
nor U23472 (N_23472,N_20029,N_20438);
and U23473 (N_23473,N_18256,N_18070);
or U23474 (N_23474,N_20346,N_18720);
or U23475 (N_23475,N_18769,N_19414);
nor U23476 (N_23476,N_20964,N_19100);
and U23477 (N_23477,N_20229,N_18431);
xnor U23478 (N_23478,N_20492,N_20658);
xnor U23479 (N_23479,N_19904,N_20239);
nor U23480 (N_23480,N_19870,N_19091);
nand U23481 (N_23481,N_18096,N_18303);
nand U23482 (N_23482,N_19555,N_18378);
and U23483 (N_23483,N_20142,N_18816);
xnor U23484 (N_23484,N_19751,N_20873);
or U23485 (N_23485,N_20710,N_18711);
or U23486 (N_23486,N_19007,N_20142);
and U23487 (N_23487,N_19463,N_19443);
and U23488 (N_23488,N_19394,N_19908);
or U23489 (N_23489,N_20157,N_20899);
or U23490 (N_23490,N_20385,N_19189);
nor U23491 (N_23491,N_20080,N_19136);
xnor U23492 (N_23492,N_20481,N_20866);
and U23493 (N_23493,N_20185,N_20731);
nand U23494 (N_23494,N_19973,N_20430);
nand U23495 (N_23495,N_18037,N_18163);
or U23496 (N_23496,N_19280,N_20416);
and U23497 (N_23497,N_18008,N_18509);
or U23498 (N_23498,N_19835,N_20986);
xor U23499 (N_23499,N_19864,N_18582);
nand U23500 (N_23500,N_18281,N_18046);
nand U23501 (N_23501,N_19783,N_18847);
nand U23502 (N_23502,N_20281,N_20338);
or U23503 (N_23503,N_19478,N_20797);
nand U23504 (N_23504,N_19402,N_20859);
nor U23505 (N_23505,N_18221,N_20462);
nor U23506 (N_23506,N_20519,N_20117);
or U23507 (N_23507,N_20208,N_18752);
xor U23508 (N_23508,N_19197,N_18078);
xnor U23509 (N_23509,N_20649,N_18276);
or U23510 (N_23510,N_18004,N_20774);
nor U23511 (N_23511,N_18376,N_19841);
or U23512 (N_23512,N_18276,N_20704);
nand U23513 (N_23513,N_20908,N_18320);
nand U23514 (N_23514,N_19664,N_18136);
and U23515 (N_23515,N_20848,N_20387);
and U23516 (N_23516,N_20033,N_19490);
and U23517 (N_23517,N_18427,N_20463);
nand U23518 (N_23518,N_18989,N_20494);
and U23519 (N_23519,N_18926,N_18031);
and U23520 (N_23520,N_18772,N_20062);
nand U23521 (N_23521,N_18975,N_20880);
and U23522 (N_23522,N_19577,N_20339);
xor U23523 (N_23523,N_20000,N_18040);
nor U23524 (N_23524,N_18120,N_20958);
and U23525 (N_23525,N_19996,N_20556);
xnor U23526 (N_23526,N_19193,N_18283);
nand U23527 (N_23527,N_19757,N_18428);
or U23528 (N_23528,N_19080,N_18535);
xnor U23529 (N_23529,N_20242,N_20405);
and U23530 (N_23530,N_19658,N_18943);
nand U23531 (N_23531,N_18017,N_18099);
nand U23532 (N_23532,N_20287,N_18977);
nand U23533 (N_23533,N_20264,N_19185);
and U23534 (N_23534,N_20127,N_19289);
nand U23535 (N_23535,N_19140,N_18891);
nand U23536 (N_23536,N_18456,N_20372);
nand U23537 (N_23537,N_19627,N_20213);
nand U23538 (N_23538,N_18015,N_20507);
or U23539 (N_23539,N_18614,N_20239);
and U23540 (N_23540,N_19795,N_20783);
nor U23541 (N_23541,N_19728,N_18020);
nand U23542 (N_23542,N_20183,N_19341);
or U23543 (N_23543,N_20220,N_19542);
nor U23544 (N_23544,N_19640,N_18503);
nor U23545 (N_23545,N_19161,N_19682);
and U23546 (N_23546,N_18191,N_19224);
xor U23547 (N_23547,N_19531,N_18179);
nor U23548 (N_23548,N_19221,N_18564);
nand U23549 (N_23549,N_20946,N_20202);
nand U23550 (N_23550,N_18213,N_18804);
and U23551 (N_23551,N_18350,N_20500);
nand U23552 (N_23552,N_19819,N_20871);
and U23553 (N_23553,N_18698,N_18040);
nor U23554 (N_23554,N_19828,N_19361);
and U23555 (N_23555,N_18650,N_20440);
or U23556 (N_23556,N_20502,N_18157);
and U23557 (N_23557,N_18044,N_19631);
xor U23558 (N_23558,N_18532,N_19821);
or U23559 (N_23559,N_19881,N_19026);
xnor U23560 (N_23560,N_18116,N_20346);
and U23561 (N_23561,N_20534,N_20413);
and U23562 (N_23562,N_20833,N_19453);
nor U23563 (N_23563,N_18119,N_18822);
xnor U23564 (N_23564,N_18590,N_18568);
nor U23565 (N_23565,N_19790,N_19252);
or U23566 (N_23566,N_20624,N_19051);
or U23567 (N_23567,N_20088,N_19462);
xor U23568 (N_23568,N_20966,N_19793);
and U23569 (N_23569,N_19928,N_20254);
or U23570 (N_23570,N_18526,N_18693);
xnor U23571 (N_23571,N_18316,N_20460);
nor U23572 (N_23572,N_18533,N_18552);
xnor U23573 (N_23573,N_20171,N_18377);
and U23574 (N_23574,N_19230,N_20368);
and U23575 (N_23575,N_20986,N_20709);
nor U23576 (N_23576,N_18682,N_19146);
nand U23577 (N_23577,N_18043,N_20573);
xor U23578 (N_23578,N_19187,N_20369);
or U23579 (N_23579,N_18817,N_18627);
or U23580 (N_23580,N_19487,N_20812);
nor U23581 (N_23581,N_18946,N_19222);
nand U23582 (N_23582,N_18662,N_20908);
or U23583 (N_23583,N_20736,N_19435);
nand U23584 (N_23584,N_19121,N_19651);
nand U23585 (N_23585,N_20440,N_19693);
or U23586 (N_23586,N_19135,N_20087);
or U23587 (N_23587,N_18352,N_20371);
or U23588 (N_23588,N_18634,N_18428);
xor U23589 (N_23589,N_18808,N_18291);
nor U23590 (N_23590,N_20285,N_20485);
nor U23591 (N_23591,N_18840,N_18067);
nor U23592 (N_23592,N_20070,N_19871);
and U23593 (N_23593,N_20968,N_18394);
xor U23594 (N_23594,N_20295,N_19591);
and U23595 (N_23595,N_19585,N_19672);
nor U23596 (N_23596,N_19352,N_20441);
nand U23597 (N_23597,N_20375,N_20661);
or U23598 (N_23598,N_20563,N_20452);
and U23599 (N_23599,N_19323,N_19824);
or U23600 (N_23600,N_20453,N_19132);
nor U23601 (N_23601,N_20496,N_19119);
or U23602 (N_23602,N_19696,N_18876);
or U23603 (N_23603,N_19724,N_18339);
xor U23604 (N_23604,N_18418,N_18083);
or U23605 (N_23605,N_20795,N_20302);
xnor U23606 (N_23606,N_18536,N_18773);
xor U23607 (N_23607,N_18232,N_20244);
xor U23608 (N_23608,N_20475,N_18682);
xnor U23609 (N_23609,N_19102,N_18276);
nor U23610 (N_23610,N_18444,N_18631);
or U23611 (N_23611,N_20832,N_20646);
nand U23612 (N_23612,N_19803,N_20653);
and U23613 (N_23613,N_20000,N_19180);
xor U23614 (N_23614,N_20778,N_18125);
or U23615 (N_23615,N_20458,N_20198);
and U23616 (N_23616,N_18496,N_18981);
nor U23617 (N_23617,N_20722,N_20484);
xnor U23618 (N_23618,N_19179,N_19402);
or U23619 (N_23619,N_20765,N_18817);
nor U23620 (N_23620,N_20994,N_20017);
nor U23621 (N_23621,N_19699,N_20848);
and U23622 (N_23622,N_20620,N_18186);
nor U23623 (N_23623,N_18937,N_20966);
nand U23624 (N_23624,N_20843,N_18424);
xor U23625 (N_23625,N_20026,N_19916);
xor U23626 (N_23626,N_20789,N_18107);
nand U23627 (N_23627,N_18142,N_18046);
and U23628 (N_23628,N_20581,N_20225);
nand U23629 (N_23629,N_18015,N_19352);
nor U23630 (N_23630,N_19884,N_20565);
and U23631 (N_23631,N_20764,N_19750);
or U23632 (N_23632,N_18610,N_18227);
and U23633 (N_23633,N_19032,N_18831);
nand U23634 (N_23634,N_18643,N_20150);
nand U23635 (N_23635,N_18037,N_20824);
or U23636 (N_23636,N_19668,N_19136);
or U23637 (N_23637,N_18821,N_18882);
xor U23638 (N_23638,N_18417,N_18491);
and U23639 (N_23639,N_20618,N_19773);
nor U23640 (N_23640,N_18416,N_20134);
xor U23641 (N_23641,N_18531,N_19160);
xnor U23642 (N_23642,N_19851,N_18437);
nor U23643 (N_23643,N_19817,N_20212);
xor U23644 (N_23644,N_18989,N_18931);
xnor U23645 (N_23645,N_20837,N_20158);
or U23646 (N_23646,N_18712,N_19306);
or U23647 (N_23647,N_18240,N_19606);
nor U23648 (N_23648,N_18801,N_19937);
and U23649 (N_23649,N_20025,N_20615);
and U23650 (N_23650,N_19366,N_18466);
nand U23651 (N_23651,N_18710,N_20969);
nand U23652 (N_23652,N_18057,N_19853);
nor U23653 (N_23653,N_19838,N_18084);
or U23654 (N_23654,N_18518,N_19324);
and U23655 (N_23655,N_19793,N_19861);
xor U23656 (N_23656,N_18099,N_18796);
or U23657 (N_23657,N_20649,N_20266);
and U23658 (N_23658,N_18291,N_19252);
or U23659 (N_23659,N_18276,N_19934);
nor U23660 (N_23660,N_20892,N_20226);
or U23661 (N_23661,N_18131,N_20013);
nor U23662 (N_23662,N_20485,N_20321);
nand U23663 (N_23663,N_20657,N_19634);
xor U23664 (N_23664,N_20511,N_19162);
nand U23665 (N_23665,N_19539,N_18012);
nand U23666 (N_23666,N_20030,N_18483);
nor U23667 (N_23667,N_20924,N_18507);
xor U23668 (N_23668,N_19713,N_18983);
nand U23669 (N_23669,N_20650,N_19561);
nor U23670 (N_23670,N_18112,N_20153);
nor U23671 (N_23671,N_20803,N_19260);
and U23672 (N_23672,N_18802,N_18085);
xnor U23673 (N_23673,N_18959,N_20186);
xor U23674 (N_23674,N_19451,N_20262);
or U23675 (N_23675,N_20750,N_20052);
nor U23676 (N_23676,N_20216,N_18557);
nand U23677 (N_23677,N_20277,N_18682);
xor U23678 (N_23678,N_18088,N_20329);
xor U23679 (N_23679,N_20013,N_19523);
nand U23680 (N_23680,N_18116,N_18678);
nor U23681 (N_23681,N_20018,N_20463);
and U23682 (N_23682,N_20370,N_19745);
or U23683 (N_23683,N_19277,N_18213);
nand U23684 (N_23684,N_18598,N_18454);
and U23685 (N_23685,N_18367,N_20211);
or U23686 (N_23686,N_20109,N_18738);
nand U23687 (N_23687,N_19803,N_20257);
nor U23688 (N_23688,N_20275,N_20072);
xor U23689 (N_23689,N_20336,N_19610);
nor U23690 (N_23690,N_19465,N_18805);
and U23691 (N_23691,N_19675,N_20417);
or U23692 (N_23692,N_19334,N_20692);
xnor U23693 (N_23693,N_18974,N_18931);
nor U23694 (N_23694,N_20524,N_20463);
and U23695 (N_23695,N_18107,N_18735);
xnor U23696 (N_23696,N_20351,N_19753);
or U23697 (N_23697,N_20433,N_20167);
or U23698 (N_23698,N_20140,N_19955);
nand U23699 (N_23699,N_20205,N_18650);
and U23700 (N_23700,N_18334,N_18738);
nand U23701 (N_23701,N_19433,N_20655);
or U23702 (N_23702,N_19740,N_18520);
and U23703 (N_23703,N_20195,N_18985);
or U23704 (N_23704,N_19241,N_19508);
nand U23705 (N_23705,N_20546,N_18110);
xnor U23706 (N_23706,N_18817,N_19971);
nor U23707 (N_23707,N_20421,N_20467);
or U23708 (N_23708,N_18179,N_20352);
nand U23709 (N_23709,N_20928,N_18231);
nor U23710 (N_23710,N_18602,N_18474);
nand U23711 (N_23711,N_18319,N_20594);
nand U23712 (N_23712,N_20648,N_20080);
xnor U23713 (N_23713,N_20202,N_20526);
nor U23714 (N_23714,N_18890,N_19152);
nor U23715 (N_23715,N_20660,N_19161);
xnor U23716 (N_23716,N_18143,N_18054);
and U23717 (N_23717,N_20130,N_18854);
or U23718 (N_23718,N_18300,N_19370);
or U23719 (N_23719,N_18823,N_20561);
nor U23720 (N_23720,N_19358,N_20174);
xor U23721 (N_23721,N_20524,N_18349);
xnor U23722 (N_23722,N_19816,N_18003);
xor U23723 (N_23723,N_19596,N_20518);
nand U23724 (N_23724,N_20635,N_18345);
xor U23725 (N_23725,N_19544,N_20922);
or U23726 (N_23726,N_20888,N_18323);
xnor U23727 (N_23727,N_19896,N_20222);
or U23728 (N_23728,N_19378,N_20458);
or U23729 (N_23729,N_19515,N_20061);
nor U23730 (N_23730,N_19082,N_19392);
nor U23731 (N_23731,N_20785,N_20927);
nor U23732 (N_23732,N_20488,N_19043);
nand U23733 (N_23733,N_20293,N_18041);
or U23734 (N_23734,N_18731,N_18975);
nand U23735 (N_23735,N_18289,N_19027);
or U23736 (N_23736,N_18481,N_20603);
or U23737 (N_23737,N_19267,N_19300);
nand U23738 (N_23738,N_20929,N_19122);
and U23739 (N_23739,N_18754,N_19233);
and U23740 (N_23740,N_19738,N_19014);
or U23741 (N_23741,N_18112,N_19897);
or U23742 (N_23742,N_19509,N_20003);
or U23743 (N_23743,N_19442,N_18925);
nand U23744 (N_23744,N_19370,N_20789);
nand U23745 (N_23745,N_18786,N_18806);
nor U23746 (N_23746,N_18763,N_18995);
nor U23747 (N_23747,N_20488,N_20132);
nor U23748 (N_23748,N_20275,N_18244);
xnor U23749 (N_23749,N_19744,N_20339);
nor U23750 (N_23750,N_19358,N_19917);
xor U23751 (N_23751,N_19660,N_19152);
nand U23752 (N_23752,N_20238,N_19757);
nand U23753 (N_23753,N_18388,N_20812);
nand U23754 (N_23754,N_18060,N_18402);
and U23755 (N_23755,N_18707,N_19244);
nor U23756 (N_23756,N_18172,N_20183);
xor U23757 (N_23757,N_20750,N_18688);
nand U23758 (N_23758,N_19064,N_19801);
or U23759 (N_23759,N_19631,N_20077);
or U23760 (N_23760,N_19930,N_19494);
and U23761 (N_23761,N_20270,N_19402);
xnor U23762 (N_23762,N_19669,N_18540);
or U23763 (N_23763,N_20629,N_19190);
nor U23764 (N_23764,N_19870,N_19648);
xnor U23765 (N_23765,N_18365,N_18785);
or U23766 (N_23766,N_18301,N_19079);
nor U23767 (N_23767,N_20052,N_18269);
xnor U23768 (N_23768,N_20712,N_18839);
nor U23769 (N_23769,N_18807,N_20971);
and U23770 (N_23770,N_20122,N_19313);
xnor U23771 (N_23771,N_18651,N_19056);
nand U23772 (N_23772,N_20102,N_19899);
nor U23773 (N_23773,N_18319,N_20169);
and U23774 (N_23774,N_20673,N_18036);
nor U23775 (N_23775,N_19174,N_19523);
nand U23776 (N_23776,N_18137,N_20025);
or U23777 (N_23777,N_20961,N_18369);
nand U23778 (N_23778,N_18590,N_18608);
and U23779 (N_23779,N_19454,N_19552);
or U23780 (N_23780,N_20889,N_18706);
and U23781 (N_23781,N_18511,N_18949);
nand U23782 (N_23782,N_18709,N_18769);
nor U23783 (N_23783,N_20172,N_19859);
xor U23784 (N_23784,N_19416,N_20001);
nor U23785 (N_23785,N_20171,N_18168);
xnor U23786 (N_23786,N_19979,N_19761);
and U23787 (N_23787,N_20597,N_19948);
and U23788 (N_23788,N_19426,N_19844);
and U23789 (N_23789,N_18546,N_18040);
nand U23790 (N_23790,N_18644,N_18406);
nor U23791 (N_23791,N_19747,N_19648);
nand U23792 (N_23792,N_19062,N_18037);
nor U23793 (N_23793,N_19856,N_20376);
and U23794 (N_23794,N_18815,N_20015);
nor U23795 (N_23795,N_18458,N_18217);
nand U23796 (N_23796,N_20671,N_19223);
and U23797 (N_23797,N_20264,N_19758);
nand U23798 (N_23798,N_19365,N_19163);
xnor U23799 (N_23799,N_20120,N_18326);
xnor U23800 (N_23800,N_19325,N_18031);
or U23801 (N_23801,N_18151,N_18399);
or U23802 (N_23802,N_19257,N_18883);
xor U23803 (N_23803,N_20987,N_19271);
nand U23804 (N_23804,N_19448,N_19226);
nor U23805 (N_23805,N_18169,N_19244);
xor U23806 (N_23806,N_18660,N_18919);
or U23807 (N_23807,N_18536,N_20630);
xnor U23808 (N_23808,N_19235,N_19105);
nor U23809 (N_23809,N_18745,N_20810);
nand U23810 (N_23810,N_19914,N_18250);
and U23811 (N_23811,N_19825,N_20317);
nor U23812 (N_23812,N_19378,N_19936);
and U23813 (N_23813,N_19868,N_18128);
xnor U23814 (N_23814,N_20934,N_19724);
xor U23815 (N_23815,N_20018,N_19232);
nand U23816 (N_23816,N_18110,N_19228);
or U23817 (N_23817,N_20306,N_20612);
or U23818 (N_23818,N_18071,N_20697);
nand U23819 (N_23819,N_19419,N_19891);
xnor U23820 (N_23820,N_18808,N_18354);
or U23821 (N_23821,N_20638,N_18424);
or U23822 (N_23822,N_18354,N_20189);
nand U23823 (N_23823,N_18535,N_19639);
xnor U23824 (N_23824,N_18172,N_18407);
nand U23825 (N_23825,N_20542,N_19498);
nor U23826 (N_23826,N_18184,N_18425);
nor U23827 (N_23827,N_20053,N_20556);
and U23828 (N_23828,N_18141,N_18447);
xor U23829 (N_23829,N_20949,N_20150);
nor U23830 (N_23830,N_18790,N_20139);
and U23831 (N_23831,N_18957,N_19618);
and U23832 (N_23832,N_20783,N_20098);
or U23833 (N_23833,N_19166,N_18202);
nor U23834 (N_23834,N_19409,N_18535);
and U23835 (N_23835,N_19809,N_20750);
or U23836 (N_23836,N_18154,N_20236);
xor U23837 (N_23837,N_18501,N_20026);
and U23838 (N_23838,N_20741,N_19127);
xor U23839 (N_23839,N_20603,N_20019);
xor U23840 (N_23840,N_19079,N_18108);
xnor U23841 (N_23841,N_20336,N_19300);
and U23842 (N_23842,N_20198,N_18909);
nor U23843 (N_23843,N_20194,N_18232);
xnor U23844 (N_23844,N_18082,N_18162);
and U23845 (N_23845,N_20226,N_18916);
xor U23846 (N_23846,N_20105,N_19560);
or U23847 (N_23847,N_20385,N_19777);
xor U23848 (N_23848,N_18213,N_18061);
nand U23849 (N_23849,N_19182,N_19217);
nand U23850 (N_23850,N_20876,N_18240);
nand U23851 (N_23851,N_18081,N_19403);
nand U23852 (N_23852,N_19998,N_19258);
or U23853 (N_23853,N_18923,N_20407);
or U23854 (N_23854,N_19468,N_18634);
xor U23855 (N_23855,N_20392,N_20763);
nand U23856 (N_23856,N_18279,N_20362);
and U23857 (N_23857,N_19074,N_20631);
or U23858 (N_23858,N_18343,N_19960);
nand U23859 (N_23859,N_20700,N_19267);
or U23860 (N_23860,N_18294,N_20051);
xnor U23861 (N_23861,N_18424,N_18217);
or U23862 (N_23862,N_19416,N_19320);
xor U23863 (N_23863,N_20203,N_19590);
nor U23864 (N_23864,N_19486,N_20753);
xnor U23865 (N_23865,N_18736,N_18314);
xnor U23866 (N_23866,N_19254,N_18973);
nor U23867 (N_23867,N_20638,N_19666);
nand U23868 (N_23868,N_20708,N_20622);
nand U23869 (N_23869,N_19696,N_18628);
and U23870 (N_23870,N_20408,N_19623);
nor U23871 (N_23871,N_20818,N_18302);
nor U23872 (N_23872,N_18528,N_20479);
nor U23873 (N_23873,N_20070,N_18212);
and U23874 (N_23874,N_19854,N_19309);
or U23875 (N_23875,N_18523,N_19632);
or U23876 (N_23876,N_18789,N_18988);
nand U23877 (N_23877,N_18754,N_20373);
or U23878 (N_23878,N_18192,N_19626);
nor U23879 (N_23879,N_19039,N_18489);
and U23880 (N_23880,N_18048,N_20318);
xnor U23881 (N_23881,N_18988,N_20436);
xor U23882 (N_23882,N_19236,N_20625);
nor U23883 (N_23883,N_18399,N_20694);
nor U23884 (N_23884,N_19487,N_19207);
xnor U23885 (N_23885,N_18699,N_18979);
and U23886 (N_23886,N_18433,N_18686);
and U23887 (N_23887,N_20024,N_18169);
and U23888 (N_23888,N_18245,N_19396);
nor U23889 (N_23889,N_19955,N_19414);
and U23890 (N_23890,N_20047,N_18397);
xor U23891 (N_23891,N_20388,N_18775);
xor U23892 (N_23892,N_19102,N_18308);
and U23893 (N_23893,N_20281,N_19792);
xor U23894 (N_23894,N_19912,N_20486);
and U23895 (N_23895,N_18266,N_19175);
nand U23896 (N_23896,N_19424,N_18131);
nor U23897 (N_23897,N_20360,N_19363);
nand U23898 (N_23898,N_18609,N_19412);
or U23899 (N_23899,N_20122,N_19333);
and U23900 (N_23900,N_19689,N_20828);
nand U23901 (N_23901,N_20423,N_18791);
and U23902 (N_23902,N_20989,N_20919);
nand U23903 (N_23903,N_19608,N_19109);
or U23904 (N_23904,N_19159,N_19895);
xor U23905 (N_23905,N_19787,N_19477);
nand U23906 (N_23906,N_20849,N_18203);
nor U23907 (N_23907,N_18490,N_20968);
nand U23908 (N_23908,N_18707,N_18257);
nor U23909 (N_23909,N_20983,N_19085);
nand U23910 (N_23910,N_18394,N_19347);
or U23911 (N_23911,N_20989,N_20666);
or U23912 (N_23912,N_20663,N_20284);
nor U23913 (N_23913,N_18879,N_19650);
nand U23914 (N_23914,N_19315,N_20901);
nand U23915 (N_23915,N_19281,N_19451);
nor U23916 (N_23916,N_18393,N_19950);
and U23917 (N_23917,N_20117,N_20702);
xnor U23918 (N_23918,N_18384,N_19933);
or U23919 (N_23919,N_20473,N_18038);
xnor U23920 (N_23920,N_19257,N_18497);
nor U23921 (N_23921,N_20232,N_19447);
or U23922 (N_23922,N_20332,N_19789);
and U23923 (N_23923,N_18459,N_20314);
and U23924 (N_23924,N_20533,N_18683);
or U23925 (N_23925,N_20876,N_18145);
nor U23926 (N_23926,N_18321,N_18233);
or U23927 (N_23927,N_18673,N_20689);
xnor U23928 (N_23928,N_19464,N_19469);
or U23929 (N_23929,N_20813,N_19925);
or U23930 (N_23930,N_19429,N_19768);
nand U23931 (N_23931,N_20187,N_18671);
nand U23932 (N_23932,N_18278,N_19696);
and U23933 (N_23933,N_20067,N_20048);
nor U23934 (N_23934,N_20928,N_18625);
and U23935 (N_23935,N_19306,N_18252);
xnor U23936 (N_23936,N_18923,N_20676);
nor U23937 (N_23937,N_18783,N_18381);
and U23938 (N_23938,N_19832,N_20371);
or U23939 (N_23939,N_18809,N_20195);
nand U23940 (N_23940,N_19967,N_18741);
nand U23941 (N_23941,N_20492,N_20776);
xor U23942 (N_23942,N_20528,N_19694);
nor U23943 (N_23943,N_20072,N_20723);
xnor U23944 (N_23944,N_19980,N_20801);
nor U23945 (N_23945,N_19586,N_18700);
or U23946 (N_23946,N_18716,N_19912);
and U23947 (N_23947,N_20236,N_20533);
nor U23948 (N_23948,N_18008,N_19115);
nand U23949 (N_23949,N_19895,N_18139);
nand U23950 (N_23950,N_18714,N_20076);
nand U23951 (N_23951,N_19776,N_20809);
nand U23952 (N_23952,N_19101,N_19001);
and U23953 (N_23953,N_20716,N_18072);
and U23954 (N_23954,N_20537,N_20340);
nor U23955 (N_23955,N_18128,N_18835);
and U23956 (N_23956,N_20322,N_20272);
nor U23957 (N_23957,N_20656,N_19999);
xnor U23958 (N_23958,N_19292,N_19296);
xor U23959 (N_23959,N_19241,N_18313);
nand U23960 (N_23960,N_19846,N_18310);
xor U23961 (N_23961,N_20956,N_20738);
nor U23962 (N_23962,N_20814,N_18824);
or U23963 (N_23963,N_18823,N_18220);
nor U23964 (N_23964,N_19662,N_18169);
nor U23965 (N_23965,N_19794,N_19814);
or U23966 (N_23966,N_20749,N_18384);
and U23967 (N_23967,N_20830,N_20192);
nor U23968 (N_23968,N_19163,N_19619);
xnor U23969 (N_23969,N_20881,N_18154);
or U23970 (N_23970,N_19314,N_18025);
nand U23971 (N_23971,N_20207,N_20523);
or U23972 (N_23972,N_19725,N_19327);
nor U23973 (N_23973,N_20083,N_19922);
or U23974 (N_23974,N_20368,N_19092);
or U23975 (N_23975,N_19714,N_18343);
or U23976 (N_23976,N_18116,N_20383);
nor U23977 (N_23977,N_19426,N_19717);
xnor U23978 (N_23978,N_20154,N_20023);
nand U23979 (N_23979,N_20048,N_19765);
xor U23980 (N_23980,N_19765,N_18235);
xnor U23981 (N_23981,N_18644,N_18016);
xor U23982 (N_23982,N_20253,N_19593);
xor U23983 (N_23983,N_18675,N_18178);
or U23984 (N_23984,N_19973,N_20578);
and U23985 (N_23985,N_20962,N_20088);
and U23986 (N_23986,N_18131,N_18702);
or U23987 (N_23987,N_18001,N_19161);
nor U23988 (N_23988,N_20166,N_20383);
nand U23989 (N_23989,N_19859,N_18463);
or U23990 (N_23990,N_20620,N_20825);
or U23991 (N_23991,N_18115,N_19546);
or U23992 (N_23992,N_19460,N_19512);
nand U23993 (N_23993,N_20712,N_19353);
nor U23994 (N_23994,N_20377,N_18148);
and U23995 (N_23995,N_20149,N_18253);
and U23996 (N_23996,N_18047,N_19591);
and U23997 (N_23997,N_19487,N_20937);
xor U23998 (N_23998,N_20671,N_18004);
xnor U23999 (N_23999,N_20957,N_19459);
nand U24000 (N_24000,N_23559,N_23280);
nand U24001 (N_24001,N_21639,N_22641);
nor U24002 (N_24002,N_23549,N_21235);
nand U24003 (N_24003,N_23548,N_23542);
xnor U24004 (N_24004,N_23192,N_23832);
nand U24005 (N_24005,N_23632,N_22247);
xnor U24006 (N_24006,N_22864,N_23801);
or U24007 (N_24007,N_21311,N_23914);
or U24008 (N_24008,N_23410,N_23581);
nor U24009 (N_24009,N_21649,N_23400);
or U24010 (N_24010,N_21121,N_21840);
nand U24011 (N_24011,N_23792,N_22455);
nor U24012 (N_24012,N_22524,N_21561);
xnor U24013 (N_24013,N_23691,N_23350);
nor U24014 (N_24014,N_21026,N_21078);
nand U24015 (N_24015,N_21550,N_22317);
and U24016 (N_24016,N_23185,N_22561);
or U24017 (N_24017,N_23932,N_23418);
nor U24018 (N_24018,N_23329,N_22358);
nand U24019 (N_24019,N_21870,N_22067);
xor U24020 (N_24020,N_23814,N_22987);
or U24021 (N_24021,N_21719,N_23461);
or U24022 (N_24022,N_23576,N_23700);
nand U24023 (N_24023,N_22632,N_21593);
and U24024 (N_24024,N_23759,N_23655);
xor U24025 (N_24025,N_22112,N_23219);
nor U24026 (N_24026,N_22242,N_22644);
or U24027 (N_24027,N_23153,N_21605);
and U24028 (N_24028,N_22459,N_21459);
or U24029 (N_24029,N_21691,N_22918);
nor U24030 (N_24030,N_23658,N_23474);
nand U24031 (N_24031,N_23292,N_22735);
and U24032 (N_24032,N_22788,N_21970);
xnor U24033 (N_24033,N_22286,N_22947);
xor U24034 (N_24034,N_22044,N_23873);
xnor U24035 (N_24035,N_22300,N_23236);
nor U24036 (N_24036,N_22109,N_21763);
xnor U24037 (N_24037,N_21864,N_23490);
nor U24038 (N_24038,N_21946,N_23864);
nor U24039 (N_24039,N_21966,N_22677);
nor U24040 (N_24040,N_21402,N_21426);
and U24041 (N_24041,N_21543,N_22239);
or U24042 (N_24042,N_22333,N_23633);
nor U24043 (N_24043,N_23448,N_23084);
and U24044 (N_24044,N_22433,N_22703);
xor U24045 (N_24045,N_21520,N_23887);
and U24046 (N_24046,N_23966,N_23313);
or U24047 (N_24047,N_22752,N_21186);
or U24048 (N_24048,N_23718,N_23685);
or U24049 (N_24049,N_21917,N_22246);
or U24050 (N_24050,N_21337,N_22651);
and U24051 (N_24051,N_23096,N_21314);
nand U24052 (N_24052,N_23834,N_21660);
nand U24053 (N_24053,N_23485,N_23821);
nand U24054 (N_24054,N_22287,N_21565);
nor U24055 (N_24055,N_22270,N_22158);
nand U24056 (N_24056,N_22315,N_21357);
nor U24057 (N_24057,N_23766,N_21780);
nand U24058 (N_24058,N_23135,N_22734);
xor U24059 (N_24059,N_23360,N_22440);
and U24060 (N_24060,N_23199,N_21274);
xnor U24061 (N_24061,N_22631,N_21906);
xor U24062 (N_24062,N_21044,N_21199);
and U24063 (N_24063,N_21369,N_21204);
or U24064 (N_24064,N_22209,N_21401);
or U24065 (N_24065,N_21872,N_22751);
and U24066 (N_24066,N_21031,N_22263);
nand U24067 (N_24067,N_23877,N_22955);
nand U24068 (N_24068,N_22537,N_22323);
and U24069 (N_24069,N_22164,N_21448);
xor U24070 (N_24070,N_22303,N_23805);
xor U24071 (N_24071,N_23808,N_22890);
nor U24072 (N_24072,N_23369,N_23958);
xor U24073 (N_24073,N_23267,N_21869);
and U24074 (N_24074,N_22380,N_21677);
xnor U24075 (N_24075,N_22028,N_23977);
nand U24076 (N_24076,N_22061,N_23183);
or U24077 (N_24077,N_21024,N_23851);
nand U24078 (N_24078,N_23279,N_21484);
or U24079 (N_24079,N_23336,N_21434);
and U24080 (N_24080,N_22810,N_22123);
nand U24081 (N_24081,N_23128,N_23340);
xor U24082 (N_24082,N_21366,N_23197);
nor U24083 (N_24083,N_21263,N_22274);
xor U24084 (N_24084,N_22971,N_23242);
or U24085 (N_24085,N_23535,N_22689);
nand U24086 (N_24086,N_23435,N_23281);
nor U24087 (N_24087,N_21331,N_23493);
and U24088 (N_24088,N_21179,N_21535);
or U24089 (N_24089,N_22359,N_23810);
nor U24090 (N_24090,N_22063,N_21379);
xor U24091 (N_24091,N_22901,N_21531);
xor U24092 (N_24092,N_23269,N_21806);
xnor U24093 (N_24093,N_22460,N_23201);
and U24094 (N_24094,N_21042,N_23600);
or U24095 (N_24095,N_22761,N_22084);
and U24096 (N_24096,N_23919,N_23909);
nor U24097 (N_24097,N_22108,N_22225);
and U24098 (N_24098,N_23889,N_23622);
and U24099 (N_24099,N_21356,N_22930);
nor U24100 (N_24100,N_23896,N_22508);
nor U24101 (N_24101,N_21422,N_22948);
nor U24102 (N_24102,N_22593,N_23890);
nand U24103 (N_24103,N_21943,N_23593);
nand U24104 (N_24104,N_21583,N_23678);
xor U24105 (N_24105,N_23129,N_21417);
and U24106 (N_24106,N_21797,N_23934);
nand U24107 (N_24107,N_23200,N_21928);
or U24108 (N_24108,N_23579,N_22075);
nand U24109 (N_24109,N_21655,N_21015);
nand U24110 (N_24110,N_22452,N_21103);
nand U24111 (N_24111,N_21932,N_23294);
or U24112 (N_24112,N_21245,N_22032);
or U24113 (N_24113,N_21232,N_21809);
and U24114 (N_24114,N_21388,N_22978);
nand U24115 (N_24115,N_22215,N_23125);
nand U24116 (N_24116,N_23041,N_22293);
and U24117 (N_24117,N_22186,N_23748);
nand U24118 (N_24118,N_22523,N_23160);
nand U24119 (N_24119,N_23905,N_21383);
and U24120 (N_24120,N_21184,N_23845);
nor U24121 (N_24121,N_21393,N_23844);
and U24122 (N_24122,N_23843,N_23346);
nor U24123 (N_24123,N_22150,N_22970);
nor U24124 (N_24124,N_21815,N_22833);
nor U24125 (N_24125,N_23211,N_21482);
nor U24126 (N_24126,N_23960,N_23970);
nand U24127 (N_24127,N_22959,N_22352);
or U24128 (N_24128,N_22395,N_23922);
nand U24129 (N_24129,N_23308,N_21166);
xnor U24130 (N_24130,N_21053,N_23708);
and U24131 (N_24131,N_21124,N_22153);
xor U24132 (N_24132,N_22914,N_23532);
xor U24133 (N_24133,N_23785,N_21156);
and U24134 (N_24134,N_23869,N_23000);
and U24135 (N_24135,N_21335,N_21123);
nor U24136 (N_24136,N_21762,N_23662);
or U24137 (N_24137,N_23626,N_21244);
or U24138 (N_24138,N_21532,N_23429);
or U24139 (N_24139,N_21304,N_22763);
xnor U24140 (N_24140,N_23587,N_21487);
or U24141 (N_24141,N_23991,N_23547);
nand U24142 (N_24142,N_21773,N_22684);
and U24143 (N_24143,N_23690,N_22113);
xnor U24144 (N_24144,N_23916,N_23293);
or U24145 (N_24145,N_21193,N_23907);
nand U24146 (N_24146,N_23610,N_22705);
nor U24147 (N_24147,N_22094,N_21570);
xor U24148 (N_24148,N_21557,N_21058);
nor U24149 (N_24149,N_22927,N_22952);
or U24150 (N_24150,N_21433,N_21170);
xnor U24151 (N_24151,N_21884,N_23252);
or U24152 (N_24152,N_22887,N_23514);
and U24153 (N_24153,N_21699,N_21206);
nand U24154 (N_24154,N_21181,N_21116);
or U24155 (N_24155,N_21038,N_23320);
xnor U24156 (N_24156,N_22596,N_21662);
xnor U24157 (N_24157,N_23636,N_21858);
xnor U24158 (N_24158,N_22767,N_22878);
and U24159 (N_24159,N_22590,N_22698);
xor U24160 (N_24160,N_22818,N_23720);
nand U24161 (N_24161,N_22128,N_23165);
nand U24162 (N_24162,N_22973,N_23120);
xnor U24163 (N_24163,N_21391,N_23799);
and U24164 (N_24164,N_22271,N_21219);
and U24165 (N_24165,N_23781,N_23617);
or U24166 (N_24166,N_21903,N_22029);
nand U24167 (N_24167,N_22964,N_22551);
xnor U24168 (N_24168,N_21622,N_21555);
nand U24169 (N_24169,N_21808,N_23679);
xnor U24170 (N_24170,N_21405,N_22111);
or U24171 (N_24171,N_23455,N_21403);
or U24172 (N_24172,N_21326,N_23762);
nor U24173 (N_24173,N_21959,N_23484);
and U24174 (N_24174,N_22608,N_21130);
nand U24175 (N_24175,N_21476,N_23453);
or U24176 (N_24176,N_23882,N_22690);
and U24177 (N_24177,N_21952,N_23059);
nor U24178 (N_24178,N_21611,N_22041);
nand U24179 (N_24179,N_23427,N_21897);
or U24180 (N_24180,N_21071,N_22776);
nor U24181 (N_24181,N_22643,N_23659);
nor U24182 (N_24182,N_22231,N_21469);
and U24183 (N_24183,N_23717,N_22100);
or U24184 (N_24184,N_23394,N_23498);
and U24185 (N_24185,N_22856,N_23897);
and U24186 (N_24186,N_21657,N_23738);
nand U24187 (N_24187,N_21297,N_22416);
or U24188 (N_24188,N_22160,N_23268);
or U24189 (N_24189,N_21941,N_21594);
xor U24190 (N_24190,N_23477,N_22257);
xor U24191 (N_24191,N_21317,N_22994);
nor U24192 (N_24192,N_22347,N_23246);
nor U24193 (N_24193,N_22665,N_22258);
nand U24194 (N_24194,N_21370,N_23906);
or U24195 (N_24195,N_23553,N_21939);
nor U24196 (N_24196,N_22943,N_23705);
nand U24197 (N_24197,N_23092,N_23591);
and U24198 (N_24198,N_22986,N_21996);
xnor U24199 (N_24199,N_21212,N_23370);
nor U24200 (N_24200,N_22288,N_22098);
or U24201 (N_24201,N_22332,N_22652);
nor U24202 (N_24202,N_22497,N_22997);
or U24203 (N_24203,N_21174,N_23789);
nand U24204 (N_24204,N_22586,N_21468);
nor U24205 (N_24205,N_23886,N_22449);
or U24206 (N_24206,N_21871,N_23812);
nor U24207 (N_24207,N_21863,N_23214);
and U24208 (N_24208,N_22791,N_23556);
nand U24209 (N_24209,N_22933,N_22789);
and U24210 (N_24210,N_21211,N_23543);
nand U24211 (N_24211,N_21319,N_21138);
or U24212 (N_24212,N_22016,N_21511);
or U24213 (N_24213,N_23392,N_21607);
nor U24214 (N_24214,N_23133,N_23085);
nand U24215 (N_24215,N_23223,N_22397);
nand U24216 (N_24216,N_22383,N_22135);
or U24217 (N_24217,N_23359,N_21127);
nor U24218 (N_24218,N_23853,N_23777);
and U24219 (N_24219,N_21257,N_22189);
nor U24220 (N_24220,N_22045,N_21187);
or U24221 (N_24221,N_21745,N_21802);
nor U24222 (N_24222,N_21473,N_23207);
and U24223 (N_24223,N_21328,N_23783);
nand U24224 (N_24224,N_22754,N_22038);
and U24225 (N_24225,N_23974,N_22476);
nor U24226 (N_24226,N_21954,N_23208);
nor U24227 (N_24227,N_23441,N_21838);
nor U24228 (N_24228,N_22381,N_23618);
nor U24229 (N_24229,N_22199,N_21982);
or U24230 (N_24230,N_21960,N_23942);
nor U24231 (N_24231,N_21614,N_21290);
nand U24232 (N_24232,N_23376,N_21107);
nand U24233 (N_24233,N_22471,N_22174);
nor U24234 (N_24234,N_23501,N_23911);
nand U24235 (N_24235,N_22893,N_21205);
or U24236 (N_24236,N_22904,N_22206);
xnor U24237 (N_24237,N_21684,N_22223);
xor U24238 (N_24238,N_23623,N_22145);
xnor U24239 (N_24239,N_22807,N_21835);
and U24240 (N_24240,N_23767,N_22097);
or U24241 (N_24241,N_23880,N_22773);
nor U24242 (N_24242,N_23443,N_23209);
nor U24243 (N_24243,N_22085,N_22653);
xnor U24244 (N_24244,N_21475,N_21013);
xnor U24245 (N_24245,N_21740,N_21330);
and U24246 (N_24246,N_22902,N_23692);
or U24247 (N_24247,N_22102,N_23285);
or U24248 (N_24248,N_23933,N_21382);
nor U24249 (N_24249,N_22027,N_21208);
nor U24250 (N_24250,N_21972,N_23684);
and U24251 (N_24251,N_22539,N_23836);
or U24252 (N_24252,N_22615,N_21651);
nor U24253 (N_24253,N_22533,N_22908);
nor U24254 (N_24254,N_22047,N_21976);
nor U24255 (N_24255,N_22033,N_23081);
or U24256 (N_24256,N_23216,N_23288);
nor U24257 (N_24257,N_22729,N_21447);
nand U24258 (N_24258,N_22191,N_22443);
xnor U24259 (N_24259,N_22007,N_21818);
nor U24260 (N_24260,N_23331,N_22444);
nor U24261 (N_24261,N_23804,N_23787);
nor U24262 (N_24262,N_23098,N_23303);
xor U24263 (N_24263,N_21949,N_22682);
nand U24264 (N_24264,N_23309,N_23523);
nand U24265 (N_24265,N_21003,N_21153);
nand U24266 (N_24266,N_21336,N_21786);
and U24267 (N_24267,N_21008,N_21288);
nor U24268 (N_24268,N_23029,N_21980);
or U24269 (N_24269,N_23315,N_21995);
or U24270 (N_24270,N_22151,N_21673);
or U24271 (N_24271,N_22388,N_21460);
nor U24272 (N_24272,N_23938,N_21985);
or U24273 (N_24273,N_23439,N_21596);
xnor U24274 (N_24274,N_23130,N_23829);
nor U24275 (N_24275,N_21788,N_23721);
or U24276 (N_24276,N_23965,N_22068);
xor U24277 (N_24277,N_21712,N_21148);
nand U24278 (N_24278,N_22697,N_22741);
or U24279 (N_24279,N_21597,N_22295);
or U24280 (N_24280,N_22351,N_22107);
nor U24281 (N_24281,N_21419,N_21425);
and U24282 (N_24282,N_23631,N_21320);
xnor U24283 (N_24283,N_23302,N_21234);
xnor U24284 (N_24284,N_21877,N_23872);
and U24285 (N_24285,N_21046,N_22552);
nor U24286 (N_24286,N_23782,N_21694);
nand U24287 (N_24287,N_23551,N_21455);
xnor U24288 (N_24288,N_22275,N_22410);
nor U24289 (N_24289,N_22666,N_21958);
xnor U24290 (N_24290,N_23412,N_21801);
or U24291 (N_24291,N_23064,N_21201);
xor U24292 (N_24292,N_23521,N_22022);
or U24293 (N_24293,N_22506,N_21559);
nand U24294 (N_24294,N_22273,N_23226);
and U24295 (N_24295,N_21720,N_23637);
nand U24296 (N_24296,N_22942,N_21832);
and U24297 (N_24297,N_21791,N_23317);
or U24298 (N_24298,N_22324,N_23695);
nor U24299 (N_24299,N_22686,N_23778);
nor U24300 (N_24300,N_21303,N_22083);
nand U24301 (N_24301,N_23127,N_23825);
nand U24302 (N_24302,N_22891,N_21868);
nand U24303 (N_24303,N_22204,N_21457);
and U24304 (N_24304,N_21521,N_23496);
nor U24305 (N_24305,N_23327,N_21165);
nand U24306 (N_24306,N_21066,N_21151);
or U24307 (N_24307,N_21774,N_21096);
and U24308 (N_24308,N_21207,N_21817);
or U24309 (N_24309,N_23117,N_21747);
nor U24310 (N_24310,N_21374,N_22924);
or U24311 (N_24311,N_22600,N_23402);
and U24312 (N_24312,N_23487,N_22346);
nand U24313 (N_24313,N_23976,N_21617);
nor U24314 (N_24314,N_23816,N_22485);
or U24315 (N_24315,N_23750,N_23102);
nor U24316 (N_24316,N_22855,N_22106);
xor U24317 (N_24317,N_21302,N_22170);
nor U24318 (N_24318,N_22367,N_23368);
nor U24319 (N_24319,N_22502,N_21432);
nor U24320 (N_24320,N_21354,N_22453);
nor U24321 (N_24321,N_23557,N_22005);
or U24322 (N_24322,N_23364,N_23053);
nand U24323 (N_24323,N_21224,N_23611);
nand U24324 (N_24324,N_22228,N_21094);
nand U24325 (N_24325,N_21630,N_22363);
nand U24326 (N_24326,N_23374,N_21140);
nor U24327 (N_24327,N_22421,N_23526);
xnor U24328 (N_24328,N_23344,N_22664);
or U24329 (N_24329,N_22177,N_21493);
nor U24330 (N_24330,N_22760,N_21579);
nor U24331 (N_24331,N_23824,N_22121);
and U24332 (N_24332,N_21256,N_23740);
nor U24333 (N_24333,N_21272,N_23703);
nand U24334 (N_24334,N_22292,N_23701);
xor U24335 (N_24335,N_23055,N_22224);
nand U24336 (N_24336,N_21343,N_21190);
nand U24337 (N_24337,N_23462,N_22046);
xnor U24338 (N_24338,N_22601,N_21502);
nor U24339 (N_24339,N_23475,N_22836);
or U24340 (N_24340,N_21977,N_21989);
or U24341 (N_24341,N_22841,N_22863);
xnor U24342 (N_24342,N_21280,N_23702);
nand U24343 (N_24343,N_21668,N_22711);
nor U24344 (N_24344,N_21516,N_22463);
nor U24345 (N_24345,N_22165,N_22728);
nor U24346 (N_24346,N_22081,N_23167);
nor U24347 (N_24347,N_21576,N_22087);
xnor U24348 (N_24348,N_22757,N_22249);
xor U24349 (N_24349,N_23635,N_22373);
nand U24350 (N_24350,N_23419,N_23654);
nand U24351 (N_24351,N_23023,N_23379);
xnor U24352 (N_24352,N_23025,N_21371);
nand U24353 (N_24353,N_22372,N_23489);
nand U24354 (N_24354,N_23287,N_23384);
nand U24355 (N_24355,N_22409,N_21727);
xnor U24356 (N_24356,N_23067,N_21057);
and U24357 (N_24357,N_22521,N_23395);
xor U24358 (N_24358,N_22992,N_22451);
nand U24359 (N_24359,N_21679,N_22956);
xor U24360 (N_24360,N_23920,N_23554);
and U24361 (N_24361,N_21230,N_22202);
nand U24362 (N_24362,N_23253,N_21196);
nand U24363 (N_24363,N_21628,N_21811);
nand U24364 (N_24364,N_23114,N_22205);
xnor U24365 (N_24365,N_22470,N_21705);
nand U24366 (N_24366,N_21002,N_22217);
nor U24367 (N_24367,N_21333,N_21601);
or U24368 (N_24368,N_23464,N_22427);
nor U24369 (N_24369,N_23002,N_22417);
nand U24370 (N_24370,N_22528,N_21498);
xnor U24371 (N_24371,N_23347,N_22584);
or U24372 (N_24372,N_21087,N_21756);
and U24373 (N_24373,N_23390,N_23594);
nand U24374 (N_24374,N_22077,N_21191);
nor U24375 (N_24375,N_22458,N_22141);
and U24376 (N_24376,N_23885,N_21120);
xnor U24377 (N_24377,N_22338,N_21608);
or U24378 (N_24378,N_21427,N_22516);
or U24379 (N_24379,N_21881,N_23529);
nor U24380 (N_24380,N_23524,N_23837);
nand U24381 (N_24381,N_23694,N_21083);
xnor U24382 (N_24382,N_21658,N_23580);
nand U24383 (N_24383,N_22979,N_22423);
xor U24384 (N_24384,N_21324,N_22616);
nor U24385 (N_24385,N_21471,N_21037);
nand U24386 (N_24386,N_23575,N_22547);
nor U24387 (N_24387,N_23314,N_23731);
or U24388 (N_24388,N_21243,N_23902);
nor U24389 (N_24389,N_22704,N_22194);
or U24390 (N_24390,N_21014,N_22486);
nor U24391 (N_24391,N_22526,N_23726);
or U24392 (N_24392,N_22411,N_23517);
and U24393 (N_24393,N_21306,N_22163);
and U24394 (N_24394,N_23358,N_21592);
or U24395 (N_24395,N_21064,N_21344);
xnor U24396 (N_24396,N_21591,N_21278);
or U24397 (N_24397,N_23110,N_23768);
nand U24398 (N_24398,N_22559,N_21968);
and U24399 (N_24399,N_22700,N_23106);
and U24400 (N_24400,N_22520,N_23075);
or U24401 (N_24401,N_21392,N_21744);
and U24402 (N_24402,N_21132,N_22732);
xnor U24403 (N_24403,N_22819,N_21937);
nand U24404 (N_24404,N_22659,N_23918);
and U24405 (N_24405,N_21005,N_21925);
or U24406 (N_24406,N_23625,N_23345);
nand U24407 (N_24407,N_21730,N_23241);
or U24408 (N_24408,N_23381,N_22161);
xnor U24409 (N_24409,N_22009,N_23052);
or U24410 (N_24410,N_21346,N_21816);
nor U24411 (N_24411,N_23854,N_23951);
xor U24412 (N_24412,N_21569,N_23234);
or U24413 (N_24413,N_22091,N_22474);
nand U24414 (N_24414,N_21865,N_22598);
nor U24415 (N_24415,N_22857,N_22718);
nor U24416 (N_24416,N_23035,N_21259);
or U24417 (N_24417,N_23420,N_22642);
xor U24418 (N_24418,N_23995,N_21777);
or U24419 (N_24419,N_23282,N_21118);
nand U24420 (N_24420,N_22238,N_23447);
xnor U24421 (N_24421,N_21819,N_23168);
nor U24422 (N_24422,N_23332,N_23038);
nand U24423 (N_24423,N_23482,N_21047);
or U24424 (N_24424,N_22505,N_22264);
nand U24425 (N_24425,N_21307,N_22326);
or U24426 (N_24426,N_22299,N_21039);
or U24427 (N_24427,N_21728,N_23457);
or U24428 (N_24428,N_22529,N_22136);
xor U24429 (N_24429,N_22604,N_21115);
or U24430 (N_24430,N_21839,N_23217);
nor U24431 (N_24431,N_22320,N_23196);
nand U24432 (N_24432,N_21564,N_23434);
and U24433 (N_24433,N_21710,N_22256);
or U24434 (N_24434,N_23349,N_21965);
and U24435 (N_24435,N_23424,N_21683);
or U24436 (N_24436,N_22441,N_21397);
nor U24437 (N_24437,N_21035,N_21152);
and U24438 (N_24438,N_22276,N_21595);
nand U24439 (N_24439,N_21642,N_23186);
nand U24440 (N_24440,N_23539,N_22157);
xor U24441 (N_24441,N_21483,N_22011);
xor U24442 (N_24442,N_22437,N_23512);
xor U24443 (N_24443,N_21027,N_21154);
nor U24444 (N_24444,N_22574,N_21552);
or U24445 (N_24445,N_21680,N_21202);
xnor U24446 (N_24446,N_21634,N_23697);
nand U24447 (N_24447,N_23088,N_22852);
nor U24448 (N_24448,N_21856,N_21713);
xor U24449 (N_24449,N_22678,N_22051);
and U24450 (N_24450,N_22765,N_23629);
or U24451 (N_24451,N_23187,N_23009);
nor U24452 (N_24452,N_21536,N_22636);
xnor U24453 (N_24453,N_21102,N_22848);
or U24454 (N_24454,N_21301,N_23458);
nand U24455 (N_24455,N_21305,N_21737);
or U24456 (N_24456,N_21180,N_22607);
xor U24457 (N_24457,N_23572,N_22585);
xnor U24458 (N_24458,N_23972,N_23833);
xor U24459 (N_24459,N_21828,N_22960);
nor U24460 (N_24460,N_23990,N_22640);
or U24461 (N_24461,N_21329,N_23486);
or U24462 (N_24462,N_22294,N_21155);
nor U24463 (N_24463,N_21969,N_23875);
nor U24464 (N_24464,N_22104,N_23661);
and U24465 (N_24465,N_22823,N_22696);
nor U24466 (N_24466,N_21359,N_23259);
nand U24467 (N_24467,N_23389,N_23599);
or U24468 (N_24468,N_22001,N_22759);
or U24469 (N_24469,N_23982,N_22656);
nand U24470 (N_24470,N_23083,N_21540);
xor U24471 (N_24471,N_22507,N_23177);
nand U24472 (N_24472,N_23624,N_22748);
nor U24473 (N_24473,N_22727,N_23578);
or U24474 (N_24474,N_21189,N_22981);
xor U24475 (N_24475,N_23734,N_21133);
nand U24476 (N_24476,N_23154,N_23251);
and U24477 (N_24477,N_23733,N_23955);
xnor U24478 (N_24478,N_21616,N_22624);
nand U24479 (N_24479,N_23416,N_21771);
and U24480 (N_24480,N_22747,N_21736);
or U24481 (N_24481,N_22389,N_23870);
xnor U24482 (N_24482,N_21505,N_22579);
or U24483 (N_24483,N_23577,N_21702);
or U24484 (N_24484,N_22798,N_21365);
nand U24485 (N_24485,N_21990,N_21472);
and U24486 (N_24486,N_23776,N_22755);
or U24487 (N_24487,N_22824,N_23601);
nor U24488 (N_24488,N_21666,N_21076);
or U24489 (N_24489,N_21162,N_23536);
nor U24490 (N_24490,N_23842,N_22309);
or U24491 (N_24491,N_22610,N_23155);
nand U24492 (N_24492,N_21309,N_22813);
nor U24493 (N_24493,N_23109,N_22390);
and U24494 (N_24494,N_23744,N_22398);
and U24495 (N_24495,N_21955,N_21604);
xor U24496 (N_24496,N_22043,N_23463);
nor U24497 (N_24497,N_23538,N_21045);
or U24498 (N_24498,N_22334,N_21528);
nor U24499 (N_24499,N_22037,N_22255);
and U24500 (N_24500,N_21798,N_23131);
xnor U24501 (N_24501,N_21355,N_23054);
nor U24502 (N_24502,N_22095,N_22922);
xor U24503 (N_24503,N_21384,N_21519);
or U24504 (N_24504,N_22906,N_23164);
or U24505 (N_24505,N_22120,N_21255);
or U24506 (N_24506,N_21325,N_23794);
xnor U24507 (N_24507,N_22442,N_23311);
xor U24508 (N_24508,N_23820,N_21022);
and U24509 (N_24509,N_21646,N_22261);
nand U24510 (N_24510,N_22466,N_23939);
xor U24511 (N_24511,N_21911,N_21879);
and U24512 (N_24512,N_23921,N_23509);
or U24513 (N_24513,N_22681,N_22420);
nor U24514 (N_24514,N_23879,N_21246);
nor U24515 (N_24515,N_21993,N_23513);
nor U24516 (N_24516,N_21222,N_23022);
nand U24517 (N_24517,N_23707,N_23005);
nor U24518 (N_24518,N_23273,N_23915);
nand U24519 (N_24519,N_23683,N_21574);
nand U24520 (N_24520,N_22240,N_22879);
nor U24521 (N_24521,N_21599,N_21523);
nor U24522 (N_24522,N_22801,N_21349);
or U24523 (N_24523,N_22467,N_21743);
nor U24524 (N_24524,N_22302,N_22553);
nand U24525 (N_24525,N_21760,N_23989);
and U24526 (N_24526,N_21778,N_23569);
xnor U24527 (N_24527,N_23984,N_23438);
and U24528 (N_24528,N_21826,N_22265);
or U24529 (N_24529,N_22144,N_21010);
nand U24530 (N_24530,N_22072,N_21831);
and U24531 (N_24531,N_21407,N_22746);
or U24532 (N_24532,N_22564,N_22861);
or U24533 (N_24533,N_23604,N_21823);
nand U24534 (N_24534,N_21940,N_23082);
nor U24535 (N_24535,N_21978,N_23649);
and U24536 (N_24536,N_21665,N_22845);
nand U24537 (N_24537,N_21362,N_21936);
nor U24538 (N_24538,N_22784,N_22804);
and U24539 (N_24539,N_22418,N_22869);
or U24540 (N_24540,N_22393,N_23488);
nor U24541 (N_24541,N_22400,N_21888);
nand U24542 (N_24542,N_21409,N_23073);
nand U24543 (N_24543,N_23423,N_21933);
and U24544 (N_24544,N_22483,N_21950);
xnor U24545 (N_24545,N_23215,N_21411);
nor U24546 (N_24546,N_23375,N_22006);
xor U24547 (N_24547,N_21470,N_23564);
or U24548 (N_24548,N_23256,N_22262);
or U24549 (N_24549,N_22296,N_22839);
nand U24550 (N_24550,N_23432,N_22672);
nor U24551 (N_24551,N_22003,N_22129);
nor U24552 (N_24552,N_23095,N_22021);
nor U24553 (N_24553,N_22445,N_21268);
and U24554 (N_24554,N_21962,N_21386);
nand U24555 (N_24555,N_21412,N_22777);
or U24556 (N_24556,N_21814,N_21441);
nand U24557 (N_24557,N_22544,N_23238);
xor U24558 (N_24558,N_22307,N_23910);
or U24559 (N_24559,N_21088,N_23265);
or U24560 (N_24560,N_21291,N_22179);
xor U24561 (N_24561,N_22571,N_23722);
xnor U24562 (N_24562,N_23465,N_22012);
or U24563 (N_24563,N_21404,N_21629);
or U24564 (N_24564,N_21142,N_21807);
xnor U24565 (N_24565,N_21258,N_21220);
or U24566 (N_24566,N_22715,N_22980);
or U24567 (N_24567,N_21390,N_21810);
nor U24568 (N_24568,N_22768,N_21061);
and U24569 (N_24569,N_21492,N_21731);
nand U24570 (N_24570,N_21456,N_22779);
xnor U24571 (N_24571,N_21108,N_21285);
and U24572 (N_24572,N_22282,N_22318);
and U24573 (N_24573,N_23752,N_21275);
or U24574 (N_24574,N_21114,N_22775);
nor U24575 (N_24575,N_23953,N_22062);
nand U24576 (N_24576,N_21690,N_22403);
and U24577 (N_24577,N_22849,N_21091);
and U24578 (N_24578,N_21104,N_23118);
nor U24579 (N_24579,N_21261,N_21316);
xor U24580 (N_24580,N_22143,N_21714);
nor U24581 (N_24581,N_22701,N_21643);
and U24582 (N_24582,N_23987,N_23003);
nand U24583 (N_24583,N_21600,N_23665);
nor U24584 (N_24584,N_22251,N_22885);
and U24585 (N_24585,N_23149,N_22337);
and U24586 (N_24586,N_21159,N_21533);
nand U24587 (N_24587,N_21910,N_22243);
and U24588 (N_24588,N_22059,N_23105);
or U24589 (N_24589,N_23760,N_23510);
or U24590 (N_24590,N_21676,N_21697);
xor U24591 (N_24591,N_22064,N_23056);
and U24592 (N_24592,N_21837,N_21631);
nor U24593 (N_24593,N_23680,N_22996);
nand U24594 (N_24594,N_21992,N_22920);
nand U24595 (N_24595,N_23950,N_22031);
nor U24596 (N_24596,N_22492,N_22313);
and U24597 (N_24597,N_22984,N_22875);
nor U24598 (N_24598,N_21381,N_21474);
and U24599 (N_24599,N_21624,N_23552);
or U24600 (N_24600,N_22127,N_21466);
xor U24601 (N_24601,N_21675,N_23043);
or U24602 (N_24602,N_22510,N_21685);
nor U24603 (N_24603,N_21241,N_23986);
nand U24604 (N_24604,N_23240,N_22439);
and U24605 (N_24605,N_23664,N_21340);
xnor U24606 (N_24606,N_23868,N_21769);
or U24607 (N_24607,N_23363,N_21678);
nor U24608 (N_24608,N_23132,N_22030);
nor U24609 (N_24609,N_23729,N_22739);
xor U24610 (N_24610,N_21883,N_23180);
and U24611 (N_24611,N_21610,N_22220);
nand U24612 (N_24612,N_21249,N_21499);
nand U24613 (N_24613,N_21266,N_21418);
and U24614 (N_24614,N_22951,N_21636);
nor U24615 (N_24615,N_22219,N_21438);
nor U24616 (N_24616,N_23584,N_21613);
xnor U24617 (N_24617,N_21553,N_23080);
nor U24618 (N_24618,N_23235,N_22342);
or U24619 (N_24619,N_22926,N_22753);
nor U24620 (N_24620,N_21568,N_21700);
xnor U24621 (N_24621,N_21439,N_23795);
nor U24622 (N_24622,N_22685,N_22790);
xnor U24623 (N_24623,N_22961,N_23595);
nor U24624 (N_24624,N_23900,N_22691);
or U24625 (N_24625,N_22938,N_22212);
and U24626 (N_24626,N_21073,N_23630);
xor U24627 (N_24627,N_21721,N_22910);
xor U24628 (N_24628,N_22621,N_23473);
and U24629 (N_24629,N_21725,N_21231);
xnor U24630 (N_24630,N_23028,N_21517);
xnor U24631 (N_24631,N_22336,N_22310);
or U24632 (N_24632,N_21880,N_21075);
nor U24633 (N_24633,N_22982,N_23802);
nor U24634 (N_24634,N_22283,N_23296);
and U24635 (N_24635,N_23755,N_21376);
or U24636 (N_24636,N_22932,N_23706);
and U24637 (N_24637,N_23797,N_23188);
xnor U24638 (N_24638,N_22594,N_21669);
nor U24639 (N_24639,N_21416,N_22872);
xnor U24640 (N_24640,N_22867,N_23666);
or U24641 (N_24641,N_23924,N_22957);
and U24642 (N_24642,N_21844,N_22850);
nor U24643 (N_24643,N_23944,N_22490);
xnor U24644 (N_24644,N_22620,N_22658);
nor U24645 (N_24645,N_23646,N_23520);
and U24646 (N_24646,N_21247,N_23827);
or U24647 (N_24647,N_21805,N_23048);
and U24648 (N_24648,N_23060,N_22532);
nand U24649 (N_24649,N_21848,N_22568);
xnor U24650 (N_24650,N_21389,N_21000);
nor U24651 (N_24651,N_22499,N_21703);
or U24652 (N_24652,N_21855,N_22572);
and U24653 (N_24653,N_21920,N_23338);
xor U24654 (N_24654,N_21824,N_21792);
and U24655 (N_24655,N_22820,N_22683);
or U24656 (N_24656,N_21506,N_22424);
or U24657 (N_24657,N_23727,N_22774);
nand U24658 (N_24658,N_21749,N_23307);
nand U24659 (N_24659,N_23403,N_22569);
or U24660 (N_24660,N_23562,N_21185);
nor U24661 (N_24661,N_22415,N_21117);
xnor U24662 (N_24662,N_23001,N_23888);
xor U24663 (N_24663,N_23874,N_21387);
nand U24664 (N_24664,N_22844,N_21916);
nor U24665 (N_24665,N_23070,N_22040);
and U24666 (N_24666,N_21742,N_22725);
and U24667 (N_24667,N_21264,N_21776);
xor U24668 (N_24668,N_23627,N_22020);
and U24669 (N_24669,N_23817,N_22557);
nor U24670 (N_24670,N_21999,N_21139);
xor U24671 (N_24671,N_22232,N_22335);
xor U24672 (N_24672,N_23849,N_22540);
nand U24673 (N_24673,N_23045,N_22625);
nor U24674 (N_24674,N_22717,N_22178);
and U24675 (N_24675,N_23198,N_22786);
nand U24676 (N_24676,N_21069,N_22024);
and U24677 (N_24677,N_23641,N_22488);
nor U24678 (N_24678,N_22723,N_21874);
or U24679 (N_24679,N_23318,N_23563);
nor U24680 (N_24680,N_21524,N_21948);
nand U24681 (N_24681,N_22408,N_23507);
and U24682 (N_24682,N_21289,N_21223);
nand U24683 (N_24683,N_21254,N_21095);
nor U24684 (N_24684,N_23652,N_22052);
xor U24685 (N_24685,N_22661,N_23442);
or U24686 (N_24686,N_21175,N_21167);
and U24687 (N_24687,N_23306,N_21772);
xor U24688 (N_24688,N_22082,N_21030);
xnor U24689 (N_24689,N_23341,N_21902);
and U24690 (N_24690,N_21887,N_21467);
xor U24691 (N_24691,N_21361,N_22599);
nand U24692 (N_24692,N_21620,N_21262);
or U24693 (N_24693,N_23615,N_23495);
xor U24694 (N_24694,N_21512,N_23996);
or U24695 (N_24695,N_21105,N_21542);
or U24696 (N_24696,N_23254,N_22921);
xor U24697 (N_24697,N_23790,N_22673);
or U24698 (N_24698,N_21873,N_22646);
or U24699 (N_24699,N_23930,N_23689);
xnor U24700 (N_24700,N_23747,N_22010);
nand U24701 (N_24701,N_21462,N_22089);
nand U24702 (N_24702,N_22958,N_23826);
nor U24703 (N_24703,N_22382,N_22093);
nor U24704 (N_24704,N_21111,N_23062);
nand U24705 (N_24705,N_22237,N_21650);
and U24706 (N_24706,N_22073,N_21490);
nand U24707 (N_24707,N_23642,N_21358);
xor U24708 (N_24708,N_23848,N_23669);
or U24709 (N_24709,N_23985,N_21585);
nor U24710 (N_24710,N_23469,N_21043);
xor U24711 (N_24711,N_21011,N_22435);
nand U24712 (N_24712,N_22669,N_21753);
nand U24713 (N_24713,N_21766,N_22812);
xor U24714 (N_24714,N_23112,N_21313);
and U24715 (N_24715,N_22827,N_21098);
xnor U24716 (N_24716,N_23634,N_22384);
xnor U24717 (N_24717,N_21081,N_23231);
xor U24718 (N_24718,N_23156,N_22138);
nor U24719 (N_24719,N_23973,N_22025);
or U24720 (N_24720,N_22706,N_22260);
and U24721 (N_24721,N_23943,N_23753);
nand U24722 (N_24722,N_23894,N_22781);
nand U24723 (N_24723,N_22949,N_21351);
or U24724 (N_24724,N_23608,N_22802);
nor U24725 (N_24725,N_23770,N_21036);
nand U24726 (N_24726,N_21203,N_21975);
nand U24727 (N_24727,N_21785,N_23756);
and U24728 (N_24728,N_21007,N_21347);
xor U24729 (N_24729,N_23213,N_22361);
and U24730 (N_24730,N_23150,N_22154);
nand U24731 (N_24731,N_23676,N_21086);
or U24732 (N_24732,N_23039,N_22983);
xnor U24733 (N_24733,N_23619,N_21442);
and U24734 (N_24734,N_22985,N_21237);
xnor U24735 (N_24735,N_22339,N_21238);
and U24736 (N_24736,N_21161,N_23195);
nand U24737 (N_24737,N_22738,N_23862);
xnor U24738 (N_24738,N_21192,N_23798);
and U24739 (N_24739,N_21322,N_22617);
nor U24740 (N_24740,N_22851,N_21287);
and U24741 (N_24741,N_22912,N_21479);
xnor U24742 (N_24742,N_23143,N_21659);
or U24743 (N_24743,N_22758,N_21143);
and U24744 (N_24744,N_22894,N_21034);
and U24745 (N_24745,N_22889,N_21671);
nand U24746 (N_24746,N_21847,N_21050);
xor U24747 (N_24747,N_22563,N_22182);
or U24748 (N_24748,N_23772,N_23505);
or U24749 (N_24749,N_21198,N_21619);
nand U24750 (N_24750,N_22454,N_21644);
xnor U24751 (N_24751,N_21501,N_23565);
xor U24752 (N_24752,N_22993,N_22929);
nand U24753 (N_24753,N_23674,N_21757);
nand U24754 (N_24754,N_22482,N_23405);
and U24755 (N_24755,N_23454,N_22362);
nand U24756 (N_24756,N_22484,N_22555);
and U24757 (N_24757,N_23971,N_21953);
xnor U24758 (N_24758,N_21944,N_23793);
xor U24759 (N_24759,N_21841,N_23881);
nor U24760 (N_24760,N_23515,N_21567);
xor U24761 (N_24761,N_23945,N_21375);
xor U24762 (N_24762,N_22580,N_22468);
nor U24763 (N_24763,N_23650,N_22130);
xor U24764 (N_24764,N_22917,N_23528);
or U24765 (N_24765,N_22525,N_22687);
xor U24766 (N_24766,N_21327,N_22822);
and U24767 (N_24767,N_23710,N_22013);
or U24768 (N_24768,N_22806,N_21221);
and U24769 (N_24769,N_21751,N_23113);
xnor U24770 (N_24770,N_23284,N_23323);
xor U24771 (N_24771,N_22173,N_21924);
nor U24772 (N_24772,N_22816,N_22501);
and U24773 (N_24773,N_23571,N_23139);
or U24774 (N_24774,N_21226,N_22749);
nand U24775 (N_24775,N_21544,N_23981);
or U24776 (N_24776,N_23249,N_23247);
or U24777 (N_24777,N_23573,N_21674);
xor U24778 (N_24778,N_21571,N_23161);
and U24779 (N_24779,N_21729,N_23479);
nand U24780 (N_24780,N_21413,N_22180);
and U24781 (N_24781,N_23034,N_23440);
or U24782 (N_24782,N_21891,N_23103);
nand U24783 (N_24783,N_22436,N_23191);
or U24784 (N_24784,N_21182,N_23283);
xnor U24785 (N_24785,N_22137,N_21062);
and U24786 (N_24786,N_22379,N_21093);
or U24787 (N_24787,N_22976,N_21637);
nand U24788 (N_24788,N_23437,N_23061);
xor U24789 (N_24789,N_22562,N_21172);
nor U24790 (N_24790,N_22268,N_23409);
and U24791 (N_24791,N_23651,N_22050);
nor U24792 (N_24792,N_22392,N_23018);
nor U24793 (N_24793,N_23602,N_23638);
and U24794 (N_24794,N_21210,N_22710);
nor U24795 (N_24795,N_22211,N_22056);
or U24796 (N_24796,N_22782,N_21923);
or U24797 (N_24797,N_23398,N_21465);
or U24798 (N_24798,N_22152,N_21926);
and U24799 (N_24799,N_23550,N_21739);
or U24800 (N_24800,N_22783,N_22892);
nor U24801 (N_24801,N_23506,N_23585);
and U24802 (N_24802,N_21912,N_23352);
xor U24803 (N_24803,N_22811,N_23983);
nand U24804 (N_24804,N_21752,N_22195);
xnor U24805 (N_24805,N_22500,N_23596);
xor U24806 (N_24806,N_22900,N_23534);
nand U24807 (N_24807,N_23301,N_21846);
or U24808 (N_24808,N_23751,N_22937);
or U24809 (N_24809,N_22431,N_22124);
nand U24810 (N_24810,N_21006,N_23754);
nor U24811 (N_24811,N_21718,N_22327);
nand U24812 (N_24812,N_21686,N_23322);
nor U24813 (N_24813,N_22355,N_22042);
nor U24814 (N_24814,N_23124,N_22277);
nor U24815 (N_24815,N_21558,N_23091);
nand U24816 (N_24816,N_22438,N_21168);
and U24817 (N_24817,N_21463,N_22865);
nand U24818 (N_24818,N_22450,N_22133);
and U24819 (N_24819,N_21641,N_23835);
nand U24820 (N_24820,N_23286,N_23590);
or U24821 (N_24821,N_21905,N_22419);
xnor U24822 (N_24822,N_23518,N_22015);
and U24823 (N_24823,N_21144,N_23144);
xor U24824 (N_24824,N_21586,N_23620);
and U24825 (N_24825,N_23540,N_22060);
or U24826 (N_24826,N_22495,N_22099);
xnor U24827 (N_24827,N_22187,N_21973);
or U24828 (N_24828,N_22764,N_21378);
nor U24829 (N_24829,N_22939,N_23558);
nor U24830 (N_24830,N_22649,N_21200);
nor U24831 (N_24831,N_23116,N_22058);
xor U24832 (N_24832,N_22794,N_23769);
nand U24833 (N_24833,N_21489,N_22216);
and U24834 (N_24834,N_21761,N_21089);
nand U24835 (N_24835,N_23237,N_23176);
xor U24836 (N_24836,N_23739,N_22944);
xor U24837 (N_24837,N_23138,N_21783);
and U24838 (N_24838,N_23609,N_22530);
and U24839 (N_24839,N_22428,N_23011);
xor U24840 (N_24840,N_23800,N_23929);
and U24841 (N_24841,N_22800,N_23019);
nor U24842 (N_24842,N_21486,N_22554);
nor U24843 (N_24843,N_23422,N_21461);
nand U24844 (N_24844,N_23531,N_21827);
nand U24845 (N_24845,N_22167,N_21163);
nand U24846 (N_24846,N_23895,N_21907);
xnor U24847 (N_24847,N_22511,N_21687);
and U24848 (N_24848,N_23391,N_23430);
nand U24849 (N_24849,N_21452,N_23964);
xnor U24850 (N_24850,N_21399,N_21429);
or U24851 (N_24851,N_21947,N_22628);
and U24852 (N_24852,N_23941,N_21001);
nand U24853 (N_24853,N_23356,N_22541);
and U24854 (N_24854,N_21787,N_23763);
and U24855 (N_24855,N_21882,N_23732);
or U24856 (N_24856,N_23956,N_22542);
xnor U24857 (N_24857,N_23162,N_22266);
and U24858 (N_24858,N_22234,N_22475);
or U24859 (N_24859,N_22829,N_21793);
nor U24860 (N_24860,N_22066,N_22583);
or U24861 (N_24861,N_21251,N_22805);
nor U24862 (N_24862,N_23784,N_23975);
and U24863 (N_24863,N_21794,N_22724);
nand U24864 (N_24864,N_23086,N_23101);
and U24865 (N_24865,N_22662,N_23451);
nor U24866 (N_24866,N_22660,N_23847);
nand U24867 (N_24867,N_21032,N_21260);
nor U24868 (N_24868,N_22250,N_21711);
xnor U24869 (N_24869,N_22965,N_23262);
xnor U24870 (N_24870,N_21551,N_22969);
nand U24871 (N_24871,N_23699,N_23735);
or U24872 (N_24872,N_23193,N_22638);
nor U24873 (N_24873,N_22828,N_22328);
and U24874 (N_24874,N_22053,N_23917);
nor U24875 (N_24875,N_21830,N_23004);
nand U24876 (N_24876,N_22931,N_21055);
and U24877 (N_24877,N_22345,N_22535);
nand U24878 (N_24878,N_21799,N_22070);
nor U24879 (N_24879,N_21253,N_21672);
nand U24880 (N_24880,N_23855,N_23290);
and U24881 (N_24881,N_21146,N_22606);
nand U24882 (N_24882,N_23786,N_23470);
and U24883 (N_24883,N_23295,N_21341);
xnor U24884 (N_24884,N_21178,N_22004);
nand U24885 (N_24885,N_21136,N_21633);
or U24886 (N_24886,N_21556,N_22990);
nor U24887 (N_24887,N_23997,N_22487);
and U24888 (N_24888,N_21451,N_22633);
and U24889 (N_24889,N_23931,N_21885);
nor U24890 (N_24890,N_22826,N_23858);
nor U24891 (N_24891,N_23401,N_21878);
xnor U24892 (N_24892,N_22925,N_22637);
xor U24893 (N_24893,N_22166,N_21077);
xor U24894 (N_24894,N_23583,N_21775);
and U24895 (N_24895,N_22731,N_22110);
xor U24896 (N_24896,N_23065,N_23170);
and U24897 (N_24897,N_23169,N_22132);
xor U24898 (N_24898,N_23174,N_22103);
nand U24899 (N_24899,N_22792,N_23988);
nand U24900 (N_24900,N_21534,N_22903);
xnor U24901 (N_24901,N_21446,N_22873);
or U24902 (N_24902,N_21692,N_22709);
or U24903 (N_24903,N_23645,N_22695);
nor U24904 (N_24904,N_22831,N_23946);
nand U24905 (N_24905,N_21746,N_21545);
nand U24906 (N_24906,N_21510,N_23525);
xnor U24907 (N_24907,N_21415,N_22375);
and U24908 (N_24908,N_21918,N_22634);
nand U24909 (N_24909,N_23230,N_21408);
or U24910 (N_24910,N_21875,N_21377);
and U24911 (N_24911,N_22699,N_21895);
or U24912 (N_24912,N_23480,N_22737);
nand U24913 (N_24913,N_23407,N_23730);
or U24914 (N_24914,N_21584,N_22192);
nand U24915 (N_24915,N_21183,N_22329);
nand U24916 (N_24916,N_21368,N_21548);
nand U24917 (N_24917,N_23452,N_21276);
xor U24918 (N_24918,N_23272,N_21218);
nor U24919 (N_24919,N_23876,N_21400);
nand U24920 (N_24920,N_22884,N_23494);
and U24921 (N_24921,N_23968,N_21508);
xnor U24922 (N_24922,N_23743,N_23502);
and U24923 (N_24923,N_21529,N_23663);
nand U24924 (N_24924,N_22227,N_22870);
xor U24925 (N_24925,N_22139,N_21312);
nor U24926 (N_24926,N_21981,N_23757);
nand U24927 (N_24927,N_23828,N_23716);
and U24928 (N_24928,N_21424,N_23239);
and U24929 (N_24929,N_21209,N_23712);
and U24930 (N_24930,N_21054,N_22172);
nor U24931 (N_24931,N_23903,N_21695);
nor U24932 (N_24932,N_21428,N_22622);
nor U24933 (N_24933,N_23588,N_21292);
xor U24934 (N_24934,N_23163,N_22378);
xor U24935 (N_24935,N_22750,N_22648);
or U24936 (N_24936,N_23998,N_23366);
xnor U24937 (N_24937,N_23688,N_23310);
xnor U24938 (N_24938,N_22076,N_22119);
nand U24939 (N_24939,N_23818,N_21458);
nand U24940 (N_24940,N_21945,N_21507);
nand U24941 (N_24941,N_23202,N_22835);
nor U24942 (N_24942,N_23406,N_22055);
or U24943 (N_24943,N_21963,N_23255);
nor U24944 (N_24944,N_23511,N_22623);
xnor U24945 (N_24945,N_21348,N_23497);
or U24946 (N_24946,N_21956,N_21706);
nand U24947 (N_24947,N_21663,N_23994);
nor U24948 (N_24948,N_22842,N_22962);
nand U24949 (N_24949,N_23926,N_21497);
and U24950 (N_24950,N_23775,N_23728);
or U24951 (N_24951,N_23040,N_21334);
nor U24952 (N_24952,N_21129,N_23936);
nand U24953 (N_24953,N_22374,N_23681);
nand U24954 (N_24954,N_22494,N_23339);
xor U24955 (N_24955,N_21021,N_22522);
nand U24956 (N_24956,N_22146,N_22817);
nor U24957 (N_24957,N_23709,N_21866);
or U24958 (N_24958,N_21784,N_22360);
xnor U24959 (N_24959,N_23937,N_22577);
nor U24960 (N_24960,N_21137,N_23159);
or U24961 (N_24961,N_22975,N_22803);
and U24962 (N_24962,N_21150,N_23806);
or U24963 (N_24963,N_22858,N_23957);
nor U24964 (N_24964,N_22159,N_22694);
xor U24965 (N_24965,N_23428,N_22676);
or U24966 (N_24966,N_22057,N_23884);
xor U24967 (N_24967,N_21974,N_23838);
nor U24968 (N_24968,N_23503,N_21495);
and U24969 (N_24969,N_23218,N_21704);
nor U24970 (N_24970,N_21126,N_23773);
xor U24971 (N_24971,N_22635,N_21197);
and U24972 (N_24972,N_22998,N_23232);
and U24973 (N_24973,N_21065,N_21562);
or U24974 (N_24974,N_22744,N_23445);
or U24975 (N_24975,N_22928,N_21025);
and U24976 (N_24976,N_22291,N_23411);
or U24977 (N_24977,N_21225,N_23456);
and U24978 (N_24978,N_21696,N_22899);
or U24979 (N_24979,N_22200,N_21967);
and U24980 (N_24980,N_21635,N_22742);
nor U24981 (N_24981,N_21195,N_23030);
or U24982 (N_24982,N_21609,N_21899);
nand U24983 (N_24983,N_23136,N_21273);
nor U24984 (N_24984,N_22650,N_22245);
xor U24985 (N_24985,N_23928,N_22126);
xnor U24986 (N_24986,N_21602,N_21141);
xor U24987 (N_24987,N_23033,N_23087);
and U24988 (N_24988,N_21547,N_22825);
nor U24989 (N_24989,N_23300,N_21796);
nor U24990 (N_24990,N_23397,N_22496);
nand U24991 (N_24991,N_22550,N_22399);
xnor U24992 (N_24992,N_23178,N_23657);
nor U24993 (N_24993,N_21716,N_21563);
xnor U24994 (N_24994,N_23046,N_22425);
nor U24995 (N_24995,N_23324,N_22675);
xor U24996 (N_24996,N_23745,N_22193);
and U24997 (N_24997,N_21323,N_22221);
and U24998 (N_24998,N_21901,N_21857);
or U24999 (N_24999,N_23145,N_21979);
and U25000 (N_25000,N_23227,N_22088);
nor U25001 (N_25001,N_22702,N_21812);
or U25002 (N_25002,N_21085,N_21915);
and U25003 (N_25003,N_22190,N_21833);
nor U25004 (N_25004,N_22670,N_21332);
nor U25005 (N_25005,N_21577,N_21339);
nor U25006 (N_25006,N_23980,N_23134);
and U25007 (N_25007,N_23522,N_22655);
xor U25008 (N_25008,N_23948,N_23467);
and U25009 (N_25009,N_23715,N_21023);
and U25010 (N_25010,N_23026,N_23758);
nor U25011 (N_25011,N_22140,N_22349);
and U25012 (N_25012,N_21723,N_23612);
xnor U25013 (N_25013,N_23068,N_22797);
nand U25014 (N_25014,N_21090,N_23173);
nand U25015 (N_25015,N_22248,N_23741);
or U25016 (N_25016,N_22253,N_21147);
nand U25017 (N_25017,N_23077,N_23644);
or U25018 (N_25018,N_23561,N_23013);
xor U25019 (N_25019,N_22647,N_23653);
or U25020 (N_25020,N_22498,N_22815);
nor U25021 (N_25021,N_22396,N_21621);
or U25022 (N_25022,N_22565,N_23963);
xnor U25023 (N_25023,N_21158,N_22344);
nand U25024 (N_25024,N_23668,N_21765);
and U25025 (N_25025,N_23421,N_23736);
nand U25026 (N_25026,N_22284,N_22235);
xor U25027 (N_25027,N_21698,N_21284);
nor U25028 (N_25028,N_23333,N_22538);
or U25029 (N_25029,N_22799,N_22548);
and U25030 (N_25030,N_22988,N_22114);
xnor U25031 (N_25031,N_23660,N_21581);
nand U25032 (N_25032,N_21522,N_21194);
nand U25033 (N_25033,N_22740,N_22534);
xnor U25034 (N_25034,N_21110,N_21653);
nor U25035 (N_25035,N_22280,N_22846);
or U25036 (N_25036,N_23530,N_21681);
nor U25037 (N_25037,N_21527,N_23090);
and U25038 (N_25038,N_22208,N_23404);
xor U25039 (N_25039,N_23819,N_21767);
nor U25040 (N_25040,N_23151,N_22874);
nor U25041 (N_25041,N_23377,N_22353);
nor U25042 (N_25042,N_22589,N_22592);
or U25043 (N_25043,N_22171,N_23122);
xor U25044 (N_25044,N_23050,N_22069);
xnor U25045 (N_25045,N_22543,N_21656);
xor U25046 (N_25046,N_23481,N_22229);
xnor U25047 (N_25047,N_22860,N_21821);
or U25048 (N_25048,N_21131,N_22366);
nand U25049 (N_25049,N_22181,N_22259);
nor U25050 (N_25050,N_21250,N_23570);
or U25051 (N_25051,N_23166,N_23714);
nand U25052 (N_25052,N_22605,N_21164);
or U25053 (N_25053,N_22019,N_23566);
xor U25054 (N_25054,N_22707,N_21267);
xnor U25055 (N_25055,N_22385,N_22406);
nand U25056 (N_25056,N_22588,N_22570);
or U25057 (N_25057,N_23999,N_21606);
and U25058 (N_25058,N_21732,N_23711);
nand U25059 (N_25059,N_21688,N_23672);
or U25060 (N_25060,N_23365,N_23811);
or U25061 (N_25061,N_22478,N_22226);
or U25062 (N_25062,N_22218,N_21627);
xor U25063 (N_25063,N_21800,N_21931);
nor U25064 (N_25064,N_21060,N_22198);
nand U25065 (N_25065,N_23516,N_21070);
xnor U25066 (N_25066,N_21537,N_23640);
xor U25067 (N_25067,N_21986,N_21640);
xor U25068 (N_25068,N_23275,N_23774);
or U25069 (N_25069,N_23846,N_22657);
and U25070 (N_25070,N_23326,N_23628);
xnor U25071 (N_25071,N_21896,N_22911);
or U25072 (N_25072,N_21724,N_23568);
or U25073 (N_25073,N_21770,N_21849);
nor U25074 (N_25074,N_21942,N_21546);
nor U25075 (N_25075,N_21119,N_22566);
nand U25076 (N_25076,N_22297,N_23372);
xnor U25077 (N_25077,N_22306,N_21099);
or U25078 (N_25078,N_21829,N_22434);
or U25079 (N_25079,N_23724,N_23670);
nor U25080 (N_25080,N_22096,N_22745);
or U25081 (N_25081,N_23527,N_22733);
nor U25082 (N_25082,N_23316,N_22519);
nand U25083 (N_25083,N_21080,N_23194);
nand U25084 (N_25084,N_22279,N_23499);
nor U25085 (N_25085,N_22945,N_22974);
and U25086 (N_25086,N_23904,N_22882);
xor U25087 (N_25087,N_21228,N_23115);
nand U25088 (N_25088,N_22331,N_21876);
xor U25089 (N_25089,N_23104,N_22905);
xnor U25090 (N_25090,N_21898,N_22469);
nor U25091 (N_25091,N_21277,N_22343);
or U25092 (N_25092,N_21177,N_23190);
xor U25093 (N_25093,N_23328,N_23276);
nand U25094 (N_25094,N_23222,N_23291);
xnor U25095 (N_25095,N_22214,N_23107);
xnor U25096 (N_25096,N_22185,N_23492);
xnor U25097 (N_25097,N_23089,N_23245);
and U25098 (N_25098,N_23100,N_21754);
xnor U25099 (N_25099,N_22793,N_21113);
or U25100 (N_25100,N_21430,N_21478);
nor U25101 (N_25101,N_21049,N_21892);
nand U25102 (N_25102,N_22808,N_21759);
nor U25103 (N_25103,N_23840,N_23908);
nand U25104 (N_25104,N_21820,N_23841);
nor U25105 (N_25105,N_23761,N_23647);
nor U25106 (N_25106,N_21233,N_21009);
or U25107 (N_25107,N_21598,N_23044);
nor U25108 (N_25108,N_21248,N_22281);
nor U25109 (N_25109,N_22558,N_23546);
nor U25110 (N_25110,N_22473,N_23555);
or U25111 (N_25111,N_22222,N_23224);
nor U25112 (N_25112,N_22573,N_23399);
nor U25113 (N_25113,N_22896,N_21227);
nand U25114 (N_25114,N_23094,N_21431);
or U25115 (N_25115,N_23471,N_23803);
and U25116 (N_25116,N_21367,N_22972);
nand U25117 (N_25117,N_21160,N_21638);
or U25118 (N_25118,N_22560,N_23182);
xor U25119 (N_25119,N_23417,N_21913);
nand U25120 (N_25120,N_23913,N_23582);
nand U25121 (N_25121,N_22602,N_22721);
xnor U25122 (N_25122,N_22609,N_22341);
nand U25123 (N_25123,N_22853,N_21851);
nor U25124 (N_25124,N_22446,N_21414);
nor U25125 (N_25125,N_23426,N_22412);
or U25126 (N_25126,N_23597,N_21488);
nand U25127 (N_25127,N_23852,N_21112);
nand U25128 (N_25128,N_23342,N_23899);
nand U25129 (N_25129,N_22886,N_23289);
nor U25130 (N_25130,N_21813,N_22462);
nand U25131 (N_25131,N_23725,N_21242);
and U25132 (N_25132,N_21957,N_21645);
or U25133 (N_25133,N_22278,N_22883);
or U25134 (N_25134,N_22394,N_21735);
or U25135 (N_25135,N_21722,N_22995);
nand U25136 (N_25136,N_23148,N_21491);
or U25137 (N_25137,N_23682,N_23431);
nand U25138 (N_25138,N_23863,N_22591);
nor U25139 (N_25139,N_22125,N_22036);
xor U25140 (N_25140,N_23058,N_21421);
or U25141 (N_25141,N_22430,N_22612);
and U25142 (N_25142,N_23491,N_23779);
and U25143 (N_25143,N_22184,N_21961);
nand U25144 (N_25144,N_23378,N_23959);
xor U25145 (N_25145,N_23823,N_21717);
nand U25146 (N_25146,N_23337,N_23206);
and U25147 (N_25147,N_21843,N_21125);
or U25148 (N_25148,N_21444,N_21998);
or U25149 (N_25149,N_22480,N_21363);
and U25150 (N_25150,N_23076,N_22368);
nor U25151 (N_25151,N_22726,N_23560);
and U25152 (N_25152,N_21935,N_23771);
and U25153 (N_25153,N_22092,N_21648);
nand U25154 (N_25154,N_23413,N_21578);
or U25155 (N_25155,N_21240,N_22935);
and U25156 (N_25156,N_23330,N_22183);
nand U25157 (N_25157,N_23746,N_22671);
xor U25158 (N_25158,N_23476,N_22626);
and U25159 (N_25159,N_22402,N_21500);
nand U25160 (N_25160,N_23687,N_22762);
nor U25161 (N_25161,N_22298,N_21145);
and U25162 (N_25162,N_23704,N_23093);
xor U25163 (N_25163,N_21443,N_21664);
and U25164 (N_25164,N_22531,N_21509);
or U25165 (N_25165,N_21904,N_23839);
xnor U25166 (N_25166,N_22155,N_23883);
nand U25167 (N_25167,N_23459,N_22340);
and U25168 (N_25168,N_23415,N_21315);
or U25169 (N_25169,N_22769,N_21701);
and U25170 (N_25170,N_23270,N_22148);
xor U25171 (N_25171,N_23172,N_22244);
xnor U25172 (N_25172,N_22639,N_22391);
xnor U25173 (N_25173,N_22210,N_23871);
and U25174 (N_25174,N_23007,N_22233);
xor U25175 (N_25175,N_23414,N_21886);
nor U25176 (N_25176,N_22854,N_21321);
or U25177 (N_25177,N_21217,N_21889);
and U25178 (N_25178,N_21514,N_22630);
and U25179 (N_25179,N_21345,N_22188);
nor U25180 (N_25180,N_21667,N_23867);
nand U25181 (N_25181,N_21423,N_22272);
and U25182 (N_25182,N_23444,N_23006);
nor U25183 (N_25183,N_23436,N_22314);
xnor U25184 (N_25184,N_23141,N_21632);
and U25185 (N_25185,N_23764,N_22176);
nand U25186 (N_25186,N_23859,N_21395);
xnor U25187 (N_25187,N_21048,N_22714);
nor U25188 (N_25188,N_21804,N_21040);
nor U25189 (N_25189,N_22479,N_21795);
nand U25190 (N_25190,N_22230,N_22880);
and U25191 (N_25191,N_22627,N_23146);
and U25192 (N_25192,N_21373,N_23220);
or U25193 (N_25193,N_22413,N_23504);
nand U25194 (N_25194,N_22941,N_23263);
nand U25195 (N_25195,N_21236,N_23713);
xnor U25196 (N_25196,N_21682,N_22269);
and U25197 (N_25197,N_21406,N_23605);
xnor U25198 (N_25198,N_21789,N_22074);
and U25199 (N_25199,N_22207,N_21921);
nand U25200 (N_25200,N_23111,N_22465);
xnor U25201 (N_25201,N_23184,N_23935);
nor U25202 (N_25202,N_21004,N_22371);
and U25203 (N_25203,N_23807,N_21372);
nor U25204 (N_25204,N_22618,N_22115);
and U25205 (N_25205,N_23947,N_23861);
nor U25206 (N_25206,N_22304,N_22252);
xnor U25207 (N_25207,N_21782,N_21464);
nor U25208 (N_25208,N_21983,N_23014);
or U25209 (N_25209,N_21169,N_21214);
and U25210 (N_25210,N_22549,N_23271);
nor U25211 (N_25211,N_22401,N_21265);
xnor U25212 (N_25212,N_22832,N_23266);
xnor U25213 (N_25213,N_21215,N_22404);
or U25214 (N_25214,N_23696,N_22837);
nand U25215 (N_25215,N_22301,N_21453);
and U25216 (N_25216,N_21790,N_22354);
xor U25217 (N_25217,N_22934,N_22319);
nor U25218 (N_25218,N_23533,N_22877);
xor U25219 (N_25219,N_23099,N_21449);
nand U25220 (N_25220,N_23388,N_21994);
xor U25221 (N_25221,N_22838,N_23157);
nor U25222 (N_25222,N_21128,N_21100);
and U25223 (N_25223,N_21282,N_22595);
xor U25224 (N_25224,N_22414,N_21420);
or U25225 (N_25225,N_23545,N_22743);
and U25226 (N_25226,N_21020,N_22876);
xor U25227 (N_25227,N_22916,N_22308);
xor U25228 (N_25228,N_22785,N_21626);
nand U25229 (N_25229,N_23788,N_21909);
or U25230 (N_25230,N_22668,N_21861);
or U25231 (N_25231,N_22587,N_21518);
and U25232 (N_25232,N_22014,N_22405);
or U25233 (N_25233,N_22909,N_22578);
and U25234 (N_25234,N_22840,N_23607);
xnor U25235 (N_25235,N_23648,N_21575);
and U25236 (N_25236,N_22365,N_23822);
or U25237 (N_25237,N_22898,N_22175);
or U25238 (N_25238,N_21436,N_21661);
xnor U25239 (N_25239,N_23923,N_22377);
or U25240 (N_25240,N_23221,N_22356);
or U25241 (N_25241,N_21525,N_21082);
nor U25242 (N_25242,N_23063,N_23257);
and U25243 (N_25243,N_22049,N_21919);
or U25244 (N_25244,N_23297,N_22897);
xor U25245 (N_25245,N_21216,N_21515);
nor U25246 (N_25246,N_21670,N_21012);
xor U25247 (N_25247,N_23274,N_22386);
nand U25248 (N_25248,N_23354,N_22090);
xnor U25249 (N_25249,N_23830,N_23478);
and U25250 (N_25250,N_22168,N_21738);
nor U25251 (N_25251,N_21239,N_23260);
or U25252 (N_25252,N_21530,N_23878);
xnor U25253 (N_25253,N_23780,N_23152);
xnor U25254 (N_25254,N_22756,N_23335);
and U25255 (N_25255,N_23866,N_23675);
nand U25256 (N_25256,N_23567,N_21173);
nor U25257 (N_25257,N_23386,N_23047);
xor U25258 (N_25258,N_21450,N_23396);
and U25259 (N_25259,N_21852,N_23057);
nor U25260 (N_25260,N_23017,N_21106);
or U25261 (N_25261,N_22477,N_23079);
nor U25262 (N_25262,N_22290,N_21171);
nor U25263 (N_25263,N_23765,N_21612);
and U25264 (N_25264,N_23204,N_22325);
nor U25265 (N_25265,N_22147,N_23233);
nand U25266 (N_25266,N_23032,N_23940);
nor U25267 (N_25267,N_23671,N_23893);
nand U25268 (N_25268,N_22963,N_23952);
and U25269 (N_25269,N_23850,N_22546);
xnor U25270 (N_25270,N_23796,N_21074);
and U25271 (N_25271,N_21029,N_21308);
nor U25272 (N_25272,N_23097,N_21494);
and U25273 (N_25273,N_21654,N_21072);
and U25274 (N_25274,N_21758,N_22871);
and U25275 (N_25275,N_23071,N_21028);
nand U25276 (N_25276,N_23203,N_23181);
and U25277 (N_25277,N_22517,N_23586);
and U25278 (N_25278,N_22919,N_21929);
or U25279 (N_25279,N_21298,N_21271);
and U25280 (N_25280,N_22162,N_21068);
nor U25281 (N_25281,N_21437,N_23598);
nand U25282 (N_25282,N_21310,N_21477);
xnor U25283 (N_25283,N_23978,N_22603);
nand U25284 (N_25284,N_21481,N_23639);
or U25285 (N_25285,N_21748,N_21134);
and U25286 (N_25286,N_23020,N_23225);
nand U25287 (N_25287,N_21987,N_21504);
and U25288 (N_25288,N_23387,N_21485);
xnor U25289 (N_25289,N_21279,N_23334);
and U25290 (N_25290,N_21019,N_22778);
xor U25291 (N_25291,N_21149,N_21850);
or U25292 (N_25292,N_23278,N_21618);
nand U25293 (N_25293,N_21084,N_21764);
nand U25294 (N_25294,N_22134,N_21033);
and U25295 (N_25295,N_21342,N_22834);
or U25296 (N_25296,N_21781,N_23809);
and U25297 (N_25297,N_21440,N_23371);
nand U25298 (N_25298,N_22567,N_22674);
nand U25299 (N_25299,N_22575,N_22667);
or U25300 (N_25300,N_23857,N_21398);
or U25301 (N_25301,N_23603,N_21293);
nor U25302 (N_25302,N_21647,N_23012);
or U25303 (N_25303,N_23015,N_22619);
or U25304 (N_25304,N_22895,N_23321);
xor U25305 (N_25305,N_22513,N_22881);
and U25306 (N_25306,N_23175,N_21281);
nand U25307 (N_25307,N_22771,N_23961);
and U25308 (N_25308,N_23066,N_23108);
and U25309 (N_25309,N_22868,N_22311);
nor U25310 (N_25310,N_23979,N_22370);
nor U25311 (N_25311,N_22322,N_22118);
nor U25312 (N_25312,N_23037,N_22923);
xnor U25313 (N_25313,N_23613,N_22429);
and U25314 (N_25314,N_22866,N_23541);
nand U25315 (N_25315,N_23010,N_23031);
or U25316 (N_25316,N_21715,N_22719);
or U25317 (N_25317,N_22913,N_22809);
or U25318 (N_25318,N_21893,N_21930);
nand U25319 (N_25319,N_21364,N_23312);
or U25320 (N_25320,N_22201,N_22663);
nor U25321 (N_25321,N_23383,N_22387);
or U25322 (N_25322,N_21709,N_21454);
or U25323 (N_25323,N_22491,N_22105);
nor U25324 (N_25324,N_23385,N_21836);
or U25325 (N_25325,N_22796,N_21860);
nand U25326 (N_25326,N_22950,N_21270);
or U25327 (N_25327,N_22536,N_21988);
xnor U25328 (N_25328,N_21964,N_22461);
or U25329 (N_25329,N_23078,N_22766);
nor U25330 (N_25330,N_23361,N_23992);
and U25331 (N_25331,N_22692,N_23016);
or U25332 (N_25332,N_23614,N_21726);
nand U25333 (N_25333,N_22156,N_22481);
and U25334 (N_25334,N_21252,N_22654);
nor U25335 (N_25335,N_22350,N_23158);
xor U25336 (N_25336,N_21707,N_23126);
nand U25337 (N_25337,N_22787,N_22357);
and U25338 (N_25338,N_22364,N_22080);
nand U25339 (N_25339,N_23351,N_22688);
xnor U25340 (N_25340,N_21360,N_21588);
nor U25341 (N_25341,N_21589,N_21295);
nor U25342 (N_25342,N_23749,N_22018);
nand U25343 (N_25343,N_21859,N_22614);
nand U25344 (N_25344,N_22330,N_21908);
nand U25345 (N_25345,N_23912,N_23021);
xnor U25346 (N_25346,N_23147,N_21480);
and U25347 (N_25347,N_22968,N_21052);
or U25348 (N_25348,N_21854,N_22078);
nand U25349 (N_25349,N_21041,N_21286);
xor U25350 (N_25350,N_22071,N_22464);
and U25351 (N_25351,N_21997,N_21652);
and U25352 (N_25352,N_21352,N_22693);
and U25353 (N_25353,N_23466,N_23865);
nand U25354 (N_25354,N_22613,N_23229);
nor U25355 (N_25355,N_22780,N_23723);
and U25356 (N_25356,N_22169,N_23305);
and U25357 (N_25357,N_21549,N_21353);
xor U25358 (N_25358,N_23737,N_22432);
nand U25359 (N_25359,N_23319,N_22023);
or U25360 (N_25360,N_21689,N_21934);
nand U25361 (N_25361,N_21526,N_22117);
nor U25362 (N_25362,N_23433,N_22054);
or U25363 (N_25363,N_23449,N_21733);
nor U25364 (N_25364,N_21539,N_22321);
and U25365 (N_25365,N_23264,N_22989);
nor U25366 (N_25366,N_23140,N_23072);
and U25367 (N_25367,N_23791,N_22503);
and U25368 (N_25368,N_22504,N_21051);
xor U25369 (N_25369,N_23304,N_21927);
xnor U25370 (N_25370,N_21176,N_23677);
and U25371 (N_25371,N_23719,N_22142);
and U25372 (N_25372,N_22597,N_21825);
xor U25373 (N_25373,N_22611,N_21296);
nor U25374 (N_25374,N_22000,N_21496);
or U25375 (N_25375,N_21135,N_23343);
and U25376 (N_25376,N_21894,N_21971);
and U25377 (N_25377,N_22236,N_22026);
and U25378 (N_25378,N_23027,N_23325);
and U25379 (N_25379,N_22821,N_22149);
xnor U25380 (N_25380,N_21410,N_21435);
nand U25381 (N_25381,N_21350,N_23348);
or U25382 (N_25382,N_22582,N_23393);
nand U25383 (N_25383,N_23425,N_21708);
and U25384 (N_25384,N_22515,N_23042);
xnor U25385 (N_25385,N_21283,N_21768);
and U25386 (N_25386,N_23446,N_23212);
xor U25387 (N_25387,N_21951,N_23686);
nand U25388 (N_25388,N_22847,N_23468);
or U25389 (N_25389,N_23891,N_23698);
or U25390 (N_25390,N_21938,N_21560);
or U25391 (N_25391,N_23367,N_21734);
nor U25392 (N_25392,N_23123,N_22285);
or U25393 (N_25393,N_23472,N_22289);
and U25394 (N_25394,N_22736,N_23299);
nor U25395 (N_25395,N_23693,N_22509);
xnor U25396 (N_25396,N_23228,N_23119);
xor U25397 (N_25397,N_23574,N_23621);
and U25398 (N_25398,N_21587,N_21750);
or U25399 (N_25399,N_21056,N_22131);
and U25400 (N_25400,N_22472,N_21922);
nand U25401 (N_25401,N_23508,N_21779);
nor U25402 (N_25402,N_22039,N_23142);
nand U25403 (N_25403,N_21623,N_23408);
nand U25404 (N_25404,N_23993,N_23244);
and U25405 (N_25405,N_22770,N_23815);
and U25406 (N_25406,N_23024,N_21338);
or U25407 (N_25407,N_22977,N_21396);
nor U25408 (N_25408,N_23656,N_21845);
nor U25409 (N_25409,N_22002,N_23036);
nor U25410 (N_25410,N_21603,N_21385);
and U25411 (N_25411,N_23049,N_21538);
nand U25412 (N_25412,N_22830,N_23592);
and U25413 (N_25413,N_21573,N_21755);
and U25414 (N_25414,N_21803,N_23179);
and U25415 (N_25415,N_22576,N_23373);
nor U25416 (N_25416,N_22448,N_23382);
xor U25417 (N_25417,N_22999,N_21318);
and U25418 (N_25418,N_23813,N_22954);
and U25419 (N_25419,N_22772,N_22991);
xor U25420 (N_25420,N_23258,N_22348);
nor U25421 (N_25421,N_21541,N_22267);
xor U25422 (N_25422,N_22795,N_23121);
or U25423 (N_25423,N_23460,N_22645);
nand U25424 (N_25424,N_22116,N_21625);
and U25425 (N_25425,N_21580,N_21867);
or U25426 (N_25426,N_22713,N_22556);
and U25427 (N_25427,N_22457,N_22936);
nor U25428 (N_25428,N_22407,N_23537);
nand U25429 (N_25429,N_22048,N_23927);
nor U25430 (N_25430,N_21122,N_21853);
xor U25431 (N_25431,N_23519,N_21554);
xnor U25432 (N_25432,N_21513,N_22079);
xnor U25433 (N_25433,N_22581,N_22196);
and U25434 (N_25434,N_21229,N_23357);
or U25435 (N_25435,N_22680,N_23261);
nor U25436 (N_25436,N_23210,N_22422);
xor U25437 (N_25437,N_22966,N_21097);
nand U25438 (N_25438,N_23243,N_21582);
nor U25439 (N_25439,N_23860,N_21109);
and U25440 (N_25440,N_22376,N_22814);
or U25441 (N_25441,N_23450,N_21572);
and U25442 (N_25442,N_22312,N_23643);
xor U25443 (N_25443,N_23277,N_21092);
nand U25444 (N_25444,N_22035,N_22101);
and U25445 (N_25445,N_23589,N_23962);
and U25446 (N_25446,N_21213,N_22316);
nand U25447 (N_25447,N_22512,N_21079);
nor U25448 (N_25448,N_22034,N_21188);
xnor U25449 (N_25449,N_23925,N_22722);
and U25450 (N_25450,N_22197,N_22967);
nand U25451 (N_25451,N_21059,N_21991);
xnor U25452 (N_25452,N_23901,N_21890);
nand U25453 (N_25453,N_22213,N_22915);
or U25454 (N_25454,N_23898,N_21566);
or U25455 (N_25455,N_22489,N_21741);
or U25456 (N_25456,N_23380,N_22241);
or U25457 (N_25457,N_22716,N_21294);
nor U25458 (N_25458,N_23500,N_22946);
nand U25459 (N_25459,N_23954,N_21914);
or U25460 (N_25460,N_22017,N_23205);
xnor U25461 (N_25461,N_23298,N_22859);
and U25462 (N_25462,N_23949,N_22545);
and U25463 (N_25463,N_21590,N_21834);
nand U25464 (N_25464,N_22086,N_23074);
xnor U25465 (N_25465,N_23353,N_22862);
xor U25466 (N_25466,N_21394,N_21299);
or U25467 (N_25467,N_22527,N_22940);
and U25468 (N_25468,N_21615,N_23250);
nor U25469 (N_25469,N_23362,N_22456);
and U25470 (N_25470,N_22907,N_21693);
nor U25471 (N_25471,N_22679,N_22730);
nand U25472 (N_25472,N_21900,N_22708);
or U25473 (N_25473,N_23069,N_21016);
or U25474 (N_25474,N_23667,N_21269);
nor U25475 (N_25475,N_23171,N_22843);
xor U25476 (N_25476,N_23606,N_23544);
or U25477 (N_25477,N_23967,N_21984);
xor U25478 (N_25478,N_22065,N_21063);
xor U25479 (N_25479,N_21445,N_21842);
and U25480 (N_25480,N_22888,N_21017);
nor U25481 (N_25481,N_23969,N_22514);
nor U25482 (N_25482,N_22122,N_23831);
or U25483 (N_25483,N_21101,N_23483);
or U25484 (N_25484,N_22426,N_23008);
and U25485 (N_25485,N_22953,N_23892);
or U25486 (N_25486,N_22369,N_21300);
xor U25487 (N_25487,N_22203,N_23355);
and U25488 (N_25488,N_21067,N_23616);
nand U25489 (N_25489,N_22254,N_21822);
xnor U25490 (N_25490,N_23051,N_21380);
or U25491 (N_25491,N_22493,N_23137);
nand U25492 (N_25492,N_22518,N_22712);
nor U25493 (N_25493,N_22447,N_22008);
nand U25494 (N_25494,N_22305,N_21503);
nor U25495 (N_25495,N_21862,N_23742);
nand U25496 (N_25496,N_21018,N_21157);
nor U25497 (N_25497,N_23856,N_23189);
nor U25498 (N_25498,N_22720,N_23673);
xor U25499 (N_25499,N_22629,N_23248);
and U25500 (N_25500,N_23436,N_23170);
and U25501 (N_25501,N_22203,N_23906);
or U25502 (N_25502,N_22304,N_21917);
xor U25503 (N_25503,N_23793,N_22375);
nand U25504 (N_25504,N_22903,N_22033);
nand U25505 (N_25505,N_23053,N_21112);
nor U25506 (N_25506,N_22395,N_22715);
nand U25507 (N_25507,N_21361,N_21358);
nor U25508 (N_25508,N_23664,N_23445);
nor U25509 (N_25509,N_23363,N_21754);
nor U25510 (N_25510,N_23854,N_22282);
nand U25511 (N_25511,N_22658,N_23025);
nand U25512 (N_25512,N_23054,N_22503);
or U25513 (N_25513,N_23779,N_22259);
nor U25514 (N_25514,N_23846,N_22404);
xor U25515 (N_25515,N_21952,N_21598);
and U25516 (N_25516,N_21706,N_21649);
nor U25517 (N_25517,N_22924,N_21377);
nand U25518 (N_25518,N_23262,N_22374);
or U25519 (N_25519,N_22652,N_21445);
xor U25520 (N_25520,N_23043,N_22928);
and U25521 (N_25521,N_23806,N_23492);
and U25522 (N_25522,N_22496,N_21311);
and U25523 (N_25523,N_21774,N_21755);
nor U25524 (N_25524,N_23411,N_22876);
and U25525 (N_25525,N_22567,N_21749);
nor U25526 (N_25526,N_23534,N_22454);
or U25527 (N_25527,N_22784,N_23205);
or U25528 (N_25528,N_23606,N_21126);
nand U25529 (N_25529,N_21421,N_23760);
and U25530 (N_25530,N_21447,N_23550);
and U25531 (N_25531,N_22977,N_23490);
nor U25532 (N_25532,N_23698,N_23621);
xnor U25533 (N_25533,N_21914,N_23619);
and U25534 (N_25534,N_21529,N_23980);
xnor U25535 (N_25535,N_22802,N_23188);
xnor U25536 (N_25536,N_23222,N_23294);
nor U25537 (N_25537,N_22159,N_21959);
xnor U25538 (N_25538,N_23954,N_22632);
and U25539 (N_25539,N_23548,N_22416);
nand U25540 (N_25540,N_21374,N_23227);
or U25541 (N_25541,N_22804,N_22604);
nand U25542 (N_25542,N_23002,N_21068);
xor U25543 (N_25543,N_22052,N_22623);
nand U25544 (N_25544,N_21909,N_21784);
nand U25545 (N_25545,N_23086,N_22297);
xnor U25546 (N_25546,N_22065,N_22784);
and U25547 (N_25547,N_21935,N_21291);
nor U25548 (N_25548,N_23544,N_21794);
or U25549 (N_25549,N_23808,N_22574);
nor U25550 (N_25550,N_22661,N_23262);
nand U25551 (N_25551,N_23919,N_23800);
nor U25552 (N_25552,N_22764,N_23085);
nand U25553 (N_25553,N_22844,N_22133);
xnor U25554 (N_25554,N_21636,N_23768);
nor U25555 (N_25555,N_21026,N_21839);
and U25556 (N_25556,N_23458,N_21246);
nand U25557 (N_25557,N_22884,N_23745);
nor U25558 (N_25558,N_21626,N_21842);
nand U25559 (N_25559,N_21425,N_22980);
nand U25560 (N_25560,N_22721,N_23179);
and U25561 (N_25561,N_22104,N_23202);
and U25562 (N_25562,N_23481,N_22399);
nand U25563 (N_25563,N_22481,N_22563);
xnor U25564 (N_25564,N_22059,N_23065);
and U25565 (N_25565,N_22538,N_21588);
xor U25566 (N_25566,N_21635,N_21499);
and U25567 (N_25567,N_21531,N_22010);
xnor U25568 (N_25568,N_22810,N_22640);
xnor U25569 (N_25569,N_21214,N_21645);
nand U25570 (N_25570,N_22550,N_23496);
xnor U25571 (N_25571,N_22658,N_23183);
nor U25572 (N_25572,N_21158,N_23629);
and U25573 (N_25573,N_22234,N_21585);
and U25574 (N_25574,N_22552,N_21846);
and U25575 (N_25575,N_21305,N_22293);
nor U25576 (N_25576,N_23877,N_23641);
xnor U25577 (N_25577,N_23730,N_21818);
and U25578 (N_25578,N_21848,N_22943);
xor U25579 (N_25579,N_23440,N_23347);
and U25580 (N_25580,N_23866,N_21059);
xor U25581 (N_25581,N_21910,N_23869);
and U25582 (N_25582,N_21928,N_22913);
xor U25583 (N_25583,N_21832,N_22550);
or U25584 (N_25584,N_21575,N_22760);
xor U25585 (N_25585,N_22744,N_22015);
nor U25586 (N_25586,N_22866,N_22933);
xnor U25587 (N_25587,N_23376,N_22253);
nor U25588 (N_25588,N_22037,N_21898);
nand U25589 (N_25589,N_23741,N_23392);
and U25590 (N_25590,N_23369,N_21747);
and U25591 (N_25591,N_23597,N_22764);
nor U25592 (N_25592,N_21442,N_23665);
and U25593 (N_25593,N_22825,N_23605);
nand U25594 (N_25594,N_22227,N_22316);
and U25595 (N_25595,N_21551,N_22370);
nor U25596 (N_25596,N_23624,N_22687);
xnor U25597 (N_25597,N_21517,N_23781);
nand U25598 (N_25598,N_23983,N_22610);
or U25599 (N_25599,N_22807,N_21530);
xnor U25600 (N_25600,N_23503,N_23380);
or U25601 (N_25601,N_22944,N_23153);
nand U25602 (N_25602,N_22026,N_23896);
nor U25603 (N_25603,N_22286,N_21252);
nor U25604 (N_25604,N_21975,N_21741);
nor U25605 (N_25605,N_21748,N_23818);
or U25606 (N_25606,N_21951,N_22292);
nand U25607 (N_25607,N_22677,N_21633);
nand U25608 (N_25608,N_21370,N_21214);
or U25609 (N_25609,N_23731,N_22328);
xnor U25610 (N_25610,N_22304,N_22701);
and U25611 (N_25611,N_22716,N_23322);
or U25612 (N_25612,N_21342,N_23312);
or U25613 (N_25613,N_21879,N_21607);
nand U25614 (N_25614,N_21297,N_22514);
nand U25615 (N_25615,N_22310,N_21864);
nand U25616 (N_25616,N_21913,N_22158);
or U25617 (N_25617,N_21344,N_22353);
nor U25618 (N_25618,N_23034,N_22575);
and U25619 (N_25619,N_23502,N_23842);
nor U25620 (N_25620,N_22293,N_23124);
or U25621 (N_25621,N_22784,N_21079);
xor U25622 (N_25622,N_22137,N_23446);
xnor U25623 (N_25623,N_22007,N_22836);
nand U25624 (N_25624,N_23224,N_23059);
xor U25625 (N_25625,N_22892,N_23427);
nor U25626 (N_25626,N_22911,N_23770);
xor U25627 (N_25627,N_21423,N_21170);
and U25628 (N_25628,N_23020,N_23952);
xnor U25629 (N_25629,N_22694,N_23443);
nor U25630 (N_25630,N_21575,N_21229);
nand U25631 (N_25631,N_21357,N_23362);
and U25632 (N_25632,N_21557,N_23866);
and U25633 (N_25633,N_22194,N_23676);
and U25634 (N_25634,N_21911,N_22727);
xor U25635 (N_25635,N_22794,N_21688);
and U25636 (N_25636,N_23288,N_22766);
nand U25637 (N_25637,N_23268,N_21700);
nor U25638 (N_25638,N_22779,N_23789);
xnor U25639 (N_25639,N_22789,N_23232);
and U25640 (N_25640,N_21264,N_22251);
xnor U25641 (N_25641,N_23501,N_21371);
nand U25642 (N_25642,N_22407,N_23975);
nor U25643 (N_25643,N_21615,N_21313);
nand U25644 (N_25644,N_21863,N_23351);
nor U25645 (N_25645,N_21145,N_23398);
nor U25646 (N_25646,N_22791,N_23295);
xor U25647 (N_25647,N_22049,N_22752);
nor U25648 (N_25648,N_21576,N_22579);
nor U25649 (N_25649,N_22650,N_21106);
or U25650 (N_25650,N_22884,N_23124);
and U25651 (N_25651,N_22486,N_21139);
nor U25652 (N_25652,N_22623,N_23268);
nand U25653 (N_25653,N_23102,N_23161);
or U25654 (N_25654,N_21726,N_21432);
or U25655 (N_25655,N_21700,N_21827);
nand U25656 (N_25656,N_23522,N_22220);
and U25657 (N_25657,N_21229,N_22439);
nand U25658 (N_25658,N_21659,N_21457);
or U25659 (N_25659,N_21493,N_23876);
xor U25660 (N_25660,N_23222,N_22973);
or U25661 (N_25661,N_23561,N_22592);
nand U25662 (N_25662,N_21729,N_22272);
and U25663 (N_25663,N_23612,N_21140);
xnor U25664 (N_25664,N_23854,N_22634);
nand U25665 (N_25665,N_21965,N_21129);
nand U25666 (N_25666,N_23721,N_22059);
nor U25667 (N_25667,N_22088,N_23834);
nand U25668 (N_25668,N_23146,N_23688);
nand U25669 (N_25669,N_22925,N_23463);
or U25670 (N_25670,N_22616,N_22153);
or U25671 (N_25671,N_23260,N_23288);
or U25672 (N_25672,N_23950,N_22738);
or U25673 (N_25673,N_22936,N_23092);
or U25674 (N_25674,N_22041,N_21353);
and U25675 (N_25675,N_23157,N_22451);
and U25676 (N_25676,N_21943,N_22171);
nor U25677 (N_25677,N_23662,N_21394);
nor U25678 (N_25678,N_21130,N_22315);
nor U25679 (N_25679,N_23773,N_23980);
nand U25680 (N_25680,N_23630,N_21892);
xnor U25681 (N_25681,N_22543,N_23094);
xor U25682 (N_25682,N_22438,N_22380);
nor U25683 (N_25683,N_22229,N_22142);
xor U25684 (N_25684,N_22604,N_22652);
nor U25685 (N_25685,N_21908,N_22176);
nor U25686 (N_25686,N_21613,N_21160);
xnor U25687 (N_25687,N_21525,N_23797);
nor U25688 (N_25688,N_21361,N_23673);
nor U25689 (N_25689,N_22215,N_22056);
or U25690 (N_25690,N_21647,N_23299);
nor U25691 (N_25691,N_21208,N_23178);
or U25692 (N_25692,N_22730,N_23014);
and U25693 (N_25693,N_21277,N_23715);
or U25694 (N_25694,N_23609,N_23184);
nand U25695 (N_25695,N_21142,N_23717);
xnor U25696 (N_25696,N_23713,N_21425);
or U25697 (N_25697,N_21056,N_22416);
or U25698 (N_25698,N_23437,N_23364);
or U25699 (N_25699,N_21415,N_21534);
nor U25700 (N_25700,N_21549,N_23303);
and U25701 (N_25701,N_21323,N_23205);
or U25702 (N_25702,N_23135,N_22339);
or U25703 (N_25703,N_22919,N_23684);
and U25704 (N_25704,N_23343,N_22695);
nor U25705 (N_25705,N_23125,N_21687);
or U25706 (N_25706,N_23859,N_23471);
nor U25707 (N_25707,N_22271,N_22253);
xor U25708 (N_25708,N_21274,N_23416);
and U25709 (N_25709,N_22779,N_21535);
nand U25710 (N_25710,N_22927,N_22019);
nor U25711 (N_25711,N_23243,N_23006);
nand U25712 (N_25712,N_23376,N_23626);
xor U25713 (N_25713,N_23724,N_21046);
nand U25714 (N_25714,N_23672,N_22049);
or U25715 (N_25715,N_21663,N_22642);
nand U25716 (N_25716,N_23981,N_22469);
and U25717 (N_25717,N_21737,N_23227);
nor U25718 (N_25718,N_21387,N_22710);
nand U25719 (N_25719,N_22004,N_23700);
and U25720 (N_25720,N_21470,N_23118);
or U25721 (N_25721,N_23706,N_21610);
nor U25722 (N_25722,N_23480,N_21500);
or U25723 (N_25723,N_22451,N_23763);
or U25724 (N_25724,N_22296,N_21079);
nand U25725 (N_25725,N_23153,N_21932);
and U25726 (N_25726,N_22168,N_22568);
and U25727 (N_25727,N_22713,N_22691);
and U25728 (N_25728,N_21732,N_22184);
and U25729 (N_25729,N_22756,N_21175);
and U25730 (N_25730,N_22360,N_23100);
xnor U25731 (N_25731,N_22345,N_21042);
nand U25732 (N_25732,N_23935,N_23363);
xnor U25733 (N_25733,N_22792,N_22361);
xnor U25734 (N_25734,N_22435,N_21872);
and U25735 (N_25735,N_21939,N_22202);
or U25736 (N_25736,N_23837,N_23325);
or U25737 (N_25737,N_21002,N_21338);
or U25738 (N_25738,N_22836,N_22910);
nor U25739 (N_25739,N_23710,N_22713);
or U25740 (N_25740,N_23165,N_22430);
and U25741 (N_25741,N_21632,N_22468);
nand U25742 (N_25742,N_22216,N_23382);
and U25743 (N_25743,N_23965,N_23798);
nand U25744 (N_25744,N_23148,N_21581);
or U25745 (N_25745,N_21554,N_22271);
xor U25746 (N_25746,N_22618,N_22614);
nand U25747 (N_25747,N_22486,N_22920);
or U25748 (N_25748,N_23040,N_23388);
nor U25749 (N_25749,N_22789,N_21137);
or U25750 (N_25750,N_22618,N_23098);
and U25751 (N_25751,N_22472,N_22939);
xnor U25752 (N_25752,N_23670,N_23669);
nor U25753 (N_25753,N_22880,N_22727);
and U25754 (N_25754,N_22103,N_23399);
xor U25755 (N_25755,N_22097,N_21537);
or U25756 (N_25756,N_21830,N_21920);
nor U25757 (N_25757,N_22099,N_23385);
nand U25758 (N_25758,N_23008,N_21442);
nor U25759 (N_25759,N_23113,N_22485);
or U25760 (N_25760,N_21882,N_22768);
nand U25761 (N_25761,N_22064,N_23173);
and U25762 (N_25762,N_23256,N_22646);
xor U25763 (N_25763,N_21111,N_22416);
or U25764 (N_25764,N_22667,N_21736);
xnor U25765 (N_25765,N_22848,N_22371);
or U25766 (N_25766,N_22275,N_23702);
or U25767 (N_25767,N_23606,N_23420);
or U25768 (N_25768,N_21150,N_21601);
and U25769 (N_25769,N_21943,N_21754);
xor U25770 (N_25770,N_23994,N_22267);
and U25771 (N_25771,N_21713,N_23381);
nand U25772 (N_25772,N_22306,N_21372);
nand U25773 (N_25773,N_23335,N_23456);
or U25774 (N_25774,N_23279,N_21164);
and U25775 (N_25775,N_22063,N_23948);
nand U25776 (N_25776,N_23857,N_22530);
nor U25777 (N_25777,N_21266,N_23860);
or U25778 (N_25778,N_23632,N_23423);
nand U25779 (N_25779,N_23526,N_21000);
nand U25780 (N_25780,N_23182,N_22603);
or U25781 (N_25781,N_23015,N_23606);
nor U25782 (N_25782,N_22395,N_22519);
xor U25783 (N_25783,N_22864,N_21538);
nor U25784 (N_25784,N_22347,N_21346);
nand U25785 (N_25785,N_23230,N_22556);
and U25786 (N_25786,N_22676,N_21347);
or U25787 (N_25787,N_23448,N_21029);
nor U25788 (N_25788,N_22453,N_21648);
nor U25789 (N_25789,N_21159,N_23585);
nor U25790 (N_25790,N_21258,N_21995);
and U25791 (N_25791,N_21745,N_21877);
and U25792 (N_25792,N_22279,N_23724);
nand U25793 (N_25793,N_21980,N_22079);
nor U25794 (N_25794,N_21770,N_21586);
or U25795 (N_25795,N_21549,N_23811);
nor U25796 (N_25796,N_21452,N_23812);
nor U25797 (N_25797,N_23396,N_22852);
and U25798 (N_25798,N_21479,N_23478);
nor U25799 (N_25799,N_21407,N_22560);
nor U25800 (N_25800,N_21956,N_21027);
and U25801 (N_25801,N_21711,N_23755);
and U25802 (N_25802,N_23326,N_21196);
xnor U25803 (N_25803,N_23456,N_21665);
xor U25804 (N_25804,N_22591,N_21186);
and U25805 (N_25805,N_22549,N_22219);
xnor U25806 (N_25806,N_22431,N_22607);
xnor U25807 (N_25807,N_22863,N_23705);
or U25808 (N_25808,N_22272,N_21453);
or U25809 (N_25809,N_21933,N_23295);
nand U25810 (N_25810,N_23950,N_23017);
nor U25811 (N_25811,N_23330,N_22057);
nor U25812 (N_25812,N_23083,N_22923);
nand U25813 (N_25813,N_21222,N_23414);
xor U25814 (N_25814,N_21871,N_21124);
and U25815 (N_25815,N_22090,N_23157);
xor U25816 (N_25816,N_23285,N_22874);
xnor U25817 (N_25817,N_22264,N_21860);
xnor U25818 (N_25818,N_21577,N_22522);
nor U25819 (N_25819,N_23014,N_23059);
nor U25820 (N_25820,N_22219,N_21813);
and U25821 (N_25821,N_23233,N_22274);
or U25822 (N_25822,N_23847,N_21104);
or U25823 (N_25823,N_22164,N_22352);
nor U25824 (N_25824,N_22895,N_22774);
nand U25825 (N_25825,N_22720,N_23945);
and U25826 (N_25826,N_21314,N_22978);
nand U25827 (N_25827,N_22219,N_21249);
nor U25828 (N_25828,N_23741,N_23142);
nand U25829 (N_25829,N_23282,N_22344);
xor U25830 (N_25830,N_22311,N_22574);
or U25831 (N_25831,N_23950,N_22420);
xor U25832 (N_25832,N_21089,N_21970);
and U25833 (N_25833,N_23792,N_22693);
or U25834 (N_25834,N_22879,N_22694);
and U25835 (N_25835,N_21563,N_21031);
nand U25836 (N_25836,N_22488,N_22839);
and U25837 (N_25837,N_22533,N_21289);
nand U25838 (N_25838,N_23629,N_23130);
nor U25839 (N_25839,N_22269,N_23055);
or U25840 (N_25840,N_21921,N_22509);
and U25841 (N_25841,N_21070,N_23761);
and U25842 (N_25842,N_23873,N_22727);
nor U25843 (N_25843,N_21740,N_23786);
nand U25844 (N_25844,N_23795,N_22596);
nand U25845 (N_25845,N_21690,N_23260);
xor U25846 (N_25846,N_21237,N_21980);
xnor U25847 (N_25847,N_21830,N_21241);
nor U25848 (N_25848,N_22449,N_23742);
nand U25849 (N_25849,N_23492,N_21214);
nor U25850 (N_25850,N_22269,N_21021);
and U25851 (N_25851,N_22090,N_21154);
nor U25852 (N_25852,N_21223,N_23509);
nor U25853 (N_25853,N_21483,N_21522);
nand U25854 (N_25854,N_22033,N_21870);
nor U25855 (N_25855,N_23585,N_21403);
or U25856 (N_25856,N_22599,N_22365);
xnor U25857 (N_25857,N_22037,N_21412);
and U25858 (N_25858,N_23953,N_21372);
and U25859 (N_25859,N_23481,N_23719);
nand U25860 (N_25860,N_22664,N_22942);
nor U25861 (N_25861,N_23243,N_23701);
xnor U25862 (N_25862,N_22904,N_23574);
xor U25863 (N_25863,N_22792,N_21618);
and U25864 (N_25864,N_21859,N_23033);
and U25865 (N_25865,N_22719,N_22063);
xor U25866 (N_25866,N_23435,N_23503);
and U25867 (N_25867,N_21745,N_21014);
and U25868 (N_25868,N_23320,N_22236);
and U25869 (N_25869,N_21795,N_22495);
or U25870 (N_25870,N_22761,N_23739);
nand U25871 (N_25871,N_23133,N_23534);
and U25872 (N_25872,N_21987,N_22318);
xor U25873 (N_25873,N_23741,N_22271);
xnor U25874 (N_25874,N_21785,N_23330);
or U25875 (N_25875,N_23106,N_22147);
or U25876 (N_25876,N_22833,N_22753);
nand U25877 (N_25877,N_21247,N_21743);
nand U25878 (N_25878,N_22008,N_21531);
and U25879 (N_25879,N_23631,N_22256);
xnor U25880 (N_25880,N_23174,N_23581);
nand U25881 (N_25881,N_21385,N_23675);
nand U25882 (N_25882,N_23069,N_22817);
and U25883 (N_25883,N_21255,N_23510);
and U25884 (N_25884,N_23806,N_23468);
nor U25885 (N_25885,N_23824,N_22695);
and U25886 (N_25886,N_22375,N_23487);
or U25887 (N_25887,N_23031,N_22132);
xor U25888 (N_25888,N_21218,N_22888);
nor U25889 (N_25889,N_23696,N_22344);
and U25890 (N_25890,N_23462,N_21303);
nor U25891 (N_25891,N_23939,N_22535);
or U25892 (N_25892,N_22336,N_21279);
or U25893 (N_25893,N_22993,N_22251);
nand U25894 (N_25894,N_22574,N_22353);
and U25895 (N_25895,N_23383,N_23114);
and U25896 (N_25896,N_21022,N_23170);
xnor U25897 (N_25897,N_22043,N_23394);
and U25898 (N_25898,N_21981,N_21994);
and U25899 (N_25899,N_21278,N_22062);
nand U25900 (N_25900,N_21633,N_23120);
and U25901 (N_25901,N_21752,N_21075);
nand U25902 (N_25902,N_21215,N_23217);
nor U25903 (N_25903,N_22686,N_22545);
xor U25904 (N_25904,N_21637,N_22392);
nor U25905 (N_25905,N_21773,N_21713);
or U25906 (N_25906,N_22245,N_21920);
nand U25907 (N_25907,N_23435,N_22216);
and U25908 (N_25908,N_23324,N_21807);
or U25909 (N_25909,N_22109,N_22762);
or U25910 (N_25910,N_22714,N_22898);
or U25911 (N_25911,N_23719,N_23070);
and U25912 (N_25912,N_23667,N_22003);
or U25913 (N_25913,N_21895,N_22930);
and U25914 (N_25914,N_23019,N_23406);
or U25915 (N_25915,N_22778,N_23024);
nand U25916 (N_25916,N_23822,N_23158);
or U25917 (N_25917,N_22220,N_22777);
or U25918 (N_25918,N_23193,N_22419);
nor U25919 (N_25919,N_22100,N_21437);
and U25920 (N_25920,N_21297,N_22471);
nand U25921 (N_25921,N_22249,N_21923);
nand U25922 (N_25922,N_21475,N_21403);
xnor U25923 (N_25923,N_21461,N_21818);
xnor U25924 (N_25924,N_23471,N_22936);
xor U25925 (N_25925,N_22921,N_23713);
or U25926 (N_25926,N_21624,N_22316);
or U25927 (N_25927,N_23647,N_21314);
nand U25928 (N_25928,N_22491,N_22906);
xnor U25929 (N_25929,N_23610,N_21479);
or U25930 (N_25930,N_22543,N_21240);
or U25931 (N_25931,N_23203,N_21566);
and U25932 (N_25932,N_23766,N_23210);
and U25933 (N_25933,N_23254,N_21573);
and U25934 (N_25934,N_21990,N_21632);
nand U25935 (N_25935,N_22909,N_23930);
and U25936 (N_25936,N_22009,N_23135);
and U25937 (N_25937,N_21563,N_23021);
nor U25938 (N_25938,N_22817,N_22685);
or U25939 (N_25939,N_21362,N_23914);
or U25940 (N_25940,N_22801,N_23899);
xor U25941 (N_25941,N_21858,N_21923);
or U25942 (N_25942,N_22406,N_23580);
and U25943 (N_25943,N_23890,N_23653);
and U25944 (N_25944,N_23077,N_23263);
xor U25945 (N_25945,N_23168,N_21117);
nand U25946 (N_25946,N_23428,N_23420);
and U25947 (N_25947,N_23290,N_23545);
xnor U25948 (N_25948,N_22520,N_23883);
xnor U25949 (N_25949,N_21077,N_21155);
nor U25950 (N_25950,N_21304,N_21977);
or U25951 (N_25951,N_22305,N_23754);
nand U25952 (N_25952,N_21821,N_23699);
xnor U25953 (N_25953,N_22318,N_23065);
or U25954 (N_25954,N_22212,N_23135);
nand U25955 (N_25955,N_21016,N_21155);
nand U25956 (N_25956,N_22217,N_22934);
nor U25957 (N_25957,N_21098,N_23764);
and U25958 (N_25958,N_21593,N_22585);
and U25959 (N_25959,N_22308,N_22899);
or U25960 (N_25960,N_22003,N_21126);
and U25961 (N_25961,N_23917,N_22254);
xor U25962 (N_25962,N_23543,N_22176);
and U25963 (N_25963,N_23117,N_21423);
or U25964 (N_25964,N_23990,N_23774);
xor U25965 (N_25965,N_22860,N_21103);
or U25966 (N_25966,N_21169,N_21077);
and U25967 (N_25967,N_23525,N_23800);
nor U25968 (N_25968,N_21001,N_23358);
nor U25969 (N_25969,N_22051,N_22407);
nor U25970 (N_25970,N_21415,N_23206);
xor U25971 (N_25971,N_23939,N_23008);
and U25972 (N_25972,N_21412,N_22544);
nand U25973 (N_25973,N_23734,N_21049);
and U25974 (N_25974,N_23122,N_21725);
nor U25975 (N_25975,N_23597,N_22781);
or U25976 (N_25976,N_22461,N_22454);
or U25977 (N_25977,N_22928,N_21947);
or U25978 (N_25978,N_22649,N_23492);
nor U25979 (N_25979,N_23734,N_21390);
xor U25980 (N_25980,N_21927,N_21874);
and U25981 (N_25981,N_22798,N_23810);
nor U25982 (N_25982,N_22526,N_21616);
nor U25983 (N_25983,N_23958,N_23254);
xor U25984 (N_25984,N_23009,N_23093);
or U25985 (N_25985,N_23405,N_23051);
and U25986 (N_25986,N_21125,N_23055);
xor U25987 (N_25987,N_22589,N_23923);
and U25988 (N_25988,N_22147,N_22455);
and U25989 (N_25989,N_23396,N_22728);
or U25990 (N_25990,N_22707,N_22653);
nor U25991 (N_25991,N_23890,N_21511);
and U25992 (N_25992,N_21998,N_21207);
or U25993 (N_25993,N_23455,N_22963);
and U25994 (N_25994,N_22678,N_23315);
or U25995 (N_25995,N_21155,N_22662);
xnor U25996 (N_25996,N_23932,N_22670);
or U25997 (N_25997,N_22953,N_21983);
nor U25998 (N_25998,N_21742,N_23618);
and U25999 (N_25999,N_23341,N_21974);
xor U26000 (N_26000,N_21973,N_22323);
nor U26001 (N_26001,N_22419,N_22016);
xnor U26002 (N_26002,N_21665,N_21387);
or U26003 (N_26003,N_23585,N_22017);
or U26004 (N_26004,N_22889,N_22724);
and U26005 (N_26005,N_22413,N_21294);
nand U26006 (N_26006,N_22716,N_21697);
and U26007 (N_26007,N_22748,N_21827);
or U26008 (N_26008,N_23322,N_22221);
or U26009 (N_26009,N_21965,N_22797);
or U26010 (N_26010,N_22520,N_23376);
and U26011 (N_26011,N_23157,N_23307);
or U26012 (N_26012,N_21132,N_23302);
nor U26013 (N_26013,N_21710,N_21778);
xor U26014 (N_26014,N_23716,N_22420);
nand U26015 (N_26015,N_21157,N_21360);
xor U26016 (N_26016,N_23367,N_21489);
nand U26017 (N_26017,N_22577,N_22926);
and U26018 (N_26018,N_23982,N_22779);
nor U26019 (N_26019,N_23472,N_23775);
nand U26020 (N_26020,N_23259,N_21144);
or U26021 (N_26021,N_21246,N_23691);
nand U26022 (N_26022,N_22338,N_21614);
xnor U26023 (N_26023,N_22606,N_23682);
nor U26024 (N_26024,N_22521,N_22558);
or U26025 (N_26025,N_22480,N_23368);
or U26026 (N_26026,N_22348,N_21981);
or U26027 (N_26027,N_21987,N_22040);
and U26028 (N_26028,N_22563,N_22646);
or U26029 (N_26029,N_23843,N_21795);
or U26030 (N_26030,N_21370,N_23103);
xnor U26031 (N_26031,N_23616,N_21903);
nor U26032 (N_26032,N_22628,N_23107);
and U26033 (N_26033,N_23513,N_23774);
and U26034 (N_26034,N_21365,N_22304);
nor U26035 (N_26035,N_22035,N_21173);
and U26036 (N_26036,N_23944,N_21813);
or U26037 (N_26037,N_22662,N_22818);
or U26038 (N_26038,N_23130,N_21924);
or U26039 (N_26039,N_22039,N_22369);
or U26040 (N_26040,N_21098,N_21850);
and U26041 (N_26041,N_23722,N_21233);
nand U26042 (N_26042,N_23811,N_23977);
and U26043 (N_26043,N_21792,N_22828);
or U26044 (N_26044,N_21513,N_21422);
nor U26045 (N_26045,N_23074,N_23737);
xnor U26046 (N_26046,N_23532,N_22797);
nand U26047 (N_26047,N_21533,N_22999);
or U26048 (N_26048,N_21701,N_23510);
and U26049 (N_26049,N_21429,N_23467);
xnor U26050 (N_26050,N_21291,N_21516);
xnor U26051 (N_26051,N_21361,N_22645);
nor U26052 (N_26052,N_22436,N_22165);
and U26053 (N_26053,N_23173,N_23528);
nor U26054 (N_26054,N_21208,N_22460);
nor U26055 (N_26055,N_23069,N_22606);
nand U26056 (N_26056,N_23152,N_23158);
or U26057 (N_26057,N_22533,N_23227);
xnor U26058 (N_26058,N_23684,N_21325);
xor U26059 (N_26059,N_23830,N_22181);
and U26060 (N_26060,N_23733,N_21282);
xor U26061 (N_26061,N_23881,N_23192);
nand U26062 (N_26062,N_21820,N_23041);
or U26063 (N_26063,N_21971,N_21387);
xnor U26064 (N_26064,N_21805,N_22094);
and U26065 (N_26065,N_23488,N_22232);
or U26066 (N_26066,N_23331,N_23940);
nor U26067 (N_26067,N_23531,N_23328);
nor U26068 (N_26068,N_23658,N_22004);
nand U26069 (N_26069,N_23400,N_22465);
xnor U26070 (N_26070,N_23673,N_23474);
and U26071 (N_26071,N_21671,N_21301);
or U26072 (N_26072,N_22021,N_21405);
nor U26073 (N_26073,N_21035,N_22868);
nand U26074 (N_26074,N_23577,N_23716);
nor U26075 (N_26075,N_22370,N_23234);
or U26076 (N_26076,N_22179,N_21344);
or U26077 (N_26077,N_21612,N_23467);
nor U26078 (N_26078,N_23637,N_21703);
nand U26079 (N_26079,N_21864,N_21931);
or U26080 (N_26080,N_21174,N_21653);
nand U26081 (N_26081,N_23757,N_23035);
or U26082 (N_26082,N_22190,N_23787);
nand U26083 (N_26083,N_23550,N_22619);
or U26084 (N_26084,N_22518,N_22397);
nand U26085 (N_26085,N_22968,N_22458);
and U26086 (N_26086,N_22918,N_23946);
xor U26087 (N_26087,N_21493,N_22611);
xor U26088 (N_26088,N_23236,N_21223);
nand U26089 (N_26089,N_22532,N_23070);
nor U26090 (N_26090,N_21649,N_21712);
nor U26091 (N_26091,N_23581,N_21076);
and U26092 (N_26092,N_23043,N_21407);
xnor U26093 (N_26093,N_22906,N_23357);
and U26094 (N_26094,N_21499,N_23206);
and U26095 (N_26095,N_21535,N_22003);
and U26096 (N_26096,N_22481,N_21743);
nor U26097 (N_26097,N_21077,N_23200);
and U26098 (N_26098,N_22810,N_23308);
nand U26099 (N_26099,N_22106,N_23359);
xnor U26100 (N_26100,N_23849,N_22964);
xnor U26101 (N_26101,N_21769,N_23893);
and U26102 (N_26102,N_23218,N_22077);
nor U26103 (N_26103,N_23209,N_23191);
xor U26104 (N_26104,N_22319,N_23961);
nor U26105 (N_26105,N_23350,N_21805);
and U26106 (N_26106,N_22739,N_23786);
nor U26107 (N_26107,N_22497,N_21863);
and U26108 (N_26108,N_21533,N_22264);
xor U26109 (N_26109,N_21120,N_23355);
or U26110 (N_26110,N_22120,N_21448);
xor U26111 (N_26111,N_22749,N_22303);
nand U26112 (N_26112,N_23406,N_22096);
and U26113 (N_26113,N_23984,N_23214);
and U26114 (N_26114,N_22146,N_22672);
and U26115 (N_26115,N_22007,N_22151);
nand U26116 (N_26116,N_22023,N_21536);
xor U26117 (N_26117,N_22728,N_22559);
and U26118 (N_26118,N_22144,N_21908);
and U26119 (N_26119,N_23857,N_22864);
nand U26120 (N_26120,N_21097,N_23217);
nand U26121 (N_26121,N_23333,N_23442);
nor U26122 (N_26122,N_21844,N_23716);
nor U26123 (N_26123,N_21490,N_23057);
and U26124 (N_26124,N_22244,N_23266);
and U26125 (N_26125,N_23479,N_23303);
xnor U26126 (N_26126,N_22407,N_22417);
xor U26127 (N_26127,N_23618,N_22514);
or U26128 (N_26128,N_23725,N_22425);
nand U26129 (N_26129,N_22300,N_22373);
and U26130 (N_26130,N_21670,N_22118);
nand U26131 (N_26131,N_21605,N_21349);
nor U26132 (N_26132,N_21788,N_21958);
and U26133 (N_26133,N_21508,N_21828);
nor U26134 (N_26134,N_23361,N_22853);
xnor U26135 (N_26135,N_23704,N_22572);
xor U26136 (N_26136,N_22626,N_23402);
or U26137 (N_26137,N_21989,N_21629);
nor U26138 (N_26138,N_22275,N_23886);
and U26139 (N_26139,N_23505,N_22323);
or U26140 (N_26140,N_22314,N_22857);
xnor U26141 (N_26141,N_22237,N_22563);
nor U26142 (N_26142,N_22856,N_23282);
nand U26143 (N_26143,N_22947,N_23797);
or U26144 (N_26144,N_22878,N_21545);
and U26145 (N_26145,N_21580,N_21516);
nand U26146 (N_26146,N_23061,N_22864);
and U26147 (N_26147,N_23993,N_22756);
nor U26148 (N_26148,N_23123,N_21033);
xor U26149 (N_26149,N_22765,N_23859);
xor U26150 (N_26150,N_22150,N_23255);
nand U26151 (N_26151,N_23454,N_21987);
or U26152 (N_26152,N_21948,N_22010);
nand U26153 (N_26153,N_22224,N_23740);
or U26154 (N_26154,N_22565,N_21471);
nand U26155 (N_26155,N_23239,N_22179);
nand U26156 (N_26156,N_21912,N_23280);
xor U26157 (N_26157,N_23224,N_21430);
xor U26158 (N_26158,N_23619,N_22457);
and U26159 (N_26159,N_22355,N_21422);
nor U26160 (N_26160,N_23533,N_23532);
and U26161 (N_26161,N_22108,N_22681);
nand U26162 (N_26162,N_21787,N_22848);
nor U26163 (N_26163,N_22751,N_22384);
nand U26164 (N_26164,N_21736,N_21858);
nor U26165 (N_26165,N_23758,N_23083);
and U26166 (N_26166,N_21066,N_22052);
nor U26167 (N_26167,N_22893,N_22660);
nor U26168 (N_26168,N_21795,N_23666);
or U26169 (N_26169,N_23182,N_21367);
or U26170 (N_26170,N_23755,N_23766);
or U26171 (N_26171,N_22410,N_22093);
or U26172 (N_26172,N_22823,N_23148);
nor U26173 (N_26173,N_21517,N_22552);
nand U26174 (N_26174,N_22034,N_23471);
nor U26175 (N_26175,N_23354,N_23843);
nor U26176 (N_26176,N_21526,N_23734);
and U26177 (N_26177,N_21680,N_22328);
or U26178 (N_26178,N_22613,N_21908);
or U26179 (N_26179,N_23204,N_22387);
nand U26180 (N_26180,N_21586,N_23088);
and U26181 (N_26181,N_21423,N_21110);
nor U26182 (N_26182,N_23569,N_22508);
nor U26183 (N_26183,N_23292,N_22066);
xnor U26184 (N_26184,N_22087,N_23341);
nand U26185 (N_26185,N_22619,N_22440);
or U26186 (N_26186,N_21923,N_22818);
nand U26187 (N_26187,N_23555,N_22253);
xnor U26188 (N_26188,N_21932,N_21817);
xor U26189 (N_26189,N_22449,N_22876);
and U26190 (N_26190,N_23383,N_23242);
and U26191 (N_26191,N_21101,N_22191);
or U26192 (N_26192,N_23967,N_21604);
nor U26193 (N_26193,N_22942,N_23900);
xnor U26194 (N_26194,N_22168,N_21094);
or U26195 (N_26195,N_21339,N_22615);
xor U26196 (N_26196,N_23427,N_21779);
and U26197 (N_26197,N_22362,N_21277);
xor U26198 (N_26198,N_21282,N_22857);
or U26199 (N_26199,N_23385,N_22457);
or U26200 (N_26200,N_21950,N_23215);
xnor U26201 (N_26201,N_22516,N_23626);
xor U26202 (N_26202,N_21094,N_22053);
and U26203 (N_26203,N_23540,N_23713);
and U26204 (N_26204,N_23587,N_23512);
nand U26205 (N_26205,N_22833,N_22741);
nand U26206 (N_26206,N_22074,N_22865);
xnor U26207 (N_26207,N_23635,N_22973);
nand U26208 (N_26208,N_23231,N_22055);
nand U26209 (N_26209,N_23360,N_23030);
and U26210 (N_26210,N_21741,N_22366);
nand U26211 (N_26211,N_22779,N_22086);
or U26212 (N_26212,N_22780,N_23413);
and U26213 (N_26213,N_21452,N_21920);
nor U26214 (N_26214,N_23966,N_22301);
nand U26215 (N_26215,N_23139,N_22724);
nor U26216 (N_26216,N_21594,N_23975);
or U26217 (N_26217,N_21727,N_22663);
and U26218 (N_26218,N_23306,N_22838);
or U26219 (N_26219,N_22663,N_23404);
nor U26220 (N_26220,N_23763,N_23308);
xnor U26221 (N_26221,N_23843,N_23155);
nand U26222 (N_26222,N_23261,N_21746);
or U26223 (N_26223,N_23684,N_23814);
and U26224 (N_26224,N_23802,N_23943);
or U26225 (N_26225,N_21012,N_23170);
nor U26226 (N_26226,N_22225,N_23589);
or U26227 (N_26227,N_21091,N_23496);
nand U26228 (N_26228,N_22416,N_21087);
nor U26229 (N_26229,N_21945,N_22465);
or U26230 (N_26230,N_21800,N_21608);
and U26231 (N_26231,N_22170,N_21950);
xor U26232 (N_26232,N_23402,N_21983);
and U26233 (N_26233,N_23134,N_22018);
xnor U26234 (N_26234,N_23935,N_21310);
or U26235 (N_26235,N_22318,N_22673);
xor U26236 (N_26236,N_22816,N_23331);
or U26237 (N_26237,N_22608,N_21713);
and U26238 (N_26238,N_21303,N_21596);
and U26239 (N_26239,N_21585,N_22096);
and U26240 (N_26240,N_23400,N_23536);
nand U26241 (N_26241,N_23578,N_21765);
or U26242 (N_26242,N_21217,N_21644);
xor U26243 (N_26243,N_21231,N_21213);
nand U26244 (N_26244,N_21210,N_21486);
nand U26245 (N_26245,N_21932,N_22601);
nand U26246 (N_26246,N_21331,N_23091);
nor U26247 (N_26247,N_21278,N_21763);
or U26248 (N_26248,N_21860,N_21131);
xor U26249 (N_26249,N_23747,N_22618);
nor U26250 (N_26250,N_21582,N_22261);
or U26251 (N_26251,N_21706,N_21278);
and U26252 (N_26252,N_23414,N_21724);
xnor U26253 (N_26253,N_23553,N_23215);
nand U26254 (N_26254,N_21296,N_23686);
and U26255 (N_26255,N_23540,N_22332);
and U26256 (N_26256,N_22535,N_21276);
nand U26257 (N_26257,N_23217,N_23921);
xor U26258 (N_26258,N_23883,N_23232);
and U26259 (N_26259,N_23019,N_23591);
nor U26260 (N_26260,N_21717,N_21546);
xnor U26261 (N_26261,N_22314,N_23011);
nand U26262 (N_26262,N_22265,N_22936);
or U26263 (N_26263,N_21581,N_22499);
and U26264 (N_26264,N_22043,N_23993);
or U26265 (N_26265,N_22188,N_22486);
and U26266 (N_26266,N_23141,N_21472);
nor U26267 (N_26267,N_22933,N_23752);
or U26268 (N_26268,N_23760,N_22258);
and U26269 (N_26269,N_23929,N_22738);
and U26270 (N_26270,N_21853,N_22964);
and U26271 (N_26271,N_23645,N_23748);
nand U26272 (N_26272,N_21984,N_23348);
xnor U26273 (N_26273,N_22133,N_22364);
nand U26274 (N_26274,N_23718,N_23268);
nand U26275 (N_26275,N_21066,N_22130);
nor U26276 (N_26276,N_23577,N_21205);
xnor U26277 (N_26277,N_21450,N_23279);
nand U26278 (N_26278,N_23722,N_23294);
nor U26279 (N_26279,N_23860,N_22027);
nor U26280 (N_26280,N_23989,N_23647);
nor U26281 (N_26281,N_23302,N_22236);
xnor U26282 (N_26282,N_21359,N_23627);
nor U26283 (N_26283,N_23634,N_22451);
xor U26284 (N_26284,N_21994,N_22374);
nand U26285 (N_26285,N_22421,N_23388);
nand U26286 (N_26286,N_23583,N_21149);
nand U26287 (N_26287,N_22549,N_23800);
or U26288 (N_26288,N_22562,N_21637);
and U26289 (N_26289,N_23570,N_21740);
nand U26290 (N_26290,N_21253,N_22702);
nor U26291 (N_26291,N_23550,N_21594);
nor U26292 (N_26292,N_21135,N_23023);
or U26293 (N_26293,N_21553,N_23716);
xor U26294 (N_26294,N_21757,N_21413);
xnor U26295 (N_26295,N_21372,N_23292);
nor U26296 (N_26296,N_22046,N_21598);
nand U26297 (N_26297,N_22400,N_23936);
nand U26298 (N_26298,N_21580,N_22131);
xor U26299 (N_26299,N_23911,N_21448);
nand U26300 (N_26300,N_22371,N_23674);
and U26301 (N_26301,N_21046,N_21738);
and U26302 (N_26302,N_23531,N_21160);
and U26303 (N_26303,N_23776,N_23094);
and U26304 (N_26304,N_21187,N_21587);
or U26305 (N_26305,N_21063,N_21618);
and U26306 (N_26306,N_22258,N_21329);
or U26307 (N_26307,N_21083,N_23708);
or U26308 (N_26308,N_22914,N_21086);
nor U26309 (N_26309,N_21556,N_22019);
or U26310 (N_26310,N_21507,N_22109);
nand U26311 (N_26311,N_22858,N_23851);
nor U26312 (N_26312,N_22420,N_22684);
and U26313 (N_26313,N_21499,N_21954);
and U26314 (N_26314,N_21858,N_21221);
or U26315 (N_26315,N_21131,N_23020);
xor U26316 (N_26316,N_22950,N_21138);
or U26317 (N_26317,N_21051,N_22823);
or U26318 (N_26318,N_22505,N_22757);
and U26319 (N_26319,N_23970,N_21172);
or U26320 (N_26320,N_21428,N_22237);
nand U26321 (N_26321,N_21866,N_22298);
nor U26322 (N_26322,N_23818,N_21557);
xnor U26323 (N_26323,N_23411,N_21157);
and U26324 (N_26324,N_22032,N_21023);
and U26325 (N_26325,N_21333,N_22080);
xnor U26326 (N_26326,N_23471,N_22366);
or U26327 (N_26327,N_21102,N_23682);
and U26328 (N_26328,N_22109,N_23128);
nand U26329 (N_26329,N_23178,N_22177);
nand U26330 (N_26330,N_23974,N_22640);
and U26331 (N_26331,N_21576,N_23662);
nor U26332 (N_26332,N_23471,N_21137);
or U26333 (N_26333,N_21071,N_23338);
xnor U26334 (N_26334,N_21615,N_22243);
nand U26335 (N_26335,N_23495,N_23792);
nand U26336 (N_26336,N_22888,N_21254);
nor U26337 (N_26337,N_22277,N_21300);
and U26338 (N_26338,N_21708,N_22408);
or U26339 (N_26339,N_21437,N_21556);
xor U26340 (N_26340,N_21828,N_23713);
nand U26341 (N_26341,N_23807,N_22345);
nor U26342 (N_26342,N_23193,N_21205);
or U26343 (N_26343,N_22351,N_23902);
nand U26344 (N_26344,N_23429,N_21944);
xor U26345 (N_26345,N_22933,N_21844);
nand U26346 (N_26346,N_22037,N_22685);
and U26347 (N_26347,N_23971,N_22620);
and U26348 (N_26348,N_21513,N_22709);
and U26349 (N_26349,N_22512,N_23838);
or U26350 (N_26350,N_21343,N_23766);
nor U26351 (N_26351,N_22615,N_21295);
or U26352 (N_26352,N_23703,N_22517);
and U26353 (N_26353,N_21722,N_23064);
nand U26354 (N_26354,N_21313,N_22716);
xor U26355 (N_26355,N_22746,N_22097);
and U26356 (N_26356,N_21840,N_23222);
nand U26357 (N_26357,N_23529,N_23244);
nor U26358 (N_26358,N_23266,N_22785);
xnor U26359 (N_26359,N_22964,N_21958);
nor U26360 (N_26360,N_21578,N_23316);
xor U26361 (N_26361,N_22374,N_21193);
and U26362 (N_26362,N_22277,N_21006);
nand U26363 (N_26363,N_22837,N_23429);
and U26364 (N_26364,N_23602,N_21477);
xor U26365 (N_26365,N_23502,N_22987);
xor U26366 (N_26366,N_21449,N_22517);
and U26367 (N_26367,N_22630,N_22711);
xor U26368 (N_26368,N_23567,N_22744);
nor U26369 (N_26369,N_23981,N_21947);
nand U26370 (N_26370,N_22571,N_21729);
xnor U26371 (N_26371,N_22885,N_22180);
and U26372 (N_26372,N_23496,N_21281);
nand U26373 (N_26373,N_23596,N_22580);
and U26374 (N_26374,N_22836,N_22660);
or U26375 (N_26375,N_22035,N_23025);
nand U26376 (N_26376,N_22780,N_21094);
nand U26377 (N_26377,N_21040,N_23232);
or U26378 (N_26378,N_21190,N_21604);
and U26379 (N_26379,N_21503,N_23825);
nand U26380 (N_26380,N_22701,N_22770);
nor U26381 (N_26381,N_23036,N_23958);
or U26382 (N_26382,N_21407,N_22951);
xor U26383 (N_26383,N_23306,N_22443);
or U26384 (N_26384,N_21513,N_22595);
xor U26385 (N_26385,N_22232,N_23712);
nand U26386 (N_26386,N_23127,N_22220);
or U26387 (N_26387,N_22535,N_23875);
nand U26388 (N_26388,N_21027,N_21113);
and U26389 (N_26389,N_21074,N_23856);
nor U26390 (N_26390,N_21475,N_21029);
nor U26391 (N_26391,N_21795,N_23672);
or U26392 (N_26392,N_21111,N_22554);
nand U26393 (N_26393,N_21012,N_23058);
nor U26394 (N_26394,N_22079,N_22735);
or U26395 (N_26395,N_22257,N_21784);
xnor U26396 (N_26396,N_23368,N_22948);
and U26397 (N_26397,N_23651,N_21569);
xnor U26398 (N_26398,N_21511,N_21256);
xor U26399 (N_26399,N_21101,N_23391);
xor U26400 (N_26400,N_21433,N_23974);
or U26401 (N_26401,N_22746,N_21839);
nand U26402 (N_26402,N_23000,N_21131);
nor U26403 (N_26403,N_21481,N_23057);
xnor U26404 (N_26404,N_22040,N_22409);
and U26405 (N_26405,N_22825,N_23124);
nor U26406 (N_26406,N_21331,N_23260);
or U26407 (N_26407,N_22963,N_23763);
or U26408 (N_26408,N_21183,N_21942);
nand U26409 (N_26409,N_23453,N_23962);
or U26410 (N_26410,N_21887,N_22683);
xor U26411 (N_26411,N_22180,N_23783);
xnor U26412 (N_26412,N_22608,N_21088);
and U26413 (N_26413,N_23530,N_22154);
and U26414 (N_26414,N_22873,N_21338);
nand U26415 (N_26415,N_21870,N_22016);
xnor U26416 (N_26416,N_22698,N_21449);
or U26417 (N_26417,N_23969,N_23321);
xor U26418 (N_26418,N_21045,N_21626);
and U26419 (N_26419,N_23567,N_23680);
nor U26420 (N_26420,N_22961,N_21347);
or U26421 (N_26421,N_22682,N_21096);
xnor U26422 (N_26422,N_21781,N_23374);
xor U26423 (N_26423,N_22373,N_22059);
nor U26424 (N_26424,N_22932,N_23535);
nand U26425 (N_26425,N_23567,N_23106);
nor U26426 (N_26426,N_21514,N_22738);
or U26427 (N_26427,N_22832,N_23772);
or U26428 (N_26428,N_23588,N_22572);
or U26429 (N_26429,N_23612,N_22100);
or U26430 (N_26430,N_22047,N_21427);
nand U26431 (N_26431,N_23900,N_21783);
xor U26432 (N_26432,N_21765,N_22688);
or U26433 (N_26433,N_23422,N_23283);
and U26434 (N_26434,N_21908,N_21774);
nor U26435 (N_26435,N_23477,N_21825);
nand U26436 (N_26436,N_22600,N_23196);
nand U26437 (N_26437,N_23191,N_21260);
xnor U26438 (N_26438,N_22924,N_22603);
or U26439 (N_26439,N_22717,N_23604);
nand U26440 (N_26440,N_22541,N_22264);
nor U26441 (N_26441,N_22361,N_21153);
or U26442 (N_26442,N_23665,N_22877);
and U26443 (N_26443,N_21703,N_21904);
or U26444 (N_26444,N_21835,N_23378);
and U26445 (N_26445,N_23058,N_22634);
nand U26446 (N_26446,N_22667,N_23403);
and U26447 (N_26447,N_23332,N_22685);
or U26448 (N_26448,N_22429,N_21273);
or U26449 (N_26449,N_22204,N_23031);
xnor U26450 (N_26450,N_22856,N_22142);
nand U26451 (N_26451,N_22818,N_22857);
xnor U26452 (N_26452,N_22013,N_23641);
nand U26453 (N_26453,N_22742,N_23383);
nand U26454 (N_26454,N_21543,N_22195);
or U26455 (N_26455,N_23217,N_23892);
or U26456 (N_26456,N_22085,N_22670);
or U26457 (N_26457,N_21297,N_23542);
nand U26458 (N_26458,N_23849,N_21482);
nand U26459 (N_26459,N_22184,N_22432);
nand U26460 (N_26460,N_22151,N_21941);
xnor U26461 (N_26461,N_23396,N_22637);
or U26462 (N_26462,N_22379,N_23873);
nor U26463 (N_26463,N_21896,N_21913);
xor U26464 (N_26464,N_21258,N_21546);
xor U26465 (N_26465,N_21071,N_22206);
nand U26466 (N_26466,N_23921,N_23136);
nand U26467 (N_26467,N_22487,N_23984);
or U26468 (N_26468,N_23928,N_23195);
or U26469 (N_26469,N_21599,N_22699);
xor U26470 (N_26470,N_22890,N_22327);
nand U26471 (N_26471,N_22451,N_23514);
nor U26472 (N_26472,N_21068,N_21560);
xnor U26473 (N_26473,N_22343,N_22581);
nand U26474 (N_26474,N_23152,N_21893);
and U26475 (N_26475,N_23451,N_23859);
and U26476 (N_26476,N_23715,N_22735);
or U26477 (N_26477,N_21985,N_21291);
nand U26478 (N_26478,N_21856,N_23030);
and U26479 (N_26479,N_21021,N_21331);
and U26480 (N_26480,N_21072,N_22635);
xnor U26481 (N_26481,N_22814,N_21252);
nor U26482 (N_26482,N_23729,N_23151);
or U26483 (N_26483,N_21018,N_23426);
nand U26484 (N_26484,N_23752,N_23865);
xnor U26485 (N_26485,N_23555,N_21056);
nand U26486 (N_26486,N_21015,N_21669);
and U26487 (N_26487,N_22911,N_23189);
nand U26488 (N_26488,N_21882,N_21671);
and U26489 (N_26489,N_21067,N_23954);
nand U26490 (N_26490,N_22081,N_23542);
xor U26491 (N_26491,N_21473,N_21150);
and U26492 (N_26492,N_21119,N_22946);
xnor U26493 (N_26493,N_22213,N_23744);
and U26494 (N_26494,N_21338,N_21709);
nand U26495 (N_26495,N_22525,N_23197);
xor U26496 (N_26496,N_21283,N_22031);
and U26497 (N_26497,N_23374,N_22068);
xnor U26498 (N_26498,N_22951,N_22491);
nor U26499 (N_26499,N_23653,N_21810);
or U26500 (N_26500,N_23525,N_22291);
or U26501 (N_26501,N_21716,N_22163);
xnor U26502 (N_26502,N_23912,N_23526);
and U26503 (N_26503,N_23421,N_22755);
and U26504 (N_26504,N_22356,N_21088);
nand U26505 (N_26505,N_23863,N_23133);
nand U26506 (N_26506,N_22988,N_21890);
and U26507 (N_26507,N_21176,N_21182);
or U26508 (N_26508,N_22099,N_23311);
xor U26509 (N_26509,N_22140,N_23790);
and U26510 (N_26510,N_22466,N_22639);
and U26511 (N_26511,N_21485,N_21701);
nor U26512 (N_26512,N_23166,N_22436);
and U26513 (N_26513,N_22935,N_22955);
nor U26514 (N_26514,N_21356,N_22964);
and U26515 (N_26515,N_21773,N_21703);
and U26516 (N_26516,N_22049,N_23794);
and U26517 (N_26517,N_21901,N_22862);
or U26518 (N_26518,N_23024,N_23652);
or U26519 (N_26519,N_21849,N_22158);
xor U26520 (N_26520,N_21337,N_22276);
and U26521 (N_26521,N_22560,N_23551);
xor U26522 (N_26522,N_22745,N_21463);
nor U26523 (N_26523,N_21393,N_23083);
nand U26524 (N_26524,N_22173,N_21965);
xnor U26525 (N_26525,N_21634,N_21374);
xor U26526 (N_26526,N_23328,N_21971);
xnor U26527 (N_26527,N_23081,N_21256);
and U26528 (N_26528,N_23952,N_23195);
nand U26529 (N_26529,N_22451,N_23838);
xnor U26530 (N_26530,N_23298,N_21588);
nand U26531 (N_26531,N_22548,N_23790);
or U26532 (N_26532,N_21257,N_23157);
nand U26533 (N_26533,N_23772,N_21180);
or U26534 (N_26534,N_23139,N_22337);
nand U26535 (N_26535,N_23359,N_22636);
and U26536 (N_26536,N_22145,N_23829);
nor U26537 (N_26537,N_23370,N_23309);
or U26538 (N_26538,N_23630,N_23542);
or U26539 (N_26539,N_23748,N_21743);
nor U26540 (N_26540,N_21503,N_22265);
and U26541 (N_26541,N_23619,N_21404);
xor U26542 (N_26542,N_21012,N_22444);
or U26543 (N_26543,N_21359,N_22233);
nor U26544 (N_26544,N_23677,N_22214);
nor U26545 (N_26545,N_21452,N_23105);
nand U26546 (N_26546,N_21295,N_22217);
or U26547 (N_26547,N_22210,N_23481);
or U26548 (N_26548,N_21507,N_22835);
nand U26549 (N_26549,N_21340,N_22492);
and U26550 (N_26550,N_23256,N_23584);
nand U26551 (N_26551,N_23857,N_22184);
xnor U26552 (N_26552,N_23371,N_21380);
xnor U26553 (N_26553,N_21084,N_21349);
xnor U26554 (N_26554,N_23923,N_23934);
xor U26555 (N_26555,N_22475,N_21663);
and U26556 (N_26556,N_23164,N_21058);
nand U26557 (N_26557,N_22234,N_21857);
nor U26558 (N_26558,N_21610,N_23857);
nand U26559 (N_26559,N_21957,N_21253);
nor U26560 (N_26560,N_22802,N_23494);
nand U26561 (N_26561,N_21406,N_21283);
nor U26562 (N_26562,N_23394,N_21670);
and U26563 (N_26563,N_23482,N_23607);
and U26564 (N_26564,N_22327,N_22873);
xnor U26565 (N_26565,N_22557,N_23828);
or U26566 (N_26566,N_22077,N_21896);
and U26567 (N_26567,N_23050,N_21749);
nor U26568 (N_26568,N_21683,N_21114);
and U26569 (N_26569,N_22436,N_23026);
nor U26570 (N_26570,N_23184,N_22028);
or U26571 (N_26571,N_23516,N_22807);
nor U26572 (N_26572,N_23067,N_23398);
nand U26573 (N_26573,N_21837,N_23302);
xor U26574 (N_26574,N_23292,N_22791);
nor U26575 (N_26575,N_22444,N_23528);
xnor U26576 (N_26576,N_21995,N_23429);
or U26577 (N_26577,N_22052,N_23358);
xor U26578 (N_26578,N_23074,N_22928);
nand U26579 (N_26579,N_23370,N_21633);
nor U26580 (N_26580,N_22518,N_23424);
nand U26581 (N_26581,N_22857,N_22118);
nand U26582 (N_26582,N_22821,N_23381);
xnor U26583 (N_26583,N_23856,N_21262);
or U26584 (N_26584,N_22813,N_23249);
xnor U26585 (N_26585,N_23873,N_21198);
nor U26586 (N_26586,N_22388,N_22386);
and U26587 (N_26587,N_21014,N_21589);
xor U26588 (N_26588,N_22522,N_23348);
or U26589 (N_26589,N_23792,N_22011);
nand U26590 (N_26590,N_21260,N_21937);
and U26591 (N_26591,N_23350,N_23808);
or U26592 (N_26592,N_23832,N_22563);
nand U26593 (N_26593,N_22404,N_22775);
or U26594 (N_26594,N_22087,N_23688);
or U26595 (N_26595,N_23434,N_23691);
xor U26596 (N_26596,N_22590,N_22375);
and U26597 (N_26597,N_23003,N_23245);
nor U26598 (N_26598,N_23479,N_22901);
xor U26599 (N_26599,N_22957,N_22408);
xnor U26600 (N_26600,N_22542,N_21775);
xnor U26601 (N_26601,N_22053,N_22059);
and U26602 (N_26602,N_21964,N_22647);
nand U26603 (N_26603,N_23475,N_22102);
nor U26604 (N_26604,N_21863,N_21088);
and U26605 (N_26605,N_22023,N_21647);
or U26606 (N_26606,N_22299,N_22875);
or U26607 (N_26607,N_23735,N_22354);
xor U26608 (N_26608,N_22298,N_22955);
xnor U26609 (N_26609,N_21028,N_21304);
nor U26610 (N_26610,N_22785,N_23385);
xnor U26611 (N_26611,N_23188,N_23476);
nor U26612 (N_26612,N_22961,N_23605);
nor U26613 (N_26613,N_23497,N_21652);
nor U26614 (N_26614,N_21239,N_21355);
xor U26615 (N_26615,N_23926,N_22503);
xnor U26616 (N_26616,N_23579,N_22261);
nor U26617 (N_26617,N_22544,N_22109);
nand U26618 (N_26618,N_23325,N_23435);
and U26619 (N_26619,N_22641,N_23768);
xor U26620 (N_26620,N_22382,N_21990);
or U26621 (N_26621,N_23442,N_21495);
xor U26622 (N_26622,N_23972,N_23078);
nor U26623 (N_26623,N_22437,N_22894);
nor U26624 (N_26624,N_23916,N_22791);
and U26625 (N_26625,N_22690,N_21615);
or U26626 (N_26626,N_23161,N_22263);
nand U26627 (N_26627,N_23546,N_22144);
and U26628 (N_26628,N_21821,N_23596);
and U26629 (N_26629,N_23233,N_21657);
nor U26630 (N_26630,N_23769,N_22450);
nor U26631 (N_26631,N_23695,N_23307);
xor U26632 (N_26632,N_22871,N_23280);
nor U26633 (N_26633,N_22207,N_21097);
and U26634 (N_26634,N_22889,N_21659);
and U26635 (N_26635,N_21928,N_21843);
nor U26636 (N_26636,N_23912,N_23315);
nand U26637 (N_26637,N_21424,N_23729);
xor U26638 (N_26638,N_23175,N_21465);
and U26639 (N_26639,N_22665,N_21586);
nor U26640 (N_26640,N_23386,N_23577);
and U26641 (N_26641,N_21506,N_23155);
nor U26642 (N_26642,N_21163,N_23115);
xor U26643 (N_26643,N_23633,N_22591);
nand U26644 (N_26644,N_23674,N_21625);
nand U26645 (N_26645,N_21671,N_23317);
nand U26646 (N_26646,N_23378,N_22234);
or U26647 (N_26647,N_23008,N_21812);
and U26648 (N_26648,N_21802,N_22550);
and U26649 (N_26649,N_22808,N_21094);
and U26650 (N_26650,N_23031,N_21098);
xor U26651 (N_26651,N_21272,N_22843);
xnor U26652 (N_26652,N_21652,N_22888);
nor U26653 (N_26653,N_21500,N_22673);
nand U26654 (N_26654,N_21736,N_23295);
or U26655 (N_26655,N_21238,N_23408);
and U26656 (N_26656,N_23832,N_23118);
nor U26657 (N_26657,N_22233,N_23029);
and U26658 (N_26658,N_21233,N_23362);
nand U26659 (N_26659,N_22474,N_22213);
xor U26660 (N_26660,N_23521,N_21120);
nor U26661 (N_26661,N_21009,N_21773);
xnor U26662 (N_26662,N_21949,N_22102);
nand U26663 (N_26663,N_22778,N_23852);
or U26664 (N_26664,N_22486,N_21768);
or U26665 (N_26665,N_22445,N_21665);
and U26666 (N_26666,N_22331,N_22781);
or U26667 (N_26667,N_21384,N_21203);
and U26668 (N_26668,N_21423,N_21708);
nor U26669 (N_26669,N_21158,N_22023);
xnor U26670 (N_26670,N_23769,N_21176);
and U26671 (N_26671,N_21069,N_21302);
nand U26672 (N_26672,N_22716,N_22808);
or U26673 (N_26673,N_21935,N_21477);
xor U26674 (N_26674,N_23094,N_23737);
xor U26675 (N_26675,N_22564,N_21735);
and U26676 (N_26676,N_23044,N_23928);
nor U26677 (N_26677,N_23923,N_22610);
nor U26678 (N_26678,N_22598,N_23594);
xor U26679 (N_26679,N_23389,N_23254);
nor U26680 (N_26680,N_22730,N_22691);
nor U26681 (N_26681,N_23789,N_23477);
nand U26682 (N_26682,N_21438,N_22763);
or U26683 (N_26683,N_22068,N_22277);
xnor U26684 (N_26684,N_22231,N_22258);
and U26685 (N_26685,N_22144,N_22054);
or U26686 (N_26686,N_22319,N_23944);
and U26687 (N_26687,N_22186,N_23007);
or U26688 (N_26688,N_21940,N_21520);
xor U26689 (N_26689,N_21745,N_21336);
and U26690 (N_26690,N_21195,N_21033);
xor U26691 (N_26691,N_23145,N_21055);
or U26692 (N_26692,N_23044,N_22990);
xnor U26693 (N_26693,N_22385,N_21270);
xor U26694 (N_26694,N_22196,N_21908);
nand U26695 (N_26695,N_22967,N_21709);
nand U26696 (N_26696,N_23533,N_22751);
nand U26697 (N_26697,N_22841,N_23236);
nor U26698 (N_26698,N_21004,N_21257);
or U26699 (N_26699,N_23582,N_23473);
nor U26700 (N_26700,N_23678,N_21730);
nor U26701 (N_26701,N_21707,N_21095);
and U26702 (N_26702,N_23663,N_23656);
nand U26703 (N_26703,N_21235,N_23694);
or U26704 (N_26704,N_22804,N_21116);
xor U26705 (N_26705,N_23785,N_22157);
or U26706 (N_26706,N_23085,N_23761);
nand U26707 (N_26707,N_23483,N_21794);
or U26708 (N_26708,N_22923,N_22550);
or U26709 (N_26709,N_23612,N_22070);
and U26710 (N_26710,N_21937,N_23321);
or U26711 (N_26711,N_22721,N_23734);
and U26712 (N_26712,N_21413,N_21821);
and U26713 (N_26713,N_23056,N_23245);
nand U26714 (N_26714,N_22155,N_23583);
and U26715 (N_26715,N_21009,N_23394);
nand U26716 (N_26716,N_21889,N_22034);
or U26717 (N_26717,N_22692,N_21402);
nor U26718 (N_26718,N_23833,N_21247);
and U26719 (N_26719,N_23404,N_21836);
and U26720 (N_26720,N_22526,N_21357);
nand U26721 (N_26721,N_23217,N_21603);
or U26722 (N_26722,N_21587,N_23825);
or U26723 (N_26723,N_23478,N_22743);
and U26724 (N_26724,N_23782,N_22868);
nand U26725 (N_26725,N_22393,N_21228);
nand U26726 (N_26726,N_21491,N_21821);
nand U26727 (N_26727,N_23911,N_23455);
and U26728 (N_26728,N_21069,N_23720);
and U26729 (N_26729,N_22395,N_23625);
xor U26730 (N_26730,N_22703,N_21668);
nor U26731 (N_26731,N_21357,N_21058);
nand U26732 (N_26732,N_22935,N_22880);
or U26733 (N_26733,N_22167,N_21744);
nor U26734 (N_26734,N_22225,N_21895);
or U26735 (N_26735,N_22257,N_23230);
xor U26736 (N_26736,N_23966,N_21947);
xnor U26737 (N_26737,N_23110,N_23368);
or U26738 (N_26738,N_21060,N_22969);
nor U26739 (N_26739,N_23014,N_22998);
nand U26740 (N_26740,N_23780,N_21176);
nand U26741 (N_26741,N_22255,N_21068);
nand U26742 (N_26742,N_23680,N_22219);
and U26743 (N_26743,N_22060,N_22290);
xor U26744 (N_26744,N_23269,N_23789);
nand U26745 (N_26745,N_21083,N_22184);
nor U26746 (N_26746,N_22668,N_22052);
or U26747 (N_26747,N_23059,N_23905);
nand U26748 (N_26748,N_23157,N_23488);
nand U26749 (N_26749,N_21584,N_23900);
nor U26750 (N_26750,N_21847,N_22419);
nand U26751 (N_26751,N_23230,N_22915);
nor U26752 (N_26752,N_22262,N_22689);
xor U26753 (N_26753,N_23407,N_22391);
and U26754 (N_26754,N_21078,N_22327);
xnor U26755 (N_26755,N_23191,N_21048);
nand U26756 (N_26756,N_22302,N_22390);
xor U26757 (N_26757,N_22506,N_22307);
and U26758 (N_26758,N_21447,N_22819);
nand U26759 (N_26759,N_23355,N_22919);
or U26760 (N_26760,N_21492,N_23962);
and U26761 (N_26761,N_22660,N_22047);
nor U26762 (N_26762,N_22555,N_23588);
nor U26763 (N_26763,N_23942,N_21377);
nand U26764 (N_26764,N_23976,N_22291);
nor U26765 (N_26765,N_21533,N_23201);
or U26766 (N_26766,N_21844,N_22979);
or U26767 (N_26767,N_21494,N_22211);
and U26768 (N_26768,N_21207,N_22632);
nor U26769 (N_26769,N_23054,N_22574);
and U26770 (N_26770,N_21764,N_21335);
nand U26771 (N_26771,N_21570,N_22898);
nand U26772 (N_26772,N_21112,N_23134);
or U26773 (N_26773,N_23460,N_23522);
xnor U26774 (N_26774,N_23086,N_23775);
xor U26775 (N_26775,N_22943,N_21760);
or U26776 (N_26776,N_21393,N_23970);
nand U26777 (N_26777,N_22340,N_21541);
or U26778 (N_26778,N_22680,N_22691);
xnor U26779 (N_26779,N_22757,N_22919);
nor U26780 (N_26780,N_23810,N_22129);
or U26781 (N_26781,N_23960,N_22439);
nand U26782 (N_26782,N_21214,N_21679);
or U26783 (N_26783,N_22431,N_22213);
xor U26784 (N_26784,N_23953,N_21351);
nand U26785 (N_26785,N_21750,N_21795);
or U26786 (N_26786,N_21245,N_23216);
nor U26787 (N_26787,N_21135,N_21131);
and U26788 (N_26788,N_23657,N_21905);
xor U26789 (N_26789,N_22851,N_22463);
nor U26790 (N_26790,N_23635,N_22843);
nor U26791 (N_26791,N_22243,N_22215);
nand U26792 (N_26792,N_22878,N_23651);
or U26793 (N_26793,N_23334,N_23359);
and U26794 (N_26794,N_23291,N_21752);
nand U26795 (N_26795,N_22458,N_22055);
and U26796 (N_26796,N_21792,N_21222);
nor U26797 (N_26797,N_23652,N_21278);
xor U26798 (N_26798,N_23877,N_21643);
nor U26799 (N_26799,N_21995,N_22340);
xor U26800 (N_26800,N_23626,N_23080);
nor U26801 (N_26801,N_22398,N_22200);
or U26802 (N_26802,N_21945,N_22712);
xor U26803 (N_26803,N_22845,N_21061);
and U26804 (N_26804,N_23232,N_21479);
nand U26805 (N_26805,N_23376,N_21671);
or U26806 (N_26806,N_22072,N_22193);
nor U26807 (N_26807,N_23821,N_22363);
nor U26808 (N_26808,N_23027,N_22602);
xnor U26809 (N_26809,N_22787,N_22733);
or U26810 (N_26810,N_21006,N_22740);
and U26811 (N_26811,N_21963,N_23257);
xnor U26812 (N_26812,N_23683,N_22205);
nand U26813 (N_26813,N_23886,N_21490);
and U26814 (N_26814,N_23589,N_23362);
nand U26815 (N_26815,N_21379,N_21101);
or U26816 (N_26816,N_23121,N_21004);
nor U26817 (N_26817,N_22479,N_21235);
nor U26818 (N_26818,N_22620,N_23941);
xor U26819 (N_26819,N_23044,N_22851);
or U26820 (N_26820,N_21969,N_23119);
xnor U26821 (N_26821,N_21580,N_21778);
nor U26822 (N_26822,N_23869,N_21088);
and U26823 (N_26823,N_23712,N_22130);
xor U26824 (N_26824,N_22348,N_22946);
or U26825 (N_26825,N_22018,N_23923);
or U26826 (N_26826,N_23908,N_22053);
nor U26827 (N_26827,N_23023,N_23903);
or U26828 (N_26828,N_22254,N_21568);
nor U26829 (N_26829,N_23350,N_21079);
or U26830 (N_26830,N_21175,N_23426);
xor U26831 (N_26831,N_23196,N_21447);
or U26832 (N_26832,N_21261,N_21250);
nor U26833 (N_26833,N_21097,N_23669);
nand U26834 (N_26834,N_21697,N_21982);
or U26835 (N_26835,N_22922,N_21483);
and U26836 (N_26836,N_22195,N_23923);
nor U26837 (N_26837,N_23394,N_22610);
or U26838 (N_26838,N_23914,N_22004);
xor U26839 (N_26839,N_21791,N_23314);
nand U26840 (N_26840,N_23552,N_22332);
and U26841 (N_26841,N_22262,N_23854);
or U26842 (N_26842,N_22768,N_21291);
or U26843 (N_26843,N_23512,N_21146);
nor U26844 (N_26844,N_21530,N_23851);
nand U26845 (N_26845,N_21299,N_23150);
nor U26846 (N_26846,N_23383,N_22223);
nand U26847 (N_26847,N_21926,N_21765);
or U26848 (N_26848,N_23488,N_23836);
nand U26849 (N_26849,N_22424,N_23198);
and U26850 (N_26850,N_21118,N_21441);
and U26851 (N_26851,N_22230,N_22553);
and U26852 (N_26852,N_21863,N_21154);
or U26853 (N_26853,N_21805,N_21461);
xor U26854 (N_26854,N_21598,N_21257);
or U26855 (N_26855,N_21272,N_21132);
nor U26856 (N_26856,N_22613,N_23655);
nor U26857 (N_26857,N_22133,N_21973);
nor U26858 (N_26858,N_23000,N_23012);
nand U26859 (N_26859,N_22803,N_21803);
or U26860 (N_26860,N_21087,N_22569);
and U26861 (N_26861,N_22279,N_22973);
nor U26862 (N_26862,N_22704,N_22328);
or U26863 (N_26863,N_22976,N_22170);
xor U26864 (N_26864,N_23901,N_23105);
or U26865 (N_26865,N_22651,N_23193);
and U26866 (N_26866,N_21734,N_23652);
xor U26867 (N_26867,N_22363,N_22592);
nand U26868 (N_26868,N_22837,N_23088);
nor U26869 (N_26869,N_23913,N_22871);
xor U26870 (N_26870,N_23684,N_21314);
or U26871 (N_26871,N_22165,N_21212);
nand U26872 (N_26872,N_22713,N_23687);
nor U26873 (N_26873,N_22816,N_22848);
and U26874 (N_26874,N_21361,N_23775);
xnor U26875 (N_26875,N_22062,N_23966);
nor U26876 (N_26876,N_23030,N_23971);
nand U26877 (N_26877,N_21625,N_23763);
nand U26878 (N_26878,N_21090,N_23750);
nand U26879 (N_26879,N_22101,N_21336);
nor U26880 (N_26880,N_23302,N_21524);
and U26881 (N_26881,N_22180,N_21639);
xor U26882 (N_26882,N_23295,N_22590);
and U26883 (N_26883,N_21724,N_23470);
xnor U26884 (N_26884,N_23596,N_22191);
nand U26885 (N_26885,N_23712,N_22789);
xor U26886 (N_26886,N_22258,N_21414);
nand U26887 (N_26887,N_23392,N_22847);
xor U26888 (N_26888,N_22141,N_22207);
xor U26889 (N_26889,N_23267,N_21684);
nand U26890 (N_26890,N_22301,N_22521);
or U26891 (N_26891,N_21925,N_23110);
nor U26892 (N_26892,N_23184,N_23126);
nor U26893 (N_26893,N_23806,N_22221);
and U26894 (N_26894,N_22641,N_22610);
or U26895 (N_26895,N_21063,N_23587);
xnor U26896 (N_26896,N_23387,N_21751);
or U26897 (N_26897,N_23569,N_23141);
or U26898 (N_26898,N_23592,N_21287);
xnor U26899 (N_26899,N_21191,N_23061);
nand U26900 (N_26900,N_21779,N_22484);
xor U26901 (N_26901,N_21196,N_21349);
and U26902 (N_26902,N_21267,N_21360);
xor U26903 (N_26903,N_21057,N_21898);
nor U26904 (N_26904,N_23105,N_23716);
or U26905 (N_26905,N_22406,N_21358);
or U26906 (N_26906,N_21041,N_22633);
and U26907 (N_26907,N_21925,N_22677);
or U26908 (N_26908,N_22634,N_21921);
xnor U26909 (N_26909,N_21457,N_23360);
and U26910 (N_26910,N_23992,N_23890);
nand U26911 (N_26911,N_22416,N_21972);
and U26912 (N_26912,N_22067,N_23215);
xor U26913 (N_26913,N_23797,N_22064);
nand U26914 (N_26914,N_22225,N_21366);
xor U26915 (N_26915,N_22012,N_22889);
xor U26916 (N_26916,N_21315,N_21174);
and U26917 (N_26917,N_22434,N_22295);
and U26918 (N_26918,N_21909,N_23968);
or U26919 (N_26919,N_21656,N_23932);
or U26920 (N_26920,N_22402,N_23339);
xor U26921 (N_26921,N_23770,N_22189);
or U26922 (N_26922,N_21802,N_23884);
xnor U26923 (N_26923,N_23686,N_21909);
or U26924 (N_26924,N_22396,N_22757);
xor U26925 (N_26925,N_23153,N_23822);
nor U26926 (N_26926,N_21121,N_23567);
xor U26927 (N_26927,N_22539,N_22951);
nand U26928 (N_26928,N_23838,N_21389);
nor U26929 (N_26929,N_22245,N_22669);
xnor U26930 (N_26930,N_21354,N_22609);
nand U26931 (N_26931,N_22512,N_22912);
nand U26932 (N_26932,N_22745,N_21167);
xnor U26933 (N_26933,N_21007,N_23528);
nor U26934 (N_26934,N_22997,N_22686);
nand U26935 (N_26935,N_22763,N_22637);
or U26936 (N_26936,N_21959,N_21585);
nand U26937 (N_26937,N_21766,N_23284);
nand U26938 (N_26938,N_22361,N_23412);
nor U26939 (N_26939,N_21830,N_22317);
xnor U26940 (N_26940,N_23168,N_22579);
or U26941 (N_26941,N_21669,N_22599);
and U26942 (N_26942,N_21198,N_23507);
or U26943 (N_26943,N_22757,N_21698);
nand U26944 (N_26944,N_23688,N_22581);
nand U26945 (N_26945,N_23285,N_23259);
and U26946 (N_26946,N_21805,N_22696);
nor U26947 (N_26947,N_22704,N_23022);
nand U26948 (N_26948,N_21083,N_21005);
and U26949 (N_26949,N_21972,N_21841);
nor U26950 (N_26950,N_22277,N_23386);
and U26951 (N_26951,N_23754,N_23078);
or U26952 (N_26952,N_23987,N_23748);
or U26953 (N_26953,N_21657,N_21875);
xnor U26954 (N_26954,N_21847,N_22416);
xor U26955 (N_26955,N_21029,N_21572);
or U26956 (N_26956,N_23802,N_23023);
nor U26957 (N_26957,N_22440,N_21964);
and U26958 (N_26958,N_23869,N_21749);
xor U26959 (N_26959,N_21198,N_23254);
nor U26960 (N_26960,N_21113,N_21383);
xor U26961 (N_26961,N_22885,N_23115);
and U26962 (N_26962,N_23335,N_22730);
nand U26963 (N_26963,N_22144,N_21680);
and U26964 (N_26964,N_22712,N_22904);
nand U26965 (N_26965,N_22558,N_21463);
nand U26966 (N_26966,N_23603,N_21091);
and U26967 (N_26967,N_21509,N_22449);
nand U26968 (N_26968,N_22653,N_22065);
or U26969 (N_26969,N_21028,N_22897);
and U26970 (N_26970,N_22149,N_23968);
nand U26971 (N_26971,N_21118,N_21215);
xor U26972 (N_26972,N_21605,N_22529);
or U26973 (N_26973,N_21633,N_21273);
nand U26974 (N_26974,N_23184,N_21292);
and U26975 (N_26975,N_23941,N_23957);
and U26976 (N_26976,N_22972,N_22606);
nand U26977 (N_26977,N_23803,N_23577);
xnor U26978 (N_26978,N_23111,N_21144);
xor U26979 (N_26979,N_21248,N_21708);
nor U26980 (N_26980,N_23071,N_23906);
or U26981 (N_26981,N_22759,N_23507);
and U26982 (N_26982,N_23132,N_23874);
or U26983 (N_26983,N_22459,N_23209);
and U26984 (N_26984,N_22117,N_22677);
xor U26985 (N_26985,N_21006,N_21277);
and U26986 (N_26986,N_23089,N_22649);
nor U26987 (N_26987,N_22559,N_21621);
nand U26988 (N_26988,N_23838,N_22516);
or U26989 (N_26989,N_21187,N_21605);
nor U26990 (N_26990,N_23809,N_23671);
or U26991 (N_26991,N_21245,N_21775);
or U26992 (N_26992,N_22956,N_21706);
xnor U26993 (N_26993,N_22867,N_22972);
nor U26994 (N_26994,N_23768,N_21673);
and U26995 (N_26995,N_22224,N_22488);
or U26996 (N_26996,N_22855,N_22911);
xor U26997 (N_26997,N_22974,N_22539);
or U26998 (N_26998,N_23321,N_21461);
nand U26999 (N_26999,N_22129,N_22265);
xnor U27000 (N_27000,N_26656,N_25656);
nor U27001 (N_27001,N_26983,N_26664);
xnor U27002 (N_27002,N_24937,N_26819);
nor U27003 (N_27003,N_25960,N_24668);
and U27004 (N_27004,N_26885,N_24911);
or U27005 (N_27005,N_25335,N_26073);
or U27006 (N_27006,N_25050,N_24477);
nor U27007 (N_27007,N_25836,N_25721);
or U27008 (N_27008,N_24346,N_24222);
xor U27009 (N_27009,N_26807,N_25563);
nor U27010 (N_27010,N_24510,N_24427);
nor U27011 (N_27011,N_24159,N_25257);
or U27012 (N_27012,N_25436,N_26641);
and U27013 (N_27013,N_26206,N_25585);
nand U27014 (N_27014,N_25916,N_24639);
nor U27015 (N_27015,N_26563,N_25028);
or U27016 (N_27016,N_26343,N_25073);
xor U27017 (N_27017,N_26064,N_24979);
nand U27018 (N_27018,N_25030,N_25822);
nor U27019 (N_27019,N_26537,N_24219);
xnor U27020 (N_27020,N_25885,N_24662);
xnor U27021 (N_27021,N_24015,N_26487);
nor U27022 (N_27022,N_25285,N_25104);
and U27023 (N_27023,N_25423,N_24268);
and U27024 (N_27024,N_26663,N_24380);
nand U27025 (N_27025,N_26801,N_26741);
xor U27026 (N_27026,N_25988,N_26418);
nor U27027 (N_27027,N_24103,N_24749);
or U27028 (N_27028,N_25823,N_24040);
nor U27029 (N_27029,N_26749,N_25473);
or U27030 (N_27030,N_25735,N_26455);
xnor U27031 (N_27031,N_24616,N_26146);
nand U27032 (N_27032,N_25930,N_25839);
nand U27033 (N_27033,N_26758,N_25550);
nand U27034 (N_27034,N_25158,N_25455);
or U27035 (N_27035,N_25990,N_25259);
nor U27036 (N_27036,N_26248,N_26264);
nor U27037 (N_27037,N_25818,N_25289);
and U27038 (N_27038,N_26800,N_25901);
xnor U27039 (N_27039,N_25250,N_26864);
xnor U27040 (N_27040,N_26934,N_26679);
and U27041 (N_27041,N_26292,N_24963);
nand U27042 (N_27042,N_25309,N_26545);
nor U27043 (N_27043,N_26133,N_26902);
and U27044 (N_27044,N_24318,N_25382);
xnor U27045 (N_27045,N_25597,N_25451);
or U27046 (N_27046,N_26125,N_26151);
xor U27047 (N_27047,N_26899,N_26592);
or U27048 (N_27048,N_25861,N_24025);
nor U27049 (N_27049,N_24468,N_24488);
xor U27050 (N_27050,N_25044,N_24323);
nand U27051 (N_27051,N_25185,N_26927);
and U27052 (N_27052,N_25182,N_24795);
nor U27053 (N_27053,N_25083,N_24415);
nor U27054 (N_27054,N_25280,N_26039);
nor U27055 (N_27055,N_25165,N_26478);
nor U27056 (N_27056,N_25790,N_26752);
xor U27057 (N_27057,N_25814,N_25704);
and U27058 (N_27058,N_26481,N_26972);
xnor U27059 (N_27059,N_25487,N_24532);
or U27060 (N_27060,N_25359,N_25346);
and U27061 (N_27061,N_24231,N_24332);
and U27062 (N_27062,N_25511,N_24029);
or U27063 (N_27063,N_24600,N_25838);
nand U27064 (N_27064,N_25594,N_26168);
xor U27065 (N_27065,N_25931,N_24754);
nand U27066 (N_27066,N_26591,N_24619);
nor U27067 (N_27067,N_26525,N_24392);
nor U27068 (N_27068,N_26070,N_25323);
nor U27069 (N_27069,N_26636,N_25903);
nand U27070 (N_27070,N_26862,N_24958);
and U27071 (N_27071,N_25040,N_25884);
nand U27072 (N_27072,N_24939,N_25048);
or U27073 (N_27073,N_26737,N_24317);
or U27074 (N_27074,N_26470,N_25488);
nor U27075 (N_27075,N_24558,N_25767);
xor U27076 (N_27076,N_26669,N_26678);
or U27077 (N_27077,N_26342,N_24178);
nand U27078 (N_27078,N_25015,N_25986);
or U27079 (N_27079,N_25649,N_25234);
xor U27080 (N_27080,N_26102,N_26281);
and U27081 (N_27081,N_24553,N_26124);
xor U27082 (N_27082,N_26409,N_25366);
xor U27083 (N_27083,N_24110,N_25776);
xnor U27084 (N_27084,N_25208,N_26345);
and U27085 (N_27085,N_24880,N_26658);
xnor U27086 (N_27086,N_25755,N_26650);
and U27087 (N_27087,N_26093,N_24202);
or U27088 (N_27088,N_24345,N_26619);
nor U27089 (N_27089,N_24854,N_24820);
nand U27090 (N_27090,N_24512,N_25624);
nor U27091 (N_27091,N_24129,N_26831);
or U27092 (N_27092,N_25342,N_25622);
or U27093 (N_27093,N_26384,N_24618);
and U27094 (N_27094,N_24076,N_25940);
or U27095 (N_27095,N_26869,N_24931);
xnor U27096 (N_27096,N_26379,N_25004);
and U27097 (N_27097,N_25019,N_25750);
or U27098 (N_27098,N_26310,N_24849);
xor U27099 (N_27099,N_24506,N_24357);
nand U27100 (N_27100,N_25315,N_24206);
and U27101 (N_27101,N_25085,N_25377);
nand U27102 (N_27102,N_25059,N_26994);
and U27103 (N_27103,N_24746,N_25218);
xnor U27104 (N_27104,N_26611,N_24727);
and U27105 (N_27105,N_24060,N_26244);
and U27106 (N_27106,N_24166,N_26405);
or U27107 (N_27107,N_24570,N_26322);
xor U27108 (N_27108,N_25586,N_24130);
nor U27109 (N_27109,N_24423,N_24478);
nor U27110 (N_27110,N_25950,N_26539);
or U27111 (N_27111,N_25422,N_26683);
or U27112 (N_27112,N_25066,N_24261);
nand U27113 (N_27113,N_26031,N_25949);
or U27114 (N_27114,N_25567,N_25754);
xnor U27115 (N_27115,N_25322,N_26984);
and U27116 (N_27116,N_24943,N_26736);
nor U27117 (N_27117,N_25592,N_26645);
and U27118 (N_27118,N_25316,N_26453);
xnor U27119 (N_27119,N_25490,N_26498);
xnor U27120 (N_27120,N_26458,N_24112);
nand U27121 (N_27121,N_26180,N_25596);
or U27122 (N_27122,N_25768,N_25363);
and U27123 (N_27123,N_26931,N_24882);
xnor U27124 (N_27124,N_24455,N_24235);
nor U27125 (N_27125,N_25731,N_24364);
xor U27126 (N_27126,N_25393,N_24243);
xnor U27127 (N_27127,N_24590,N_24004);
and U27128 (N_27128,N_25039,N_24888);
nand U27129 (N_27129,N_25527,N_26744);
nand U27130 (N_27130,N_26260,N_25661);
nor U27131 (N_27131,N_26193,N_25094);
nand U27132 (N_27132,N_26456,N_24155);
or U27133 (N_27133,N_24960,N_26940);
and U27134 (N_27134,N_24709,N_25320);
or U27135 (N_27135,N_25896,N_24733);
nor U27136 (N_27136,N_25432,N_26840);
nand U27137 (N_27137,N_25389,N_25482);
and U27138 (N_27138,N_24424,N_25435);
xor U27139 (N_27139,N_26859,N_26370);
nand U27140 (N_27140,N_24999,N_26485);
nor U27141 (N_27141,N_26414,N_24615);
nand U27142 (N_27142,N_26060,N_25474);
or U27143 (N_27143,N_25225,N_26794);
and U27144 (N_27144,N_25395,N_26337);
nand U27145 (N_27145,N_25114,N_24414);
or U27146 (N_27146,N_26078,N_24355);
nand U27147 (N_27147,N_25404,N_26399);
xnor U27148 (N_27148,N_25466,N_25353);
or U27149 (N_27149,N_25054,N_26044);
and U27150 (N_27150,N_25708,N_26305);
or U27151 (N_27151,N_25715,N_24843);
xor U27152 (N_27152,N_24870,N_26547);
nor U27153 (N_27153,N_25464,N_26171);
nand U27154 (N_27154,N_26430,N_26085);
xor U27155 (N_27155,N_24201,N_24751);
nand U27156 (N_27156,N_24578,N_26142);
xnor U27157 (N_27157,N_25305,N_26394);
xor U27158 (N_27158,N_26770,N_26585);
nand U27159 (N_27159,N_26989,N_26556);
nand U27160 (N_27160,N_25443,N_25747);
xnor U27161 (N_27161,N_25888,N_24818);
or U27162 (N_27162,N_25993,N_25440);
xor U27163 (N_27163,N_26668,N_26375);
xnor U27164 (N_27164,N_24139,N_26190);
and U27165 (N_27165,N_26195,N_24366);
or U27166 (N_27166,N_24951,N_25340);
or U27167 (N_27167,N_26564,N_25425);
or U27168 (N_27168,N_26858,N_26063);
xor U27169 (N_27169,N_26883,N_24731);
and U27170 (N_27170,N_25573,N_24518);
nand U27171 (N_27171,N_24347,N_26482);
xnor U27172 (N_27172,N_26835,N_26480);
xor U27173 (N_27173,N_25100,N_24724);
nand U27174 (N_27174,N_26640,N_26299);
xor U27175 (N_27175,N_24292,N_25235);
and U27176 (N_27176,N_25079,N_24714);
xnor U27177 (N_27177,N_25113,N_24428);
or U27178 (N_27178,N_24856,N_26250);
nand U27179 (N_27179,N_26030,N_26170);
and U27180 (N_27180,N_26763,N_24790);
nor U27181 (N_27181,N_25133,N_25697);
nor U27182 (N_27182,N_25918,N_25426);
xor U27183 (N_27183,N_25530,N_25557);
xor U27184 (N_27184,N_24565,N_26287);
and U27185 (N_27185,N_26968,N_25992);
nor U27186 (N_27186,N_26369,N_24371);
nand U27187 (N_27187,N_24990,N_25064);
xnor U27188 (N_27188,N_24124,N_24555);
or U27189 (N_27189,N_25175,N_24383);
xnor U27190 (N_27190,N_26357,N_24150);
xnor U27191 (N_27191,N_25043,N_26410);
nand U27192 (N_27192,N_24629,N_25484);
or U27193 (N_27193,N_25688,N_24324);
xnor U27194 (N_27194,N_25303,N_25271);
xor U27195 (N_27195,N_26526,N_24370);
and U27196 (N_27196,N_25685,N_24322);
xnor U27197 (N_27197,N_24230,N_25061);
xnor U27198 (N_27198,N_26340,N_26602);
or U27199 (N_27199,N_25765,N_25506);
nor U27200 (N_27200,N_24598,N_26175);
and U27201 (N_27201,N_26542,N_24788);
nand U27202 (N_27202,N_26049,N_26684);
nor U27203 (N_27203,N_24961,N_24100);
or U27204 (N_27204,N_26432,N_26870);
and U27205 (N_27205,N_25817,N_25576);
xnor U27206 (N_27206,N_25087,N_25304);
nor U27207 (N_27207,N_25878,N_26075);
or U27208 (N_27208,N_24403,N_25429);
nand U27209 (N_27209,N_25621,N_24906);
nor U27210 (N_27210,N_25101,N_25779);
and U27211 (N_27211,N_25266,N_25716);
nor U27212 (N_27212,N_26690,N_26372);
nand U27213 (N_27213,N_26492,N_26224);
nand U27214 (N_27214,N_25135,N_24650);
xnor U27215 (N_27215,N_26086,N_26423);
xor U27216 (N_27216,N_24592,N_24752);
nand U27217 (N_27217,N_25778,N_24624);
nor U27218 (N_27218,N_24607,N_25760);
or U27219 (N_27219,N_26944,N_24390);
nand U27220 (N_27220,N_25543,N_26953);
nand U27221 (N_27221,N_24812,N_26134);
nor U27222 (N_27222,N_24376,N_25198);
nand U27223 (N_27223,N_26903,N_24011);
and U27224 (N_27224,N_26079,N_26301);
nor U27225 (N_27225,N_26554,N_25883);
or U27226 (N_27226,N_25577,N_24059);
nor U27227 (N_27227,N_24244,N_26757);
nor U27228 (N_27228,N_24576,N_25179);
and U27229 (N_27229,N_26583,N_26576);
xnor U27230 (N_27230,N_26397,N_24012);
nand U27231 (N_27231,N_26980,N_25739);
nand U27232 (N_27232,N_25086,N_25841);
nand U27233 (N_27233,N_25427,N_26852);
or U27234 (N_27234,N_26336,N_26601);
nand U27235 (N_27235,N_24688,N_24877);
or U27236 (N_27236,N_26661,N_24815);
xor U27237 (N_27237,N_26028,N_24726);
nand U27238 (N_27238,N_25651,N_25437);
and U27239 (N_27239,N_25991,N_25869);
nand U27240 (N_27240,N_24435,N_26966);
xor U27241 (N_27241,N_25772,N_25223);
and U27242 (N_27242,N_25994,N_26303);
xor U27243 (N_27243,N_24045,N_26797);
nor U27244 (N_27244,N_25997,N_24096);
nor U27245 (N_27245,N_24338,N_25021);
or U27246 (N_27246,N_24548,N_25889);
or U27247 (N_27247,N_26255,N_24282);
xor U27248 (N_27248,N_25411,N_25169);
xor U27249 (N_27249,N_24036,N_26251);
nand U27250 (N_27250,N_24504,N_26326);
xnor U27251 (N_27251,N_26766,N_24115);
or U27252 (N_27252,N_25345,N_24388);
xor U27253 (N_27253,N_26330,N_24702);
xor U27254 (N_27254,N_24881,N_26892);
and U27255 (N_27255,N_25671,N_24396);
xor U27256 (N_27256,N_25391,N_26383);
nor U27257 (N_27257,N_25695,N_24509);
nand U27258 (N_27258,N_25684,N_25191);
nor U27259 (N_27259,N_24687,N_25682);
nand U27260 (N_27260,N_24145,N_25240);
or U27261 (N_27261,N_25080,N_24902);
or U27262 (N_27262,N_25801,N_25452);
nor U27263 (N_27263,N_24678,N_24883);
or U27264 (N_27264,N_25745,N_26693);
nand U27265 (N_27265,N_24511,N_24407);
and U27266 (N_27266,N_26388,N_26227);
nand U27267 (N_27267,N_24101,N_24940);
nand U27268 (N_27268,N_24360,N_26876);
nand U27269 (N_27269,N_24944,N_24462);
and U27270 (N_27270,N_24467,N_26176);
nand U27271 (N_27271,N_26138,N_26448);
and U27272 (N_27272,N_25270,N_26694);
xnor U27273 (N_27273,N_26768,N_25536);
nor U27274 (N_27274,N_25262,N_26426);
and U27275 (N_27275,N_24343,N_26841);
nand U27276 (N_27276,N_24711,N_26197);
nand U27277 (N_27277,N_25770,N_25385);
and U27278 (N_27278,N_26446,N_25007);
xor U27279 (N_27279,N_24801,N_25691);
xnor U27280 (N_27280,N_24568,N_25851);
and U27281 (N_27281,N_25144,N_25663);
and U27282 (N_27282,N_24665,N_26726);
nand U27283 (N_27283,N_25789,N_25176);
nand U27284 (N_27284,N_26377,N_25927);
nand U27285 (N_27285,N_26089,N_24051);
and U27286 (N_27286,N_24573,N_24251);
nand U27287 (N_27287,N_24846,N_24766);
or U27288 (N_27288,N_24156,N_25381);
or U27289 (N_27289,N_25917,N_24238);
or U27290 (N_27290,N_25512,N_24194);
nor U27291 (N_27291,N_25036,N_24102);
xnor U27292 (N_27292,N_25729,N_26135);
or U27293 (N_27293,N_24748,N_25867);
nor U27294 (N_27294,N_26703,N_24917);
xor U27295 (N_27295,N_26643,N_26024);
xnor U27296 (N_27296,N_26291,N_25204);
nor U27297 (N_27297,N_24104,N_25648);
nand U27298 (N_27298,N_24262,N_24168);
nor U27299 (N_27299,N_25909,N_26895);
xor U27300 (N_27300,N_24701,N_26930);
nor U27301 (N_27301,N_26762,N_25654);
or U27302 (N_27302,N_26905,N_25753);
nor U27303 (N_27303,N_24485,N_24273);
nor U27304 (N_27304,N_25633,N_25063);
and U27305 (N_27305,N_24740,N_25496);
nor U27306 (N_27306,N_25367,N_25650);
nand U27307 (N_27307,N_25792,N_24526);
and U27308 (N_27308,N_24158,N_24184);
nor U27309 (N_27309,N_24919,N_24476);
xnor U27310 (N_27310,N_25141,N_26932);
xor U27311 (N_27311,N_24704,N_25026);
nand U27312 (N_27312,N_26220,N_25400);
and U27313 (N_27313,N_26567,N_25072);
nor U27314 (N_27314,N_24493,N_24779);
nor U27315 (N_27315,N_24637,N_24456);
or U27316 (N_27316,N_24452,N_26366);
nor U27317 (N_27317,N_26472,N_26698);
nand U27318 (N_27318,N_24368,N_24369);
xnor U27319 (N_27319,N_24429,N_24020);
and U27320 (N_27320,N_24806,N_24128);
and U27321 (N_27321,N_25293,N_26033);
nor U27322 (N_27322,N_24792,N_25439);
nor U27323 (N_27323,N_24609,N_24807);
nand U27324 (N_27324,N_24442,N_26471);
nand U27325 (N_27325,N_24413,N_24461);
and U27326 (N_27326,N_24628,N_26155);
xnor U27327 (N_27327,N_26850,N_24387);
nand U27328 (N_27328,N_26475,N_24621);
or U27329 (N_27329,N_25572,N_25636);
nand U27330 (N_27330,N_25955,N_24564);
nand U27331 (N_27331,N_26952,N_26211);
and U27332 (N_27332,N_26181,N_24196);
xnor U27333 (N_27333,N_26697,N_24786);
xnor U27334 (N_27334,N_25812,N_24861);
xnor U27335 (N_27335,N_24667,N_24460);
xnor U27336 (N_27336,N_26925,N_25614);
and U27337 (N_27337,N_26507,N_24361);
nor U27338 (N_27338,N_24533,N_26574);
or U27339 (N_27339,N_25607,N_24250);
nand U27340 (N_27340,N_25540,N_26167);
nand U27341 (N_27341,N_26112,N_24777);
or U27342 (N_27342,N_25447,N_25816);
or U27343 (N_27343,N_24897,N_24562);
nor U27344 (N_27344,N_25160,N_25161);
xor U27345 (N_27345,N_24402,N_24271);
nor U27346 (N_27346,N_24860,N_25479);
nor U27347 (N_27347,N_26416,N_26177);
and U27348 (N_27348,N_26381,N_26532);
nor U27349 (N_27349,N_25001,N_26404);
and U27350 (N_27350,N_25388,N_25922);
xor U27351 (N_27351,N_24329,N_26243);
nor U27352 (N_27352,N_25970,N_26047);
or U27353 (N_27353,N_25683,N_24984);
or U27354 (N_27354,N_25372,N_26214);
nor U27355 (N_27355,N_24125,N_24082);
nor U27356 (N_27356,N_24254,N_24337);
nor U27357 (N_27357,N_24671,N_24116);
nor U27358 (N_27358,N_26438,N_24247);
nor U27359 (N_27359,N_24647,N_24947);
nand U27360 (N_27360,N_24137,N_25219);
nand U27361 (N_27361,N_25774,N_25402);
nor U27362 (N_27362,N_26385,N_25678);
xor U27363 (N_27363,N_25355,N_24126);
nand U27364 (N_27364,N_26374,N_24108);
or U27365 (N_27365,N_25127,N_24813);
xnor U27366 (N_27366,N_25310,N_26692);
xor U27367 (N_27367,N_26897,N_24430);
nor U27368 (N_27368,N_24018,N_25249);
and U27369 (N_27369,N_25620,N_25053);
nor U27370 (N_27370,N_25016,N_24715);
nor U27371 (N_27371,N_24094,N_24031);
xor U27372 (N_27372,N_26530,N_25207);
and U27373 (N_27373,N_24655,N_24022);
and U27374 (N_27374,N_26502,N_24622);
and U27375 (N_27375,N_26077,N_24585);
xnor U27376 (N_27376,N_24470,N_24342);
or U27377 (N_27377,N_24448,N_25166);
or U27378 (N_27378,N_25498,N_26313);
or U27379 (N_27379,N_24320,N_25000);
or U27380 (N_27380,N_24956,N_25926);
and U27381 (N_27381,N_24287,N_26083);
nand U27382 (N_27382,N_24669,N_24459);
and U27383 (N_27383,N_25687,N_24188);
nand U27384 (N_27384,N_26868,N_26116);
or U27385 (N_27385,N_24105,N_26958);
and U27386 (N_27386,N_24087,N_24024);
or U27387 (N_27387,N_26734,N_24758);
nor U27388 (N_27388,N_24418,N_26199);
and U27389 (N_27389,N_25583,N_25842);
and U27390 (N_27390,N_24062,N_26445);
or U27391 (N_27391,N_26731,N_24541);
nor U27392 (N_27392,N_25174,N_26578);
nand U27393 (N_27393,N_24341,N_25291);
and U27394 (N_27394,N_25740,N_24301);
nor U27395 (N_27395,N_26769,N_25863);
nor U27396 (N_27396,N_24875,N_25494);
nand U27397 (N_27397,N_25775,N_25424);
xor U27398 (N_27398,N_25507,N_25153);
xnor U27399 (N_27399,N_25813,N_25590);
nand U27400 (N_27400,N_24569,N_26058);
or U27401 (N_27401,N_24484,N_26657);
or U27402 (N_27402,N_26778,N_25416);
nand U27403 (N_27403,N_24398,N_25757);
nand U27404 (N_27404,N_24177,N_26237);
and U27405 (N_27405,N_24953,N_24379);
nand U27406 (N_27406,N_25787,N_25741);
nand U27407 (N_27407,N_25122,N_26950);
nor U27408 (N_27408,N_26393,N_24039);
and U27409 (N_27409,N_25508,N_24646);
nand U27410 (N_27410,N_25460,N_25503);
xnor U27411 (N_27411,N_24088,N_24674);
nand U27412 (N_27412,N_24508,N_24771);
nand U27413 (N_27413,N_26879,N_25800);
or U27414 (N_27414,N_24068,N_25211);
nor U27415 (N_27415,N_26017,N_25606);
and U27416 (N_27416,N_25184,N_25037);
nor U27417 (N_27417,N_24679,N_26050);
and U27418 (N_27418,N_25628,N_24385);
or U27419 (N_27419,N_26750,N_25568);
nor U27420 (N_27420,N_25873,N_25358);
and U27421 (N_27421,N_26121,N_24998);
xor U27422 (N_27422,N_25780,N_25971);
and U27423 (N_27423,N_24146,N_26854);
or U27424 (N_27424,N_25216,N_26558);
nor U27425 (N_27425,N_24874,N_24141);
or U27426 (N_27426,N_24010,N_26117);
nor U27427 (N_27427,N_24938,N_26904);
nor U27428 (N_27428,N_24153,N_24651);
or U27429 (N_27429,N_26610,N_26202);
nor U27430 (N_27430,N_26739,N_24181);
or U27431 (N_27431,N_26837,N_24695);
and U27432 (N_27432,N_26725,N_25111);
or U27433 (N_27433,N_24930,N_25977);
nor U27434 (N_27434,N_26184,N_26436);
xor U27435 (N_27435,N_25870,N_25777);
xnor U27436 (N_27436,N_25398,N_26926);
xnor U27437 (N_27437,N_26920,N_26522);
nand U27438 (N_27438,N_24474,N_25237);
xor U27439 (N_27439,N_25008,N_26246);
nor U27440 (N_27440,N_26524,N_25170);
and U27441 (N_27441,N_26939,N_26666);
nor U27442 (N_27442,N_25613,N_26293);
or U27443 (N_27443,N_25337,N_26270);
or U27444 (N_27444,N_24492,N_24069);
nor U27445 (N_27445,N_25420,N_24743);
and U27446 (N_27446,N_26252,N_24255);
nor U27447 (N_27447,N_26579,N_24694);
or U27448 (N_27448,N_24842,N_25545);
xor U27449 (N_27449,N_25706,N_24315);
nor U27450 (N_27450,N_26154,N_24725);
nand U27451 (N_27451,N_26978,N_24197);
and U27452 (N_27452,N_25513,N_25055);
and U27453 (N_27453,N_26976,N_24374);
nand U27454 (N_27454,N_25071,N_25587);
or U27455 (N_27455,N_26829,N_26160);
nor U27456 (N_27456,N_26391,N_26594);
xor U27457 (N_27457,N_25020,N_25475);
nor U27458 (N_27458,N_25049,N_26126);
nor U27459 (N_27459,N_26511,N_24584);
and U27460 (N_27460,N_25296,N_26013);
nand U27461 (N_27461,N_24982,N_26973);
nand U27462 (N_27462,N_24378,N_26598);
and U27463 (N_27463,N_24910,N_24421);
nand U27464 (N_27464,N_24784,N_25042);
xnor U27465 (N_27465,N_24079,N_26857);
xor U27466 (N_27466,N_26921,N_24642);
xor U27467 (N_27467,N_26347,N_25632);
nand U27468 (N_27468,N_25657,N_24959);
nand U27469 (N_27469,N_25689,N_26802);
xor U27470 (N_27470,N_25268,N_24965);
xnor U27471 (N_27471,N_25705,N_24234);
and U27472 (N_27472,N_25603,N_25953);
nor U27473 (N_27473,N_25876,N_26667);
or U27474 (N_27474,N_25564,N_25928);
or U27475 (N_27475,N_25921,N_26584);
or U27476 (N_27476,N_25478,N_26285);
xnor U27477 (N_27477,N_25961,N_26479);
nor U27478 (N_27478,N_24524,N_25941);
xor U27479 (N_27479,N_26531,N_26833);
or U27480 (N_27480,N_24450,N_25840);
nor U27481 (N_27481,N_25062,N_24325);
or U27482 (N_27482,N_26463,N_25676);
or U27483 (N_27483,N_24835,N_25306);
or U27484 (N_27484,N_26639,N_26911);
or U27485 (N_27485,N_26842,N_26396);
and U27486 (N_27486,N_24353,N_24540);
nand U27487 (N_27487,N_24957,N_24966);
or U27488 (N_27488,N_25441,N_24972);
nand U27489 (N_27489,N_25858,N_25277);
nand U27490 (N_27490,N_25091,N_25319);
and U27491 (N_27491,N_24226,N_24213);
nor U27492 (N_27492,N_24187,N_26331);
nand U27493 (N_27493,N_26137,N_26359);
and U27494 (N_27494,N_26907,N_26900);
nor U27495 (N_27495,N_26424,N_26182);
xor U27496 (N_27496,N_26501,N_26543);
and U27497 (N_27497,N_26915,N_24408);
or U27498 (N_27498,N_25384,N_25292);
xnor U27499 (N_27499,N_25793,N_25022);
nor U27500 (N_27500,N_24593,N_24041);
nor U27501 (N_27501,N_25421,N_26462);
nor U27502 (N_27502,N_26200,N_26304);
or U27503 (N_27503,N_25089,N_24992);
and U27504 (N_27504,N_24502,N_25092);
or U27505 (N_27505,N_24279,N_25502);
nor U27506 (N_27506,N_26977,N_26056);
and U27507 (N_27507,N_26887,N_26685);
and U27508 (N_27508,N_26843,N_26041);
xor U27509 (N_27509,N_25565,N_24176);
xor U27510 (N_27510,N_24149,N_25963);
and U27511 (N_27511,N_24719,N_26130);
or U27512 (N_27512,N_24469,N_26386);
nor U27513 (N_27513,N_26474,N_25915);
xnor U27514 (N_27514,N_24433,N_24871);
nand U27515 (N_27515,N_24117,N_26630);
nand U27516 (N_27516,N_24969,N_26395);
or U27517 (N_27517,N_26091,N_26699);
nor U27518 (N_27518,N_25205,N_25908);
nor U27519 (N_27519,N_25515,N_24297);
nor U27520 (N_27520,N_24974,N_25520);
or U27521 (N_27521,N_26551,N_24797);
xnor U27522 (N_27522,N_26365,N_26942);
nor U27523 (N_27523,N_26625,N_24422);
xor U27524 (N_27524,N_26234,N_24498);
and U27525 (N_27525,N_25253,N_25177);
or U27526 (N_27526,N_24935,N_26018);
and U27527 (N_27527,N_25333,N_25875);
and U27528 (N_27528,N_25137,N_26101);
xnor U27529 (N_27529,N_25407,N_26004);
nand U27530 (N_27530,N_26269,N_25699);
nand U27531 (N_27531,N_26228,N_25276);
nand U27532 (N_27532,N_26354,N_26705);
nor U27533 (N_27533,N_24192,N_26732);
and U27534 (N_27534,N_25213,N_24144);
and U27535 (N_27535,N_26748,N_25431);
nor U27536 (N_27536,N_25217,N_25756);
xnor U27537 (N_27537,N_26527,N_25625);
nor U27538 (N_27538,N_25919,N_24789);
nor U27539 (N_27539,N_26993,N_24863);
or U27540 (N_27540,N_26568,N_26027);
or U27541 (N_27541,N_24803,N_24723);
and U27542 (N_27542,N_26913,N_26296);
or U27543 (N_27543,N_26662,N_24419);
xnor U27544 (N_27544,N_25764,N_24095);
nand U27545 (N_27545,N_24107,N_26817);
nand U27546 (N_27546,N_26933,N_25701);
xor U27547 (N_27547,N_26371,N_24827);
nor U27548 (N_27548,N_25599,N_25338);
or U27549 (N_27549,N_26586,N_26235);
or U27550 (N_27550,N_25645,N_24527);
nand U27551 (N_27551,N_25295,N_25032);
xnor U27552 (N_27552,N_26320,N_25962);
and U27553 (N_27553,N_26593,N_26622);
and U27554 (N_27554,N_26552,N_25522);
nand U27555 (N_27555,N_24934,N_26443);
and U27556 (N_27556,N_25312,N_26729);
nand U27557 (N_27557,N_25379,N_25944);
nand U27558 (N_27558,N_24458,N_26136);
nand U27559 (N_27559,N_24349,N_25396);
nand U27560 (N_27560,N_24599,N_26431);
and U27561 (N_27561,N_25251,N_25525);
xor U27562 (N_27562,N_24926,N_26755);
or U27563 (N_27563,N_25958,N_26439);
and U27564 (N_27564,N_26290,N_26107);
or U27565 (N_27565,N_25692,N_25084);
nor U27566 (N_27566,N_24823,N_26286);
xor U27567 (N_27567,N_26187,N_24109);
and U27568 (N_27568,N_26790,N_25414);
or U27569 (N_27569,N_25445,N_24248);
or U27570 (N_27570,N_25611,N_26131);
xnor U27571 (N_27571,N_24252,N_26995);
and U27572 (N_27572,N_24073,N_24259);
or U27573 (N_27573,N_26888,N_26295);
or U27574 (N_27574,N_25635,N_25149);
nand U27575 (N_27575,N_26258,N_26680);
xnor U27576 (N_27576,N_25453,N_24967);
nor U27577 (N_27577,N_25588,N_25535);
xor U27578 (N_27578,N_26449,N_26886);
xor U27579 (N_27579,N_26057,N_25349);
xor U27580 (N_27580,N_25227,N_26889);
and U27581 (N_27581,N_26959,N_24348);
nor U27582 (N_27582,N_25832,N_26398);
or U27583 (N_27583,N_24840,N_24265);
xnor U27584 (N_27584,N_24898,N_24805);
or U27585 (N_27585,N_26451,N_26569);
or U27586 (N_27586,N_24334,N_25344);
and U27587 (N_27587,N_25107,N_24365);
or U27588 (N_27588,N_25328,N_24114);
nand U27589 (N_27589,N_26508,N_26623);
nor U27590 (N_27590,N_25698,N_26420);
xor U27591 (N_27591,N_24229,N_24057);
nor U27592 (N_27592,N_26087,N_25202);
and U27593 (N_27593,N_24272,N_24933);
and U27594 (N_27594,N_26824,N_26210);
xor U27595 (N_27595,N_25806,N_24280);
nor U27596 (N_27596,N_25965,N_25136);
or U27597 (N_27597,N_25486,N_26987);
or U27598 (N_27598,N_26642,N_25696);
or U27599 (N_27599,N_25034,N_25575);
and U27600 (N_27600,N_25308,N_26781);
or U27601 (N_27601,N_26247,N_24443);
or U27602 (N_27602,N_26652,N_26830);
and U27603 (N_27603,N_24180,N_24617);
or U27604 (N_27604,N_24521,N_25673);
nand U27605 (N_27605,N_24483,N_24986);
nand U27606 (N_27606,N_26428,N_26129);
nand U27607 (N_27607,N_26590,N_26742);
or U27608 (N_27608,N_26795,N_24008);
nand U27609 (N_27609,N_25758,N_24833);
and U27610 (N_27610,N_26673,N_25442);
nor U27611 (N_27611,N_24528,N_25826);
nand U27612 (N_27612,N_26894,N_24978);
or U27613 (N_27613,N_24636,N_26122);
or U27614 (N_27614,N_24586,N_24233);
xor U27615 (N_27615,N_24375,N_25732);
nand U27616 (N_27616,N_25119,N_24829);
nor U27617 (N_27617,N_24717,N_26327);
nand U27618 (N_27618,N_26687,N_26442);
nand U27619 (N_27619,N_26026,N_24552);
nand U27620 (N_27620,N_25804,N_24876);
nor U27621 (N_27621,N_26528,N_25737);
or U27622 (N_27622,N_25088,N_25300);
or U27623 (N_27623,N_24741,N_24739);
nand U27624 (N_27624,N_26382,N_26948);
nand U27625 (N_27625,N_25945,N_25848);
nor U27626 (N_27626,N_24927,N_25052);
nand U27627 (N_27627,N_25882,N_26881);
nand U27628 (N_27628,N_24730,N_24831);
nand U27629 (N_27629,N_26464,N_24716);
or U27630 (N_27630,N_25246,N_25313);
and U27631 (N_27631,N_24924,N_24253);
and U27632 (N_27632,N_26062,N_24580);
nor U27633 (N_27633,N_26861,N_24852);
xor U27634 (N_27634,N_25428,N_25670);
xor U27635 (N_27635,N_24915,N_26194);
nor U27636 (N_27636,N_25761,N_25341);
xor U27637 (N_27637,N_25852,N_26380);
and U27638 (N_27638,N_26367,N_25279);
nor U27639 (N_27639,N_24002,N_25751);
nand U27640 (N_27640,N_24067,N_25786);
or U27641 (N_27641,N_24453,N_26346);
and U27642 (N_27642,N_26321,N_24240);
nand U27643 (N_27643,N_26402,N_24755);
and U27644 (N_27644,N_24864,N_26738);
and U27645 (N_27645,N_25877,N_25631);
xor U27646 (N_27646,N_25700,N_26038);
xnor U27647 (N_27647,N_24602,N_26157);
nor U27648 (N_27648,N_25710,N_26081);
nor U27649 (N_27649,N_26720,N_24074);
and U27650 (N_27650,N_26924,N_25966);
or U27651 (N_27651,N_26435,N_24574);
xor U27652 (N_27652,N_25112,N_24258);
xor U27653 (N_27653,N_25974,N_25868);
nor U27654 (N_27654,N_25552,N_25912);
and U27655 (N_27655,N_25419,N_25068);
and U27656 (N_27656,N_26695,N_26604);
nand U27657 (N_27657,N_26466,N_25433);
and U27658 (N_27658,N_25601,N_26536);
nand U27659 (N_27659,N_24119,N_25387);
nor U27660 (N_27660,N_24825,N_25203);
and U27661 (N_27661,N_25148,N_24989);
nor U27662 (N_27662,N_26483,N_25749);
nand U27663 (N_27663,N_26496,N_24249);
xor U27664 (N_27664,N_25644,N_24896);
and U27665 (N_27665,N_24200,N_24030);
nand U27666 (N_27666,N_25403,N_26562);
nor U27667 (N_27667,N_24913,N_24594);
nor U27668 (N_27668,N_24001,N_26580);
nand U27669 (N_27669,N_24211,N_24722);
xnor U27670 (N_27670,N_25334,N_25267);
and U27671 (N_27671,N_24393,N_25168);
and U27672 (N_27672,N_26140,N_26233);
xor U27673 (N_27673,N_25327,N_25132);
or U27674 (N_27674,N_24439,N_26048);
nor U27675 (N_27675,N_24588,N_24326);
and U27676 (N_27676,N_25899,N_24535);
or U27677 (N_27677,N_26332,N_26163);
or U27678 (N_27678,N_26759,N_25006);
xor U27679 (N_27679,N_24692,N_25976);
nand U27680 (N_27680,N_26262,N_24327);
xor U27681 (N_27681,N_26427,N_24952);
xor U27682 (N_27682,N_25459,N_25014);
xnor U27683 (N_27683,N_25640,N_25093);
nand U27684 (N_27684,N_25664,N_24445);
nand U27685 (N_27685,N_26059,N_25711);
nand U27686 (N_27686,N_24633,N_26390);
nand U27687 (N_27687,N_26792,N_25057);
xnor U27688 (N_27688,N_24163,N_24773);
nor U27689 (N_27689,N_26929,N_24685);
and U27690 (N_27690,N_25667,N_25605);
nor U27691 (N_27691,N_26519,N_24764);
or U27692 (N_27692,N_24859,N_25252);
and U27693 (N_27693,N_24775,N_24804);
or U27694 (N_27694,N_24648,N_25717);
and U27695 (N_27695,N_26815,N_25643);
and U27696 (N_27696,N_26974,N_26045);
nor U27697 (N_27697,N_24091,N_26486);
xnor U27698 (N_27698,N_26620,N_24276);
and U27699 (N_27699,N_26413,N_26315);
and U27700 (N_27700,N_25409,N_25046);
xor U27701 (N_27701,N_24363,N_25462);
and U27702 (N_27702,N_25924,N_24099);
nand U27703 (N_27703,N_26407,N_26012);
xor U27704 (N_27704,N_26328,N_26144);
or U27705 (N_27705,N_26653,N_25890);
xnor U27706 (N_27706,N_26893,N_26230);
or U27707 (N_27707,N_24718,N_24577);
or U27708 (N_27708,N_24625,N_24098);
nand U27709 (N_27709,N_25477,N_26069);
or U27710 (N_27710,N_24410,N_24772);
or U27711 (N_27711,N_26773,N_24157);
or U27712 (N_27712,N_25998,N_25412);
xor U27713 (N_27713,N_25558,N_26717);
nor U27714 (N_27714,N_24298,N_24055);
xnor U27715 (N_27715,N_25866,N_24895);
and U27716 (N_27716,N_26499,N_24855);
or U27717 (N_27717,N_24899,N_24663);
nor U27718 (N_27718,N_24643,N_24970);
or U27719 (N_27719,N_24014,N_25183);
nor U27720 (N_27720,N_24808,N_26051);
nand U27721 (N_27721,N_26847,N_24405);
nand U27722 (N_27722,N_25531,N_25138);
xor U27723 (N_27723,N_26297,N_26760);
or U27724 (N_27724,N_26222,N_24649);
xor U27725 (N_27725,N_26450,N_25031);
xor U27726 (N_27726,N_26872,N_24826);
nand U27727 (N_27727,N_26616,N_24237);
nand U27728 (N_27728,N_25196,N_25415);
or U27729 (N_27729,N_24171,N_25481);
nor U27730 (N_27730,N_24800,N_25733);
nor U27731 (N_27731,N_25476,N_24005);
xnor U27732 (N_27732,N_25980,N_24946);
nor U27733 (N_27733,N_25591,N_24132);
nor U27734 (N_27734,N_24505,N_26714);
nor U27735 (N_27735,N_26818,N_25058);
nand U27736 (N_27736,N_26433,N_26023);
nor U27737 (N_27737,N_25045,N_25274);
and U27738 (N_27738,N_25215,N_24027);
or U27739 (N_27739,N_24162,N_26169);
xnor U27740 (N_27740,N_26675,N_24319);
nand U27741 (N_27741,N_26836,N_25833);
or U27742 (N_27742,N_26672,N_25150);
or U27743 (N_27743,N_24411,N_26822);
nand U27744 (N_27744,N_25470,N_25579);
nor U27745 (N_27745,N_25364,N_26599);
or U27746 (N_27746,N_26826,N_26935);
nor U27747 (N_27747,N_25951,N_24397);
xnor U27748 (N_27748,N_26096,N_24083);
xor U27749 (N_27749,N_25109,N_25714);
and U27750 (N_27750,N_26707,N_25467);
or U27751 (N_27751,N_24097,N_26730);
nand U27752 (N_27752,N_24121,N_24359);
and U27753 (N_27753,N_24514,N_24866);
or U27754 (N_27754,N_26565,N_24500);
xnor U27755 (N_27755,N_26954,N_26655);
and U27756 (N_27756,N_26275,N_25378);
nand U27757 (N_27757,N_26637,N_26922);
nor U27758 (N_27758,N_25410,N_26882);
and U27759 (N_27759,N_26014,N_25604);
and U27760 (N_27760,N_25471,N_25336);
nor U27761 (N_27761,N_25108,N_25139);
and U27762 (N_27762,N_24776,N_26509);
xor U27763 (N_27763,N_25637,N_25615);
nand U27764 (N_27764,N_26141,N_24848);
and U27765 (N_27765,N_24841,N_25538);
xor U27766 (N_27766,N_25595,N_26596);
and U27767 (N_27767,N_26986,N_25214);
nor U27768 (N_27768,N_24700,N_26808);
nand U27769 (N_27769,N_24212,N_26353);
and U27770 (N_27770,N_26408,N_24987);
and U27771 (N_27771,N_26985,N_24734);
or U27772 (N_27772,N_25551,N_26677);
nor U27773 (N_27773,N_24760,N_25897);
and U27774 (N_27774,N_25843,N_24209);
and U27775 (N_27775,N_24546,N_25830);
nand U27776 (N_27776,N_25247,N_26866);
and U27777 (N_27777,N_26783,N_24285);
nand U27778 (N_27778,N_25060,N_25666);
nand U27779 (N_27779,N_24160,N_24571);
nor U27780 (N_27780,N_26309,N_24053);
nor U27781 (N_27781,N_24705,N_24757);
xnor U27782 (N_27782,N_26654,N_26360);
nand U27783 (N_27783,N_24023,N_25748);
xnor U27784 (N_27784,N_26516,N_26185);
xor U27785 (N_27785,N_26118,N_25612);
and U27786 (N_27786,N_24274,N_25581);
or U27787 (N_27787,N_26476,N_24447);
and U27788 (N_27788,N_24519,N_25893);
nand U27789 (N_27789,N_25634,N_26029);
or U27790 (N_27790,N_24340,N_26090);
nand U27791 (N_27791,N_25788,N_24908);
and U27792 (N_27792,N_25369,N_26632);
or U27793 (N_27793,N_25067,N_25394);
or U27794 (N_27794,N_25147,N_25430);
xnor U27795 (N_27795,N_24290,N_25626);
nor U27796 (N_27796,N_26676,N_24603);
nor U27797 (N_27797,N_26437,N_26615);
nand U27798 (N_27798,N_24995,N_26825);
nand U27799 (N_27799,N_24676,N_25162);
nand U27800 (N_27800,N_24017,N_24501);
nand U27801 (N_27801,N_25972,N_25324);
nand U27802 (N_27802,N_24809,N_25642);
xor U27803 (N_27803,N_26878,N_26844);
xnor U27804 (N_27804,N_26148,N_25461);
and U27805 (N_27805,N_24173,N_24303);
or U27806 (N_27806,N_24154,N_26158);
nor U27807 (N_27807,N_26025,N_25831);
nor U27808 (N_27808,N_25450,N_26271);
or U27809 (N_27809,N_24638,N_25937);
and U27810 (N_27810,N_26221,N_26816);
nand U27811 (N_27811,N_25326,N_26534);
and U27812 (N_27812,N_25163,N_24151);
xor U27813 (N_27813,N_24869,N_26627);
xor U27814 (N_27814,N_24199,N_25533);
or U27815 (N_27815,N_26906,N_24283);
nand U27816 (N_27816,N_25516,N_24495);
and U27817 (N_27817,N_26207,N_25469);
or U27818 (N_27818,N_26043,N_26356);
nand U27819 (N_27819,N_25766,N_25229);
nor U27820 (N_27820,N_26823,N_25548);
or U27821 (N_27821,N_25534,N_24682);
and U27822 (N_27822,N_25589,N_26421);
xor U27823 (N_27823,N_26603,N_25655);
or U27824 (N_27824,N_24845,N_26898);
and U27825 (N_27825,N_24246,N_24389);
xor U27826 (N_27826,N_25730,N_26495);
or U27827 (N_27827,N_26282,N_26261);
nor U27828 (N_27828,N_24377,N_25935);
xor U27829 (N_27829,N_26459,N_25097);
and U27830 (N_27830,N_25383,N_24819);
and U27831 (N_27831,N_25862,N_26988);
xnor U27832 (N_27832,N_25472,N_24763);
nor U27833 (N_27833,N_25807,N_26875);
or U27834 (N_27834,N_25602,N_26946);
and U27835 (N_27835,N_24923,N_26415);
and U27836 (N_27836,N_24893,N_26191);
xor U27837 (N_27837,N_25297,N_25985);
and U27838 (N_27838,N_26647,N_24307);
nor U27839 (N_27839,N_24006,N_24286);
or U27840 (N_27840,N_24583,N_26009);
xnor U27841 (N_27841,N_25738,N_26621);
nand U27842 (N_27842,N_25702,N_25898);
xor U27843 (N_27843,N_24983,N_26333);
nand U27844 (N_27844,N_25881,N_24185);
nor U27845 (N_27845,N_26635,N_24131);
xnor U27846 (N_27846,N_25854,N_25562);
or U27847 (N_27847,N_24865,N_26704);
or U27848 (N_27848,N_26771,N_25850);
nor U27849 (N_27849,N_24401,N_26628);
and U27850 (N_27850,N_25199,N_26003);
nand U27851 (N_27851,N_25226,N_24744);
xnor U27852 (N_27852,N_25090,N_26213);
or U27853 (N_27853,N_24799,N_24547);
and U27854 (N_27854,N_25012,N_26276);
nand U27855 (N_27855,N_26965,N_24778);
and U27856 (N_27856,N_25154,N_25434);
nand U27857 (N_27857,N_24582,N_26457);
nor U27858 (N_27858,N_25120,N_24170);
and U27859 (N_27859,N_26775,N_26205);
nand U27860 (N_27860,N_26709,N_25194);
nand U27861 (N_27861,N_24905,N_26307);
nand U27862 (N_27862,N_25029,N_26713);
or U27863 (N_27863,N_24677,N_26810);
nor U27864 (N_27864,N_25076,N_25938);
xnor U27865 (N_27865,N_26242,N_24466);
nand U27866 (N_27866,N_26497,N_24696);
nor U27867 (N_27867,N_26254,N_26477);
xnor U27868 (N_27868,N_24215,N_24853);
xor U27869 (N_27869,N_25347,N_25483);
nor U27870 (N_27870,N_26349,N_25314);
nor U27871 (N_27871,N_24208,N_25523);
or U27872 (N_27872,N_26145,N_24497);
or U27873 (N_27873,N_24542,N_24228);
nor U27874 (N_27874,N_26780,N_26204);
nand U27875 (N_27875,N_25500,N_25559);
nand U27876 (N_27876,N_25173,N_24186);
nand U27877 (N_27877,N_24928,N_26080);
nor U27878 (N_27878,N_24078,N_24567);
or U27879 (N_27879,N_25907,N_25669);
nor U27880 (N_27880,N_25357,N_25569);
xnor U27881 (N_27881,N_26002,N_24968);
nand U27882 (N_27882,N_25041,N_26820);
nand U27883 (N_27883,N_26947,N_24260);
nand U27884 (N_27884,N_26557,N_25895);
xor U27885 (N_27885,N_25009,N_24991);
xnor U27886 (N_27886,N_25978,N_26828);
nor U27887 (N_27887,N_24544,N_24281);
nand U27888 (N_27888,N_24216,N_26969);
and U27889 (N_27889,N_24033,N_25835);
or U27890 (N_27890,N_24457,N_24333);
or U27891 (N_27891,N_25023,N_25005);
and U27892 (N_27892,N_26173,N_26429);
and U27893 (N_27893,N_25239,N_24444);
or U27894 (N_27894,N_25674,N_24641);
xnor U27895 (N_27895,N_25146,N_25796);
and U27896 (N_27896,N_26351,N_24113);
nor U27897 (N_27897,N_25152,N_25197);
or U27898 (N_27898,N_24314,N_24737);
nand U27899 (N_27899,N_26799,N_24684);
and U27900 (N_27900,N_25380,N_25013);
or U27901 (N_27901,N_26318,N_26053);
and U27902 (N_27902,N_25456,N_24683);
or U27903 (N_27903,N_25892,N_26506);
xnor U27904 (N_27904,N_25130,N_25553);
nor U27905 (N_27905,N_24781,N_24077);
or U27906 (N_27906,N_24693,N_26022);
xor U27907 (N_27907,N_24660,N_25561);
xnor U27908 (N_27908,N_25743,N_25846);
and U27909 (N_27909,N_25752,N_25282);
or U27910 (N_27910,N_25724,N_26034);
nor U27911 (N_27911,N_24471,N_25995);
nor U27912 (N_27912,N_24720,N_25815);
nor U27913 (N_27913,N_25521,N_24916);
and U27914 (N_27914,N_24305,N_24623);
and U27915 (N_27915,N_25106,N_25281);
nand U27916 (N_27916,N_24198,N_25231);
or U27917 (N_27917,N_24047,N_24048);
xor U27918 (N_27918,N_26348,N_24032);
nor U27919 (N_27919,N_25544,N_26629);
and U27920 (N_27920,N_24284,N_24089);
nand U27921 (N_27921,N_24308,N_24135);
nor U27922 (N_27922,N_26804,N_24316);
xnor U27923 (N_27923,N_24672,N_26011);
xor U27924 (N_27924,N_25362,N_25514);
or U27925 (N_27925,N_24358,N_25224);
and U27926 (N_27926,N_26541,N_24210);
and U27927 (N_27927,N_24644,N_25401);
nor U27928 (N_27928,N_26099,N_24486);
nor U27929 (N_27929,N_24918,N_25798);
and U27930 (N_27930,N_26040,N_26406);
or U27931 (N_27931,N_26229,N_26517);
xor U27932 (N_27932,N_26434,N_24084);
nand U27933 (N_27933,N_26245,N_24620);
nor U27934 (N_27934,N_26937,N_25290);
and U27935 (N_27935,N_26700,N_26324);
and U27936 (N_27936,N_25947,N_25734);
nand U27937 (N_27937,N_26649,N_25526);
xnor U27938 (N_27938,N_25159,N_25082);
nand U27939 (N_27939,N_25825,N_25723);
or U27940 (N_27940,N_24768,N_26503);
nand U27941 (N_27941,N_26094,N_26997);
nand U27942 (N_27942,N_26681,N_25791);
and U27943 (N_27943,N_24127,N_25703);
nand U27944 (N_27944,N_26358,N_25641);
and U27945 (N_27945,N_26368,N_26283);
or U27946 (N_27946,N_25348,N_25145);
xnor U27947 (N_27947,N_25769,N_26066);
nor U27948 (N_27948,N_24742,N_26923);
nand U27949 (N_27949,N_25056,N_24894);
xnor U27950 (N_27950,N_24381,N_24277);
and U27951 (N_27951,N_24993,N_24066);
nor U27952 (N_27952,N_24612,N_24732);
nor U27953 (N_27953,N_26161,N_26761);
nor U27954 (N_27954,N_25560,N_24409);
and U27955 (N_27955,N_25134,N_24224);
or U27956 (N_27956,N_25156,N_24165);
nand U27957 (N_27957,N_25725,N_24007);
xnor U27958 (N_27958,N_25272,N_26606);
or U27959 (N_27959,N_25195,N_25679);
nor U27960 (N_27960,N_26341,N_26806);
xor U27961 (N_27961,N_25616,N_24839);
and U27962 (N_27962,N_25283,N_26196);
nor U27963 (N_27963,N_24133,N_24172);
nand U27964 (N_27964,N_26774,N_25709);
nor U27965 (N_27965,N_24416,N_24656);
xnor U27966 (N_27966,N_25957,N_24120);
nand U27967 (N_27967,N_26711,N_25571);
xor U27968 (N_27968,N_24830,N_24596);
and U27969 (N_27969,N_24556,N_26082);
nor U27970 (N_27970,N_25261,N_25365);
or U27971 (N_27971,N_25914,N_26728);
nand U27972 (N_27972,N_24892,N_25675);
nor U27973 (N_27973,N_26447,N_24291);
nor U27974 (N_27974,N_24106,N_26240);
or U27975 (N_27975,N_26648,N_24543);
or U27976 (N_27976,N_25555,N_24382);
nand U27977 (N_27977,N_24335,N_25155);
or U27978 (N_27978,N_25744,N_26618);
nand U27979 (N_27979,N_26873,N_25904);
or U27980 (N_27980,N_24331,N_25244);
nor U27981 (N_27981,N_25623,N_26779);
xor U27982 (N_27982,N_24545,N_24783);
xor U27983 (N_27983,N_24191,N_25351);
and U27984 (N_27984,N_24912,N_25495);
nor U27985 (N_27985,N_25124,N_26727);
xor U27986 (N_27986,N_26871,N_26805);
or U27987 (N_27987,N_26132,N_24858);
nand U27988 (N_27988,N_24437,N_24138);
nand U27989 (N_27989,N_26743,N_26514);
or U27990 (N_27990,N_25936,N_25886);
xnor U27991 (N_27991,N_24356,N_26863);
nand U27992 (N_27992,N_24697,N_26054);
nor U27993 (N_27993,N_25652,N_25762);
nor U27994 (N_27994,N_26152,N_26747);
nand U27995 (N_27995,N_26238,N_24454);
or U27996 (N_27996,N_26814,N_24955);
or U27997 (N_27997,N_26605,N_26890);
nor U27998 (N_27998,N_25025,N_25532);
xor U27999 (N_27999,N_26813,N_24903);
nor U28000 (N_28000,N_26626,N_24275);
and U28001 (N_28001,N_26263,N_25350);
nand U28002 (N_28002,N_24964,N_26174);
xor U28003 (N_28003,N_25243,N_24009);
nor U28004 (N_28004,N_25258,N_24537);
nor U28005 (N_28005,N_26570,N_24161);
nor U28006 (N_28006,N_25694,N_26266);
or U28007 (N_28007,N_26412,N_25010);
or U28008 (N_28008,N_24203,N_26120);
nand U28009 (N_28009,N_24811,N_25126);
nor U28010 (N_28010,N_25537,N_25746);
xnor U28011 (N_28011,N_24464,N_26914);
xnor U28012 (N_28012,N_24652,N_26166);
nor U28013 (N_28013,N_25929,N_25547);
xor U28014 (N_28014,N_24522,N_26253);
xor U28015 (N_28015,N_26325,N_25956);
or U28016 (N_28016,N_24626,N_24675);
and U28017 (N_28017,N_24785,N_26493);
xor U28018 (N_28018,N_24635,N_25672);
and U28019 (N_28019,N_24517,N_24572);
or U28020 (N_28020,N_26721,N_26019);
xor U28021 (N_28021,N_24266,N_24921);
xnor U28022 (N_28022,N_25549,N_25686);
nand U28023 (N_28023,N_25390,N_25095);
nor U28024 (N_28024,N_26581,N_24891);
nor U28025 (N_28025,N_26839,N_25582);
nand U28026 (N_28026,N_25418,N_25318);
and U28027 (N_28027,N_26179,N_26208);
nor U28028 (N_28028,N_26735,N_26488);
nor U28029 (N_28029,N_26378,N_25844);
or U28030 (N_28030,N_24071,N_25954);
xnor U28031 (N_28031,N_26105,N_26928);
xnor U28032 (N_28032,N_24306,N_24530);
and U28033 (N_28033,N_24802,N_26504);
and U28034 (N_28034,N_26219,N_26867);
and U28035 (N_28035,N_26362,N_26949);
and U28036 (N_28036,N_24386,N_25828);
and U28037 (N_28037,N_26231,N_24520);
xor U28038 (N_28038,N_25241,N_24557);
xnor U28039 (N_28039,N_26572,N_26338);
or U28040 (N_28040,N_24645,N_24836);
xnor U28041 (N_28041,N_25853,N_26361);
xor U28042 (N_28042,N_26573,N_26088);
nand U28043 (N_28043,N_26150,N_25719);
xnor U28044 (N_28044,N_26334,N_25343);
and U28045 (N_28045,N_24713,N_25969);
or U28046 (N_28046,N_24904,N_26884);
xor U28047 (N_28047,N_25458,N_24981);
or U28048 (N_28048,N_26232,N_24013);
nor U28049 (N_28049,N_25879,N_26733);
and U28050 (N_28050,N_24703,N_25255);
nor U28051 (N_28051,N_26785,N_26311);
nor U28052 (N_28052,N_24054,N_25541);
or U28053 (N_28053,N_24631,N_25574);
and U28054 (N_28054,N_24523,N_25989);
nor U28055 (N_28055,N_24728,N_24434);
and U28056 (N_28056,N_24949,N_24780);
nand U28057 (N_28057,N_26007,N_26308);
xnor U28058 (N_28058,N_24834,N_24479);
and U28059 (N_28059,N_25578,N_26788);
or U28060 (N_28060,N_24080,N_26874);
nor U28061 (N_28061,N_25811,N_25987);
nor U28062 (N_28062,N_24313,N_26100);
nand U28063 (N_28063,N_24605,N_25151);
and U28064 (N_28064,N_24844,N_25959);
nor U28065 (N_28065,N_24566,N_25373);
nand U28066 (N_28066,N_25098,N_24300);
xor U28067 (N_28067,N_26691,N_25979);
xor U28068 (N_28068,N_24205,N_24753);
xnor U28069 (N_28069,N_25035,N_25859);
and U28070 (N_28070,N_26329,N_26469);
nor U28071 (N_28071,N_25361,N_26149);
or U28072 (N_28072,N_25906,N_24037);
nand U28073 (N_28073,N_24143,N_26198);
nor U28074 (N_28074,N_25232,N_25078);
xnor U28075 (N_28075,N_24821,N_25805);
xor U28076 (N_28076,N_26128,N_24140);
nor U28077 (N_28077,N_26417,N_24997);
xnor U28078 (N_28078,N_24123,N_24507);
nand U28079 (N_28079,N_26373,N_25463);
nor U28080 (N_28080,N_26845,N_25123);
xnor U28081 (N_28081,N_25948,N_26164);
nor U28082 (N_28082,N_24451,N_25809);
nor U28083 (N_28083,N_25913,N_25186);
nor U28084 (N_28084,N_25417,N_24670);
or U28085 (N_28085,N_26461,N_24111);
xnor U28086 (N_28086,N_24666,N_26425);
nor U28087 (N_28087,N_25902,N_24310);
nor U28088 (N_28088,N_24339,N_24559);
nor U28089 (N_28089,N_26319,N_24691);
or U28090 (N_28090,N_26723,N_26624);
xnor U28091 (N_28091,N_24661,N_26520);
or U28092 (N_28092,N_24217,N_24640);
or U28093 (N_28093,N_26473,N_25736);
nor U28094 (N_28094,N_25011,N_25386);
nand U28095 (N_28095,N_25584,N_24525);
xor U28096 (N_28096,N_26489,N_24529);
or U28097 (N_28097,N_25529,N_26577);
xnor U28098 (N_28098,N_24950,N_24372);
nand U28099 (N_28099,N_26798,N_24884);
xnor U28100 (N_28100,N_24167,N_25920);
or U28101 (N_28101,N_24817,N_25598);
and U28102 (N_28102,N_25834,N_24729);
xor U28103 (N_28103,N_25923,N_26998);
nand U28104 (N_28104,N_26999,N_25763);
or U28105 (N_28105,N_26908,N_25795);
or U28106 (N_28106,N_25275,N_25397);
nand U28107 (N_28107,N_25727,N_24767);
xor U28108 (N_28108,N_26139,N_25212);
or U28109 (N_28109,N_24890,N_25593);
or U28110 (N_28110,N_26225,N_24373);
nor U28111 (N_28111,N_26609,N_24399);
nor U28112 (N_28112,N_26712,N_26951);
and U28113 (N_28113,N_24791,N_25081);
or U28114 (N_28114,N_24782,N_24092);
nand U28115 (N_28115,N_26000,N_25307);
and U28116 (N_28116,N_25117,N_25375);
or U28117 (N_28117,N_24035,N_26991);
or U28118 (N_28118,N_24681,N_25742);
and U28119 (N_28119,N_25311,N_24086);
nor U28120 (N_28120,N_25718,N_24046);
nor U28121 (N_28121,N_25797,N_25254);
xor U28122 (N_28122,N_24657,N_25933);
xnor U28123 (N_28123,N_25265,N_26561);
and U28124 (N_28124,N_26278,N_26880);
nor U28125 (N_28125,N_24736,N_24878);
xnor U28126 (N_28126,N_26856,N_25501);
or U28127 (N_28127,N_24822,N_26696);
nor U28128 (N_28128,N_24996,N_25299);
nand U28129 (N_28129,N_25785,N_25287);
or U28130 (N_28130,N_24597,N_24658);
and U28131 (N_28131,N_24735,N_26274);
or U28132 (N_28132,N_25096,N_24236);
nor U28133 (N_28133,N_25646,N_26767);
or U28134 (N_28134,N_26201,N_26990);
or U28135 (N_28135,N_26716,N_25298);
xnor U28136 (N_28136,N_26172,N_26689);
xnor U28137 (N_28137,N_25794,N_24034);
nor U28138 (N_28138,N_25847,N_25505);
and U28139 (N_28139,N_26919,N_24932);
xnor U28140 (N_28140,N_26651,N_24481);
or U28141 (N_28141,N_25996,N_26701);
or U28142 (N_28142,N_25074,N_24070);
nor U28143 (N_28143,N_26967,N_26162);
and U28144 (N_28144,N_26098,N_26392);
nor U28145 (N_28145,N_26156,N_24406);
nor U28146 (N_28146,N_26827,N_26865);
and U28147 (N_28147,N_24973,N_24465);
nor U28148 (N_28148,N_25121,N_25286);
nand U28149 (N_28149,N_25810,N_26718);
and U28150 (N_28150,N_25288,N_24828);
nor U28151 (N_28151,N_26745,N_24304);
nand U28152 (N_28152,N_26722,N_26363);
xor U28153 (N_28153,N_25003,N_24516);
nor U28154 (N_28154,N_26422,N_25802);
nand U28155 (N_28155,N_25405,N_24309);
nand U28156 (N_28156,N_25465,N_26035);
nor U28157 (N_28157,N_24321,N_26223);
or U28158 (N_28158,N_24440,N_25681);
nand U28159 (N_28159,N_25051,N_25115);
and U28160 (N_28160,N_24056,N_26178);
xor U28161 (N_28161,N_24659,N_24554);
xor U28162 (N_28162,N_26226,N_26834);
nand U28163 (N_28163,N_24118,N_26979);
xnor U28164 (N_28164,N_26682,N_24328);
nand U28165 (N_28165,N_25172,N_26644);
xor U28166 (N_28166,N_26119,N_24985);
nand U28167 (N_28167,N_26267,N_24914);
nor U28168 (N_28168,N_24148,N_26764);
xnor U28169 (N_28169,N_24042,N_26671);
nor U28170 (N_28170,N_24706,N_26008);
and U28171 (N_28171,N_24929,N_24475);
and U28172 (N_28172,N_26510,N_25799);
and U28173 (N_28173,N_25264,N_25808);
nand U28174 (N_28174,N_24886,N_24551);
and U28175 (N_28175,N_24242,N_25659);
nand U28176 (N_28176,N_25542,N_26803);
nor U28177 (N_28177,N_25609,N_24220);
xor U28178 (N_28178,N_25783,N_24630);
nand U28179 (N_28179,N_24611,N_24278);
nor U28180 (N_28180,N_26097,N_25131);
nand U28181 (N_28181,N_26317,N_24296);
or U28182 (N_28182,N_25726,N_24245);
nand U28183 (N_28183,N_24868,N_25018);
nor U28184 (N_28184,N_26335,N_24352);
nand U28185 (N_28185,N_24183,N_25891);
nor U28186 (N_28186,N_26559,N_26848);
nor U28187 (N_28187,N_24016,N_25339);
nor U28188 (N_28188,N_26015,N_24962);
nor U28189 (N_28189,N_25566,N_24490);
or U28190 (N_28190,N_25017,N_26387);
or U28191 (N_28191,N_25024,N_26945);
nor U28192 (N_28192,N_24223,N_24175);
nor U28193 (N_28193,N_24227,N_25665);
xnor U28194 (N_28194,N_25856,N_24204);
and U28195 (N_28195,N_24686,N_24000);
and U28196 (N_28196,N_25449,N_26249);
xnor U28197 (N_28197,N_24613,N_24606);
and U28198 (N_28198,N_26971,N_25925);
and U28199 (N_28199,N_26265,N_25864);
nand U28200 (N_28200,N_24289,N_25371);
nand U28201 (N_28201,N_26183,N_24400);
nand U28202 (N_28202,N_25210,N_26513);
or U28203 (N_28203,N_24072,N_25630);
nand U28204 (N_28204,N_26279,N_26708);
and U28205 (N_28205,N_26970,N_26020);
and U28206 (N_28206,N_26239,N_26512);
or U28207 (N_28207,N_25376,N_25653);
xnor U28208 (N_28208,N_26484,N_24049);
nor U28209 (N_28209,N_26052,N_26560);
nand U28210 (N_28210,N_25894,N_26746);
or U28211 (N_28211,N_24980,N_24179);
and U28212 (N_28212,N_26032,N_26111);
xnor U28213 (N_28213,N_26715,N_24214);
or U28214 (N_28214,N_25392,N_25943);
nor U28215 (N_28215,N_25781,N_26916);
nor U28216 (N_28216,N_26411,N_25493);
and U28217 (N_28217,N_25556,N_26113);
and U28218 (N_28218,N_25302,N_25102);
nor U28219 (N_28219,N_26550,N_24232);
and U28220 (N_28220,N_24604,N_25973);
and U28221 (N_28221,N_26787,N_25982);
and U28222 (N_28222,N_25803,N_25722);
and U28223 (N_28223,N_25999,N_25027);
and U28224 (N_28224,N_25627,N_26036);
nor U28225 (N_28225,N_25354,N_26896);
xnor U28226 (N_28226,N_26006,N_26964);
nor U28227 (N_28227,N_24575,N_26838);
xnor U28228 (N_28228,N_26772,N_25570);
xor U28229 (N_28229,N_25284,N_24765);
xnor U28230 (N_28230,N_26901,N_24207);
xor U28231 (N_28231,N_25874,N_25233);
or U28232 (N_28232,N_24463,N_25554);
nand U28233 (N_28233,N_24920,N_25331);
nand U28234 (N_28234,N_26288,N_25837);
nor U28235 (N_28235,N_26877,N_24591);
nand U28236 (N_28236,N_26465,N_25446);
or U28237 (N_28237,N_24122,N_24473);
and U28238 (N_28238,N_26608,N_26364);
and U28239 (N_28239,N_26280,N_24061);
nand U28240 (N_28240,N_25157,N_26010);
nor U28241 (N_28241,N_24550,N_26614);
and U28242 (N_28242,N_24761,N_25485);
xor U28243 (N_28243,N_26273,N_26789);
or U28244 (N_28244,N_26284,N_25278);
xor U28245 (N_28245,N_25639,N_24241);
nand U28246 (N_28246,N_25820,N_26891);
xnor U28247 (N_28247,N_25206,N_25448);
and U28248 (N_28248,N_26538,N_24446);
or U28249 (N_28249,N_25105,N_24065);
and U28250 (N_28250,N_24838,N_24404);
nor U28251 (N_28251,N_24019,N_26071);
xnor U28252 (N_28252,N_25629,N_26670);
nor U28253 (N_28253,N_26909,N_25330);
and U28254 (N_28254,N_24595,N_26613);
nand U28255 (N_28255,N_26444,N_25408);
or U28256 (N_28256,N_25517,N_25038);
or U28257 (N_28257,N_26960,N_26533);
xnor U28258 (N_28258,N_26272,N_24794);
nand U28259 (N_28259,N_24850,N_26074);
xnor U28260 (N_28260,N_26236,N_26740);
xnor U28261 (N_28261,N_24312,N_24922);
xnor U28262 (N_28262,N_25905,N_25209);
or U28263 (N_28263,N_24721,N_26851);
or U28264 (N_28264,N_25201,N_24664);
xor U28265 (N_28265,N_25819,N_26491);
nand U28266 (N_28266,N_26912,N_24503);
and U28267 (N_28267,N_25872,N_25200);
xor U28268 (N_28268,N_24587,N_24745);
and U28269 (N_28269,N_25880,N_25638);
nand U28270 (N_28270,N_25143,N_25647);
xnor U28271 (N_28271,N_26257,N_26312);
and U28272 (N_28272,N_25524,N_24436);
nand U28273 (N_28273,N_24708,N_26633);
xor U28274 (N_28274,N_25188,N_25860);
or U28275 (N_28275,N_26189,N_24756);
xnor U28276 (N_28276,N_26165,N_26756);
xnor U28277 (N_28277,N_26314,N_25910);
or U28278 (N_28278,N_26786,N_24798);
or U28279 (N_28279,N_25981,N_25824);
nand U28280 (N_28280,N_25713,N_25821);
nor U28281 (N_28281,N_25069,N_26268);
nand U28282 (N_28282,N_24264,N_25260);
or U28283 (N_28283,N_26535,N_25444);
xnor U28284 (N_28284,N_26595,N_26123);
and U28285 (N_28285,N_25360,N_26587);
nor U28286 (N_28286,N_24941,N_25939);
nor U28287 (N_28287,N_24712,N_26686);
nor U28288 (N_28288,N_26791,N_26555);
or U28289 (N_28289,N_26114,N_24627);
and U28290 (N_28290,N_26719,N_25125);
nor U28291 (N_28291,N_25849,N_25294);
or U28292 (N_28292,N_26216,N_25236);
or U28293 (N_28293,N_26544,N_24412);
and U28294 (N_28294,N_26617,N_25518);
or U28295 (N_28295,N_26109,N_26212);
and U28296 (N_28296,N_26917,N_24239);
xnor U28297 (N_28297,N_26115,N_25827);
and U28298 (N_28298,N_24549,N_24539);
and U28299 (N_28299,N_26936,N_24164);
xnor U28300 (N_28300,N_25193,N_25167);
and U28301 (N_28301,N_26110,N_26638);
and U28302 (N_28302,N_25829,N_24302);
and U28303 (N_28303,N_26918,N_24311);
nor U28304 (N_28304,N_25242,N_26515);
nor U28305 (N_28305,N_26540,N_25504);
nor U28306 (N_28306,N_26186,N_26460);
nor U28307 (N_28307,N_24193,N_26494);
nand U28308 (N_28308,N_26588,N_25245);
xnor U28309 (N_28309,N_24857,N_25273);
nand U28310 (N_28310,N_24293,N_25413);
xnor U28311 (N_28311,N_26302,N_26631);
and U28312 (N_28312,N_24654,N_26065);
or U28313 (N_28313,N_24085,N_24945);
nor U28314 (N_28314,N_25181,N_25075);
xor U28315 (N_28315,N_24043,N_24195);
and U28316 (N_28316,N_25608,N_25099);
and U28317 (N_28317,N_25116,N_25964);
xnor U28318 (N_28318,N_26467,N_25406);
or U28319 (N_28319,N_26108,N_24793);
nand U28320 (N_28320,N_24190,N_25946);
and U28321 (N_28321,N_26241,N_25784);
nand U28322 (N_28322,N_26549,N_26981);
and U28323 (N_28323,N_24090,N_24887);
nand U28324 (N_28324,N_25658,N_24489);
and U28325 (N_28325,N_24909,N_24769);
xor U28326 (N_28326,N_25887,N_25519);
nor U28327 (N_28327,N_26777,N_24136);
and U28328 (N_28328,N_24269,N_26751);
xnor U28329 (N_28329,N_24690,N_24942);
nor U28330 (N_28330,N_26832,N_24064);
nor U28331 (N_28331,N_25178,N_25865);
and U28332 (N_28332,N_24052,N_26674);
and U28333 (N_28333,N_24563,N_25668);
and U28334 (N_28334,N_24221,N_26992);
nor U28335 (N_28335,N_25190,N_25900);
nor U28336 (N_28336,N_24994,N_24218);
nand U28337 (N_28337,N_26441,N_25728);
nor U28338 (N_28338,N_24954,N_24075);
nor U28339 (N_28339,N_24796,N_25164);
and U28340 (N_28340,N_26962,N_24851);
and U28341 (N_28341,N_26846,N_25690);
and U28342 (N_28342,N_24608,N_24256);
nand U28343 (N_28343,N_25238,N_26095);
and U28344 (N_28344,N_26529,N_26521);
or U28345 (N_28345,N_24294,N_25374);
nor U28346 (N_28346,N_26468,N_24330);
nor U28347 (N_28347,N_26811,N_26566);
nor U28348 (N_28348,N_24907,N_24634);
xnor U28349 (N_28349,N_24689,N_26982);
nand U28350 (N_28350,N_25617,N_24350);
or U28351 (N_28351,N_26796,N_26352);
or U28352 (N_28352,N_25047,N_26192);
xor U28353 (N_28353,N_26597,N_24515);
nor U28354 (N_28354,N_25230,N_26855);
xnor U28355 (N_28355,N_26218,N_25619);
nand U28356 (N_28356,N_24081,N_25180);
nand U28357 (N_28357,N_24225,N_26103);
or U28358 (N_28358,N_26809,N_26344);
nor U28359 (N_28359,N_25352,N_26765);
and U28360 (N_28360,N_26634,N_24257);
nor U28361 (N_28361,N_25857,N_26072);
nand U28362 (N_28362,N_25065,N_26277);
and U28363 (N_28363,N_25499,N_26957);
nor U28364 (N_28364,N_24021,N_24134);
and U28365 (N_28365,N_24976,N_26849);
xor U28366 (N_28366,N_25855,N_25773);
xor U28367 (N_28367,N_26753,N_25142);
nand U28368 (N_28368,N_25248,N_26938);
and U28369 (N_28369,N_25033,N_26104);
nand U28370 (N_28370,N_24837,N_26665);
xnor U28371 (N_28371,N_24750,N_25468);
nor U28372 (N_28372,N_26037,N_26259);
or U28373 (N_28373,N_25712,N_24538);
nor U28374 (N_28374,N_24336,N_26042);
or U28375 (N_28375,N_24093,N_25662);
nor U28376 (N_28376,N_24900,N_24710);
or U28377 (N_28377,N_24063,N_26706);
xnor U28378 (N_28378,N_25332,N_25610);
xor U28379 (N_28379,N_25911,N_26860);
and U28380 (N_28380,N_24431,N_26553);
xor U28381 (N_28381,N_26821,N_26084);
nor U28382 (N_28382,N_26306,N_25228);
nand U28383 (N_28383,N_24425,N_25677);
nor U28384 (N_28384,N_24174,N_26350);
nor U28385 (N_28385,N_25368,N_24680);
nor U28386 (N_28386,N_25356,N_24901);
and U28387 (N_28387,N_25317,N_24267);
xnor U28388 (N_28388,N_26956,N_24395);
nor U28389 (N_28389,N_24367,N_24614);
or U28390 (N_28390,N_24698,N_26376);
nor U28391 (N_28391,N_24971,N_25189);
or U28392 (N_28392,N_26910,N_25932);
or U28393 (N_28393,N_26941,N_24438);
xor U28394 (N_28394,N_26505,N_25301);
or U28395 (N_28395,N_26215,N_25759);
or U28396 (N_28396,N_25509,N_25968);
nand U28397 (N_28397,N_26055,N_26106);
nor U28398 (N_28398,N_26159,N_25077);
nand U28399 (N_28399,N_26256,N_24432);
nand U28400 (N_28400,N_26961,N_24872);
and U28401 (N_28401,N_25983,N_24847);
nand U28402 (N_28402,N_26589,N_25399);
xor U28403 (N_28403,N_24759,N_24579);
nand U28404 (N_28404,N_25187,N_25693);
nor U28405 (N_28405,N_26612,N_24496);
xor U28406 (N_28406,N_26776,N_26575);
and U28407 (N_28407,N_25222,N_25438);
and U28408 (N_28408,N_24026,N_25680);
nor U28409 (N_28409,N_25489,N_24536);
nor U28410 (N_28410,N_25070,N_25118);
and U28411 (N_28411,N_26046,N_24814);
nor U28412 (N_28412,N_24560,N_26188);
xnor U28413 (N_28413,N_25942,N_24601);
and U28414 (N_28414,N_24354,N_25845);
xor U28415 (N_28415,N_25329,N_25952);
and U28416 (N_28416,N_26996,N_24152);
nand U28417 (N_28417,N_24531,N_26209);
nand U28418 (N_28418,N_24420,N_26660);
nand U28419 (N_28419,N_25934,N_25546);
and U28420 (N_28420,N_24747,N_26076);
xnor U28421 (N_28421,N_26289,N_25269);
nand U28422 (N_28422,N_25618,N_24263);
and U28423 (N_28423,N_24513,N_26571);
or U28424 (N_28424,N_24362,N_26147);
nand U28425 (N_28425,N_24610,N_25975);
nor U28426 (N_28426,N_24426,N_25492);
or U28427 (N_28427,N_24288,N_25480);
xnor U28428 (N_28428,N_25110,N_26323);
or U28429 (N_28429,N_24977,N_25510);
nor U28430 (N_28430,N_25600,N_26389);
and U28431 (N_28431,N_26523,N_25129);
or U28432 (N_28432,N_25967,N_25871);
xnor U28433 (N_28433,N_26419,N_24058);
nand U28434 (N_28434,N_26546,N_24044);
xnor U28435 (N_28435,N_24344,N_24885);
or U28436 (N_28436,N_25128,N_24774);
nor U28437 (N_28437,N_26127,N_25457);
nor U28438 (N_28438,N_25370,N_24351);
nand U28439 (N_28439,N_24632,N_24673);
or U28440 (N_28440,N_26600,N_26754);
nor U28441 (N_28441,N_26955,N_25256);
xor U28442 (N_28442,N_26607,N_25497);
or U28443 (N_28443,N_26316,N_26298);
xnor U28444 (N_28444,N_24810,N_24295);
nor U28445 (N_28445,N_24182,N_24417);
or U28446 (N_28446,N_24384,N_24487);
nand U28447 (N_28447,N_24879,N_25325);
nor U28448 (N_28448,N_24589,N_24889);
or U28449 (N_28449,N_25454,N_25220);
and U28450 (N_28450,N_26500,N_24449);
and U28451 (N_28451,N_26490,N_25140);
nor U28452 (N_28452,N_24824,N_24494);
or U28453 (N_28453,N_24653,N_26355);
xnor U28454 (N_28454,N_26784,N_26963);
nor U28455 (N_28455,N_26143,N_24948);
nand U28456 (N_28456,N_25528,N_26518);
and U28457 (N_28457,N_25321,N_24561);
nand U28458 (N_28458,N_26659,N_24988);
xor U28459 (N_28459,N_24762,N_24270);
or U28460 (N_28460,N_24936,N_26853);
nand U28461 (N_28461,N_24873,N_26452);
nand U28462 (N_28462,N_26582,N_26454);
nand U28463 (N_28463,N_26943,N_24581);
nand U28464 (N_28464,N_25720,N_24441);
or U28465 (N_28465,N_24787,N_26016);
or U28466 (N_28466,N_26294,N_26005);
nor U28467 (N_28467,N_24707,N_24699);
nand U28468 (N_28468,N_26688,N_24770);
and U28469 (N_28469,N_25103,N_25263);
nand U28470 (N_28470,N_26217,N_24832);
nor U28471 (N_28471,N_25660,N_24189);
nor U28472 (N_28472,N_26153,N_26061);
xnor U28473 (N_28473,N_26548,N_25491);
xor U28474 (N_28474,N_25192,N_26203);
nor U28475 (N_28475,N_24147,N_25771);
xnor U28476 (N_28476,N_24472,N_24480);
xnor U28477 (N_28477,N_24862,N_24975);
nor U28478 (N_28478,N_24169,N_26975);
or U28479 (N_28479,N_26782,N_25002);
nor U28480 (N_28480,N_26092,N_24028);
nor U28481 (N_28481,N_24299,N_24003);
or U28482 (N_28482,N_25984,N_26021);
or U28483 (N_28483,N_25580,N_26702);
nor U28484 (N_28484,N_26710,N_25171);
nand U28485 (N_28485,N_24738,N_25782);
xnor U28486 (N_28486,N_26440,N_26401);
xor U28487 (N_28487,N_24394,N_24482);
nand U28488 (N_28488,N_24534,N_26793);
nand U28489 (N_28489,N_24491,N_26403);
nand U28490 (N_28490,N_24391,N_24816);
nor U28491 (N_28491,N_26646,N_26300);
xnor U28492 (N_28492,N_24925,N_25539);
nor U28493 (N_28493,N_24038,N_26001);
nor U28494 (N_28494,N_24050,N_24142);
or U28495 (N_28495,N_26068,N_26339);
nand U28496 (N_28496,N_24867,N_25221);
nand U28497 (N_28497,N_26400,N_25707);
or U28498 (N_28498,N_26067,N_24499);
xor U28499 (N_28499,N_26812,N_26724);
nor U28500 (N_28500,N_25524,N_24421);
and U28501 (N_28501,N_26440,N_24833);
and U28502 (N_28502,N_25070,N_25972);
or U28503 (N_28503,N_26106,N_26223);
nor U28504 (N_28504,N_26850,N_26831);
nor U28505 (N_28505,N_24559,N_25198);
or U28506 (N_28506,N_26888,N_26751);
or U28507 (N_28507,N_25843,N_24963);
nand U28508 (N_28508,N_25984,N_26091);
or U28509 (N_28509,N_26449,N_25245);
or U28510 (N_28510,N_25814,N_25799);
or U28511 (N_28511,N_26092,N_25202);
xor U28512 (N_28512,N_24428,N_26906);
and U28513 (N_28513,N_26080,N_24606);
and U28514 (N_28514,N_24127,N_26378);
nor U28515 (N_28515,N_24680,N_26299);
or U28516 (N_28516,N_24218,N_24101);
xor U28517 (N_28517,N_25636,N_26215);
and U28518 (N_28518,N_24046,N_25890);
or U28519 (N_28519,N_26867,N_25829);
or U28520 (N_28520,N_25853,N_24969);
nand U28521 (N_28521,N_25905,N_25201);
xor U28522 (N_28522,N_26732,N_24155);
nor U28523 (N_28523,N_26195,N_26039);
xnor U28524 (N_28524,N_25124,N_25306);
nor U28525 (N_28525,N_26753,N_26372);
nor U28526 (N_28526,N_25836,N_26899);
nand U28527 (N_28527,N_24257,N_24121);
nand U28528 (N_28528,N_26609,N_25843);
or U28529 (N_28529,N_24307,N_25964);
xnor U28530 (N_28530,N_24442,N_26636);
or U28531 (N_28531,N_24334,N_24652);
and U28532 (N_28532,N_26167,N_26969);
and U28533 (N_28533,N_25419,N_24667);
xor U28534 (N_28534,N_25232,N_25370);
nand U28535 (N_28535,N_24200,N_26654);
nor U28536 (N_28536,N_26510,N_24522);
or U28537 (N_28537,N_26291,N_25888);
xor U28538 (N_28538,N_26968,N_25951);
xnor U28539 (N_28539,N_25424,N_26825);
and U28540 (N_28540,N_24077,N_26513);
and U28541 (N_28541,N_26965,N_24728);
xor U28542 (N_28542,N_26396,N_25861);
and U28543 (N_28543,N_25064,N_24944);
nand U28544 (N_28544,N_26309,N_24579);
and U28545 (N_28545,N_24910,N_24576);
xor U28546 (N_28546,N_24420,N_25139);
nor U28547 (N_28547,N_24933,N_24209);
and U28548 (N_28548,N_26577,N_26603);
nand U28549 (N_28549,N_25964,N_25301);
or U28550 (N_28550,N_24320,N_24645);
or U28551 (N_28551,N_25725,N_25948);
nor U28552 (N_28552,N_24202,N_25240);
nand U28553 (N_28553,N_24319,N_24562);
nand U28554 (N_28554,N_24577,N_25529);
xor U28555 (N_28555,N_24523,N_24749);
nand U28556 (N_28556,N_24678,N_24654);
or U28557 (N_28557,N_24983,N_24879);
xor U28558 (N_28558,N_25488,N_25592);
xor U28559 (N_28559,N_26508,N_24845);
nor U28560 (N_28560,N_26874,N_25955);
and U28561 (N_28561,N_25925,N_26470);
or U28562 (N_28562,N_25536,N_24422);
nor U28563 (N_28563,N_26830,N_24876);
nor U28564 (N_28564,N_26363,N_26294);
or U28565 (N_28565,N_24436,N_25250);
xnor U28566 (N_28566,N_24548,N_26237);
xor U28567 (N_28567,N_26842,N_25170);
or U28568 (N_28568,N_24075,N_26565);
xor U28569 (N_28569,N_26079,N_26871);
nor U28570 (N_28570,N_25129,N_26645);
nor U28571 (N_28571,N_25686,N_26826);
nand U28572 (N_28572,N_26137,N_26794);
nand U28573 (N_28573,N_25080,N_26261);
or U28574 (N_28574,N_25673,N_25323);
nor U28575 (N_28575,N_26787,N_25087);
nor U28576 (N_28576,N_26442,N_24869);
or U28577 (N_28577,N_25446,N_26516);
or U28578 (N_28578,N_26992,N_24345);
and U28579 (N_28579,N_25488,N_24166);
or U28580 (N_28580,N_25447,N_24633);
and U28581 (N_28581,N_24740,N_25873);
nor U28582 (N_28582,N_26235,N_24531);
nand U28583 (N_28583,N_25489,N_24815);
and U28584 (N_28584,N_26061,N_24347);
nand U28585 (N_28585,N_24675,N_24791);
and U28586 (N_28586,N_24063,N_24193);
xnor U28587 (N_28587,N_26448,N_25836);
and U28588 (N_28588,N_24669,N_26846);
nand U28589 (N_28589,N_24499,N_25303);
xor U28590 (N_28590,N_24293,N_24446);
nand U28591 (N_28591,N_24060,N_24335);
and U28592 (N_28592,N_24190,N_25374);
nand U28593 (N_28593,N_24636,N_24040);
xnor U28594 (N_28594,N_24865,N_24437);
nand U28595 (N_28595,N_24294,N_25075);
and U28596 (N_28596,N_25549,N_25386);
nor U28597 (N_28597,N_25391,N_24385);
xnor U28598 (N_28598,N_26993,N_26155);
and U28599 (N_28599,N_25515,N_25925);
nand U28600 (N_28600,N_24135,N_25279);
nand U28601 (N_28601,N_25083,N_26004);
nor U28602 (N_28602,N_26873,N_25867);
and U28603 (N_28603,N_24353,N_26447);
and U28604 (N_28604,N_26558,N_24724);
and U28605 (N_28605,N_26741,N_24364);
nand U28606 (N_28606,N_25167,N_25003);
nor U28607 (N_28607,N_24586,N_26903);
or U28608 (N_28608,N_26567,N_24166);
and U28609 (N_28609,N_25244,N_24470);
or U28610 (N_28610,N_24417,N_26557);
or U28611 (N_28611,N_25765,N_25822);
nor U28612 (N_28612,N_25084,N_26252);
nor U28613 (N_28613,N_24361,N_24922);
or U28614 (N_28614,N_26871,N_25498);
nor U28615 (N_28615,N_24896,N_25192);
nor U28616 (N_28616,N_25242,N_26844);
nor U28617 (N_28617,N_24297,N_24180);
and U28618 (N_28618,N_25517,N_24968);
nand U28619 (N_28619,N_25508,N_24018);
nor U28620 (N_28620,N_25261,N_26881);
xnor U28621 (N_28621,N_26177,N_25970);
xor U28622 (N_28622,N_24029,N_26655);
xor U28623 (N_28623,N_25077,N_25798);
or U28624 (N_28624,N_26573,N_25600);
nand U28625 (N_28625,N_24972,N_25051);
nand U28626 (N_28626,N_25817,N_24195);
xor U28627 (N_28627,N_25330,N_26966);
nand U28628 (N_28628,N_24824,N_25590);
or U28629 (N_28629,N_25402,N_25974);
nand U28630 (N_28630,N_26422,N_26948);
or U28631 (N_28631,N_24872,N_26888);
or U28632 (N_28632,N_26401,N_24346);
or U28633 (N_28633,N_24323,N_25460);
xor U28634 (N_28634,N_25556,N_25568);
and U28635 (N_28635,N_24289,N_26052);
nand U28636 (N_28636,N_24409,N_26158);
nor U28637 (N_28637,N_24341,N_26954);
or U28638 (N_28638,N_26540,N_24050);
or U28639 (N_28639,N_24845,N_26957);
or U28640 (N_28640,N_24869,N_25264);
xor U28641 (N_28641,N_25195,N_24857);
xor U28642 (N_28642,N_24787,N_25884);
or U28643 (N_28643,N_25683,N_24472);
and U28644 (N_28644,N_24624,N_26536);
nor U28645 (N_28645,N_25106,N_26694);
nand U28646 (N_28646,N_25659,N_25168);
or U28647 (N_28647,N_26662,N_26401);
nand U28648 (N_28648,N_26562,N_26966);
and U28649 (N_28649,N_25055,N_26857);
or U28650 (N_28650,N_25105,N_24283);
or U28651 (N_28651,N_24876,N_26988);
xnor U28652 (N_28652,N_25891,N_24271);
nand U28653 (N_28653,N_24823,N_24008);
or U28654 (N_28654,N_25731,N_26173);
xnor U28655 (N_28655,N_24837,N_26612);
or U28656 (N_28656,N_24149,N_24354);
and U28657 (N_28657,N_24968,N_26104);
xor U28658 (N_28658,N_25177,N_24685);
and U28659 (N_28659,N_26089,N_24530);
nor U28660 (N_28660,N_24557,N_26592);
xor U28661 (N_28661,N_25033,N_26290);
xnor U28662 (N_28662,N_26455,N_24324);
and U28663 (N_28663,N_25223,N_25829);
nand U28664 (N_28664,N_26983,N_26413);
and U28665 (N_28665,N_24041,N_26104);
xnor U28666 (N_28666,N_24097,N_24688);
nor U28667 (N_28667,N_24746,N_26120);
and U28668 (N_28668,N_24464,N_25445);
xnor U28669 (N_28669,N_26647,N_24940);
and U28670 (N_28670,N_26161,N_26319);
or U28671 (N_28671,N_26787,N_26658);
nor U28672 (N_28672,N_25028,N_25304);
xor U28673 (N_28673,N_25579,N_26653);
nor U28674 (N_28674,N_25320,N_25946);
or U28675 (N_28675,N_24447,N_26907);
nor U28676 (N_28676,N_26683,N_24660);
or U28677 (N_28677,N_25855,N_24310);
and U28678 (N_28678,N_24397,N_25911);
xor U28679 (N_28679,N_25642,N_24717);
xor U28680 (N_28680,N_26312,N_25406);
xor U28681 (N_28681,N_26486,N_25810);
or U28682 (N_28682,N_24553,N_25949);
and U28683 (N_28683,N_24977,N_24479);
nand U28684 (N_28684,N_24779,N_24366);
or U28685 (N_28685,N_26386,N_24303);
and U28686 (N_28686,N_26393,N_25735);
nor U28687 (N_28687,N_26597,N_24379);
or U28688 (N_28688,N_25652,N_26743);
or U28689 (N_28689,N_25453,N_24347);
and U28690 (N_28690,N_24943,N_26536);
nor U28691 (N_28691,N_26359,N_26007);
nor U28692 (N_28692,N_26881,N_26756);
nor U28693 (N_28693,N_25370,N_25198);
and U28694 (N_28694,N_24714,N_25895);
nor U28695 (N_28695,N_26042,N_25466);
and U28696 (N_28696,N_24133,N_26926);
nand U28697 (N_28697,N_25997,N_24215);
nand U28698 (N_28698,N_25777,N_24742);
nand U28699 (N_28699,N_26437,N_24616);
nor U28700 (N_28700,N_24089,N_26744);
xor U28701 (N_28701,N_25471,N_25951);
xnor U28702 (N_28702,N_25569,N_24510);
or U28703 (N_28703,N_26588,N_26420);
nand U28704 (N_28704,N_25533,N_24960);
nand U28705 (N_28705,N_26402,N_25319);
or U28706 (N_28706,N_26497,N_24457);
xor U28707 (N_28707,N_26894,N_24282);
nor U28708 (N_28708,N_24708,N_24322);
and U28709 (N_28709,N_25315,N_25016);
and U28710 (N_28710,N_26397,N_25370);
and U28711 (N_28711,N_26394,N_25149);
or U28712 (N_28712,N_24146,N_25027);
nor U28713 (N_28713,N_24549,N_24738);
and U28714 (N_28714,N_25980,N_25749);
xor U28715 (N_28715,N_26216,N_25028);
and U28716 (N_28716,N_26574,N_26158);
and U28717 (N_28717,N_25102,N_25459);
nand U28718 (N_28718,N_25593,N_26287);
or U28719 (N_28719,N_25267,N_24071);
nor U28720 (N_28720,N_24789,N_26606);
nand U28721 (N_28721,N_26737,N_24705);
nand U28722 (N_28722,N_24479,N_26667);
and U28723 (N_28723,N_24674,N_24272);
and U28724 (N_28724,N_25864,N_24135);
xnor U28725 (N_28725,N_26073,N_25567);
nor U28726 (N_28726,N_26590,N_26745);
xnor U28727 (N_28727,N_26660,N_24393);
xnor U28728 (N_28728,N_26831,N_25129);
xnor U28729 (N_28729,N_25796,N_26219);
nand U28730 (N_28730,N_26177,N_24598);
xor U28731 (N_28731,N_24432,N_25152);
or U28732 (N_28732,N_24218,N_25111);
and U28733 (N_28733,N_25637,N_25015);
nor U28734 (N_28734,N_25631,N_24376);
nor U28735 (N_28735,N_26252,N_25303);
and U28736 (N_28736,N_24916,N_26014);
nand U28737 (N_28737,N_25791,N_26563);
or U28738 (N_28738,N_26774,N_25479);
nand U28739 (N_28739,N_25007,N_26506);
and U28740 (N_28740,N_24929,N_26574);
or U28741 (N_28741,N_25563,N_26957);
nor U28742 (N_28742,N_24618,N_24569);
or U28743 (N_28743,N_24168,N_26762);
nand U28744 (N_28744,N_25338,N_26946);
and U28745 (N_28745,N_26338,N_26847);
or U28746 (N_28746,N_25382,N_25515);
and U28747 (N_28747,N_26129,N_26132);
nor U28748 (N_28748,N_24883,N_26077);
xor U28749 (N_28749,N_26871,N_24991);
or U28750 (N_28750,N_26649,N_24913);
nor U28751 (N_28751,N_24135,N_25425);
nor U28752 (N_28752,N_26674,N_24384);
nor U28753 (N_28753,N_25847,N_26380);
xor U28754 (N_28754,N_26247,N_26759);
nor U28755 (N_28755,N_25671,N_24149);
or U28756 (N_28756,N_25670,N_25031);
nor U28757 (N_28757,N_26626,N_26386);
and U28758 (N_28758,N_26397,N_26795);
or U28759 (N_28759,N_24906,N_26244);
nand U28760 (N_28760,N_25926,N_26516);
nor U28761 (N_28761,N_25920,N_24469);
nand U28762 (N_28762,N_25577,N_26133);
or U28763 (N_28763,N_24306,N_26998);
xnor U28764 (N_28764,N_25482,N_24716);
and U28765 (N_28765,N_26983,N_25307);
or U28766 (N_28766,N_25577,N_25309);
nor U28767 (N_28767,N_26341,N_25184);
and U28768 (N_28768,N_24616,N_26160);
nand U28769 (N_28769,N_25290,N_24339);
nand U28770 (N_28770,N_26905,N_24238);
and U28771 (N_28771,N_26163,N_26942);
and U28772 (N_28772,N_24246,N_25753);
or U28773 (N_28773,N_26398,N_26223);
nand U28774 (N_28774,N_26740,N_25128);
nor U28775 (N_28775,N_24502,N_25708);
and U28776 (N_28776,N_25490,N_24958);
and U28777 (N_28777,N_26784,N_24482);
xnor U28778 (N_28778,N_25934,N_26534);
nor U28779 (N_28779,N_26627,N_24083);
or U28780 (N_28780,N_26547,N_26440);
and U28781 (N_28781,N_24906,N_26301);
or U28782 (N_28782,N_24744,N_26288);
xor U28783 (N_28783,N_25712,N_26150);
and U28784 (N_28784,N_24964,N_24159);
xor U28785 (N_28785,N_25455,N_24030);
or U28786 (N_28786,N_26642,N_24912);
or U28787 (N_28787,N_26085,N_26812);
nor U28788 (N_28788,N_26163,N_24366);
nor U28789 (N_28789,N_26952,N_26337);
or U28790 (N_28790,N_25590,N_24459);
nand U28791 (N_28791,N_26251,N_26668);
nand U28792 (N_28792,N_24803,N_25961);
and U28793 (N_28793,N_24001,N_25203);
or U28794 (N_28794,N_24075,N_26745);
xor U28795 (N_28795,N_26170,N_26389);
or U28796 (N_28796,N_25665,N_25249);
nor U28797 (N_28797,N_24455,N_25911);
nand U28798 (N_28798,N_24114,N_26052);
nor U28799 (N_28799,N_25879,N_25275);
nand U28800 (N_28800,N_25451,N_25424);
xnor U28801 (N_28801,N_26542,N_24021);
and U28802 (N_28802,N_24692,N_24062);
nor U28803 (N_28803,N_26091,N_25864);
and U28804 (N_28804,N_26119,N_24141);
xor U28805 (N_28805,N_25488,N_26066);
or U28806 (N_28806,N_26798,N_26497);
nand U28807 (N_28807,N_24058,N_25442);
xnor U28808 (N_28808,N_24887,N_25933);
nand U28809 (N_28809,N_26175,N_24691);
or U28810 (N_28810,N_25635,N_26126);
or U28811 (N_28811,N_25867,N_25123);
nor U28812 (N_28812,N_26062,N_24131);
or U28813 (N_28813,N_26256,N_24729);
nand U28814 (N_28814,N_24762,N_25772);
and U28815 (N_28815,N_25924,N_24073);
or U28816 (N_28816,N_26390,N_26564);
and U28817 (N_28817,N_25004,N_25712);
or U28818 (N_28818,N_24708,N_25098);
xnor U28819 (N_28819,N_24546,N_24287);
nor U28820 (N_28820,N_25300,N_25420);
nand U28821 (N_28821,N_25716,N_25698);
and U28822 (N_28822,N_24442,N_24690);
or U28823 (N_28823,N_26099,N_26954);
xnor U28824 (N_28824,N_25735,N_25240);
or U28825 (N_28825,N_25647,N_26580);
xnor U28826 (N_28826,N_25899,N_25394);
and U28827 (N_28827,N_24632,N_24298);
nand U28828 (N_28828,N_26910,N_24722);
and U28829 (N_28829,N_26986,N_24165);
and U28830 (N_28830,N_26746,N_25680);
nor U28831 (N_28831,N_25245,N_26004);
or U28832 (N_28832,N_25018,N_24084);
or U28833 (N_28833,N_26149,N_26978);
xnor U28834 (N_28834,N_25397,N_25425);
nand U28835 (N_28835,N_24826,N_26877);
and U28836 (N_28836,N_24781,N_24148);
and U28837 (N_28837,N_24519,N_25046);
xor U28838 (N_28838,N_26737,N_24079);
and U28839 (N_28839,N_24550,N_24621);
or U28840 (N_28840,N_24077,N_24355);
nor U28841 (N_28841,N_24314,N_24357);
nor U28842 (N_28842,N_25037,N_26820);
and U28843 (N_28843,N_25309,N_26306);
nand U28844 (N_28844,N_25265,N_25090);
xor U28845 (N_28845,N_26270,N_25819);
xnor U28846 (N_28846,N_25388,N_26737);
xnor U28847 (N_28847,N_25722,N_24540);
nand U28848 (N_28848,N_25065,N_25561);
xnor U28849 (N_28849,N_24213,N_26620);
nand U28850 (N_28850,N_26970,N_25853);
nor U28851 (N_28851,N_25563,N_24547);
or U28852 (N_28852,N_25728,N_24071);
and U28853 (N_28853,N_25610,N_26947);
or U28854 (N_28854,N_25069,N_25496);
and U28855 (N_28855,N_25575,N_24191);
nor U28856 (N_28856,N_25239,N_24214);
and U28857 (N_28857,N_26224,N_24351);
and U28858 (N_28858,N_24957,N_25720);
nor U28859 (N_28859,N_25737,N_25016);
xor U28860 (N_28860,N_25700,N_24780);
nor U28861 (N_28861,N_24104,N_25829);
xnor U28862 (N_28862,N_25550,N_24677);
and U28863 (N_28863,N_25160,N_24396);
nor U28864 (N_28864,N_25841,N_24522);
nand U28865 (N_28865,N_25902,N_24720);
nor U28866 (N_28866,N_26167,N_25428);
or U28867 (N_28867,N_26532,N_26821);
and U28868 (N_28868,N_25295,N_26564);
nand U28869 (N_28869,N_25276,N_24915);
nor U28870 (N_28870,N_25457,N_25494);
and U28871 (N_28871,N_26184,N_24091);
and U28872 (N_28872,N_26490,N_26253);
and U28873 (N_28873,N_24633,N_26425);
nor U28874 (N_28874,N_26307,N_24691);
nor U28875 (N_28875,N_24163,N_26557);
nand U28876 (N_28876,N_26025,N_26884);
and U28877 (N_28877,N_26312,N_24468);
nor U28878 (N_28878,N_25253,N_24260);
nand U28879 (N_28879,N_26206,N_24010);
nor U28880 (N_28880,N_26091,N_25285);
or U28881 (N_28881,N_25907,N_26704);
or U28882 (N_28882,N_24524,N_25543);
or U28883 (N_28883,N_24367,N_25701);
and U28884 (N_28884,N_26490,N_26421);
and U28885 (N_28885,N_25197,N_25687);
nor U28886 (N_28886,N_25531,N_25863);
or U28887 (N_28887,N_24639,N_26980);
xnor U28888 (N_28888,N_25896,N_24452);
and U28889 (N_28889,N_25027,N_24582);
or U28890 (N_28890,N_26286,N_24790);
or U28891 (N_28891,N_26313,N_26842);
or U28892 (N_28892,N_24304,N_26611);
xor U28893 (N_28893,N_24777,N_25225);
xnor U28894 (N_28894,N_25471,N_24773);
xor U28895 (N_28895,N_26484,N_25490);
or U28896 (N_28896,N_25342,N_26309);
or U28897 (N_28897,N_26904,N_26802);
or U28898 (N_28898,N_25554,N_25390);
nand U28899 (N_28899,N_24326,N_25476);
and U28900 (N_28900,N_26221,N_24302);
or U28901 (N_28901,N_24983,N_25601);
xnor U28902 (N_28902,N_25328,N_24550);
or U28903 (N_28903,N_24725,N_26679);
nand U28904 (N_28904,N_25432,N_25583);
and U28905 (N_28905,N_25609,N_25183);
or U28906 (N_28906,N_25529,N_24293);
and U28907 (N_28907,N_24095,N_25882);
or U28908 (N_28908,N_25157,N_26245);
and U28909 (N_28909,N_26403,N_26670);
and U28910 (N_28910,N_26325,N_24839);
and U28911 (N_28911,N_24301,N_24055);
xor U28912 (N_28912,N_24993,N_24627);
nand U28913 (N_28913,N_26793,N_25783);
or U28914 (N_28914,N_25695,N_24967);
xor U28915 (N_28915,N_24982,N_25123);
xnor U28916 (N_28916,N_24348,N_26205);
nand U28917 (N_28917,N_26106,N_24051);
nor U28918 (N_28918,N_24640,N_25882);
xor U28919 (N_28919,N_25924,N_25243);
nand U28920 (N_28920,N_25377,N_25140);
xor U28921 (N_28921,N_24602,N_25097);
xor U28922 (N_28922,N_25041,N_26385);
xor U28923 (N_28923,N_25544,N_25906);
or U28924 (N_28924,N_25244,N_26687);
and U28925 (N_28925,N_25086,N_25605);
and U28926 (N_28926,N_26341,N_25989);
or U28927 (N_28927,N_24367,N_25612);
and U28928 (N_28928,N_26583,N_26316);
nor U28929 (N_28929,N_24102,N_26316);
or U28930 (N_28930,N_26812,N_26309);
nor U28931 (N_28931,N_25631,N_24684);
nor U28932 (N_28932,N_24100,N_25365);
and U28933 (N_28933,N_25594,N_25180);
and U28934 (N_28934,N_24409,N_25621);
nand U28935 (N_28935,N_26680,N_25312);
nand U28936 (N_28936,N_25548,N_24751);
or U28937 (N_28937,N_26513,N_26406);
nand U28938 (N_28938,N_24084,N_24962);
nor U28939 (N_28939,N_26984,N_26759);
xor U28940 (N_28940,N_24437,N_25599);
nand U28941 (N_28941,N_25459,N_25991);
and U28942 (N_28942,N_24036,N_26737);
or U28943 (N_28943,N_25925,N_25910);
nand U28944 (N_28944,N_25227,N_24485);
xor U28945 (N_28945,N_24904,N_26223);
nand U28946 (N_28946,N_26173,N_25812);
and U28947 (N_28947,N_26209,N_25945);
nor U28948 (N_28948,N_25797,N_26306);
or U28949 (N_28949,N_26502,N_24035);
nand U28950 (N_28950,N_25720,N_24249);
and U28951 (N_28951,N_25066,N_24950);
nor U28952 (N_28952,N_25496,N_26289);
and U28953 (N_28953,N_26314,N_26572);
nor U28954 (N_28954,N_26677,N_25650);
nor U28955 (N_28955,N_26857,N_24512);
xor U28956 (N_28956,N_25167,N_25250);
or U28957 (N_28957,N_26230,N_24847);
and U28958 (N_28958,N_25518,N_25995);
xnor U28959 (N_28959,N_26715,N_24821);
nand U28960 (N_28960,N_26188,N_24246);
or U28961 (N_28961,N_25822,N_26839);
nand U28962 (N_28962,N_25483,N_24131);
or U28963 (N_28963,N_25142,N_25861);
nand U28964 (N_28964,N_25644,N_25308);
nor U28965 (N_28965,N_25785,N_26347);
and U28966 (N_28966,N_24208,N_24533);
or U28967 (N_28967,N_26560,N_26932);
xnor U28968 (N_28968,N_24913,N_24734);
nand U28969 (N_28969,N_26195,N_24716);
or U28970 (N_28970,N_25154,N_25208);
and U28971 (N_28971,N_26990,N_24129);
xor U28972 (N_28972,N_24223,N_24308);
and U28973 (N_28973,N_25679,N_26189);
nor U28974 (N_28974,N_25974,N_26842);
nand U28975 (N_28975,N_26308,N_25958);
or U28976 (N_28976,N_25673,N_26000);
and U28977 (N_28977,N_24361,N_24508);
xor U28978 (N_28978,N_24807,N_24588);
nor U28979 (N_28979,N_25624,N_25956);
or U28980 (N_28980,N_24485,N_26911);
nand U28981 (N_28981,N_25585,N_26317);
xor U28982 (N_28982,N_25005,N_24630);
nor U28983 (N_28983,N_25394,N_25398);
or U28984 (N_28984,N_24067,N_24103);
or U28985 (N_28985,N_25455,N_25474);
nor U28986 (N_28986,N_26305,N_24785);
nand U28987 (N_28987,N_25502,N_26148);
and U28988 (N_28988,N_25016,N_26271);
and U28989 (N_28989,N_25927,N_26191);
nor U28990 (N_28990,N_26179,N_26130);
nand U28991 (N_28991,N_24383,N_25288);
xnor U28992 (N_28992,N_24630,N_24552);
xor U28993 (N_28993,N_25221,N_26913);
nor U28994 (N_28994,N_26867,N_26298);
xor U28995 (N_28995,N_25222,N_24031);
xor U28996 (N_28996,N_24648,N_26502);
and U28997 (N_28997,N_26255,N_26940);
xnor U28998 (N_28998,N_26790,N_24320);
nand U28999 (N_28999,N_25462,N_24437);
or U29000 (N_29000,N_26286,N_25312);
xor U29001 (N_29001,N_26621,N_26619);
nor U29002 (N_29002,N_26050,N_26564);
xnor U29003 (N_29003,N_24029,N_24464);
and U29004 (N_29004,N_26796,N_24995);
nor U29005 (N_29005,N_26235,N_24005);
nand U29006 (N_29006,N_24114,N_26035);
and U29007 (N_29007,N_25447,N_25891);
nor U29008 (N_29008,N_26955,N_24859);
nand U29009 (N_29009,N_26669,N_25426);
or U29010 (N_29010,N_24575,N_26378);
nor U29011 (N_29011,N_26945,N_25728);
nand U29012 (N_29012,N_25270,N_24472);
xor U29013 (N_29013,N_24672,N_25495);
or U29014 (N_29014,N_26893,N_24147);
and U29015 (N_29015,N_25525,N_25035);
and U29016 (N_29016,N_24180,N_25831);
or U29017 (N_29017,N_26770,N_26273);
nor U29018 (N_29018,N_25068,N_25652);
nor U29019 (N_29019,N_26616,N_26792);
nor U29020 (N_29020,N_24468,N_24928);
or U29021 (N_29021,N_25318,N_26157);
or U29022 (N_29022,N_25734,N_26150);
nor U29023 (N_29023,N_26293,N_24525);
xnor U29024 (N_29024,N_24366,N_25814);
nor U29025 (N_29025,N_24498,N_25379);
nand U29026 (N_29026,N_26530,N_24667);
or U29027 (N_29027,N_24928,N_26638);
nor U29028 (N_29028,N_26036,N_26669);
xnor U29029 (N_29029,N_26692,N_26457);
nand U29030 (N_29030,N_26651,N_25726);
xnor U29031 (N_29031,N_24997,N_24113);
nor U29032 (N_29032,N_25724,N_25733);
or U29033 (N_29033,N_24200,N_25712);
nand U29034 (N_29034,N_25142,N_26785);
or U29035 (N_29035,N_24314,N_26387);
or U29036 (N_29036,N_26604,N_26392);
xor U29037 (N_29037,N_26561,N_25234);
and U29038 (N_29038,N_25425,N_25871);
or U29039 (N_29039,N_26590,N_25493);
nand U29040 (N_29040,N_24382,N_24327);
or U29041 (N_29041,N_24812,N_24298);
nand U29042 (N_29042,N_24904,N_26623);
or U29043 (N_29043,N_25059,N_24664);
and U29044 (N_29044,N_26798,N_25634);
and U29045 (N_29045,N_25704,N_26542);
nor U29046 (N_29046,N_26672,N_24323);
xor U29047 (N_29047,N_24352,N_26014);
nand U29048 (N_29048,N_26919,N_26839);
or U29049 (N_29049,N_26579,N_24107);
and U29050 (N_29050,N_26875,N_26851);
nor U29051 (N_29051,N_26308,N_25337);
or U29052 (N_29052,N_25446,N_25736);
nor U29053 (N_29053,N_24649,N_24107);
nand U29054 (N_29054,N_25226,N_26531);
or U29055 (N_29055,N_24338,N_24558);
and U29056 (N_29056,N_24167,N_26022);
and U29057 (N_29057,N_26444,N_24241);
nor U29058 (N_29058,N_26268,N_26616);
or U29059 (N_29059,N_25280,N_24171);
nor U29060 (N_29060,N_26244,N_26248);
nor U29061 (N_29061,N_24356,N_26722);
nand U29062 (N_29062,N_26191,N_24743);
or U29063 (N_29063,N_24863,N_26655);
nand U29064 (N_29064,N_25016,N_26226);
xor U29065 (N_29065,N_24871,N_24854);
nand U29066 (N_29066,N_24178,N_24741);
or U29067 (N_29067,N_26763,N_25665);
or U29068 (N_29068,N_24509,N_24894);
nand U29069 (N_29069,N_24165,N_26717);
and U29070 (N_29070,N_25229,N_24038);
and U29071 (N_29071,N_25104,N_25759);
nor U29072 (N_29072,N_25520,N_25496);
xnor U29073 (N_29073,N_25032,N_24049);
or U29074 (N_29074,N_26455,N_26116);
xnor U29075 (N_29075,N_24367,N_25550);
or U29076 (N_29076,N_25952,N_25892);
nand U29077 (N_29077,N_24034,N_25423);
nand U29078 (N_29078,N_24904,N_24952);
and U29079 (N_29079,N_25349,N_24777);
xnor U29080 (N_29080,N_24954,N_26089);
xnor U29081 (N_29081,N_25282,N_25039);
and U29082 (N_29082,N_25154,N_26654);
nor U29083 (N_29083,N_24316,N_25572);
xor U29084 (N_29084,N_25640,N_26264);
and U29085 (N_29085,N_26081,N_26500);
or U29086 (N_29086,N_25340,N_25026);
nor U29087 (N_29087,N_26265,N_26869);
or U29088 (N_29088,N_26227,N_25880);
and U29089 (N_29089,N_24172,N_24418);
xnor U29090 (N_29090,N_25407,N_24102);
or U29091 (N_29091,N_25726,N_24505);
and U29092 (N_29092,N_26751,N_25021);
nor U29093 (N_29093,N_26247,N_25654);
xor U29094 (N_29094,N_26604,N_24119);
and U29095 (N_29095,N_25510,N_24384);
and U29096 (N_29096,N_25476,N_24860);
nor U29097 (N_29097,N_26187,N_26128);
xnor U29098 (N_29098,N_24498,N_24325);
and U29099 (N_29099,N_24588,N_24217);
nand U29100 (N_29100,N_26396,N_26018);
nand U29101 (N_29101,N_25045,N_26999);
or U29102 (N_29102,N_26057,N_26373);
xnor U29103 (N_29103,N_24772,N_25118);
xnor U29104 (N_29104,N_26940,N_26845);
xor U29105 (N_29105,N_26244,N_26460);
or U29106 (N_29106,N_25801,N_25661);
and U29107 (N_29107,N_25063,N_24049);
or U29108 (N_29108,N_26426,N_26623);
xor U29109 (N_29109,N_26045,N_26069);
or U29110 (N_29110,N_25254,N_25389);
xor U29111 (N_29111,N_25509,N_24280);
nor U29112 (N_29112,N_24784,N_24418);
nand U29113 (N_29113,N_24992,N_26407);
nor U29114 (N_29114,N_25079,N_24348);
or U29115 (N_29115,N_25924,N_26394);
nand U29116 (N_29116,N_26502,N_24170);
or U29117 (N_29117,N_26018,N_26091);
or U29118 (N_29118,N_26580,N_26822);
and U29119 (N_29119,N_25816,N_26335);
or U29120 (N_29120,N_24970,N_25569);
nand U29121 (N_29121,N_25110,N_24583);
xnor U29122 (N_29122,N_25349,N_25005);
nand U29123 (N_29123,N_25043,N_25015);
or U29124 (N_29124,N_25147,N_26458);
nand U29125 (N_29125,N_24923,N_24872);
nor U29126 (N_29126,N_25873,N_24806);
and U29127 (N_29127,N_24709,N_24238);
and U29128 (N_29128,N_26479,N_24023);
xor U29129 (N_29129,N_24219,N_26772);
nand U29130 (N_29130,N_26096,N_26819);
nor U29131 (N_29131,N_24534,N_25111);
and U29132 (N_29132,N_26851,N_25616);
nor U29133 (N_29133,N_25715,N_24262);
xor U29134 (N_29134,N_25133,N_26496);
nand U29135 (N_29135,N_25818,N_25462);
or U29136 (N_29136,N_26823,N_26857);
and U29137 (N_29137,N_26415,N_26299);
and U29138 (N_29138,N_25316,N_24905);
nand U29139 (N_29139,N_24803,N_26803);
nand U29140 (N_29140,N_26151,N_25613);
or U29141 (N_29141,N_25773,N_25758);
or U29142 (N_29142,N_26922,N_24202);
or U29143 (N_29143,N_26242,N_24524);
or U29144 (N_29144,N_24981,N_26243);
xnor U29145 (N_29145,N_25501,N_25388);
xor U29146 (N_29146,N_24549,N_26799);
nor U29147 (N_29147,N_24150,N_26701);
and U29148 (N_29148,N_24265,N_24274);
or U29149 (N_29149,N_24493,N_25586);
nand U29150 (N_29150,N_24239,N_24918);
xnor U29151 (N_29151,N_25440,N_25095);
xor U29152 (N_29152,N_26259,N_25899);
or U29153 (N_29153,N_24559,N_25865);
nor U29154 (N_29154,N_24350,N_26490);
nand U29155 (N_29155,N_24572,N_25035);
xnor U29156 (N_29156,N_25264,N_25929);
nand U29157 (N_29157,N_24625,N_24978);
and U29158 (N_29158,N_25456,N_26686);
nor U29159 (N_29159,N_24663,N_26432);
or U29160 (N_29160,N_24107,N_24878);
nand U29161 (N_29161,N_26773,N_26935);
xor U29162 (N_29162,N_26569,N_25090);
xnor U29163 (N_29163,N_25220,N_25187);
nand U29164 (N_29164,N_25266,N_24770);
nand U29165 (N_29165,N_26288,N_25791);
nand U29166 (N_29166,N_26942,N_26440);
or U29167 (N_29167,N_24758,N_25613);
and U29168 (N_29168,N_26046,N_24259);
nor U29169 (N_29169,N_25770,N_25336);
nand U29170 (N_29170,N_26768,N_26802);
and U29171 (N_29171,N_24573,N_24446);
nor U29172 (N_29172,N_25518,N_24914);
and U29173 (N_29173,N_26866,N_24228);
and U29174 (N_29174,N_24992,N_26520);
nand U29175 (N_29175,N_26101,N_25740);
nand U29176 (N_29176,N_26947,N_26887);
and U29177 (N_29177,N_24540,N_25875);
and U29178 (N_29178,N_25004,N_25438);
and U29179 (N_29179,N_25644,N_24381);
nand U29180 (N_29180,N_26249,N_26526);
or U29181 (N_29181,N_25558,N_26017);
nor U29182 (N_29182,N_24203,N_24377);
xor U29183 (N_29183,N_26512,N_24251);
xor U29184 (N_29184,N_25276,N_24609);
xnor U29185 (N_29185,N_25587,N_24144);
and U29186 (N_29186,N_25649,N_25709);
and U29187 (N_29187,N_25000,N_25651);
nand U29188 (N_29188,N_25042,N_24471);
nor U29189 (N_29189,N_25217,N_25397);
xnor U29190 (N_29190,N_24179,N_24535);
nor U29191 (N_29191,N_26887,N_24398);
or U29192 (N_29192,N_25451,N_24469);
xnor U29193 (N_29193,N_26816,N_25288);
nor U29194 (N_29194,N_25226,N_26008);
nand U29195 (N_29195,N_25400,N_25459);
nor U29196 (N_29196,N_26446,N_26290);
xor U29197 (N_29197,N_26722,N_24308);
nor U29198 (N_29198,N_26273,N_26848);
nand U29199 (N_29199,N_25325,N_26023);
nand U29200 (N_29200,N_24742,N_25353);
or U29201 (N_29201,N_26895,N_25440);
nand U29202 (N_29202,N_24400,N_24218);
xor U29203 (N_29203,N_26033,N_26982);
xnor U29204 (N_29204,N_25844,N_24443);
and U29205 (N_29205,N_24798,N_26481);
or U29206 (N_29206,N_26450,N_26671);
or U29207 (N_29207,N_26482,N_26479);
or U29208 (N_29208,N_26596,N_25797);
or U29209 (N_29209,N_24518,N_26770);
xor U29210 (N_29210,N_26548,N_26844);
nor U29211 (N_29211,N_25991,N_24431);
or U29212 (N_29212,N_24976,N_24440);
xnor U29213 (N_29213,N_26909,N_26713);
xnor U29214 (N_29214,N_25241,N_24226);
and U29215 (N_29215,N_26925,N_26367);
or U29216 (N_29216,N_25478,N_25420);
nor U29217 (N_29217,N_24099,N_26744);
nor U29218 (N_29218,N_24189,N_24469);
nor U29219 (N_29219,N_26229,N_26506);
or U29220 (N_29220,N_24290,N_26213);
or U29221 (N_29221,N_25181,N_26235);
and U29222 (N_29222,N_26368,N_25616);
or U29223 (N_29223,N_26398,N_26007);
nand U29224 (N_29224,N_25060,N_25287);
nor U29225 (N_29225,N_26615,N_25006);
xnor U29226 (N_29226,N_26225,N_25038);
nor U29227 (N_29227,N_26214,N_24868);
nand U29228 (N_29228,N_26420,N_25509);
xnor U29229 (N_29229,N_24670,N_24284);
or U29230 (N_29230,N_25135,N_26488);
nand U29231 (N_29231,N_26670,N_25847);
and U29232 (N_29232,N_25083,N_26624);
nor U29233 (N_29233,N_26495,N_26064);
and U29234 (N_29234,N_24146,N_26656);
and U29235 (N_29235,N_24943,N_25635);
xor U29236 (N_29236,N_24976,N_24301);
nor U29237 (N_29237,N_25060,N_25434);
and U29238 (N_29238,N_26353,N_24803);
or U29239 (N_29239,N_24823,N_24601);
xor U29240 (N_29240,N_26221,N_26050);
and U29241 (N_29241,N_25525,N_26014);
or U29242 (N_29242,N_25569,N_26488);
nor U29243 (N_29243,N_24924,N_25468);
xor U29244 (N_29244,N_26199,N_25977);
xor U29245 (N_29245,N_26278,N_26704);
and U29246 (N_29246,N_24135,N_26182);
nand U29247 (N_29247,N_26391,N_25933);
nand U29248 (N_29248,N_25818,N_25719);
nor U29249 (N_29249,N_26226,N_24662);
and U29250 (N_29250,N_25682,N_26130);
nand U29251 (N_29251,N_25357,N_25059);
nor U29252 (N_29252,N_26139,N_26155);
nand U29253 (N_29253,N_24768,N_24831);
and U29254 (N_29254,N_25386,N_26972);
xor U29255 (N_29255,N_25149,N_25211);
nand U29256 (N_29256,N_24737,N_26924);
xor U29257 (N_29257,N_24968,N_24952);
or U29258 (N_29258,N_26242,N_26598);
and U29259 (N_29259,N_26355,N_26044);
and U29260 (N_29260,N_24545,N_24096);
nor U29261 (N_29261,N_26029,N_26161);
xor U29262 (N_29262,N_24581,N_25157);
nand U29263 (N_29263,N_26872,N_26883);
nor U29264 (N_29264,N_24725,N_25544);
and U29265 (N_29265,N_24609,N_26228);
nand U29266 (N_29266,N_25745,N_24027);
xnor U29267 (N_29267,N_26170,N_25482);
and U29268 (N_29268,N_25904,N_25695);
or U29269 (N_29269,N_25214,N_25287);
xor U29270 (N_29270,N_25801,N_24171);
nand U29271 (N_29271,N_24614,N_26022);
and U29272 (N_29272,N_26767,N_25709);
nor U29273 (N_29273,N_26674,N_24827);
and U29274 (N_29274,N_24106,N_26545);
or U29275 (N_29275,N_26875,N_25362);
nor U29276 (N_29276,N_25059,N_24523);
xor U29277 (N_29277,N_25779,N_26601);
xor U29278 (N_29278,N_25561,N_25040);
nor U29279 (N_29279,N_26909,N_25249);
or U29280 (N_29280,N_24279,N_24382);
nor U29281 (N_29281,N_26420,N_26788);
nand U29282 (N_29282,N_24729,N_24683);
nor U29283 (N_29283,N_26392,N_26145);
and U29284 (N_29284,N_25534,N_25795);
nand U29285 (N_29285,N_24665,N_24212);
nand U29286 (N_29286,N_24355,N_25564);
or U29287 (N_29287,N_24922,N_25382);
xor U29288 (N_29288,N_24667,N_26554);
or U29289 (N_29289,N_26831,N_25697);
nor U29290 (N_29290,N_24101,N_24582);
nor U29291 (N_29291,N_24455,N_26417);
and U29292 (N_29292,N_26954,N_24652);
and U29293 (N_29293,N_25506,N_25850);
nor U29294 (N_29294,N_26140,N_26635);
or U29295 (N_29295,N_26310,N_25667);
nor U29296 (N_29296,N_25314,N_25067);
xnor U29297 (N_29297,N_26022,N_25027);
and U29298 (N_29298,N_26226,N_25059);
nor U29299 (N_29299,N_24187,N_25605);
xnor U29300 (N_29300,N_24655,N_24027);
nor U29301 (N_29301,N_25851,N_26859);
and U29302 (N_29302,N_26559,N_25109);
xor U29303 (N_29303,N_26807,N_25304);
nand U29304 (N_29304,N_24083,N_24346);
nor U29305 (N_29305,N_26325,N_26258);
and U29306 (N_29306,N_24131,N_24021);
or U29307 (N_29307,N_25150,N_24135);
and U29308 (N_29308,N_24268,N_26043);
nand U29309 (N_29309,N_24223,N_26582);
nor U29310 (N_29310,N_26885,N_24185);
or U29311 (N_29311,N_25010,N_24362);
and U29312 (N_29312,N_26238,N_26594);
or U29313 (N_29313,N_25637,N_25767);
nor U29314 (N_29314,N_25251,N_25466);
nor U29315 (N_29315,N_24722,N_26422);
nor U29316 (N_29316,N_24923,N_25674);
nor U29317 (N_29317,N_26635,N_25899);
and U29318 (N_29318,N_25510,N_25022);
nand U29319 (N_29319,N_25703,N_26126);
nor U29320 (N_29320,N_25091,N_24975);
and U29321 (N_29321,N_25736,N_24532);
or U29322 (N_29322,N_26942,N_24140);
xor U29323 (N_29323,N_25644,N_24326);
or U29324 (N_29324,N_24125,N_24734);
nor U29325 (N_29325,N_26205,N_24302);
and U29326 (N_29326,N_26409,N_26333);
nor U29327 (N_29327,N_24286,N_24222);
nor U29328 (N_29328,N_25888,N_26608);
nor U29329 (N_29329,N_26906,N_24219);
nand U29330 (N_29330,N_24727,N_25611);
nor U29331 (N_29331,N_26533,N_24558);
nor U29332 (N_29332,N_25853,N_26918);
and U29333 (N_29333,N_26236,N_24491);
or U29334 (N_29334,N_26274,N_26798);
nand U29335 (N_29335,N_24620,N_24063);
nand U29336 (N_29336,N_26037,N_26511);
nand U29337 (N_29337,N_26192,N_25853);
nor U29338 (N_29338,N_25005,N_26522);
nand U29339 (N_29339,N_26835,N_24574);
nand U29340 (N_29340,N_26914,N_25668);
nor U29341 (N_29341,N_26285,N_24394);
and U29342 (N_29342,N_25291,N_26749);
nor U29343 (N_29343,N_25702,N_24631);
xor U29344 (N_29344,N_26210,N_24535);
nor U29345 (N_29345,N_25622,N_26338);
xor U29346 (N_29346,N_24241,N_26460);
and U29347 (N_29347,N_24791,N_25791);
and U29348 (N_29348,N_26365,N_26959);
xor U29349 (N_29349,N_25577,N_25490);
xor U29350 (N_29350,N_24510,N_25089);
xor U29351 (N_29351,N_24134,N_25476);
or U29352 (N_29352,N_25992,N_24264);
nor U29353 (N_29353,N_25677,N_25361);
nand U29354 (N_29354,N_26264,N_24659);
nand U29355 (N_29355,N_24396,N_24868);
xnor U29356 (N_29356,N_25876,N_24298);
or U29357 (N_29357,N_26979,N_26694);
or U29358 (N_29358,N_24147,N_26082);
and U29359 (N_29359,N_24424,N_24704);
xnor U29360 (N_29360,N_24579,N_25180);
xor U29361 (N_29361,N_25964,N_24773);
nor U29362 (N_29362,N_25210,N_24582);
nand U29363 (N_29363,N_24181,N_26351);
and U29364 (N_29364,N_25005,N_26373);
nor U29365 (N_29365,N_26746,N_26474);
nand U29366 (N_29366,N_25731,N_24471);
and U29367 (N_29367,N_24699,N_26521);
nor U29368 (N_29368,N_25757,N_26027);
xor U29369 (N_29369,N_25427,N_26391);
xnor U29370 (N_29370,N_25333,N_25924);
nor U29371 (N_29371,N_26911,N_25876);
or U29372 (N_29372,N_26835,N_24067);
nand U29373 (N_29373,N_25127,N_24439);
nor U29374 (N_29374,N_26724,N_26214);
and U29375 (N_29375,N_26267,N_26992);
nor U29376 (N_29376,N_26326,N_25459);
and U29377 (N_29377,N_24301,N_24674);
nor U29378 (N_29378,N_25690,N_26648);
and U29379 (N_29379,N_26995,N_25867);
xor U29380 (N_29380,N_25514,N_26809);
and U29381 (N_29381,N_24542,N_24721);
nor U29382 (N_29382,N_24821,N_24413);
or U29383 (N_29383,N_26655,N_25692);
or U29384 (N_29384,N_26339,N_26689);
nand U29385 (N_29385,N_24936,N_25116);
or U29386 (N_29386,N_25945,N_25900);
xor U29387 (N_29387,N_24393,N_24373);
xnor U29388 (N_29388,N_24268,N_26418);
and U29389 (N_29389,N_26488,N_25213);
xnor U29390 (N_29390,N_26607,N_24088);
nor U29391 (N_29391,N_26614,N_26978);
and U29392 (N_29392,N_26109,N_24840);
and U29393 (N_29393,N_26817,N_24386);
xnor U29394 (N_29394,N_24417,N_25805);
nand U29395 (N_29395,N_26227,N_24892);
xor U29396 (N_29396,N_25718,N_26062);
or U29397 (N_29397,N_26220,N_25763);
or U29398 (N_29398,N_25546,N_26467);
xnor U29399 (N_29399,N_26274,N_26190);
nor U29400 (N_29400,N_24221,N_25821);
nor U29401 (N_29401,N_24023,N_25252);
nand U29402 (N_29402,N_25927,N_24348);
and U29403 (N_29403,N_26118,N_26623);
and U29404 (N_29404,N_26305,N_25299);
nand U29405 (N_29405,N_26436,N_25199);
xnor U29406 (N_29406,N_25327,N_25576);
nor U29407 (N_29407,N_24788,N_24750);
nand U29408 (N_29408,N_25820,N_26048);
and U29409 (N_29409,N_25267,N_25230);
nor U29410 (N_29410,N_25547,N_24933);
nor U29411 (N_29411,N_26882,N_24711);
nand U29412 (N_29412,N_24509,N_26261);
nand U29413 (N_29413,N_25193,N_24125);
or U29414 (N_29414,N_24690,N_25494);
nor U29415 (N_29415,N_24999,N_24026);
nor U29416 (N_29416,N_25954,N_26186);
xor U29417 (N_29417,N_24681,N_26735);
xor U29418 (N_29418,N_26354,N_24966);
xnor U29419 (N_29419,N_26208,N_24790);
xnor U29420 (N_29420,N_25821,N_26886);
and U29421 (N_29421,N_25691,N_26984);
and U29422 (N_29422,N_25217,N_24788);
and U29423 (N_29423,N_26921,N_25220);
xor U29424 (N_29424,N_25103,N_26784);
or U29425 (N_29425,N_26241,N_25237);
or U29426 (N_29426,N_26808,N_24054);
nor U29427 (N_29427,N_26104,N_25002);
xnor U29428 (N_29428,N_26944,N_26793);
nand U29429 (N_29429,N_26385,N_24000);
or U29430 (N_29430,N_24598,N_25107);
nor U29431 (N_29431,N_25119,N_26925);
xor U29432 (N_29432,N_25057,N_24061);
nor U29433 (N_29433,N_24585,N_24142);
nand U29434 (N_29434,N_24795,N_24127);
nand U29435 (N_29435,N_24180,N_26765);
xor U29436 (N_29436,N_25052,N_25478);
and U29437 (N_29437,N_26431,N_26228);
xnor U29438 (N_29438,N_25896,N_24464);
and U29439 (N_29439,N_25014,N_25412);
xnor U29440 (N_29440,N_24483,N_26017);
or U29441 (N_29441,N_25541,N_24582);
nor U29442 (N_29442,N_25386,N_25954);
and U29443 (N_29443,N_24355,N_24177);
xnor U29444 (N_29444,N_26460,N_25197);
nand U29445 (N_29445,N_25639,N_24192);
xor U29446 (N_29446,N_26826,N_24739);
xor U29447 (N_29447,N_26293,N_26131);
and U29448 (N_29448,N_24785,N_24156);
and U29449 (N_29449,N_26583,N_24176);
or U29450 (N_29450,N_25692,N_25891);
or U29451 (N_29451,N_25458,N_24329);
nand U29452 (N_29452,N_25412,N_26816);
nor U29453 (N_29453,N_25103,N_25156);
nand U29454 (N_29454,N_25024,N_24809);
or U29455 (N_29455,N_26425,N_25652);
and U29456 (N_29456,N_24453,N_25859);
or U29457 (N_29457,N_26341,N_26859);
nor U29458 (N_29458,N_24086,N_24238);
and U29459 (N_29459,N_24946,N_24669);
xnor U29460 (N_29460,N_26116,N_26733);
nor U29461 (N_29461,N_25533,N_26094);
or U29462 (N_29462,N_26662,N_26996);
and U29463 (N_29463,N_25724,N_26992);
or U29464 (N_29464,N_26110,N_26161);
and U29465 (N_29465,N_24330,N_24309);
or U29466 (N_29466,N_25397,N_26207);
nand U29467 (N_29467,N_24178,N_24499);
xnor U29468 (N_29468,N_26457,N_25123);
or U29469 (N_29469,N_26239,N_25916);
xnor U29470 (N_29470,N_24895,N_25752);
and U29471 (N_29471,N_24787,N_24689);
nor U29472 (N_29472,N_26289,N_26166);
nor U29473 (N_29473,N_24899,N_25969);
xnor U29474 (N_29474,N_25630,N_25186);
nor U29475 (N_29475,N_24852,N_24066);
and U29476 (N_29476,N_25007,N_25432);
xnor U29477 (N_29477,N_25077,N_24543);
nor U29478 (N_29478,N_26510,N_24299);
xor U29479 (N_29479,N_26514,N_26373);
nand U29480 (N_29480,N_25490,N_24750);
nor U29481 (N_29481,N_26059,N_26067);
nor U29482 (N_29482,N_26384,N_26075);
nor U29483 (N_29483,N_25679,N_25092);
nor U29484 (N_29484,N_24639,N_25443);
nand U29485 (N_29485,N_24742,N_25292);
xnor U29486 (N_29486,N_26445,N_25451);
xor U29487 (N_29487,N_24691,N_26006);
and U29488 (N_29488,N_24783,N_25250);
nand U29489 (N_29489,N_24541,N_24019);
xor U29490 (N_29490,N_26341,N_24172);
or U29491 (N_29491,N_24697,N_25310);
nand U29492 (N_29492,N_26188,N_26680);
and U29493 (N_29493,N_26856,N_25819);
xnor U29494 (N_29494,N_26820,N_24511);
or U29495 (N_29495,N_25134,N_24177);
xnor U29496 (N_29496,N_26466,N_25032);
and U29497 (N_29497,N_26759,N_24926);
or U29498 (N_29498,N_26925,N_24900);
nand U29499 (N_29499,N_25992,N_26936);
nand U29500 (N_29500,N_24494,N_25300);
nand U29501 (N_29501,N_26606,N_25866);
and U29502 (N_29502,N_25839,N_24408);
nor U29503 (N_29503,N_26536,N_24524);
and U29504 (N_29504,N_25127,N_24111);
nor U29505 (N_29505,N_24205,N_24519);
nor U29506 (N_29506,N_26076,N_24392);
nand U29507 (N_29507,N_24216,N_24436);
nor U29508 (N_29508,N_25906,N_25351);
or U29509 (N_29509,N_25770,N_26682);
nand U29510 (N_29510,N_25733,N_24094);
nand U29511 (N_29511,N_24734,N_26441);
xnor U29512 (N_29512,N_25160,N_25211);
xnor U29513 (N_29513,N_25036,N_24273);
nand U29514 (N_29514,N_25061,N_26070);
and U29515 (N_29515,N_26897,N_26326);
and U29516 (N_29516,N_24737,N_25027);
nor U29517 (N_29517,N_24091,N_24461);
and U29518 (N_29518,N_26196,N_24584);
xnor U29519 (N_29519,N_26601,N_24345);
nand U29520 (N_29520,N_24864,N_24208);
nor U29521 (N_29521,N_26144,N_25279);
and U29522 (N_29522,N_24946,N_26960);
nor U29523 (N_29523,N_24567,N_25997);
or U29524 (N_29524,N_24526,N_26083);
nor U29525 (N_29525,N_25072,N_24228);
or U29526 (N_29526,N_25723,N_24646);
nand U29527 (N_29527,N_26209,N_26099);
or U29528 (N_29528,N_24873,N_24592);
nand U29529 (N_29529,N_24456,N_25166);
xnor U29530 (N_29530,N_26808,N_26320);
or U29531 (N_29531,N_24494,N_25199);
and U29532 (N_29532,N_25826,N_25925);
xor U29533 (N_29533,N_24985,N_24626);
xor U29534 (N_29534,N_25488,N_26075);
xnor U29535 (N_29535,N_25284,N_25827);
nor U29536 (N_29536,N_26083,N_26912);
and U29537 (N_29537,N_24145,N_26717);
or U29538 (N_29538,N_24160,N_26137);
nand U29539 (N_29539,N_24819,N_24488);
xor U29540 (N_29540,N_25328,N_25163);
nor U29541 (N_29541,N_25390,N_25418);
nor U29542 (N_29542,N_26626,N_24698);
or U29543 (N_29543,N_25751,N_26180);
nor U29544 (N_29544,N_24137,N_26954);
or U29545 (N_29545,N_25968,N_25650);
or U29546 (N_29546,N_24738,N_26801);
xnor U29547 (N_29547,N_25325,N_26253);
or U29548 (N_29548,N_26853,N_24773);
nor U29549 (N_29549,N_24464,N_24544);
nand U29550 (N_29550,N_25960,N_26068);
xnor U29551 (N_29551,N_26129,N_25076);
and U29552 (N_29552,N_25041,N_24596);
nor U29553 (N_29553,N_26066,N_25991);
or U29554 (N_29554,N_24598,N_25392);
and U29555 (N_29555,N_26244,N_25179);
nand U29556 (N_29556,N_25689,N_26135);
nor U29557 (N_29557,N_25358,N_25330);
xor U29558 (N_29558,N_25653,N_26110);
nor U29559 (N_29559,N_25771,N_24387);
nand U29560 (N_29560,N_26113,N_26332);
and U29561 (N_29561,N_24341,N_25564);
nor U29562 (N_29562,N_25692,N_24917);
nor U29563 (N_29563,N_26824,N_24387);
xnor U29564 (N_29564,N_26711,N_25596);
and U29565 (N_29565,N_26365,N_25134);
or U29566 (N_29566,N_26184,N_25715);
xnor U29567 (N_29567,N_24019,N_25519);
nand U29568 (N_29568,N_24730,N_25201);
nand U29569 (N_29569,N_26533,N_25635);
nand U29570 (N_29570,N_26610,N_24572);
nand U29571 (N_29571,N_26823,N_25734);
nor U29572 (N_29572,N_25406,N_26447);
xnor U29573 (N_29573,N_26787,N_26070);
nand U29574 (N_29574,N_24682,N_25833);
xnor U29575 (N_29575,N_26723,N_26482);
and U29576 (N_29576,N_26016,N_26886);
nand U29577 (N_29577,N_25756,N_25562);
nor U29578 (N_29578,N_25183,N_25844);
or U29579 (N_29579,N_25324,N_25144);
xnor U29580 (N_29580,N_25426,N_24319);
nand U29581 (N_29581,N_24887,N_25421);
xor U29582 (N_29582,N_25845,N_26878);
nor U29583 (N_29583,N_24501,N_26574);
or U29584 (N_29584,N_24460,N_24278);
and U29585 (N_29585,N_26883,N_24814);
or U29586 (N_29586,N_26516,N_26229);
nor U29587 (N_29587,N_25936,N_25483);
or U29588 (N_29588,N_26872,N_25081);
xnor U29589 (N_29589,N_25475,N_26104);
nand U29590 (N_29590,N_26416,N_24142);
or U29591 (N_29591,N_25330,N_26784);
or U29592 (N_29592,N_26209,N_24447);
xor U29593 (N_29593,N_26409,N_24114);
nor U29594 (N_29594,N_25333,N_26175);
or U29595 (N_29595,N_25985,N_24749);
nand U29596 (N_29596,N_25123,N_26666);
xnor U29597 (N_29597,N_26784,N_24480);
nand U29598 (N_29598,N_25889,N_25666);
nand U29599 (N_29599,N_26269,N_24749);
xnor U29600 (N_29600,N_25313,N_26684);
nor U29601 (N_29601,N_24043,N_25883);
nor U29602 (N_29602,N_25453,N_26445);
or U29603 (N_29603,N_26052,N_25286);
nand U29604 (N_29604,N_25008,N_25018);
nand U29605 (N_29605,N_26896,N_26676);
and U29606 (N_29606,N_24660,N_26929);
nand U29607 (N_29607,N_25397,N_25102);
nor U29608 (N_29608,N_26650,N_24600);
and U29609 (N_29609,N_25212,N_25395);
xnor U29610 (N_29610,N_26635,N_25660);
nand U29611 (N_29611,N_26929,N_25991);
or U29612 (N_29612,N_26304,N_25817);
nand U29613 (N_29613,N_24880,N_24359);
xor U29614 (N_29614,N_26062,N_25963);
and U29615 (N_29615,N_24755,N_26961);
and U29616 (N_29616,N_25876,N_26292);
and U29617 (N_29617,N_25989,N_26241);
and U29618 (N_29618,N_24455,N_26174);
nand U29619 (N_29619,N_26837,N_24407);
nor U29620 (N_29620,N_26800,N_24209);
nor U29621 (N_29621,N_26093,N_26864);
xnor U29622 (N_29622,N_24789,N_25691);
and U29623 (N_29623,N_24469,N_26940);
nand U29624 (N_29624,N_25801,N_25389);
xor U29625 (N_29625,N_26729,N_24305);
and U29626 (N_29626,N_25931,N_25437);
nand U29627 (N_29627,N_25869,N_24025);
nand U29628 (N_29628,N_25959,N_26665);
and U29629 (N_29629,N_26935,N_24191);
xnor U29630 (N_29630,N_26374,N_24820);
xor U29631 (N_29631,N_24502,N_24855);
nor U29632 (N_29632,N_25351,N_24824);
and U29633 (N_29633,N_26448,N_26931);
or U29634 (N_29634,N_25990,N_24354);
nand U29635 (N_29635,N_26162,N_24231);
nor U29636 (N_29636,N_25542,N_24524);
nor U29637 (N_29637,N_25773,N_26219);
or U29638 (N_29638,N_26391,N_24460);
or U29639 (N_29639,N_26635,N_26527);
and U29640 (N_29640,N_26450,N_24795);
or U29641 (N_29641,N_24468,N_25104);
xnor U29642 (N_29642,N_25654,N_25508);
nand U29643 (N_29643,N_26478,N_24877);
xnor U29644 (N_29644,N_26439,N_25725);
nand U29645 (N_29645,N_25265,N_26852);
xnor U29646 (N_29646,N_26628,N_24311);
xnor U29647 (N_29647,N_25490,N_25544);
and U29648 (N_29648,N_26047,N_26728);
and U29649 (N_29649,N_25829,N_26144);
nor U29650 (N_29650,N_24652,N_25463);
nor U29651 (N_29651,N_24021,N_26706);
and U29652 (N_29652,N_24407,N_24649);
xnor U29653 (N_29653,N_26319,N_25654);
xnor U29654 (N_29654,N_26571,N_24158);
and U29655 (N_29655,N_24652,N_25537);
or U29656 (N_29656,N_24129,N_26284);
nand U29657 (N_29657,N_25014,N_25463);
nor U29658 (N_29658,N_26334,N_24472);
nand U29659 (N_29659,N_26620,N_25018);
nand U29660 (N_29660,N_25454,N_24215);
nand U29661 (N_29661,N_25979,N_24149);
xor U29662 (N_29662,N_24670,N_25744);
nand U29663 (N_29663,N_24635,N_25321);
xor U29664 (N_29664,N_24743,N_25859);
and U29665 (N_29665,N_24818,N_24745);
nand U29666 (N_29666,N_25510,N_25033);
and U29667 (N_29667,N_26934,N_25964);
nand U29668 (N_29668,N_24673,N_25019);
nand U29669 (N_29669,N_25703,N_24906);
nand U29670 (N_29670,N_25672,N_24407);
or U29671 (N_29671,N_24945,N_24409);
nand U29672 (N_29672,N_25775,N_25422);
xnor U29673 (N_29673,N_25107,N_24030);
nor U29674 (N_29674,N_26839,N_24428);
xor U29675 (N_29675,N_26926,N_25231);
xnor U29676 (N_29676,N_25010,N_24409);
and U29677 (N_29677,N_25029,N_25968);
or U29678 (N_29678,N_25430,N_24905);
nor U29679 (N_29679,N_26327,N_24368);
or U29680 (N_29680,N_26467,N_26081);
and U29681 (N_29681,N_26321,N_25956);
and U29682 (N_29682,N_25856,N_25105);
nor U29683 (N_29683,N_24525,N_24359);
or U29684 (N_29684,N_24668,N_24029);
nand U29685 (N_29685,N_24031,N_26594);
nor U29686 (N_29686,N_24753,N_25883);
nor U29687 (N_29687,N_24127,N_26980);
nand U29688 (N_29688,N_24164,N_25044);
and U29689 (N_29689,N_25907,N_24380);
nand U29690 (N_29690,N_26831,N_24086);
xor U29691 (N_29691,N_26794,N_24121);
and U29692 (N_29692,N_24718,N_25254);
nor U29693 (N_29693,N_26147,N_26413);
and U29694 (N_29694,N_25444,N_25200);
nor U29695 (N_29695,N_24091,N_25931);
nor U29696 (N_29696,N_24190,N_26466);
nand U29697 (N_29697,N_24098,N_24396);
nor U29698 (N_29698,N_26447,N_24638);
xnor U29699 (N_29699,N_25609,N_25323);
xor U29700 (N_29700,N_26280,N_26320);
xnor U29701 (N_29701,N_25016,N_26847);
and U29702 (N_29702,N_25041,N_26780);
nand U29703 (N_29703,N_25369,N_26182);
nand U29704 (N_29704,N_26156,N_26877);
nor U29705 (N_29705,N_25330,N_26366);
xor U29706 (N_29706,N_26193,N_25342);
and U29707 (N_29707,N_26269,N_26998);
nor U29708 (N_29708,N_24919,N_25237);
nand U29709 (N_29709,N_26297,N_26389);
nand U29710 (N_29710,N_25228,N_26004);
or U29711 (N_29711,N_24876,N_24330);
nor U29712 (N_29712,N_26909,N_25485);
and U29713 (N_29713,N_25528,N_26241);
or U29714 (N_29714,N_24853,N_26327);
and U29715 (N_29715,N_24355,N_25575);
xor U29716 (N_29716,N_24851,N_25574);
xnor U29717 (N_29717,N_25383,N_24711);
or U29718 (N_29718,N_25886,N_24196);
nand U29719 (N_29719,N_26544,N_26159);
xnor U29720 (N_29720,N_26809,N_25008);
or U29721 (N_29721,N_26336,N_26853);
or U29722 (N_29722,N_24575,N_26124);
or U29723 (N_29723,N_24982,N_26498);
nand U29724 (N_29724,N_26704,N_25903);
xor U29725 (N_29725,N_26721,N_25455);
nor U29726 (N_29726,N_24396,N_25763);
and U29727 (N_29727,N_24074,N_24025);
or U29728 (N_29728,N_25971,N_25842);
nor U29729 (N_29729,N_25983,N_26490);
nor U29730 (N_29730,N_26181,N_24929);
and U29731 (N_29731,N_26125,N_24755);
or U29732 (N_29732,N_26700,N_25889);
and U29733 (N_29733,N_25306,N_26444);
and U29734 (N_29734,N_25104,N_24999);
nor U29735 (N_29735,N_25876,N_25329);
or U29736 (N_29736,N_25879,N_25689);
and U29737 (N_29737,N_25057,N_25093);
nand U29738 (N_29738,N_26415,N_26790);
nand U29739 (N_29739,N_24726,N_26845);
or U29740 (N_29740,N_24478,N_24123);
xor U29741 (N_29741,N_24269,N_25141);
nor U29742 (N_29742,N_26008,N_25520);
xor U29743 (N_29743,N_24135,N_25980);
and U29744 (N_29744,N_25909,N_25778);
or U29745 (N_29745,N_24807,N_26419);
xor U29746 (N_29746,N_24843,N_26251);
xor U29747 (N_29747,N_26554,N_24234);
nor U29748 (N_29748,N_24892,N_25708);
or U29749 (N_29749,N_24342,N_25403);
or U29750 (N_29750,N_25094,N_24458);
and U29751 (N_29751,N_26968,N_24120);
nor U29752 (N_29752,N_24652,N_25172);
nor U29753 (N_29753,N_26392,N_24301);
or U29754 (N_29754,N_24775,N_24742);
or U29755 (N_29755,N_24927,N_25662);
nor U29756 (N_29756,N_26956,N_24418);
and U29757 (N_29757,N_26411,N_26259);
nand U29758 (N_29758,N_24796,N_25279);
xor U29759 (N_29759,N_24498,N_24373);
nand U29760 (N_29760,N_24400,N_25499);
or U29761 (N_29761,N_26332,N_24058);
nand U29762 (N_29762,N_26102,N_24505);
nand U29763 (N_29763,N_25870,N_26845);
nor U29764 (N_29764,N_26514,N_24473);
nand U29765 (N_29765,N_25895,N_25002);
nor U29766 (N_29766,N_24701,N_24103);
and U29767 (N_29767,N_24987,N_25704);
nor U29768 (N_29768,N_26555,N_25427);
and U29769 (N_29769,N_25353,N_25719);
xnor U29770 (N_29770,N_24919,N_24345);
or U29771 (N_29771,N_26530,N_25954);
xnor U29772 (N_29772,N_25239,N_24563);
nor U29773 (N_29773,N_26997,N_24213);
nand U29774 (N_29774,N_24161,N_26411);
xor U29775 (N_29775,N_24770,N_25119);
or U29776 (N_29776,N_25472,N_25254);
or U29777 (N_29777,N_26096,N_24177);
or U29778 (N_29778,N_25743,N_26057);
nor U29779 (N_29779,N_25128,N_26469);
xor U29780 (N_29780,N_26462,N_25728);
nand U29781 (N_29781,N_25630,N_25592);
or U29782 (N_29782,N_24165,N_24371);
xor U29783 (N_29783,N_24525,N_24023);
xor U29784 (N_29784,N_25868,N_25629);
or U29785 (N_29785,N_26858,N_25751);
nand U29786 (N_29786,N_26826,N_26451);
nand U29787 (N_29787,N_24772,N_24180);
nor U29788 (N_29788,N_24293,N_25102);
xnor U29789 (N_29789,N_25712,N_24369);
xor U29790 (N_29790,N_26028,N_26726);
or U29791 (N_29791,N_25200,N_24437);
and U29792 (N_29792,N_25880,N_26751);
nor U29793 (N_29793,N_26380,N_25824);
nand U29794 (N_29794,N_25105,N_25950);
nand U29795 (N_29795,N_24929,N_26862);
or U29796 (N_29796,N_24711,N_25586);
and U29797 (N_29797,N_25186,N_24471);
and U29798 (N_29798,N_25155,N_24550);
xor U29799 (N_29799,N_25617,N_25181);
nand U29800 (N_29800,N_25821,N_25621);
and U29801 (N_29801,N_25284,N_26077);
nor U29802 (N_29802,N_24718,N_24272);
and U29803 (N_29803,N_26942,N_26527);
and U29804 (N_29804,N_24118,N_26471);
nor U29805 (N_29805,N_24659,N_26414);
and U29806 (N_29806,N_26018,N_25860);
xnor U29807 (N_29807,N_26401,N_25631);
nor U29808 (N_29808,N_25633,N_24447);
or U29809 (N_29809,N_25867,N_25064);
xnor U29810 (N_29810,N_26743,N_24091);
xor U29811 (N_29811,N_24239,N_26617);
or U29812 (N_29812,N_25228,N_26462);
nor U29813 (N_29813,N_26301,N_26201);
nand U29814 (N_29814,N_25453,N_25862);
and U29815 (N_29815,N_25246,N_25222);
nand U29816 (N_29816,N_24210,N_24838);
or U29817 (N_29817,N_24557,N_25970);
and U29818 (N_29818,N_25554,N_26230);
xor U29819 (N_29819,N_24780,N_24229);
nand U29820 (N_29820,N_26581,N_26934);
xor U29821 (N_29821,N_25886,N_24508);
or U29822 (N_29822,N_25710,N_24812);
xnor U29823 (N_29823,N_24251,N_25828);
nand U29824 (N_29824,N_24509,N_25142);
nand U29825 (N_29825,N_25117,N_24241);
or U29826 (N_29826,N_24715,N_25422);
nor U29827 (N_29827,N_24380,N_24364);
xor U29828 (N_29828,N_25140,N_25162);
nor U29829 (N_29829,N_25626,N_25482);
xnor U29830 (N_29830,N_25772,N_25542);
nor U29831 (N_29831,N_25817,N_25105);
and U29832 (N_29832,N_24770,N_25528);
xnor U29833 (N_29833,N_24271,N_25459);
and U29834 (N_29834,N_24569,N_24924);
or U29835 (N_29835,N_25875,N_26211);
xor U29836 (N_29836,N_25034,N_26442);
and U29837 (N_29837,N_24441,N_25269);
nand U29838 (N_29838,N_26981,N_25949);
and U29839 (N_29839,N_26453,N_24289);
nand U29840 (N_29840,N_24358,N_24429);
nand U29841 (N_29841,N_26568,N_25856);
nand U29842 (N_29842,N_25263,N_24936);
nor U29843 (N_29843,N_26476,N_24059);
nor U29844 (N_29844,N_24411,N_24421);
and U29845 (N_29845,N_25217,N_24159);
nand U29846 (N_29846,N_24173,N_26833);
nand U29847 (N_29847,N_26396,N_24100);
or U29848 (N_29848,N_25846,N_26247);
and U29849 (N_29849,N_25390,N_25154);
nand U29850 (N_29850,N_24333,N_24339);
nand U29851 (N_29851,N_26931,N_24355);
nor U29852 (N_29852,N_26357,N_25803);
nand U29853 (N_29853,N_25111,N_24339);
or U29854 (N_29854,N_26337,N_25895);
nand U29855 (N_29855,N_26886,N_26819);
xor U29856 (N_29856,N_25082,N_24933);
nand U29857 (N_29857,N_26612,N_24718);
and U29858 (N_29858,N_26879,N_25480);
xnor U29859 (N_29859,N_24898,N_26285);
nor U29860 (N_29860,N_26491,N_25529);
nand U29861 (N_29861,N_26703,N_25717);
or U29862 (N_29862,N_25629,N_26221);
and U29863 (N_29863,N_26904,N_26402);
xnor U29864 (N_29864,N_25994,N_26508);
and U29865 (N_29865,N_25051,N_24564);
nor U29866 (N_29866,N_24747,N_25564);
and U29867 (N_29867,N_26185,N_26713);
or U29868 (N_29868,N_24409,N_26755);
nor U29869 (N_29869,N_24214,N_26006);
or U29870 (N_29870,N_24417,N_26709);
xor U29871 (N_29871,N_26174,N_25138);
xor U29872 (N_29872,N_24975,N_24737);
xor U29873 (N_29873,N_26853,N_24197);
or U29874 (N_29874,N_25421,N_24235);
or U29875 (N_29875,N_24282,N_24750);
nand U29876 (N_29876,N_25676,N_26129);
nand U29877 (N_29877,N_24434,N_25163);
nand U29878 (N_29878,N_24181,N_25899);
nor U29879 (N_29879,N_24038,N_24204);
xnor U29880 (N_29880,N_25813,N_24667);
or U29881 (N_29881,N_24161,N_24367);
or U29882 (N_29882,N_26405,N_25679);
xor U29883 (N_29883,N_24986,N_24385);
and U29884 (N_29884,N_24986,N_26155);
or U29885 (N_29885,N_25328,N_25392);
and U29886 (N_29886,N_24453,N_26689);
nor U29887 (N_29887,N_26514,N_24190);
xnor U29888 (N_29888,N_25423,N_24395);
nor U29889 (N_29889,N_26079,N_25362);
nor U29890 (N_29890,N_24746,N_24437);
and U29891 (N_29891,N_25125,N_26645);
or U29892 (N_29892,N_25547,N_26574);
or U29893 (N_29893,N_25061,N_25617);
or U29894 (N_29894,N_24067,N_24308);
and U29895 (N_29895,N_25789,N_26939);
or U29896 (N_29896,N_26109,N_24856);
nand U29897 (N_29897,N_25460,N_25687);
xnor U29898 (N_29898,N_24466,N_24191);
xor U29899 (N_29899,N_24825,N_25221);
xnor U29900 (N_29900,N_24367,N_26013);
nand U29901 (N_29901,N_26320,N_25507);
xnor U29902 (N_29902,N_25362,N_24956);
nand U29903 (N_29903,N_26538,N_25795);
and U29904 (N_29904,N_26688,N_25867);
nor U29905 (N_29905,N_25670,N_24769);
nor U29906 (N_29906,N_26263,N_25169);
nand U29907 (N_29907,N_26054,N_25826);
xor U29908 (N_29908,N_24714,N_26044);
xnor U29909 (N_29909,N_25199,N_26424);
xnor U29910 (N_29910,N_24140,N_25630);
and U29911 (N_29911,N_24621,N_25051);
nand U29912 (N_29912,N_24439,N_24050);
nor U29913 (N_29913,N_24228,N_25918);
nor U29914 (N_29914,N_25471,N_26559);
xor U29915 (N_29915,N_25952,N_24900);
and U29916 (N_29916,N_25736,N_25550);
xnor U29917 (N_29917,N_25146,N_26404);
and U29918 (N_29918,N_24029,N_24175);
and U29919 (N_29919,N_26445,N_24982);
and U29920 (N_29920,N_25737,N_25815);
nand U29921 (N_29921,N_26593,N_26690);
xor U29922 (N_29922,N_25267,N_25541);
nor U29923 (N_29923,N_24814,N_26045);
nand U29924 (N_29924,N_26940,N_25875);
and U29925 (N_29925,N_25046,N_24176);
or U29926 (N_29926,N_24444,N_26920);
and U29927 (N_29927,N_24589,N_26650);
nand U29928 (N_29928,N_25951,N_25540);
and U29929 (N_29929,N_26569,N_24273);
and U29930 (N_29930,N_24241,N_25036);
nand U29931 (N_29931,N_26308,N_26832);
and U29932 (N_29932,N_25933,N_24435);
and U29933 (N_29933,N_24432,N_25345);
or U29934 (N_29934,N_24624,N_26628);
nand U29935 (N_29935,N_26875,N_26640);
and U29936 (N_29936,N_25535,N_26064);
nand U29937 (N_29937,N_26934,N_24920);
xor U29938 (N_29938,N_25865,N_26361);
or U29939 (N_29939,N_25938,N_25369);
xor U29940 (N_29940,N_26571,N_25448);
nand U29941 (N_29941,N_26304,N_26801);
nand U29942 (N_29942,N_26858,N_26041);
and U29943 (N_29943,N_26856,N_25716);
xnor U29944 (N_29944,N_24740,N_25368);
and U29945 (N_29945,N_26989,N_26516);
nand U29946 (N_29946,N_26962,N_26318);
or U29947 (N_29947,N_24708,N_24807);
nand U29948 (N_29948,N_26228,N_26341);
nand U29949 (N_29949,N_26604,N_25344);
or U29950 (N_29950,N_25558,N_26501);
or U29951 (N_29951,N_24734,N_26119);
or U29952 (N_29952,N_24020,N_25565);
xor U29953 (N_29953,N_26555,N_24134);
xnor U29954 (N_29954,N_25658,N_25372);
xnor U29955 (N_29955,N_26873,N_24396);
nand U29956 (N_29956,N_24648,N_24974);
xnor U29957 (N_29957,N_26927,N_26230);
nor U29958 (N_29958,N_25571,N_26346);
nor U29959 (N_29959,N_24036,N_26435);
nand U29960 (N_29960,N_26948,N_26662);
and U29961 (N_29961,N_26376,N_24237);
and U29962 (N_29962,N_26861,N_26257);
or U29963 (N_29963,N_25417,N_24837);
xnor U29964 (N_29964,N_24769,N_26891);
and U29965 (N_29965,N_24154,N_24270);
xnor U29966 (N_29966,N_26615,N_25365);
xor U29967 (N_29967,N_24635,N_25824);
nand U29968 (N_29968,N_25347,N_26039);
nor U29969 (N_29969,N_25715,N_26490);
nor U29970 (N_29970,N_24434,N_26852);
or U29971 (N_29971,N_25229,N_25233);
nand U29972 (N_29972,N_26573,N_24142);
nor U29973 (N_29973,N_25297,N_24810);
or U29974 (N_29974,N_25151,N_24646);
and U29975 (N_29975,N_25226,N_24720);
nand U29976 (N_29976,N_26907,N_26726);
xor U29977 (N_29977,N_26091,N_24678);
and U29978 (N_29978,N_26508,N_24425);
nand U29979 (N_29979,N_25805,N_24851);
or U29980 (N_29980,N_24619,N_24550);
and U29981 (N_29981,N_26423,N_26378);
or U29982 (N_29982,N_24035,N_24602);
or U29983 (N_29983,N_24672,N_25947);
or U29984 (N_29984,N_25073,N_25762);
xnor U29985 (N_29985,N_24079,N_25063);
xnor U29986 (N_29986,N_25858,N_26525);
and U29987 (N_29987,N_26025,N_26500);
or U29988 (N_29988,N_26095,N_24267);
nor U29989 (N_29989,N_25217,N_26585);
xnor U29990 (N_29990,N_26429,N_26227);
or U29991 (N_29991,N_26046,N_26103);
or U29992 (N_29992,N_24506,N_26294);
xor U29993 (N_29993,N_25157,N_26075);
or U29994 (N_29994,N_26429,N_24102);
or U29995 (N_29995,N_26613,N_25657);
xor U29996 (N_29996,N_24287,N_25763);
and U29997 (N_29997,N_26559,N_24905);
or U29998 (N_29998,N_26488,N_25378);
and U29999 (N_29999,N_25563,N_26793);
and UO_0 (O_0,N_27855,N_28422);
nand UO_1 (O_1,N_27880,N_27979);
xnor UO_2 (O_2,N_28335,N_28187);
nand UO_3 (O_3,N_27126,N_28973);
nand UO_4 (O_4,N_28153,N_29294);
and UO_5 (O_5,N_27869,N_27189);
and UO_6 (O_6,N_29590,N_28084);
or UO_7 (O_7,N_28429,N_27325);
xnor UO_8 (O_8,N_28051,N_28950);
or UO_9 (O_9,N_27987,N_27616);
xor UO_10 (O_10,N_28216,N_28206);
and UO_11 (O_11,N_28538,N_27174);
nor UO_12 (O_12,N_28173,N_29463);
nor UO_13 (O_13,N_28557,N_28363);
or UO_14 (O_14,N_28552,N_28336);
and UO_15 (O_15,N_27463,N_29082);
or UO_16 (O_16,N_27974,N_29290);
xnor UO_17 (O_17,N_27814,N_29604);
or UO_18 (O_18,N_27474,N_27194);
xnor UO_19 (O_19,N_27466,N_28318);
or UO_20 (O_20,N_29796,N_28381);
nand UO_21 (O_21,N_28822,N_29882);
nor UO_22 (O_22,N_28582,N_28456);
xor UO_23 (O_23,N_27503,N_29887);
nor UO_24 (O_24,N_28971,N_27231);
xor UO_25 (O_25,N_29602,N_29824);
xnor UO_26 (O_26,N_29751,N_29659);
xnor UO_27 (O_27,N_28604,N_27227);
and UO_28 (O_28,N_27635,N_29099);
and UO_29 (O_29,N_28281,N_27796);
and UO_30 (O_30,N_28262,N_28674);
nor UO_31 (O_31,N_27274,N_28887);
or UO_32 (O_32,N_29809,N_27394);
xor UO_33 (O_33,N_28465,N_27183);
or UO_34 (O_34,N_28509,N_28221);
nor UO_35 (O_35,N_29425,N_27822);
or UO_36 (O_36,N_29398,N_28475);
or UO_37 (O_37,N_28151,N_29213);
nor UO_38 (O_38,N_29093,N_28589);
nand UO_39 (O_39,N_29741,N_28925);
nand UO_40 (O_40,N_29505,N_28022);
or UO_41 (O_41,N_27809,N_27072);
and UO_42 (O_42,N_29841,N_28614);
xor UO_43 (O_43,N_27175,N_29978);
nand UO_44 (O_44,N_28792,N_28577);
or UO_45 (O_45,N_27788,N_27592);
and UO_46 (O_46,N_27465,N_28935);
xnor UO_47 (O_47,N_29847,N_27560);
and UO_48 (O_48,N_28595,N_27576);
nor UO_49 (O_49,N_28949,N_29932);
xnor UO_50 (O_50,N_27820,N_27035);
and UO_51 (O_51,N_28389,N_29456);
xor UO_52 (O_52,N_28105,N_29064);
and UO_53 (O_53,N_29493,N_28908);
nor UO_54 (O_54,N_29601,N_27362);
nor UO_55 (O_55,N_27150,N_27190);
and UO_56 (O_56,N_29710,N_29970);
and UO_57 (O_57,N_29906,N_27352);
nor UO_58 (O_58,N_29490,N_27600);
or UO_59 (O_59,N_27654,N_27764);
or UO_60 (O_60,N_27714,N_28127);
or UO_61 (O_61,N_29790,N_28806);
and UO_62 (O_62,N_29447,N_29444);
or UO_63 (O_63,N_28823,N_28057);
nand UO_64 (O_64,N_28521,N_28612);
or UO_65 (O_65,N_28053,N_28957);
or UO_66 (O_66,N_28564,N_27455);
or UO_67 (O_67,N_27017,N_27122);
nor UO_68 (O_68,N_28341,N_28669);
and UO_69 (O_69,N_27957,N_29948);
and UO_70 (O_70,N_29016,N_29135);
or UO_71 (O_71,N_28987,N_28406);
xor UO_72 (O_72,N_28914,N_29062);
nor UO_73 (O_73,N_27490,N_29465);
and UO_74 (O_74,N_29990,N_27716);
nor UO_75 (O_75,N_27574,N_27514);
nor UO_76 (O_76,N_29524,N_29578);
nand UO_77 (O_77,N_28349,N_29791);
nand UO_78 (O_78,N_29792,N_27525);
and UO_79 (O_79,N_29944,N_28214);
nand UO_80 (O_80,N_29875,N_29512);
nand UO_81 (O_81,N_27236,N_28321);
or UO_82 (O_82,N_29794,N_28442);
nand UO_83 (O_83,N_28458,N_28631);
or UO_84 (O_84,N_27262,N_27609);
and UO_85 (O_85,N_28686,N_27830);
nor UO_86 (O_86,N_29683,N_28558);
nand UO_87 (O_87,N_27916,N_28453);
nor UO_88 (O_88,N_29739,N_29318);
nor UO_89 (O_89,N_29765,N_29316);
and UO_90 (O_90,N_27043,N_28068);
or UO_91 (O_91,N_29032,N_29283);
xor UO_92 (O_92,N_27684,N_29730);
nor UO_93 (O_93,N_27143,N_28154);
nor UO_94 (O_94,N_28506,N_27747);
nand UO_95 (O_95,N_29357,N_29542);
or UO_96 (O_96,N_28817,N_29892);
xnor UO_97 (O_97,N_28942,N_28872);
nand UO_98 (O_98,N_28625,N_27843);
or UO_99 (O_99,N_29289,N_29757);
nand UO_100 (O_100,N_29795,N_27159);
or UO_101 (O_101,N_28890,N_27518);
nor UO_102 (O_102,N_29368,N_29306);
xnor UO_103 (O_103,N_27831,N_27892);
or UO_104 (O_104,N_29565,N_27046);
or UO_105 (O_105,N_28437,N_28164);
xnor UO_106 (O_106,N_28457,N_27279);
nor UO_107 (O_107,N_29605,N_27295);
nor UO_108 (O_108,N_29558,N_27483);
and UO_109 (O_109,N_27431,N_29781);
nor UO_110 (O_110,N_29469,N_27965);
nor UO_111 (O_111,N_28947,N_29335);
nand UO_112 (O_112,N_29334,N_29185);
or UO_113 (O_113,N_28049,N_27475);
and UO_114 (O_114,N_28487,N_27137);
xor UO_115 (O_115,N_28342,N_29196);
or UO_116 (O_116,N_28292,N_29001);
and UO_117 (O_117,N_28192,N_27409);
nand UO_118 (O_118,N_27462,N_29343);
nand UO_119 (O_119,N_28072,N_29127);
and UO_120 (O_120,N_28092,N_29534);
xor UO_121 (O_121,N_27424,N_29609);
or UO_122 (O_122,N_29467,N_27778);
nor UO_123 (O_123,N_29162,N_29307);
xnor UO_124 (O_124,N_28649,N_28140);
nand UO_125 (O_125,N_28137,N_28428);
xor UO_126 (O_126,N_28114,N_27558);
nor UO_127 (O_127,N_27945,N_29347);
or UO_128 (O_128,N_27223,N_27547);
xor UO_129 (O_129,N_28383,N_28832);
nor UO_130 (O_130,N_29884,N_27550);
nand UO_131 (O_131,N_29636,N_28409);
xnor UO_132 (O_132,N_27495,N_29375);
or UO_133 (O_133,N_29551,N_27901);
nor UO_134 (O_134,N_27938,N_27149);
nor UO_135 (O_135,N_28374,N_27007);
nor UO_136 (O_136,N_27739,N_27829);
xor UO_137 (O_137,N_28998,N_27636);
nand UO_138 (O_138,N_28923,N_27339);
nor UO_139 (O_139,N_27057,N_27070);
and UO_140 (O_140,N_28377,N_29938);
nor UO_141 (O_141,N_29896,N_28673);
nor UO_142 (O_142,N_28352,N_28941);
and UO_143 (O_143,N_28619,N_27058);
or UO_144 (O_144,N_28002,N_28041);
nand UO_145 (O_145,N_27589,N_27834);
or UO_146 (O_146,N_27811,N_28853);
and UO_147 (O_147,N_29432,N_28061);
nor UO_148 (O_148,N_28955,N_29385);
nor UO_149 (O_149,N_28917,N_27508);
xor UO_150 (O_150,N_28211,N_28867);
or UO_151 (O_151,N_27594,N_27177);
xnor UO_152 (O_152,N_27204,N_29638);
or UO_153 (O_153,N_28005,N_29059);
xor UO_154 (O_154,N_29308,N_29771);
nor UO_155 (O_155,N_27498,N_27299);
nor UO_156 (O_156,N_27812,N_29296);
xnor UO_157 (O_157,N_28520,N_29759);
nor UO_158 (O_158,N_27876,N_27668);
or UO_159 (O_159,N_27675,N_29982);
and UO_160 (O_160,N_29407,N_29525);
xor UO_161 (O_161,N_27597,N_27264);
or UO_162 (O_162,N_27792,N_29243);
and UO_163 (O_163,N_27346,N_29063);
nand UO_164 (O_164,N_29876,N_27398);
or UO_165 (O_165,N_29395,N_27403);
or UO_166 (O_166,N_28497,N_27320);
xnor UO_167 (O_167,N_29428,N_28338);
nand UO_168 (O_168,N_27519,N_29483);
or UO_169 (O_169,N_29198,N_27791);
nand UO_170 (O_170,N_28358,N_27363);
xnor UO_171 (O_171,N_29777,N_28440);
nand UO_172 (O_172,N_27089,N_28616);
xor UO_173 (O_173,N_27036,N_27453);
xnor UO_174 (O_174,N_29391,N_29258);
nor UO_175 (O_175,N_27691,N_28459);
and UO_176 (O_176,N_29762,N_29802);
xor UO_177 (O_177,N_28572,N_28907);
nand UO_178 (O_178,N_28510,N_28030);
xnor UO_179 (O_179,N_29798,N_29533);
nand UO_180 (O_180,N_28020,N_28166);
or UO_181 (O_181,N_27828,N_27022);
and UO_182 (O_182,N_28545,N_29141);
or UO_183 (O_183,N_29136,N_28160);
or UO_184 (O_184,N_29509,N_29359);
or UO_185 (O_185,N_27327,N_27208);
or UO_186 (O_186,N_27765,N_29842);
nor UO_187 (O_187,N_29380,N_27507);
and UO_188 (O_188,N_28663,N_28851);
nor UO_189 (O_189,N_28985,N_28896);
and UO_190 (O_190,N_27585,N_27566);
and UO_191 (O_191,N_29203,N_28431);
nor UO_192 (O_192,N_28500,N_28136);
xor UO_193 (O_193,N_29562,N_27847);
nor UO_194 (O_194,N_29164,N_28514);
or UO_195 (O_195,N_27485,N_29550);
or UO_196 (O_196,N_27815,N_29071);
xor UO_197 (O_197,N_28085,N_27117);
or UO_198 (O_198,N_28977,N_28778);
nor UO_199 (O_199,N_29338,N_29039);
and UO_200 (O_200,N_29228,N_29439);
nand UO_201 (O_201,N_29635,N_27201);
and UO_202 (O_202,N_29251,N_27003);
xnor UO_203 (O_203,N_28253,N_29641);
and UO_204 (O_204,N_29329,N_28375);
xor UO_205 (O_205,N_27337,N_28791);
nand UO_206 (O_206,N_28074,N_29773);
nand UO_207 (O_207,N_29124,N_29173);
or UO_208 (O_208,N_29508,N_27061);
nor UO_209 (O_209,N_29580,N_29331);
or UO_210 (O_210,N_27124,N_29042);
or UO_211 (O_211,N_28567,N_28159);
nor UO_212 (O_212,N_27493,N_27782);
xor UO_213 (O_213,N_29626,N_28225);
or UO_214 (O_214,N_27021,N_28910);
nor UO_215 (O_215,N_29592,N_29879);
and UO_216 (O_216,N_27571,N_27599);
nand UO_217 (O_217,N_27048,N_27915);
xnor UO_218 (O_218,N_28800,N_29497);
nor UO_219 (O_219,N_29206,N_27094);
xnor UO_220 (O_220,N_27735,N_29891);
nor UO_221 (O_221,N_27138,N_28764);
nor UO_222 (O_222,N_27780,N_29889);
xor UO_223 (O_223,N_29713,N_28097);
or UO_224 (O_224,N_27724,N_28541);
and UO_225 (O_225,N_29914,N_27018);
xor UO_226 (O_226,N_27312,N_27596);
nor UO_227 (O_227,N_29188,N_28134);
xor UO_228 (O_228,N_27752,N_27091);
nand UO_229 (O_229,N_29917,N_28780);
or UO_230 (O_230,N_27947,N_28018);
and UO_231 (O_231,N_28812,N_28714);
xor UO_232 (O_232,N_28869,N_29890);
nor UO_233 (O_233,N_28069,N_28740);
xor UO_234 (O_234,N_28360,N_28297);
or UO_235 (O_235,N_27008,N_27435);
and UO_236 (O_236,N_29106,N_27912);
nand UO_237 (O_237,N_29256,N_28986);
xor UO_238 (O_238,N_28819,N_29121);
nor UO_239 (O_239,N_29690,N_27309);
xnor UO_240 (O_240,N_29051,N_27631);
and UO_241 (O_241,N_28592,N_28613);
nand UO_242 (O_242,N_27775,N_29210);
xor UO_243 (O_243,N_28969,N_27893);
and UO_244 (O_244,N_28718,N_29442);
nor UO_245 (O_245,N_28814,N_28331);
xor UO_246 (O_246,N_29648,N_29342);
nor UO_247 (O_247,N_29707,N_28449);
nor UO_248 (O_248,N_29653,N_27545);
nor UO_249 (O_249,N_28413,N_28676);
nand UO_250 (O_250,N_27929,N_28568);
nor UO_251 (O_251,N_27106,N_29787);
nor UO_252 (O_252,N_27064,N_29718);
nand UO_253 (O_253,N_27188,N_27981);
and UO_254 (O_254,N_29496,N_28099);
or UO_255 (O_255,N_29346,N_28280);
nor UO_256 (O_256,N_29088,N_28464);
or UO_257 (O_257,N_29764,N_28432);
nand UO_258 (O_258,N_29968,N_29133);
nand UO_259 (O_259,N_27863,N_27405);
and UO_260 (O_260,N_27578,N_28641);
or UO_261 (O_261,N_29011,N_29814);
nor UO_262 (O_262,N_28028,N_28899);
and UO_263 (O_263,N_27395,N_27364);
nand UO_264 (O_264,N_29895,N_27397);
xnor UO_265 (O_265,N_27242,N_28642);
or UO_266 (O_266,N_29284,N_29597);
nor UO_267 (O_267,N_28968,N_28007);
or UO_268 (O_268,N_29446,N_27146);
nand UO_269 (O_269,N_28016,N_27185);
or UO_270 (O_270,N_27696,N_28855);
xnor UO_271 (O_271,N_29817,N_27891);
nor UO_272 (O_272,N_28761,N_27639);
nor UO_273 (O_273,N_27345,N_28001);
or UO_274 (O_274,N_27492,N_27410);
xor UO_275 (O_275,N_29214,N_27013);
or UO_276 (O_276,N_27034,N_29293);
nand UO_277 (O_277,N_28524,N_27854);
or UO_278 (O_278,N_28461,N_29390);
nor UO_279 (O_279,N_29721,N_27155);
nor UO_280 (O_280,N_29725,N_28943);
and UO_281 (O_281,N_27727,N_28738);
nand UO_282 (O_282,N_27818,N_27224);
nand UO_283 (O_283,N_29285,N_28646);
and UO_284 (O_284,N_28039,N_28043);
and UO_285 (O_285,N_29888,N_28798);
nand UO_286 (O_286,N_27538,N_29547);
and UO_287 (O_287,N_29504,N_27567);
or UO_288 (O_288,N_29367,N_27206);
and UO_289 (O_289,N_29231,N_28783);
nand UO_290 (O_290,N_29409,N_28760);
xnor UO_291 (O_291,N_29235,N_28387);
xor UO_292 (O_292,N_29129,N_29441);
nor UO_293 (O_293,N_28197,N_28285);
or UO_294 (O_294,N_27548,N_28893);
nand UO_295 (O_295,N_29351,N_28199);
nor UO_296 (O_296,N_29568,N_28665);
nor UO_297 (O_297,N_29176,N_29652);
nor UO_298 (O_298,N_27484,N_27428);
nand UO_299 (O_299,N_27993,N_27569);
nor UO_300 (O_300,N_28838,N_28593);
nand UO_301 (O_301,N_28622,N_27321);
or UO_302 (O_302,N_27918,N_28742);
xor UO_303 (O_303,N_27877,N_27099);
or UO_304 (O_304,N_29157,N_27120);
nand UO_305 (O_305,N_29820,N_27991);
nand UO_306 (O_306,N_27366,N_29072);
and UO_307 (O_307,N_27167,N_29950);
xor UO_308 (O_308,N_29557,N_28366);
nor UO_309 (O_309,N_29302,N_27010);
xor UO_310 (O_310,N_27068,N_29193);
nor UO_311 (O_311,N_27249,N_29860);
nand UO_312 (O_312,N_28438,N_28999);
or UO_313 (O_313,N_29480,N_28198);
and UO_314 (O_314,N_29159,N_27510);
nand UO_315 (O_315,N_29386,N_29946);
nand UO_316 (O_316,N_27667,N_28873);
nand UO_317 (O_317,N_29170,N_27817);
xor UO_318 (O_318,N_28630,N_27549);
xnor UO_319 (O_319,N_28797,N_29478);
and UO_320 (O_320,N_28145,N_27479);
and UO_321 (O_321,N_28484,N_29705);
nand UO_322 (O_322,N_28547,N_29190);
and UO_323 (O_323,N_29957,N_27128);
nor UO_324 (O_324,N_27618,N_27874);
xnor UO_325 (O_325,N_29819,N_27865);
or UO_326 (O_326,N_28540,N_28570);
or UO_327 (O_327,N_28130,N_29411);
or UO_328 (O_328,N_28073,N_27878);
or UO_329 (O_329,N_28975,N_27628);
nand UO_330 (O_330,N_29598,N_29988);
xor UO_331 (O_331,N_29865,N_28284);
xor UO_332 (O_332,N_27731,N_29680);
or UO_333 (O_333,N_28444,N_29614);
xor UO_334 (O_334,N_27723,N_27678);
nand UO_335 (O_335,N_28116,N_27688);
nand UO_336 (O_336,N_27433,N_29619);
nor UO_337 (O_337,N_27999,N_29309);
xnor UO_338 (O_338,N_28010,N_29920);
nor UO_339 (O_339,N_27743,N_29315);
nor UO_340 (O_340,N_28122,N_28433);
or UO_341 (O_341,N_29100,N_28208);
or UO_342 (O_342,N_28393,N_28576);
xor UO_343 (O_343,N_28584,N_27712);
or UO_344 (O_344,N_28905,N_29528);
and UO_345 (O_345,N_27709,N_28109);
nor UO_346 (O_346,N_29564,N_29918);
nor UO_347 (O_347,N_28356,N_29736);
and UO_348 (O_348,N_28201,N_27084);
nor UO_349 (O_349,N_29225,N_27996);
nor UO_350 (O_350,N_27166,N_29181);
nor UO_351 (O_351,N_29953,N_27838);
and UO_352 (O_352,N_29958,N_28242);
xor UO_353 (O_353,N_29379,N_27319);
nor UO_354 (O_354,N_27305,N_27728);
or UO_355 (O_355,N_28060,N_27041);
or UO_356 (O_356,N_28367,N_27740);
and UO_357 (O_357,N_27448,N_28378);
xor UO_358 (O_358,N_29234,N_29273);
nor UO_359 (O_359,N_28729,N_29056);
and UO_360 (O_360,N_28255,N_28322);
and UO_361 (O_361,N_27645,N_29134);
or UO_362 (O_362,N_27973,N_29731);
xor UO_363 (O_363,N_27537,N_27357);
nand UO_364 (O_364,N_28274,N_29947);
or UO_365 (O_365,N_29142,N_27436);
nor UO_366 (O_366,N_28106,N_27808);
nand UO_367 (O_367,N_28055,N_27643);
and UO_368 (O_368,N_27954,N_27109);
nand UO_369 (O_369,N_29049,N_28291);
xnor UO_370 (O_370,N_29069,N_27480);
nor UO_371 (O_371,N_28699,N_28499);
nor UO_372 (O_372,N_27162,N_28328);
and UO_373 (O_373,N_27977,N_27079);
nand UO_374 (O_374,N_27533,N_29007);
and UO_375 (O_375,N_28289,N_27706);
and UO_376 (O_376,N_29660,N_29595);
nand UO_377 (O_377,N_28959,N_28410);
xnor UO_378 (O_378,N_28194,N_29570);
nor UO_379 (O_379,N_28997,N_28082);
nand UO_380 (O_380,N_28648,N_28989);
or UO_381 (O_381,N_28048,N_27750);
nand UO_382 (O_382,N_29855,N_27807);
and UO_383 (O_383,N_27404,N_27681);
nor UO_384 (O_384,N_27887,N_29433);
and UO_385 (O_385,N_28575,N_27280);
and UO_386 (O_386,N_28306,N_28354);
and UO_387 (O_387,N_27603,N_27470);
xor UO_388 (O_388,N_28024,N_29146);
or UO_389 (O_389,N_29111,N_27238);
xnor UO_390 (O_390,N_27927,N_29928);
and UO_391 (O_391,N_29934,N_29327);
xnor UO_392 (O_392,N_28156,N_29826);
or UO_393 (O_393,N_27130,N_27145);
nor UO_394 (O_394,N_28270,N_29963);
and UO_395 (O_395,N_29406,N_28228);
or UO_396 (O_396,N_28861,N_27456);
or UO_397 (O_397,N_28139,N_29555);
nand UO_398 (O_398,N_28587,N_27897);
or UO_399 (O_399,N_28035,N_28310);
nand UO_400 (O_400,N_29460,N_28209);
nor UO_401 (O_401,N_29054,N_28118);
nand UO_402 (O_402,N_29232,N_28725);
nor UO_403 (O_403,N_29576,N_27434);
xnor UO_404 (O_404,N_28301,N_28561);
and UO_405 (O_405,N_29734,N_28585);
and UO_406 (O_406,N_28566,N_29872);
nand UO_407 (O_407,N_29085,N_27575);
xnor UO_408 (O_408,N_29607,N_29147);
nor UO_409 (O_409,N_27350,N_27252);
and UO_410 (O_410,N_29581,N_27193);
nand UO_411 (O_411,N_28535,N_27923);
nor UO_412 (O_412,N_29837,N_27388);
and UO_413 (O_413,N_29022,N_28300);
nor UO_414 (O_414,N_29749,N_27922);
or UO_415 (O_415,N_29935,N_29077);
nand UO_416 (O_416,N_28878,N_29215);
nand UO_417 (O_417,N_28235,N_28277);
nand UO_418 (O_418,N_28532,N_27982);
xnor UO_419 (O_419,N_27755,N_29271);
and UO_420 (O_420,N_28357,N_29114);
nand UO_421 (O_421,N_29748,N_27420);
or UO_422 (O_422,N_29588,N_27445);
and UO_423 (O_423,N_27284,N_28003);
or UO_424 (O_424,N_28848,N_27920);
nand UO_425 (O_425,N_27650,N_29009);
and UO_426 (O_426,N_29663,N_27692);
nand UO_427 (O_427,N_28758,N_28064);
xnor UO_428 (O_428,N_28189,N_29171);
and UO_429 (O_429,N_28371,N_28994);
xnor UO_430 (O_430,N_29221,N_27367);
and UO_431 (O_431,N_29599,N_28078);
or UO_432 (O_432,N_27400,N_29012);
and UO_433 (O_433,N_28058,N_27802);
and UO_434 (O_434,N_27827,N_27263);
or UO_435 (O_435,N_27486,N_28799);
and UO_436 (O_436,N_27777,N_27073);
nor UO_437 (O_437,N_27859,N_28750);
or UO_438 (O_438,N_28183,N_28835);
xor UO_439 (O_439,N_27411,N_29924);
and UO_440 (O_440,N_27103,N_29037);
nand UO_441 (O_441,N_28144,N_28477);
nor UO_442 (O_442,N_27531,N_27816);
nor UO_443 (O_443,N_28675,N_28793);
nor UO_444 (O_444,N_29167,N_27179);
xor UO_445 (O_445,N_28621,N_29040);
xnor UO_446 (O_446,N_28709,N_28922);
and UO_447 (O_447,N_29295,N_29584);
nor UO_448 (O_448,N_27332,N_29417);
xnor UO_449 (O_449,N_29627,N_27783);
xnor UO_450 (O_450,N_29515,N_27399);
xnor UO_451 (O_451,N_29254,N_28844);
nand UO_452 (O_452,N_27027,N_27077);
and UO_453 (O_453,N_29322,N_28653);
xor UO_454 (O_454,N_29416,N_27972);
nand UO_455 (O_455,N_28617,N_29745);
nand UO_456 (O_456,N_28390,N_28528);
or UO_457 (O_457,N_27211,N_29628);
and UO_458 (O_458,N_28932,N_28483);
nor UO_459 (O_459,N_28644,N_29518);
nand UO_460 (O_460,N_27568,N_29211);
nand UO_461 (O_461,N_28876,N_28385);
or UO_462 (O_462,N_29392,N_29337);
xnor UO_463 (O_463,N_27590,N_29775);
nor UO_464 (O_464,N_28830,N_29929);
nand UO_465 (O_465,N_27302,N_29028);
or UO_466 (O_466,N_28207,N_27303);
and UO_467 (O_467,N_28370,N_28239);
xnor UO_468 (O_468,N_27506,N_29219);
and UO_469 (O_469,N_28185,N_27255);
nand UO_470 (O_470,N_27736,N_27734);
xor UO_471 (O_471,N_27232,N_27666);
nand UO_472 (O_472,N_29615,N_29191);
nand UO_473 (O_473,N_29204,N_28178);
and UO_474 (O_474,N_28781,N_29816);
nand UO_475 (O_475,N_27772,N_27552);
nor UO_476 (O_476,N_27200,N_28278);
xor UO_477 (O_477,N_29014,N_29989);
or UO_478 (O_478,N_29836,N_29959);
nor UO_479 (O_479,N_29361,N_29424);
nand UO_480 (O_480,N_29931,N_28809);
nor UO_481 (O_481,N_27000,N_29669);
xnor UO_482 (O_482,N_29856,N_28480);
or UO_483 (O_483,N_27660,N_29276);
xnor UO_484 (O_484,N_27115,N_28895);
and UO_485 (O_485,N_28293,N_27665);
and UO_486 (O_486,N_29087,N_29073);
nand UO_487 (O_487,N_28681,N_27697);
xor UO_488 (O_488,N_27835,N_27195);
xnor UO_489 (O_489,N_29596,N_27541);
or UO_490 (O_490,N_28113,N_28288);
nand UO_491 (O_491,N_28845,N_29864);
or UO_492 (O_492,N_28021,N_29153);
or UO_493 (O_493,N_27413,N_28737);
and UO_494 (O_494,N_29649,N_27761);
nor UO_495 (O_495,N_27119,N_28143);
and UO_496 (O_496,N_27649,N_28450);
or UO_497 (O_497,N_29760,N_29259);
and UO_498 (O_498,N_27317,N_29697);
xor UO_499 (O_499,N_28150,N_29637);
nand UO_500 (O_500,N_27924,N_28610);
nand UO_501 (O_501,N_27862,N_27459);
or UO_502 (O_502,N_27412,N_29706);
nor UO_503 (O_503,N_29647,N_28694);
and UO_504 (O_504,N_29332,N_28327);
xor UO_505 (O_505,N_28337,N_27886);
xor UO_506 (O_506,N_29319,N_29954);
xor UO_507 (O_507,N_28933,N_28004);
and UO_508 (O_508,N_29616,N_28515);
nand UO_509 (O_509,N_27156,N_28254);
nand UO_510 (O_510,N_27801,N_28672);
and UO_511 (O_511,N_29236,N_27088);
and UO_512 (O_512,N_27447,N_28287);
and UO_513 (O_513,N_29940,N_29152);
or UO_514 (O_514,N_28779,N_27451);
nor UO_515 (O_515,N_28807,N_28243);
nor UO_516 (O_516,N_28379,N_28972);
nor UO_517 (O_517,N_28571,N_27781);
xnor UO_518 (O_518,N_28888,N_29880);
nor UO_519 (O_519,N_28634,N_29843);
nand UO_520 (O_520,N_29101,N_27423);
nand UO_521 (O_521,N_29536,N_29247);
or UO_522 (O_522,N_29827,N_29930);
nor UO_523 (O_523,N_29571,N_27160);
or UO_524 (O_524,N_29737,N_28530);
and UO_525 (O_525,N_29326,N_27066);
xnor UO_526 (O_526,N_28019,N_27396);
xor UO_527 (O_527,N_28754,N_28990);
nor UO_528 (O_528,N_28081,N_29898);
nand UO_529 (O_529,N_27970,N_29182);
xor UO_530 (O_530,N_29374,N_29901);
or UO_531 (O_531,N_28948,N_27360);
or UO_532 (O_532,N_28701,N_29716);
and UO_533 (O_533,N_29255,N_29603);
nor UO_534 (O_534,N_29224,N_27819);
nor UO_535 (O_535,N_29109,N_29067);
and UO_536 (O_536,N_27113,N_29674);
and UO_537 (O_537,N_28931,N_29092);
or UO_538 (O_538,N_27006,N_29569);
nor UO_539 (O_539,N_28656,N_28875);
and UO_540 (O_540,N_28924,N_28227);
and UO_541 (O_541,N_27943,N_28298);
nand UO_542 (O_542,N_28014,N_28219);
and UO_543 (O_543,N_28915,N_28944);
and UO_544 (O_544,N_29105,N_28494);
or UO_545 (O_545,N_28495,N_28596);
nand UO_546 (O_546,N_29464,N_29418);
nor UO_547 (O_547,N_28871,N_28025);
or UO_548 (O_548,N_29404,N_27478);
or UO_549 (O_549,N_29498,N_29832);
and UO_550 (O_550,N_29662,N_29268);
nor UO_551 (O_551,N_27546,N_27062);
or UO_552 (O_552,N_27326,N_29358);
or UO_553 (O_553,N_27803,N_28573);
or UO_554 (O_554,N_29753,N_28463);
nand UO_555 (O_555,N_27852,N_27906);
nand UO_556 (O_556,N_27329,N_29178);
or UO_557 (O_557,N_28044,N_27646);
or UO_558 (O_558,N_29986,N_29500);
nand UO_559 (O_559,N_27960,N_29297);
and UO_560 (O_560,N_28544,N_27429);
or UO_561 (O_561,N_29560,N_27392);
xnor UO_562 (O_562,N_28874,N_27257);
nor UO_563 (O_563,N_28498,N_28650);
and UO_564 (O_564,N_28346,N_27521);
and UO_565 (O_565,N_28045,N_27577);
nand UO_566 (O_566,N_28751,N_27215);
and UO_567 (O_567,N_28307,N_29727);
nand UO_568 (O_568,N_29369,N_28067);
xor UO_569 (O_569,N_28726,N_27873);
or UO_570 (O_570,N_28283,N_27297);
and UO_571 (O_571,N_28857,N_28279);
xnor UO_572 (O_572,N_28042,N_29853);
or UO_573 (O_573,N_29878,N_27349);
xnor UO_574 (O_574,N_29844,N_28347);
or UO_575 (O_575,N_27967,N_28089);
or UO_576 (O_576,N_28785,N_28258);
nand UO_577 (O_577,N_29752,N_27657);
and UO_578 (O_578,N_29086,N_29511);
nand UO_579 (O_579,N_28898,N_29320);
nor UO_580 (O_580,N_29722,N_28103);
xnor UO_581 (O_581,N_29102,N_27213);
nor UO_582 (O_582,N_29549,N_29382);
xnor UO_583 (O_583,N_28926,N_27375);
and UO_584 (O_584,N_28687,N_27151);
nand UO_585 (O_585,N_28056,N_28756);
or UO_586 (O_586,N_28963,N_28420);
or UO_587 (O_587,N_27677,N_28138);
or UO_588 (O_588,N_29671,N_28316);
nand UO_589 (O_589,N_27144,N_29961);
or UO_590 (O_590,N_29070,N_29743);
and UO_591 (O_591,N_28423,N_29645);
xnor UO_592 (O_592,N_27343,N_29066);
and UO_593 (O_593,N_29554,N_28901);
or UO_594 (O_594,N_27551,N_29941);
xor UO_595 (O_595,N_28640,N_28107);
xnor UO_596 (O_596,N_27347,N_27028);
and UO_597 (O_597,N_29212,N_27340);
and UO_598 (O_598,N_27795,N_27438);
nor UO_599 (O_599,N_29695,N_28938);
xor UO_600 (O_600,N_27842,N_28482);
xnor UO_601 (O_601,N_28286,N_27686);
or UO_602 (O_602,N_29624,N_28868);
nor UO_603 (O_603,N_29150,N_28353);
xor UO_604 (O_604,N_27306,N_28152);
xor UO_605 (O_605,N_28195,N_27528);
xor UO_606 (O_606,N_27700,N_28174);
xor UO_607 (O_607,N_27276,N_27254);
or UO_608 (O_608,N_29241,N_27198);
nor UO_609 (O_609,N_28079,N_29983);
nor UO_610 (O_610,N_27365,N_28493);
or UO_611 (O_611,N_28680,N_27080);
xor UO_612 (O_612,N_28664,N_29119);
or UO_613 (O_613,N_27563,N_27376);
nor UO_614 (O_614,N_27882,N_27037);
nand UO_615 (O_615,N_27024,N_29089);
and UO_616 (O_616,N_27093,N_28268);
and UO_617 (O_617,N_27172,N_27373);
nand UO_618 (O_618,N_27333,N_29027);
nand UO_619 (O_619,N_27919,N_27427);
nor UO_620 (O_620,N_29199,N_28565);
nand UO_621 (O_621,N_27372,N_27625);
xor UO_622 (O_622,N_29384,N_27648);
nor UO_623 (O_623,N_27212,N_29854);
xor UO_624 (O_624,N_28351,N_28607);
nor UO_625 (O_625,N_29149,N_28369);
nand UO_626 (O_626,N_28569,N_29195);
nor UO_627 (O_627,N_29378,N_28682);
nor UO_628 (O_628,N_27572,N_27670);
nand UO_629 (O_629,N_27142,N_29910);
nand UO_630 (O_630,N_27038,N_29955);
xor UO_631 (O_631,N_27270,N_27861);
nor UO_632 (O_632,N_28047,N_27836);
and UO_633 (O_633,N_28344,N_27173);
nand UO_634 (O_634,N_29783,N_27380);
nand UO_635 (O_635,N_27233,N_27621);
or UO_636 (O_636,N_29481,N_27002);
or UO_637 (O_637,N_29838,N_27440);
and UO_638 (O_638,N_29942,N_29328);
nand UO_639 (O_639,N_28101,N_28992);
nand UO_640 (O_640,N_27751,N_27065);
or UO_641 (O_641,N_27244,N_27019);
nand UO_642 (O_642,N_29415,N_28556);
nor UO_643 (O_643,N_29026,N_28364);
xnor UO_644 (O_644,N_27307,N_29813);
nand UO_645 (O_645,N_29714,N_28919);
and UO_646 (O_646,N_28157,N_29393);
and UO_647 (O_647,N_29679,N_28802);
xor UO_648 (O_648,N_29699,N_27135);
nand UO_649 (O_649,N_28418,N_27417);
or UO_650 (O_650,N_29926,N_28606);
xor UO_651 (O_651,N_29263,N_27356);
nand UO_652 (O_652,N_29161,N_28479);
xnor UO_653 (O_653,N_28412,N_28334);
and UO_654 (O_654,N_28952,N_27557);
and UO_655 (O_655,N_27497,N_27132);
and UO_656 (O_656,N_28692,N_28794);
or UO_657 (O_657,N_27180,N_27769);
nor UO_658 (O_658,N_28244,N_29443);
nand UO_659 (O_659,N_29519,N_28359);
and UO_660 (O_660,N_27182,N_27797);
xor UO_661 (O_661,N_29956,N_28993);
and UO_662 (O_662,N_28052,N_28745);
xnor UO_663 (O_663,N_28980,N_29353);
or UO_664 (O_664,N_29981,N_27799);
nor UO_665 (O_665,N_29107,N_27932);
xor UO_666 (O_666,N_27586,N_29644);
xnor UO_667 (O_667,N_29687,N_29482);
xnor UO_668 (O_668,N_27757,N_28320);
xnor UO_669 (O_669,N_28722,N_28401);
xnor UO_670 (O_670,N_29006,N_28600);
nor UO_671 (O_671,N_29726,N_29815);
nand UO_672 (O_672,N_27701,N_29700);
and UO_673 (O_673,N_27905,N_28065);
nor UO_674 (O_674,N_29692,N_28711);
nand UO_675 (O_675,N_27237,N_28323);
or UO_676 (O_676,N_27604,N_28533);
nand UO_677 (O_677,N_29915,N_29396);
nor UO_678 (O_678,N_27903,N_29470);
nor UO_679 (O_679,N_28721,N_29080);
xnor UO_680 (O_680,N_29996,N_28825);
xor UO_681 (O_681,N_28936,N_28141);
or UO_682 (O_682,N_29747,N_29510);
nand UO_683 (O_683,N_27632,N_27216);
xnor UO_684 (O_684,N_29381,N_29506);
xnor UO_685 (O_685,N_28771,N_29230);
xor UO_686 (O_686,N_27230,N_29998);
and UO_687 (O_687,N_27766,N_27591);
and UO_688 (O_688,N_29646,N_29279);
xor UO_689 (O_689,N_28891,N_27464);
nand UO_690 (O_690,N_29462,N_28314);
nand UO_691 (O_691,N_28077,N_28266);
or UO_692 (O_692,N_29115,N_27259);
nor UO_693 (O_693,N_29689,N_28330);
and UO_694 (O_694,N_27529,N_29402);
nor UO_695 (O_695,N_28038,N_27371);
xor UO_696 (O_696,N_29189,N_29421);
nand UO_697 (O_697,N_28679,N_29702);
and UO_698 (O_698,N_29613,N_27939);
and UO_699 (O_699,N_28441,N_29905);
and UO_700 (O_700,N_28503,N_28609);
xnor UO_701 (O_701,N_28847,N_29967);
or UO_702 (O_702,N_28471,N_29282);
and UO_703 (O_703,N_27239,N_29436);
nand UO_704 (O_704,N_29048,N_28504);
or UO_705 (O_705,N_29239,N_28961);
nor UO_706 (O_706,N_29656,N_28176);
and UO_707 (O_707,N_27821,N_29767);
xnor UO_708 (O_708,N_27853,N_27023);
nand UO_709 (O_709,N_29197,N_28094);
xor UO_710 (O_710,N_27832,N_29237);
nand UO_711 (O_711,N_29526,N_29186);
nor UO_712 (O_712,N_28264,N_29287);
and UO_713 (O_713,N_28117,N_27687);
and UO_714 (O_714,N_28251,N_28637);
nand UO_715 (O_715,N_27672,N_27205);
and UO_716 (O_716,N_28615,N_28488);
or UO_717 (O_717,N_27899,N_27271);
xnor UO_718 (O_718,N_27437,N_29194);
nand UO_719 (O_719,N_27860,N_29449);
nand UO_720 (O_720,N_29720,N_29240);
xnor UO_721 (O_721,N_28815,N_29991);
and UO_722 (O_722,N_29420,N_27060);
nand UO_723 (O_723,N_27102,N_27348);
xnor UO_724 (O_724,N_27773,N_29175);
nor UO_725 (O_725,N_28840,N_29352);
xnor UO_726 (O_726,N_29354,N_28583);
and UO_727 (O_727,N_27745,N_28034);
nor UO_728 (O_728,N_27989,N_27994);
nand UO_729 (O_729,N_29589,N_28704);
nand UO_730 (O_730,N_27473,N_28996);
nand UO_731 (O_731,N_28563,N_27118);
nand UO_732 (O_732,N_29894,N_29728);
xnor UO_733 (O_733,N_29657,N_27784);
nand UO_734 (O_734,N_28636,N_27148);
or UO_735 (O_735,N_28626,N_28215);
nand UO_736 (O_736,N_27730,N_29805);
xor UO_737 (O_737,N_28525,N_29611);
nor UO_738 (O_738,N_29522,N_28690);
nor UO_739 (O_739,N_27491,N_28424);
and UO_740 (O_740,N_27512,N_27526);
nor UO_741 (O_741,N_27588,N_28708);
nor UO_742 (O_742,N_27914,N_27315);
or UO_743 (O_743,N_28193,N_28960);
xnor UO_744 (O_744,N_29431,N_29413);
and UO_745 (O_745,N_27898,N_27642);
nand UO_746 (O_746,N_29750,N_29020);
xnor UO_747 (O_747,N_27564,N_29774);
nand UO_748 (O_748,N_28309,N_29266);
xnor UO_749 (O_749,N_28661,N_28267);
or UO_750 (O_750,N_29499,N_29015);
nor UO_751 (O_751,N_28885,N_28502);
or UO_752 (O_752,N_28599,N_28180);
nor UO_753 (O_753,N_28365,N_27653);
nor UO_754 (O_754,N_27140,N_29793);
xor UO_755 (O_755,N_28093,N_27718);
xor UO_756 (O_756,N_29997,N_29172);
xor UO_757 (O_757,N_29013,N_29365);
xnor UO_758 (O_758,N_27573,N_27457);
nand UO_759 (O_759,N_28693,N_29539);
nor UO_760 (O_760,N_29587,N_27948);
or UO_761 (O_761,N_28689,N_27275);
or UO_762 (O_762,N_27840,N_29846);
or UO_763 (O_763,N_27744,N_27226);
nor UO_764 (O_764,N_27944,N_27097);
and UO_765 (O_765,N_29103,N_27983);
and UO_766 (O_766,N_28902,N_29301);
nand UO_767 (O_767,N_27133,N_28516);
or UO_768 (O_768,N_29494,N_28315);
or UO_769 (O_769,N_27516,N_28303);
and UO_770 (O_770,N_28852,N_27199);
nor UO_771 (O_771,N_29041,N_27582);
or UO_772 (O_772,N_28033,N_27934);
xnor UO_773 (O_773,N_27833,N_29050);
and UO_774 (O_774,N_28308,N_28531);
nand UO_775 (O_775,N_29985,N_28404);
xor UO_776 (O_776,N_28982,N_27620);
nand UO_777 (O_777,N_28181,N_29123);
nand UO_778 (O_778,N_29691,N_29448);
nand UO_779 (O_779,N_27925,N_28128);
or UO_780 (O_780,N_28467,N_29631);
or UO_781 (O_781,N_28037,N_27704);
xnor UO_782 (O_782,N_27517,N_27968);
xor UO_783 (O_783,N_28829,N_27505);
and UO_784 (O_784,N_29873,N_29098);
nand UO_785 (O_785,N_28177,N_29964);
nand UO_786 (O_786,N_28304,N_27310);
nand UO_787 (O_787,N_29921,N_28376);
and UO_788 (O_788,N_27441,N_29625);
or UO_789 (O_789,N_27884,N_28755);
or UO_790 (O_790,N_27896,N_29693);
xor UO_791 (O_791,N_27785,N_28324);
and UO_792 (O_792,N_27634,N_27504);
nand UO_793 (O_793,N_28485,N_29643);
and UO_794 (O_794,N_28313,N_27004);
xnor UO_795 (O_795,N_29476,N_28850);
xnor UO_796 (O_796,N_27674,N_29005);
or UO_797 (O_797,N_28408,N_29632);
and UO_798 (O_798,N_28169,N_27361);
nand UO_799 (O_799,N_27015,N_29874);
nand UO_800 (O_800,N_29746,N_28131);
and UO_801 (O_801,N_27178,N_27472);
xnor UO_802 (O_802,N_29845,N_29076);
nand UO_803 (O_803,N_29586,N_28833);
nor UO_804 (O_804,N_28396,N_28719);
or UO_805 (O_805,N_27846,N_29292);
nor UO_806 (O_806,N_28854,N_28723);
nor UO_807 (O_807,N_27662,N_27753);
or UO_808 (O_808,N_29140,N_27288);
xnor UO_809 (O_809,N_27956,N_29538);
nand UO_810 (O_810,N_27902,N_29912);
xor UO_811 (O_811,N_28731,N_27131);
or UO_812 (O_812,N_27656,N_29772);
nand UO_813 (O_813,N_28965,N_29561);
xnor UO_814 (O_814,N_28611,N_29514);
xor UO_815 (O_815,N_29937,N_29227);
nand UO_816 (O_816,N_27881,N_27894);
nand UO_817 (O_817,N_29169,N_28883);
or UO_818 (O_818,N_28527,N_28749);
xnor UO_819 (O_819,N_29763,N_28115);
or UO_820 (O_820,N_27680,N_29274);
or UO_821 (O_821,N_29818,N_28032);
nor UO_822 (O_822,N_27690,N_28548);
or UO_823 (O_823,N_28230,N_29992);
or UO_824 (O_824,N_29936,N_29949);
nand UO_825 (O_825,N_27153,N_29804);
and UO_826 (O_826,N_29620,N_28311);
nand UO_827 (O_827,N_28678,N_27936);
xor UO_828 (O_828,N_29806,N_27168);
nor UO_829 (O_829,N_27287,N_27565);
nor UO_830 (O_830,N_28302,N_27341);
or UO_831 (O_831,N_29517,N_29715);
xnor UO_832 (O_832,N_29678,N_28759);
or UO_833 (O_833,N_29249,N_27837);
or UO_834 (O_834,N_28647,N_28362);
xnor UO_835 (O_835,N_28210,N_28537);
and UO_836 (O_836,N_28712,N_27240);
nand UO_837 (O_837,N_28000,N_27432);
nor UO_838 (O_838,N_28928,N_29364);
or UO_839 (O_839,N_27532,N_28299);
xor UO_840 (O_840,N_28511,N_28862);
or UO_841 (O_841,N_27300,N_27539);
nor UO_842 (O_842,N_29900,N_28172);
xnor UO_843 (O_843,N_28087,N_29502);
or UO_844 (O_844,N_28076,N_28818);
and UO_845 (O_845,N_29002,N_27952);
nand UO_846 (O_846,N_28350,N_28015);
nand UO_847 (O_847,N_29866,N_29546);
xor UO_848 (O_848,N_28911,N_29466);
xor UO_849 (O_849,N_28953,N_27487);
or UO_850 (O_850,N_28981,N_27221);
nand UO_851 (O_851,N_27849,N_29553);
or UO_852 (O_852,N_27078,N_28200);
nor UO_853 (O_853,N_29556,N_27047);
nor UO_854 (O_854,N_29952,N_27689);
nand UO_855 (O_855,N_27793,N_28730);
nand UO_856 (O_856,N_28772,N_29630);
xnor UO_857 (O_857,N_27241,N_27556);
xnor UO_858 (O_858,N_28090,N_27823);
nor UO_859 (O_859,N_29582,N_28474);
nand UO_860 (O_860,N_27962,N_29719);
or UO_861 (O_861,N_27351,N_29812);
nor UO_862 (O_862,N_29345,N_28695);
xnor UO_863 (O_863,N_28163,N_28720);
and UO_864 (O_864,N_27866,N_29811);
xor UO_865 (O_865,N_28108,N_29733);
or UO_866 (O_866,N_27489,N_29744);
xor UO_867 (O_867,N_29083,N_28744);
nor UO_868 (O_868,N_27086,N_27978);
or UO_869 (O_869,N_29640,N_29664);
or UO_870 (O_870,N_27502,N_29084);
nor UO_871 (O_871,N_27071,N_28667);
or UO_872 (O_872,N_28294,N_27917);
nand UO_873 (O_873,N_27454,N_27946);
or UO_874 (O_874,N_29665,N_29363);
nor UO_875 (O_875,N_28446,N_27087);
nand UO_876 (O_876,N_27051,N_27116);
nand UO_877 (O_877,N_29673,N_29886);
or UO_878 (O_878,N_27900,N_27014);
nand UO_879 (O_879,N_28123,N_29999);
xor UO_880 (O_880,N_27527,N_28080);
or UO_881 (O_881,N_29366,N_27553);
nor UO_882 (O_882,N_29160,N_28290);
and UO_883 (O_883,N_27318,N_28560);
xnor UO_884 (O_884,N_29377,N_29701);
nand UO_885 (O_885,N_28008,N_27850);
xor UO_886 (O_886,N_29238,N_28513);
xor UO_887 (O_887,N_27449,N_29971);
nor UO_888 (O_888,N_29330,N_27170);
or UO_889 (O_889,N_27813,N_27031);
or UO_890 (O_890,N_29870,N_27655);
nor UO_891 (O_891,N_27540,N_29491);
and UO_892 (O_892,N_29972,N_29681);
xnor UO_893 (O_893,N_27872,N_27075);
and UO_894 (O_894,N_28234,N_28762);
or UO_895 (O_895,N_28826,N_28843);
nand UO_896 (O_896,N_28380,N_27110);
nand UO_897 (O_897,N_29623,N_28202);
nor UO_898 (O_898,N_28391,N_27415);
xor UO_899 (O_899,N_28063,N_27595);
nand UO_900 (O_900,N_29312,N_27738);
nand UO_901 (O_901,N_28436,N_29995);
nand UO_902 (O_902,N_28752,N_27513);
or UO_903 (O_903,N_29144,N_29047);
xor UO_904 (O_904,N_27386,N_29471);
xnor UO_905 (O_905,N_28810,N_29711);
nor UO_906 (O_906,N_28550,N_29053);
nor UO_907 (O_907,N_29766,N_29000);
xor UO_908 (O_908,N_27076,N_28715);
xor UO_909 (O_909,N_27955,N_27895);
nor UO_910 (O_910,N_27930,N_28940);
nand UO_911 (O_911,N_27370,N_28734);
or UO_912 (O_912,N_29537,N_27052);
and UO_913 (O_913,N_27841,N_28426);
and UO_914 (O_914,N_28241,N_29810);
and UO_915 (O_915,N_29246,N_28702);
nand UO_916 (O_916,N_28858,N_27063);
or UO_917 (O_917,N_29849,N_27251);
or UO_918 (O_918,N_29113,N_27971);
xor UO_919 (O_919,N_29229,N_28361);
nand UO_920 (O_920,N_28578,N_29321);
nor UO_921 (O_921,N_27406,N_27669);
xor UO_922 (O_922,N_28269,N_29125);
nand UO_923 (O_923,N_29139,N_27544);
or UO_924 (O_924,N_27127,N_29994);
nor UO_925 (O_925,N_28562,N_27617);
xnor UO_926 (O_926,N_27450,N_28884);
nand UO_927 (O_927,N_29021,N_28448);
xnor UO_928 (O_928,N_29226,N_28392);
nor UO_929 (O_929,N_28605,N_28624);
xor UO_930 (O_930,N_27598,N_28317);
xor UO_931 (O_931,N_27460,N_28031);
nor UO_932 (O_932,N_29387,N_29184);
or UO_933 (O_933,N_27385,N_28075);
or UO_934 (O_934,N_28594,N_29797);
xor UO_935 (O_935,N_29857,N_27703);
xor UO_936 (O_936,N_29675,N_27439);
and UO_937 (O_937,N_29291,N_29606);
or UO_938 (O_938,N_28158,N_27858);
nor UO_939 (O_939,N_29486,N_29907);
and UO_940 (O_940,N_29755,N_27904);
and UO_941 (O_941,N_29676,N_29852);
and UO_942 (O_942,N_29911,N_28706);
and UO_943 (O_943,N_29323,N_29388);
xor UO_944 (O_944,N_28824,N_28223);
or UO_945 (O_945,N_28939,N_29200);
nand UO_946 (O_946,N_27344,N_28329);
or UO_947 (O_947,N_28691,N_28135);
xor UO_948 (O_948,N_27209,N_27105);
or UO_949 (O_949,N_28951,N_29137);
and UO_950 (O_950,N_27272,N_28472);
or UO_951 (O_951,N_28340,N_27191);
or UO_952 (O_952,N_28892,N_28703);
xor UO_953 (O_953,N_28273,N_27638);
or UO_954 (O_954,N_29769,N_29724);
nand UO_955 (O_955,N_27005,N_27452);
nand UO_956 (O_956,N_29939,N_28276);
xor UO_957 (O_957,N_29403,N_28618);
and UO_958 (O_958,N_27384,N_28017);
nor UO_959 (O_959,N_29487,N_29801);
nand UO_960 (O_960,N_29729,N_28407);
nand UO_961 (O_961,N_29610,N_27786);
xor UO_962 (O_962,N_29858,N_29394);
nand UO_963 (O_963,N_28382,N_28546);
or UO_964 (O_964,N_29097,N_28343);
nand UO_965 (O_965,N_27311,N_28816);
nor UO_966 (O_966,N_27085,N_29541);
nand UO_967 (O_967,N_27418,N_28534);
xor UO_968 (O_968,N_28237,N_28421);
and UO_969 (O_969,N_28132,N_29712);
nand UO_970 (O_970,N_29350,N_28713);
nor UO_971 (O_971,N_28086,N_27698);
xnor UO_972 (O_972,N_27986,N_27520);
or UO_973 (O_973,N_27268,N_29848);
or UO_974 (O_974,N_27111,N_27157);
xnor UO_975 (O_975,N_28782,N_27468);
xor UO_976 (O_976,N_27839,N_28491);
or UO_977 (O_977,N_27767,N_29183);
and UO_978 (O_978,N_28275,N_27482);
or UO_979 (O_979,N_27611,N_28226);
and UO_980 (O_980,N_28542,N_28769);
nor UO_981 (O_981,N_29600,N_29303);
nand UO_982 (O_982,N_27787,N_29267);
and UO_983 (O_983,N_27067,N_29242);
or UO_984 (O_984,N_28395,N_27746);
xor UO_985 (O_985,N_28054,N_29577);
nor UO_986 (O_986,N_29723,N_29341);
nor UO_987 (O_987,N_28629,N_29822);
or UO_988 (O_988,N_27296,N_29429);
nor UO_989 (O_989,N_29356,N_27651);
nand UO_990 (O_990,N_28104,N_27641);
nor UO_991 (O_991,N_27682,N_29435);
xnor UO_992 (O_992,N_28549,N_28419);
nor UO_993 (O_993,N_29023,N_29566);
nand UO_994 (O_994,N_28768,N_27250);
or UO_995 (O_995,N_29672,N_29148);
and UO_996 (O_996,N_28966,N_27419);
nor UO_997 (O_997,N_28434,N_27658);
xor UO_998 (O_998,N_29943,N_29126);
xor UO_999 (O_999,N_27806,N_29808);
and UO_1000 (O_1000,N_27933,N_28125);
and UO_1001 (O_1001,N_27401,N_28733);
nand UO_1002 (O_1002,N_27581,N_29220);
xnor UO_1003 (O_1003,N_28828,N_27602);
and UO_1004 (O_1004,N_27269,N_28655);
nor UO_1005 (O_1005,N_29179,N_27579);
xnor UO_1006 (O_1006,N_27134,N_29548);
and UO_1007 (O_1007,N_29575,N_29192);
xor UO_1008 (O_1008,N_29400,N_28906);
nor UO_1009 (O_1009,N_27379,N_28581);
and UO_1010 (O_1010,N_29233,N_29800);
or UO_1011 (O_1011,N_29264,N_27107);
nor UO_1012 (O_1012,N_28995,N_28543);
nor UO_1013 (O_1013,N_27100,N_27708);
and UO_1014 (O_1014,N_27218,N_29807);
nand UO_1015 (O_1015,N_28222,N_29010);
nand UO_1016 (O_1016,N_29452,N_28455);
nor UO_1017 (O_1017,N_28405,N_27256);
or UO_1018 (O_1018,N_28231,N_28247);
nor UO_1019 (O_1019,N_29974,N_27011);
nor UO_1020 (O_1020,N_29789,N_27121);
and UO_1021 (O_1021,N_27054,N_28523);
nand UO_1022 (O_1022,N_27779,N_28705);
xor UO_1023 (O_1023,N_27030,N_28945);
nor UO_1024 (O_1024,N_28260,N_27220);
or UO_1025 (O_1025,N_28657,N_29567);
xnor UO_1026 (O_1026,N_27147,N_28635);
xnor UO_1027 (O_1027,N_27614,N_29029);
and UO_1028 (O_1028,N_28023,N_29180);
xnor UO_1029 (O_1029,N_27535,N_29572);
xnor UO_1030 (O_1030,N_27615,N_29655);
nor UO_1031 (O_1031,N_28466,N_28555);
or UO_1032 (O_1032,N_29430,N_27848);
nor UO_1033 (O_1033,N_28930,N_27733);
nor UO_1034 (O_1034,N_28789,N_28462);
xor UO_1035 (O_1035,N_29017,N_27805);
xor UO_1036 (O_1036,N_29018,N_29768);
nor UO_1037 (O_1037,N_28149,N_27857);
xor UO_1038 (O_1038,N_27713,N_27314);
nor UO_1039 (O_1039,N_27381,N_29883);
and UO_1040 (O_1040,N_28095,N_28179);
and UO_1041 (O_1041,N_27074,N_28481);
and UO_1042 (O_1042,N_29654,N_27378);
or UO_1043 (O_1043,N_27219,N_27984);
nor UO_1044 (O_1044,N_28168,N_28238);
or UO_1045 (O_1045,N_27940,N_29916);
or UO_1046 (O_1046,N_27258,N_28191);
or UO_1047 (O_1047,N_27243,N_27158);
or UO_1048 (O_1048,N_27969,N_28111);
nor UO_1049 (O_1049,N_29698,N_27950);
or UO_1050 (O_1050,N_29272,N_27580);
nand UO_1051 (O_1051,N_28059,N_28439);
nand UO_1052 (O_1052,N_27217,N_28688);
nor UO_1053 (O_1053,N_27444,N_29438);
or UO_1054 (O_1054,N_27608,N_29046);
xnor UO_1055 (O_1055,N_28512,N_27112);
xor UO_1056 (O_1056,N_29209,N_28696);
or UO_1057 (O_1057,N_28454,N_27707);
xor UO_1058 (O_1058,N_27584,N_28909);
xnor UO_1059 (O_1059,N_29658,N_27033);
and UO_1060 (O_1060,N_28598,N_27039);
xor UO_1061 (O_1061,N_29075,N_27096);
xnor UO_1062 (O_1062,N_27511,N_28220);
or UO_1063 (O_1063,N_27210,N_29980);
xnor UO_1064 (O_1064,N_29052,N_28724);
nand UO_1065 (O_1065,N_27702,N_29453);
nand UO_1066 (O_1066,N_29168,N_29742);
and UO_1067 (O_1067,N_28880,N_27020);
nand UO_1068 (O_1068,N_29440,N_27559);
xnor UO_1069 (O_1069,N_29280,N_29034);
or UO_1070 (O_1070,N_28813,N_28345);
or UO_1071 (O_1071,N_28245,N_29617);
nor UO_1072 (O_1072,N_27494,N_27016);
and UO_1073 (O_1073,N_28962,N_27496);
xor UO_1074 (O_1074,N_29507,N_27998);
and UO_1075 (O_1075,N_27322,N_29684);
nor UO_1076 (O_1076,N_27671,N_27711);
nand UO_1077 (O_1077,N_29543,N_28536);
nor UO_1078 (O_1078,N_29851,N_29666);
and UO_1079 (O_1079,N_29732,N_28796);
or UO_1080 (O_1080,N_29399,N_27699);
nor UO_1081 (O_1081,N_29573,N_28050);
and UO_1082 (O_1082,N_29217,N_28476);
and UO_1083 (O_1083,N_27937,N_27368);
or UO_1084 (O_1084,N_27601,N_28881);
and UO_1085 (O_1085,N_29112,N_28677);
nand UO_1086 (O_1086,N_27387,N_28171);
nor UO_1087 (O_1087,N_28388,N_28903);
nor UO_1088 (O_1088,N_27587,N_29138);
nand UO_1089 (O_1089,N_29340,N_27235);
nor UO_1090 (O_1090,N_28246,N_28517);
nor UO_1091 (O_1091,N_27909,N_27393);
nor UO_1092 (O_1092,N_28743,N_29779);
xnor UO_1093 (O_1093,N_29629,N_29840);
xor UO_1094 (O_1094,N_28460,N_29419);
nand UO_1095 (O_1095,N_27095,N_27710);
and UO_1096 (O_1096,N_28766,N_28062);
nor UO_1097 (O_1097,N_27804,N_28217);
or UO_1098 (O_1098,N_28508,N_27961);
and UO_1099 (O_1099,N_28282,N_28811);
or UO_1100 (O_1100,N_28196,N_28490);
nand UO_1101 (O_1101,N_29738,N_29520);
xor UO_1102 (O_1102,N_28305,N_29313);
xor UO_1103 (O_1103,N_27369,N_28684);
nor UO_1104 (O_1104,N_28639,N_29530);
nand UO_1105 (O_1105,N_27055,N_28747);
nand UO_1106 (O_1106,N_28697,N_29608);
nand UO_1107 (O_1107,N_29893,N_27214);
or UO_1108 (O_1108,N_28451,N_27184);
and UO_1109 (O_1109,N_29154,N_29612);
nand UO_1110 (O_1110,N_27389,N_29299);
nor UO_1111 (O_1111,N_29158,N_29786);
xnor UO_1112 (O_1112,N_27661,N_28820);
and UO_1113 (O_1113,N_28846,N_29965);
nor UO_1114 (O_1114,N_27953,N_27695);
xnor UO_1115 (O_1115,N_27561,N_29445);
or UO_1116 (O_1116,N_28271,N_29776);
and UO_1117 (O_1117,N_28601,N_27253);
xor UO_1118 (O_1118,N_29594,N_29559);
nor UO_1119 (O_1119,N_29074,N_29155);
nand UO_1120 (O_1120,N_27098,N_27633);
and UO_1121 (O_1121,N_27629,N_28040);
nand UO_1122 (O_1122,N_27042,N_27910);
or UO_1123 (O_1123,N_28492,N_27324);
and UO_1124 (O_1124,N_28518,N_28889);
or UO_1125 (O_1125,N_28836,N_27338);
or UO_1126 (O_1126,N_27885,N_27870);
nor UO_1127 (O_1127,N_28232,N_29975);
xnor UO_1128 (O_1128,N_28551,N_29861);
nor UO_1129 (O_1129,N_29278,N_28333);
or UO_1130 (O_1130,N_28190,N_28805);
or UO_1131 (O_1131,N_29523,N_28397);
xor UO_1132 (O_1132,N_29128,N_29208);
nand UO_1133 (O_1133,N_29038,N_28098);
nor UO_1134 (O_1134,N_27619,N_28859);
nor UO_1135 (O_1135,N_28553,N_27798);
or UO_1136 (O_1136,N_29685,N_28579);
xnor UO_1137 (O_1137,N_28580,N_29951);
and UO_1138 (O_1138,N_27081,N_29833);
nand UO_1139 (O_1139,N_29788,N_29945);
or UO_1140 (O_1140,N_28671,N_27606);
or UO_1141 (O_1141,N_27583,N_27562);
xor UO_1142 (O_1142,N_27754,N_29835);
or UO_1143 (O_1143,N_28927,N_29222);
or UO_1144 (O_1144,N_27719,N_28013);
or UO_1145 (O_1145,N_28027,N_27958);
nor UO_1146 (O_1146,N_29130,N_29275);
nand UO_1147 (O_1147,N_29925,N_28148);
and UO_1148 (O_1148,N_28224,N_29869);
and UO_1149 (O_1149,N_29682,N_28100);
nand UO_1150 (O_1150,N_28918,N_29281);
and UO_1151 (O_1151,N_27500,N_28700);
nand UO_1152 (O_1152,N_28735,N_27053);
xnor UO_1153 (O_1153,N_29650,N_29250);
and UO_1154 (O_1154,N_27685,N_27613);
xor UO_1155 (O_1155,N_27292,N_29410);
and UO_1156 (O_1156,N_27050,N_28124);
nor UO_1157 (O_1157,N_29055,N_29223);
or UO_1158 (O_1158,N_27390,N_28312);
xnor UO_1159 (O_1159,N_28620,N_28841);
and UO_1160 (O_1160,N_28319,N_27012);
and UO_1161 (O_1161,N_27247,N_28877);
nor UO_1162 (O_1162,N_27794,N_27992);
or UO_1163 (O_1163,N_28112,N_29244);
and UO_1164 (O_1164,N_29834,N_27790);
nand UO_1165 (O_1165,N_28597,N_28866);
nand UO_1166 (O_1166,N_28654,N_27673);
or UO_1167 (O_1167,N_28958,N_27964);
nor UO_1168 (O_1168,N_28970,N_27637);
nand UO_1169 (O_1169,N_27825,N_29455);
nor UO_1170 (O_1170,N_28628,N_28175);
nand UO_1171 (O_1171,N_27009,N_27607);
and UO_1172 (O_1172,N_29305,N_28519);
nand UO_1173 (O_1173,N_29535,N_28775);
xor UO_1174 (O_1174,N_29993,N_27358);
and UO_1175 (O_1175,N_28250,N_27985);
and UO_1176 (O_1176,N_28643,N_29008);
nor UO_1177 (O_1177,N_28856,N_27308);
xor UO_1178 (O_1178,N_27291,N_28736);
and UO_1179 (O_1179,N_27756,N_29688);
or UO_1180 (O_1180,N_29579,N_29516);
or UO_1181 (O_1181,N_29686,N_28662);
and UO_1182 (O_1182,N_28717,N_28588);
xnor UO_1183 (O_1183,N_27542,N_28976);
nand UO_1184 (O_1184,N_27921,N_29831);
or UO_1185 (O_1185,N_29899,N_29317);
and UO_1186 (O_1186,N_28256,N_27139);
nor UO_1187 (O_1187,N_28205,N_29253);
or UO_1188 (O_1188,N_29881,N_28332);
nand UO_1189 (O_1189,N_28870,N_28496);
nand UO_1190 (O_1190,N_29373,N_27328);
or UO_1191 (O_1191,N_27391,N_27114);
or UO_1192 (O_1192,N_29922,N_27044);
or UO_1193 (O_1193,N_29333,N_27298);
xor UO_1194 (O_1194,N_28710,N_29068);
nor UO_1195 (O_1195,N_28916,N_29877);
or UO_1196 (O_1196,N_27335,N_27748);
or UO_1197 (O_1197,N_28658,N_27593);
nand UO_1198 (O_1198,N_27261,N_29405);
nor UO_1199 (O_1199,N_28608,N_29091);
nand UO_1200 (O_1200,N_28821,N_27725);
xnor UO_1201 (O_1201,N_28988,N_28897);
xnor UO_1202 (O_1202,N_28767,N_29120);
xnor UO_1203 (O_1203,N_28133,N_28670);
and UO_1204 (O_1204,N_29108,N_27679);
nor UO_1205 (O_1205,N_29044,N_27377);
and UO_1206 (O_1206,N_27092,N_29670);
nor UO_1207 (O_1207,N_27851,N_29043);
or UO_1208 (O_1208,N_29708,N_27421);
nor UO_1209 (O_1209,N_28006,N_27267);
xor UO_1210 (O_1210,N_27408,N_28739);
or UO_1211 (O_1211,N_27029,N_28526);
nand UO_1212 (O_1212,N_29458,N_28120);
nand UO_1213 (O_1213,N_27323,N_27186);
nor UO_1214 (O_1214,N_28501,N_29252);
or UO_1215 (O_1215,N_28071,N_28469);
nand UO_1216 (O_1216,N_28348,N_29094);
nor UO_1217 (O_1217,N_28529,N_28842);
or UO_1218 (O_1218,N_29336,N_29145);
nand UO_1219 (O_1219,N_27331,N_28801);
nor UO_1220 (O_1220,N_27069,N_27488);
xnor UO_1221 (O_1221,N_28394,N_29492);
or UO_1222 (O_1222,N_29202,N_29218);
xor UO_1223 (O_1223,N_28204,N_29165);
nor UO_1224 (O_1224,N_27304,N_29850);
or UO_1225 (O_1225,N_27890,N_27467);
xnor UO_1226 (O_1226,N_29372,N_27382);
nand UO_1227 (O_1227,N_28913,N_28757);
xnor UO_1228 (O_1228,N_28803,N_27313);
nand UO_1229 (O_1229,N_29205,N_28746);
and UO_1230 (O_1230,N_28083,N_28325);
nor UO_1231 (O_1231,N_28026,N_27800);
and UO_1232 (O_1232,N_29717,N_27975);
or UO_1233 (O_1233,N_28632,N_29633);
nand UO_1234 (O_1234,N_27129,N_28091);
and UO_1235 (O_1235,N_27026,N_27762);
or UO_1236 (O_1236,N_27443,N_28574);
xor UO_1237 (O_1237,N_28505,N_27768);
nand UO_1238 (O_1238,N_27402,N_29003);
or UO_1239 (O_1239,N_28727,N_27245);
xor UO_1240 (O_1240,N_27963,N_28430);
and UO_1241 (O_1241,N_28070,N_27336);
nand UO_1242 (O_1242,N_27741,N_28946);
nor UO_1243 (O_1243,N_27383,N_27845);
or UO_1244 (O_1244,N_29859,N_28295);
xnor UO_1245 (O_1245,N_28770,N_28400);
nand UO_1246 (O_1246,N_29132,N_29756);
nand UO_1247 (O_1247,N_29245,N_27760);
nand UO_1248 (O_1248,N_28170,N_28146);
nor UO_1249 (O_1249,N_29667,N_29969);
and UO_1250 (O_1250,N_27676,N_28468);
or UO_1251 (O_1251,N_28920,N_28339);
nand UO_1252 (O_1252,N_29110,N_29163);
xor UO_1253 (O_1253,N_29030,N_29261);
xnor UO_1254 (O_1254,N_29116,N_29058);
and UO_1255 (O_1255,N_27187,N_28904);
nand UO_1256 (O_1256,N_27524,N_29585);
or UO_1257 (O_1257,N_29862,N_28425);
or UO_1258 (O_1258,N_29735,N_28184);
nor UO_1259 (O_1259,N_29593,N_28929);
and UO_1260 (O_1260,N_27913,N_27995);
xor UO_1261 (O_1261,N_28403,N_29437);
or UO_1262 (O_1262,N_28886,N_27980);
and UO_1263 (O_1263,N_29348,N_28954);
and UO_1264 (O_1264,N_28590,N_27523);
and UO_1265 (O_1265,N_27045,N_27515);
nand UO_1266 (O_1266,N_28233,N_28559);
or UO_1267 (O_1267,N_27108,N_29839);
and UO_1268 (O_1268,N_28659,N_29288);
or UO_1269 (O_1269,N_29909,N_27889);
nor UO_1270 (O_1270,N_28402,N_27059);
and UO_1271 (O_1271,N_29187,N_28435);
nor UO_1272 (O_1272,N_27824,N_28834);
or UO_1273 (O_1273,N_29785,N_27286);
xor UO_1274 (O_1274,N_29057,N_29639);
or UO_1275 (O_1275,N_27202,N_28763);
or UO_1276 (O_1276,N_29122,N_29545);
or UO_1277 (O_1277,N_27001,N_29269);
xnor UO_1278 (O_1278,N_28129,N_27171);
xor UO_1279 (O_1279,N_29422,N_27203);
nor UO_1280 (O_1280,N_27826,N_29355);
xor UO_1281 (O_1281,N_29475,N_28046);
nand UO_1282 (O_1282,N_29304,N_29216);
nand UO_1283 (O_1283,N_27623,N_27630);
or UO_1284 (O_1284,N_28252,N_28698);
nor UO_1285 (O_1285,N_28539,N_29799);
or UO_1286 (O_1286,N_27090,N_27407);
nor UO_1287 (O_1287,N_28265,N_29201);
nor UO_1288 (O_1288,N_27951,N_29019);
xnor UO_1289 (O_1289,N_28102,N_28119);
nor UO_1290 (O_1290,N_27988,N_29095);
and UO_1291 (O_1291,N_27720,N_29529);
nand UO_1292 (O_1292,N_28165,N_29495);
nor UO_1293 (O_1293,N_28864,N_29661);
xnor UO_1294 (O_1294,N_29065,N_29489);
nand UO_1295 (O_1295,N_28478,N_27737);
xor UO_1296 (O_1296,N_28257,N_29260);
or UO_1297 (O_1297,N_27867,N_28964);
xor UO_1298 (O_1298,N_28623,N_29310);
and UO_1299 (O_1299,N_29025,N_27471);
and UO_1300 (O_1300,N_27141,N_27871);
nand UO_1301 (O_1301,N_27770,N_27425);
or UO_1302 (O_1302,N_28249,N_27659);
nor UO_1303 (O_1303,N_27683,N_27290);
and UO_1304 (O_1304,N_27422,N_28373);
and UO_1305 (O_1305,N_29521,N_27942);
or UO_1306 (O_1306,N_28921,N_28707);
nand UO_1307 (O_1307,N_29923,N_27330);
and UO_1308 (O_1308,N_27907,N_29897);
and UO_1309 (O_1309,N_28638,N_28066);
nand UO_1310 (O_1310,N_29457,N_29574);
or UO_1311 (O_1311,N_29060,N_27868);
nor UO_1312 (O_1312,N_28991,N_28956);
xnor UO_1313 (O_1313,N_28967,N_28355);
xor UO_1314 (O_1314,N_29540,N_27626);
xor UO_1315 (O_1315,N_27293,N_27931);
nor UO_1316 (O_1316,N_29642,N_28808);
xnor UO_1317 (O_1317,N_29709,N_27941);
xnor UO_1318 (O_1318,N_27446,N_27759);
xnor UO_1319 (O_1319,N_27844,N_29829);
xor UO_1320 (O_1320,N_28384,N_28795);
or UO_1321 (O_1321,N_27749,N_28666);
nand UO_1322 (O_1322,N_27458,N_28240);
nand UO_1323 (O_1323,N_27949,N_28627);
or UO_1324 (O_1324,N_27083,N_27197);
and UO_1325 (O_1325,N_29973,N_28096);
and UO_1326 (O_1326,N_27509,N_28447);
xnor UO_1327 (O_1327,N_29913,N_28900);
nand UO_1328 (O_1328,N_29544,N_29286);
xor UO_1329 (O_1329,N_29311,N_29434);
nand UO_1330 (O_1330,N_27248,N_27196);
or UO_1331 (O_1331,N_29459,N_29503);
nand UO_1332 (O_1332,N_29166,N_29552);
nand UO_1333 (O_1333,N_28602,N_29151);
nor UO_1334 (O_1334,N_27265,N_29962);
nor UO_1335 (O_1335,N_29414,N_29033);
and UO_1336 (O_1336,N_29118,N_29265);
nand UO_1337 (O_1337,N_28186,N_27353);
or UO_1338 (O_1338,N_27136,N_27705);
nand UO_1339 (O_1339,N_29618,N_27928);
xor UO_1340 (O_1340,N_27430,N_28784);
nor UO_1341 (O_1341,N_29031,N_28765);
or UO_1342 (O_1342,N_27354,N_29371);
and UO_1343 (O_1343,N_28728,N_29668);
xnor UO_1344 (O_1344,N_27163,N_29677);
and UO_1345 (O_1345,N_28776,N_29344);
and UO_1346 (O_1346,N_29401,N_27281);
nand UO_1347 (O_1347,N_29821,N_29427);
nand UO_1348 (O_1348,N_28121,N_28860);
xnor UO_1349 (O_1349,N_29477,N_27888);
nand UO_1350 (O_1350,N_28212,N_29484);
or UO_1351 (O_1351,N_28651,N_27192);
nand UO_1352 (O_1352,N_29412,N_29376);
nand UO_1353 (O_1353,N_28011,N_29339);
xor UO_1354 (O_1354,N_29257,N_28263);
xor UO_1355 (O_1355,N_29927,N_29325);
xnor UO_1356 (O_1356,N_28147,N_27334);
nand UO_1357 (O_1357,N_28865,N_27875);
and UO_1358 (O_1358,N_29174,N_29314);
xnor UO_1359 (O_1359,N_27664,N_28788);
or UO_1360 (O_1360,N_28603,N_28879);
nor UO_1361 (O_1361,N_29454,N_29061);
nor UO_1362 (O_1362,N_27911,N_28182);
nor UO_1363 (O_1363,N_28741,N_28236);
nor UO_1364 (O_1364,N_27997,N_27610);
nand UO_1365 (O_1365,N_29761,N_27554);
xor UO_1366 (O_1366,N_27294,N_29976);
nor UO_1367 (O_1367,N_28417,N_27416);
or UO_1368 (O_1368,N_29527,N_28934);
and UO_1369 (O_1369,N_28894,N_27477);
and UO_1370 (O_1370,N_29904,N_28586);
nand UO_1371 (O_1371,N_29977,N_28009);
and UO_1372 (O_1372,N_28372,N_28668);
xnor UO_1373 (O_1373,N_28411,N_28984);
nor UO_1374 (O_1374,N_29979,N_27273);
xor UO_1375 (O_1375,N_29324,N_28162);
or UO_1376 (O_1376,N_29468,N_29583);
and UO_1377 (O_1377,N_28507,N_28660);
xor UO_1378 (O_1378,N_28774,N_28029);
nor UO_1379 (O_1379,N_29563,N_29960);
nand UO_1380 (O_1380,N_29362,N_29651);
and UO_1381 (O_1381,N_27693,N_27176);
xnor UO_1382 (O_1382,N_28683,N_27810);
or UO_1383 (O_1383,N_27729,N_28445);
and UO_1384 (O_1384,N_28645,N_29867);
and UO_1385 (O_1385,N_27316,N_29622);
xnor UO_1386 (O_1386,N_27025,N_28473);
nor UO_1387 (O_1387,N_27879,N_29177);
nor UO_1388 (O_1388,N_29621,N_27722);
nand UO_1389 (O_1389,N_28790,N_27990);
and UO_1390 (O_1390,N_29488,N_29863);
nor UO_1391 (O_1391,N_29513,N_27164);
and UO_1392 (O_1392,N_27152,N_27246);
and UO_1393 (O_1393,N_28452,N_28161);
and UO_1394 (O_1394,N_27663,N_27222);
xnor UO_1395 (O_1395,N_29248,N_27082);
nand UO_1396 (O_1396,N_29803,N_27161);
nor UO_1397 (O_1397,N_27260,N_27789);
nor UO_1398 (O_1398,N_27461,N_27481);
and UO_1399 (O_1399,N_29828,N_29045);
or UO_1400 (O_1400,N_29408,N_28974);
and UO_1401 (O_1401,N_28837,N_29987);
nand UO_1402 (O_1402,N_28978,N_28229);
nand UO_1403 (O_1403,N_29383,N_28489);
and UO_1404 (O_1404,N_29984,N_28155);
and UO_1405 (O_1405,N_29902,N_27374);
or UO_1406 (O_1406,N_27742,N_27154);
and UO_1407 (O_1407,N_27555,N_27926);
xor UO_1408 (O_1408,N_29143,N_28036);
xnor UO_1409 (O_1409,N_28261,N_28591);
nor UO_1410 (O_1410,N_27732,N_29871);
nor UO_1411 (O_1411,N_27605,N_29778);
or UO_1412 (O_1412,N_29825,N_27627);
nor UO_1413 (O_1413,N_27721,N_27976);
nor UO_1414 (O_1414,N_27414,N_27125);
nor UO_1415 (O_1415,N_27266,N_29397);
xnor UO_1416 (O_1416,N_27234,N_27530);
and UO_1417 (O_1417,N_28716,N_29501);
nor UO_1418 (O_1418,N_29479,N_29298);
or UO_1419 (O_1419,N_29036,N_27225);
xnor UO_1420 (O_1420,N_27543,N_27908);
xor UO_1421 (O_1421,N_27049,N_28470);
xnor UO_1422 (O_1422,N_27570,N_29090);
nor UO_1423 (O_1423,N_27040,N_29300);
xor UO_1424 (O_1424,N_27935,N_27123);
nor UO_1425 (O_1425,N_29830,N_29754);
and UO_1426 (O_1426,N_29696,N_28386);
xor UO_1427 (O_1427,N_29704,N_27289);
or UO_1428 (O_1428,N_27522,N_27104);
nor UO_1429 (O_1429,N_27442,N_28753);
and UO_1430 (O_1430,N_28110,N_29885);
and UO_1431 (O_1431,N_28685,N_28486);
or UO_1432 (O_1432,N_29349,N_29919);
xor UO_1433 (O_1433,N_28088,N_29450);
and UO_1434 (O_1434,N_29035,N_29634);
or UO_1435 (O_1435,N_29024,N_27301);
xor UO_1436 (O_1436,N_28839,N_27469);
nand UO_1437 (O_1437,N_28787,N_28522);
and UO_1438 (O_1438,N_28831,N_29270);
xnor UO_1439 (O_1439,N_28777,N_29472);
nor UO_1440 (O_1440,N_29903,N_29277);
nor UO_1441 (O_1441,N_28827,N_28912);
nand UO_1442 (O_1442,N_29423,N_27285);
or UO_1443 (O_1443,N_28849,N_27694);
and UO_1444 (O_1444,N_28398,N_28142);
or UO_1445 (O_1445,N_28554,N_28427);
xor UO_1446 (O_1446,N_27426,N_28786);
nand UO_1447 (O_1447,N_28259,N_27032);
xnor UO_1448 (O_1448,N_27864,N_29370);
xor UO_1449 (O_1449,N_29823,N_28804);
xor UO_1450 (O_1450,N_29933,N_29131);
xor UO_1451 (O_1451,N_29207,N_29532);
and UO_1452 (O_1452,N_28326,N_29461);
nand UO_1453 (O_1453,N_28652,N_29758);
nand UO_1454 (O_1454,N_28126,N_28633);
nand UO_1455 (O_1455,N_29473,N_29451);
or UO_1456 (O_1456,N_27763,N_28012);
nand UO_1457 (O_1457,N_27181,N_27359);
nand UO_1458 (O_1458,N_29081,N_28368);
nor UO_1459 (O_1459,N_29966,N_27355);
nand UO_1460 (O_1460,N_27647,N_27652);
or UO_1461 (O_1461,N_28416,N_27534);
nand UO_1462 (O_1462,N_27758,N_27717);
nor UO_1463 (O_1463,N_27640,N_27726);
xor UO_1464 (O_1464,N_28167,N_29078);
xnor UO_1465 (O_1465,N_29117,N_27499);
or UO_1466 (O_1466,N_27165,N_28748);
and UO_1467 (O_1467,N_28443,N_27283);
nor UO_1468 (O_1468,N_28863,N_27883);
or UO_1469 (O_1469,N_27056,N_29591);
xor UO_1470 (O_1470,N_29360,N_28983);
xor UO_1471 (O_1471,N_27959,N_29389);
xor UO_1472 (O_1472,N_28272,N_29694);
and UO_1473 (O_1473,N_28732,N_29096);
nand UO_1474 (O_1474,N_27101,N_27169);
and UO_1475 (O_1475,N_28415,N_29908);
xor UO_1476 (O_1476,N_27612,N_28979);
nand UO_1477 (O_1477,N_27228,N_29531);
or UO_1478 (O_1478,N_29782,N_27966);
nand UO_1479 (O_1479,N_28213,N_27856);
xnor UO_1480 (O_1480,N_27622,N_27476);
xnor UO_1481 (O_1481,N_27644,N_28218);
and UO_1482 (O_1482,N_29156,N_28773);
nand UO_1483 (O_1483,N_29004,N_28399);
and UO_1484 (O_1484,N_27776,N_28188);
or UO_1485 (O_1485,N_28937,N_29703);
nand UO_1486 (O_1486,N_29485,N_27277);
and UO_1487 (O_1487,N_29780,N_28203);
and UO_1488 (O_1488,N_27771,N_29868);
nor UO_1489 (O_1489,N_27207,N_29770);
and UO_1490 (O_1490,N_28414,N_28882);
nor UO_1491 (O_1491,N_29104,N_27278);
or UO_1492 (O_1492,N_29784,N_27229);
nor UO_1493 (O_1493,N_28296,N_27774);
nand UO_1494 (O_1494,N_29740,N_27536);
nand UO_1495 (O_1495,N_29262,N_29079);
nor UO_1496 (O_1496,N_27624,N_27715);
nor UO_1497 (O_1497,N_27342,N_29426);
xnor UO_1498 (O_1498,N_27282,N_29474);
xor UO_1499 (O_1499,N_28248,N_27501);
nor UO_1500 (O_1500,N_29201,N_28247);
nand UO_1501 (O_1501,N_27560,N_29190);
xnor UO_1502 (O_1502,N_27000,N_28508);
xor UO_1503 (O_1503,N_28683,N_27288);
nand UO_1504 (O_1504,N_27776,N_29233);
nor UO_1505 (O_1505,N_29121,N_27667);
and UO_1506 (O_1506,N_28794,N_29484);
and UO_1507 (O_1507,N_28074,N_29297);
and UO_1508 (O_1508,N_28819,N_29383);
nor UO_1509 (O_1509,N_29022,N_27949);
or UO_1510 (O_1510,N_28964,N_29741);
and UO_1511 (O_1511,N_28116,N_29424);
nor UO_1512 (O_1512,N_29287,N_28123);
nor UO_1513 (O_1513,N_29128,N_27657);
xnor UO_1514 (O_1514,N_27898,N_28562);
and UO_1515 (O_1515,N_29397,N_27507);
or UO_1516 (O_1516,N_27636,N_28192);
or UO_1517 (O_1517,N_29604,N_28188);
nand UO_1518 (O_1518,N_27942,N_28150);
xnor UO_1519 (O_1519,N_29309,N_28512);
nand UO_1520 (O_1520,N_29529,N_29516);
nand UO_1521 (O_1521,N_27864,N_27541);
and UO_1522 (O_1522,N_28489,N_28333);
or UO_1523 (O_1523,N_28597,N_27402);
xnor UO_1524 (O_1524,N_28841,N_28552);
and UO_1525 (O_1525,N_28294,N_28876);
and UO_1526 (O_1526,N_28028,N_28758);
and UO_1527 (O_1527,N_27408,N_27668);
xnor UO_1528 (O_1528,N_27434,N_28562);
nor UO_1529 (O_1529,N_29318,N_28381);
nand UO_1530 (O_1530,N_28952,N_27987);
xor UO_1531 (O_1531,N_29818,N_27269);
nor UO_1532 (O_1532,N_27362,N_29059);
xor UO_1533 (O_1533,N_29346,N_29995);
xor UO_1534 (O_1534,N_27129,N_28677);
and UO_1535 (O_1535,N_28852,N_29024);
nand UO_1536 (O_1536,N_28452,N_29356);
and UO_1537 (O_1537,N_28735,N_29550);
nor UO_1538 (O_1538,N_29447,N_28770);
nor UO_1539 (O_1539,N_28020,N_27559);
nand UO_1540 (O_1540,N_29242,N_29916);
or UO_1541 (O_1541,N_29721,N_29501);
nor UO_1542 (O_1542,N_27794,N_28969);
xnor UO_1543 (O_1543,N_28437,N_28953);
nor UO_1544 (O_1544,N_27462,N_27374);
nand UO_1545 (O_1545,N_27656,N_29246);
or UO_1546 (O_1546,N_28301,N_27360);
xnor UO_1547 (O_1547,N_27561,N_28283);
or UO_1548 (O_1548,N_28887,N_29962);
nor UO_1549 (O_1549,N_29135,N_28512);
or UO_1550 (O_1550,N_27089,N_28337);
and UO_1551 (O_1551,N_28281,N_28752);
nand UO_1552 (O_1552,N_28988,N_27686);
and UO_1553 (O_1553,N_27088,N_27603);
nand UO_1554 (O_1554,N_27142,N_28056);
xor UO_1555 (O_1555,N_29403,N_28922);
nand UO_1556 (O_1556,N_29046,N_29744);
or UO_1557 (O_1557,N_28168,N_29266);
xor UO_1558 (O_1558,N_28194,N_27391);
xor UO_1559 (O_1559,N_29725,N_28910);
xor UO_1560 (O_1560,N_29055,N_29180);
nand UO_1561 (O_1561,N_29260,N_28160);
and UO_1562 (O_1562,N_29040,N_29550);
nor UO_1563 (O_1563,N_29451,N_29096);
nand UO_1564 (O_1564,N_27370,N_27509);
or UO_1565 (O_1565,N_28300,N_29757);
nand UO_1566 (O_1566,N_27718,N_29010);
xor UO_1567 (O_1567,N_27355,N_29334);
nand UO_1568 (O_1568,N_28028,N_29704);
or UO_1569 (O_1569,N_29605,N_27272);
and UO_1570 (O_1570,N_28942,N_29170);
and UO_1571 (O_1571,N_27207,N_28762);
and UO_1572 (O_1572,N_29524,N_27416);
nor UO_1573 (O_1573,N_28682,N_28961);
and UO_1574 (O_1574,N_27980,N_27699);
nor UO_1575 (O_1575,N_27811,N_28638);
nand UO_1576 (O_1576,N_27057,N_28608);
or UO_1577 (O_1577,N_28333,N_29224);
or UO_1578 (O_1578,N_29963,N_29193);
nor UO_1579 (O_1579,N_27783,N_28679);
nor UO_1580 (O_1580,N_27393,N_27692);
xor UO_1581 (O_1581,N_28721,N_29047);
or UO_1582 (O_1582,N_28151,N_27229);
nand UO_1583 (O_1583,N_28314,N_27850);
nand UO_1584 (O_1584,N_27228,N_27745);
xor UO_1585 (O_1585,N_29622,N_29321);
and UO_1586 (O_1586,N_29405,N_28145);
and UO_1587 (O_1587,N_29184,N_28752);
xnor UO_1588 (O_1588,N_27200,N_27515);
nor UO_1589 (O_1589,N_27896,N_27837);
and UO_1590 (O_1590,N_29497,N_27715);
xnor UO_1591 (O_1591,N_27350,N_29652);
nor UO_1592 (O_1592,N_28469,N_29713);
or UO_1593 (O_1593,N_27771,N_29060);
xnor UO_1594 (O_1594,N_27100,N_28086);
or UO_1595 (O_1595,N_28262,N_29281);
xor UO_1596 (O_1596,N_27137,N_27789);
xnor UO_1597 (O_1597,N_29354,N_27663);
and UO_1598 (O_1598,N_27104,N_28668);
nand UO_1599 (O_1599,N_28234,N_28219);
xor UO_1600 (O_1600,N_27159,N_27790);
xor UO_1601 (O_1601,N_29025,N_27035);
nor UO_1602 (O_1602,N_27113,N_27680);
nand UO_1603 (O_1603,N_28521,N_28681);
nor UO_1604 (O_1604,N_27860,N_28628);
and UO_1605 (O_1605,N_28044,N_27869);
or UO_1606 (O_1606,N_28253,N_29643);
and UO_1607 (O_1607,N_29673,N_29469);
nor UO_1608 (O_1608,N_29605,N_29089);
nand UO_1609 (O_1609,N_28293,N_27817);
and UO_1610 (O_1610,N_27764,N_29483);
or UO_1611 (O_1611,N_29304,N_28157);
xnor UO_1612 (O_1612,N_27924,N_29749);
nor UO_1613 (O_1613,N_29542,N_27536);
nor UO_1614 (O_1614,N_27614,N_28731);
or UO_1615 (O_1615,N_28043,N_28997);
and UO_1616 (O_1616,N_28022,N_28432);
nand UO_1617 (O_1617,N_29313,N_29984);
nand UO_1618 (O_1618,N_27764,N_28799);
and UO_1619 (O_1619,N_29724,N_28231);
nand UO_1620 (O_1620,N_27199,N_28108);
or UO_1621 (O_1621,N_27545,N_28203);
nor UO_1622 (O_1622,N_29047,N_27365);
xnor UO_1623 (O_1623,N_27028,N_28512);
and UO_1624 (O_1624,N_27151,N_29890);
nand UO_1625 (O_1625,N_28674,N_27232);
xnor UO_1626 (O_1626,N_27071,N_27204);
and UO_1627 (O_1627,N_29792,N_29251);
and UO_1628 (O_1628,N_28871,N_29193);
nand UO_1629 (O_1629,N_29715,N_28588);
xnor UO_1630 (O_1630,N_27103,N_27217);
xnor UO_1631 (O_1631,N_27967,N_27947);
or UO_1632 (O_1632,N_27262,N_27630);
nor UO_1633 (O_1633,N_27083,N_28817);
and UO_1634 (O_1634,N_29769,N_28503);
nand UO_1635 (O_1635,N_28525,N_27185);
or UO_1636 (O_1636,N_29998,N_27183);
nand UO_1637 (O_1637,N_27463,N_27252);
nor UO_1638 (O_1638,N_27400,N_28476);
or UO_1639 (O_1639,N_27688,N_28717);
and UO_1640 (O_1640,N_28533,N_28222);
nor UO_1641 (O_1641,N_27034,N_28464);
xor UO_1642 (O_1642,N_28877,N_29175);
or UO_1643 (O_1643,N_27171,N_29830);
xor UO_1644 (O_1644,N_29406,N_28208);
nor UO_1645 (O_1645,N_29837,N_27249);
nor UO_1646 (O_1646,N_28200,N_28705);
nor UO_1647 (O_1647,N_27320,N_29951);
nor UO_1648 (O_1648,N_28287,N_29550);
xor UO_1649 (O_1649,N_29802,N_28100);
or UO_1650 (O_1650,N_29385,N_29220);
xnor UO_1651 (O_1651,N_27255,N_29267);
or UO_1652 (O_1652,N_27562,N_29423);
and UO_1653 (O_1653,N_28389,N_28214);
xnor UO_1654 (O_1654,N_27398,N_28678);
xor UO_1655 (O_1655,N_28976,N_28996);
xor UO_1656 (O_1656,N_29773,N_29632);
xnor UO_1657 (O_1657,N_28107,N_28035);
or UO_1658 (O_1658,N_27167,N_28864);
nand UO_1659 (O_1659,N_28441,N_29886);
xor UO_1660 (O_1660,N_29144,N_27083);
nand UO_1661 (O_1661,N_27736,N_27081);
or UO_1662 (O_1662,N_27557,N_29492);
nor UO_1663 (O_1663,N_28575,N_28435);
and UO_1664 (O_1664,N_28938,N_29270);
nand UO_1665 (O_1665,N_29545,N_29221);
xnor UO_1666 (O_1666,N_27245,N_29745);
xor UO_1667 (O_1667,N_29916,N_27077);
nor UO_1668 (O_1668,N_28247,N_27337);
and UO_1669 (O_1669,N_29325,N_27317);
or UO_1670 (O_1670,N_28405,N_28355);
nor UO_1671 (O_1671,N_29043,N_28318);
and UO_1672 (O_1672,N_29491,N_29686);
nor UO_1673 (O_1673,N_29981,N_28716);
nand UO_1674 (O_1674,N_27352,N_27300);
nand UO_1675 (O_1675,N_29748,N_29336);
and UO_1676 (O_1676,N_29463,N_28211);
or UO_1677 (O_1677,N_28506,N_29602);
nor UO_1678 (O_1678,N_28262,N_27003);
xor UO_1679 (O_1679,N_27687,N_27445);
or UO_1680 (O_1680,N_27714,N_28416);
nor UO_1681 (O_1681,N_29678,N_29447);
nor UO_1682 (O_1682,N_27188,N_28396);
xor UO_1683 (O_1683,N_27690,N_28351);
and UO_1684 (O_1684,N_28196,N_28357);
or UO_1685 (O_1685,N_27888,N_28766);
nand UO_1686 (O_1686,N_28961,N_28761);
or UO_1687 (O_1687,N_29037,N_29917);
xor UO_1688 (O_1688,N_28499,N_28762);
xnor UO_1689 (O_1689,N_27335,N_29365);
or UO_1690 (O_1690,N_29473,N_27495);
xor UO_1691 (O_1691,N_28468,N_28818);
nand UO_1692 (O_1692,N_28638,N_27997);
nor UO_1693 (O_1693,N_28598,N_27214);
and UO_1694 (O_1694,N_29405,N_29491);
or UO_1695 (O_1695,N_28642,N_28315);
xnor UO_1696 (O_1696,N_27608,N_29332);
and UO_1697 (O_1697,N_28683,N_29058);
nand UO_1698 (O_1698,N_29982,N_27028);
and UO_1699 (O_1699,N_28891,N_27089);
xor UO_1700 (O_1700,N_27121,N_28245);
xor UO_1701 (O_1701,N_29841,N_28024);
nand UO_1702 (O_1702,N_27722,N_29836);
xor UO_1703 (O_1703,N_29297,N_28099);
xnor UO_1704 (O_1704,N_28647,N_28387);
or UO_1705 (O_1705,N_27498,N_29836);
xor UO_1706 (O_1706,N_29219,N_28738);
and UO_1707 (O_1707,N_29223,N_27415);
or UO_1708 (O_1708,N_29744,N_27057);
nor UO_1709 (O_1709,N_28080,N_27009);
xnor UO_1710 (O_1710,N_28655,N_27022);
nor UO_1711 (O_1711,N_27141,N_29520);
nand UO_1712 (O_1712,N_27024,N_28158);
xnor UO_1713 (O_1713,N_27217,N_29812);
xor UO_1714 (O_1714,N_29693,N_29057);
or UO_1715 (O_1715,N_28308,N_27215);
xor UO_1716 (O_1716,N_28799,N_29806);
and UO_1717 (O_1717,N_29502,N_28562);
or UO_1718 (O_1718,N_27694,N_28816);
and UO_1719 (O_1719,N_28961,N_29762);
xnor UO_1720 (O_1720,N_29167,N_27396);
or UO_1721 (O_1721,N_29145,N_28587);
or UO_1722 (O_1722,N_28666,N_28029);
nor UO_1723 (O_1723,N_29902,N_29336);
xnor UO_1724 (O_1724,N_29996,N_27499);
nor UO_1725 (O_1725,N_28942,N_28905);
nor UO_1726 (O_1726,N_28682,N_29727);
or UO_1727 (O_1727,N_27206,N_29643);
or UO_1728 (O_1728,N_29522,N_27575);
xnor UO_1729 (O_1729,N_27007,N_29806);
or UO_1730 (O_1730,N_28659,N_27608);
and UO_1731 (O_1731,N_28714,N_28998);
or UO_1732 (O_1732,N_27274,N_28774);
or UO_1733 (O_1733,N_28108,N_27662);
nand UO_1734 (O_1734,N_27740,N_28268);
and UO_1735 (O_1735,N_29794,N_28508);
nand UO_1736 (O_1736,N_29413,N_29854);
and UO_1737 (O_1737,N_27627,N_29514);
nand UO_1738 (O_1738,N_27262,N_27612);
xnor UO_1739 (O_1739,N_28717,N_28506);
nor UO_1740 (O_1740,N_29227,N_27862);
and UO_1741 (O_1741,N_27155,N_29691);
xor UO_1742 (O_1742,N_28125,N_27096);
or UO_1743 (O_1743,N_27809,N_29196);
nor UO_1744 (O_1744,N_27957,N_27724);
nor UO_1745 (O_1745,N_28162,N_29452);
nor UO_1746 (O_1746,N_27932,N_27018);
and UO_1747 (O_1747,N_28417,N_27668);
nand UO_1748 (O_1748,N_29418,N_28233);
nand UO_1749 (O_1749,N_27852,N_28444);
and UO_1750 (O_1750,N_28601,N_27598);
nor UO_1751 (O_1751,N_27823,N_28186);
or UO_1752 (O_1752,N_27819,N_29172);
or UO_1753 (O_1753,N_29329,N_27701);
xor UO_1754 (O_1754,N_27743,N_28582);
nand UO_1755 (O_1755,N_28430,N_28455);
and UO_1756 (O_1756,N_29256,N_29614);
and UO_1757 (O_1757,N_27630,N_28761);
and UO_1758 (O_1758,N_27736,N_29336);
xnor UO_1759 (O_1759,N_29167,N_28201);
xor UO_1760 (O_1760,N_29713,N_27816);
xnor UO_1761 (O_1761,N_27589,N_28898);
or UO_1762 (O_1762,N_29064,N_28251);
or UO_1763 (O_1763,N_29867,N_27307);
nand UO_1764 (O_1764,N_28805,N_27719);
nor UO_1765 (O_1765,N_29956,N_28431);
and UO_1766 (O_1766,N_28205,N_29742);
and UO_1767 (O_1767,N_29000,N_27944);
or UO_1768 (O_1768,N_27436,N_29732);
or UO_1769 (O_1769,N_27033,N_28161);
nor UO_1770 (O_1770,N_28735,N_29235);
nand UO_1771 (O_1771,N_28570,N_29397);
nor UO_1772 (O_1772,N_28437,N_28315);
nor UO_1773 (O_1773,N_28872,N_29537);
nand UO_1774 (O_1774,N_27566,N_29889);
xor UO_1775 (O_1775,N_28875,N_27014);
nand UO_1776 (O_1776,N_27536,N_28873);
or UO_1777 (O_1777,N_29226,N_28008);
nand UO_1778 (O_1778,N_28425,N_29749);
xnor UO_1779 (O_1779,N_29524,N_27897);
nor UO_1780 (O_1780,N_27418,N_28916);
xor UO_1781 (O_1781,N_29997,N_27158);
nor UO_1782 (O_1782,N_29713,N_27966);
nor UO_1783 (O_1783,N_27646,N_27074);
nand UO_1784 (O_1784,N_29866,N_27127);
nor UO_1785 (O_1785,N_29793,N_27364);
and UO_1786 (O_1786,N_28164,N_28371);
or UO_1787 (O_1787,N_28848,N_28417);
nor UO_1788 (O_1788,N_29817,N_28727);
nor UO_1789 (O_1789,N_27181,N_27694);
and UO_1790 (O_1790,N_27467,N_28211);
xor UO_1791 (O_1791,N_27098,N_29584);
xor UO_1792 (O_1792,N_29619,N_29708);
xnor UO_1793 (O_1793,N_29885,N_29515);
nand UO_1794 (O_1794,N_29138,N_29257);
and UO_1795 (O_1795,N_29950,N_27293);
xor UO_1796 (O_1796,N_29782,N_29278);
and UO_1797 (O_1797,N_27128,N_28763);
and UO_1798 (O_1798,N_29013,N_27221);
or UO_1799 (O_1799,N_29889,N_29331);
nor UO_1800 (O_1800,N_29003,N_29664);
xor UO_1801 (O_1801,N_28294,N_27803);
nor UO_1802 (O_1802,N_28121,N_28805);
nor UO_1803 (O_1803,N_28179,N_29231);
xnor UO_1804 (O_1804,N_28492,N_28452);
xnor UO_1805 (O_1805,N_28093,N_27691);
nand UO_1806 (O_1806,N_27705,N_29693);
xor UO_1807 (O_1807,N_27899,N_28369);
nand UO_1808 (O_1808,N_29557,N_27282);
nor UO_1809 (O_1809,N_27453,N_27165);
nor UO_1810 (O_1810,N_29296,N_29564);
xor UO_1811 (O_1811,N_29484,N_29838);
nand UO_1812 (O_1812,N_27850,N_28789);
or UO_1813 (O_1813,N_29747,N_29200);
xor UO_1814 (O_1814,N_28383,N_29138);
nor UO_1815 (O_1815,N_27416,N_28429);
nand UO_1816 (O_1816,N_27094,N_28007);
and UO_1817 (O_1817,N_28332,N_29404);
nor UO_1818 (O_1818,N_28120,N_27595);
nand UO_1819 (O_1819,N_28255,N_29347);
or UO_1820 (O_1820,N_28962,N_29550);
or UO_1821 (O_1821,N_28373,N_28090);
nor UO_1822 (O_1822,N_28172,N_27179);
xnor UO_1823 (O_1823,N_29451,N_28513);
or UO_1824 (O_1824,N_27025,N_28580);
and UO_1825 (O_1825,N_27125,N_27948);
nand UO_1826 (O_1826,N_27210,N_29205);
xnor UO_1827 (O_1827,N_27734,N_29019);
xor UO_1828 (O_1828,N_29621,N_27354);
nand UO_1829 (O_1829,N_27601,N_29193);
nor UO_1830 (O_1830,N_27813,N_28885);
xnor UO_1831 (O_1831,N_28249,N_27960);
xnor UO_1832 (O_1832,N_27328,N_27190);
nor UO_1833 (O_1833,N_28470,N_29441);
nand UO_1834 (O_1834,N_29162,N_28920);
nand UO_1835 (O_1835,N_29169,N_28790);
nand UO_1836 (O_1836,N_28804,N_27171);
nand UO_1837 (O_1837,N_27026,N_28409);
and UO_1838 (O_1838,N_29588,N_28211);
xor UO_1839 (O_1839,N_29523,N_28565);
nor UO_1840 (O_1840,N_28084,N_27852);
or UO_1841 (O_1841,N_28945,N_29589);
xnor UO_1842 (O_1842,N_27654,N_27157);
nand UO_1843 (O_1843,N_29823,N_28635);
nor UO_1844 (O_1844,N_29762,N_28348);
or UO_1845 (O_1845,N_29685,N_29203);
and UO_1846 (O_1846,N_28890,N_29311);
nand UO_1847 (O_1847,N_28546,N_28109);
xnor UO_1848 (O_1848,N_28575,N_27881);
or UO_1849 (O_1849,N_29667,N_29310);
and UO_1850 (O_1850,N_29240,N_29896);
nand UO_1851 (O_1851,N_27040,N_28035);
xor UO_1852 (O_1852,N_27996,N_28322);
xor UO_1853 (O_1853,N_28451,N_28253);
nand UO_1854 (O_1854,N_27322,N_29547);
or UO_1855 (O_1855,N_29585,N_27786);
nand UO_1856 (O_1856,N_28880,N_28481);
and UO_1857 (O_1857,N_29483,N_27624);
xor UO_1858 (O_1858,N_28824,N_28365);
xor UO_1859 (O_1859,N_29295,N_29319);
and UO_1860 (O_1860,N_27368,N_28793);
nor UO_1861 (O_1861,N_27895,N_27126);
nand UO_1862 (O_1862,N_27505,N_28876);
nor UO_1863 (O_1863,N_27036,N_28993);
xnor UO_1864 (O_1864,N_27302,N_28678);
nand UO_1865 (O_1865,N_28919,N_27694);
nor UO_1866 (O_1866,N_27017,N_27720);
and UO_1867 (O_1867,N_29818,N_27126);
xnor UO_1868 (O_1868,N_27711,N_28694);
or UO_1869 (O_1869,N_27935,N_28229);
nand UO_1870 (O_1870,N_28450,N_28979);
and UO_1871 (O_1871,N_29455,N_27762);
or UO_1872 (O_1872,N_29150,N_27452);
nand UO_1873 (O_1873,N_28190,N_27356);
nor UO_1874 (O_1874,N_27027,N_27376);
nand UO_1875 (O_1875,N_29287,N_29330);
nor UO_1876 (O_1876,N_29679,N_27142);
xnor UO_1877 (O_1877,N_29410,N_29431);
xor UO_1878 (O_1878,N_29456,N_27577);
xnor UO_1879 (O_1879,N_28979,N_29677);
or UO_1880 (O_1880,N_27667,N_29705);
and UO_1881 (O_1881,N_28949,N_27935);
nor UO_1882 (O_1882,N_29353,N_27168);
nand UO_1883 (O_1883,N_27107,N_27602);
nand UO_1884 (O_1884,N_27541,N_28712);
nand UO_1885 (O_1885,N_29278,N_27058);
nand UO_1886 (O_1886,N_27318,N_29258);
and UO_1887 (O_1887,N_27261,N_28060);
nor UO_1888 (O_1888,N_28861,N_27008);
xnor UO_1889 (O_1889,N_27317,N_27005);
nand UO_1890 (O_1890,N_27590,N_27350);
nor UO_1891 (O_1891,N_27679,N_28741);
xor UO_1892 (O_1892,N_29256,N_27815);
xnor UO_1893 (O_1893,N_29463,N_28589);
xnor UO_1894 (O_1894,N_28740,N_29618);
or UO_1895 (O_1895,N_27219,N_27878);
and UO_1896 (O_1896,N_27152,N_29497);
xor UO_1897 (O_1897,N_29351,N_29931);
and UO_1898 (O_1898,N_28996,N_29862);
xor UO_1899 (O_1899,N_29372,N_27360);
or UO_1900 (O_1900,N_28352,N_29866);
xor UO_1901 (O_1901,N_29383,N_29816);
nor UO_1902 (O_1902,N_29797,N_28461);
xor UO_1903 (O_1903,N_27140,N_28981);
xor UO_1904 (O_1904,N_28872,N_27535);
and UO_1905 (O_1905,N_27330,N_27408);
nor UO_1906 (O_1906,N_28036,N_28581);
xnor UO_1907 (O_1907,N_27891,N_28990);
xnor UO_1908 (O_1908,N_29826,N_29271);
xor UO_1909 (O_1909,N_27341,N_29308);
nand UO_1910 (O_1910,N_29722,N_27438);
nand UO_1911 (O_1911,N_27697,N_27412);
and UO_1912 (O_1912,N_27423,N_27817);
xor UO_1913 (O_1913,N_28107,N_27537);
or UO_1914 (O_1914,N_27571,N_29326);
nand UO_1915 (O_1915,N_27076,N_28508);
or UO_1916 (O_1916,N_27311,N_27630);
nand UO_1917 (O_1917,N_27603,N_27586);
or UO_1918 (O_1918,N_29805,N_29678);
nand UO_1919 (O_1919,N_29197,N_29379);
and UO_1920 (O_1920,N_27910,N_27471);
nand UO_1921 (O_1921,N_29157,N_28132);
nand UO_1922 (O_1922,N_29997,N_27346);
nor UO_1923 (O_1923,N_28970,N_29560);
or UO_1924 (O_1924,N_29367,N_27927);
and UO_1925 (O_1925,N_29682,N_27823);
xor UO_1926 (O_1926,N_29215,N_27369);
and UO_1927 (O_1927,N_27386,N_29034);
xnor UO_1928 (O_1928,N_29472,N_28058);
nor UO_1929 (O_1929,N_29715,N_27045);
nand UO_1930 (O_1930,N_28832,N_28916);
or UO_1931 (O_1931,N_29391,N_28229);
xnor UO_1932 (O_1932,N_27964,N_29174);
nor UO_1933 (O_1933,N_28930,N_27588);
xor UO_1934 (O_1934,N_28988,N_27826);
nand UO_1935 (O_1935,N_27156,N_29383);
nand UO_1936 (O_1936,N_27822,N_27665);
nand UO_1937 (O_1937,N_27097,N_27875);
nand UO_1938 (O_1938,N_28522,N_27343);
or UO_1939 (O_1939,N_27489,N_29683);
xor UO_1940 (O_1940,N_29202,N_27996);
or UO_1941 (O_1941,N_29771,N_28078);
nor UO_1942 (O_1942,N_28044,N_28422);
xor UO_1943 (O_1943,N_29088,N_27803);
or UO_1944 (O_1944,N_27630,N_28549);
nor UO_1945 (O_1945,N_28993,N_28328);
nand UO_1946 (O_1946,N_29330,N_27965);
or UO_1947 (O_1947,N_28323,N_27212);
nor UO_1948 (O_1948,N_28979,N_28826);
or UO_1949 (O_1949,N_27717,N_28261);
or UO_1950 (O_1950,N_27005,N_29068);
or UO_1951 (O_1951,N_28521,N_29686);
xnor UO_1952 (O_1952,N_28400,N_27142);
or UO_1953 (O_1953,N_29625,N_28111);
nand UO_1954 (O_1954,N_27229,N_27982);
nand UO_1955 (O_1955,N_28277,N_28104);
xnor UO_1956 (O_1956,N_29707,N_29369);
nor UO_1957 (O_1957,N_28123,N_27986);
xor UO_1958 (O_1958,N_29355,N_29103);
nand UO_1959 (O_1959,N_27291,N_29325);
nor UO_1960 (O_1960,N_28828,N_27619);
nor UO_1961 (O_1961,N_27778,N_27692);
nand UO_1962 (O_1962,N_28924,N_28826);
or UO_1963 (O_1963,N_29716,N_29901);
or UO_1964 (O_1964,N_27604,N_28336);
nand UO_1965 (O_1965,N_29726,N_28799);
nor UO_1966 (O_1966,N_29021,N_27692);
xnor UO_1967 (O_1967,N_29096,N_29033);
and UO_1968 (O_1968,N_28363,N_29435);
nand UO_1969 (O_1969,N_29641,N_28958);
nand UO_1970 (O_1970,N_29988,N_28945);
and UO_1971 (O_1971,N_28898,N_29169);
nand UO_1972 (O_1972,N_28171,N_28834);
or UO_1973 (O_1973,N_27995,N_27719);
xor UO_1974 (O_1974,N_27727,N_27808);
nand UO_1975 (O_1975,N_27406,N_28086);
and UO_1976 (O_1976,N_28289,N_27576);
and UO_1977 (O_1977,N_28373,N_27927);
and UO_1978 (O_1978,N_27481,N_29873);
or UO_1979 (O_1979,N_28226,N_27414);
and UO_1980 (O_1980,N_28252,N_29524);
nand UO_1981 (O_1981,N_27273,N_29602);
or UO_1982 (O_1982,N_29143,N_27501);
and UO_1983 (O_1983,N_28372,N_27297);
nor UO_1984 (O_1984,N_28201,N_29993);
or UO_1985 (O_1985,N_27734,N_27146);
or UO_1986 (O_1986,N_27925,N_27726);
or UO_1987 (O_1987,N_28611,N_27695);
and UO_1988 (O_1988,N_28358,N_28106);
xor UO_1989 (O_1989,N_27593,N_27974);
nor UO_1990 (O_1990,N_29816,N_27018);
nor UO_1991 (O_1991,N_28045,N_28700);
and UO_1992 (O_1992,N_28224,N_27958);
nand UO_1993 (O_1993,N_27597,N_28988);
and UO_1994 (O_1994,N_28490,N_28066);
nor UO_1995 (O_1995,N_27848,N_29019);
nor UO_1996 (O_1996,N_28702,N_28696);
and UO_1997 (O_1997,N_29502,N_28487);
nand UO_1998 (O_1998,N_28071,N_29284);
nor UO_1999 (O_1999,N_28923,N_28906);
xnor UO_2000 (O_2000,N_27028,N_28973);
nand UO_2001 (O_2001,N_29775,N_29921);
or UO_2002 (O_2002,N_27692,N_28703);
nor UO_2003 (O_2003,N_29152,N_28616);
xor UO_2004 (O_2004,N_27049,N_27285);
or UO_2005 (O_2005,N_28395,N_28252);
xnor UO_2006 (O_2006,N_27761,N_28745);
and UO_2007 (O_2007,N_27938,N_27005);
and UO_2008 (O_2008,N_27494,N_27306);
or UO_2009 (O_2009,N_28037,N_29481);
nand UO_2010 (O_2010,N_29348,N_28498);
and UO_2011 (O_2011,N_29743,N_29470);
or UO_2012 (O_2012,N_29304,N_28360);
nand UO_2013 (O_2013,N_27005,N_27875);
and UO_2014 (O_2014,N_27450,N_28832);
and UO_2015 (O_2015,N_27231,N_29993);
or UO_2016 (O_2016,N_27276,N_29535);
and UO_2017 (O_2017,N_28783,N_29762);
or UO_2018 (O_2018,N_27023,N_29801);
xnor UO_2019 (O_2019,N_27615,N_28898);
nand UO_2020 (O_2020,N_28733,N_29387);
nor UO_2021 (O_2021,N_28778,N_29199);
nand UO_2022 (O_2022,N_28445,N_28471);
and UO_2023 (O_2023,N_29160,N_27685);
nand UO_2024 (O_2024,N_28242,N_28116);
xnor UO_2025 (O_2025,N_28481,N_27050);
and UO_2026 (O_2026,N_29786,N_27638);
xnor UO_2027 (O_2027,N_29348,N_27572);
or UO_2028 (O_2028,N_28351,N_29893);
nand UO_2029 (O_2029,N_27555,N_27774);
xnor UO_2030 (O_2030,N_27885,N_29225);
nor UO_2031 (O_2031,N_28299,N_28087);
nand UO_2032 (O_2032,N_29943,N_29136);
or UO_2033 (O_2033,N_29323,N_27253);
xor UO_2034 (O_2034,N_28941,N_28937);
nand UO_2035 (O_2035,N_27852,N_29090);
nand UO_2036 (O_2036,N_28933,N_29998);
nor UO_2037 (O_2037,N_28963,N_28155);
and UO_2038 (O_2038,N_29602,N_27652);
nand UO_2039 (O_2039,N_27153,N_28868);
or UO_2040 (O_2040,N_27780,N_28846);
nor UO_2041 (O_2041,N_27600,N_28026);
or UO_2042 (O_2042,N_28116,N_27842);
nand UO_2043 (O_2043,N_27248,N_27184);
and UO_2044 (O_2044,N_28931,N_27108);
xnor UO_2045 (O_2045,N_27322,N_29213);
nor UO_2046 (O_2046,N_29106,N_27636);
and UO_2047 (O_2047,N_27618,N_29460);
xor UO_2048 (O_2048,N_28905,N_27939);
nand UO_2049 (O_2049,N_29409,N_28397);
nand UO_2050 (O_2050,N_29642,N_29339);
or UO_2051 (O_2051,N_29012,N_27701);
or UO_2052 (O_2052,N_29819,N_28119);
nand UO_2053 (O_2053,N_29087,N_29769);
and UO_2054 (O_2054,N_29158,N_27854);
xnor UO_2055 (O_2055,N_29478,N_28776);
nor UO_2056 (O_2056,N_27601,N_28655);
or UO_2057 (O_2057,N_29821,N_28809);
nand UO_2058 (O_2058,N_27819,N_27439);
or UO_2059 (O_2059,N_29035,N_28298);
and UO_2060 (O_2060,N_29446,N_28530);
and UO_2061 (O_2061,N_28276,N_28869);
or UO_2062 (O_2062,N_29312,N_27637);
xor UO_2063 (O_2063,N_29563,N_29415);
or UO_2064 (O_2064,N_27492,N_29484);
nor UO_2065 (O_2065,N_28440,N_29980);
nand UO_2066 (O_2066,N_27193,N_28583);
or UO_2067 (O_2067,N_27900,N_29798);
or UO_2068 (O_2068,N_29856,N_29861);
and UO_2069 (O_2069,N_29663,N_29277);
xnor UO_2070 (O_2070,N_27842,N_27685);
nand UO_2071 (O_2071,N_28629,N_29742);
nor UO_2072 (O_2072,N_28138,N_28159);
nand UO_2073 (O_2073,N_29436,N_27271);
xor UO_2074 (O_2074,N_28305,N_27416);
nor UO_2075 (O_2075,N_28904,N_29046);
nand UO_2076 (O_2076,N_27140,N_29482);
or UO_2077 (O_2077,N_27073,N_27715);
xor UO_2078 (O_2078,N_27568,N_29153);
or UO_2079 (O_2079,N_29153,N_28126);
nor UO_2080 (O_2080,N_29980,N_27553);
and UO_2081 (O_2081,N_28930,N_28264);
xnor UO_2082 (O_2082,N_27828,N_27518);
nand UO_2083 (O_2083,N_29297,N_29807);
and UO_2084 (O_2084,N_28093,N_29020);
xor UO_2085 (O_2085,N_29098,N_28299);
or UO_2086 (O_2086,N_27043,N_27438);
nor UO_2087 (O_2087,N_28899,N_29352);
or UO_2088 (O_2088,N_27244,N_27105);
or UO_2089 (O_2089,N_27529,N_28190);
nand UO_2090 (O_2090,N_27344,N_27531);
nand UO_2091 (O_2091,N_29072,N_29607);
nand UO_2092 (O_2092,N_27582,N_27343);
and UO_2093 (O_2093,N_28214,N_28404);
and UO_2094 (O_2094,N_28681,N_28186);
nand UO_2095 (O_2095,N_29958,N_28193);
or UO_2096 (O_2096,N_29716,N_28237);
xor UO_2097 (O_2097,N_28673,N_28757);
xor UO_2098 (O_2098,N_29098,N_27406);
xnor UO_2099 (O_2099,N_29143,N_27950);
and UO_2100 (O_2100,N_29451,N_29982);
and UO_2101 (O_2101,N_28424,N_28340);
or UO_2102 (O_2102,N_27925,N_27288);
and UO_2103 (O_2103,N_28599,N_28661);
nor UO_2104 (O_2104,N_27685,N_28663);
nand UO_2105 (O_2105,N_29616,N_29128);
and UO_2106 (O_2106,N_28659,N_27134);
or UO_2107 (O_2107,N_27952,N_28778);
nor UO_2108 (O_2108,N_27067,N_28193);
nand UO_2109 (O_2109,N_29206,N_27914);
nand UO_2110 (O_2110,N_27441,N_29247);
and UO_2111 (O_2111,N_29836,N_28736);
or UO_2112 (O_2112,N_27942,N_29710);
or UO_2113 (O_2113,N_29027,N_27866);
nand UO_2114 (O_2114,N_29448,N_29830);
xor UO_2115 (O_2115,N_29873,N_28605);
and UO_2116 (O_2116,N_28769,N_29790);
and UO_2117 (O_2117,N_27017,N_29595);
nor UO_2118 (O_2118,N_28159,N_27157);
xor UO_2119 (O_2119,N_28952,N_28912);
xor UO_2120 (O_2120,N_27730,N_27311);
or UO_2121 (O_2121,N_27157,N_27203);
xor UO_2122 (O_2122,N_29601,N_28266);
xor UO_2123 (O_2123,N_27057,N_28449);
nor UO_2124 (O_2124,N_29685,N_29127);
nor UO_2125 (O_2125,N_28101,N_28724);
nor UO_2126 (O_2126,N_29208,N_27232);
xor UO_2127 (O_2127,N_29463,N_27014);
nand UO_2128 (O_2128,N_28973,N_28787);
nand UO_2129 (O_2129,N_28135,N_29724);
and UO_2130 (O_2130,N_28215,N_29058);
xnor UO_2131 (O_2131,N_29517,N_29757);
or UO_2132 (O_2132,N_29536,N_27320);
xor UO_2133 (O_2133,N_27560,N_29789);
xor UO_2134 (O_2134,N_29413,N_27877);
nor UO_2135 (O_2135,N_27036,N_29943);
or UO_2136 (O_2136,N_29607,N_29356);
nor UO_2137 (O_2137,N_28531,N_28935);
nor UO_2138 (O_2138,N_29380,N_29347);
and UO_2139 (O_2139,N_29394,N_28472);
xnor UO_2140 (O_2140,N_27341,N_29870);
and UO_2141 (O_2141,N_27980,N_29994);
nand UO_2142 (O_2142,N_29933,N_29325);
and UO_2143 (O_2143,N_27469,N_29212);
xor UO_2144 (O_2144,N_28756,N_29588);
and UO_2145 (O_2145,N_28880,N_29684);
nor UO_2146 (O_2146,N_27100,N_28053);
or UO_2147 (O_2147,N_27721,N_28176);
xnor UO_2148 (O_2148,N_28592,N_27634);
nand UO_2149 (O_2149,N_29959,N_28250);
or UO_2150 (O_2150,N_28995,N_27691);
and UO_2151 (O_2151,N_27384,N_29579);
nor UO_2152 (O_2152,N_29598,N_29135);
or UO_2153 (O_2153,N_28062,N_28787);
nand UO_2154 (O_2154,N_29438,N_27512);
nor UO_2155 (O_2155,N_27692,N_27810);
xor UO_2156 (O_2156,N_28775,N_29779);
xor UO_2157 (O_2157,N_28068,N_29346);
nor UO_2158 (O_2158,N_29441,N_28828);
xnor UO_2159 (O_2159,N_29784,N_27479);
and UO_2160 (O_2160,N_28205,N_28473);
nor UO_2161 (O_2161,N_27956,N_28467);
xnor UO_2162 (O_2162,N_29436,N_29132);
and UO_2163 (O_2163,N_29838,N_28976);
nor UO_2164 (O_2164,N_29141,N_27987);
xnor UO_2165 (O_2165,N_28273,N_27738);
and UO_2166 (O_2166,N_28044,N_27845);
nand UO_2167 (O_2167,N_27779,N_29364);
and UO_2168 (O_2168,N_29278,N_27162);
or UO_2169 (O_2169,N_27615,N_29246);
xnor UO_2170 (O_2170,N_28525,N_29719);
xor UO_2171 (O_2171,N_29579,N_29801);
nand UO_2172 (O_2172,N_27707,N_28017);
nor UO_2173 (O_2173,N_27462,N_28831);
nor UO_2174 (O_2174,N_28450,N_28040);
or UO_2175 (O_2175,N_28770,N_29346);
xnor UO_2176 (O_2176,N_29564,N_29112);
nand UO_2177 (O_2177,N_29271,N_27847);
and UO_2178 (O_2178,N_28692,N_29379);
and UO_2179 (O_2179,N_28966,N_28718);
nor UO_2180 (O_2180,N_27507,N_28997);
xor UO_2181 (O_2181,N_27717,N_28032);
xor UO_2182 (O_2182,N_29360,N_28528);
xor UO_2183 (O_2183,N_29549,N_29258);
and UO_2184 (O_2184,N_28978,N_29657);
or UO_2185 (O_2185,N_28070,N_27768);
nand UO_2186 (O_2186,N_29793,N_29383);
nand UO_2187 (O_2187,N_29961,N_28062);
or UO_2188 (O_2188,N_27833,N_29233);
xnor UO_2189 (O_2189,N_27983,N_28175);
nor UO_2190 (O_2190,N_29487,N_27003);
xnor UO_2191 (O_2191,N_29392,N_29203);
xor UO_2192 (O_2192,N_28062,N_27510);
or UO_2193 (O_2193,N_28375,N_28824);
and UO_2194 (O_2194,N_27413,N_28437);
or UO_2195 (O_2195,N_28621,N_27112);
xor UO_2196 (O_2196,N_27066,N_27797);
nand UO_2197 (O_2197,N_28235,N_27098);
nand UO_2198 (O_2198,N_27572,N_29001);
or UO_2199 (O_2199,N_28552,N_29236);
nand UO_2200 (O_2200,N_29848,N_27020);
nor UO_2201 (O_2201,N_27624,N_28133);
nor UO_2202 (O_2202,N_27352,N_29834);
or UO_2203 (O_2203,N_27211,N_28047);
xnor UO_2204 (O_2204,N_28309,N_28279);
or UO_2205 (O_2205,N_27201,N_27739);
and UO_2206 (O_2206,N_28591,N_29118);
nor UO_2207 (O_2207,N_29639,N_28779);
nand UO_2208 (O_2208,N_29593,N_28520);
or UO_2209 (O_2209,N_27660,N_29612);
or UO_2210 (O_2210,N_29136,N_29731);
and UO_2211 (O_2211,N_28076,N_28065);
or UO_2212 (O_2212,N_28294,N_28055);
xnor UO_2213 (O_2213,N_28302,N_27827);
and UO_2214 (O_2214,N_28710,N_28870);
nor UO_2215 (O_2215,N_28787,N_29573);
nor UO_2216 (O_2216,N_27636,N_27522);
or UO_2217 (O_2217,N_27776,N_28004);
xor UO_2218 (O_2218,N_28389,N_27682);
and UO_2219 (O_2219,N_27453,N_27473);
nor UO_2220 (O_2220,N_28714,N_28275);
nor UO_2221 (O_2221,N_29390,N_29572);
nor UO_2222 (O_2222,N_28111,N_29070);
and UO_2223 (O_2223,N_29487,N_27488);
and UO_2224 (O_2224,N_29849,N_27651);
nor UO_2225 (O_2225,N_28412,N_29139);
nor UO_2226 (O_2226,N_29164,N_28023);
or UO_2227 (O_2227,N_29104,N_27232);
nand UO_2228 (O_2228,N_29479,N_28752);
nand UO_2229 (O_2229,N_27117,N_27827);
xnor UO_2230 (O_2230,N_27050,N_29538);
or UO_2231 (O_2231,N_28119,N_27561);
nand UO_2232 (O_2232,N_28485,N_28997);
nor UO_2233 (O_2233,N_27696,N_29173);
or UO_2234 (O_2234,N_28056,N_29982);
xor UO_2235 (O_2235,N_27686,N_28193);
or UO_2236 (O_2236,N_29833,N_28173);
nor UO_2237 (O_2237,N_27700,N_28033);
or UO_2238 (O_2238,N_27965,N_28247);
or UO_2239 (O_2239,N_28278,N_29107);
and UO_2240 (O_2240,N_28028,N_28296);
xnor UO_2241 (O_2241,N_28019,N_29885);
nor UO_2242 (O_2242,N_28599,N_27071);
nor UO_2243 (O_2243,N_29421,N_28741);
xor UO_2244 (O_2244,N_29266,N_28278);
xnor UO_2245 (O_2245,N_27397,N_28550);
and UO_2246 (O_2246,N_27647,N_28253);
nand UO_2247 (O_2247,N_27706,N_28637);
and UO_2248 (O_2248,N_28252,N_29463);
nor UO_2249 (O_2249,N_28331,N_28224);
xor UO_2250 (O_2250,N_29966,N_28829);
xor UO_2251 (O_2251,N_28443,N_28512);
nor UO_2252 (O_2252,N_29002,N_27141);
or UO_2253 (O_2253,N_28807,N_28433);
and UO_2254 (O_2254,N_27673,N_29219);
or UO_2255 (O_2255,N_27579,N_27529);
or UO_2256 (O_2256,N_28755,N_28245);
nor UO_2257 (O_2257,N_27261,N_28937);
nor UO_2258 (O_2258,N_28792,N_27173);
nand UO_2259 (O_2259,N_29343,N_28844);
xor UO_2260 (O_2260,N_28963,N_28964);
nand UO_2261 (O_2261,N_28946,N_28646);
nor UO_2262 (O_2262,N_29948,N_29319);
and UO_2263 (O_2263,N_29215,N_29229);
or UO_2264 (O_2264,N_28445,N_27938);
nor UO_2265 (O_2265,N_29617,N_28275);
xor UO_2266 (O_2266,N_29627,N_27039);
nand UO_2267 (O_2267,N_27211,N_29591);
and UO_2268 (O_2268,N_28003,N_28183);
and UO_2269 (O_2269,N_29634,N_27057);
nor UO_2270 (O_2270,N_28596,N_29895);
xnor UO_2271 (O_2271,N_28874,N_29979);
nand UO_2272 (O_2272,N_27925,N_28147);
xnor UO_2273 (O_2273,N_27665,N_29854);
nand UO_2274 (O_2274,N_28063,N_28780);
nor UO_2275 (O_2275,N_27074,N_29868);
and UO_2276 (O_2276,N_28945,N_28272);
or UO_2277 (O_2277,N_29644,N_27542);
and UO_2278 (O_2278,N_27072,N_29973);
nand UO_2279 (O_2279,N_28278,N_27247);
xor UO_2280 (O_2280,N_29929,N_28717);
and UO_2281 (O_2281,N_28243,N_29687);
nor UO_2282 (O_2282,N_27442,N_28899);
nor UO_2283 (O_2283,N_27886,N_29635);
or UO_2284 (O_2284,N_29552,N_27536);
nand UO_2285 (O_2285,N_29314,N_28458);
nand UO_2286 (O_2286,N_29730,N_28981);
nor UO_2287 (O_2287,N_27367,N_28623);
and UO_2288 (O_2288,N_28486,N_29266);
nor UO_2289 (O_2289,N_28288,N_27519);
and UO_2290 (O_2290,N_28941,N_29437);
xor UO_2291 (O_2291,N_27240,N_28351);
or UO_2292 (O_2292,N_28171,N_28303);
nor UO_2293 (O_2293,N_28422,N_27942);
or UO_2294 (O_2294,N_28391,N_27102);
and UO_2295 (O_2295,N_27329,N_29927);
and UO_2296 (O_2296,N_28482,N_27167);
nor UO_2297 (O_2297,N_27151,N_29620);
nand UO_2298 (O_2298,N_27619,N_29779);
nor UO_2299 (O_2299,N_27006,N_27272);
nand UO_2300 (O_2300,N_28975,N_28626);
or UO_2301 (O_2301,N_29450,N_28067);
nor UO_2302 (O_2302,N_27778,N_27470);
nor UO_2303 (O_2303,N_29096,N_27225);
and UO_2304 (O_2304,N_29906,N_28600);
xor UO_2305 (O_2305,N_28873,N_27733);
xnor UO_2306 (O_2306,N_29796,N_28962);
nand UO_2307 (O_2307,N_29805,N_27849);
or UO_2308 (O_2308,N_29362,N_28766);
and UO_2309 (O_2309,N_29575,N_28517);
nand UO_2310 (O_2310,N_29825,N_29096);
nor UO_2311 (O_2311,N_27891,N_29867);
nand UO_2312 (O_2312,N_28461,N_29803);
and UO_2313 (O_2313,N_27686,N_28183);
xor UO_2314 (O_2314,N_27487,N_29588);
xor UO_2315 (O_2315,N_29576,N_29547);
nand UO_2316 (O_2316,N_29238,N_29898);
nor UO_2317 (O_2317,N_28257,N_29146);
xnor UO_2318 (O_2318,N_27157,N_27061);
and UO_2319 (O_2319,N_27901,N_27087);
or UO_2320 (O_2320,N_29536,N_27143);
nor UO_2321 (O_2321,N_27363,N_27268);
or UO_2322 (O_2322,N_27985,N_27446);
nand UO_2323 (O_2323,N_29151,N_28517);
and UO_2324 (O_2324,N_28641,N_28177);
nand UO_2325 (O_2325,N_29895,N_28325);
or UO_2326 (O_2326,N_29528,N_29867);
xor UO_2327 (O_2327,N_28283,N_28678);
nor UO_2328 (O_2328,N_28852,N_29616);
and UO_2329 (O_2329,N_29031,N_28962);
xor UO_2330 (O_2330,N_27073,N_29677);
and UO_2331 (O_2331,N_29868,N_27906);
or UO_2332 (O_2332,N_28192,N_28323);
and UO_2333 (O_2333,N_29060,N_28677);
nand UO_2334 (O_2334,N_29407,N_27704);
or UO_2335 (O_2335,N_27862,N_27001);
nor UO_2336 (O_2336,N_28516,N_27970);
nand UO_2337 (O_2337,N_27169,N_29165);
or UO_2338 (O_2338,N_27102,N_29224);
or UO_2339 (O_2339,N_29583,N_29537);
nor UO_2340 (O_2340,N_27619,N_29232);
or UO_2341 (O_2341,N_27933,N_29816);
and UO_2342 (O_2342,N_28277,N_28681);
and UO_2343 (O_2343,N_27068,N_29590);
or UO_2344 (O_2344,N_27420,N_28706);
or UO_2345 (O_2345,N_27623,N_28895);
xnor UO_2346 (O_2346,N_29454,N_27791);
nand UO_2347 (O_2347,N_28581,N_27381);
nor UO_2348 (O_2348,N_28834,N_29911);
nor UO_2349 (O_2349,N_27895,N_28913);
and UO_2350 (O_2350,N_27019,N_27439);
nor UO_2351 (O_2351,N_29813,N_28063);
or UO_2352 (O_2352,N_27616,N_27465);
xnor UO_2353 (O_2353,N_28185,N_28967);
xor UO_2354 (O_2354,N_28966,N_28594);
and UO_2355 (O_2355,N_27851,N_28916);
or UO_2356 (O_2356,N_28929,N_28592);
nor UO_2357 (O_2357,N_28065,N_27005);
xnor UO_2358 (O_2358,N_29086,N_27091);
or UO_2359 (O_2359,N_28540,N_28014);
xnor UO_2360 (O_2360,N_28372,N_29229);
xor UO_2361 (O_2361,N_29730,N_28271);
nor UO_2362 (O_2362,N_28996,N_29362);
or UO_2363 (O_2363,N_29906,N_28861);
xnor UO_2364 (O_2364,N_29590,N_28253);
or UO_2365 (O_2365,N_27223,N_29491);
or UO_2366 (O_2366,N_27173,N_28026);
or UO_2367 (O_2367,N_28973,N_28635);
xor UO_2368 (O_2368,N_29915,N_28269);
or UO_2369 (O_2369,N_29723,N_28544);
and UO_2370 (O_2370,N_29165,N_28252);
and UO_2371 (O_2371,N_29461,N_28564);
nand UO_2372 (O_2372,N_29394,N_27986);
or UO_2373 (O_2373,N_27782,N_29088);
nor UO_2374 (O_2374,N_29959,N_28228);
or UO_2375 (O_2375,N_28120,N_28345);
nand UO_2376 (O_2376,N_29802,N_28702);
or UO_2377 (O_2377,N_29535,N_27932);
nand UO_2378 (O_2378,N_27986,N_27285);
nor UO_2379 (O_2379,N_28110,N_29070);
xnor UO_2380 (O_2380,N_29159,N_29409);
nand UO_2381 (O_2381,N_29860,N_27456);
nor UO_2382 (O_2382,N_27259,N_27433);
nand UO_2383 (O_2383,N_28505,N_28210);
nor UO_2384 (O_2384,N_29958,N_28640);
xnor UO_2385 (O_2385,N_28275,N_28248);
or UO_2386 (O_2386,N_28551,N_29476);
nand UO_2387 (O_2387,N_28676,N_29791);
nor UO_2388 (O_2388,N_28528,N_28045);
and UO_2389 (O_2389,N_27672,N_29148);
and UO_2390 (O_2390,N_29833,N_27825);
or UO_2391 (O_2391,N_27565,N_28989);
and UO_2392 (O_2392,N_29865,N_29267);
and UO_2393 (O_2393,N_29825,N_29849);
and UO_2394 (O_2394,N_29946,N_27098);
and UO_2395 (O_2395,N_29340,N_28707);
xor UO_2396 (O_2396,N_28924,N_27315);
or UO_2397 (O_2397,N_27038,N_27231);
nor UO_2398 (O_2398,N_27999,N_27281);
or UO_2399 (O_2399,N_28410,N_27366);
nand UO_2400 (O_2400,N_28310,N_28955);
nor UO_2401 (O_2401,N_29435,N_28722);
and UO_2402 (O_2402,N_28475,N_29561);
and UO_2403 (O_2403,N_29579,N_28999);
and UO_2404 (O_2404,N_29921,N_29035);
and UO_2405 (O_2405,N_29518,N_28031);
and UO_2406 (O_2406,N_28524,N_29462);
nor UO_2407 (O_2407,N_28251,N_27255);
and UO_2408 (O_2408,N_28838,N_29662);
nor UO_2409 (O_2409,N_29062,N_28273);
and UO_2410 (O_2410,N_28415,N_28708);
xor UO_2411 (O_2411,N_28170,N_28107);
and UO_2412 (O_2412,N_28853,N_29249);
xor UO_2413 (O_2413,N_28280,N_27350);
or UO_2414 (O_2414,N_29036,N_27534);
or UO_2415 (O_2415,N_27731,N_27572);
and UO_2416 (O_2416,N_27946,N_27230);
xor UO_2417 (O_2417,N_27175,N_29656);
xnor UO_2418 (O_2418,N_27273,N_27812);
nand UO_2419 (O_2419,N_28393,N_29464);
nand UO_2420 (O_2420,N_29472,N_28580);
and UO_2421 (O_2421,N_28547,N_28467);
and UO_2422 (O_2422,N_28713,N_29191);
or UO_2423 (O_2423,N_28585,N_27118);
and UO_2424 (O_2424,N_27210,N_27845);
nand UO_2425 (O_2425,N_28493,N_28643);
nand UO_2426 (O_2426,N_27204,N_28130);
nand UO_2427 (O_2427,N_28107,N_27809);
xnor UO_2428 (O_2428,N_28505,N_27630);
nor UO_2429 (O_2429,N_29287,N_29407);
nor UO_2430 (O_2430,N_27996,N_27943);
nand UO_2431 (O_2431,N_28061,N_28501);
nand UO_2432 (O_2432,N_29782,N_28781);
or UO_2433 (O_2433,N_28667,N_29479);
or UO_2434 (O_2434,N_27892,N_27703);
or UO_2435 (O_2435,N_27636,N_27183);
xor UO_2436 (O_2436,N_28829,N_27726);
nand UO_2437 (O_2437,N_27528,N_27540);
and UO_2438 (O_2438,N_29528,N_29707);
xor UO_2439 (O_2439,N_27957,N_28213);
and UO_2440 (O_2440,N_29689,N_27728);
nor UO_2441 (O_2441,N_29662,N_29877);
nor UO_2442 (O_2442,N_28430,N_28968);
and UO_2443 (O_2443,N_28513,N_29340);
or UO_2444 (O_2444,N_28943,N_29151);
nor UO_2445 (O_2445,N_29406,N_29043);
or UO_2446 (O_2446,N_28228,N_29430);
and UO_2447 (O_2447,N_27063,N_29085);
or UO_2448 (O_2448,N_28066,N_28913);
nor UO_2449 (O_2449,N_29738,N_27538);
or UO_2450 (O_2450,N_27641,N_29313);
xnor UO_2451 (O_2451,N_28838,N_28074);
xor UO_2452 (O_2452,N_27307,N_29266);
xnor UO_2453 (O_2453,N_28823,N_28257);
xor UO_2454 (O_2454,N_29884,N_28403);
nor UO_2455 (O_2455,N_27586,N_29416);
and UO_2456 (O_2456,N_27504,N_28355);
or UO_2457 (O_2457,N_27089,N_28399);
xnor UO_2458 (O_2458,N_28048,N_28204);
and UO_2459 (O_2459,N_28843,N_29069);
nor UO_2460 (O_2460,N_28810,N_29909);
nand UO_2461 (O_2461,N_29931,N_28028);
nor UO_2462 (O_2462,N_27426,N_29436);
nand UO_2463 (O_2463,N_27467,N_29044);
nand UO_2464 (O_2464,N_27078,N_27988);
nand UO_2465 (O_2465,N_27106,N_27100);
nor UO_2466 (O_2466,N_28876,N_27041);
nand UO_2467 (O_2467,N_28430,N_28063);
nand UO_2468 (O_2468,N_27722,N_28187);
and UO_2469 (O_2469,N_28374,N_27791);
xnor UO_2470 (O_2470,N_29322,N_27933);
nand UO_2471 (O_2471,N_29555,N_28665);
nand UO_2472 (O_2472,N_28902,N_28479);
nand UO_2473 (O_2473,N_27667,N_29624);
nand UO_2474 (O_2474,N_29170,N_27115);
nor UO_2475 (O_2475,N_27061,N_29201);
and UO_2476 (O_2476,N_28337,N_28387);
or UO_2477 (O_2477,N_27814,N_28176);
xor UO_2478 (O_2478,N_28118,N_29639);
nand UO_2479 (O_2479,N_27123,N_28729);
and UO_2480 (O_2480,N_27855,N_28309);
nand UO_2481 (O_2481,N_29042,N_27423);
or UO_2482 (O_2482,N_27393,N_28127);
nor UO_2483 (O_2483,N_27754,N_28392);
nor UO_2484 (O_2484,N_29275,N_28052);
nand UO_2485 (O_2485,N_28221,N_29273);
nand UO_2486 (O_2486,N_29958,N_28646);
or UO_2487 (O_2487,N_27739,N_29342);
or UO_2488 (O_2488,N_28086,N_27258);
or UO_2489 (O_2489,N_28952,N_29619);
nor UO_2490 (O_2490,N_28903,N_28687);
xnor UO_2491 (O_2491,N_29731,N_27094);
and UO_2492 (O_2492,N_27870,N_28487);
nand UO_2493 (O_2493,N_28836,N_29731);
or UO_2494 (O_2494,N_27736,N_28578);
or UO_2495 (O_2495,N_28871,N_27354);
nand UO_2496 (O_2496,N_28663,N_28866);
xnor UO_2497 (O_2497,N_29031,N_29951);
or UO_2498 (O_2498,N_29150,N_29492);
or UO_2499 (O_2499,N_27124,N_29748);
or UO_2500 (O_2500,N_27720,N_27990);
or UO_2501 (O_2501,N_29499,N_27929);
xor UO_2502 (O_2502,N_27104,N_29455);
and UO_2503 (O_2503,N_29967,N_28800);
nand UO_2504 (O_2504,N_27664,N_28542);
and UO_2505 (O_2505,N_29283,N_29686);
and UO_2506 (O_2506,N_28219,N_27604);
and UO_2507 (O_2507,N_28109,N_27996);
and UO_2508 (O_2508,N_27198,N_27418);
nand UO_2509 (O_2509,N_29883,N_28001);
and UO_2510 (O_2510,N_28920,N_29109);
nand UO_2511 (O_2511,N_28073,N_29289);
nor UO_2512 (O_2512,N_29824,N_29969);
or UO_2513 (O_2513,N_29654,N_28412);
or UO_2514 (O_2514,N_27368,N_27474);
and UO_2515 (O_2515,N_29108,N_28848);
and UO_2516 (O_2516,N_27974,N_28041);
and UO_2517 (O_2517,N_29246,N_28337);
nor UO_2518 (O_2518,N_28295,N_28518);
nor UO_2519 (O_2519,N_29398,N_28261);
nor UO_2520 (O_2520,N_28188,N_28998);
nor UO_2521 (O_2521,N_27789,N_27661);
xnor UO_2522 (O_2522,N_28543,N_29473);
or UO_2523 (O_2523,N_29638,N_29836);
xor UO_2524 (O_2524,N_28529,N_27956);
or UO_2525 (O_2525,N_28405,N_28726);
nor UO_2526 (O_2526,N_29416,N_28382);
or UO_2527 (O_2527,N_28309,N_28513);
nand UO_2528 (O_2528,N_28416,N_27758);
nand UO_2529 (O_2529,N_28695,N_27751);
nand UO_2530 (O_2530,N_28721,N_29863);
nor UO_2531 (O_2531,N_29932,N_29552);
nor UO_2532 (O_2532,N_29104,N_29874);
or UO_2533 (O_2533,N_27130,N_29229);
nand UO_2534 (O_2534,N_27357,N_28826);
xor UO_2535 (O_2535,N_28639,N_28220);
or UO_2536 (O_2536,N_27260,N_28064);
nand UO_2537 (O_2537,N_27992,N_27343);
nand UO_2538 (O_2538,N_29648,N_28870);
nor UO_2539 (O_2539,N_28817,N_29729);
nor UO_2540 (O_2540,N_28379,N_29197);
and UO_2541 (O_2541,N_29156,N_28357);
nand UO_2542 (O_2542,N_27637,N_28156);
or UO_2543 (O_2543,N_29265,N_29683);
nor UO_2544 (O_2544,N_28777,N_27647);
nand UO_2545 (O_2545,N_27091,N_29123);
nor UO_2546 (O_2546,N_29688,N_27009);
nand UO_2547 (O_2547,N_27899,N_28406);
xor UO_2548 (O_2548,N_28396,N_29800);
xor UO_2549 (O_2549,N_29856,N_29842);
xor UO_2550 (O_2550,N_27580,N_27492);
xor UO_2551 (O_2551,N_29762,N_29616);
nor UO_2552 (O_2552,N_27486,N_28671);
and UO_2553 (O_2553,N_28425,N_28763);
and UO_2554 (O_2554,N_27930,N_27061);
nand UO_2555 (O_2555,N_29653,N_28426);
and UO_2556 (O_2556,N_29974,N_29722);
and UO_2557 (O_2557,N_27014,N_28101);
and UO_2558 (O_2558,N_27961,N_29239);
xnor UO_2559 (O_2559,N_28164,N_27709);
or UO_2560 (O_2560,N_29654,N_27055);
or UO_2561 (O_2561,N_27271,N_28362);
nand UO_2562 (O_2562,N_28067,N_27706);
nand UO_2563 (O_2563,N_29112,N_27049);
nand UO_2564 (O_2564,N_29938,N_27828);
or UO_2565 (O_2565,N_28877,N_28100);
and UO_2566 (O_2566,N_29258,N_29589);
nand UO_2567 (O_2567,N_29766,N_29500);
nand UO_2568 (O_2568,N_29466,N_27969);
xor UO_2569 (O_2569,N_29938,N_27236);
and UO_2570 (O_2570,N_29928,N_27649);
nor UO_2571 (O_2571,N_27514,N_27622);
xor UO_2572 (O_2572,N_28586,N_28765);
nor UO_2573 (O_2573,N_28277,N_27715);
nand UO_2574 (O_2574,N_27890,N_29164);
xnor UO_2575 (O_2575,N_29136,N_29710);
nor UO_2576 (O_2576,N_29678,N_28672);
and UO_2577 (O_2577,N_27313,N_28217);
or UO_2578 (O_2578,N_27046,N_27336);
or UO_2579 (O_2579,N_29184,N_29664);
nand UO_2580 (O_2580,N_28765,N_28585);
or UO_2581 (O_2581,N_27238,N_27175);
xnor UO_2582 (O_2582,N_29003,N_27633);
and UO_2583 (O_2583,N_27768,N_29426);
xnor UO_2584 (O_2584,N_27122,N_28428);
nand UO_2585 (O_2585,N_27940,N_27267);
and UO_2586 (O_2586,N_28647,N_27041);
nand UO_2587 (O_2587,N_29057,N_28344);
xor UO_2588 (O_2588,N_28359,N_29665);
and UO_2589 (O_2589,N_29261,N_27079);
and UO_2590 (O_2590,N_27005,N_29556);
nand UO_2591 (O_2591,N_27733,N_27260);
nor UO_2592 (O_2592,N_29595,N_28987);
xnor UO_2593 (O_2593,N_27897,N_28975);
and UO_2594 (O_2594,N_27284,N_28828);
or UO_2595 (O_2595,N_28728,N_28326);
and UO_2596 (O_2596,N_29712,N_28952);
nor UO_2597 (O_2597,N_29400,N_28474);
and UO_2598 (O_2598,N_28170,N_28570);
or UO_2599 (O_2599,N_27379,N_29181);
nor UO_2600 (O_2600,N_29773,N_28262);
nor UO_2601 (O_2601,N_28450,N_28514);
nand UO_2602 (O_2602,N_27194,N_27392);
or UO_2603 (O_2603,N_29325,N_29096);
nor UO_2604 (O_2604,N_29229,N_29947);
and UO_2605 (O_2605,N_27875,N_27708);
nand UO_2606 (O_2606,N_29393,N_27799);
xnor UO_2607 (O_2607,N_27890,N_28528);
or UO_2608 (O_2608,N_28190,N_29482);
nand UO_2609 (O_2609,N_29333,N_27022);
xnor UO_2610 (O_2610,N_29750,N_29024);
nor UO_2611 (O_2611,N_29767,N_27508);
nand UO_2612 (O_2612,N_27155,N_27806);
nor UO_2613 (O_2613,N_29898,N_29659);
nand UO_2614 (O_2614,N_28787,N_27062);
nor UO_2615 (O_2615,N_29545,N_29655);
nor UO_2616 (O_2616,N_27067,N_29326);
and UO_2617 (O_2617,N_27711,N_27353);
and UO_2618 (O_2618,N_29485,N_27457);
or UO_2619 (O_2619,N_29288,N_28399);
xor UO_2620 (O_2620,N_28278,N_29458);
nor UO_2621 (O_2621,N_28217,N_29720);
nor UO_2622 (O_2622,N_29372,N_29238);
or UO_2623 (O_2623,N_29691,N_29278);
or UO_2624 (O_2624,N_29838,N_28507);
nor UO_2625 (O_2625,N_29976,N_29824);
and UO_2626 (O_2626,N_29074,N_27844);
xor UO_2627 (O_2627,N_28963,N_28999);
nor UO_2628 (O_2628,N_29854,N_28508);
nor UO_2629 (O_2629,N_29068,N_28331);
nor UO_2630 (O_2630,N_27752,N_27649);
and UO_2631 (O_2631,N_27741,N_29951);
nand UO_2632 (O_2632,N_29891,N_29378);
nor UO_2633 (O_2633,N_28430,N_27617);
nor UO_2634 (O_2634,N_27273,N_28452);
nand UO_2635 (O_2635,N_27750,N_28162);
and UO_2636 (O_2636,N_28522,N_28094);
and UO_2637 (O_2637,N_29751,N_29465);
or UO_2638 (O_2638,N_27649,N_29074);
xor UO_2639 (O_2639,N_27856,N_27298);
nand UO_2640 (O_2640,N_27126,N_27727);
nand UO_2641 (O_2641,N_29228,N_27301);
nand UO_2642 (O_2642,N_29168,N_28228);
xor UO_2643 (O_2643,N_28291,N_29807);
xor UO_2644 (O_2644,N_27801,N_28219);
and UO_2645 (O_2645,N_27587,N_27105);
or UO_2646 (O_2646,N_27648,N_28650);
or UO_2647 (O_2647,N_27789,N_27386);
nor UO_2648 (O_2648,N_29569,N_28175);
and UO_2649 (O_2649,N_27791,N_27452);
or UO_2650 (O_2650,N_28719,N_29738);
xor UO_2651 (O_2651,N_29438,N_28198);
nand UO_2652 (O_2652,N_27455,N_29874);
xnor UO_2653 (O_2653,N_27454,N_28251);
xor UO_2654 (O_2654,N_28130,N_27747);
or UO_2655 (O_2655,N_28324,N_27519);
and UO_2656 (O_2656,N_27242,N_28755);
xor UO_2657 (O_2657,N_29443,N_27834);
or UO_2658 (O_2658,N_29943,N_27589);
nor UO_2659 (O_2659,N_27303,N_28662);
and UO_2660 (O_2660,N_27929,N_29681);
and UO_2661 (O_2661,N_29833,N_29652);
xnor UO_2662 (O_2662,N_28587,N_28083);
nor UO_2663 (O_2663,N_29654,N_27794);
or UO_2664 (O_2664,N_28548,N_28719);
and UO_2665 (O_2665,N_27808,N_28869);
nand UO_2666 (O_2666,N_27463,N_28773);
nand UO_2667 (O_2667,N_27496,N_28084);
and UO_2668 (O_2668,N_28776,N_29959);
nand UO_2669 (O_2669,N_27476,N_28834);
or UO_2670 (O_2670,N_28134,N_27687);
nor UO_2671 (O_2671,N_29068,N_29872);
nand UO_2672 (O_2672,N_29688,N_27968);
and UO_2673 (O_2673,N_28673,N_27987);
xnor UO_2674 (O_2674,N_28527,N_29591);
nor UO_2675 (O_2675,N_27452,N_27913);
xnor UO_2676 (O_2676,N_29598,N_27391);
and UO_2677 (O_2677,N_29896,N_29478);
xnor UO_2678 (O_2678,N_27216,N_29339);
and UO_2679 (O_2679,N_28395,N_29056);
nor UO_2680 (O_2680,N_27335,N_27722);
nor UO_2681 (O_2681,N_29567,N_29963);
nand UO_2682 (O_2682,N_29636,N_27859);
nand UO_2683 (O_2683,N_29221,N_27170);
and UO_2684 (O_2684,N_27330,N_27574);
nor UO_2685 (O_2685,N_27228,N_27355);
or UO_2686 (O_2686,N_29438,N_29464);
nor UO_2687 (O_2687,N_28346,N_28619);
nor UO_2688 (O_2688,N_27500,N_28831);
nand UO_2689 (O_2689,N_29298,N_29026);
and UO_2690 (O_2690,N_27784,N_29123);
and UO_2691 (O_2691,N_27073,N_28880);
or UO_2692 (O_2692,N_29585,N_29041);
nor UO_2693 (O_2693,N_28298,N_27088);
or UO_2694 (O_2694,N_29785,N_28056);
nor UO_2695 (O_2695,N_29863,N_29280);
nand UO_2696 (O_2696,N_27987,N_27885);
nor UO_2697 (O_2697,N_28879,N_27246);
nand UO_2698 (O_2698,N_29075,N_28522);
nand UO_2699 (O_2699,N_28965,N_28984);
and UO_2700 (O_2700,N_28051,N_29906);
nand UO_2701 (O_2701,N_29204,N_28776);
or UO_2702 (O_2702,N_27471,N_29874);
or UO_2703 (O_2703,N_29886,N_28137);
nand UO_2704 (O_2704,N_28573,N_27518);
nor UO_2705 (O_2705,N_27398,N_29172);
or UO_2706 (O_2706,N_29830,N_27146);
xnor UO_2707 (O_2707,N_27823,N_28124);
nand UO_2708 (O_2708,N_27904,N_29612);
or UO_2709 (O_2709,N_29850,N_29433);
nand UO_2710 (O_2710,N_29364,N_29134);
nand UO_2711 (O_2711,N_28556,N_27001);
xnor UO_2712 (O_2712,N_29922,N_28289);
and UO_2713 (O_2713,N_27123,N_29033);
and UO_2714 (O_2714,N_28920,N_28233);
or UO_2715 (O_2715,N_29469,N_27802);
xor UO_2716 (O_2716,N_28688,N_28509);
or UO_2717 (O_2717,N_28354,N_28781);
nor UO_2718 (O_2718,N_28758,N_27147);
and UO_2719 (O_2719,N_28857,N_29470);
nor UO_2720 (O_2720,N_29662,N_29502);
nor UO_2721 (O_2721,N_29430,N_27306);
xnor UO_2722 (O_2722,N_27272,N_28063);
and UO_2723 (O_2723,N_27461,N_27723);
or UO_2724 (O_2724,N_27492,N_29336);
and UO_2725 (O_2725,N_27921,N_27677);
xor UO_2726 (O_2726,N_27707,N_28281);
or UO_2727 (O_2727,N_27961,N_27553);
or UO_2728 (O_2728,N_28534,N_28806);
nor UO_2729 (O_2729,N_27623,N_27107);
and UO_2730 (O_2730,N_29968,N_27230);
and UO_2731 (O_2731,N_29182,N_27412);
xnor UO_2732 (O_2732,N_28783,N_29515);
nor UO_2733 (O_2733,N_28940,N_27040);
xnor UO_2734 (O_2734,N_29818,N_29752);
xor UO_2735 (O_2735,N_29894,N_28317);
and UO_2736 (O_2736,N_27569,N_29974);
nor UO_2737 (O_2737,N_27168,N_29834);
and UO_2738 (O_2738,N_27569,N_27259);
and UO_2739 (O_2739,N_27924,N_28542);
nand UO_2740 (O_2740,N_27774,N_29585);
xnor UO_2741 (O_2741,N_28944,N_29594);
or UO_2742 (O_2742,N_28706,N_28552);
or UO_2743 (O_2743,N_29791,N_27245);
and UO_2744 (O_2744,N_27362,N_28083);
and UO_2745 (O_2745,N_27620,N_27163);
or UO_2746 (O_2746,N_28487,N_27252);
and UO_2747 (O_2747,N_29934,N_29897);
nand UO_2748 (O_2748,N_29749,N_28499);
nand UO_2749 (O_2749,N_28325,N_29397);
and UO_2750 (O_2750,N_28028,N_29777);
nor UO_2751 (O_2751,N_27591,N_29815);
nor UO_2752 (O_2752,N_28106,N_29545);
nand UO_2753 (O_2753,N_27038,N_27503);
and UO_2754 (O_2754,N_28653,N_27344);
or UO_2755 (O_2755,N_27737,N_28099);
and UO_2756 (O_2756,N_29165,N_28673);
nor UO_2757 (O_2757,N_27034,N_28555);
and UO_2758 (O_2758,N_27266,N_29336);
nor UO_2759 (O_2759,N_29303,N_27606);
xnor UO_2760 (O_2760,N_27695,N_28400);
or UO_2761 (O_2761,N_27695,N_29989);
or UO_2762 (O_2762,N_29379,N_27822);
and UO_2763 (O_2763,N_28689,N_29765);
nand UO_2764 (O_2764,N_28184,N_29505);
xor UO_2765 (O_2765,N_29761,N_27976);
and UO_2766 (O_2766,N_28930,N_27665);
and UO_2767 (O_2767,N_29398,N_29564);
nor UO_2768 (O_2768,N_29864,N_29384);
or UO_2769 (O_2769,N_28334,N_29077);
nand UO_2770 (O_2770,N_27372,N_28963);
nand UO_2771 (O_2771,N_27763,N_28764);
xnor UO_2772 (O_2772,N_27869,N_28066);
nor UO_2773 (O_2773,N_27341,N_29313);
xnor UO_2774 (O_2774,N_28098,N_27906);
nand UO_2775 (O_2775,N_28901,N_28725);
nand UO_2776 (O_2776,N_29228,N_27660);
or UO_2777 (O_2777,N_29623,N_28476);
xor UO_2778 (O_2778,N_28605,N_28421);
and UO_2779 (O_2779,N_28601,N_27257);
or UO_2780 (O_2780,N_27833,N_28221);
nand UO_2781 (O_2781,N_27355,N_28605);
or UO_2782 (O_2782,N_29147,N_28759);
nor UO_2783 (O_2783,N_29789,N_29102);
xor UO_2784 (O_2784,N_29687,N_29080);
and UO_2785 (O_2785,N_28112,N_28525);
nor UO_2786 (O_2786,N_28528,N_28224);
or UO_2787 (O_2787,N_27830,N_27241);
xnor UO_2788 (O_2788,N_27756,N_27016);
xnor UO_2789 (O_2789,N_29960,N_29384);
xnor UO_2790 (O_2790,N_27819,N_28077);
and UO_2791 (O_2791,N_27544,N_29160);
and UO_2792 (O_2792,N_28734,N_28428);
xor UO_2793 (O_2793,N_28464,N_29101);
xnor UO_2794 (O_2794,N_28961,N_28589);
or UO_2795 (O_2795,N_29540,N_28731);
nor UO_2796 (O_2796,N_29416,N_29256);
nor UO_2797 (O_2797,N_29322,N_29950);
xnor UO_2798 (O_2798,N_29491,N_29519);
or UO_2799 (O_2799,N_29380,N_27656);
and UO_2800 (O_2800,N_29379,N_29410);
and UO_2801 (O_2801,N_29378,N_28314);
and UO_2802 (O_2802,N_27190,N_28768);
and UO_2803 (O_2803,N_29389,N_27073);
xnor UO_2804 (O_2804,N_27339,N_27970);
and UO_2805 (O_2805,N_28472,N_28987);
or UO_2806 (O_2806,N_29290,N_27984);
or UO_2807 (O_2807,N_27814,N_27402);
and UO_2808 (O_2808,N_27307,N_27787);
or UO_2809 (O_2809,N_28914,N_28511);
nor UO_2810 (O_2810,N_29882,N_28569);
nor UO_2811 (O_2811,N_29193,N_27794);
and UO_2812 (O_2812,N_27654,N_28464);
xnor UO_2813 (O_2813,N_28191,N_29878);
nand UO_2814 (O_2814,N_29035,N_29081);
xnor UO_2815 (O_2815,N_27248,N_28403);
or UO_2816 (O_2816,N_29211,N_27309);
xor UO_2817 (O_2817,N_27687,N_28251);
and UO_2818 (O_2818,N_27803,N_28936);
nor UO_2819 (O_2819,N_27771,N_29502);
nor UO_2820 (O_2820,N_28608,N_29121);
or UO_2821 (O_2821,N_28786,N_27040);
or UO_2822 (O_2822,N_28491,N_27241);
and UO_2823 (O_2823,N_28307,N_29543);
nor UO_2824 (O_2824,N_28823,N_29836);
xor UO_2825 (O_2825,N_29326,N_28290);
xnor UO_2826 (O_2826,N_29032,N_28178);
xnor UO_2827 (O_2827,N_29045,N_27832);
xor UO_2828 (O_2828,N_29213,N_28438);
or UO_2829 (O_2829,N_29989,N_28411);
or UO_2830 (O_2830,N_28101,N_27402);
or UO_2831 (O_2831,N_27614,N_29617);
nand UO_2832 (O_2832,N_27402,N_28228);
and UO_2833 (O_2833,N_27543,N_29273);
or UO_2834 (O_2834,N_28225,N_27477);
and UO_2835 (O_2835,N_28453,N_27760);
xnor UO_2836 (O_2836,N_29238,N_27628);
nor UO_2837 (O_2837,N_28909,N_28610);
nand UO_2838 (O_2838,N_29029,N_28067);
and UO_2839 (O_2839,N_29361,N_27032);
or UO_2840 (O_2840,N_29282,N_28662);
nand UO_2841 (O_2841,N_27985,N_28792);
and UO_2842 (O_2842,N_28158,N_27109);
or UO_2843 (O_2843,N_27172,N_29142);
and UO_2844 (O_2844,N_27559,N_29819);
or UO_2845 (O_2845,N_27292,N_27294);
and UO_2846 (O_2846,N_27971,N_27285);
nor UO_2847 (O_2847,N_29972,N_29742);
xnor UO_2848 (O_2848,N_28159,N_28441);
or UO_2849 (O_2849,N_27302,N_29310);
nand UO_2850 (O_2850,N_27686,N_27340);
nor UO_2851 (O_2851,N_27639,N_27702);
and UO_2852 (O_2852,N_28767,N_28670);
xnor UO_2853 (O_2853,N_28181,N_28365);
or UO_2854 (O_2854,N_27790,N_28252);
nor UO_2855 (O_2855,N_28534,N_29284);
nor UO_2856 (O_2856,N_29253,N_29331);
nor UO_2857 (O_2857,N_28844,N_27311);
nor UO_2858 (O_2858,N_29532,N_27543);
and UO_2859 (O_2859,N_27012,N_27875);
nand UO_2860 (O_2860,N_29758,N_28066);
xnor UO_2861 (O_2861,N_29760,N_27210);
or UO_2862 (O_2862,N_27773,N_28143);
or UO_2863 (O_2863,N_27504,N_27020);
xnor UO_2864 (O_2864,N_28860,N_29533);
or UO_2865 (O_2865,N_28051,N_29410);
xnor UO_2866 (O_2866,N_28751,N_29032);
or UO_2867 (O_2867,N_28469,N_27879);
nand UO_2868 (O_2868,N_28318,N_29419);
nor UO_2869 (O_2869,N_28057,N_28433);
nor UO_2870 (O_2870,N_28667,N_28418);
nand UO_2871 (O_2871,N_27916,N_29143);
xor UO_2872 (O_2872,N_28031,N_29889);
or UO_2873 (O_2873,N_27711,N_28313);
xnor UO_2874 (O_2874,N_28260,N_27592);
nand UO_2875 (O_2875,N_29763,N_29877);
xor UO_2876 (O_2876,N_27827,N_27770);
and UO_2877 (O_2877,N_27901,N_29823);
or UO_2878 (O_2878,N_28407,N_27750);
or UO_2879 (O_2879,N_29747,N_28993);
nor UO_2880 (O_2880,N_27055,N_29397);
nor UO_2881 (O_2881,N_27502,N_29387);
nor UO_2882 (O_2882,N_27047,N_27352);
nand UO_2883 (O_2883,N_27851,N_27768);
and UO_2884 (O_2884,N_27700,N_28611);
nand UO_2885 (O_2885,N_27591,N_28253);
nand UO_2886 (O_2886,N_27453,N_28608);
nand UO_2887 (O_2887,N_28131,N_27255);
or UO_2888 (O_2888,N_28466,N_27319);
nor UO_2889 (O_2889,N_29890,N_28754);
nor UO_2890 (O_2890,N_28427,N_28140);
or UO_2891 (O_2891,N_29871,N_27046);
nand UO_2892 (O_2892,N_28490,N_27469);
and UO_2893 (O_2893,N_27721,N_27620);
nor UO_2894 (O_2894,N_27533,N_29047);
nor UO_2895 (O_2895,N_29379,N_29494);
xnor UO_2896 (O_2896,N_28144,N_27117);
or UO_2897 (O_2897,N_29322,N_28427);
and UO_2898 (O_2898,N_29028,N_28124);
nor UO_2899 (O_2899,N_27857,N_27233);
nand UO_2900 (O_2900,N_27380,N_27246);
nor UO_2901 (O_2901,N_28244,N_29734);
or UO_2902 (O_2902,N_27485,N_27641);
nor UO_2903 (O_2903,N_27999,N_27427);
or UO_2904 (O_2904,N_27851,N_27579);
nand UO_2905 (O_2905,N_28336,N_29892);
nand UO_2906 (O_2906,N_28886,N_27791);
and UO_2907 (O_2907,N_28516,N_28889);
xor UO_2908 (O_2908,N_27514,N_29445);
or UO_2909 (O_2909,N_28492,N_28284);
nand UO_2910 (O_2910,N_29987,N_29396);
nor UO_2911 (O_2911,N_29037,N_27515);
and UO_2912 (O_2912,N_27773,N_27024);
nor UO_2913 (O_2913,N_27298,N_29448);
or UO_2914 (O_2914,N_29772,N_27249);
xnor UO_2915 (O_2915,N_29894,N_27022);
nand UO_2916 (O_2916,N_29516,N_27157);
xnor UO_2917 (O_2917,N_29902,N_29944);
xnor UO_2918 (O_2918,N_28309,N_27610);
and UO_2919 (O_2919,N_27508,N_27919);
or UO_2920 (O_2920,N_29767,N_28500);
xor UO_2921 (O_2921,N_29893,N_29246);
and UO_2922 (O_2922,N_29153,N_29790);
nor UO_2923 (O_2923,N_29383,N_28678);
nor UO_2924 (O_2924,N_29242,N_29813);
and UO_2925 (O_2925,N_29615,N_27561);
nand UO_2926 (O_2926,N_27576,N_28717);
or UO_2927 (O_2927,N_28930,N_27363);
or UO_2928 (O_2928,N_29908,N_28510);
xor UO_2929 (O_2929,N_27126,N_29359);
xnor UO_2930 (O_2930,N_29689,N_28053);
nor UO_2931 (O_2931,N_28460,N_27946);
nand UO_2932 (O_2932,N_27181,N_28804);
xor UO_2933 (O_2933,N_29950,N_29126);
and UO_2934 (O_2934,N_29484,N_27184);
and UO_2935 (O_2935,N_27737,N_27615);
xnor UO_2936 (O_2936,N_27357,N_28182);
nand UO_2937 (O_2937,N_29251,N_27270);
xor UO_2938 (O_2938,N_28782,N_29639);
or UO_2939 (O_2939,N_28045,N_29674);
and UO_2940 (O_2940,N_27989,N_29593);
nor UO_2941 (O_2941,N_29639,N_28379);
or UO_2942 (O_2942,N_28792,N_28754);
or UO_2943 (O_2943,N_29638,N_28895);
nand UO_2944 (O_2944,N_28363,N_29863);
nand UO_2945 (O_2945,N_28029,N_28886);
xnor UO_2946 (O_2946,N_27780,N_29249);
or UO_2947 (O_2947,N_28066,N_28250);
nor UO_2948 (O_2948,N_28678,N_27672);
nor UO_2949 (O_2949,N_28169,N_28841);
xnor UO_2950 (O_2950,N_28650,N_27811);
nand UO_2951 (O_2951,N_27188,N_28996);
or UO_2952 (O_2952,N_29986,N_29287);
nand UO_2953 (O_2953,N_29004,N_27615);
nor UO_2954 (O_2954,N_29533,N_27096);
nor UO_2955 (O_2955,N_29204,N_27989);
and UO_2956 (O_2956,N_27217,N_27740);
xnor UO_2957 (O_2957,N_28655,N_29348);
nand UO_2958 (O_2958,N_28549,N_28284);
xor UO_2959 (O_2959,N_28537,N_29542);
xnor UO_2960 (O_2960,N_28460,N_27413);
and UO_2961 (O_2961,N_28054,N_27832);
and UO_2962 (O_2962,N_28622,N_29087);
nand UO_2963 (O_2963,N_27180,N_27675);
nand UO_2964 (O_2964,N_28032,N_27235);
and UO_2965 (O_2965,N_27046,N_29016);
and UO_2966 (O_2966,N_27277,N_29575);
or UO_2967 (O_2967,N_27373,N_28935);
nand UO_2968 (O_2968,N_29747,N_28931);
nand UO_2969 (O_2969,N_27377,N_28630);
xnor UO_2970 (O_2970,N_27117,N_28949);
nor UO_2971 (O_2971,N_29532,N_27716);
and UO_2972 (O_2972,N_27277,N_27850);
or UO_2973 (O_2973,N_27973,N_28307);
or UO_2974 (O_2974,N_28569,N_27867);
nor UO_2975 (O_2975,N_28017,N_28536);
or UO_2976 (O_2976,N_28043,N_29303);
or UO_2977 (O_2977,N_27921,N_28806);
and UO_2978 (O_2978,N_28958,N_28904);
nor UO_2979 (O_2979,N_29792,N_28652);
nand UO_2980 (O_2980,N_29470,N_28765);
xor UO_2981 (O_2981,N_27921,N_27086);
nor UO_2982 (O_2982,N_28810,N_29636);
or UO_2983 (O_2983,N_29801,N_28457);
and UO_2984 (O_2984,N_29005,N_28492);
nor UO_2985 (O_2985,N_28247,N_28531);
or UO_2986 (O_2986,N_27461,N_28063);
or UO_2987 (O_2987,N_27890,N_28663);
nand UO_2988 (O_2988,N_28067,N_27133);
xnor UO_2989 (O_2989,N_28536,N_29342);
nor UO_2990 (O_2990,N_28665,N_29995);
or UO_2991 (O_2991,N_29942,N_27041);
nor UO_2992 (O_2992,N_28065,N_28710);
xor UO_2993 (O_2993,N_27187,N_28312);
nand UO_2994 (O_2994,N_28268,N_27521);
and UO_2995 (O_2995,N_29078,N_28474);
nor UO_2996 (O_2996,N_29787,N_29758);
xor UO_2997 (O_2997,N_28703,N_29386);
xor UO_2998 (O_2998,N_29581,N_29945);
or UO_2999 (O_2999,N_27077,N_28414);
nor UO_3000 (O_3000,N_28821,N_29492);
nor UO_3001 (O_3001,N_28894,N_27428);
nand UO_3002 (O_3002,N_27198,N_29839);
and UO_3003 (O_3003,N_27823,N_29405);
or UO_3004 (O_3004,N_27713,N_29199);
xor UO_3005 (O_3005,N_27045,N_28871);
or UO_3006 (O_3006,N_27783,N_28479);
or UO_3007 (O_3007,N_28660,N_29829);
xnor UO_3008 (O_3008,N_28008,N_28026);
xnor UO_3009 (O_3009,N_28037,N_27007);
nor UO_3010 (O_3010,N_27334,N_29055);
and UO_3011 (O_3011,N_29964,N_28222);
nand UO_3012 (O_3012,N_28933,N_27187);
xnor UO_3013 (O_3013,N_27344,N_28136);
nand UO_3014 (O_3014,N_27097,N_27209);
xor UO_3015 (O_3015,N_28180,N_29289);
or UO_3016 (O_3016,N_28381,N_27735);
xor UO_3017 (O_3017,N_29832,N_27739);
nor UO_3018 (O_3018,N_28588,N_27599);
nand UO_3019 (O_3019,N_27318,N_28225);
or UO_3020 (O_3020,N_27115,N_28533);
or UO_3021 (O_3021,N_29306,N_28819);
nand UO_3022 (O_3022,N_29282,N_27720);
xor UO_3023 (O_3023,N_29497,N_28060);
nand UO_3024 (O_3024,N_28489,N_28681);
or UO_3025 (O_3025,N_28411,N_28202);
nand UO_3026 (O_3026,N_27226,N_29441);
and UO_3027 (O_3027,N_28970,N_28050);
xor UO_3028 (O_3028,N_27169,N_28315);
or UO_3029 (O_3029,N_29074,N_27997);
nor UO_3030 (O_3030,N_28380,N_29996);
or UO_3031 (O_3031,N_28624,N_28918);
nand UO_3032 (O_3032,N_28648,N_29849);
nor UO_3033 (O_3033,N_28534,N_28178);
and UO_3034 (O_3034,N_27073,N_27049);
and UO_3035 (O_3035,N_27747,N_27783);
or UO_3036 (O_3036,N_27240,N_29146);
nand UO_3037 (O_3037,N_28140,N_28188);
and UO_3038 (O_3038,N_29703,N_28029);
nand UO_3039 (O_3039,N_29564,N_27929);
nand UO_3040 (O_3040,N_28931,N_29535);
and UO_3041 (O_3041,N_27473,N_28788);
and UO_3042 (O_3042,N_29649,N_28815);
xnor UO_3043 (O_3043,N_28670,N_29339);
and UO_3044 (O_3044,N_29860,N_28325);
nor UO_3045 (O_3045,N_27384,N_28405);
nand UO_3046 (O_3046,N_27669,N_29397);
nand UO_3047 (O_3047,N_28107,N_29591);
or UO_3048 (O_3048,N_28108,N_27478);
or UO_3049 (O_3049,N_29706,N_29707);
nor UO_3050 (O_3050,N_29394,N_27985);
nand UO_3051 (O_3051,N_29957,N_28741);
nor UO_3052 (O_3052,N_27663,N_27574);
nor UO_3053 (O_3053,N_29931,N_28867);
xnor UO_3054 (O_3054,N_29256,N_29985);
and UO_3055 (O_3055,N_27335,N_27739);
nor UO_3056 (O_3056,N_28983,N_29604);
nor UO_3057 (O_3057,N_27203,N_27022);
and UO_3058 (O_3058,N_28028,N_28879);
nor UO_3059 (O_3059,N_28318,N_28820);
and UO_3060 (O_3060,N_29224,N_29800);
nor UO_3061 (O_3061,N_28448,N_29765);
nor UO_3062 (O_3062,N_27852,N_28146);
xnor UO_3063 (O_3063,N_27120,N_29669);
and UO_3064 (O_3064,N_28035,N_29774);
and UO_3065 (O_3065,N_28788,N_29075);
nor UO_3066 (O_3066,N_27024,N_29908);
nor UO_3067 (O_3067,N_28405,N_27564);
or UO_3068 (O_3068,N_29109,N_27531);
or UO_3069 (O_3069,N_29394,N_28816);
or UO_3070 (O_3070,N_28571,N_29655);
xor UO_3071 (O_3071,N_29635,N_29038);
or UO_3072 (O_3072,N_28654,N_28019);
xor UO_3073 (O_3073,N_28068,N_28821);
xor UO_3074 (O_3074,N_28297,N_27438);
nand UO_3075 (O_3075,N_28719,N_27201);
nor UO_3076 (O_3076,N_29170,N_29218);
nand UO_3077 (O_3077,N_27883,N_29212);
nor UO_3078 (O_3078,N_29431,N_29956);
xor UO_3079 (O_3079,N_27049,N_27117);
nand UO_3080 (O_3080,N_29669,N_29016);
xor UO_3081 (O_3081,N_28837,N_28334);
and UO_3082 (O_3082,N_29818,N_27446);
xnor UO_3083 (O_3083,N_29366,N_28972);
or UO_3084 (O_3084,N_29058,N_28398);
nand UO_3085 (O_3085,N_29076,N_29530);
nor UO_3086 (O_3086,N_27102,N_29776);
nand UO_3087 (O_3087,N_29847,N_29592);
and UO_3088 (O_3088,N_27934,N_27341);
nor UO_3089 (O_3089,N_29509,N_27181);
or UO_3090 (O_3090,N_29260,N_29360);
nand UO_3091 (O_3091,N_28379,N_28816);
and UO_3092 (O_3092,N_27036,N_28845);
xor UO_3093 (O_3093,N_28387,N_28377);
or UO_3094 (O_3094,N_28228,N_29410);
or UO_3095 (O_3095,N_29493,N_29481);
or UO_3096 (O_3096,N_29059,N_29722);
nor UO_3097 (O_3097,N_27048,N_28929);
nor UO_3098 (O_3098,N_27580,N_28252);
nand UO_3099 (O_3099,N_27266,N_27403);
or UO_3100 (O_3100,N_29867,N_29010);
and UO_3101 (O_3101,N_29433,N_27882);
nor UO_3102 (O_3102,N_27431,N_28206);
xor UO_3103 (O_3103,N_27953,N_27530);
xor UO_3104 (O_3104,N_29205,N_27044);
nor UO_3105 (O_3105,N_29791,N_28343);
nand UO_3106 (O_3106,N_28728,N_27376);
or UO_3107 (O_3107,N_29070,N_29683);
or UO_3108 (O_3108,N_29889,N_29736);
or UO_3109 (O_3109,N_29496,N_27577);
nand UO_3110 (O_3110,N_28658,N_29915);
and UO_3111 (O_3111,N_27686,N_29510);
or UO_3112 (O_3112,N_27080,N_29437);
xor UO_3113 (O_3113,N_29703,N_29385);
xnor UO_3114 (O_3114,N_28046,N_29913);
or UO_3115 (O_3115,N_27551,N_28890);
or UO_3116 (O_3116,N_27470,N_27040);
nand UO_3117 (O_3117,N_27061,N_29794);
nand UO_3118 (O_3118,N_28495,N_28651);
and UO_3119 (O_3119,N_28137,N_27520);
nand UO_3120 (O_3120,N_29926,N_29230);
or UO_3121 (O_3121,N_28738,N_28501);
nor UO_3122 (O_3122,N_29309,N_27088);
nor UO_3123 (O_3123,N_29700,N_28210);
xor UO_3124 (O_3124,N_28194,N_28481);
or UO_3125 (O_3125,N_27100,N_29035);
xnor UO_3126 (O_3126,N_28820,N_27207);
and UO_3127 (O_3127,N_28902,N_27326);
nand UO_3128 (O_3128,N_29155,N_27151);
or UO_3129 (O_3129,N_27826,N_27994);
nor UO_3130 (O_3130,N_29237,N_29139);
and UO_3131 (O_3131,N_27321,N_28911);
or UO_3132 (O_3132,N_28674,N_28990);
xnor UO_3133 (O_3133,N_27053,N_27755);
xor UO_3134 (O_3134,N_27941,N_28660);
or UO_3135 (O_3135,N_28725,N_28259);
nor UO_3136 (O_3136,N_29958,N_29417);
and UO_3137 (O_3137,N_29510,N_29982);
or UO_3138 (O_3138,N_28055,N_28229);
xnor UO_3139 (O_3139,N_29802,N_28329);
nand UO_3140 (O_3140,N_27181,N_27944);
nand UO_3141 (O_3141,N_28262,N_29154);
xnor UO_3142 (O_3142,N_28920,N_29042);
xor UO_3143 (O_3143,N_27880,N_28575);
and UO_3144 (O_3144,N_29726,N_29028);
nand UO_3145 (O_3145,N_28176,N_27470);
nor UO_3146 (O_3146,N_28598,N_28209);
or UO_3147 (O_3147,N_28532,N_28397);
nand UO_3148 (O_3148,N_28730,N_27007);
and UO_3149 (O_3149,N_27965,N_28935);
or UO_3150 (O_3150,N_28123,N_27988);
or UO_3151 (O_3151,N_28198,N_28283);
and UO_3152 (O_3152,N_27738,N_28084);
or UO_3153 (O_3153,N_29788,N_27490);
nand UO_3154 (O_3154,N_28871,N_27436);
xnor UO_3155 (O_3155,N_28793,N_27880);
xnor UO_3156 (O_3156,N_28712,N_28550);
or UO_3157 (O_3157,N_27415,N_29020);
or UO_3158 (O_3158,N_27315,N_27027);
xnor UO_3159 (O_3159,N_29097,N_27670);
or UO_3160 (O_3160,N_29829,N_28839);
or UO_3161 (O_3161,N_27386,N_28690);
nand UO_3162 (O_3162,N_27170,N_28660);
or UO_3163 (O_3163,N_28071,N_27910);
and UO_3164 (O_3164,N_27142,N_28576);
nor UO_3165 (O_3165,N_29251,N_29752);
and UO_3166 (O_3166,N_29170,N_27383);
xnor UO_3167 (O_3167,N_27940,N_29102);
nor UO_3168 (O_3168,N_27100,N_29939);
or UO_3169 (O_3169,N_27210,N_28069);
nand UO_3170 (O_3170,N_29057,N_28857);
xor UO_3171 (O_3171,N_29524,N_27652);
or UO_3172 (O_3172,N_27878,N_28412);
or UO_3173 (O_3173,N_29638,N_28008);
and UO_3174 (O_3174,N_27643,N_29419);
or UO_3175 (O_3175,N_29640,N_28775);
or UO_3176 (O_3176,N_27189,N_28282);
nand UO_3177 (O_3177,N_27353,N_28799);
xnor UO_3178 (O_3178,N_27605,N_27263);
nor UO_3179 (O_3179,N_29950,N_27063);
or UO_3180 (O_3180,N_27910,N_27064);
xnor UO_3181 (O_3181,N_27023,N_29610);
or UO_3182 (O_3182,N_27114,N_29898);
nand UO_3183 (O_3183,N_29902,N_28385);
or UO_3184 (O_3184,N_27402,N_27200);
and UO_3185 (O_3185,N_27752,N_27371);
nor UO_3186 (O_3186,N_29788,N_28417);
or UO_3187 (O_3187,N_29981,N_27902);
nor UO_3188 (O_3188,N_29244,N_28723);
and UO_3189 (O_3189,N_28217,N_27130);
or UO_3190 (O_3190,N_28205,N_27825);
xor UO_3191 (O_3191,N_28643,N_28186);
and UO_3192 (O_3192,N_28338,N_27658);
xnor UO_3193 (O_3193,N_28031,N_27486);
nand UO_3194 (O_3194,N_29705,N_28013);
or UO_3195 (O_3195,N_29903,N_28721);
nand UO_3196 (O_3196,N_27868,N_27490);
nor UO_3197 (O_3197,N_28324,N_27927);
nand UO_3198 (O_3198,N_29684,N_27546);
and UO_3199 (O_3199,N_29861,N_27466);
xor UO_3200 (O_3200,N_29796,N_28625);
nor UO_3201 (O_3201,N_28388,N_29159);
and UO_3202 (O_3202,N_28419,N_27627);
and UO_3203 (O_3203,N_28986,N_27174);
or UO_3204 (O_3204,N_28938,N_28318);
and UO_3205 (O_3205,N_27665,N_29564);
nor UO_3206 (O_3206,N_29333,N_27849);
nor UO_3207 (O_3207,N_29182,N_29460);
xnor UO_3208 (O_3208,N_28338,N_27715);
or UO_3209 (O_3209,N_29563,N_29650);
nor UO_3210 (O_3210,N_29669,N_28368);
or UO_3211 (O_3211,N_29878,N_27076);
nand UO_3212 (O_3212,N_27783,N_29102);
or UO_3213 (O_3213,N_28097,N_28532);
nand UO_3214 (O_3214,N_27871,N_29256);
nand UO_3215 (O_3215,N_27572,N_29891);
or UO_3216 (O_3216,N_27152,N_28538);
nor UO_3217 (O_3217,N_29700,N_28441);
and UO_3218 (O_3218,N_29702,N_28309);
and UO_3219 (O_3219,N_29838,N_29391);
xnor UO_3220 (O_3220,N_28667,N_29771);
nand UO_3221 (O_3221,N_28915,N_29740);
xor UO_3222 (O_3222,N_27550,N_28347);
or UO_3223 (O_3223,N_27415,N_28693);
and UO_3224 (O_3224,N_28860,N_28040);
and UO_3225 (O_3225,N_28426,N_29874);
nand UO_3226 (O_3226,N_27428,N_29923);
and UO_3227 (O_3227,N_27058,N_28382);
or UO_3228 (O_3228,N_29902,N_28416);
or UO_3229 (O_3229,N_29155,N_29776);
or UO_3230 (O_3230,N_27856,N_28484);
nor UO_3231 (O_3231,N_27385,N_28223);
nor UO_3232 (O_3232,N_29868,N_27785);
and UO_3233 (O_3233,N_29605,N_28497);
xor UO_3234 (O_3234,N_28446,N_28880);
nand UO_3235 (O_3235,N_27452,N_28902);
xor UO_3236 (O_3236,N_27982,N_29521);
and UO_3237 (O_3237,N_29786,N_29277);
or UO_3238 (O_3238,N_29944,N_27774);
and UO_3239 (O_3239,N_28500,N_29260);
nand UO_3240 (O_3240,N_29039,N_29336);
xor UO_3241 (O_3241,N_27513,N_27472);
nor UO_3242 (O_3242,N_29305,N_27689);
or UO_3243 (O_3243,N_28502,N_29086);
nand UO_3244 (O_3244,N_28658,N_27952);
and UO_3245 (O_3245,N_28546,N_28916);
or UO_3246 (O_3246,N_29008,N_28945);
xor UO_3247 (O_3247,N_27554,N_28015);
and UO_3248 (O_3248,N_28000,N_29449);
nand UO_3249 (O_3249,N_27648,N_28269);
nor UO_3250 (O_3250,N_29797,N_27790);
nand UO_3251 (O_3251,N_29685,N_29982);
nand UO_3252 (O_3252,N_27701,N_28421);
or UO_3253 (O_3253,N_29863,N_28286);
and UO_3254 (O_3254,N_29418,N_28502);
and UO_3255 (O_3255,N_27177,N_28935);
and UO_3256 (O_3256,N_27785,N_27499);
nor UO_3257 (O_3257,N_28447,N_27356);
and UO_3258 (O_3258,N_29700,N_29417);
and UO_3259 (O_3259,N_29820,N_29697);
and UO_3260 (O_3260,N_29339,N_28924);
nor UO_3261 (O_3261,N_27557,N_29735);
or UO_3262 (O_3262,N_28463,N_27659);
xor UO_3263 (O_3263,N_29710,N_28245);
nand UO_3264 (O_3264,N_28707,N_29525);
and UO_3265 (O_3265,N_29654,N_28122);
and UO_3266 (O_3266,N_29805,N_29944);
or UO_3267 (O_3267,N_29079,N_28836);
xnor UO_3268 (O_3268,N_27770,N_29507);
nor UO_3269 (O_3269,N_29539,N_27564);
nand UO_3270 (O_3270,N_29750,N_29247);
and UO_3271 (O_3271,N_28777,N_28476);
xor UO_3272 (O_3272,N_28733,N_29236);
and UO_3273 (O_3273,N_28662,N_27645);
nor UO_3274 (O_3274,N_28896,N_29885);
xor UO_3275 (O_3275,N_27326,N_27644);
or UO_3276 (O_3276,N_27816,N_27508);
and UO_3277 (O_3277,N_29169,N_28136);
nor UO_3278 (O_3278,N_29726,N_28801);
nor UO_3279 (O_3279,N_28436,N_28464);
nor UO_3280 (O_3280,N_29568,N_28714);
and UO_3281 (O_3281,N_27221,N_27339);
nor UO_3282 (O_3282,N_27737,N_29418);
or UO_3283 (O_3283,N_28848,N_27907);
nand UO_3284 (O_3284,N_27334,N_28911);
nand UO_3285 (O_3285,N_27756,N_27073);
or UO_3286 (O_3286,N_27918,N_27041);
and UO_3287 (O_3287,N_29836,N_27803);
xnor UO_3288 (O_3288,N_28977,N_28547);
xor UO_3289 (O_3289,N_29506,N_27955);
nand UO_3290 (O_3290,N_27504,N_29032);
and UO_3291 (O_3291,N_27054,N_27639);
xnor UO_3292 (O_3292,N_27973,N_29715);
xnor UO_3293 (O_3293,N_28953,N_27432);
nand UO_3294 (O_3294,N_27796,N_29003);
nand UO_3295 (O_3295,N_27596,N_29206);
xor UO_3296 (O_3296,N_28948,N_28167);
and UO_3297 (O_3297,N_28367,N_28162);
and UO_3298 (O_3298,N_27181,N_28604);
xor UO_3299 (O_3299,N_27737,N_27145);
or UO_3300 (O_3300,N_27717,N_29649);
nor UO_3301 (O_3301,N_27300,N_27446);
xnor UO_3302 (O_3302,N_28830,N_27846);
or UO_3303 (O_3303,N_27228,N_27661);
xnor UO_3304 (O_3304,N_27666,N_28391);
and UO_3305 (O_3305,N_29959,N_28829);
and UO_3306 (O_3306,N_28381,N_27445);
nand UO_3307 (O_3307,N_27557,N_29473);
or UO_3308 (O_3308,N_27572,N_28702);
and UO_3309 (O_3309,N_28558,N_29799);
or UO_3310 (O_3310,N_29275,N_27360);
nand UO_3311 (O_3311,N_29596,N_27638);
and UO_3312 (O_3312,N_27436,N_28389);
and UO_3313 (O_3313,N_29658,N_27565);
nand UO_3314 (O_3314,N_27430,N_27816);
nor UO_3315 (O_3315,N_28412,N_27367);
and UO_3316 (O_3316,N_28960,N_27152);
and UO_3317 (O_3317,N_28736,N_29943);
nand UO_3318 (O_3318,N_28270,N_27549);
xnor UO_3319 (O_3319,N_29117,N_27209);
and UO_3320 (O_3320,N_27240,N_27239);
nand UO_3321 (O_3321,N_27992,N_29534);
nand UO_3322 (O_3322,N_27981,N_28051);
and UO_3323 (O_3323,N_27874,N_27177);
nand UO_3324 (O_3324,N_29538,N_29933);
or UO_3325 (O_3325,N_29301,N_28647);
or UO_3326 (O_3326,N_28368,N_28012);
nand UO_3327 (O_3327,N_28839,N_27920);
nand UO_3328 (O_3328,N_29686,N_28877);
nand UO_3329 (O_3329,N_28814,N_27948);
xor UO_3330 (O_3330,N_27540,N_27717);
nand UO_3331 (O_3331,N_27320,N_28385);
nor UO_3332 (O_3332,N_29338,N_29617);
and UO_3333 (O_3333,N_29248,N_29801);
and UO_3334 (O_3334,N_29396,N_28746);
xnor UO_3335 (O_3335,N_27975,N_27476);
nand UO_3336 (O_3336,N_28741,N_27600);
nor UO_3337 (O_3337,N_28403,N_27883);
and UO_3338 (O_3338,N_28123,N_27278);
or UO_3339 (O_3339,N_29221,N_27808);
nor UO_3340 (O_3340,N_27382,N_28993);
xnor UO_3341 (O_3341,N_29284,N_29604);
nor UO_3342 (O_3342,N_29253,N_29287);
and UO_3343 (O_3343,N_28526,N_28921);
or UO_3344 (O_3344,N_27273,N_29398);
nor UO_3345 (O_3345,N_28257,N_27244);
nand UO_3346 (O_3346,N_27379,N_27846);
nor UO_3347 (O_3347,N_29429,N_29544);
nor UO_3348 (O_3348,N_27916,N_29533);
xnor UO_3349 (O_3349,N_29250,N_29880);
or UO_3350 (O_3350,N_29277,N_29312);
or UO_3351 (O_3351,N_27552,N_27738);
nor UO_3352 (O_3352,N_29354,N_28890);
and UO_3353 (O_3353,N_29999,N_27878);
nor UO_3354 (O_3354,N_27669,N_29985);
and UO_3355 (O_3355,N_28990,N_28691);
xnor UO_3356 (O_3356,N_28533,N_29899);
nor UO_3357 (O_3357,N_27330,N_29732);
or UO_3358 (O_3358,N_27226,N_27521);
nor UO_3359 (O_3359,N_27821,N_28681);
nor UO_3360 (O_3360,N_29966,N_28343);
and UO_3361 (O_3361,N_29645,N_28539);
nor UO_3362 (O_3362,N_27898,N_29916);
nor UO_3363 (O_3363,N_28495,N_27025);
nor UO_3364 (O_3364,N_27753,N_29070);
or UO_3365 (O_3365,N_29067,N_27465);
or UO_3366 (O_3366,N_27635,N_27336);
xor UO_3367 (O_3367,N_28158,N_27360);
or UO_3368 (O_3368,N_29749,N_29886);
nand UO_3369 (O_3369,N_28461,N_28975);
xnor UO_3370 (O_3370,N_27749,N_27461);
and UO_3371 (O_3371,N_27059,N_27786);
nand UO_3372 (O_3372,N_28375,N_27141);
and UO_3373 (O_3373,N_27078,N_29225);
and UO_3374 (O_3374,N_29486,N_28328);
nor UO_3375 (O_3375,N_28959,N_27395);
and UO_3376 (O_3376,N_28832,N_28816);
xor UO_3377 (O_3377,N_29705,N_28331);
nand UO_3378 (O_3378,N_28754,N_27467);
nand UO_3379 (O_3379,N_27395,N_29551);
and UO_3380 (O_3380,N_29419,N_29182);
and UO_3381 (O_3381,N_27083,N_27789);
xor UO_3382 (O_3382,N_29159,N_29687);
or UO_3383 (O_3383,N_28414,N_27083);
or UO_3384 (O_3384,N_28007,N_29491);
xor UO_3385 (O_3385,N_29930,N_28848);
xor UO_3386 (O_3386,N_28438,N_29368);
nand UO_3387 (O_3387,N_27978,N_28875);
or UO_3388 (O_3388,N_27869,N_28215);
xnor UO_3389 (O_3389,N_28775,N_28269);
and UO_3390 (O_3390,N_27741,N_29142);
nand UO_3391 (O_3391,N_27585,N_27375);
nand UO_3392 (O_3392,N_27108,N_27009);
or UO_3393 (O_3393,N_28313,N_28023);
and UO_3394 (O_3394,N_28436,N_28840);
nor UO_3395 (O_3395,N_28479,N_29377);
or UO_3396 (O_3396,N_28349,N_29265);
xnor UO_3397 (O_3397,N_29113,N_28044);
xor UO_3398 (O_3398,N_29489,N_27076);
and UO_3399 (O_3399,N_27255,N_27150);
nor UO_3400 (O_3400,N_29176,N_28522);
xnor UO_3401 (O_3401,N_28955,N_27481);
and UO_3402 (O_3402,N_27316,N_27581);
nand UO_3403 (O_3403,N_27549,N_28042);
nand UO_3404 (O_3404,N_27579,N_27208);
nand UO_3405 (O_3405,N_29520,N_28782);
xnor UO_3406 (O_3406,N_28220,N_27253);
and UO_3407 (O_3407,N_27384,N_29252);
xor UO_3408 (O_3408,N_29683,N_29379);
xor UO_3409 (O_3409,N_29495,N_29223);
and UO_3410 (O_3410,N_29680,N_28914);
and UO_3411 (O_3411,N_28618,N_27335);
and UO_3412 (O_3412,N_29361,N_27994);
nor UO_3413 (O_3413,N_28799,N_27017);
or UO_3414 (O_3414,N_27543,N_28557);
or UO_3415 (O_3415,N_28582,N_29444);
nor UO_3416 (O_3416,N_27546,N_28751);
nand UO_3417 (O_3417,N_29987,N_28363);
nor UO_3418 (O_3418,N_28635,N_27275);
xor UO_3419 (O_3419,N_27489,N_27877);
xnor UO_3420 (O_3420,N_29420,N_28956);
nor UO_3421 (O_3421,N_28811,N_29715);
or UO_3422 (O_3422,N_28738,N_29687);
nand UO_3423 (O_3423,N_29409,N_28816);
or UO_3424 (O_3424,N_29456,N_29174);
nor UO_3425 (O_3425,N_28979,N_29725);
nor UO_3426 (O_3426,N_28925,N_28000);
xor UO_3427 (O_3427,N_29806,N_28471);
nand UO_3428 (O_3428,N_29539,N_28620);
and UO_3429 (O_3429,N_28848,N_28794);
nor UO_3430 (O_3430,N_28694,N_28960);
xor UO_3431 (O_3431,N_28089,N_28886);
nor UO_3432 (O_3432,N_27929,N_27411);
and UO_3433 (O_3433,N_28498,N_29720);
nand UO_3434 (O_3434,N_29458,N_28105);
xor UO_3435 (O_3435,N_27938,N_27490);
nand UO_3436 (O_3436,N_29329,N_29717);
nand UO_3437 (O_3437,N_29986,N_27445);
and UO_3438 (O_3438,N_29188,N_27999);
nand UO_3439 (O_3439,N_29862,N_28186);
or UO_3440 (O_3440,N_27515,N_27228);
or UO_3441 (O_3441,N_29114,N_27483);
nand UO_3442 (O_3442,N_29379,N_27775);
nand UO_3443 (O_3443,N_27511,N_28806);
or UO_3444 (O_3444,N_29300,N_29867);
or UO_3445 (O_3445,N_28645,N_29957);
nor UO_3446 (O_3446,N_27836,N_29530);
nand UO_3447 (O_3447,N_27220,N_28630);
xnor UO_3448 (O_3448,N_28230,N_29663);
or UO_3449 (O_3449,N_28032,N_29622);
and UO_3450 (O_3450,N_27818,N_27883);
xnor UO_3451 (O_3451,N_29089,N_27139);
nor UO_3452 (O_3452,N_29728,N_27333);
xnor UO_3453 (O_3453,N_29860,N_28311);
and UO_3454 (O_3454,N_27666,N_27857);
nand UO_3455 (O_3455,N_27607,N_29549);
nand UO_3456 (O_3456,N_27289,N_28220);
xnor UO_3457 (O_3457,N_27869,N_27324);
and UO_3458 (O_3458,N_29743,N_29639);
nor UO_3459 (O_3459,N_28136,N_27100);
xnor UO_3460 (O_3460,N_27639,N_28018);
xnor UO_3461 (O_3461,N_29248,N_28602);
nor UO_3462 (O_3462,N_27514,N_29136);
xor UO_3463 (O_3463,N_29335,N_28768);
or UO_3464 (O_3464,N_28898,N_29031);
nand UO_3465 (O_3465,N_27420,N_28184);
nand UO_3466 (O_3466,N_29890,N_28590);
nor UO_3467 (O_3467,N_27134,N_27315);
and UO_3468 (O_3468,N_29305,N_27291);
nand UO_3469 (O_3469,N_28051,N_27052);
or UO_3470 (O_3470,N_28498,N_29351);
xor UO_3471 (O_3471,N_29653,N_29717);
nand UO_3472 (O_3472,N_29372,N_27403);
nand UO_3473 (O_3473,N_27544,N_29629);
xnor UO_3474 (O_3474,N_27833,N_27286);
nor UO_3475 (O_3475,N_28545,N_28179);
and UO_3476 (O_3476,N_29014,N_27982);
xnor UO_3477 (O_3477,N_28321,N_28665);
nor UO_3478 (O_3478,N_27410,N_29031);
nor UO_3479 (O_3479,N_29911,N_27930);
nand UO_3480 (O_3480,N_29489,N_27105);
nand UO_3481 (O_3481,N_27936,N_29626);
xor UO_3482 (O_3482,N_28454,N_28529);
nand UO_3483 (O_3483,N_27267,N_27956);
xnor UO_3484 (O_3484,N_29433,N_29486);
or UO_3485 (O_3485,N_29584,N_27972);
nand UO_3486 (O_3486,N_28387,N_29716);
nor UO_3487 (O_3487,N_27522,N_29558);
and UO_3488 (O_3488,N_29769,N_28460);
nand UO_3489 (O_3489,N_29033,N_29863);
or UO_3490 (O_3490,N_27102,N_28037);
xnor UO_3491 (O_3491,N_27043,N_27743);
xor UO_3492 (O_3492,N_27742,N_28618);
xnor UO_3493 (O_3493,N_29730,N_29548);
xnor UO_3494 (O_3494,N_27872,N_29631);
nand UO_3495 (O_3495,N_27628,N_27778);
xor UO_3496 (O_3496,N_27168,N_28101);
nand UO_3497 (O_3497,N_27836,N_27496);
nor UO_3498 (O_3498,N_27946,N_27356);
nor UO_3499 (O_3499,N_27713,N_27932);
endmodule