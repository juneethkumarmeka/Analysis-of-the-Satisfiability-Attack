module basic_1000_10000_1500_4_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_459,In_335);
and U1 (N_1,In_679,In_672);
and U2 (N_2,In_363,In_485);
nand U3 (N_3,In_911,In_396);
or U4 (N_4,In_268,In_352);
nor U5 (N_5,In_512,In_467);
nand U6 (N_6,In_217,In_638);
and U7 (N_7,In_424,In_4);
and U8 (N_8,In_148,In_431);
and U9 (N_9,In_558,In_443);
nand U10 (N_10,In_676,In_616);
xnor U11 (N_11,In_514,In_782);
and U12 (N_12,In_91,In_601);
nor U13 (N_13,In_24,In_765);
and U14 (N_14,In_804,In_16);
and U15 (N_15,In_72,In_416);
nor U16 (N_16,In_341,In_312);
nand U17 (N_17,In_429,In_328);
nor U18 (N_18,In_26,In_550);
nor U19 (N_19,In_496,In_783);
nand U20 (N_20,In_873,In_735);
or U21 (N_21,In_504,In_325);
or U22 (N_22,In_654,In_271);
nor U23 (N_23,In_288,In_45);
and U24 (N_24,In_366,In_880);
nor U25 (N_25,In_207,In_825);
or U26 (N_26,In_808,In_40);
or U27 (N_27,In_499,In_215);
and U28 (N_28,In_297,In_618);
nand U29 (N_29,In_213,In_139);
nor U30 (N_30,In_289,In_517);
and U31 (N_31,In_492,In_607);
nor U32 (N_32,In_145,In_802);
or U33 (N_33,In_827,In_188);
nor U34 (N_34,In_175,In_318);
nand U35 (N_35,In_615,In_342);
nand U36 (N_36,In_187,In_623);
or U37 (N_37,In_681,In_817);
and U38 (N_38,In_264,In_275);
nor U39 (N_39,In_260,In_578);
or U40 (N_40,In_892,In_53);
nor U41 (N_41,In_430,In_47);
and U42 (N_42,In_852,In_540);
nand U43 (N_43,In_794,In_771);
or U44 (N_44,In_59,In_994);
nor U45 (N_45,In_956,In_242);
nor U46 (N_46,In_78,In_869);
xnor U47 (N_47,In_847,In_214);
and U48 (N_48,In_85,In_690);
nor U49 (N_49,In_724,In_929);
or U50 (N_50,In_400,In_32);
and U51 (N_51,In_395,In_426);
or U52 (N_52,In_487,In_980);
nand U53 (N_53,In_351,In_563);
and U54 (N_54,In_893,In_52);
or U55 (N_55,In_889,In_602);
or U56 (N_56,In_954,In_147);
and U57 (N_57,In_585,In_151);
or U58 (N_58,In_593,In_523);
nand U59 (N_59,In_294,In_274);
or U60 (N_60,In_9,In_773);
or U61 (N_61,In_455,In_247);
and U62 (N_62,In_249,In_181);
nor U63 (N_63,In_624,In_451);
nor U64 (N_64,In_453,In_739);
or U65 (N_65,In_678,In_530);
or U66 (N_66,In_870,In_167);
nor U67 (N_67,In_256,In_991);
nor U68 (N_68,In_711,In_903);
nand U69 (N_69,In_749,In_643);
and U70 (N_70,In_904,In_874);
and U71 (N_71,In_486,In_266);
nor U72 (N_72,In_968,In_924);
and U73 (N_73,In_914,In_526);
or U74 (N_74,In_830,In_522);
nor U75 (N_75,In_544,In_600);
nor U76 (N_76,In_969,In_251);
nand U77 (N_77,In_806,In_406);
nor U78 (N_78,In_932,In_941);
and U79 (N_79,In_245,In_770);
and U80 (N_80,In_916,In_134);
or U81 (N_81,In_382,In_344);
and U82 (N_82,In_419,In_810);
or U83 (N_83,In_629,In_358);
nor U84 (N_84,In_218,In_388);
nor U85 (N_85,In_117,In_74);
or U86 (N_86,In_49,In_883);
nand U87 (N_87,In_500,In_938);
or U88 (N_88,In_595,In_273);
nand U89 (N_89,In_712,In_90);
nor U90 (N_90,In_42,In_421);
or U91 (N_91,In_478,In_983);
or U92 (N_92,In_964,In_34);
or U93 (N_93,In_494,In_51);
nor U94 (N_94,In_476,In_906);
nor U95 (N_95,In_977,In_963);
nand U96 (N_96,In_515,In_412);
nor U97 (N_97,In_803,In_714);
and U98 (N_98,In_743,In_591);
and U99 (N_99,In_726,In_594);
or U100 (N_100,In_118,In_308);
and U101 (N_101,In_97,In_706);
and U102 (N_102,In_891,In_882);
or U103 (N_103,In_283,In_390);
nor U104 (N_104,In_915,In_740);
or U105 (N_105,In_166,In_354);
and U106 (N_106,In_686,In_734);
nand U107 (N_107,In_990,In_68);
or U108 (N_108,In_716,In_70);
nor U109 (N_109,In_15,In_502);
or U110 (N_110,In_713,In_458);
and U111 (N_111,In_107,In_89);
and U112 (N_112,In_627,In_570);
nand U113 (N_113,In_310,In_641);
or U114 (N_114,In_322,In_140);
or U115 (N_115,In_848,In_821);
nand U116 (N_116,In_884,In_463);
nand U117 (N_117,In_933,In_332);
and U118 (N_118,In_555,In_119);
and U119 (N_119,In_781,In_282);
nand U120 (N_120,In_754,In_656);
or U121 (N_121,In_392,In_910);
and U122 (N_122,In_890,In_864);
nor U123 (N_123,In_674,In_805);
or U124 (N_124,In_746,In_295);
and U125 (N_125,In_795,In_186);
nor U126 (N_126,In_748,In_133);
nand U127 (N_127,In_509,In_926);
or U128 (N_128,In_222,In_12);
and U129 (N_129,In_225,In_583);
nor U130 (N_130,In_265,In_131);
and U131 (N_131,In_520,In_291);
and U132 (N_132,In_784,In_966);
nor U133 (N_133,In_490,In_603);
or U134 (N_134,In_507,In_420);
nand U135 (N_135,In_612,In_105);
or U136 (N_136,In_423,In_646);
or U137 (N_137,In_73,In_248);
or U138 (N_138,In_564,In_621);
nor U139 (N_139,In_501,In_173);
and U140 (N_140,In_647,In_313);
or U141 (N_141,In_359,In_35);
nand U142 (N_142,In_800,In_587);
or U143 (N_143,In_691,In_315);
or U144 (N_144,In_338,In_785);
nand U145 (N_145,In_87,In_226);
or U146 (N_146,In_239,In_116);
nand U147 (N_147,In_56,In_997);
and U148 (N_148,In_136,In_142);
xor U149 (N_149,In_340,In_123);
and U150 (N_150,In_320,In_143);
and U151 (N_151,In_719,In_745);
nor U152 (N_152,In_409,In_861);
or U153 (N_153,In_162,In_920);
or U154 (N_154,In_436,In_566);
or U155 (N_155,In_872,In_150);
or U156 (N_156,In_54,In_818);
nor U157 (N_157,In_732,In_447);
nand U158 (N_158,In_384,In_285);
and U159 (N_159,In_168,In_981);
nand U160 (N_160,In_721,In_144);
and U161 (N_161,In_940,In_547);
or U162 (N_162,In_820,In_832);
and U163 (N_163,In_546,In_900);
or U164 (N_164,In_841,In_270);
nand U165 (N_165,In_684,In_263);
nor U166 (N_166,In_66,In_157);
nand U167 (N_167,In_855,In_449);
nor U168 (N_168,In_865,In_650);
nand U169 (N_169,In_25,In_863);
xnor U170 (N_170,In_491,In_71);
or U171 (N_171,In_552,In_528);
nor U172 (N_172,In_183,In_577);
or U173 (N_173,In_422,In_524);
or U174 (N_174,In_480,In_859);
nand U175 (N_175,In_586,In_856);
nand U176 (N_176,In_461,In_702);
xor U177 (N_177,In_277,In_200);
or U178 (N_178,In_921,In_508);
nand U179 (N_179,In_115,In_599);
and U180 (N_180,In_441,In_100);
or U181 (N_181,In_323,In_55);
and U182 (N_182,In_975,In_829);
and U183 (N_183,In_521,In_633);
nand U184 (N_184,In_75,In_293);
or U185 (N_185,In_747,In_844);
nand U186 (N_186,In_696,In_448);
nor U187 (N_187,In_238,In_94);
nor U188 (N_188,In_645,In_185);
or U189 (N_189,In_878,In_81);
and U190 (N_190,In_457,In_907);
and U191 (N_191,In_231,In_164);
nand U192 (N_192,In_797,In_815);
and U193 (N_193,In_758,In_337);
and U194 (N_194,In_327,In_667);
nand U195 (N_195,In_464,In_23);
nand U196 (N_196,In_895,In_261);
and U197 (N_197,In_871,In_919);
nand U198 (N_198,In_3,In_573);
nor U199 (N_199,In_571,In_43);
and U200 (N_200,In_896,In_179);
and U201 (N_201,In_39,In_978);
nand U202 (N_202,In_619,In_840);
nand U203 (N_203,In_651,In_755);
or U204 (N_204,In_776,In_553);
nand U205 (N_205,In_965,In_877);
nand U206 (N_206,In_57,In_279);
nand U207 (N_207,In_640,In_398);
nor U208 (N_208,In_854,In_372);
nand U209 (N_209,In_303,In_495);
nand U210 (N_210,In_201,In_163);
nand U211 (N_211,In_210,In_582);
nand U212 (N_212,In_756,In_673);
nor U213 (N_213,In_22,In_302);
or U214 (N_214,In_816,In_554);
or U215 (N_215,In_428,In_703);
nand U216 (N_216,In_17,In_535);
and U217 (N_217,In_2,In_913);
nand U218 (N_218,In_838,In_171);
nand U219 (N_219,In_999,In_113);
and U220 (N_220,In_622,In_246);
xor U221 (N_221,In_664,In_159);
nand U222 (N_222,In_741,In_330);
nor U223 (N_223,In_208,In_88);
and U224 (N_224,In_809,In_733);
nor U225 (N_225,In_833,In_127);
nor U226 (N_226,In_10,In_280);
or U227 (N_227,In_109,In_284);
nor U228 (N_228,In_787,In_18);
and U229 (N_229,In_93,In_620);
nor U230 (N_230,In_205,In_172);
or U231 (N_231,In_232,In_321);
or U232 (N_232,In_826,In_763);
nand U233 (N_233,In_596,In_61);
nor U234 (N_234,In_391,In_767);
and U235 (N_235,In_567,In_760);
or U236 (N_236,In_738,In_19);
nand U237 (N_237,In_154,In_692);
nor U238 (N_238,In_375,In_106);
nor U239 (N_239,In_757,In_551);
nand U240 (N_240,In_37,In_402);
nand U241 (N_241,In_697,In_584);
nor U242 (N_242,In_69,In_837);
and U243 (N_243,In_206,In_862);
nand U244 (N_244,In_780,In_202);
or U245 (N_245,In_959,In_834);
or U246 (N_246,In_170,In_102);
or U247 (N_247,In_184,In_717);
nand U248 (N_248,In_949,In_510);
xor U249 (N_249,In_474,In_65);
nand U250 (N_250,In_927,In_946);
and U251 (N_251,In_197,In_744);
nand U252 (N_252,In_945,In_132);
nand U253 (N_253,In_807,In_793);
and U254 (N_254,In_588,In_452);
and U255 (N_255,In_683,In_385);
nor U256 (N_256,In_709,In_377);
nor U257 (N_257,In_287,In_434);
nor U258 (N_258,In_425,In_44);
nor U259 (N_259,In_575,In_176);
nor U260 (N_260,In_326,In_298);
or U261 (N_261,In_814,In_153);
or U262 (N_262,In_637,In_533);
and U263 (N_263,In_936,In_92);
or U264 (N_264,In_427,In_648);
nand U265 (N_265,In_20,In_41);
nand U266 (N_266,In_403,In_408);
nor U267 (N_267,In_345,In_418);
and U268 (N_268,In_775,In_152);
and U269 (N_269,In_894,In_982);
and U270 (N_270,In_935,In_475);
nand U271 (N_271,In_715,In_301);
nand U272 (N_272,In_300,In_7);
or U273 (N_273,In_989,In_652);
nand U274 (N_274,In_851,In_155);
nor U275 (N_275,In_364,In_636);
or U276 (N_276,In_897,In_948);
nand U277 (N_277,In_227,In_158);
nand U278 (N_278,In_952,In_866);
and U279 (N_279,In_468,In_708);
nand U280 (N_280,In_343,In_482);
nor U281 (N_281,In_369,In_876);
nand U282 (N_282,In_146,In_8);
nor U283 (N_283,In_761,In_126);
nand U284 (N_284,In_376,In_137);
or U285 (N_285,In_190,In_138);
xor U286 (N_286,In_525,In_367);
xnor U287 (N_287,In_174,In_296);
nor U288 (N_288,In_737,In_565);
and U289 (N_289,In_233,In_576);
nor U290 (N_290,In_460,In_542);
or U291 (N_291,In_886,In_62);
or U292 (N_292,In_680,In_110);
nor U293 (N_293,In_6,In_488);
nor U294 (N_294,In_483,In_701);
nor U295 (N_295,In_29,In_687);
nor U296 (N_296,In_108,In_842);
or U297 (N_297,In_779,In_259);
nand U298 (N_298,In_671,In_608);
nand U299 (N_299,In_631,In_710);
nand U300 (N_300,In_628,In_898);
nor U301 (N_301,In_511,In_357);
nor U302 (N_302,In_822,In_254);
nor U303 (N_303,In_722,In_845);
and U304 (N_304,In_662,In_456);
nor U305 (N_305,In_698,In_195);
and U306 (N_306,In_923,In_286);
nor U307 (N_307,In_630,In_433);
xor U308 (N_308,In_356,In_617);
nor U309 (N_309,In_128,In_812);
nor U310 (N_310,In_489,In_48);
or U311 (N_311,In_262,In_389);
or U312 (N_312,In_568,In_958);
and U313 (N_313,In_473,In_828);
nand U314 (N_314,In_967,In_331);
nor U315 (N_315,In_665,In_543);
nand U316 (N_316,In_953,In_875);
nor U317 (N_317,In_435,In_518);
or U318 (N_318,In_442,In_413);
nor U319 (N_319,In_731,In_979);
nor U320 (N_320,In_574,In_944);
nand U321 (N_321,In_347,In_998);
and U322 (N_322,In_901,In_751);
nand U323 (N_323,In_789,In_36);
nor U324 (N_324,In_657,In_130);
or U325 (N_325,In_272,In_58);
or U326 (N_326,In_417,In_292);
or U327 (N_327,In_446,In_120);
nand U328 (N_328,In_885,In_212);
or U329 (N_329,In_5,In_768);
nor U330 (N_330,In_194,In_639);
xnor U331 (N_331,In_850,In_21);
or U332 (N_332,In_970,In_267);
nand U333 (N_333,In_677,In_378);
or U334 (N_334,In_700,In_67);
nor U335 (N_335,In_196,In_439);
nand U336 (N_336,In_614,In_723);
nor U337 (N_337,In_498,In_182);
and U338 (N_338,In_947,In_819);
nor U339 (N_339,In_393,In_655);
and U340 (N_340,In_305,In_529);
nand U341 (N_341,In_532,In_560);
and U342 (N_342,In_549,In_561);
nor U343 (N_343,In_705,In_193);
or U344 (N_344,In_221,In_943);
and U345 (N_345,In_813,In_937);
or U346 (N_346,In_778,In_960);
and U347 (N_347,In_250,In_198);
nor U348 (N_348,In_505,In_831);
or U349 (N_349,In_635,In_604);
nor U350 (N_350,In_481,In_169);
nand U351 (N_351,In_365,In_83);
nand U352 (N_352,In_304,In_613);
and U353 (N_353,In_27,In_465);
nand U354 (N_354,In_811,In_592);
nand U355 (N_355,In_971,In_466);
and U356 (N_356,In_996,In_14);
nand U357 (N_357,In_278,In_368);
and U358 (N_358,In_902,In_580);
nand U359 (N_359,In_868,In_661);
or U360 (N_360,In_96,In_370);
and U361 (N_361,In_995,In_727);
and U362 (N_362,In_432,In_668);
nor U363 (N_363,In_203,In_404);
nand U364 (N_364,In_234,In_497);
or U365 (N_365,In_644,In_33);
nand U366 (N_366,In_13,In_986);
or U367 (N_367,In_685,In_209);
and U368 (N_368,In_707,In_559);
nand U369 (N_369,In_383,In_135);
nor U370 (N_370,In_742,In_762);
nand U371 (N_371,In_887,In_791);
nor U372 (N_372,In_753,In_230);
nor U373 (N_373,In_216,In_394);
and U374 (N_374,In_371,In_792);
nand U375 (N_375,In_976,In_414);
and U376 (N_376,In_632,In_76);
and U377 (N_377,In_539,In_860);
nor U378 (N_378,In_857,In_317);
or U379 (N_379,In_228,In_984);
or U380 (N_380,In_440,In_670);
nand U381 (N_381,In_224,In_899);
nand U382 (N_382,In_111,In_255);
or U383 (N_383,In_688,In_649);
and U384 (N_384,In_407,In_663);
or U385 (N_385,In_114,In_161);
nor U386 (N_386,In_450,In_538);
nand U387 (N_387,In_788,In_579);
and U388 (N_388,In_454,In_477);
and U389 (N_389,In_545,In_240);
and U390 (N_390,In_125,In_930);
nand U391 (N_391,In_379,In_634);
or U392 (N_392,In_470,In_177);
nand U393 (N_393,In_374,In_84);
nor U394 (N_394,In_839,In_858);
and U395 (N_395,In_824,In_349);
nor U396 (N_396,In_104,In_598);
nand U397 (N_397,In_165,In_973);
nand U398 (N_398,In_659,In_581);
nand U399 (N_399,In_63,In_316);
or U400 (N_400,In_401,In_471);
or U401 (N_401,In_361,In_957);
nor U402 (N_402,In_269,In_950);
nand U403 (N_403,In_189,In_399);
nor U404 (N_404,In_493,In_752);
and U405 (N_405,In_124,In_642);
xor U406 (N_406,In_972,In_122);
and U407 (N_407,In_556,In_355);
nand U408 (N_408,In_503,In_849);
nand U409 (N_409,In_694,In_241);
and U410 (N_410,In_82,In_766);
or U411 (N_411,In_38,In_922);
nand U412 (N_412,In_334,In_772);
nand U413 (N_413,In_333,In_1);
nor U414 (N_414,In_103,In_191);
nand U415 (N_415,In_360,In_728);
and U416 (N_416,In_993,In_536);
or U417 (N_417,In_843,In_777);
and U418 (N_418,In_362,In_86);
nor U419 (N_419,In_597,In_386);
and U420 (N_420,In_699,In_479);
nand U421 (N_421,In_309,In_31);
nand U422 (N_422,In_888,In_625);
and U423 (N_423,In_387,In_77);
and U424 (N_424,In_314,In_934);
or U425 (N_425,In_557,In_660);
nand U426 (N_426,In_590,In_750);
or U427 (N_427,In_626,In_484);
nor U428 (N_428,In_918,In_50);
and U429 (N_429,In_799,In_879);
and U430 (N_430,In_257,In_955);
and U431 (N_431,In_204,In_373);
or U432 (N_432,In_237,In_675);
nor U433 (N_433,In_846,In_101);
and U434 (N_434,In_112,In_801);
or U435 (N_435,In_192,In_736);
nand U436 (N_436,In_867,In_606);
nor U437 (N_437,In_836,In_444);
nand U438 (N_438,In_987,In_415);
and U439 (N_439,In_541,In_764);
nand U440 (N_440,In_324,In_730);
nor U441 (N_441,In_462,In_689);
nand U442 (N_442,In_786,In_759);
and U443 (N_443,In_244,In_258);
nor U444 (N_444,In_669,In_307);
nor U445 (N_445,In_531,In_410);
nand U446 (N_446,In_411,In_199);
nand U447 (N_447,In_306,In_506);
nand U448 (N_448,In_79,In_942);
xor U449 (N_449,In_569,In_925);
nor U450 (N_450,In_99,In_516);
nand U451 (N_451,In_774,In_796);
nor U452 (N_452,In_985,In_380);
nor U453 (N_453,In_64,In_835);
nor U454 (N_454,In_605,In_243);
nor U455 (N_455,In_534,In_60);
nor U456 (N_456,In_438,In_95);
nand U457 (N_457,In_823,In_729);
nor U458 (N_458,In_704,In_769);
nand U459 (N_459,In_682,In_961);
or U460 (N_460,In_229,In_472);
or U461 (N_461,In_235,In_917);
nor U462 (N_462,In_611,In_988);
or U463 (N_463,In_653,In_311);
and U464 (N_464,In_223,In_572);
nor U465 (N_465,In_381,In_339);
nand U466 (N_466,In_329,In_974);
and U467 (N_467,In_513,In_527);
nand U468 (N_468,In_253,In_905);
nor U469 (N_469,In_912,In_28);
nand U470 (N_470,In_609,In_445);
or U471 (N_471,In_951,In_336);
nor U472 (N_472,In_178,In_211);
or U473 (N_473,In_469,In_160);
nor U474 (N_474,In_276,In_437);
nor U475 (N_475,In_350,In_353);
nor U476 (N_476,In_589,In_962);
or U477 (N_477,In_180,In_939);
and U478 (N_478,In_798,In_562);
and U479 (N_479,In_346,In_98);
nor U480 (N_480,In_281,In_519);
and U481 (N_481,In_909,In_853);
and U482 (N_482,In_928,In_658);
and U483 (N_483,In_397,In_129);
nor U484 (N_484,In_908,In_537);
and U485 (N_485,In_80,In_121);
nand U486 (N_486,In_405,In_881);
or U487 (N_487,In_992,In_149);
nor U488 (N_488,In_666,In_790);
and U489 (N_489,In_30,In_610);
and U490 (N_490,In_0,In_720);
nand U491 (N_491,In_319,In_718);
and U492 (N_492,In_46,In_219);
nand U493 (N_493,In_220,In_299);
nor U494 (N_494,In_290,In_11);
and U495 (N_495,In_156,In_548);
nand U496 (N_496,In_725,In_931);
nand U497 (N_497,In_348,In_693);
nand U498 (N_498,In_236,In_141);
nor U499 (N_499,In_252,In_695);
nand U500 (N_500,In_920,In_846);
nor U501 (N_501,In_545,In_104);
and U502 (N_502,In_819,In_148);
or U503 (N_503,In_201,In_225);
and U504 (N_504,In_124,In_448);
nor U505 (N_505,In_116,In_77);
or U506 (N_506,In_250,In_774);
and U507 (N_507,In_892,In_31);
nor U508 (N_508,In_404,In_741);
or U509 (N_509,In_392,In_675);
nand U510 (N_510,In_347,In_864);
nand U511 (N_511,In_160,In_848);
or U512 (N_512,In_437,In_412);
nor U513 (N_513,In_760,In_814);
nor U514 (N_514,In_186,In_698);
and U515 (N_515,In_164,In_265);
nor U516 (N_516,In_967,In_175);
and U517 (N_517,In_463,In_698);
or U518 (N_518,In_925,In_568);
nand U519 (N_519,In_784,In_741);
nand U520 (N_520,In_332,In_708);
nor U521 (N_521,In_122,In_505);
nor U522 (N_522,In_105,In_923);
and U523 (N_523,In_860,In_123);
and U524 (N_524,In_770,In_410);
and U525 (N_525,In_792,In_269);
nand U526 (N_526,In_435,In_434);
nand U527 (N_527,In_333,In_505);
nand U528 (N_528,In_224,In_340);
and U529 (N_529,In_517,In_410);
or U530 (N_530,In_784,In_186);
nand U531 (N_531,In_455,In_454);
nand U532 (N_532,In_947,In_13);
or U533 (N_533,In_334,In_712);
nor U534 (N_534,In_630,In_406);
and U535 (N_535,In_476,In_992);
or U536 (N_536,In_548,In_450);
or U537 (N_537,In_954,In_742);
nand U538 (N_538,In_964,In_733);
and U539 (N_539,In_306,In_806);
nand U540 (N_540,In_444,In_446);
xor U541 (N_541,In_945,In_668);
nor U542 (N_542,In_34,In_234);
and U543 (N_543,In_948,In_693);
and U544 (N_544,In_815,In_326);
nor U545 (N_545,In_213,In_532);
nor U546 (N_546,In_229,In_660);
nand U547 (N_547,In_550,In_887);
and U548 (N_548,In_285,In_725);
and U549 (N_549,In_841,In_949);
nor U550 (N_550,In_176,In_810);
nor U551 (N_551,In_668,In_647);
or U552 (N_552,In_639,In_609);
and U553 (N_553,In_737,In_768);
and U554 (N_554,In_180,In_831);
and U555 (N_555,In_936,In_968);
nand U556 (N_556,In_477,In_433);
or U557 (N_557,In_105,In_508);
or U558 (N_558,In_780,In_689);
and U559 (N_559,In_320,In_120);
nor U560 (N_560,In_569,In_736);
and U561 (N_561,In_531,In_817);
nand U562 (N_562,In_652,In_405);
nor U563 (N_563,In_154,In_690);
nand U564 (N_564,In_792,In_793);
nand U565 (N_565,In_560,In_745);
or U566 (N_566,In_917,In_225);
nand U567 (N_567,In_497,In_276);
and U568 (N_568,In_949,In_720);
or U569 (N_569,In_704,In_460);
nand U570 (N_570,In_403,In_255);
nor U571 (N_571,In_972,In_786);
nor U572 (N_572,In_523,In_123);
or U573 (N_573,In_960,In_296);
nand U574 (N_574,In_901,In_246);
nor U575 (N_575,In_929,In_975);
nor U576 (N_576,In_847,In_562);
or U577 (N_577,In_104,In_103);
nor U578 (N_578,In_118,In_556);
nand U579 (N_579,In_769,In_496);
and U580 (N_580,In_881,In_462);
nand U581 (N_581,In_72,In_767);
or U582 (N_582,In_613,In_95);
nor U583 (N_583,In_383,In_155);
and U584 (N_584,In_76,In_2);
nand U585 (N_585,In_383,In_248);
or U586 (N_586,In_485,In_3);
nor U587 (N_587,In_466,In_148);
nor U588 (N_588,In_603,In_609);
and U589 (N_589,In_906,In_529);
nand U590 (N_590,In_356,In_241);
nand U591 (N_591,In_415,In_12);
and U592 (N_592,In_918,In_825);
nand U593 (N_593,In_483,In_462);
nand U594 (N_594,In_65,In_259);
nand U595 (N_595,In_954,In_758);
nand U596 (N_596,In_875,In_654);
nor U597 (N_597,In_196,In_892);
nand U598 (N_598,In_697,In_52);
nand U599 (N_599,In_876,In_167);
nand U600 (N_600,In_115,In_506);
and U601 (N_601,In_603,In_924);
nor U602 (N_602,In_857,In_448);
nor U603 (N_603,In_605,In_606);
nor U604 (N_604,In_681,In_474);
nand U605 (N_605,In_531,In_376);
nand U606 (N_606,In_179,In_717);
and U607 (N_607,In_691,In_128);
or U608 (N_608,In_451,In_937);
or U609 (N_609,In_784,In_526);
or U610 (N_610,In_694,In_449);
and U611 (N_611,In_376,In_725);
and U612 (N_612,In_451,In_809);
nand U613 (N_613,In_683,In_576);
xor U614 (N_614,In_156,In_728);
or U615 (N_615,In_376,In_803);
or U616 (N_616,In_942,In_482);
or U617 (N_617,In_220,In_733);
and U618 (N_618,In_284,In_747);
nor U619 (N_619,In_1,In_590);
or U620 (N_620,In_606,In_553);
and U621 (N_621,In_244,In_633);
nor U622 (N_622,In_623,In_961);
or U623 (N_623,In_225,In_36);
nor U624 (N_624,In_612,In_688);
nand U625 (N_625,In_274,In_735);
nor U626 (N_626,In_264,In_844);
and U627 (N_627,In_115,In_749);
nand U628 (N_628,In_691,In_155);
and U629 (N_629,In_457,In_394);
or U630 (N_630,In_874,In_415);
nand U631 (N_631,In_828,In_617);
nand U632 (N_632,In_573,In_703);
nor U633 (N_633,In_787,In_488);
and U634 (N_634,In_625,In_744);
or U635 (N_635,In_278,In_733);
or U636 (N_636,In_25,In_240);
or U637 (N_637,In_450,In_998);
and U638 (N_638,In_636,In_357);
and U639 (N_639,In_104,In_276);
nand U640 (N_640,In_709,In_823);
and U641 (N_641,In_966,In_947);
and U642 (N_642,In_721,In_907);
and U643 (N_643,In_74,In_875);
nor U644 (N_644,In_632,In_558);
nand U645 (N_645,In_765,In_145);
or U646 (N_646,In_684,In_544);
nor U647 (N_647,In_509,In_979);
nand U648 (N_648,In_205,In_692);
nand U649 (N_649,In_786,In_710);
or U650 (N_650,In_686,In_366);
nand U651 (N_651,In_972,In_230);
nand U652 (N_652,In_526,In_637);
or U653 (N_653,In_873,In_792);
nor U654 (N_654,In_16,In_846);
nor U655 (N_655,In_127,In_810);
nor U656 (N_656,In_252,In_785);
or U657 (N_657,In_158,In_74);
or U658 (N_658,In_524,In_526);
nor U659 (N_659,In_126,In_826);
and U660 (N_660,In_705,In_162);
nand U661 (N_661,In_312,In_107);
or U662 (N_662,In_664,In_74);
nor U663 (N_663,In_277,In_398);
and U664 (N_664,In_394,In_849);
nand U665 (N_665,In_515,In_908);
and U666 (N_666,In_965,In_67);
or U667 (N_667,In_580,In_76);
and U668 (N_668,In_952,In_313);
nor U669 (N_669,In_840,In_469);
nor U670 (N_670,In_217,In_278);
and U671 (N_671,In_647,In_987);
nand U672 (N_672,In_244,In_323);
nor U673 (N_673,In_730,In_467);
nand U674 (N_674,In_153,In_815);
or U675 (N_675,In_518,In_353);
and U676 (N_676,In_876,In_23);
nand U677 (N_677,In_15,In_392);
or U678 (N_678,In_742,In_138);
or U679 (N_679,In_690,In_974);
nand U680 (N_680,In_118,In_982);
nand U681 (N_681,In_407,In_299);
and U682 (N_682,In_182,In_806);
nor U683 (N_683,In_734,In_963);
nand U684 (N_684,In_987,In_961);
nand U685 (N_685,In_695,In_145);
or U686 (N_686,In_417,In_287);
or U687 (N_687,In_677,In_644);
or U688 (N_688,In_786,In_756);
or U689 (N_689,In_974,In_646);
or U690 (N_690,In_784,In_375);
nand U691 (N_691,In_580,In_334);
or U692 (N_692,In_907,In_197);
nand U693 (N_693,In_950,In_84);
and U694 (N_694,In_42,In_319);
nand U695 (N_695,In_288,In_504);
and U696 (N_696,In_533,In_127);
nor U697 (N_697,In_933,In_327);
xnor U698 (N_698,In_198,In_324);
or U699 (N_699,In_543,In_998);
nor U700 (N_700,In_96,In_351);
nand U701 (N_701,In_479,In_774);
or U702 (N_702,In_917,In_269);
or U703 (N_703,In_321,In_439);
and U704 (N_704,In_724,In_210);
and U705 (N_705,In_500,In_412);
and U706 (N_706,In_481,In_142);
or U707 (N_707,In_474,In_33);
or U708 (N_708,In_326,In_205);
and U709 (N_709,In_807,In_298);
nand U710 (N_710,In_944,In_475);
and U711 (N_711,In_277,In_302);
nor U712 (N_712,In_470,In_678);
nor U713 (N_713,In_539,In_567);
nor U714 (N_714,In_804,In_198);
or U715 (N_715,In_180,In_150);
or U716 (N_716,In_46,In_347);
nand U717 (N_717,In_85,In_740);
nor U718 (N_718,In_104,In_959);
nor U719 (N_719,In_901,In_980);
nand U720 (N_720,In_227,In_697);
or U721 (N_721,In_733,In_616);
or U722 (N_722,In_934,In_461);
or U723 (N_723,In_292,In_720);
nand U724 (N_724,In_177,In_856);
or U725 (N_725,In_30,In_387);
nor U726 (N_726,In_3,In_320);
nand U727 (N_727,In_631,In_913);
nand U728 (N_728,In_338,In_824);
nand U729 (N_729,In_341,In_644);
nand U730 (N_730,In_76,In_889);
nand U731 (N_731,In_337,In_966);
or U732 (N_732,In_939,In_369);
nand U733 (N_733,In_549,In_250);
nor U734 (N_734,In_665,In_57);
or U735 (N_735,In_170,In_147);
and U736 (N_736,In_32,In_536);
or U737 (N_737,In_870,In_270);
nor U738 (N_738,In_812,In_107);
nor U739 (N_739,In_166,In_30);
or U740 (N_740,In_452,In_764);
nor U741 (N_741,In_643,In_67);
nor U742 (N_742,In_181,In_957);
and U743 (N_743,In_878,In_50);
or U744 (N_744,In_446,In_418);
and U745 (N_745,In_317,In_732);
nor U746 (N_746,In_341,In_499);
and U747 (N_747,In_517,In_185);
and U748 (N_748,In_54,In_950);
and U749 (N_749,In_639,In_698);
nor U750 (N_750,In_511,In_243);
or U751 (N_751,In_829,In_596);
xnor U752 (N_752,In_926,In_672);
nor U753 (N_753,In_635,In_96);
and U754 (N_754,In_966,In_748);
nand U755 (N_755,In_202,In_207);
and U756 (N_756,In_932,In_960);
nor U757 (N_757,In_801,In_959);
and U758 (N_758,In_940,In_611);
and U759 (N_759,In_317,In_125);
and U760 (N_760,In_529,In_767);
and U761 (N_761,In_750,In_959);
nand U762 (N_762,In_134,In_460);
and U763 (N_763,In_521,In_695);
or U764 (N_764,In_980,In_597);
and U765 (N_765,In_145,In_334);
nand U766 (N_766,In_575,In_940);
or U767 (N_767,In_786,In_240);
nand U768 (N_768,In_187,In_470);
nor U769 (N_769,In_457,In_742);
nor U770 (N_770,In_741,In_100);
nor U771 (N_771,In_458,In_120);
nand U772 (N_772,In_318,In_653);
nand U773 (N_773,In_759,In_3);
or U774 (N_774,In_580,In_716);
xnor U775 (N_775,In_633,In_775);
nor U776 (N_776,In_144,In_72);
nand U777 (N_777,In_268,In_302);
and U778 (N_778,In_397,In_679);
and U779 (N_779,In_368,In_228);
or U780 (N_780,In_657,In_569);
nand U781 (N_781,In_881,In_243);
or U782 (N_782,In_607,In_68);
or U783 (N_783,In_276,In_81);
nor U784 (N_784,In_757,In_583);
nor U785 (N_785,In_928,In_102);
nor U786 (N_786,In_55,In_928);
and U787 (N_787,In_350,In_697);
nand U788 (N_788,In_90,In_704);
nand U789 (N_789,In_133,In_462);
nor U790 (N_790,In_55,In_427);
and U791 (N_791,In_63,In_383);
nand U792 (N_792,In_460,In_961);
nand U793 (N_793,In_770,In_734);
nand U794 (N_794,In_825,In_640);
and U795 (N_795,In_760,In_29);
nor U796 (N_796,In_344,In_99);
nand U797 (N_797,In_20,In_949);
nand U798 (N_798,In_977,In_486);
nor U799 (N_799,In_221,In_511);
nand U800 (N_800,In_497,In_208);
nor U801 (N_801,In_745,In_339);
or U802 (N_802,In_20,In_707);
or U803 (N_803,In_318,In_515);
nand U804 (N_804,In_432,In_967);
nor U805 (N_805,In_593,In_562);
nor U806 (N_806,In_34,In_522);
nor U807 (N_807,In_867,In_499);
nand U808 (N_808,In_546,In_176);
nor U809 (N_809,In_304,In_416);
xnor U810 (N_810,In_29,In_987);
or U811 (N_811,In_592,In_438);
nand U812 (N_812,In_77,In_231);
nand U813 (N_813,In_973,In_661);
and U814 (N_814,In_661,In_313);
nor U815 (N_815,In_76,In_652);
and U816 (N_816,In_207,In_476);
or U817 (N_817,In_194,In_51);
nand U818 (N_818,In_765,In_793);
nand U819 (N_819,In_515,In_444);
nand U820 (N_820,In_442,In_597);
or U821 (N_821,In_920,In_315);
nor U822 (N_822,In_71,In_418);
nor U823 (N_823,In_794,In_486);
nor U824 (N_824,In_25,In_590);
nor U825 (N_825,In_970,In_398);
and U826 (N_826,In_647,In_679);
or U827 (N_827,In_697,In_450);
and U828 (N_828,In_11,In_939);
and U829 (N_829,In_771,In_256);
and U830 (N_830,In_219,In_603);
nand U831 (N_831,In_41,In_669);
and U832 (N_832,In_261,In_583);
or U833 (N_833,In_603,In_482);
and U834 (N_834,In_916,In_959);
and U835 (N_835,In_140,In_836);
or U836 (N_836,In_628,In_244);
nor U837 (N_837,In_46,In_925);
nand U838 (N_838,In_250,In_146);
or U839 (N_839,In_801,In_396);
and U840 (N_840,In_626,In_140);
or U841 (N_841,In_212,In_404);
nand U842 (N_842,In_532,In_896);
or U843 (N_843,In_420,In_707);
nand U844 (N_844,In_894,In_207);
nor U845 (N_845,In_940,In_410);
nand U846 (N_846,In_844,In_700);
or U847 (N_847,In_457,In_856);
nand U848 (N_848,In_934,In_408);
and U849 (N_849,In_229,In_133);
nor U850 (N_850,In_512,In_360);
nor U851 (N_851,In_745,In_269);
nand U852 (N_852,In_10,In_734);
nor U853 (N_853,In_139,In_808);
and U854 (N_854,In_318,In_726);
nand U855 (N_855,In_406,In_67);
and U856 (N_856,In_594,In_450);
nor U857 (N_857,In_697,In_687);
or U858 (N_858,In_687,In_1);
or U859 (N_859,In_921,In_745);
nor U860 (N_860,In_768,In_925);
nor U861 (N_861,In_957,In_286);
or U862 (N_862,In_762,In_465);
and U863 (N_863,In_684,In_555);
nand U864 (N_864,In_331,In_214);
nand U865 (N_865,In_655,In_183);
nor U866 (N_866,In_132,In_28);
nor U867 (N_867,In_352,In_609);
nor U868 (N_868,In_889,In_766);
or U869 (N_869,In_675,In_86);
nor U870 (N_870,In_555,In_553);
or U871 (N_871,In_553,In_542);
or U872 (N_872,In_649,In_966);
or U873 (N_873,In_162,In_166);
nor U874 (N_874,In_751,In_808);
or U875 (N_875,In_45,In_328);
nor U876 (N_876,In_558,In_299);
or U877 (N_877,In_726,In_326);
nor U878 (N_878,In_486,In_685);
nor U879 (N_879,In_752,In_746);
and U880 (N_880,In_208,In_253);
nand U881 (N_881,In_608,In_220);
or U882 (N_882,In_470,In_860);
and U883 (N_883,In_117,In_506);
or U884 (N_884,In_409,In_404);
and U885 (N_885,In_937,In_67);
nand U886 (N_886,In_2,In_327);
and U887 (N_887,In_769,In_691);
or U888 (N_888,In_246,In_956);
or U889 (N_889,In_493,In_98);
nand U890 (N_890,In_780,In_445);
and U891 (N_891,In_596,In_437);
and U892 (N_892,In_722,In_637);
or U893 (N_893,In_484,In_859);
and U894 (N_894,In_865,In_281);
or U895 (N_895,In_918,In_669);
and U896 (N_896,In_836,In_70);
nor U897 (N_897,In_9,In_806);
or U898 (N_898,In_930,In_203);
nand U899 (N_899,In_703,In_974);
nor U900 (N_900,In_438,In_679);
or U901 (N_901,In_576,In_702);
nor U902 (N_902,In_450,In_943);
nand U903 (N_903,In_865,In_419);
or U904 (N_904,In_836,In_600);
or U905 (N_905,In_986,In_381);
nor U906 (N_906,In_131,In_293);
nor U907 (N_907,In_843,In_640);
xnor U908 (N_908,In_890,In_199);
or U909 (N_909,In_819,In_894);
or U910 (N_910,In_857,In_404);
nor U911 (N_911,In_308,In_825);
nor U912 (N_912,In_216,In_371);
nor U913 (N_913,In_888,In_624);
or U914 (N_914,In_735,In_846);
or U915 (N_915,In_574,In_805);
nor U916 (N_916,In_234,In_232);
nand U917 (N_917,In_581,In_548);
or U918 (N_918,In_759,In_866);
nor U919 (N_919,In_231,In_984);
and U920 (N_920,In_349,In_379);
and U921 (N_921,In_169,In_279);
and U922 (N_922,In_902,In_340);
nand U923 (N_923,In_626,In_955);
or U924 (N_924,In_944,In_568);
nand U925 (N_925,In_531,In_503);
and U926 (N_926,In_831,In_651);
and U927 (N_927,In_310,In_376);
and U928 (N_928,In_859,In_781);
or U929 (N_929,In_288,In_170);
and U930 (N_930,In_487,In_114);
nor U931 (N_931,In_834,In_753);
and U932 (N_932,In_853,In_75);
nor U933 (N_933,In_311,In_919);
or U934 (N_934,In_725,In_945);
and U935 (N_935,In_511,In_320);
nor U936 (N_936,In_818,In_395);
nand U937 (N_937,In_299,In_369);
nor U938 (N_938,In_322,In_143);
or U939 (N_939,In_401,In_604);
nand U940 (N_940,In_364,In_965);
or U941 (N_941,In_940,In_963);
nor U942 (N_942,In_297,In_72);
nor U943 (N_943,In_799,In_184);
nand U944 (N_944,In_506,In_266);
nand U945 (N_945,In_311,In_625);
nand U946 (N_946,In_755,In_107);
nand U947 (N_947,In_258,In_246);
nor U948 (N_948,In_868,In_21);
nor U949 (N_949,In_804,In_458);
xnor U950 (N_950,In_142,In_832);
nor U951 (N_951,In_396,In_336);
and U952 (N_952,In_654,In_530);
or U953 (N_953,In_393,In_222);
nand U954 (N_954,In_641,In_837);
nor U955 (N_955,In_334,In_98);
or U956 (N_956,In_306,In_941);
nand U957 (N_957,In_653,In_119);
nand U958 (N_958,In_313,In_457);
nand U959 (N_959,In_531,In_801);
and U960 (N_960,In_699,In_539);
and U961 (N_961,In_489,In_768);
and U962 (N_962,In_956,In_4);
nor U963 (N_963,In_781,In_574);
nor U964 (N_964,In_254,In_652);
nand U965 (N_965,In_117,In_865);
or U966 (N_966,In_65,In_307);
and U967 (N_967,In_360,In_896);
nand U968 (N_968,In_619,In_781);
nor U969 (N_969,In_886,In_128);
nor U970 (N_970,In_158,In_763);
and U971 (N_971,In_981,In_188);
and U972 (N_972,In_461,In_547);
or U973 (N_973,In_558,In_871);
and U974 (N_974,In_626,In_333);
nor U975 (N_975,In_55,In_780);
and U976 (N_976,In_921,In_352);
nand U977 (N_977,In_234,In_397);
and U978 (N_978,In_542,In_165);
nand U979 (N_979,In_52,In_182);
nand U980 (N_980,In_617,In_931);
or U981 (N_981,In_997,In_730);
or U982 (N_982,In_529,In_733);
nand U983 (N_983,In_809,In_852);
or U984 (N_984,In_895,In_664);
nor U985 (N_985,In_458,In_188);
nor U986 (N_986,In_500,In_731);
or U987 (N_987,In_703,In_54);
or U988 (N_988,In_518,In_542);
and U989 (N_989,In_518,In_740);
nor U990 (N_990,In_546,In_137);
nand U991 (N_991,In_155,In_893);
or U992 (N_992,In_199,In_698);
and U993 (N_993,In_353,In_140);
xnor U994 (N_994,In_801,In_271);
nor U995 (N_995,In_241,In_538);
or U996 (N_996,In_239,In_343);
nor U997 (N_997,In_6,In_52);
and U998 (N_998,In_977,In_226);
nor U999 (N_999,In_813,In_1);
nor U1000 (N_1000,In_11,In_151);
nand U1001 (N_1001,In_156,In_902);
nand U1002 (N_1002,In_609,In_794);
nor U1003 (N_1003,In_749,In_339);
or U1004 (N_1004,In_160,In_433);
nand U1005 (N_1005,In_608,In_712);
nand U1006 (N_1006,In_424,In_525);
and U1007 (N_1007,In_453,In_944);
or U1008 (N_1008,In_434,In_638);
or U1009 (N_1009,In_67,In_528);
and U1010 (N_1010,In_940,In_818);
nor U1011 (N_1011,In_721,In_828);
or U1012 (N_1012,In_519,In_557);
nor U1013 (N_1013,In_356,In_521);
nand U1014 (N_1014,In_510,In_267);
or U1015 (N_1015,In_412,In_622);
nor U1016 (N_1016,In_258,In_822);
and U1017 (N_1017,In_162,In_863);
and U1018 (N_1018,In_829,In_948);
or U1019 (N_1019,In_295,In_830);
nor U1020 (N_1020,In_96,In_273);
and U1021 (N_1021,In_920,In_748);
or U1022 (N_1022,In_183,In_761);
nand U1023 (N_1023,In_608,In_144);
nor U1024 (N_1024,In_742,In_752);
or U1025 (N_1025,In_103,In_678);
and U1026 (N_1026,In_448,In_586);
nor U1027 (N_1027,In_372,In_399);
nor U1028 (N_1028,In_731,In_77);
nor U1029 (N_1029,In_757,In_992);
and U1030 (N_1030,In_384,In_257);
nand U1031 (N_1031,In_461,In_720);
and U1032 (N_1032,In_652,In_554);
nand U1033 (N_1033,In_274,In_129);
nor U1034 (N_1034,In_386,In_290);
nand U1035 (N_1035,In_617,In_611);
nand U1036 (N_1036,In_113,In_64);
nand U1037 (N_1037,In_315,In_34);
or U1038 (N_1038,In_841,In_961);
or U1039 (N_1039,In_752,In_53);
and U1040 (N_1040,In_311,In_354);
and U1041 (N_1041,In_690,In_657);
and U1042 (N_1042,In_797,In_396);
nor U1043 (N_1043,In_963,In_878);
nand U1044 (N_1044,In_507,In_89);
nand U1045 (N_1045,In_330,In_994);
xor U1046 (N_1046,In_427,In_387);
and U1047 (N_1047,In_727,In_981);
or U1048 (N_1048,In_223,In_301);
nor U1049 (N_1049,In_787,In_335);
or U1050 (N_1050,In_384,In_452);
nand U1051 (N_1051,In_93,In_299);
or U1052 (N_1052,In_787,In_548);
or U1053 (N_1053,In_196,In_852);
and U1054 (N_1054,In_295,In_550);
and U1055 (N_1055,In_326,In_981);
nand U1056 (N_1056,In_819,In_642);
nor U1057 (N_1057,In_234,In_213);
nand U1058 (N_1058,In_84,In_601);
nor U1059 (N_1059,In_104,In_811);
or U1060 (N_1060,In_121,In_846);
and U1061 (N_1061,In_394,In_308);
nand U1062 (N_1062,In_368,In_195);
or U1063 (N_1063,In_57,In_572);
or U1064 (N_1064,In_455,In_463);
nor U1065 (N_1065,In_802,In_528);
and U1066 (N_1066,In_462,In_909);
nor U1067 (N_1067,In_867,In_773);
nand U1068 (N_1068,In_643,In_544);
nor U1069 (N_1069,In_728,In_329);
nor U1070 (N_1070,In_28,In_79);
nor U1071 (N_1071,In_569,In_415);
or U1072 (N_1072,In_294,In_194);
and U1073 (N_1073,In_534,In_855);
nand U1074 (N_1074,In_654,In_296);
or U1075 (N_1075,In_902,In_657);
nor U1076 (N_1076,In_360,In_560);
nor U1077 (N_1077,In_808,In_1);
nand U1078 (N_1078,In_167,In_504);
nor U1079 (N_1079,In_819,In_993);
nor U1080 (N_1080,In_85,In_909);
nor U1081 (N_1081,In_791,In_815);
and U1082 (N_1082,In_853,In_786);
nand U1083 (N_1083,In_104,In_477);
and U1084 (N_1084,In_605,In_146);
nand U1085 (N_1085,In_540,In_315);
and U1086 (N_1086,In_79,In_419);
nor U1087 (N_1087,In_81,In_803);
nand U1088 (N_1088,In_9,In_306);
nor U1089 (N_1089,In_959,In_578);
and U1090 (N_1090,In_189,In_599);
and U1091 (N_1091,In_688,In_641);
nor U1092 (N_1092,In_621,In_347);
or U1093 (N_1093,In_898,In_850);
or U1094 (N_1094,In_945,In_71);
nor U1095 (N_1095,In_677,In_651);
and U1096 (N_1096,In_177,In_527);
nor U1097 (N_1097,In_242,In_474);
nand U1098 (N_1098,In_158,In_26);
nor U1099 (N_1099,In_633,In_234);
nand U1100 (N_1100,In_709,In_233);
nor U1101 (N_1101,In_196,In_242);
and U1102 (N_1102,In_767,In_593);
or U1103 (N_1103,In_614,In_981);
or U1104 (N_1104,In_754,In_93);
or U1105 (N_1105,In_727,In_188);
or U1106 (N_1106,In_260,In_908);
or U1107 (N_1107,In_912,In_321);
and U1108 (N_1108,In_443,In_743);
or U1109 (N_1109,In_266,In_694);
nor U1110 (N_1110,In_515,In_673);
or U1111 (N_1111,In_177,In_809);
nand U1112 (N_1112,In_918,In_279);
and U1113 (N_1113,In_752,In_980);
or U1114 (N_1114,In_442,In_842);
nor U1115 (N_1115,In_813,In_617);
nor U1116 (N_1116,In_219,In_864);
nor U1117 (N_1117,In_737,In_650);
nand U1118 (N_1118,In_734,In_37);
nor U1119 (N_1119,In_533,In_938);
nand U1120 (N_1120,In_439,In_839);
and U1121 (N_1121,In_64,In_398);
nand U1122 (N_1122,In_26,In_576);
or U1123 (N_1123,In_279,In_14);
nor U1124 (N_1124,In_551,In_455);
nand U1125 (N_1125,In_48,In_417);
and U1126 (N_1126,In_680,In_810);
or U1127 (N_1127,In_805,In_914);
nor U1128 (N_1128,In_329,In_62);
and U1129 (N_1129,In_690,In_562);
xnor U1130 (N_1130,In_473,In_408);
xor U1131 (N_1131,In_870,In_604);
nor U1132 (N_1132,In_171,In_366);
and U1133 (N_1133,In_971,In_335);
nand U1134 (N_1134,In_379,In_53);
and U1135 (N_1135,In_676,In_87);
or U1136 (N_1136,In_353,In_670);
nor U1137 (N_1137,In_306,In_356);
or U1138 (N_1138,In_161,In_56);
or U1139 (N_1139,In_398,In_535);
and U1140 (N_1140,In_735,In_67);
or U1141 (N_1141,In_5,In_90);
and U1142 (N_1142,In_30,In_869);
nor U1143 (N_1143,In_780,In_904);
nor U1144 (N_1144,In_355,In_705);
and U1145 (N_1145,In_538,In_523);
nor U1146 (N_1146,In_473,In_175);
nor U1147 (N_1147,In_632,In_824);
nand U1148 (N_1148,In_139,In_146);
and U1149 (N_1149,In_288,In_910);
nand U1150 (N_1150,In_246,In_862);
and U1151 (N_1151,In_776,In_727);
and U1152 (N_1152,In_691,In_887);
or U1153 (N_1153,In_498,In_82);
and U1154 (N_1154,In_884,In_261);
or U1155 (N_1155,In_43,In_704);
nand U1156 (N_1156,In_996,In_698);
and U1157 (N_1157,In_547,In_43);
and U1158 (N_1158,In_235,In_502);
and U1159 (N_1159,In_858,In_54);
nor U1160 (N_1160,In_332,In_153);
nand U1161 (N_1161,In_816,In_441);
and U1162 (N_1162,In_760,In_7);
nand U1163 (N_1163,In_572,In_63);
nand U1164 (N_1164,In_88,In_240);
nand U1165 (N_1165,In_637,In_153);
nand U1166 (N_1166,In_814,In_738);
nand U1167 (N_1167,In_736,In_150);
and U1168 (N_1168,In_237,In_74);
nor U1169 (N_1169,In_846,In_606);
nand U1170 (N_1170,In_937,In_50);
nor U1171 (N_1171,In_209,In_928);
and U1172 (N_1172,In_379,In_512);
or U1173 (N_1173,In_433,In_837);
and U1174 (N_1174,In_474,In_403);
nor U1175 (N_1175,In_529,In_671);
and U1176 (N_1176,In_513,In_576);
and U1177 (N_1177,In_376,In_810);
or U1178 (N_1178,In_251,In_668);
nand U1179 (N_1179,In_103,In_461);
nand U1180 (N_1180,In_59,In_792);
nand U1181 (N_1181,In_665,In_580);
nand U1182 (N_1182,In_188,In_651);
and U1183 (N_1183,In_777,In_512);
nand U1184 (N_1184,In_695,In_727);
or U1185 (N_1185,In_361,In_204);
nand U1186 (N_1186,In_877,In_827);
nor U1187 (N_1187,In_825,In_884);
or U1188 (N_1188,In_415,In_925);
or U1189 (N_1189,In_852,In_89);
nand U1190 (N_1190,In_107,In_585);
or U1191 (N_1191,In_29,In_168);
nor U1192 (N_1192,In_848,In_486);
and U1193 (N_1193,In_779,In_680);
nor U1194 (N_1194,In_688,In_660);
and U1195 (N_1195,In_520,In_27);
nand U1196 (N_1196,In_313,In_197);
or U1197 (N_1197,In_29,In_758);
nor U1198 (N_1198,In_510,In_636);
nand U1199 (N_1199,In_363,In_66);
or U1200 (N_1200,In_348,In_447);
nand U1201 (N_1201,In_203,In_14);
or U1202 (N_1202,In_671,In_438);
and U1203 (N_1203,In_835,In_561);
and U1204 (N_1204,In_997,In_320);
nor U1205 (N_1205,In_183,In_748);
or U1206 (N_1206,In_94,In_99);
nor U1207 (N_1207,In_982,In_823);
and U1208 (N_1208,In_796,In_75);
nand U1209 (N_1209,In_538,In_579);
and U1210 (N_1210,In_293,In_618);
and U1211 (N_1211,In_213,In_784);
nor U1212 (N_1212,In_500,In_540);
nand U1213 (N_1213,In_650,In_560);
nor U1214 (N_1214,In_725,In_439);
nor U1215 (N_1215,In_696,In_14);
xnor U1216 (N_1216,In_251,In_916);
nand U1217 (N_1217,In_287,In_478);
and U1218 (N_1218,In_743,In_543);
nor U1219 (N_1219,In_326,In_751);
nor U1220 (N_1220,In_440,In_358);
nor U1221 (N_1221,In_832,In_409);
nor U1222 (N_1222,In_685,In_409);
nand U1223 (N_1223,In_645,In_505);
and U1224 (N_1224,In_784,In_761);
nand U1225 (N_1225,In_16,In_881);
and U1226 (N_1226,In_786,In_229);
and U1227 (N_1227,In_318,In_460);
nand U1228 (N_1228,In_541,In_886);
nor U1229 (N_1229,In_205,In_543);
nand U1230 (N_1230,In_618,In_256);
nand U1231 (N_1231,In_9,In_368);
nor U1232 (N_1232,In_685,In_834);
or U1233 (N_1233,In_880,In_264);
nand U1234 (N_1234,In_50,In_456);
nor U1235 (N_1235,In_971,In_771);
nand U1236 (N_1236,In_235,In_57);
nand U1237 (N_1237,In_365,In_671);
and U1238 (N_1238,In_384,In_160);
nor U1239 (N_1239,In_454,In_449);
nor U1240 (N_1240,In_143,In_432);
and U1241 (N_1241,In_396,In_481);
nand U1242 (N_1242,In_887,In_388);
nor U1243 (N_1243,In_905,In_115);
and U1244 (N_1244,In_1,In_493);
nor U1245 (N_1245,In_778,In_169);
or U1246 (N_1246,In_118,In_422);
nor U1247 (N_1247,In_701,In_446);
xnor U1248 (N_1248,In_824,In_744);
and U1249 (N_1249,In_173,In_523);
nor U1250 (N_1250,In_121,In_802);
and U1251 (N_1251,In_485,In_797);
nor U1252 (N_1252,In_211,In_795);
nor U1253 (N_1253,In_352,In_535);
nand U1254 (N_1254,In_87,In_885);
nand U1255 (N_1255,In_746,In_404);
nand U1256 (N_1256,In_378,In_63);
nand U1257 (N_1257,In_206,In_153);
nor U1258 (N_1258,In_758,In_388);
or U1259 (N_1259,In_364,In_7);
nor U1260 (N_1260,In_31,In_961);
nand U1261 (N_1261,In_421,In_308);
or U1262 (N_1262,In_873,In_651);
nor U1263 (N_1263,In_417,In_26);
nor U1264 (N_1264,In_205,In_243);
and U1265 (N_1265,In_12,In_674);
or U1266 (N_1266,In_689,In_32);
or U1267 (N_1267,In_754,In_386);
nor U1268 (N_1268,In_745,In_546);
nand U1269 (N_1269,In_647,In_160);
nor U1270 (N_1270,In_700,In_900);
or U1271 (N_1271,In_385,In_231);
nor U1272 (N_1272,In_830,In_357);
nand U1273 (N_1273,In_429,In_184);
and U1274 (N_1274,In_959,In_753);
nor U1275 (N_1275,In_59,In_361);
and U1276 (N_1276,In_51,In_872);
and U1277 (N_1277,In_194,In_140);
nand U1278 (N_1278,In_89,In_457);
nand U1279 (N_1279,In_575,In_800);
nor U1280 (N_1280,In_598,In_189);
or U1281 (N_1281,In_248,In_599);
and U1282 (N_1282,In_403,In_881);
or U1283 (N_1283,In_216,In_105);
and U1284 (N_1284,In_191,In_301);
nor U1285 (N_1285,In_305,In_228);
or U1286 (N_1286,In_502,In_985);
nor U1287 (N_1287,In_409,In_589);
nor U1288 (N_1288,In_928,In_935);
nor U1289 (N_1289,In_702,In_200);
nor U1290 (N_1290,In_621,In_121);
and U1291 (N_1291,In_135,In_388);
nand U1292 (N_1292,In_610,In_936);
or U1293 (N_1293,In_497,In_744);
nor U1294 (N_1294,In_660,In_353);
or U1295 (N_1295,In_499,In_375);
nor U1296 (N_1296,In_826,In_409);
and U1297 (N_1297,In_619,In_268);
nor U1298 (N_1298,In_278,In_758);
or U1299 (N_1299,In_426,In_646);
nor U1300 (N_1300,In_501,In_383);
or U1301 (N_1301,In_874,In_484);
nand U1302 (N_1302,In_841,In_521);
nand U1303 (N_1303,In_425,In_805);
or U1304 (N_1304,In_78,In_705);
nand U1305 (N_1305,In_403,In_639);
or U1306 (N_1306,In_500,In_69);
or U1307 (N_1307,In_239,In_147);
nand U1308 (N_1308,In_656,In_564);
nor U1309 (N_1309,In_116,In_42);
and U1310 (N_1310,In_326,In_673);
nor U1311 (N_1311,In_904,In_764);
nand U1312 (N_1312,In_520,In_836);
nor U1313 (N_1313,In_339,In_284);
and U1314 (N_1314,In_68,In_376);
xor U1315 (N_1315,In_762,In_153);
or U1316 (N_1316,In_97,In_486);
nand U1317 (N_1317,In_233,In_753);
or U1318 (N_1318,In_287,In_938);
and U1319 (N_1319,In_826,In_434);
nor U1320 (N_1320,In_453,In_654);
or U1321 (N_1321,In_441,In_320);
nor U1322 (N_1322,In_482,In_522);
nor U1323 (N_1323,In_828,In_216);
or U1324 (N_1324,In_794,In_213);
or U1325 (N_1325,In_244,In_257);
and U1326 (N_1326,In_319,In_154);
xor U1327 (N_1327,In_873,In_136);
nand U1328 (N_1328,In_20,In_421);
nor U1329 (N_1329,In_220,In_627);
or U1330 (N_1330,In_502,In_936);
and U1331 (N_1331,In_14,In_610);
nand U1332 (N_1332,In_880,In_779);
and U1333 (N_1333,In_880,In_353);
nor U1334 (N_1334,In_376,In_529);
nor U1335 (N_1335,In_573,In_870);
nor U1336 (N_1336,In_373,In_900);
or U1337 (N_1337,In_895,In_932);
nor U1338 (N_1338,In_714,In_845);
nor U1339 (N_1339,In_679,In_321);
and U1340 (N_1340,In_93,In_982);
or U1341 (N_1341,In_464,In_820);
and U1342 (N_1342,In_905,In_706);
and U1343 (N_1343,In_803,In_901);
and U1344 (N_1344,In_625,In_233);
nor U1345 (N_1345,In_195,In_123);
nor U1346 (N_1346,In_906,In_221);
or U1347 (N_1347,In_977,In_939);
or U1348 (N_1348,In_26,In_55);
nand U1349 (N_1349,In_650,In_174);
nor U1350 (N_1350,In_258,In_78);
nand U1351 (N_1351,In_622,In_648);
nor U1352 (N_1352,In_688,In_841);
and U1353 (N_1353,In_624,In_776);
and U1354 (N_1354,In_538,In_981);
or U1355 (N_1355,In_136,In_545);
nor U1356 (N_1356,In_572,In_262);
or U1357 (N_1357,In_289,In_530);
or U1358 (N_1358,In_434,In_263);
nand U1359 (N_1359,In_916,In_62);
nand U1360 (N_1360,In_740,In_435);
nor U1361 (N_1361,In_11,In_770);
nor U1362 (N_1362,In_884,In_419);
nor U1363 (N_1363,In_48,In_282);
nand U1364 (N_1364,In_975,In_343);
and U1365 (N_1365,In_409,In_995);
or U1366 (N_1366,In_751,In_840);
nand U1367 (N_1367,In_770,In_652);
and U1368 (N_1368,In_917,In_345);
and U1369 (N_1369,In_564,In_113);
nor U1370 (N_1370,In_846,In_890);
or U1371 (N_1371,In_752,In_625);
nand U1372 (N_1372,In_411,In_921);
nand U1373 (N_1373,In_887,In_403);
nor U1374 (N_1374,In_892,In_351);
and U1375 (N_1375,In_353,In_960);
or U1376 (N_1376,In_271,In_551);
nor U1377 (N_1377,In_267,In_205);
or U1378 (N_1378,In_922,In_361);
and U1379 (N_1379,In_598,In_165);
and U1380 (N_1380,In_719,In_806);
or U1381 (N_1381,In_330,In_99);
and U1382 (N_1382,In_771,In_506);
nor U1383 (N_1383,In_623,In_714);
nor U1384 (N_1384,In_669,In_714);
and U1385 (N_1385,In_272,In_300);
nand U1386 (N_1386,In_852,In_226);
and U1387 (N_1387,In_231,In_5);
nand U1388 (N_1388,In_535,In_174);
or U1389 (N_1389,In_549,In_241);
nand U1390 (N_1390,In_713,In_984);
or U1391 (N_1391,In_739,In_817);
nand U1392 (N_1392,In_866,In_249);
and U1393 (N_1393,In_874,In_147);
or U1394 (N_1394,In_135,In_511);
nor U1395 (N_1395,In_116,In_949);
nand U1396 (N_1396,In_89,In_149);
or U1397 (N_1397,In_284,In_492);
and U1398 (N_1398,In_312,In_301);
and U1399 (N_1399,In_798,In_476);
and U1400 (N_1400,In_551,In_898);
or U1401 (N_1401,In_605,In_40);
nor U1402 (N_1402,In_663,In_782);
nand U1403 (N_1403,In_273,In_795);
nand U1404 (N_1404,In_386,In_581);
and U1405 (N_1405,In_771,In_588);
and U1406 (N_1406,In_562,In_364);
nand U1407 (N_1407,In_699,In_952);
and U1408 (N_1408,In_69,In_827);
and U1409 (N_1409,In_688,In_550);
and U1410 (N_1410,In_621,In_866);
and U1411 (N_1411,In_946,In_924);
nor U1412 (N_1412,In_140,In_83);
nand U1413 (N_1413,In_382,In_909);
nand U1414 (N_1414,In_196,In_503);
nor U1415 (N_1415,In_997,In_742);
nor U1416 (N_1416,In_151,In_844);
or U1417 (N_1417,In_984,In_892);
or U1418 (N_1418,In_685,In_659);
or U1419 (N_1419,In_326,In_518);
or U1420 (N_1420,In_715,In_809);
nor U1421 (N_1421,In_188,In_712);
nand U1422 (N_1422,In_502,In_35);
nor U1423 (N_1423,In_626,In_654);
nand U1424 (N_1424,In_915,In_627);
nor U1425 (N_1425,In_714,In_979);
nand U1426 (N_1426,In_561,In_726);
or U1427 (N_1427,In_357,In_519);
or U1428 (N_1428,In_209,In_88);
nand U1429 (N_1429,In_934,In_668);
and U1430 (N_1430,In_448,In_158);
and U1431 (N_1431,In_306,In_197);
and U1432 (N_1432,In_88,In_227);
nor U1433 (N_1433,In_308,In_742);
and U1434 (N_1434,In_672,In_791);
nand U1435 (N_1435,In_74,In_443);
nand U1436 (N_1436,In_267,In_959);
or U1437 (N_1437,In_352,In_594);
nor U1438 (N_1438,In_472,In_974);
and U1439 (N_1439,In_16,In_37);
and U1440 (N_1440,In_284,In_269);
nand U1441 (N_1441,In_939,In_107);
or U1442 (N_1442,In_510,In_788);
or U1443 (N_1443,In_349,In_884);
nor U1444 (N_1444,In_547,In_412);
or U1445 (N_1445,In_980,In_177);
or U1446 (N_1446,In_126,In_402);
nor U1447 (N_1447,In_628,In_977);
and U1448 (N_1448,In_630,In_859);
or U1449 (N_1449,In_898,In_925);
nor U1450 (N_1450,In_706,In_376);
and U1451 (N_1451,In_500,In_405);
nor U1452 (N_1452,In_477,In_668);
or U1453 (N_1453,In_607,In_458);
nand U1454 (N_1454,In_44,In_536);
nand U1455 (N_1455,In_566,In_681);
nand U1456 (N_1456,In_243,In_735);
nor U1457 (N_1457,In_339,In_225);
nor U1458 (N_1458,In_213,In_119);
nand U1459 (N_1459,In_795,In_171);
nor U1460 (N_1460,In_405,In_760);
and U1461 (N_1461,In_947,In_926);
nor U1462 (N_1462,In_516,In_857);
nand U1463 (N_1463,In_338,In_304);
or U1464 (N_1464,In_796,In_777);
and U1465 (N_1465,In_734,In_543);
or U1466 (N_1466,In_15,In_94);
or U1467 (N_1467,In_231,In_893);
nor U1468 (N_1468,In_651,In_966);
or U1469 (N_1469,In_545,In_712);
nand U1470 (N_1470,In_508,In_836);
or U1471 (N_1471,In_194,In_560);
and U1472 (N_1472,In_636,In_784);
and U1473 (N_1473,In_651,In_92);
nor U1474 (N_1474,In_447,In_35);
nor U1475 (N_1475,In_604,In_156);
nor U1476 (N_1476,In_81,In_661);
and U1477 (N_1477,In_819,In_347);
nand U1478 (N_1478,In_410,In_68);
and U1479 (N_1479,In_704,In_637);
nor U1480 (N_1480,In_35,In_183);
nand U1481 (N_1481,In_909,In_133);
nand U1482 (N_1482,In_198,In_402);
xor U1483 (N_1483,In_838,In_578);
nor U1484 (N_1484,In_895,In_780);
nand U1485 (N_1485,In_19,In_909);
and U1486 (N_1486,In_444,In_80);
or U1487 (N_1487,In_830,In_666);
nand U1488 (N_1488,In_32,In_241);
or U1489 (N_1489,In_866,In_864);
and U1490 (N_1490,In_497,In_614);
or U1491 (N_1491,In_501,In_831);
nor U1492 (N_1492,In_823,In_331);
and U1493 (N_1493,In_482,In_257);
nor U1494 (N_1494,In_691,In_21);
or U1495 (N_1495,In_141,In_951);
and U1496 (N_1496,In_449,In_292);
xnor U1497 (N_1497,In_278,In_188);
nand U1498 (N_1498,In_363,In_411);
nand U1499 (N_1499,In_753,In_921);
and U1500 (N_1500,In_591,In_648);
nand U1501 (N_1501,In_821,In_553);
and U1502 (N_1502,In_946,In_881);
and U1503 (N_1503,In_531,In_867);
and U1504 (N_1504,In_523,In_861);
and U1505 (N_1505,In_988,In_430);
or U1506 (N_1506,In_200,In_397);
and U1507 (N_1507,In_168,In_514);
or U1508 (N_1508,In_198,In_270);
and U1509 (N_1509,In_477,In_789);
nor U1510 (N_1510,In_562,In_31);
or U1511 (N_1511,In_232,In_435);
nor U1512 (N_1512,In_762,In_44);
and U1513 (N_1513,In_132,In_850);
nor U1514 (N_1514,In_571,In_874);
nand U1515 (N_1515,In_269,In_293);
nand U1516 (N_1516,In_914,In_744);
or U1517 (N_1517,In_670,In_915);
and U1518 (N_1518,In_29,In_583);
and U1519 (N_1519,In_90,In_604);
nand U1520 (N_1520,In_491,In_134);
nand U1521 (N_1521,In_447,In_634);
or U1522 (N_1522,In_383,In_819);
and U1523 (N_1523,In_202,In_697);
or U1524 (N_1524,In_646,In_849);
and U1525 (N_1525,In_329,In_722);
and U1526 (N_1526,In_950,In_898);
nor U1527 (N_1527,In_943,In_186);
and U1528 (N_1528,In_570,In_24);
nor U1529 (N_1529,In_843,In_947);
or U1530 (N_1530,In_719,In_774);
or U1531 (N_1531,In_257,In_81);
nand U1532 (N_1532,In_549,In_566);
nor U1533 (N_1533,In_455,In_784);
and U1534 (N_1534,In_600,In_138);
or U1535 (N_1535,In_49,In_538);
nand U1536 (N_1536,In_857,In_503);
and U1537 (N_1537,In_96,In_205);
or U1538 (N_1538,In_378,In_201);
and U1539 (N_1539,In_183,In_697);
nand U1540 (N_1540,In_505,In_89);
and U1541 (N_1541,In_996,In_744);
or U1542 (N_1542,In_195,In_746);
and U1543 (N_1543,In_99,In_275);
or U1544 (N_1544,In_476,In_761);
or U1545 (N_1545,In_582,In_68);
nand U1546 (N_1546,In_206,In_847);
nor U1547 (N_1547,In_352,In_61);
or U1548 (N_1548,In_911,In_968);
or U1549 (N_1549,In_415,In_990);
and U1550 (N_1550,In_49,In_976);
or U1551 (N_1551,In_953,In_419);
or U1552 (N_1552,In_614,In_898);
or U1553 (N_1553,In_137,In_815);
and U1554 (N_1554,In_74,In_976);
and U1555 (N_1555,In_454,In_419);
nand U1556 (N_1556,In_883,In_969);
or U1557 (N_1557,In_811,In_886);
nand U1558 (N_1558,In_155,In_345);
nand U1559 (N_1559,In_710,In_566);
or U1560 (N_1560,In_879,In_838);
and U1561 (N_1561,In_486,In_69);
or U1562 (N_1562,In_267,In_83);
nor U1563 (N_1563,In_317,In_356);
nand U1564 (N_1564,In_502,In_761);
and U1565 (N_1565,In_527,In_396);
and U1566 (N_1566,In_419,In_732);
and U1567 (N_1567,In_142,In_87);
and U1568 (N_1568,In_275,In_218);
and U1569 (N_1569,In_120,In_544);
or U1570 (N_1570,In_871,In_554);
nand U1571 (N_1571,In_740,In_278);
nand U1572 (N_1572,In_651,In_956);
nand U1573 (N_1573,In_631,In_603);
nor U1574 (N_1574,In_488,In_183);
nor U1575 (N_1575,In_664,In_554);
nand U1576 (N_1576,In_822,In_766);
nor U1577 (N_1577,In_495,In_154);
and U1578 (N_1578,In_42,In_600);
nand U1579 (N_1579,In_556,In_695);
nor U1580 (N_1580,In_381,In_547);
nand U1581 (N_1581,In_49,In_872);
nor U1582 (N_1582,In_479,In_664);
nand U1583 (N_1583,In_3,In_226);
or U1584 (N_1584,In_618,In_113);
or U1585 (N_1585,In_684,In_111);
nor U1586 (N_1586,In_919,In_589);
and U1587 (N_1587,In_261,In_174);
nor U1588 (N_1588,In_590,In_270);
or U1589 (N_1589,In_761,In_473);
nand U1590 (N_1590,In_782,In_762);
and U1591 (N_1591,In_849,In_195);
or U1592 (N_1592,In_331,In_396);
nor U1593 (N_1593,In_729,In_342);
nor U1594 (N_1594,In_995,In_208);
nand U1595 (N_1595,In_826,In_701);
and U1596 (N_1596,In_572,In_369);
and U1597 (N_1597,In_215,In_451);
nand U1598 (N_1598,In_73,In_49);
or U1599 (N_1599,In_27,In_170);
or U1600 (N_1600,In_191,In_271);
xor U1601 (N_1601,In_143,In_390);
and U1602 (N_1602,In_0,In_168);
nor U1603 (N_1603,In_118,In_297);
nand U1604 (N_1604,In_357,In_649);
nand U1605 (N_1605,In_116,In_941);
nor U1606 (N_1606,In_382,In_645);
nor U1607 (N_1607,In_129,In_179);
nand U1608 (N_1608,In_648,In_838);
or U1609 (N_1609,In_37,In_229);
or U1610 (N_1610,In_556,In_308);
or U1611 (N_1611,In_986,In_239);
or U1612 (N_1612,In_871,In_628);
nand U1613 (N_1613,In_613,In_272);
and U1614 (N_1614,In_262,In_831);
nand U1615 (N_1615,In_788,In_961);
and U1616 (N_1616,In_511,In_306);
xor U1617 (N_1617,In_830,In_179);
nor U1618 (N_1618,In_62,In_127);
nand U1619 (N_1619,In_99,In_809);
and U1620 (N_1620,In_183,In_787);
nand U1621 (N_1621,In_941,In_780);
and U1622 (N_1622,In_695,In_412);
and U1623 (N_1623,In_787,In_539);
nor U1624 (N_1624,In_159,In_629);
nand U1625 (N_1625,In_976,In_100);
nor U1626 (N_1626,In_532,In_36);
nand U1627 (N_1627,In_736,In_131);
nand U1628 (N_1628,In_288,In_924);
or U1629 (N_1629,In_547,In_244);
and U1630 (N_1630,In_245,In_332);
nor U1631 (N_1631,In_45,In_409);
nand U1632 (N_1632,In_622,In_736);
nand U1633 (N_1633,In_948,In_337);
nor U1634 (N_1634,In_958,In_438);
xor U1635 (N_1635,In_333,In_715);
nor U1636 (N_1636,In_166,In_700);
and U1637 (N_1637,In_580,In_206);
and U1638 (N_1638,In_864,In_934);
nand U1639 (N_1639,In_121,In_364);
nand U1640 (N_1640,In_237,In_851);
nor U1641 (N_1641,In_585,In_154);
nor U1642 (N_1642,In_921,In_797);
or U1643 (N_1643,In_247,In_241);
nor U1644 (N_1644,In_482,In_399);
or U1645 (N_1645,In_922,In_231);
and U1646 (N_1646,In_449,In_9);
or U1647 (N_1647,In_158,In_101);
nor U1648 (N_1648,In_628,In_936);
and U1649 (N_1649,In_726,In_810);
and U1650 (N_1650,In_972,In_213);
and U1651 (N_1651,In_378,In_542);
nor U1652 (N_1652,In_825,In_667);
nand U1653 (N_1653,In_590,In_634);
nor U1654 (N_1654,In_964,In_955);
nor U1655 (N_1655,In_328,In_574);
nor U1656 (N_1656,In_367,In_144);
nor U1657 (N_1657,In_391,In_318);
and U1658 (N_1658,In_98,In_140);
nor U1659 (N_1659,In_227,In_609);
nor U1660 (N_1660,In_711,In_103);
nand U1661 (N_1661,In_848,In_141);
or U1662 (N_1662,In_617,In_439);
and U1663 (N_1663,In_955,In_12);
or U1664 (N_1664,In_671,In_684);
and U1665 (N_1665,In_636,In_788);
nand U1666 (N_1666,In_751,In_545);
nand U1667 (N_1667,In_514,In_522);
nand U1668 (N_1668,In_145,In_793);
or U1669 (N_1669,In_138,In_78);
or U1670 (N_1670,In_87,In_739);
nor U1671 (N_1671,In_584,In_991);
nor U1672 (N_1672,In_714,In_399);
nor U1673 (N_1673,In_691,In_698);
nor U1674 (N_1674,In_638,In_232);
nand U1675 (N_1675,In_827,In_385);
nor U1676 (N_1676,In_114,In_382);
or U1677 (N_1677,In_5,In_336);
or U1678 (N_1678,In_956,In_733);
nor U1679 (N_1679,In_819,In_6);
nor U1680 (N_1680,In_259,In_928);
nor U1681 (N_1681,In_915,In_663);
and U1682 (N_1682,In_369,In_844);
or U1683 (N_1683,In_336,In_907);
nor U1684 (N_1684,In_464,In_341);
or U1685 (N_1685,In_431,In_632);
or U1686 (N_1686,In_445,In_772);
and U1687 (N_1687,In_762,In_382);
and U1688 (N_1688,In_860,In_164);
nor U1689 (N_1689,In_233,In_832);
nand U1690 (N_1690,In_66,In_638);
nor U1691 (N_1691,In_186,In_799);
and U1692 (N_1692,In_500,In_62);
nand U1693 (N_1693,In_888,In_400);
nand U1694 (N_1694,In_147,In_931);
and U1695 (N_1695,In_323,In_336);
or U1696 (N_1696,In_740,In_239);
nand U1697 (N_1697,In_760,In_742);
and U1698 (N_1698,In_957,In_804);
nand U1699 (N_1699,In_71,In_892);
and U1700 (N_1700,In_768,In_624);
nor U1701 (N_1701,In_647,In_197);
and U1702 (N_1702,In_608,In_810);
nor U1703 (N_1703,In_884,In_339);
and U1704 (N_1704,In_555,In_497);
or U1705 (N_1705,In_818,In_643);
nor U1706 (N_1706,In_514,In_716);
nand U1707 (N_1707,In_708,In_700);
and U1708 (N_1708,In_426,In_820);
and U1709 (N_1709,In_774,In_510);
nand U1710 (N_1710,In_471,In_582);
xnor U1711 (N_1711,In_817,In_461);
nand U1712 (N_1712,In_606,In_291);
or U1713 (N_1713,In_472,In_352);
and U1714 (N_1714,In_399,In_282);
and U1715 (N_1715,In_399,In_967);
and U1716 (N_1716,In_272,In_22);
or U1717 (N_1717,In_328,In_77);
and U1718 (N_1718,In_434,In_20);
nand U1719 (N_1719,In_557,In_914);
or U1720 (N_1720,In_683,In_78);
or U1721 (N_1721,In_890,In_231);
nor U1722 (N_1722,In_646,In_5);
or U1723 (N_1723,In_55,In_970);
or U1724 (N_1724,In_599,In_768);
or U1725 (N_1725,In_977,In_24);
or U1726 (N_1726,In_491,In_669);
nand U1727 (N_1727,In_623,In_478);
nand U1728 (N_1728,In_140,In_101);
nand U1729 (N_1729,In_879,In_120);
nor U1730 (N_1730,In_572,In_221);
and U1731 (N_1731,In_52,In_402);
and U1732 (N_1732,In_469,In_926);
nand U1733 (N_1733,In_615,In_62);
nand U1734 (N_1734,In_970,In_96);
or U1735 (N_1735,In_221,In_561);
and U1736 (N_1736,In_52,In_469);
nand U1737 (N_1737,In_470,In_841);
nand U1738 (N_1738,In_414,In_343);
or U1739 (N_1739,In_555,In_768);
nor U1740 (N_1740,In_576,In_198);
and U1741 (N_1741,In_342,In_768);
nor U1742 (N_1742,In_770,In_673);
nand U1743 (N_1743,In_897,In_236);
and U1744 (N_1744,In_71,In_329);
or U1745 (N_1745,In_106,In_597);
nand U1746 (N_1746,In_893,In_82);
nand U1747 (N_1747,In_1,In_654);
or U1748 (N_1748,In_496,In_564);
nand U1749 (N_1749,In_563,In_480);
or U1750 (N_1750,In_549,In_245);
nor U1751 (N_1751,In_888,In_752);
nand U1752 (N_1752,In_652,In_502);
nor U1753 (N_1753,In_930,In_32);
and U1754 (N_1754,In_793,In_146);
or U1755 (N_1755,In_3,In_965);
and U1756 (N_1756,In_81,In_169);
or U1757 (N_1757,In_298,In_165);
nand U1758 (N_1758,In_657,In_262);
or U1759 (N_1759,In_454,In_990);
or U1760 (N_1760,In_145,In_700);
nand U1761 (N_1761,In_538,In_475);
nor U1762 (N_1762,In_674,In_957);
and U1763 (N_1763,In_336,In_119);
or U1764 (N_1764,In_533,In_216);
nand U1765 (N_1765,In_886,In_195);
nor U1766 (N_1766,In_28,In_466);
nor U1767 (N_1767,In_559,In_841);
and U1768 (N_1768,In_363,In_833);
and U1769 (N_1769,In_9,In_4);
or U1770 (N_1770,In_937,In_865);
nand U1771 (N_1771,In_313,In_566);
or U1772 (N_1772,In_998,In_519);
and U1773 (N_1773,In_538,In_60);
and U1774 (N_1774,In_134,In_566);
and U1775 (N_1775,In_194,In_823);
nand U1776 (N_1776,In_820,In_508);
or U1777 (N_1777,In_703,In_877);
xor U1778 (N_1778,In_749,In_336);
and U1779 (N_1779,In_345,In_812);
nand U1780 (N_1780,In_608,In_878);
and U1781 (N_1781,In_292,In_667);
and U1782 (N_1782,In_800,In_65);
or U1783 (N_1783,In_933,In_404);
nor U1784 (N_1784,In_864,In_659);
nand U1785 (N_1785,In_927,In_935);
nor U1786 (N_1786,In_683,In_113);
nand U1787 (N_1787,In_827,In_28);
nand U1788 (N_1788,In_747,In_297);
or U1789 (N_1789,In_512,In_436);
nor U1790 (N_1790,In_535,In_908);
nand U1791 (N_1791,In_297,In_170);
or U1792 (N_1792,In_576,In_214);
or U1793 (N_1793,In_656,In_258);
and U1794 (N_1794,In_338,In_895);
or U1795 (N_1795,In_52,In_602);
and U1796 (N_1796,In_0,In_759);
nand U1797 (N_1797,In_800,In_335);
and U1798 (N_1798,In_105,In_239);
or U1799 (N_1799,In_787,In_865);
nor U1800 (N_1800,In_997,In_155);
and U1801 (N_1801,In_280,In_887);
nor U1802 (N_1802,In_697,In_311);
nand U1803 (N_1803,In_781,In_737);
and U1804 (N_1804,In_195,In_662);
nand U1805 (N_1805,In_649,In_399);
nand U1806 (N_1806,In_4,In_912);
nor U1807 (N_1807,In_67,In_248);
and U1808 (N_1808,In_325,In_931);
or U1809 (N_1809,In_789,In_310);
and U1810 (N_1810,In_205,In_956);
nor U1811 (N_1811,In_80,In_180);
and U1812 (N_1812,In_163,In_621);
and U1813 (N_1813,In_179,In_635);
nand U1814 (N_1814,In_343,In_741);
xnor U1815 (N_1815,In_26,In_829);
nor U1816 (N_1816,In_391,In_596);
and U1817 (N_1817,In_646,In_942);
nand U1818 (N_1818,In_97,In_96);
or U1819 (N_1819,In_900,In_734);
and U1820 (N_1820,In_344,In_270);
or U1821 (N_1821,In_986,In_957);
and U1822 (N_1822,In_82,In_169);
nand U1823 (N_1823,In_821,In_714);
nand U1824 (N_1824,In_9,In_977);
or U1825 (N_1825,In_526,In_799);
or U1826 (N_1826,In_68,In_49);
nand U1827 (N_1827,In_488,In_103);
or U1828 (N_1828,In_205,In_412);
nor U1829 (N_1829,In_556,In_271);
nand U1830 (N_1830,In_793,In_285);
nor U1831 (N_1831,In_274,In_609);
or U1832 (N_1832,In_280,In_430);
and U1833 (N_1833,In_143,In_227);
nor U1834 (N_1834,In_370,In_65);
and U1835 (N_1835,In_581,In_304);
nor U1836 (N_1836,In_297,In_271);
nor U1837 (N_1837,In_141,In_384);
or U1838 (N_1838,In_703,In_475);
and U1839 (N_1839,In_667,In_978);
nor U1840 (N_1840,In_847,In_859);
and U1841 (N_1841,In_444,In_241);
nor U1842 (N_1842,In_11,In_531);
nor U1843 (N_1843,In_350,In_880);
nand U1844 (N_1844,In_714,In_520);
or U1845 (N_1845,In_239,In_842);
nor U1846 (N_1846,In_166,In_722);
or U1847 (N_1847,In_88,In_788);
nor U1848 (N_1848,In_581,In_870);
nand U1849 (N_1849,In_514,In_255);
or U1850 (N_1850,In_19,In_591);
or U1851 (N_1851,In_856,In_362);
nand U1852 (N_1852,In_196,In_641);
and U1853 (N_1853,In_694,In_156);
and U1854 (N_1854,In_764,In_560);
nand U1855 (N_1855,In_561,In_49);
nor U1856 (N_1856,In_875,In_788);
or U1857 (N_1857,In_365,In_207);
and U1858 (N_1858,In_283,In_984);
and U1859 (N_1859,In_573,In_27);
nor U1860 (N_1860,In_507,In_611);
and U1861 (N_1861,In_948,In_224);
and U1862 (N_1862,In_395,In_342);
and U1863 (N_1863,In_857,In_182);
nand U1864 (N_1864,In_275,In_191);
nor U1865 (N_1865,In_907,In_835);
or U1866 (N_1866,In_413,In_20);
nand U1867 (N_1867,In_378,In_902);
nor U1868 (N_1868,In_402,In_398);
nor U1869 (N_1869,In_313,In_181);
or U1870 (N_1870,In_771,In_668);
nor U1871 (N_1871,In_225,In_351);
or U1872 (N_1872,In_574,In_265);
nand U1873 (N_1873,In_895,In_578);
nand U1874 (N_1874,In_142,In_576);
nand U1875 (N_1875,In_447,In_43);
and U1876 (N_1876,In_130,In_286);
and U1877 (N_1877,In_511,In_784);
and U1878 (N_1878,In_799,In_80);
nor U1879 (N_1879,In_985,In_878);
nor U1880 (N_1880,In_814,In_423);
nand U1881 (N_1881,In_609,In_396);
nor U1882 (N_1882,In_864,In_243);
and U1883 (N_1883,In_775,In_771);
or U1884 (N_1884,In_514,In_778);
nand U1885 (N_1885,In_489,In_996);
or U1886 (N_1886,In_334,In_56);
nor U1887 (N_1887,In_130,In_442);
or U1888 (N_1888,In_241,In_80);
and U1889 (N_1889,In_530,In_643);
nand U1890 (N_1890,In_531,In_849);
or U1891 (N_1891,In_127,In_341);
nand U1892 (N_1892,In_131,In_830);
and U1893 (N_1893,In_588,In_708);
or U1894 (N_1894,In_133,In_577);
or U1895 (N_1895,In_792,In_590);
nand U1896 (N_1896,In_375,In_305);
nand U1897 (N_1897,In_149,In_778);
and U1898 (N_1898,In_909,In_585);
and U1899 (N_1899,In_279,In_17);
or U1900 (N_1900,In_531,In_301);
nor U1901 (N_1901,In_775,In_585);
or U1902 (N_1902,In_579,In_624);
or U1903 (N_1903,In_933,In_156);
xor U1904 (N_1904,In_6,In_196);
and U1905 (N_1905,In_304,In_275);
and U1906 (N_1906,In_344,In_929);
nand U1907 (N_1907,In_3,In_496);
or U1908 (N_1908,In_429,In_582);
and U1909 (N_1909,In_102,In_869);
or U1910 (N_1910,In_391,In_271);
xor U1911 (N_1911,In_748,In_841);
or U1912 (N_1912,In_224,In_55);
or U1913 (N_1913,In_371,In_282);
or U1914 (N_1914,In_564,In_753);
nand U1915 (N_1915,In_557,In_438);
nand U1916 (N_1916,In_220,In_559);
nand U1917 (N_1917,In_6,In_568);
nand U1918 (N_1918,In_303,In_176);
nand U1919 (N_1919,In_535,In_780);
nor U1920 (N_1920,In_281,In_107);
and U1921 (N_1921,In_270,In_908);
nor U1922 (N_1922,In_366,In_637);
and U1923 (N_1923,In_205,In_492);
or U1924 (N_1924,In_449,In_992);
nand U1925 (N_1925,In_385,In_801);
nand U1926 (N_1926,In_587,In_164);
nor U1927 (N_1927,In_693,In_947);
nand U1928 (N_1928,In_480,In_697);
nand U1929 (N_1929,In_830,In_989);
nand U1930 (N_1930,In_415,In_586);
or U1931 (N_1931,In_377,In_734);
xnor U1932 (N_1932,In_935,In_286);
and U1933 (N_1933,In_385,In_799);
nand U1934 (N_1934,In_11,In_544);
or U1935 (N_1935,In_479,In_909);
and U1936 (N_1936,In_483,In_191);
nand U1937 (N_1937,In_496,In_982);
nor U1938 (N_1938,In_840,In_649);
or U1939 (N_1939,In_137,In_773);
or U1940 (N_1940,In_488,In_562);
and U1941 (N_1941,In_749,In_601);
nand U1942 (N_1942,In_625,In_990);
and U1943 (N_1943,In_984,In_65);
or U1944 (N_1944,In_72,In_389);
or U1945 (N_1945,In_869,In_932);
nand U1946 (N_1946,In_976,In_572);
or U1947 (N_1947,In_856,In_731);
nand U1948 (N_1948,In_293,In_433);
or U1949 (N_1949,In_849,In_803);
and U1950 (N_1950,In_452,In_110);
or U1951 (N_1951,In_595,In_837);
or U1952 (N_1952,In_930,In_554);
nand U1953 (N_1953,In_848,In_200);
nand U1954 (N_1954,In_230,In_715);
and U1955 (N_1955,In_168,In_358);
or U1956 (N_1956,In_292,In_129);
nand U1957 (N_1957,In_380,In_312);
and U1958 (N_1958,In_691,In_756);
and U1959 (N_1959,In_328,In_526);
nand U1960 (N_1960,In_935,In_211);
or U1961 (N_1961,In_110,In_744);
or U1962 (N_1962,In_356,In_755);
and U1963 (N_1963,In_776,In_366);
nor U1964 (N_1964,In_264,In_906);
or U1965 (N_1965,In_673,In_174);
nand U1966 (N_1966,In_906,In_258);
or U1967 (N_1967,In_143,In_877);
nand U1968 (N_1968,In_331,In_766);
nor U1969 (N_1969,In_924,In_733);
and U1970 (N_1970,In_35,In_403);
or U1971 (N_1971,In_335,In_39);
or U1972 (N_1972,In_877,In_646);
or U1973 (N_1973,In_73,In_831);
and U1974 (N_1974,In_257,In_643);
or U1975 (N_1975,In_160,In_667);
and U1976 (N_1976,In_480,In_371);
nor U1977 (N_1977,In_171,In_476);
and U1978 (N_1978,In_295,In_502);
or U1979 (N_1979,In_276,In_420);
nor U1980 (N_1980,In_15,In_833);
and U1981 (N_1981,In_994,In_183);
or U1982 (N_1982,In_53,In_523);
or U1983 (N_1983,In_203,In_801);
nor U1984 (N_1984,In_579,In_617);
nand U1985 (N_1985,In_435,In_261);
and U1986 (N_1986,In_11,In_103);
nand U1987 (N_1987,In_55,In_948);
nor U1988 (N_1988,In_109,In_636);
or U1989 (N_1989,In_24,In_292);
or U1990 (N_1990,In_166,In_615);
nand U1991 (N_1991,In_591,In_330);
xnor U1992 (N_1992,In_383,In_673);
nand U1993 (N_1993,In_224,In_1);
nand U1994 (N_1994,In_443,In_62);
and U1995 (N_1995,In_56,In_667);
nand U1996 (N_1996,In_204,In_794);
nor U1997 (N_1997,In_488,In_380);
nor U1998 (N_1998,In_111,In_422);
and U1999 (N_1999,In_265,In_429);
or U2000 (N_2000,In_999,In_235);
nor U2001 (N_2001,In_82,In_983);
and U2002 (N_2002,In_160,In_850);
xnor U2003 (N_2003,In_8,In_423);
nand U2004 (N_2004,In_782,In_444);
or U2005 (N_2005,In_668,In_935);
nor U2006 (N_2006,In_87,In_550);
nor U2007 (N_2007,In_829,In_839);
nand U2008 (N_2008,In_922,In_983);
nand U2009 (N_2009,In_188,In_86);
or U2010 (N_2010,In_957,In_590);
or U2011 (N_2011,In_602,In_197);
or U2012 (N_2012,In_190,In_287);
and U2013 (N_2013,In_401,In_646);
nor U2014 (N_2014,In_85,In_950);
nand U2015 (N_2015,In_261,In_448);
or U2016 (N_2016,In_375,In_457);
or U2017 (N_2017,In_504,In_402);
nand U2018 (N_2018,In_189,In_211);
and U2019 (N_2019,In_149,In_12);
nor U2020 (N_2020,In_735,In_740);
nand U2021 (N_2021,In_990,In_654);
nand U2022 (N_2022,In_813,In_491);
or U2023 (N_2023,In_676,In_763);
or U2024 (N_2024,In_710,In_897);
and U2025 (N_2025,In_244,In_874);
and U2026 (N_2026,In_361,In_669);
nand U2027 (N_2027,In_548,In_174);
or U2028 (N_2028,In_272,In_199);
or U2029 (N_2029,In_243,In_239);
and U2030 (N_2030,In_123,In_522);
and U2031 (N_2031,In_864,In_207);
or U2032 (N_2032,In_590,In_565);
nand U2033 (N_2033,In_919,In_412);
and U2034 (N_2034,In_1,In_527);
nor U2035 (N_2035,In_38,In_650);
nand U2036 (N_2036,In_475,In_465);
and U2037 (N_2037,In_246,In_941);
nand U2038 (N_2038,In_606,In_134);
nand U2039 (N_2039,In_990,In_464);
or U2040 (N_2040,In_16,In_323);
or U2041 (N_2041,In_588,In_69);
and U2042 (N_2042,In_346,In_495);
nor U2043 (N_2043,In_931,In_753);
nor U2044 (N_2044,In_790,In_976);
and U2045 (N_2045,In_426,In_371);
or U2046 (N_2046,In_831,In_925);
or U2047 (N_2047,In_586,In_663);
or U2048 (N_2048,In_717,In_432);
nor U2049 (N_2049,In_398,In_465);
nand U2050 (N_2050,In_375,In_917);
and U2051 (N_2051,In_219,In_618);
or U2052 (N_2052,In_702,In_21);
and U2053 (N_2053,In_471,In_681);
nand U2054 (N_2054,In_737,In_189);
nand U2055 (N_2055,In_267,In_982);
xor U2056 (N_2056,In_779,In_893);
and U2057 (N_2057,In_831,In_159);
nor U2058 (N_2058,In_212,In_436);
or U2059 (N_2059,In_689,In_589);
and U2060 (N_2060,In_481,In_935);
nand U2061 (N_2061,In_621,In_381);
and U2062 (N_2062,In_229,In_407);
nor U2063 (N_2063,In_981,In_172);
or U2064 (N_2064,In_327,In_179);
or U2065 (N_2065,In_977,In_215);
nor U2066 (N_2066,In_415,In_89);
nor U2067 (N_2067,In_867,In_736);
nand U2068 (N_2068,In_803,In_907);
or U2069 (N_2069,In_138,In_77);
nor U2070 (N_2070,In_779,In_999);
or U2071 (N_2071,In_22,In_470);
or U2072 (N_2072,In_478,In_56);
nor U2073 (N_2073,In_117,In_446);
nor U2074 (N_2074,In_399,In_23);
and U2075 (N_2075,In_836,In_532);
nor U2076 (N_2076,In_759,In_995);
nor U2077 (N_2077,In_961,In_350);
and U2078 (N_2078,In_794,In_774);
nor U2079 (N_2079,In_505,In_346);
and U2080 (N_2080,In_935,In_257);
nand U2081 (N_2081,In_550,In_630);
nand U2082 (N_2082,In_680,In_539);
nand U2083 (N_2083,In_360,In_373);
nand U2084 (N_2084,In_375,In_654);
nand U2085 (N_2085,In_459,In_188);
nand U2086 (N_2086,In_474,In_624);
nor U2087 (N_2087,In_506,In_802);
and U2088 (N_2088,In_321,In_739);
or U2089 (N_2089,In_972,In_652);
and U2090 (N_2090,In_551,In_267);
or U2091 (N_2091,In_897,In_464);
nand U2092 (N_2092,In_979,In_421);
or U2093 (N_2093,In_960,In_511);
nor U2094 (N_2094,In_55,In_633);
nand U2095 (N_2095,In_346,In_626);
or U2096 (N_2096,In_910,In_664);
nor U2097 (N_2097,In_462,In_860);
nor U2098 (N_2098,In_465,In_502);
nor U2099 (N_2099,In_996,In_214);
nor U2100 (N_2100,In_361,In_138);
nand U2101 (N_2101,In_280,In_721);
nand U2102 (N_2102,In_960,In_658);
nand U2103 (N_2103,In_416,In_740);
and U2104 (N_2104,In_82,In_885);
nor U2105 (N_2105,In_398,In_506);
or U2106 (N_2106,In_953,In_305);
nor U2107 (N_2107,In_459,In_789);
and U2108 (N_2108,In_600,In_636);
or U2109 (N_2109,In_152,In_640);
or U2110 (N_2110,In_933,In_361);
and U2111 (N_2111,In_621,In_322);
and U2112 (N_2112,In_414,In_684);
and U2113 (N_2113,In_470,In_435);
and U2114 (N_2114,In_883,In_600);
nor U2115 (N_2115,In_119,In_161);
nor U2116 (N_2116,In_221,In_674);
nand U2117 (N_2117,In_743,In_306);
nor U2118 (N_2118,In_928,In_871);
nor U2119 (N_2119,In_273,In_686);
or U2120 (N_2120,In_223,In_110);
nor U2121 (N_2121,In_549,In_4);
nand U2122 (N_2122,In_591,In_109);
nor U2123 (N_2123,In_429,In_832);
nor U2124 (N_2124,In_546,In_236);
nand U2125 (N_2125,In_867,In_335);
nor U2126 (N_2126,In_657,In_26);
nor U2127 (N_2127,In_247,In_985);
nor U2128 (N_2128,In_851,In_300);
and U2129 (N_2129,In_285,In_764);
nor U2130 (N_2130,In_886,In_526);
nand U2131 (N_2131,In_845,In_33);
and U2132 (N_2132,In_596,In_910);
nand U2133 (N_2133,In_695,In_704);
or U2134 (N_2134,In_528,In_984);
and U2135 (N_2135,In_0,In_600);
nand U2136 (N_2136,In_255,In_430);
or U2137 (N_2137,In_742,In_357);
nand U2138 (N_2138,In_228,In_738);
nor U2139 (N_2139,In_247,In_662);
and U2140 (N_2140,In_131,In_557);
nand U2141 (N_2141,In_400,In_967);
nor U2142 (N_2142,In_519,In_533);
or U2143 (N_2143,In_607,In_66);
or U2144 (N_2144,In_127,In_160);
nor U2145 (N_2145,In_769,In_135);
nand U2146 (N_2146,In_650,In_891);
or U2147 (N_2147,In_605,In_104);
nor U2148 (N_2148,In_100,In_131);
and U2149 (N_2149,In_260,In_11);
nor U2150 (N_2150,In_879,In_166);
or U2151 (N_2151,In_174,In_134);
nand U2152 (N_2152,In_899,In_560);
and U2153 (N_2153,In_31,In_439);
and U2154 (N_2154,In_548,In_673);
nand U2155 (N_2155,In_177,In_541);
and U2156 (N_2156,In_676,In_316);
and U2157 (N_2157,In_918,In_20);
or U2158 (N_2158,In_968,In_504);
nor U2159 (N_2159,In_48,In_623);
nand U2160 (N_2160,In_52,In_919);
or U2161 (N_2161,In_550,In_220);
xnor U2162 (N_2162,In_327,In_341);
or U2163 (N_2163,In_772,In_623);
or U2164 (N_2164,In_542,In_344);
and U2165 (N_2165,In_445,In_446);
nor U2166 (N_2166,In_43,In_485);
nor U2167 (N_2167,In_656,In_138);
and U2168 (N_2168,In_478,In_790);
and U2169 (N_2169,In_668,In_198);
nand U2170 (N_2170,In_696,In_131);
nand U2171 (N_2171,In_276,In_19);
nor U2172 (N_2172,In_339,In_549);
or U2173 (N_2173,In_377,In_868);
nand U2174 (N_2174,In_926,In_259);
nand U2175 (N_2175,In_421,In_61);
and U2176 (N_2176,In_170,In_1);
and U2177 (N_2177,In_55,In_336);
nand U2178 (N_2178,In_307,In_602);
nand U2179 (N_2179,In_933,In_602);
and U2180 (N_2180,In_622,In_658);
and U2181 (N_2181,In_203,In_264);
and U2182 (N_2182,In_874,In_414);
nand U2183 (N_2183,In_909,In_38);
or U2184 (N_2184,In_280,In_801);
nor U2185 (N_2185,In_281,In_706);
or U2186 (N_2186,In_185,In_145);
and U2187 (N_2187,In_297,In_384);
and U2188 (N_2188,In_248,In_394);
nor U2189 (N_2189,In_146,In_588);
nand U2190 (N_2190,In_495,In_409);
or U2191 (N_2191,In_993,In_624);
and U2192 (N_2192,In_782,In_360);
or U2193 (N_2193,In_72,In_680);
and U2194 (N_2194,In_845,In_110);
nand U2195 (N_2195,In_922,In_851);
nand U2196 (N_2196,In_31,In_797);
and U2197 (N_2197,In_584,In_349);
or U2198 (N_2198,In_519,In_342);
nor U2199 (N_2199,In_597,In_369);
nor U2200 (N_2200,In_625,In_453);
and U2201 (N_2201,In_754,In_436);
and U2202 (N_2202,In_494,In_152);
nand U2203 (N_2203,In_339,In_818);
and U2204 (N_2204,In_228,In_732);
or U2205 (N_2205,In_227,In_194);
nor U2206 (N_2206,In_692,In_191);
nor U2207 (N_2207,In_937,In_822);
nor U2208 (N_2208,In_680,In_484);
or U2209 (N_2209,In_100,In_281);
or U2210 (N_2210,In_231,In_874);
and U2211 (N_2211,In_432,In_321);
nor U2212 (N_2212,In_921,In_731);
nand U2213 (N_2213,In_25,In_845);
or U2214 (N_2214,In_753,In_533);
nand U2215 (N_2215,In_768,In_605);
nand U2216 (N_2216,In_667,In_29);
nand U2217 (N_2217,In_461,In_666);
and U2218 (N_2218,In_806,In_359);
or U2219 (N_2219,In_864,In_184);
nor U2220 (N_2220,In_675,In_74);
and U2221 (N_2221,In_213,In_929);
or U2222 (N_2222,In_607,In_782);
nand U2223 (N_2223,In_602,In_984);
or U2224 (N_2224,In_345,In_488);
and U2225 (N_2225,In_978,In_342);
and U2226 (N_2226,In_998,In_642);
or U2227 (N_2227,In_889,In_615);
or U2228 (N_2228,In_940,In_858);
nand U2229 (N_2229,In_254,In_733);
or U2230 (N_2230,In_477,In_805);
nand U2231 (N_2231,In_191,In_722);
nor U2232 (N_2232,In_812,In_575);
and U2233 (N_2233,In_553,In_655);
or U2234 (N_2234,In_640,In_653);
or U2235 (N_2235,In_169,In_507);
or U2236 (N_2236,In_316,In_799);
or U2237 (N_2237,In_176,In_687);
nand U2238 (N_2238,In_132,In_604);
nor U2239 (N_2239,In_99,In_453);
nor U2240 (N_2240,In_465,In_969);
and U2241 (N_2241,In_476,In_89);
and U2242 (N_2242,In_227,In_278);
and U2243 (N_2243,In_33,In_843);
or U2244 (N_2244,In_229,In_689);
or U2245 (N_2245,In_684,In_828);
nor U2246 (N_2246,In_549,In_92);
and U2247 (N_2247,In_653,In_31);
and U2248 (N_2248,In_107,In_846);
and U2249 (N_2249,In_12,In_810);
or U2250 (N_2250,In_829,In_377);
nand U2251 (N_2251,In_695,In_201);
nand U2252 (N_2252,In_732,In_220);
nor U2253 (N_2253,In_439,In_761);
nor U2254 (N_2254,In_834,In_343);
and U2255 (N_2255,In_334,In_539);
nand U2256 (N_2256,In_605,In_777);
and U2257 (N_2257,In_557,In_192);
xor U2258 (N_2258,In_851,In_973);
nand U2259 (N_2259,In_271,In_993);
or U2260 (N_2260,In_258,In_748);
nor U2261 (N_2261,In_732,In_122);
and U2262 (N_2262,In_324,In_637);
nand U2263 (N_2263,In_307,In_29);
or U2264 (N_2264,In_871,In_467);
nor U2265 (N_2265,In_646,In_565);
or U2266 (N_2266,In_184,In_175);
or U2267 (N_2267,In_991,In_511);
nand U2268 (N_2268,In_118,In_865);
or U2269 (N_2269,In_695,In_259);
and U2270 (N_2270,In_930,In_390);
nand U2271 (N_2271,In_128,In_300);
nor U2272 (N_2272,In_926,In_393);
nand U2273 (N_2273,In_803,In_283);
and U2274 (N_2274,In_843,In_811);
nand U2275 (N_2275,In_322,In_885);
or U2276 (N_2276,In_351,In_386);
nor U2277 (N_2277,In_518,In_813);
and U2278 (N_2278,In_367,In_975);
or U2279 (N_2279,In_281,In_772);
nor U2280 (N_2280,In_309,In_601);
nor U2281 (N_2281,In_764,In_80);
nand U2282 (N_2282,In_929,In_481);
or U2283 (N_2283,In_443,In_634);
and U2284 (N_2284,In_62,In_641);
or U2285 (N_2285,In_105,In_457);
and U2286 (N_2286,In_785,In_737);
nor U2287 (N_2287,In_418,In_130);
nand U2288 (N_2288,In_970,In_872);
nor U2289 (N_2289,In_174,In_268);
nor U2290 (N_2290,In_98,In_112);
and U2291 (N_2291,In_356,In_832);
or U2292 (N_2292,In_438,In_562);
and U2293 (N_2293,In_939,In_748);
nor U2294 (N_2294,In_352,In_505);
and U2295 (N_2295,In_580,In_861);
nor U2296 (N_2296,In_187,In_966);
nor U2297 (N_2297,In_696,In_201);
nand U2298 (N_2298,In_906,In_421);
nand U2299 (N_2299,In_594,In_838);
or U2300 (N_2300,In_757,In_652);
nor U2301 (N_2301,In_208,In_399);
and U2302 (N_2302,In_498,In_614);
nand U2303 (N_2303,In_337,In_658);
nor U2304 (N_2304,In_563,In_950);
or U2305 (N_2305,In_37,In_748);
and U2306 (N_2306,In_103,In_854);
or U2307 (N_2307,In_163,In_485);
or U2308 (N_2308,In_763,In_954);
nand U2309 (N_2309,In_459,In_400);
nand U2310 (N_2310,In_26,In_522);
and U2311 (N_2311,In_686,In_54);
or U2312 (N_2312,In_913,In_884);
nand U2313 (N_2313,In_84,In_997);
nor U2314 (N_2314,In_676,In_594);
and U2315 (N_2315,In_576,In_722);
or U2316 (N_2316,In_159,In_262);
or U2317 (N_2317,In_523,In_602);
nor U2318 (N_2318,In_328,In_140);
nor U2319 (N_2319,In_830,In_675);
and U2320 (N_2320,In_609,In_835);
and U2321 (N_2321,In_496,In_852);
or U2322 (N_2322,In_609,In_671);
or U2323 (N_2323,In_116,In_124);
nand U2324 (N_2324,In_633,In_755);
or U2325 (N_2325,In_172,In_329);
nor U2326 (N_2326,In_145,In_480);
or U2327 (N_2327,In_105,In_284);
nand U2328 (N_2328,In_375,In_876);
and U2329 (N_2329,In_315,In_205);
or U2330 (N_2330,In_203,In_556);
or U2331 (N_2331,In_790,In_78);
and U2332 (N_2332,In_706,In_558);
nor U2333 (N_2333,In_275,In_493);
nand U2334 (N_2334,In_319,In_887);
and U2335 (N_2335,In_797,In_777);
nand U2336 (N_2336,In_143,In_185);
nor U2337 (N_2337,In_679,In_428);
nor U2338 (N_2338,In_544,In_905);
nor U2339 (N_2339,In_961,In_486);
nand U2340 (N_2340,In_431,In_383);
and U2341 (N_2341,In_264,In_91);
or U2342 (N_2342,In_190,In_746);
or U2343 (N_2343,In_641,In_989);
or U2344 (N_2344,In_966,In_8);
nand U2345 (N_2345,In_771,In_102);
and U2346 (N_2346,In_237,In_604);
or U2347 (N_2347,In_517,In_345);
nand U2348 (N_2348,In_294,In_423);
nor U2349 (N_2349,In_431,In_615);
and U2350 (N_2350,In_202,In_616);
nor U2351 (N_2351,In_168,In_253);
and U2352 (N_2352,In_921,In_595);
or U2353 (N_2353,In_347,In_184);
nand U2354 (N_2354,In_620,In_898);
nand U2355 (N_2355,In_968,In_916);
nand U2356 (N_2356,In_464,In_306);
nor U2357 (N_2357,In_212,In_846);
nor U2358 (N_2358,In_516,In_706);
or U2359 (N_2359,In_518,In_257);
xnor U2360 (N_2360,In_748,In_357);
nor U2361 (N_2361,In_368,In_127);
or U2362 (N_2362,In_142,In_941);
nor U2363 (N_2363,In_906,In_368);
and U2364 (N_2364,In_505,In_254);
and U2365 (N_2365,In_431,In_15);
nor U2366 (N_2366,In_991,In_919);
or U2367 (N_2367,In_99,In_692);
nand U2368 (N_2368,In_489,In_581);
and U2369 (N_2369,In_133,In_85);
nor U2370 (N_2370,In_703,In_563);
nor U2371 (N_2371,In_682,In_376);
and U2372 (N_2372,In_492,In_851);
nor U2373 (N_2373,In_715,In_582);
nand U2374 (N_2374,In_472,In_339);
nand U2375 (N_2375,In_153,In_899);
nand U2376 (N_2376,In_296,In_689);
or U2377 (N_2377,In_734,In_840);
nor U2378 (N_2378,In_45,In_839);
and U2379 (N_2379,In_120,In_791);
or U2380 (N_2380,In_531,In_537);
or U2381 (N_2381,In_6,In_641);
nor U2382 (N_2382,In_683,In_456);
nor U2383 (N_2383,In_277,In_733);
nand U2384 (N_2384,In_275,In_923);
nand U2385 (N_2385,In_965,In_990);
nand U2386 (N_2386,In_176,In_646);
xnor U2387 (N_2387,In_240,In_449);
or U2388 (N_2388,In_32,In_34);
or U2389 (N_2389,In_16,In_479);
and U2390 (N_2390,In_506,In_881);
and U2391 (N_2391,In_165,In_243);
or U2392 (N_2392,In_854,In_670);
nand U2393 (N_2393,In_120,In_420);
nor U2394 (N_2394,In_235,In_814);
and U2395 (N_2395,In_158,In_205);
nand U2396 (N_2396,In_627,In_672);
and U2397 (N_2397,In_989,In_141);
and U2398 (N_2398,In_136,In_44);
nor U2399 (N_2399,In_247,In_124);
or U2400 (N_2400,In_917,In_897);
nor U2401 (N_2401,In_708,In_487);
xor U2402 (N_2402,In_649,In_359);
nand U2403 (N_2403,In_393,In_404);
nor U2404 (N_2404,In_838,In_507);
or U2405 (N_2405,In_662,In_442);
and U2406 (N_2406,In_518,In_459);
nor U2407 (N_2407,In_732,In_430);
nor U2408 (N_2408,In_618,In_355);
nor U2409 (N_2409,In_899,In_347);
and U2410 (N_2410,In_161,In_655);
nand U2411 (N_2411,In_586,In_331);
nand U2412 (N_2412,In_254,In_825);
or U2413 (N_2413,In_891,In_906);
and U2414 (N_2414,In_127,In_724);
nand U2415 (N_2415,In_385,In_821);
nand U2416 (N_2416,In_466,In_564);
nand U2417 (N_2417,In_682,In_182);
and U2418 (N_2418,In_848,In_909);
nand U2419 (N_2419,In_60,In_567);
nor U2420 (N_2420,In_880,In_746);
and U2421 (N_2421,In_932,In_617);
or U2422 (N_2422,In_757,In_450);
nor U2423 (N_2423,In_843,In_614);
nor U2424 (N_2424,In_677,In_130);
nor U2425 (N_2425,In_119,In_980);
nand U2426 (N_2426,In_620,In_755);
and U2427 (N_2427,In_940,In_970);
or U2428 (N_2428,In_366,In_890);
or U2429 (N_2429,In_638,In_608);
nand U2430 (N_2430,In_851,In_227);
or U2431 (N_2431,In_953,In_748);
xnor U2432 (N_2432,In_498,In_407);
nand U2433 (N_2433,In_494,In_132);
or U2434 (N_2434,In_67,In_108);
or U2435 (N_2435,In_208,In_519);
or U2436 (N_2436,In_500,In_886);
nor U2437 (N_2437,In_616,In_347);
and U2438 (N_2438,In_153,In_314);
and U2439 (N_2439,In_482,In_894);
nor U2440 (N_2440,In_778,In_544);
nor U2441 (N_2441,In_537,In_91);
or U2442 (N_2442,In_469,In_866);
nor U2443 (N_2443,In_387,In_79);
nor U2444 (N_2444,In_169,In_796);
or U2445 (N_2445,In_688,In_126);
and U2446 (N_2446,In_445,In_263);
and U2447 (N_2447,In_668,In_34);
and U2448 (N_2448,In_222,In_59);
and U2449 (N_2449,In_686,In_587);
or U2450 (N_2450,In_739,In_687);
nor U2451 (N_2451,In_660,In_987);
and U2452 (N_2452,In_311,In_611);
xnor U2453 (N_2453,In_711,In_365);
nor U2454 (N_2454,In_815,In_569);
and U2455 (N_2455,In_503,In_661);
and U2456 (N_2456,In_562,In_221);
nor U2457 (N_2457,In_78,In_427);
or U2458 (N_2458,In_705,In_568);
or U2459 (N_2459,In_382,In_398);
or U2460 (N_2460,In_539,In_811);
nand U2461 (N_2461,In_8,In_608);
and U2462 (N_2462,In_236,In_756);
and U2463 (N_2463,In_442,In_464);
nor U2464 (N_2464,In_415,In_736);
and U2465 (N_2465,In_860,In_492);
nand U2466 (N_2466,In_406,In_733);
nand U2467 (N_2467,In_804,In_300);
or U2468 (N_2468,In_253,In_421);
and U2469 (N_2469,In_64,In_51);
nor U2470 (N_2470,In_686,In_15);
nor U2471 (N_2471,In_83,In_814);
and U2472 (N_2472,In_780,In_562);
nor U2473 (N_2473,In_997,In_525);
nor U2474 (N_2474,In_573,In_469);
or U2475 (N_2475,In_853,In_826);
and U2476 (N_2476,In_67,In_531);
nor U2477 (N_2477,In_415,In_472);
nand U2478 (N_2478,In_478,In_582);
and U2479 (N_2479,In_863,In_928);
or U2480 (N_2480,In_838,In_221);
nand U2481 (N_2481,In_186,In_923);
nor U2482 (N_2482,In_60,In_942);
nor U2483 (N_2483,In_955,In_952);
nand U2484 (N_2484,In_641,In_520);
nand U2485 (N_2485,In_992,In_85);
and U2486 (N_2486,In_906,In_703);
nor U2487 (N_2487,In_382,In_345);
and U2488 (N_2488,In_645,In_871);
or U2489 (N_2489,In_701,In_148);
and U2490 (N_2490,In_150,In_248);
or U2491 (N_2491,In_232,In_982);
nor U2492 (N_2492,In_785,In_705);
or U2493 (N_2493,In_935,In_472);
and U2494 (N_2494,In_600,In_377);
or U2495 (N_2495,In_842,In_464);
or U2496 (N_2496,In_448,In_138);
or U2497 (N_2497,In_591,In_290);
or U2498 (N_2498,In_584,In_592);
nor U2499 (N_2499,In_66,In_550);
nand U2500 (N_2500,N_519,N_1167);
nand U2501 (N_2501,N_1057,N_2081);
and U2502 (N_2502,N_372,N_655);
or U2503 (N_2503,N_188,N_1697);
and U2504 (N_2504,N_1574,N_217);
and U2505 (N_2505,N_1474,N_2300);
nor U2506 (N_2506,N_1831,N_2324);
and U2507 (N_2507,N_864,N_2062);
nand U2508 (N_2508,N_288,N_2007);
nand U2509 (N_2509,N_133,N_1271);
and U2510 (N_2510,N_1048,N_1412);
nand U2511 (N_2511,N_1949,N_177);
xor U2512 (N_2512,N_76,N_1861);
or U2513 (N_2513,N_1052,N_745);
xnor U2514 (N_2514,N_2432,N_2206);
and U2515 (N_2515,N_1422,N_2499);
or U2516 (N_2516,N_978,N_220);
or U2517 (N_2517,N_977,N_1514);
nor U2518 (N_2518,N_1985,N_621);
nand U2519 (N_2519,N_1022,N_878);
nor U2520 (N_2520,N_1282,N_2258);
nor U2521 (N_2521,N_326,N_1088);
nor U2522 (N_2522,N_1044,N_1812);
and U2523 (N_2523,N_501,N_141);
nand U2524 (N_2524,N_1187,N_411);
nand U2525 (N_2525,N_1951,N_713);
nor U2526 (N_2526,N_2080,N_75);
nand U2527 (N_2527,N_72,N_2183);
or U2528 (N_2528,N_1847,N_272);
and U2529 (N_2529,N_2078,N_2240);
nand U2530 (N_2530,N_685,N_189);
nor U2531 (N_2531,N_2110,N_1999);
nand U2532 (N_2532,N_1318,N_763);
nand U2533 (N_2533,N_144,N_602);
or U2534 (N_2534,N_2233,N_608);
and U2535 (N_2535,N_812,N_122);
or U2536 (N_2536,N_1256,N_1881);
and U2537 (N_2537,N_2120,N_1533);
and U2538 (N_2538,N_164,N_610);
nor U2539 (N_2539,N_476,N_1767);
or U2540 (N_2540,N_1281,N_793);
nand U2541 (N_2541,N_159,N_2459);
or U2542 (N_2542,N_820,N_2125);
and U2543 (N_2543,N_1801,N_277);
and U2544 (N_2544,N_172,N_2409);
nor U2545 (N_2545,N_2219,N_1552);
nor U2546 (N_2546,N_2428,N_1210);
and U2547 (N_2547,N_1077,N_2225);
and U2548 (N_2548,N_96,N_2061);
nor U2549 (N_2549,N_284,N_798);
and U2550 (N_2550,N_1150,N_429);
nor U2551 (N_2551,N_2412,N_104);
and U2552 (N_2552,N_2145,N_193);
nor U2553 (N_2553,N_437,N_2151);
nand U2554 (N_2554,N_673,N_1229);
nand U2555 (N_2555,N_841,N_2108);
nand U2556 (N_2556,N_1042,N_2245);
and U2557 (N_2557,N_1089,N_2241);
nand U2558 (N_2558,N_2445,N_1395);
nor U2559 (N_2559,N_1065,N_253);
and U2560 (N_2560,N_2435,N_1369);
nor U2561 (N_2561,N_2380,N_628);
and U2562 (N_2562,N_1434,N_119);
nand U2563 (N_2563,N_1862,N_261);
nor U2564 (N_2564,N_2138,N_1916);
or U2565 (N_2565,N_1452,N_860);
nand U2566 (N_2566,N_174,N_2292);
nor U2567 (N_2567,N_1062,N_1279);
and U2568 (N_2568,N_212,N_503);
nor U2569 (N_2569,N_1682,N_2457);
and U2570 (N_2570,N_1523,N_1188);
nand U2571 (N_2571,N_2228,N_347);
and U2572 (N_2572,N_1711,N_1437);
and U2573 (N_2573,N_1982,N_1358);
nand U2574 (N_2574,N_699,N_1472);
and U2575 (N_2575,N_1567,N_138);
and U2576 (N_2576,N_1858,N_246);
or U2577 (N_2577,N_1185,N_1888);
nor U2578 (N_2578,N_1764,N_83);
or U2579 (N_2579,N_556,N_89);
or U2580 (N_2580,N_1816,N_959);
and U2581 (N_2581,N_35,N_891);
or U2582 (N_2582,N_611,N_1687);
and U2583 (N_2583,N_361,N_1011);
nor U2584 (N_2584,N_786,N_4);
and U2585 (N_2585,N_109,N_774);
nor U2586 (N_2586,N_822,N_642);
or U2587 (N_2587,N_759,N_2033);
and U2588 (N_2588,N_373,N_923);
nand U2589 (N_2589,N_1417,N_792);
and U2590 (N_2590,N_2496,N_2488);
nand U2591 (N_2591,N_2319,N_607);
nor U2592 (N_2592,N_1327,N_987);
and U2593 (N_2593,N_805,N_1186);
and U2594 (N_2594,N_2484,N_1810);
nor U2595 (N_2595,N_2360,N_2337);
nor U2596 (N_2596,N_1918,N_1835);
and U2597 (N_2597,N_91,N_1938);
nand U2598 (N_2598,N_1575,N_2472);
nor U2599 (N_2599,N_2397,N_784);
nand U2600 (N_2600,N_1499,N_1691);
nor U2601 (N_2601,N_557,N_1069);
and U2602 (N_2602,N_2103,N_2246);
and U2603 (N_2603,N_604,N_1490);
nand U2604 (N_2604,N_1481,N_1934);
or U2605 (N_2605,N_2466,N_1197);
and U2606 (N_2606,N_1205,N_892);
and U2607 (N_2607,N_531,N_1286);
nor U2608 (N_2608,N_574,N_2167);
nand U2609 (N_2609,N_1194,N_909);
and U2610 (N_2610,N_1366,N_1730);
or U2611 (N_2611,N_524,N_1432);
nor U2612 (N_2612,N_409,N_2439);
and U2613 (N_2613,N_167,N_768);
nor U2614 (N_2614,N_1675,N_1598);
nand U2615 (N_2615,N_134,N_550);
or U2616 (N_2616,N_788,N_251);
nor U2617 (N_2617,N_1624,N_2127);
nor U2618 (N_2618,N_815,N_2329);
nand U2619 (N_2619,N_1445,N_2053);
or U2620 (N_2620,N_1275,N_1664);
and U2621 (N_2621,N_386,N_579);
nor U2622 (N_2622,N_150,N_823);
and U2623 (N_2623,N_2383,N_2220);
and U2624 (N_2624,N_1750,N_1321);
nor U2625 (N_2625,N_1943,N_2441);
nor U2626 (N_2626,N_2042,N_1662);
and U2627 (N_2627,N_1181,N_1280);
and U2628 (N_2628,N_181,N_306);
nand U2629 (N_2629,N_1776,N_529);
nand U2630 (N_2630,N_1377,N_2199);
and U2631 (N_2631,N_2214,N_1371);
or U2632 (N_2632,N_2447,N_755);
nor U2633 (N_2633,N_472,N_1253);
nor U2634 (N_2634,N_593,N_200);
nand U2635 (N_2635,N_1726,N_435);
and U2636 (N_2636,N_1343,N_1457);
nand U2637 (N_2637,N_1571,N_1727);
or U2638 (N_2638,N_225,N_568);
nor U2639 (N_2639,N_450,N_1517);
nor U2640 (N_2640,N_1720,N_975);
and U2641 (N_2641,N_1549,N_1928);
nor U2642 (N_2642,N_1794,N_1689);
nor U2643 (N_2643,N_1311,N_2079);
nand U2644 (N_2644,N_56,N_2271);
or U2645 (N_2645,N_3,N_1171);
or U2646 (N_2646,N_1957,N_1442);
nand U2647 (N_2647,N_203,N_634);
nand U2648 (N_2648,N_1799,N_7);
and U2649 (N_2649,N_1820,N_1696);
nand U2650 (N_2650,N_1360,N_2209);
nor U2651 (N_2651,N_1977,N_118);
nand U2652 (N_2652,N_2384,N_88);
nand U2653 (N_2653,N_1262,N_1768);
nand U2654 (N_2654,N_1606,N_77);
or U2655 (N_2655,N_453,N_2342);
nor U2656 (N_2656,N_2216,N_599);
nor U2657 (N_2657,N_474,N_2421);
or U2658 (N_2658,N_744,N_1905);
and U2659 (N_2659,N_2226,N_1561);
and U2660 (N_2660,N_273,N_2281);
and U2661 (N_2661,N_2201,N_1272);
nand U2662 (N_2662,N_2026,N_1220);
nor U2663 (N_2663,N_1558,N_1805);
nand U2664 (N_2664,N_237,N_2440);
nor U2665 (N_2665,N_406,N_2469);
nand U2666 (N_2666,N_365,N_551);
nor U2667 (N_2667,N_697,N_2481);
or U2668 (N_2668,N_155,N_407);
nor U2669 (N_2669,N_795,N_2067);
or U2670 (N_2670,N_120,N_1607);
nand U2671 (N_2671,N_1100,N_709);
or U2672 (N_2672,N_693,N_1324);
or U2673 (N_2673,N_2390,N_395);
or U2674 (N_2674,N_374,N_1121);
or U2675 (N_2675,N_2109,N_581);
nand U2676 (N_2676,N_323,N_1619);
or U2677 (N_2677,N_2172,N_528);
nor U2678 (N_2678,N_1459,N_1397);
nand U2679 (N_2679,N_543,N_2287);
and U2680 (N_2680,N_2003,N_378);
and U2681 (N_2681,N_2204,N_868);
or U2682 (N_2682,N_298,N_662);
nor U2683 (N_2683,N_496,N_244);
or U2684 (N_2684,N_2465,N_2394);
nand U2685 (N_2685,N_1030,N_2088);
and U2686 (N_2686,N_1355,N_2133);
nor U2687 (N_2687,N_2313,N_269);
nand U2688 (N_2688,N_511,N_684);
nand U2689 (N_2689,N_2143,N_708);
nor U2690 (N_2690,N_1202,N_2419);
or U2691 (N_2691,N_92,N_2197);
nor U2692 (N_2692,N_1008,N_1853);
and U2693 (N_2693,N_1512,N_2302);
nand U2694 (N_2694,N_10,N_1793);
and U2695 (N_2695,N_1015,N_14);
or U2696 (N_2696,N_151,N_1078);
and U2697 (N_2697,N_451,N_2413);
or U2698 (N_2698,N_2414,N_43);
or U2699 (N_2699,N_1569,N_771);
and U2700 (N_2700,N_31,N_444);
nand U2701 (N_2701,N_530,N_1317);
or U2702 (N_2702,N_1570,N_2372);
and U2703 (N_2703,N_1666,N_2091);
nor U2704 (N_2704,N_111,N_1560);
or U2705 (N_2705,N_1214,N_1972);
nor U2706 (N_2706,N_441,N_45);
or U2707 (N_2707,N_2369,N_2063);
nand U2708 (N_2708,N_821,N_452);
and U2709 (N_2709,N_1811,N_2203);
nor U2710 (N_2710,N_606,N_854);
nor U2711 (N_2711,N_401,N_1705);
and U2712 (N_2712,N_1582,N_250);
nor U2713 (N_2713,N_2244,N_1364);
or U2714 (N_2714,N_887,N_157);
or U2715 (N_2715,N_1637,N_1813);
and U2716 (N_2716,N_2021,N_1900);
or U2717 (N_2717,N_668,N_1163);
and U2718 (N_2718,N_281,N_304);
or U2719 (N_2719,N_2014,N_1832);
or U2720 (N_2720,N_758,N_2236);
or U2721 (N_2721,N_2396,N_2051);
nor U2722 (N_2722,N_463,N_485);
or U2723 (N_2723,N_675,N_1906);
nor U2724 (N_2724,N_772,N_894);
or U2725 (N_2725,N_187,N_2297);
nand U2726 (N_2726,N_690,N_303);
and U2727 (N_2727,N_2353,N_523);
or U2728 (N_2728,N_641,N_1838);
nor U2729 (N_2729,N_191,N_1268);
or U2730 (N_2730,N_2198,N_1204);
nor U2731 (N_2731,N_799,N_1314);
nand U2732 (N_2732,N_1012,N_1329);
and U2733 (N_2733,N_687,N_572);
and U2734 (N_2734,N_2309,N_2087);
nand U2735 (N_2735,N_827,N_2314);
or U2736 (N_2736,N_29,N_436);
or U2737 (N_2737,N_17,N_1230);
nand U2738 (N_2738,N_1394,N_1710);
nor U2739 (N_2739,N_845,N_1718);
nand U2740 (N_2740,N_1631,N_2237);
or U2741 (N_2741,N_1864,N_414);
nor U2742 (N_2742,N_1755,N_2057);
and U2743 (N_2743,N_1867,N_1049);
and U2744 (N_2744,N_1962,N_293);
nor U2745 (N_2745,N_766,N_55);
or U2746 (N_2746,N_2264,N_2029);
nand U2747 (N_2747,N_1592,N_1741);
or U2748 (N_2748,N_38,N_499);
or U2749 (N_2749,N_695,N_352);
and U2750 (N_2750,N_1632,N_2490);
nand U2751 (N_2751,N_804,N_595);
nor U2752 (N_2752,N_2211,N_1372);
or U2753 (N_2753,N_291,N_2102);
or U2754 (N_2754,N_830,N_129);
nand U2755 (N_2755,N_743,N_2196);
or U2756 (N_2756,N_224,N_388);
nand U2757 (N_2757,N_481,N_2162);
nand U2758 (N_2758,N_908,N_1251);
or U2759 (N_2759,N_169,N_649);
nand U2760 (N_2760,N_2142,N_176);
and U2761 (N_2761,N_1541,N_2429);
or U2762 (N_2762,N_922,N_1611);
nor U2763 (N_2763,N_1291,N_1760);
nor U2764 (N_2764,N_737,N_175);
or U2765 (N_2765,N_492,N_2134);
and U2766 (N_2766,N_863,N_1161);
nand U2767 (N_2767,N_522,N_748);
nand U2768 (N_2768,N_1368,N_665);
nor U2769 (N_2769,N_2186,N_1094);
and U2770 (N_2770,N_506,N_1981);
or U2771 (N_2771,N_1531,N_121);
nor U2772 (N_2772,N_1990,N_2482);
nor U2773 (N_2773,N_1245,N_565);
nand U2774 (N_2774,N_1200,N_166);
or U2775 (N_2775,N_1717,N_1148);
nand U2776 (N_2776,N_1869,N_888);
or U2777 (N_2777,N_479,N_1158);
nor U2778 (N_2778,N_1460,N_210);
or U2779 (N_2779,N_545,N_1419);
nand U2780 (N_2780,N_1555,N_920);
and U2781 (N_2781,N_1028,N_1276);
or U2782 (N_2782,N_1852,N_2437);
nor U2783 (N_2783,N_202,N_2178);
or U2784 (N_2784,N_2164,N_1115);
and U2785 (N_2785,N_445,N_1586);
nand U2786 (N_2786,N_1660,N_1375);
and U2787 (N_2787,N_2480,N_893);
nand U2788 (N_2788,N_1380,N_2345);
or U2789 (N_2789,N_1609,N_1403);
nand U2790 (N_2790,N_1353,N_1529);
or U2791 (N_2791,N_2075,N_185);
nor U2792 (N_2792,N_2296,N_1123);
or U2793 (N_2793,N_2181,N_1783);
nor U2794 (N_2794,N_2463,N_1312);
xnor U2795 (N_2795,N_1930,N_1034);
or U2796 (N_2796,N_1244,N_482);
xnor U2797 (N_2797,N_1883,N_578);
or U2798 (N_2798,N_103,N_8);
and U2799 (N_2799,N_1504,N_1667);
nand U2800 (N_2800,N_1299,N_609);
nor U2801 (N_2801,N_389,N_2251);
or U2802 (N_2802,N_493,N_1952);
nor U2803 (N_2803,N_1897,N_1699);
and U2804 (N_2804,N_9,N_900);
and U2805 (N_2805,N_1551,N_1734);
nor U2806 (N_2806,N_2011,N_65);
or U2807 (N_2807,N_1149,N_1643);
nor U2808 (N_2808,N_2016,N_747);
nand U2809 (N_2809,N_1747,N_1237);
or U2810 (N_2810,N_1336,N_1104);
or U2811 (N_2811,N_1998,N_1240);
or U2812 (N_2812,N_2467,N_976);
nand U2813 (N_2813,N_953,N_2450);
and U2814 (N_2814,N_1941,N_2462);
nand U2815 (N_2815,N_1665,N_471);
nand U2816 (N_2816,N_1651,N_1345);
nor U2817 (N_2817,N_2210,N_1216);
or U2818 (N_2818,N_727,N_1578);
or U2819 (N_2819,N_1503,N_2250);
nor U2820 (N_2820,N_1703,N_2315);
or U2821 (N_2821,N_294,N_1648);
nand U2822 (N_2822,N_915,N_2037);
and U2823 (N_2823,N_39,N_1192);
and U2824 (N_2824,N_190,N_186);
nor U2825 (N_2825,N_1076,N_521);
nor U2826 (N_2826,N_171,N_1382);
nand U2827 (N_2827,N_2034,N_2008);
and U2828 (N_2828,N_126,N_2338);
and U2829 (N_2829,N_643,N_686);
nand U2830 (N_2830,N_1615,N_1290);
and U2831 (N_2831,N_287,N_2351);
nor U2832 (N_2832,N_1047,N_364);
nor U2833 (N_2833,N_584,N_2060);
nand U2834 (N_2834,N_1772,N_1802);
or U2835 (N_2835,N_320,N_1505);
and U2836 (N_2836,N_1842,N_1146);
and U2837 (N_2837,N_622,N_2365);
or U2838 (N_2838,N_615,N_2059);
nor U2839 (N_2839,N_391,N_2239);
nand U2840 (N_2840,N_2420,N_769);
or U2841 (N_2841,N_110,N_2243);
nor U2842 (N_2842,N_1762,N_325);
nor U2843 (N_2843,N_1885,N_623);
and U2844 (N_2844,N_552,N_535);
nor U2845 (N_2845,N_997,N_787);
nor U2846 (N_2846,N_1628,N_1289);
or U2847 (N_2847,N_837,N_15);
nor U2848 (N_2848,N_1545,N_934);
or U2849 (N_2849,N_930,N_1182);
nor U2850 (N_2850,N_1828,N_1009);
and U2851 (N_2851,N_1173,N_2492);
or U2852 (N_2852,N_1819,N_2378);
nor U2853 (N_2853,N_32,N_100);
and U2854 (N_2854,N_1633,N_1581);
or U2855 (N_2855,N_800,N_1453);
xnor U2856 (N_2856,N_2076,N_1780);
or U2857 (N_2857,N_42,N_1613);
nor U2858 (N_2858,N_1258,N_2320);
nand U2859 (N_2859,N_1892,N_938);
and U2860 (N_2860,N_717,N_1630);
or U2861 (N_2861,N_1242,N_2389);
and U2862 (N_2862,N_258,N_1273);
or U2863 (N_2863,N_33,N_999);
or U2864 (N_2864,N_566,N_1131);
nor U2865 (N_2865,N_1482,N_1993);
and U2866 (N_2866,N_1647,N_1099);
nor U2867 (N_2867,N_1084,N_505);
and U2868 (N_2868,N_1213,N_1654);
nor U2869 (N_2869,N_2165,N_580);
and U2870 (N_2870,N_2161,N_906);
or U2871 (N_2871,N_2153,N_2128);
and U2872 (N_2872,N_1976,N_2404);
nor U2873 (N_2873,N_1702,N_263);
nor U2874 (N_2874,N_954,N_97);
or U2875 (N_2875,N_1223,N_718);
and U2876 (N_2876,N_271,N_931);
xnor U2877 (N_2877,N_2208,N_152);
nor U2878 (N_2878,N_95,N_1501);
or U2879 (N_2879,N_1784,N_1528);
or U2880 (N_2880,N_1421,N_1925);
nor U2881 (N_2881,N_1797,N_1940);
and U2882 (N_2882,N_382,N_1912);
nor U2883 (N_2883,N_765,N_427);
nor U2884 (N_2884,N_1536,N_1880);
nand U2885 (N_2885,N_696,N_1969);
nor U2886 (N_2886,N_853,N_880);
nor U2887 (N_2887,N_2283,N_268);
nor U2888 (N_2888,N_1754,N_2015);
nand U2889 (N_2889,N_467,N_1248);
and U2890 (N_2890,N_738,N_858);
or U2891 (N_2891,N_1645,N_248);
nor U2892 (N_2892,N_1098,N_2438);
xnor U2893 (N_2893,N_852,N_1920);
nand U2894 (N_2894,N_1095,N_886);
or U2895 (N_2895,N_694,N_455);
or U2896 (N_2896,N_430,N_1338);
or U2897 (N_2897,N_1845,N_652);
or U2898 (N_2898,N_679,N_1913);
and U2899 (N_2899,N_948,N_539);
or U2900 (N_2900,N_148,N_846);
and U2901 (N_2901,N_1707,N_1789);
nand U2902 (N_2902,N_1626,N_2285);
or U2903 (N_2903,N_733,N_1807);
nor U2904 (N_2904,N_2327,N_791);
nor U2905 (N_2905,N_921,N_2402);
nand U2906 (N_2906,N_195,N_731);
nand U2907 (N_2907,N_542,N_2072);
nor U2908 (N_2908,N_883,N_153);
or U2909 (N_2909,N_416,N_242);
nand U2910 (N_2910,N_1729,N_1850);
and U2911 (N_2911,N_1328,N_881);
nor U2912 (N_2912,N_721,N_631);
nand U2913 (N_2913,N_2265,N_1629);
or U2914 (N_2914,N_266,N_1320);
or U2915 (N_2915,N_344,N_495);
and U2916 (N_2916,N_6,N_2443);
nor U2917 (N_2917,N_1339,N_1255);
nor U2918 (N_2918,N_2111,N_207);
nor U2919 (N_2919,N_1310,N_773);
nand U2920 (N_2920,N_968,N_2366);
nor U2921 (N_2921,N_1463,N_803);
nand U2922 (N_2922,N_726,N_1054);
and U2923 (N_2923,N_1386,N_1958);
nand U2924 (N_2924,N_71,N_36);
nor U2925 (N_2925,N_1614,N_2318);
and U2926 (N_2926,N_2024,N_671);
nor U2927 (N_2927,N_2321,N_1224);
nor U2928 (N_2928,N_1695,N_2160);
or U2929 (N_2929,N_1500,N_617);
nand U2930 (N_2930,N_1201,N_939);
and U2931 (N_2931,N_1752,N_1330);
and U2932 (N_2932,N_192,N_2215);
and U2933 (N_2933,N_1354,N_2227);
nand U2934 (N_2934,N_371,N_1715);
and U2935 (N_2935,N_2023,N_422);
and U2936 (N_2936,N_739,N_1863);
nor U2937 (N_2937,N_567,N_1899);
and U2938 (N_2938,N_1112,N_392);
and U2939 (N_2939,N_1684,N_562);
nor U2940 (N_2940,N_127,N_2129);
nor U2941 (N_2941,N_1506,N_627);
nor U2942 (N_2942,N_1122,N_783);
and U2943 (N_2943,N_1184,N_257);
or U2944 (N_2944,N_1454,N_442);
nor U2945 (N_2945,N_1239,N_285);
or U2946 (N_2946,N_723,N_2303);
nor U2947 (N_2947,N_829,N_239);
nand U2948 (N_2948,N_2494,N_69);
and U2949 (N_2949,N_2232,N_1458);
nor U2950 (N_2950,N_1388,N_1027);
or U2951 (N_2951,N_494,N_1841);
and U2952 (N_2952,N_1189,N_1059);
or U2953 (N_2953,N_1092,N_945);
nor U2954 (N_2954,N_2046,N_674);
and U2955 (N_2955,N_2044,N_514);
nor U2956 (N_2956,N_1968,N_1128);
nor U2957 (N_2957,N_2368,N_197);
or U2958 (N_2958,N_1870,N_969);
nand U2959 (N_2959,N_1413,N_1250);
nor U2960 (N_2960,N_1191,N_956);
or U2961 (N_2961,N_2294,N_1960);
or U2962 (N_2962,N_1020,N_972);
or U2963 (N_2963,N_1036,N_1479);
or U2964 (N_2964,N_1946,N_1562);
or U2965 (N_2965,N_468,N_1243);
nand U2966 (N_2966,N_1680,N_992);
or U2967 (N_2967,N_2100,N_66);
or U2968 (N_2968,N_1898,N_2487);
and U2969 (N_2969,N_1293,N_1018);
and U2970 (N_2970,N_1130,N_2180);
or U2971 (N_2971,N_1671,N_1176);
or U2972 (N_2972,N_311,N_213);
nand U2973 (N_2973,N_926,N_321);
nand U2974 (N_2974,N_569,N_227);
nand U2975 (N_2975,N_1406,N_912);
or U2976 (N_2976,N_102,N_443);
and U2977 (N_2977,N_2089,N_736);
or U2978 (N_2978,N_2114,N_1775);
nand U2979 (N_2979,N_1014,N_1378);
nor U2980 (N_2980,N_1238,N_1051);
or U2981 (N_2981,N_1809,N_657);
and U2982 (N_2982,N_2334,N_123);
nand U2983 (N_2983,N_1137,N_813);
and U2984 (N_2984,N_677,N_1919);
or U2985 (N_2985,N_1509,N_282);
or U2986 (N_2986,N_2306,N_334);
and U2987 (N_2987,N_2273,N_252);
nand U2988 (N_2988,N_1519,N_586);
nor U2989 (N_2989,N_1407,N_2074);
nor U2990 (N_2990,N_704,N_1491);
nor U2991 (N_2991,N_910,N_262);
and U2992 (N_2992,N_826,N_16);
or U2993 (N_2993,N_2234,N_917);
or U2994 (N_2994,N_2263,N_354);
and U2995 (N_2995,N_1933,N_1485);
and U2996 (N_2996,N_113,N_2478);
or U2997 (N_2997,N_681,N_1332);
nor U2998 (N_2998,N_818,N_2139);
nor U2999 (N_2999,N_1359,N_902);
nand U3000 (N_3000,N_797,N_1379);
nand U3001 (N_3001,N_1341,N_1672);
nand U3002 (N_3002,N_855,N_808);
nand U3003 (N_3003,N_458,N_1441);
or U3004 (N_3004,N_238,N_626);
and U3005 (N_3005,N_1759,N_2054);
nor U3006 (N_3006,N_1296,N_1564);
or U3007 (N_3007,N_1929,N_1818);
or U3008 (N_3008,N_336,N_233);
nand U3009 (N_3009,N_1733,N_828);
nand U3010 (N_3010,N_1742,N_204);
nand U3011 (N_3011,N_1932,N_486);
and U3012 (N_3012,N_1132,N_859);
and U3013 (N_3013,N_1524,N_201);
nor U3014 (N_3014,N_232,N_1124);
or U3015 (N_3015,N_847,N_206);
nor U3016 (N_3016,N_1644,N_1585);
nand U3017 (N_3017,N_2101,N_2433);
nor U3018 (N_3018,N_1636,N_842);
or U3019 (N_3019,N_1956,N_2290);
nand U3020 (N_3020,N_296,N_1874);
nor U3021 (N_3021,N_1806,N_460);
or U3022 (N_3022,N_1208,N_1356);
and U3023 (N_3023,N_1693,N_1537);
nand U3024 (N_3024,N_1959,N_1978);
nor U3025 (N_3025,N_369,N_2391);
and U3026 (N_3026,N_1868,N_2461);
or U3027 (N_3027,N_1170,N_275);
and U3028 (N_3028,N_691,N_1233);
or U3029 (N_3029,N_80,N_754);
nor U3030 (N_3030,N_879,N_1154);
and U3031 (N_3031,N_2479,N_12);
nor U3032 (N_3032,N_1964,N_456);
or U3033 (N_3033,N_597,N_2122);
or U3034 (N_3034,N_2043,N_1489);
nand U3035 (N_3035,N_1840,N_2493);
or U3036 (N_3036,N_1235,N_1438);
and U3037 (N_3037,N_2491,N_1971);
nor U3038 (N_3038,N_833,N_682);
and U3039 (N_3039,N_1436,N_1532);
and U3040 (N_3040,N_79,N_1766);
nand U3041 (N_3041,N_240,N_2191);
nand U3042 (N_3042,N_260,N_131);
nor U3043 (N_3043,N_431,N_762);
nor U3044 (N_3044,N_1325,N_142);
nand U3045 (N_3045,N_417,N_1821);
nor U3046 (N_3046,N_488,N_1005);
nor U3047 (N_3047,N_2086,N_2036);
and U3048 (N_3048,N_2065,N_866);
and U3049 (N_3049,N_2261,N_2468);
and U3050 (N_3050,N_1851,N_1010);
nand U3051 (N_3051,N_2410,N_756);
nor U3052 (N_3052,N_381,N_2274);
nor U3053 (N_3053,N_2364,N_1787);
nand U3054 (N_3054,N_1085,N_2221);
nor U3055 (N_3055,N_2477,N_2040);
or U3056 (N_3056,N_703,N_1348);
nor U3057 (N_3057,N_1056,N_835);
nand U3058 (N_3058,N_1713,N_2212);
and U3059 (N_3059,N_48,N_47);
and U3060 (N_3060,N_577,N_1021);
or U3061 (N_3061,N_1579,N_989);
nor U3062 (N_3062,N_625,N_979);
and U3063 (N_3063,N_715,N_21);
nand U3064 (N_3064,N_67,N_1963);
nor U3065 (N_3065,N_300,N_1294);
or U3066 (N_3066,N_1013,N_487);
nor U3067 (N_3067,N_1974,N_86);
nand U3068 (N_3068,N_2349,N_82);
and U3069 (N_3069,N_2448,N_2486);
or U3070 (N_3070,N_1270,N_1587);
or U3071 (N_3071,N_2411,N_1231);
or U3072 (N_3072,N_53,N_1659);
nand U3073 (N_3073,N_1127,N_780);
nor U3074 (N_3074,N_2350,N_457);
or U3075 (N_3075,N_265,N_614);
nor U3076 (N_3076,N_664,N_1212);
and U3077 (N_3077,N_898,N_432);
nor U3078 (N_3078,N_454,N_440);
nor U3079 (N_3079,N_1304,N_413);
or U3080 (N_3080,N_2085,N_1119);
or U3081 (N_3081,N_1988,N_1183);
nand U3082 (N_3082,N_1595,N_11);
nand U3083 (N_3083,N_1737,N_398);
or U3084 (N_3084,N_2379,N_1053);
and U3085 (N_3085,N_1017,N_973);
nand U3086 (N_3086,N_2371,N_2177);
and U3087 (N_3087,N_1190,N_849);
and U3088 (N_3088,N_1873,N_247);
nand U3089 (N_3089,N_351,N_1249);
nand U3090 (N_3090,N_40,N_146);
and U3091 (N_3091,N_1465,N_1979);
and U3092 (N_3092,N_1168,N_1384);
nand U3093 (N_3093,N_749,N_1423);
nand U3094 (N_3094,N_19,N_1103);
nand U3095 (N_3095,N_2047,N_850);
nor U3096 (N_3096,N_2200,N_955);
nor U3097 (N_3097,N_1749,N_1830);
nor U3098 (N_3098,N_2398,N_970);
or U3099 (N_3099,N_563,N_811);
nand U3100 (N_3100,N_73,N_1824);
or U3101 (N_3101,N_1677,N_1690);
nor U3102 (N_3102,N_2123,N_1265);
or U3103 (N_3103,N_1439,N_477);
and U3104 (N_3104,N_1241,N_896);
nand U3105 (N_3105,N_1498,N_465);
nor U3106 (N_3106,N_1992,N_1091);
and U3107 (N_3107,N_1082,N_865);
nand U3108 (N_3108,N_1886,N_875);
or U3109 (N_3109,N_1527,N_612);
or U3110 (N_3110,N_1178,N_752);
or U3111 (N_3111,N_135,N_1756);
nand U3112 (N_3112,N_362,N_2010);
and U3113 (N_3113,N_1950,N_1884);
xor U3114 (N_3114,N_1073,N_1577);
or U3115 (N_3115,N_809,N_1763);
or U3116 (N_3116,N_439,N_2066);
nand U3117 (N_3117,N_832,N_1315);
nand U3118 (N_3118,N_276,N_2357);
nand U3119 (N_3119,N_2056,N_526);
or U3120 (N_3120,N_1944,N_1510);
and U3121 (N_3121,N_712,N_1518);
or U3122 (N_3122,N_1826,N_1086);
nor U3123 (N_3123,N_2174,N_1922);
nand U3124 (N_3124,N_870,N_2070);
nand U3125 (N_3125,N_659,N_555);
nand U3126 (N_3126,N_1424,N_37);
or U3127 (N_3127,N_957,N_2427);
nor U3128 (N_3128,N_54,N_1470);
or U3129 (N_3129,N_1937,N_1284);
nor U3130 (N_3130,N_947,N_583);
nor U3131 (N_3131,N_249,N_724);
nand U3132 (N_3132,N_1374,N_1144);
nor U3133 (N_3133,N_2431,N_705);
or U3134 (N_3134,N_408,N_461);
nand U3135 (N_3135,N_1234,N_914);
and U3136 (N_3136,N_1849,N_2276);
or U3137 (N_3137,N_2247,N_2301);
nor U3138 (N_3138,N_980,N_1743);
nand U3139 (N_3139,N_2474,N_308);
or U3140 (N_3140,N_1777,N_1945);
nand U3141 (N_3141,N_2092,N_750);
nor U3142 (N_3142,N_981,N_2069);
nand U3143 (N_3143,N_1911,N_2105);
nand U3144 (N_3144,N_582,N_1177);
nor U3145 (N_3145,N_1016,N_116);
nor U3146 (N_3146,N_2038,N_801);
nor U3147 (N_3147,N_630,N_63);
or U3148 (N_3148,N_1456,N_1563);
nor U3149 (N_3149,N_1815,N_497);
nand U3150 (N_3150,N_867,N_270);
and U3151 (N_3151,N_2158,N_2392);
or U3152 (N_3152,N_370,N_1625);
and U3153 (N_3153,N_2146,N_22);
nand U3154 (N_3154,N_1839,N_1125);
and U3155 (N_3155,N_796,N_576);
or U3156 (N_3156,N_564,N_502);
nor U3157 (N_3157,N_357,N_504);
nand U3158 (N_3158,N_1891,N_355);
nand U3159 (N_3159,N_383,N_2403);
nand U3160 (N_3160,N_1493,N_0);
and U3161 (N_3161,N_720,N_1);
nor U3162 (N_3162,N_1393,N_507);
nor U3163 (N_3163,N_834,N_1803);
nor U3164 (N_3164,N_68,N_1591);
or U3165 (N_3165,N_943,N_1000);
or U3166 (N_3166,N_322,N_1425);
and U3167 (N_3167,N_1169,N_729);
nand U3168 (N_3168,N_1526,N_1334);
nor U3169 (N_3169,N_339,N_1954);
and U3170 (N_3170,N_518,N_1566);
and U3171 (N_3171,N_2256,N_1790);
nand U3172 (N_3172,N_2195,N_194);
or U3173 (N_3173,N_464,N_1475);
or U3174 (N_3174,N_2238,N_420);
nor U3175 (N_3175,N_346,N_525);
and U3176 (N_3176,N_2275,N_2018);
nor U3177 (N_3177,N_342,N_2179);
nand U3178 (N_3178,N_517,N_115);
and U3179 (N_3179,N_301,N_2118);
nor U3180 (N_3180,N_1774,N_490);
nor U3181 (N_3181,N_941,N_137);
nand U3182 (N_3182,N_824,N_107);
and U3183 (N_3183,N_1083,N_1274);
nor U3184 (N_3184,N_1308,N_2312);
nand U3185 (N_3185,N_1448,N_639);
nor U3186 (N_3186,N_647,N_1430);
nand U3187 (N_3187,N_1175,N_1254);
nor U3188 (N_3188,N_1404,N_18);
or U3189 (N_3189,N_1079,N_1004);
nand U3190 (N_3190,N_761,N_1264);
and U3191 (N_3191,N_2408,N_605);
and U3192 (N_3192,N_1431,N_1723);
nor U3193 (N_3193,N_2121,N_2205);
and U3194 (N_3194,N_790,N_1657);
nand U3195 (N_3195,N_2407,N_2282);
nand U3196 (N_3196,N_1006,N_428);
nor U3197 (N_3197,N_278,N_469);
and U3198 (N_3198,N_2148,N_1995);
nor U3199 (N_3199,N_1496,N_393);
xor U3200 (N_3200,N_862,N_85);
or U3201 (N_3201,N_1894,N_165);
or U3202 (N_3202,N_1745,N_74);
or U3203 (N_3203,N_1305,N_1319);
nand U3204 (N_3204,N_534,N_590);
and U3205 (N_3205,N_1159,N_1520);
or U3206 (N_3206,N_816,N_1604);
or U3207 (N_3207,N_1283,N_1970);
or U3208 (N_3208,N_2323,N_211);
or U3209 (N_3209,N_289,N_940);
or U3210 (N_3210,N_99,N_2343);
or U3211 (N_3211,N_484,N_1347);
nor U3212 (N_3212,N_1365,N_1097);
and U3213 (N_3213,N_2190,N_1050);
nand U3214 (N_3214,N_1823,N_596);
nor U3215 (N_3215,N_1116,N_2095);
nor U3216 (N_3216,N_1466,N_2299);
nand U3217 (N_3217,N_1138,N_1222);
and U3218 (N_3218,N_139,N_28);
and U3219 (N_3219,N_2173,N_2361);
and U3220 (N_3220,N_2331,N_60);
nand U3221 (N_3221,N_1907,N_1716);
and U3222 (N_3222,N_1860,N_1686);
and U3223 (N_3223,N_716,N_692);
nor U3224 (N_3224,N_651,N_633);
and U3225 (N_3225,N_2268,N_658);
xor U3226 (N_3226,N_1714,N_594);
nand U3227 (N_3227,N_1688,N_329);
and U3228 (N_3228,N_1117,N_1994);
and U3229 (N_3229,N_984,N_2149);
or U3230 (N_3230,N_872,N_2335);
and U3231 (N_3231,N_1895,N_1770);
nor U3232 (N_3232,N_236,N_802);
nor U3233 (N_3233,N_960,N_1288);
or U3234 (N_3234,N_1225,N_706);
nor U3235 (N_3235,N_585,N_961);
and U3236 (N_3236,N_2449,N_1902);
nor U3237 (N_3237,N_215,N_1904);
nand U3238 (N_3238,N_546,N_1584);
or U3239 (N_3239,N_932,N_1307);
or U3240 (N_3240,N_2097,N_1261);
and U3241 (N_3241,N_1935,N_1464);
or U3242 (N_3242,N_2340,N_962);
nor U3243 (N_3243,N_2064,N_757);
and U3244 (N_3244,N_5,N_1471);
or U3245 (N_3245,N_1580,N_1198);
or U3246 (N_3246,N_899,N_314);
nand U3247 (N_3247,N_1179,N_632);
and U3248 (N_3248,N_245,N_2012);
nor U3249 (N_3249,N_2434,N_2202);
nor U3250 (N_3250,N_2270,N_588);
and U3251 (N_3251,N_1634,N_510);
or U3252 (N_3252,N_547,N_2159);
nand U3253 (N_3253,N_209,N_2231);
nand U3254 (N_3254,N_770,N_1292);
nor U3255 (N_3255,N_1335,N_2377);
nand U3256 (N_3256,N_638,N_279);
nand U3257 (N_3257,N_1844,N_985);
nand U3258 (N_3258,N_1610,N_433);
and U3259 (N_3259,N_2497,N_2430);
nor U3260 (N_3260,N_1450,N_509);
nand U3261 (N_3261,N_1135,N_2257);
and U3262 (N_3262,N_2401,N_1101);
and U3263 (N_3263,N_1530,N_933);
and U3264 (N_3264,N_1032,N_1663);
nand U3265 (N_3265,N_2405,N_64);
nor U3266 (N_3266,N_1399,N_515);
or U3267 (N_3267,N_1685,N_2362);
and U3268 (N_3268,N_2262,N_1987);
nor U3269 (N_3269,N_1623,N_663);
or U3270 (N_3270,N_1193,N_1102);
nand U3271 (N_3271,N_264,N_2071);
and U3272 (N_3272,N_2104,N_1829);
nor U3273 (N_3273,N_305,N_1350);
nand U3274 (N_3274,N_660,N_1857);
or U3275 (N_3275,N_2288,N_1572);
nor U3276 (N_3276,N_1837,N_1433);
nand U3277 (N_3277,N_646,N_2192);
nand U3278 (N_3278,N_1642,N_2253);
and U3279 (N_3279,N_814,N_2352);
or U3280 (N_3280,N_400,N_1416);
nor U3281 (N_3281,N_2004,N_1494);
or U3282 (N_3282,N_2310,N_571);
xor U3283 (N_3283,N_1893,N_553);
and U3284 (N_3284,N_143,N_838);
or U3285 (N_3285,N_598,N_2168);
or U3286 (N_3286,N_741,N_2393);
nor U3287 (N_3287,N_2370,N_1323);
or U3288 (N_3288,N_1513,N_2355);
nand U3289 (N_3289,N_2456,N_1298);
nor U3290 (N_3290,N_34,N_1984);
and U3291 (N_3291,N_241,N_2325);
nor U3292 (N_3292,N_1263,N_1081);
nand U3293 (N_3293,N_2277,N_2354);
or U3294 (N_3294,N_1387,N_1331);
nand U3295 (N_3295,N_680,N_1683);
or U3296 (N_3296,N_877,N_2344);
and U3297 (N_3297,N_178,N_180);
nor U3298 (N_3298,N_648,N_1931);
nand U3299 (N_3299,N_1109,N_2289);
xor U3300 (N_3300,N_24,N_1694);
nor U3301 (N_3301,N_1405,N_1246);
nor U3302 (N_3302,N_1195,N_183);
and U3303 (N_3303,N_1303,N_897);
nor U3304 (N_3304,N_1565,N_231);
nor U3305 (N_3305,N_2485,N_1769);
nand U3306 (N_3306,N_857,N_810);
nor U3307 (N_3307,N_1160,N_722);
and U3308 (N_3308,N_1302,N_2259);
nand U3309 (N_3309,N_1836,N_410);
nand U3310 (N_3310,N_2154,N_2417);
or U3311 (N_3311,N_1708,N_1480);
or U3312 (N_3312,N_1196,N_1781);
nand U3313 (N_3313,N_2452,N_434);
or U3314 (N_3314,N_1120,N_1655);
or U3315 (N_3315,N_1351,N_423);
xor U3316 (N_3316,N_234,N_1674);
or U3317 (N_3317,N_218,N_1040);
or U3318 (N_3318,N_1573,N_1400);
or U3319 (N_3319,N_589,N_644);
and U3320 (N_3320,N_2436,N_1617);
or U3321 (N_3321,N_2248,N_324);
and U3322 (N_3322,N_1917,N_199);
nand U3323 (N_3323,N_2280,N_1559);
and U3324 (N_3324,N_57,N_1966);
nor U3325 (N_3325,N_1996,N_223);
and U3326 (N_3326,N_366,N_1398);
nand U3327 (N_3327,N_2235,N_998);
and U3328 (N_3328,N_2150,N_2322);
nand U3329 (N_3329,N_376,N_1947);
or U3330 (N_3330,N_952,N_929);
nand U3331 (N_3331,N_1043,N_964);
nor U3332 (N_3332,N_1019,N_2367);
or U3333 (N_3333,N_1540,N_1166);
or U3334 (N_3334,N_1605,N_1024);
and U3335 (N_3335,N_650,N_1539);
nor U3336 (N_3336,N_1877,N_2126);
or U3337 (N_3337,N_1739,N_162);
or U3338 (N_3338,N_483,N_1408);
nor U3339 (N_3339,N_678,N_2032);
nand U3340 (N_3340,N_2006,N_1638);
nor U3341 (N_3341,N_384,N_666);
nand U3342 (N_3342,N_500,N_1297);
or U3343 (N_3343,N_205,N_656);
nand U3344 (N_3344,N_1068,N_51);
nor U3345 (N_3345,N_404,N_688);
nor U3346 (N_3346,N_106,N_1340);
and U3347 (N_3347,N_2222,N_1550);
nor U3348 (N_3348,N_1444,N_1383);
and U3349 (N_3349,N_983,N_1865);
or U3350 (N_3350,N_2455,N_1646);
nor U3351 (N_3351,N_2298,N_672);
and U3352 (N_3352,N_670,N_533);
or U3353 (N_3353,N_844,N_358);
and U3354 (N_3354,N_1983,N_950);
nor U3355 (N_3355,N_2279,N_1843);
nor U3356 (N_3356,N_1980,N_2375);
nand U3357 (N_3357,N_1502,N_1226);
or U3358 (N_3358,N_124,N_2082);
and U3359 (N_3359,N_996,N_661);
nand U3360 (N_3360,N_1157,N_1827);
or U3361 (N_3361,N_1467,N_2176);
or U3362 (N_3362,N_1342,N_1141);
nor U3363 (N_3363,N_1105,N_78);
or U3364 (N_3364,N_1455,N_1247);
nor U3365 (N_3365,N_214,N_1066);
or U3366 (N_3366,N_356,N_1446);
nor U3367 (N_3367,N_396,N_1538);
or U3368 (N_3368,N_226,N_1118);
nor U3369 (N_3369,N_548,N_2382);
or U3370 (N_3370,N_2035,N_2117);
nand U3371 (N_3371,N_2278,N_1381);
nand U3372 (N_3372,N_1521,N_2426);
or U3373 (N_3373,N_2224,N_701);
nand U3374 (N_3374,N_951,N_114);
nand U3375 (N_3375,N_2017,N_1590);
nor U3376 (N_3376,N_1218,N_516);
and U3377 (N_3377,N_1126,N_928);
or U3378 (N_3378,N_2495,N_2009);
nor U3379 (N_3379,N_2460,N_1074);
nand U3380 (N_3380,N_2140,N_1924);
nor U3381 (N_3381,N_1055,N_1621);
or U3382 (N_3382,N_1495,N_1923);
nor U3383 (N_3383,N_1622,N_740);
nand U3384 (N_3384,N_1724,N_170);
nand U3385 (N_3385,N_1641,N_1295);
nor U3386 (N_3386,N_1447,N_1072);
nor U3387 (N_3387,N_290,N_2341);
nand U3388 (N_3388,N_2113,N_1435);
nand U3389 (N_3389,N_1656,N_1701);
nor U3390 (N_3390,N_1757,N_1903);
xnor U3391 (N_3391,N_274,N_1890);
nand U3392 (N_3392,N_884,N_1596);
nor U3393 (N_3393,N_1542,N_1535);
nor U3394 (N_3394,N_1164,N_1058);
nand U3395 (N_3395,N_307,N_2185);
and U3396 (N_3396,N_2182,N_2316);
nand U3397 (N_3397,N_2028,N_81);
or U3398 (N_3398,N_861,N_318);
nor U3399 (N_3399,N_1588,N_2252);
nand U3400 (N_3400,N_2002,N_1989);
or U3401 (N_3401,N_1199,N_2135);
nand U3402 (N_3402,N_1402,N_1887);
or U3403 (N_3403,N_1346,N_377);
and U3404 (N_3404,N_52,N_1953);
nor U3405 (N_3405,N_1497,N_1817);
nand U3406 (N_3406,N_1910,N_991);
and U3407 (N_3407,N_2399,N_319);
or U3408 (N_3408,N_1751,N_1469);
nor U3409 (N_3409,N_243,N_903);
or U3410 (N_3410,N_1219,N_1326);
and U3411 (N_3411,N_676,N_873);
or U3412 (N_3412,N_856,N_196);
nor U3413 (N_3413,N_2163,N_2000);
nor U3414 (N_3414,N_132,N_1418);
nand U3415 (N_3415,N_466,N_101);
and U3416 (N_3416,N_2218,N_117);
and U3417 (N_3417,N_1915,N_317);
and U3418 (N_3418,N_1771,N_2107);
and U3419 (N_3419,N_394,N_348);
nand U3420 (N_3420,N_794,N_925);
or U3421 (N_3421,N_1473,N_2106);
nor U3422 (N_3422,N_1732,N_338);
nand U3423 (N_3423,N_819,N_2099);
or U3424 (N_3424,N_2030,N_710);
and U3425 (N_3425,N_2049,N_363);
and U3426 (N_3426,N_1025,N_1428);
nand U3427 (N_3427,N_331,N_2156);
nand U3428 (N_3428,N_1060,N_1901);
nor U3429 (N_3429,N_1544,N_1309);
nor U3430 (N_3430,N_2423,N_836);
nor U3431 (N_3431,N_629,N_616);
nor U3432 (N_3432,N_1483,N_2045);
or U3433 (N_3433,N_2454,N_1599);
and U3434 (N_3434,N_390,N_904);
nor U3435 (N_3435,N_1449,N_1914);
or U3436 (N_3436,N_986,N_2249);
and U3437 (N_3437,N_1389,N_327);
nor U3438 (N_3438,N_1866,N_1153);
and U3439 (N_3439,N_23,N_2346);
nand U3440 (N_3440,N_1414,N_1896);
xor U3441 (N_3441,N_782,N_698);
nand U3442 (N_3442,N_337,N_1129);
nor U3443 (N_3443,N_108,N_1583);
and U3444 (N_3444,N_1221,N_591);
and U3445 (N_3445,N_1612,N_1391);
nor U3446 (N_3446,N_498,N_94);
and U3447 (N_3447,N_70,N_1778);
or U3448 (N_3448,N_967,N_1277);
nand U3449 (N_3449,N_882,N_1786);
nor U3450 (N_3450,N_2027,N_1142);
nor U3451 (N_3451,N_49,N_2207);
nand U3452 (N_3452,N_2170,N_2184);
xor U3453 (N_3453,N_41,N_20);
or U3454 (N_3454,N_1206,N_1211);
nand U3455 (N_3455,N_958,N_1410);
nor U3456 (N_3456,N_775,N_937);
nand U3457 (N_3457,N_62,N_2400);
and U3458 (N_3458,N_2022,N_965);
and U3459 (N_3459,N_1740,N_570);
or U3460 (N_3460,N_1209,N_328);
and U3461 (N_3461,N_2374,N_2444);
nor U3462 (N_3462,N_549,N_927);
or U3463 (N_3463,N_1882,N_1785);
nor U3464 (N_3464,N_559,N_1846);
or U3465 (N_3465,N_767,N_491);
or U3466 (N_3466,N_1939,N_1420);
nand U3467 (N_3467,N_840,N_2336);
and U3468 (N_3468,N_1507,N_313);
nand U3469 (N_3469,N_966,N_1601);
nand U3470 (N_3470,N_2305,N_2386);
nor U3471 (N_3471,N_1029,N_1543);
nor U3472 (N_3472,N_267,N_2031);
nand U3473 (N_3473,N_1728,N_219);
or U3474 (N_3474,N_1534,N_1782);
and U3475 (N_3475,N_587,N_746);
xnor U3476 (N_3476,N_1215,N_603);
nor U3477 (N_3477,N_839,N_2446);
or U3478 (N_3478,N_2141,N_1670);
nor U3479 (N_3479,N_1848,N_1722);
or U3480 (N_3480,N_1627,N_1165);
and U3481 (N_3481,N_2048,N_2347);
and U3482 (N_3482,N_147,N_995);
nand U3483 (N_3483,N_619,N_702);
nor U3484 (N_3484,N_1145,N_1376);
or U3485 (N_3485,N_254,N_335);
nor U3486 (N_3486,N_1908,N_2223);
nor U3487 (N_3487,N_130,N_59);
or U3488 (N_3488,N_87,N_1736);
or U3489 (N_3489,N_1075,N_2358);
nor U3490 (N_3490,N_1744,N_2470);
nand U3491 (N_3491,N_1071,N_1554);
or U3492 (N_3492,N_2376,N_2328);
nand U3493 (N_3493,N_1147,N_26);
or U3494 (N_3494,N_1961,N_1252);
or U3495 (N_3495,N_1761,N_876);
nor U3496 (N_3496,N_2093,N_1063);
and U3497 (N_3497,N_1668,N_1207);
nor U3498 (N_3498,N_1678,N_158);
nor U3499 (N_3499,N_1967,N_554);
or U3500 (N_3500,N_911,N_424);
nor U3501 (N_3501,N_2333,N_2266);
nor U3502 (N_3502,N_2254,N_105);
and U3503 (N_3503,N_1640,N_1834);
or U3504 (N_3504,N_725,N_916);
or U3505 (N_3505,N_1156,N_163);
or U3506 (N_3506,N_645,N_359);
and U3507 (N_3507,N_1871,N_13);
or U3508 (N_3508,N_2068,N_470);
nand U3509 (N_3509,N_473,N_1267);
xnor U3510 (N_3510,N_1889,N_2157);
or U3511 (N_3511,N_421,N_1203);
or U3512 (N_3512,N_1955,N_136);
and U3513 (N_3513,N_2112,N_789);
and U3514 (N_3514,N_1227,N_1362);
nand U3515 (N_3515,N_2147,N_2166);
or U3516 (N_3516,N_1392,N_1385);
nand U3517 (N_3517,N_1411,N_2);
and U3518 (N_3518,N_1478,N_1415);
or U3519 (N_3519,N_2442,N_1712);
and U3520 (N_3520,N_1031,N_385);
nand U3521 (N_3521,N_654,N_532);
and U3522 (N_3522,N_98,N_379);
nor U3523 (N_3523,N_1136,N_601);
and U3524 (N_3524,N_1064,N_309);
or U3525 (N_3525,N_93,N_1287);
or U3526 (N_3526,N_777,N_1033);
and U3527 (N_3527,N_742,N_1522);
nor U3528 (N_3528,N_1748,N_1322);
and U3529 (N_3529,N_1589,N_128);
or U3530 (N_3530,N_2131,N_1991);
nor U3531 (N_3531,N_1001,N_1260);
nand U3532 (N_3532,N_1635,N_228);
nor U3533 (N_3533,N_2039,N_1023);
or U3534 (N_3534,N_901,N_1301);
and U3535 (N_3535,N_90,N_2295);
nor U3536 (N_3536,N_1825,N_785);
nor U3537 (N_3537,N_168,N_1525);
nand U3538 (N_3538,N_1553,N_2013);
or U3539 (N_3539,N_831,N_734);
nor U3540 (N_3540,N_2242,N_292);
nand U3541 (N_3541,N_1735,N_711);
nand U3542 (N_3542,N_61,N_2025);
nand U3543 (N_3543,N_1337,N_513);
and U3544 (N_3544,N_156,N_2213);
nand U3545 (N_3545,N_2052,N_2489);
or U3546 (N_3546,N_895,N_1487);
nor U3547 (N_3547,N_1608,N_1548);
nand U3548 (N_3548,N_1986,N_871);
and U3549 (N_3549,N_2144,N_890);
nand U3550 (N_3550,N_1616,N_332);
nand U3551 (N_3551,N_667,N_1172);
nor U3552 (N_3552,N_50,N_375);
and U3553 (N_3553,N_2332,N_415);
nor U3554 (N_3554,N_2356,N_1673);
nand U3555 (N_3555,N_669,N_618);
or U3556 (N_3556,N_44,N_480);
nand U3557 (N_3557,N_982,N_1488);
or U3558 (N_3558,N_1035,N_2130);
and U3559 (N_3559,N_2304,N_1429);
nand U3560 (N_3560,N_179,N_689);
and U3561 (N_3561,N_1427,N_730);
nand U3562 (N_3562,N_255,N_575);
nand U3563 (N_3563,N_1814,N_2395);
and U3564 (N_3564,N_946,N_1108);
or U3565 (N_3565,N_1669,N_2077);
nand U3566 (N_3566,N_1639,N_2272);
or U3567 (N_3567,N_2073,N_1758);
or U3568 (N_3568,N_425,N_2317);
or U3569 (N_3569,N_988,N_1594);
nand U3570 (N_3570,N_368,N_1856);
nor U3571 (N_3571,N_624,N_1361);
nand U3572 (N_3572,N_2260,N_700);
xnor U3573 (N_3573,N_46,N_1003);
and U3574 (N_3574,N_426,N_2406);
nand U3575 (N_3575,N_1067,N_1316);
nand U3576 (N_3576,N_1093,N_235);
or U3577 (N_3577,N_1965,N_345);
nor U3578 (N_3578,N_963,N_1462);
nand U3579 (N_3579,N_1706,N_216);
and U3580 (N_3580,N_1822,N_2422);
or U3581 (N_3581,N_2339,N_2348);
or U3582 (N_3582,N_412,N_620);
nand U3583 (N_3583,N_145,N_1344);
and U3584 (N_3584,N_719,N_760);
and U3585 (N_3585,N_1266,N_330);
nor U3586 (N_3586,N_198,N_1973);
nor U3587 (N_3587,N_2005,N_2476);
or U3588 (N_3588,N_1070,N_2458);
or U3589 (N_3589,N_1151,N_2115);
nand U3590 (N_3590,N_1180,N_1269);
nor U3591 (N_3591,N_1859,N_2311);
and U3592 (N_3592,N_2124,N_1878);
nor U3593 (N_3593,N_27,N_1791);
or U3594 (N_3594,N_561,N_221);
nor U3595 (N_3595,N_653,N_2152);
and U3596 (N_3596,N_935,N_341);
and U3597 (N_3597,N_512,N_310);
and U3598 (N_3598,N_1927,N_1597);
and U3599 (N_3599,N_140,N_592);
nor U3600 (N_3600,N_778,N_1652);
and U3601 (N_3601,N_1773,N_312);
and U3602 (N_3602,N_1921,N_1547);
and U3603 (N_3603,N_1352,N_1390);
nor U3604 (N_3604,N_1134,N_971);
nor U3605 (N_3605,N_2193,N_380);
nor U3606 (N_3606,N_1557,N_1468);
nand U3607 (N_3607,N_2425,N_1045);
nor U3608 (N_3608,N_907,N_1236);
or U3609 (N_3609,N_367,N_636);
or U3610 (N_3610,N_1401,N_1306);
nand U3611 (N_3611,N_2385,N_1798);
and U3612 (N_3612,N_1833,N_2098);
and U3613 (N_3613,N_25,N_1618);
nand U3614 (N_3614,N_1709,N_1725);
xor U3615 (N_3615,N_295,N_735);
nand U3616 (N_3616,N_1804,N_397);
nand U3617 (N_3617,N_573,N_2171);
nor U3618 (N_3618,N_751,N_1997);
or U3619 (N_3619,N_1650,N_2119);
nor U3620 (N_3620,N_1409,N_340);
and U3621 (N_3621,N_843,N_1516);
nor U3622 (N_3622,N_1700,N_1113);
and U3623 (N_3623,N_508,N_1508);
nand U3624 (N_3624,N_1721,N_2363);
or U3625 (N_3625,N_1026,N_2229);
or U3626 (N_3626,N_1872,N_776);
nor U3627 (N_3627,N_333,N_544);
and U3628 (N_3628,N_1096,N_1443);
nor U3629 (N_3629,N_560,N_1746);
and U3630 (N_3630,N_1426,N_527);
or U3631 (N_3631,N_2286,N_1061);
nand U3632 (N_3632,N_1975,N_2415);
or U3633 (N_3633,N_2293,N_1139);
or U3634 (N_3634,N_753,N_817);
or U3635 (N_3635,N_1133,N_402);
and U3636 (N_3636,N_1602,N_84);
nor U3637 (N_3637,N_438,N_125);
or U3638 (N_3638,N_1511,N_182);
nor U3639 (N_3639,N_919,N_1038);
nor U3640 (N_3640,N_1002,N_994);
nor U3641 (N_3641,N_447,N_1114);
xor U3642 (N_3642,N_2020,N_1492);
nand U3643 (N_3643,N_1046,N_1370);
or U3644 (N_3644,N_2475,N_2387);
and U3645 (N_3645,N_944,N_520);
nand U3646 (N_3646,N_353,N_2416);
nand U3647 (N_3647,N_541,N_637);
and U3648 (N_3648,N_1333,N_732);
or U3649 (N_3649,N_2308,N_350);
or U3650 (N_3650,N_874,N_2155);
nand U3651 (N_3651,N_387,N_924);
nand U3652 (N_3652,N_1396,N_2188);
nand U3653 (N_3653,N_2498,N_2326);
or U3654 (N_3654,N_2187,N_1788);
and U3655 (N_3655,N_558,N_1556);
nand U3656 (N_3656,N_1792,N_259);
or U3657 (N_3657,N_1107,N_1349);
nor U3658 (N_3658,N_1875,N_399);
and U3659 (N_3659,N_1278,N_58);
and U3660 (N_3660,N_1477,N_1855);
nand U3661 (N_3661,N_2001,N_2169);
or U3662 (N_3662,N_1909,N_1440);
and U3663 (N_3663,N_1152,N_459);
nor U3664 (N_3664,N_315,N_2096);
or U3665 (N_3665,N_1110,N_448);
or U3666 (N_3666,N_2255,N_1313);
and U3667 (N_3667,N_1568,N_1779);
nand U3668 (N_3668,N_2330,N_2084);
and U3669 (N_3669,N_462,N_208);
nand U3670 (N_3670,N_2083,N_2175);
nand U3671 (N_3671,N_2453,N_1111);
nor U3672 (N_3672,N_2424,N_1300);
or U3673 (N_3673,N_806,N_1698);
nor U3674 (N_3674,N_640,N_256);
nand U3675 (N_3675,N_1257,N_286);
and U3676 (N_3676,N_1658,N_184);
nor U3677 (N_3677,N_825,N_540);
or U3678 (N_3678,N_2094,N_707);
and U3679 (N_3679,N_974,N_489);
and U3680 (N_3680,N_764,N_302);
nor U3681 (N_3681,N_230,N_2471);
nand U3682 (N_3682,N_1753,N_2090);
and U3683 (N_3683,N_2388,N_160);
and U3684 (N_3684,N_613,N_2267);
or U3685 (N_3685,N_2217,N_2307);
or U3686 (N_3686,N_1373,N_1731);
nor U3687 (N_3687,N_1461,N_154);
nor U3688 (N_3688,N_1363,N_1486);
nor U3689 (N_3689,N_993,N_1090);
or U3690 (N_3690,N_2194,N_2451);
nor U3691 (N_3691,N_283,N_1217);
or U3692 (N_3692,N_936,N_2381);
nor U3693 (N_3693,N_1704,N_1039);
nand U3694 (N_3694,N_1879,N_1041);
nor U3695 (N_3695,N_1692,N_316);
and U3696 (N_3696,N_1087,N_2230);
nand U3697 (N_3697,N_1037,N_446);
or U3698 (N_3698,N_173,N_1653);
and U3699 (N_3699,N_475,N_905);
nand U3700 (N_3700,N_1765,N_889);
and U3701 (N_3701,N_1476,N_635);
nand U3702 (N_3702,N_149,N_1936);
nand U3703 (N_3703,N_538,N_2269);
nand U3704 (N_3704,N_1357,N_781);
nand U3705 (N_3705,N_1661,N_536);
nand U3706 (N_3706,N_1800,N_1796);
and U3707 (N_3707,N_779,N_1080);
and U3708 (N_3708,N_1232,N_403);
or U3709 (N_3709,N_913,N_419);
nor U3710 (N_3710,N_1676,N_1795);
or U3711 (N_3711,N_2373,N_1620);
and U3712 (N_3712,N_1106,N_2284);
nor U3713 (N_3713,N_1451,N_1259);
and U3714 (N_3714,N_2483,N_949);
or U3715 (N_3715,N_360,N_942);
or U3716 (N_3716,N_1719,N_1681);
nor U3717 (N_3717,N_2136,N_683);
xor U3718 (N_3718,N_229,N_1367);
nand U3719 (N_3719,N_222,N_1546);
or U3720 (N_3720,N_990,N_1515);
or U3721 (N_3721,N_1484,N_1649);
or U3722 (N_3722,N_1228,N_1876);
nor U3723 (N_3723,N_2189,N_1808);
nor U3724 (N_3724,N_297,N_728);
nand U3725 (N_3725,N_1854,N_2132);
and U3726 (N_3726,N_405,N_343);
and U3727 (N_3727,N_1162,N_349);
or U3728 (N_3728,N_1603,N_1926);
nand U3729 (N_3729,N_30,N_1155);
nor U3730 (N_3730,N_1679,N_2116);
nand U3731 (N_3731,N_537,N_299);
nor U3732 (N_3732,N_1174,N_1285);
or U3733 (N_3733,N_1143,N_848);
and U3734 (N_3734,N_2050,N_1948);
and U3735 (N_3735,N_2473,N_2041);
nand U3736 (N_3736,N_869,N_280);
nand U3737 (N_3737,N_1576,N_1593);
and U3738 (N_3738,N_1738,N_418);
or U3739 (N_3739,N_885,N_478);
or U3740 (N_3740,N_851,N_600);
nand U3741 (N_3741,N_807,N_2137);
and U3742 (N_3742,N_2464,N_1600);
nand U3743 (N_3743,N_714,N_449);
and U3744 (N_3744,N_2418,N_161);
nor U3745 (N_3745,N_2019,N_918);
nor U3746 (N_3746,N_2055,N_1140);
or U3747 (N_3747,N_2359,N_1007);
and U3748 (N_3748,N_112,N_1942);
or U3749 (N_3749,N_2058,N_2291);
or U3750 (N_3750,N_1718,N_426);
nor U3751 (N_3751,N_607,N_536);
and U3752 (N_3752,N_1219,N_1760);
and U3753 (N_3753,N_2426,N_364);
nand U3754 (N_3754,N_1624,N_1471);
nand U3755 (N_3755,N_1785,N_728);
and U3756 (N_3756,N_1212,N_380);
nor U3757 (N_3757,N_1765,N_1445);
nand U3758 (N_3758,N_1557,N_2261);
xor U3759 (N_3759,N_1982,N_1252);
nor U3760 (N_3760,N_1530,N_1292);
nand U3761 (N_3761,N_281,N_1224);
nor U3762 (N_3762,N_162,N_63);
and U3763 (N_3763,N_716,N_1844);
and U3764 (N_3764,N_1666,N_149);
nand U3765 (N_3765,N_980,N_925);
or U3766 (N_3766,N_1428,N_2073);
nand U3767 (N_3767,N_2274,N_312);
and U3768 (N_3768,N_406,N_636);
nand U3769 (N_3769,N_55,N_1592);
and U3770 (N_3770,N_158,N_829);
nand U3771 (N_3771,N_1140,N_942);
and U3772 (N_3772,N_903,N_793);
and U3773 (N_3773,N_2116,N_1757);
nand U3774 (N_3774,N_1296,N_2415);
nand U3775 (N_3775,N_1228,N_2333);
nand U3776 (N_3776,N_1237,N_2156);
and U3777 (N_3777,N_1213,N_1535);
xnor U3778 (N_3778,N_1652,N_1079);
nand U3779 (N_3779,N_939,N_1246);
and U3780 (N_3780,N_1506,N_1932);
nand U3781 (N_3781,N_1775,N_1338);
nand U3782 (N_3782,N_1357,N_1915);
or U3783 (N_3783,N_1544,N_1062);
nor U3784 (N_3784,N_88,N_1323);
nand U3785 (N_3785,N_1010,N_1641);
nor U3786 (N_3786,N_1231,N_84);
and U3787 (N_3787,N_1438,N_1691);
nor U3788 (N_3788,N_2137,N_319);
nor U3789 (N_3789,N_611,N_1413);
or U3790 (N_3790,N_1336,N_1543);
or U3791 (N_3791,N_1247,N_1163);
or U3792 (N_3792,N_1716,N_1533);
or U3793 (N_3793,N_2067,N_683);
nand U3794 (N_3794,N_2242,N_95);
nand U3795 (N_3795,N_1834,N_2353);
nor U3796 (N_3796,N_890,N_2261);
nor U3797 (N_3797,N_2098,N_2);
nor U3798 (N_3798,N_1082,N_1789);
nand U3799 (N_3799,N_752,N_598);
nand U3800 (N_3800,N_2067,N_2193);
nand U3801 (N_3801,N_508,N_1070);
or U3802 (N_3802,N_1943,N_352);
or U3803 (N_3803,N_1185,N_686);
and U3804 (N_3804,N_1695,N_2447);
nor U3805 (N_3805,N_1645,N_1371);
or U3806 (N_3806,N_347,N_25);
and U3807 (N_3807,N_2431,N_669);
nor U3808 (N_3808,N_916,N_1674);
and U3809 (N_3809,N_1981,N_679);
and U3810 (N_3810,N_1778,N_2091);
nand U3811 (N_3811,N_365,N_74);
and U3812 (N_3812,N_1422,N_1309);
xor U3813 (N_3813,N_2152,N_1608);
nor U3814 (N_3814,N_2314,N_636);
nor U3815 (N_3815,N_71,N_807);
and U3816 (N_3816,N_2105,N_1901);
and U3817 (N_3817,N_1477,N_1063);
or U3818 (N_3818,N_908,N_2392);
or U3819 (N_3819,N_1722,N_748);
nand U3820 (N_3820,N_28,N_1177);
nand U3821 (N_3821,N_544,N_1272);
nand U3822 (N_3822,N_846,N_1149);
or U3823 (N_3823,N_1361,N_2366);
and U3824 (N_3824,N_1367,N_1257);
nor U3825 (N_3825,N_1306,N_366);
nor U3826 (N_3826,N_579,N_737);
nor U3827 (N_3827,N_901,N_1033);
nand U3828 (N_3828,N_55,N_2219);
nand U3829 (N_3829,N_1614,N_2139);
nor U3830 (N_3830,N_447,N_2413);
or U3831 (N_3831,N_1403,N_2427);
and U3832 (N_3832,N_1425,N_1842);
and U3833 (N_3833,N_2392,N_1234);
or U3834 (N_3834,N_78,N_2424);
or U3835 (N_3835,N_665,N_568);
or U3836 (N_3836,N_2305,N_2036);
or U3837 (N_3837,N_2070,N_2204);
or U3838 (N_3838,N_133,N_10);
and U3839 (N_3839,N_1829,N_23);
nand U3840 (N_3840,N_678,N_2120);
nand U3841 (N_3841,N_111,N_363);
and U3842 (N_3842,N_583,N_1738);
and U3843 (N_3843,N_1661,N_1792);
or U3844 (N_3844,N_1817,N_1838);
nand U3845 (N_3845,N_526,N_2162);
or U3846 (N_3846,N_2191,N_273);
nor U3847 (N_3847,N_1299,N_337);
nor U3848 (N_3848,N_1800,N_2173);
nand U3849 (N_3849,N_2272,N_1416);
nor U3850 (N_3850,N_2151,N_538);
nand U3851 (N_3851,N_1505,N_367);
nand U3852 (N_3852,N_590,N_707);
and U3853 (N_3853,N_1630,N_1759);
or U3854 (N_3854,N_949,N_602);
or U3855 (N_3855,N_131,N_1974);
and U3856 (N_3856,N_1189,N_311);
or U3857 (N_3857,N_338,N_1565);
nand U3858 (N_3858,N_472,N_1909);
nor U3859 (N_3859,N_490,N_2337);
and U3860 (N_3860,N_1690,N_501);
and U3861 (N_3861,N_1336,N_2145);
or U3862 (N_3862,N_1504,N_980);
and U3863 (N_3863,N_1397,N_2075);
nand U3864 (N_3864,N_2459,N_1653);
nand U3865 (N_3865,N_2332,N_327);
nor U3866 (N_3866,N_197,N_2221);
nor U3867 (N_3867,N_1625,N_1138);
or U3868 (N_3868,N_885,N_373);
and U3869 (N_3869,N_2408,N_1887);
and U3870 (N_3870,N_1431,N_147);
nor U3871 (N_3871,N_1780,N_2311);
nor U3872 (N_3872,N_2239,N_452);
or U3873 (N_3873,N_399,N_577);
and U3874 (N_3874,N_679,N_1905);
and U3875 (N_3875,N_1139,N_1957);
nand U3876 (N_3876,N_192,N_257);
or U3877 (N_3877,N_1007,N_334);
nor U3878 (N_3878,N_2438,N_1537);
or U3879 (N_3879,N_1329,N_1013);
nand U3880 (N_3880,N_1241,N_704);
nand U3881 (N_3881,N_2095,N_2192);
and U3882 (N_3882,N_1892,N_1511);
nor U3883 (N_3883,N_1716,N_986);
and U3884 (N_3884,N_2211,N_1704);
and U3885 (N_3885,N_1255,N_463);
nand U3886 (N_3886,N_1736,N_1997);
and U3887 (N_3887,N_2160,N_1209);
and U3888 (N_3888,N_1439,N_590);
or U3889 (N_3889,N_1939,N_564);
and U3890 (N_3890,N_602,N_371);
nand U3891 (N_3891,N_129,N_1647);
nor U3892 (N_3892,N_2297,N_2376);
and U3893 (N_3893,N_505,N_1276);
nor U3894 (N_3894,N_996,N_135);
and U3895 (N_3895,N_2216,N_1405);
or U3896 (N_3896,N_2294,N_1260);
or U3897 (N_3897,N_279,N_753);
or U3898 (N_3898,N_1071,N_857);
nand U3899 (N_3899,N_1717,N_2444);
and U3900 (N_3900,N_2393,N_1947);
nand U3901 (N_3901,N_727,N_14);
nor U3902 (N_3902,N_488,N_1189);
or U3903 (N_3903,N_1530,N_206);
nor U3904 (N_3904,N_1649,N_1099);
and U3905 (N_3905,N_173,N_154);
nand U3906 (N_3906,N_2480,N_137);
or U3907 (N_3907,N_1867,N_1951);
or U3908 (N_3908,N_190,N_1777);
and U3909 (N_3909,N_2262,N_2291);
nand U3910 (N_3910,N_2001,N_508);
and U3911 (N_3911,N_32,N_926);
or U3912 (N_3912,N_310,N_2481);
or U3913 (N_3913,N_1034,N_1111);
nor U3914 (N_3914,N_211,N_1616);
nand U3915 (N_3915,N_255,N_346);
and U3916 (N_3916,N_1374,N_1943);
and U3917 (N_3917,N_281,N_381);
nand U3918 (N_3918,N_1950,N_2433);
nand U3919 (N_3919,N_1088,N_2120);
and U3920 (N_3920,N_286,N_1743);
nand U3921 (N_3921,N_2132,N_1575);
and U3922 (N_3922,N_1799,N_523);
and U3923 (N_3923,N_1033,N_1609);
and U3924 (N_3924,N_1993,N_1863);
or U3925 (N_3925,N_2465,N_1989);
nor U3926 (N_3926,N_265,N_782);
nand U3927 (N_3927,N_803,N_1049);
nor U3928 (N_3928,N_788,N_89);
or U3929 (N_3929,N_885,N_1092);
or U3930 (N_3930,N_118,N_2062);
nand U3931 (N_3931,N_420,N_1513);
and U3932 (N_3932,N_2357,N_2205);
and U3933 (N_3933,N_906,N_1896);
and U3934 (N_3934,N_1657,N_1199);
nand U3935 (N_3935,N_1585,N_982);
and U3936 (N_3936,N_339,N_2088);
and U3937 (N_3937,N_2455,N_238);
or U3938 (N_3938,N_553,N_825);
nand U3939 (N_3939,N_1526,N_644);
and U3940 (N_3940,N_2154,N_1465);
and U3941 (N_3941,N_2321,N_654);
and U3942 (N_3942,N_711,N_380);
and U3943 (N_3943,N_1384,N_1382);
nor U3944 (N_3944,N_216,N_1609);
nand U3945 (N_3945,N_1180,N_2207);
nor U3946 (N_3946,N_1854,N_1795);
nor U3947 (N_3947,N_1586,N_1018);
and U3948 (N_3948,N_1084,N_1851);
and U3949 (N_3949,N_2299,N_530);
or U3950 (N_3950,N_1781,N_1996);
and U3951 (N_3951,N_2118,N_2478);
and U3952 (N_3952,N_193,N_1818);
nor U3953 (N_3953,N_1867,N_988);
nand U3954 (N_3954,N_1733,N_427);
and U3955 (N_3955,N_2311,N_260);
and U3956 (N_3956,N_2150,N_1054);
or U3957 (N_3957,N_2161,N_626);
or U3958 (N_3958,N_16,N_1658);
and U3959 (N_3959,N_1609,N_778);
nand U3960 (N_3960,N_985,N_2276);
and U3961 (N_3961,N_2071,N_1421);
and U3962 (N_3962,N_517,N_205);
and U3963 (N_3963,N_362,N_2146);
nand U3964 (N_3964,N_1249,N_1799);
or U3965 (N_3965,N_727,N_434);
or U3966 (N_3966,N_2127,N_1485);
and U3967 (N_3967,N_2432,N_218);
nand U3968 (N_3968,N_693,N_1552);
and U3969 (N_3969,N_877,N_2175);
nor U3970 (N_3970,N_359,N_1074);
nand U3971 (N_3971,N_1288,N_1885);
and U3972 (N_3972,N_2080,N_874);
nor U3973 (N_3973,N_1766,N_1450);
nor U3974 (N_3974,N_1156,N_244);
nand U3975 (N_3975,N_302,N_1161);
nor U3976 (N_3976,N_245,N_2150);
and U3977 (N_3977,N_1585,N_1400);
nor U3978 (N_3978,N_1518,N_1103);
nor U3979 (N_3979,N_198,N_581);
and U3980 (N_3980,N_218,N_604);
nor U3981 (N_3981,N_1210,N_445);
or U3982 (N_3982,N_958,N_2388);
nand U3983 (N_3983,N_1042,N_364);
nand U3984 (N_3984,N_2291,N_587);
nor U3985 (N_3985,N_579,N_751);
nand U3986 (N_3986,N_740,N_17);
nor U3987 (N_3987,N_1906,N_212);
and U3988 (N_3988,N_2322,N_257);
nand U3989 (N_3989,N_513,N_775);
and U3990 (N_3990,N_2374,N_320);
or U3991 (N_3991,N_980,N_687);
nand U3992 (N_3992,N_436,N_1435);
or U3993 (N_3993,N_1503,N_743);
and U3994 (N_3994,N_1317,N_881);
nor U3995 (N_3995,N_2158,N_1625);
and U3996 (N_3996,N_2106,N_178);
or U3997 (N_3997,N_2325,N_2);
and U3998 (N_3998,N_2345,N_1972);
or U3999 (N_3999,N_650,N_1173);
and U4000 (N_4000,N_1820,N_416);
nor U4001 (N_4001,N_2422,N_74);
nor U4002 (N_4002,N_873,N_1512);
nand U4003 (N_4003,N_2149,N_2494);
and U4004 (N_4004,N_2221,N_2334);
nand U4005 (N_4005,N_884,N_1646);
and U4006 (N_4006,N_2425,N_712);
nor U4007 (N_4007,N_1804,N_78);
nand U4008 (N_4008,N_2313,N_2453);
or U4009 (N_4009,N_1363,N_2376);
nor U4010 (N_4010,N_338,N_1682);
xnor U4011 (N_4011,N_2182,N_423);
nand U4012 (N_4012,N_1058,N_212);
nor U4013 (N_4013,N_2316,N_2399);
nand U4014 (N_4014,N_462,N_2149);
and U4015 (N_4015,N_2377,N_888);
or U4016 (N_4016,N_460,N_1991);
nor U4017 (N_4017,N_1464,N_1457);
nor U4018 (N_4018,N_1997,N_2084);
and U4019 (N_4019,N_1609,N_182);
and U4020 (N_4020,N_1032,N_688);
nor U4021 (N_4021,N_2199,N_467);
or U4022 (N_4022,N_1131,N_1776);
or U4023 (N_4023,N_2497,N_1521);
or U4024 (N_4024,N_1705,N_92);
nor U4025 (N_4025,N_104,N_2497);
nor U4026 (N_4026,N_1780,N_203);
and U4027 (N_4027,N_2145,N_1651);
nand U4028 (N_4028,N_2226,N_1966);
nand U4029 (N_4029,N_481,N_413);
or U4030 (N_4030,N_2458,N_147);
nor U4031 (N_4031,N_1303,N_1957);
nand U4032 (N_4032,N_715,N_2049);
or U4033 (N_4033,N_1576,N_984);
or U4034 (N_4034,N_468,N_76);
and U4035 (N_4035,N_1175,N_1315);
nand U4036 (N_4036,N_1878,N_2411);
and U4037 (N_4037,N_282,N_1793);
nand U4038 (N_4038,N_894,N_1584);
and U4039 (N_4039,N_138,N_954);
nor U4040 (N_4040,N_489,N_673);
or U4041 (N_4041,N_1436,N_1860);
nand U4042 (N_4042,N_2206,N_19);
nor U4043 (N_4043,N_316,N_311);
nor U4044 (N_4044,N_1987,N_2015);
and U4045 (N_4045,N_926,N_2088);
or U4046 (N_4046,N_1990,N_1776);
nand U4047 (N_4047,N_1021,N_247);
or U4048 (N_4048,N_1132,N_907);
and U4049 (N_4049,N_2023,N_97);
nor U4050 (N_4050,N_2338,N_606);
or U4051 (N_4051,N_1615,N_2358);
and U4052 (N_4052,N_1219,N_1290);
and U4053 (N_4053,N_115,N_1748);
or U4054 (N_4054,N_392,N_1254);
nor U4055 (N_4055,N_250,N_1103);
and U4056 (N_4056,N_1486,N_2492);
nand U4057 (N_4057,N_342,N_481);
or U4058 (N_4058,N_1602,N_704);
nand U4059 (N_4059,N_1277,N_1998);
nand U4060 (N_4060,N_875,N_1600);
or U4061 (N_4061,N_1995,N_1416);
or U4062 (N_4062,N_201,N_610);
or U4063 (N_4063,N_920,N_508);
or U4064 (N_4064,N_1908,N_733);
and U4065 (N_4065,N_454,N_617);
nand U4066 (N_4066,N_786,N_757);
nor U4067 (N_4067,N_1550,N_470);
nor U4068 (N_4068,N_283,N_1079);
or U4069 (N_4069,N_1211,N_715);
nand U4070 (N_4070,N_702,N_2446);
or U4071 (N_4071,N_1749,N_416);
nand U4072 (N_4072,N_1941,N_238);
or U4073 (N_4073,N_537,N_181);
and U4074 (N_4074,N_1145,N_1439);
and U4075 (N_4075,N_1755,N_2497);
and U4076 (N_4076,N_1071,N_1777);
or U4077 (N_4077,N_1782,N_921);
or U4078 (N_4078,N_1647,N_858);
or U4079 (N_4079,N_240,N_408);
and U4080 (N_4080,N_557,N_2304);
nor U4081 (N_4081,N_2337,N_2183);
and U4082 (N_4082,N_1530,N_1462);
or U4083 (N_4083,N_924,N_2350);
or U4084 (N_4084,N_1972,N_1579);
nand U4085 (N_4085,N_429,N_403);
nor U4086 (N_4086,N_1701,N_967);
nor U4087 (N_4087,N_2163,N_470);
and U4088 (N_4088,N_880,N_61);
or U4089 (N_4089,N_308,N_1876);
nand U4090 (N_4090,N_46,N_2099);
and U4091 (N_4091,N_579,N_956);
and U4092 (N_4092,N_588,N_10);
nand U4093 (N_4093,N_1265,N_15);
and U4094 (N_4094,N_1865,N_1338);
and U4095 (N_4095,N_2313,N_1730);
or U4096 (N_4096,N_50,N_1062);
nor U4097 (N_4097,N_1960,N_1378);
nand U4098 (N_4098,N_2236,N_1719);
or U4099 (N_4099,N_1046,N_845);
and U4100 (N_4100,N_1702,N_1866);
and U4101 (N_4101,N_1038,N_2497);
nand U4102 (N_4102,N_2279,N_119);
and U4103 (N_4103,N_2224,N_2377);
nand U4104 (N_4104,N_1211,N_593);
or U4105 (N_4105,N_453,N_1028);
nand U4106 (N_4106,N_1316,N_731);
nand U4107 (N_4107,N_1049,N_2262);
or U4108 (N_4108,N_2019,N_2364);
nor U4109 (N_4109,N_1165,N_2184);
nor U4110 (N_4110,N_2311,N_2120);
or U4111 (N_4111,N_596,N_2128);
nand U4112 (N_4112,N_357,N_50);
and U4113 (N_4113,N_785,N_1286);
and U4114 (N_4114,N_2428,N_2013);
and U4115 (N_4115,N_1444,N_2263);
or U4116 (N_4116,N_294,N_1835);
nand U4117 (N_4117,N_2060,N_1968);
and U4118 (N_4118,N_1793,N_491);
or U4119 (N_4119,N_113,N_266);
and U4120 (N_4120,N_2120,N_670);
and U4121 (N_4121,N_925,N_313);
nor U4122 (N_4122,N_1094,N_669);
or U4123 (N_4123,N_2019,N_545);
and U4124 (N_4124,N_1629,N_586);
xor U4125 (N_4125,N_129,N_1429);
nand U4126 (N_4126,N_1337,N_1640);
nor U4127 (N_4127,N_1161,N_1474);
nor U4128 (N_4128,N_102,N_1918);
or U4129 (N_4129,N_388,N_572);
or U4130 (N_4130,N_1264,N_1062);
and U4131 (N_4131,N_1453,N_1777);
xor U4132 (N_4132,N_1383,N_1150);
and U4133 (N_4133,N_2364,N_947);
nor U4134 (N_4134,N_1306,N_1390);
nor U4135 (N_4135,N_821,N_448);
or U4136 (N_4136,N_512,N_2061);
nor U4137 (N_4137,N_2226,N_1454);
nand U4138 (N_4138,N_263,N_2141);
and U4139 (N_4139,N_138,N_616);
and U4140 (N_4140,N_426,N_2384);
and U4141 (N_4141,N_757,N_1154);
and U4142 (N_4142,N_1114,N_1935);
nor U4143 (N_4143,N_2079,N_382);
or U4144 (N_4144,N_678,N_1411);
and U4145 (N_4145,N_1043,N_1567);
and U4146 (N_4146,N_2263,N_1906);
nor U4147 (N_4147,N_258,N_955);
or U4148 (N_4148,N_1642,N_631);
and U4149 (N_4149,N_319,N_1729);
and U4150 (N_4150,N_1323,N_52);
or U4151 (N_4151,N_516,N_1783);
nor U4152 (N_4152,N_1713,N_2030);
nor U4153 (N_4153,N_1093,N_2108);
nor U4154 (N_4154,N_2197,N_2161);
and U4155 (N_4155,N_951,N_2097);
nand U4156 (N_4156,N_382,N_1954);
and U4157 (N_4157,N_700,N_885);
nand U4158 (N_4158,N_1364,N_1676);
nor U4159 (N_4159,N_283,N_1913);
nor U4160 (N_4160,N_273,N_413);
and U4161 (N_4161,N_1851,N_2325);
or U4162 (N_4162,N_1853,N_1102);
and U4163 (N_4163,N_1183,N_962);
or U4164 (N_4164,N_585,N_1563);
or U4165 (N_4165,N_1234,N_2286);
and U4166 (N_4166,N_204,N_1624);
nand U4167 (N_4167,N_2159,N_1083);
nand U4168 (N_4168,N_2147,N_783);
or U4169 (N_4169,N_736,N_967);
and U4170 (N_4170,N_2085,N_386);
nand U4171 (N_4171,N_1238,N_2428);
nor U4172 (N_4172,N_1008,N_464);
and U4173 (N_4173,N_2071,N_1326);
nor U4174 (N_4174,N_1077,N_52);
or U4175 (N_4175,N_702,N_1603);
nor U4176 (N_4176,N_1193,N_448);
or U4177 (N_4177,N_2409,N_62);
nor U4178 (N_4178,N_1188,N_1317);
and U4179 (N_4179,N_366,N_1855);
nor U4180 (N_4180,N_1845,N_1265);
or U4181 (N_4181,N_2357,N_533);
and U4182 (N_4182,N_832,N_60);
nor U4183 (N_4183,N_23,N_1828);
xor U4184 (N_4184,N_471,N_748);
nand U4185 (N_4185,N_1709,N_2241);
nor U4186 (N_4186,N_2384,N_1047);
nand U4187 (N_4187,N_304,N_754);
and U4188 (N_4188,N_1615,N_1391);
or U4189 (N_4189,N_67,N_1255);
or U4190 (N_4190,N_1595,N_1896);
and U4191 (N_4191,N_2321,N_117);
and U4192 (N_4192,N_1603,N_2148);
nand U4193 (N_4193,N_2258,N_2286);
nor U4194 (N_4194,N_2124,N_919);
xnor U4195 (N_4195,N_2248,N_99);
xor U4196 (N_4196,N_1603,N_441);
nand U4197 (N_4197,N_1181,N_2057);
or U4198 (N_4198,N_784,N_467);
and U4199 (N_4199,N_1051,N_1281);
and U4200 (N_4200,N_821,N_1910);
nand U4201 (N_4201,N_2136,N_541);
nor U4202 (N_4202,N_2339,N_2267);
and U4203 (N_4203,N_64,N_2198);
and U4204 (N_4204,N_697,N_2489);
nor U4205 (N_4205,N_2428,N_1444);
xnor U4206 (N_4206,N_960,N_1565);
or U4207 (N_4207,N_654,N_1416);
nor U4208 (N_4208,N_287,N_633);
nand U4209 (N_4209,N_1618,N_431);
or U4210 (N_4210,N_261,N_1435);
nand U4211 (N_4211,N_1206,N_659);
nor U4212 (N_4212,N_1929,N_1737);
or U4213 (N_4213,N_1092,N_1943);
nor U4214 (N_4214,N_1225,N_2182);
or U4215 (N_4215,N_543,N_2266);
and U4216 (N_4216,N_1149,N_746);
nor U4217 (N_4217,N_261,N_2383);
and U4218 (N_4218,N_2249,N_251);
nor U4219 (N_4219,N_55,N_180);
or U4220 (N_4220,N_442,N_135);
nand U4221 (N_4221,N_1894,N_506);
nand U4222 (N_4222,N_2419,N_564);
or U4223 (N_4223,N_1850,N_1855);
and U4224 (N_4224,N_26,N_2453);
nand U4225 (N_4225,N_1886,N_2449);
or U4226 (N_4226,N_499,N_1151);
or U4227 (N_4227,N_2419,N_586);
or U4228 (N_4228,N_2205,N_1749);
or U4229 (N_4229,N_2429,N_1260);
nand U4230 (N_4230,N_1659,N_1020);
nor U4231 (N_4231,N_1087,N_1346);
nor U4232 (N_4232,N_1761,N_2154);
or U4233 (N_4233,N_190,N_592);
and U4234 (N_4234,N_566,N_901);
or U4235 (N_4235,N_111,N_1431);
nor U4236 (N_4236,N_1210,N_2230);
or U4237 (N_4237,N_1911,N_1885);
nor U4238 (N_4238,N_1275,N_783);
nor U4239 (N_4239,N_1979,N_2066);
nand U4240 (N_4240,N_119,N_351);
or U4241 (N_4241,N_1392,N_425);
and U4242 (N_4242,N_2149,N_1606);
nor U4243 (N_4243,N_1821,N_1778);
nor U4244 (N_4244,N_1496,N_155);
or U4245 (N_4245,N_1416,N_1944);
and U4246 (N_4246,N_1072,N_2362);
nand U4247 (N_4247,N_438,N_388);
or U4248 (N_4248,N_2215,N_544);
or U4249 (N_4249,N_1445,N_1728);
and U4250 (N_4250,N_352,N_1425);
or U4251 (N_4251,N_1623,N_1237);
or U4252 (N_4252,N_118,N_2295);
or U4253 (N_4253,N_1295,N_1611);
nand U4254 (N_4254,N_1606,N_19);
or U4255 (N_4255,N_813,N_194);
and U4256 (N_4256,N_667,N_2421);
or U4257 (N_4257,N_2118,N_2425);
nor U4258 (N_4258,N_1436,N_401);
or U4259 (N_4259,N_923,N_1525);
and U4260 (N_4260,N_2068,N_40);
or U4261 (N_4261,N_1118,N_702);
nor U4262 (N_4262,N_910,N_324);
and U4263 (N_4263,N_1081,N_79);
nand U4264 (N_4264,N_991,N_2050);
nor U4265 (N_4265,N_2208,N_1642);
and U4266 (N_4266,N_129,N_743);
nor U4267 (N_4267,N_970,N_1992);
and U4268 (N_4268,N_2001,N_85);
nor U4269 (N_4269,N_2207,N_1002);
or U4270 (N_4270,N_2339,N_888);
nand U4271 (N_4271,N_2480,N_1643);
or U4272 (N_4272,N_1820,N_2136);
and U4273 (N_4273,N_1899,N_1973);
or U4274 (N_4274,N_2268,N_337);
and U4275 (N_4275,N_1305,N_262);
nor U4276 (N_4276,N_2422,N_984);
nor U4277 (N_4277,N_2338,N_1786);
nor U4278 (N_4278,N_2467,N_2179);
and U4279 (N_4279,N_1323,N_1716);
or U4280 (N_4280,N_1795,N_803);
or U4281 (N_4281,N_818,N_305);
nor U4282 (N_4282,N_226,N_1829);
or U4283 (N_4283,N_892,N_396);
or U4284 (N_4284,N_857,N_1633);
and U4285 (N_4285,N_2194,N_2144);
nor U4286 (N_4286,N_1172,N_1819);
and U4287 (N_4287,N_120,N_489);
nand U4288 (N_4288,N_741,N_1746);
or U4289 (N_4289,N_1605,N_1895);
and U4290 (N_4290,N_2025,N_766);
or U4291 (N_4291,N_1675,N_2112);
nor U4292 (N_4292,N_585,N_2271);
or U4293 (N_4293,N_838,N_452);
and U4294 (N_4294,N_1878,N_2362);
nor U4295 (N_4295,N_1414,N_780);
nand U4296 (N_4296,N_1728,N_1162);
nor U4297 (N_4297,N_2194,N_1850);
or U4298 (N_4298,N_1270,N_710);
nand U4299 (N_4299,N_837,N_1517);
or U4300 (N_4300,N_1833,N_1142);
nand U4301 (N_4301,N_1024,N_592);
or U4302 (N_4302,N_1831,N_2137);
or U4303 (N_4303,N_1275,N_693);
or U4304 (N_4304,N_1111,N_284);
and U4305 (N_4305,N_862,N_1074);
or U4306 (N_4306,N_240,N_8);
and U4307 (N_4307,N_279,N_1798);
nor U4308 (N_4308,N_1371,N_2492);
or U4309 (N_4309,N_2426,N_1161);
or U4310 (N_4310,N_1580,N_2130);
or U4311 (N_4311,N_838,N_573);
nor U4312 (N_4312,N_1182,N_1579);
or U4313 (N_4313,N_2340,N_48);
or U4314 (N_4314,N_953,N_1014);
nand U4315 (N_4315,N_1031,N_750);
or U4316 (N_4316,N_2043,N_1446);
and U4317 (N_4317,N_361,N_1054);
nor U4318 (N_4318,N_2058,N_522);
and U4319 (N_4319,N_963,N_1309);
and U4320 (N_4320,N_2210,N_1923);
nand U4321 (N_4321,N_283,N_1336);
and U4322 (N_4322,N_199,N_1345);
or U4323 (N_4323,N_1994,N_2179);
nor U4324 (N_4324,N_2277,N_34);
and U4325 (N_4325,N_2104,N_484);
nor U4326 (N_4326,N_179,N_348);
and U4327 (N_4327,N_1055,N_1820);
nand U4328 (N_4328,N_1488,N_2083);
nor U4329 (N_4329,N_174,N_1737);
or U4330 (N_4330,N_2136,N_2429);
or U4331 (N_4331,N_1686,N_300);
nand U4332 (N_4332,N_2073,N_1136);
nand U4333 (N_4333,N_483,N_1067);
nand U4334 (N_4334,N_984,N_1176);
or U4335 (N_4335,N_1333,N_1865);
nor U4336 (N_4336,N_2011,N_681);
and U4337 (N_4337,N_2370,N_1239);
nor U4338 (N_4338,N_407,N_295);
and U4339 (N_4339,N_946,N_1644);
nand U4340 (N_4340,N_2,N_1557);
nor U4341 (N_4341,N_1671,N_381);
and U4342 (N_4342,N_368,N_718);
nor U4343 (N_4343,N_1816,N_666);
nand U4344 (N_4344,N_2160,N_586);
nor U4345 (N_4345,N_1998,N_1822);
nand U4346 (N_4346,N_1406,N_993);
nor U4347 (N_4347,N_988,N_1023);
nor U4348 (N_4348,N_1855,N_1709);
nand U4349 (N_4349,N_17,N_2021);
nor U4350 (N_4350,N_623,N_2146);
or U4351 (N_4351,N_1958,N_653);
and U4352 (N_4352,N_1245,N_928);
nor U4353 (N_4353,N_726,N_2033);
and U4354 (N_4354,N_1784,N_679);
nand U4355 (N_4355,N_468,N_1726);
and U4356 (N_4356,N_200,N_1565);
and U4357 (N_4357,N_1565,N_1996);
and U4358 (N_4358,N_1654,N_1590);
nor U4359 (N_4359,N_964,N_1342);
nand U4360 (N_4360,N_230,N_1301);
nor U4361 (N_4361,N_160,N_348);
or U4362 (N_4362,N_741,N_2270);
nand U4363 (N_4363,N_2163,N_1315);
nor U4364 (N_4364,N_214,N_2348);
nand U4365 (N_4365,N_1782,N_1015);
or U4366 (N_4366,N_308,N_623);
nand U4367 (N_4367,N_705,N_1331);
nor U4368 (N_4368,N_33,N_651);
or U4369 (N_4369,N_844,N_2295);
or U4370 (N_4370,N_2080,N_980);
nor U4371 (N_4371,N_1602,N_2088);
or U4372 (N_4372,N_1733,N_2471);
nand U4373 (N_4373,N_2055,N_1580);
nor U4374 (N_4374,N_1912,N_1130);
nand U4375 (N_4375,N_1117,N_1628);
nor U4376 (N_4376,N_1659,N_2172);
nor U4377 (N_4377,N_1344,N_1975);
and U4378 (N_4378,N_1248,N_957);
nand U4379 (N_4379,N_85,N_1182);
nor U4380 (N_4380,N_1800,N_1899);
nor U4381 (N_4381,N_363,N_1916);
nand U4382 (N_4382,N_1915,N_2168);
nor U4383 (N_4383,N_671,N_1039);
nor U4384 (N_4384,N_271,N_963);
nand U4385 (N_4385,N_1400,N_1779);
nand U4386 (N_4386,N_1642,N_1025);
nor U4387 (N_4387,N_856,N_711);
nand U4388 (N_4388,N_1846,N_1129);
and U4389 (N_4389,N_71,N_1471);
and U4390 (N_4390,N_1294,N_1597);
nor U4391 (N_4391,N_888,N_493);
or U4392 (N_4392,N_1818,N_2257);
or U4393 (N_4393,N_1420,N_2085);
and U4394 (N_4394,N_1931,N_436);
nor U4395 (N_4395,N_1885,N_1104);
nand U4396 (N_4396,N_682,N_2335);
nand U4397 (N_4397,N_162,N_1334);
or U4398 (N_4398,N_83,N_2328);
nand U4399 (N_4399,N_2236,N_2218);
and U4400 (N_4400,N_1764,N_1241);
and U4401 (N_4401,N_702,N_1827);
nor U4402 (N_4402,N_1304,N_279);
or U4403 (N_4403,N_101,N_1745);
nor U4404 (N_4404,N_395,N_1906);
and U4405 (N_4405,N_2126,N_2108);
or U4406 (N_4406,N_958,N_632);
and U4407 (N_4407,N_4,N_1905);
and U4408 (N_4408,N_2191,N_153);
nor U4409 (N_4409,N_781,N_214);
and U4410 (N_4410,N_227,N_410);
nor U4411 (N_4411,N_1244,N_2404);
nand U4412 (N_4412,N_1533,N_2345);
nand U4413 (N_4413,N_1290,N_250);
nand U4414 (N_4414,N_1150,N_2335);
nand U4415 (N_4415,N_714,N_2092);
and U4416 (N_4416,N_2030,N_2093);
nor U4417 (N_4417,N_487,N_1906);
and U4418 (N_4418,N_911,N_499);
nor U4419 (N_4419,N_1635,N_918);
nand U4420 (N_4420,N_1908,N_1122);
or U4421 (N_4421,N_69,N_978);
nor U4422 (N_4422,N_290,N_1127);
nand U4423 (N_4423,N_1867,N_923);
nor U4424 (N_4424,N_161,N_34);
or U4425 (N_4425,N_2173,N_718);
and U4426 (N_4426,N_317,N_538);
nand U4427 (N_4427,N_808,N_1806);
nand U4428 (N_4428,N_283,N_606);
nand U4429 (N_4429,N_376,N_2034);
or U4430 (N_4430,N_700,N_1898);
or U4431 (N_4431,N_431,N_996);
nor U4432 (N_4432,N_354,N_1597);
and U4433 (N_4433,N_166,N_1697);
and U4434 (N_4434,N_1044,N_1601);
or U4435 (N_4435,N_894,N_188);
or U4436 (N_4436,N_1355,N_2200);
or U4437 (N_4437,N_2260,N_1903);
nand U4438 (N_4438,N_6,N_2403);
nand U4439 (N_4439,N_343,N_1801);
nand U4440 (N_4440,N_647,N_404);
and U4441 (N_4441,N_1607,N_1822);
nand U4442 (N_4442,N_1907,N_961);
nand U4443 (N_4443,N_920,N_1906);
nand U4444 (N_4444,N_692,N_31);
or U4445 (N_4445,N_1231,N_136);
or U4446 (N_4446,N_621,N_1559);
nor U4447 (N_4447,N_29,N_1570);
nand U4448 (N_4448,N_2003,N_110);
and U4449 (N_4449,N_497,N_2264);
nand U4450 (N_4450,N_2085,N_2280);
nor U4451 (N_4451,N_283,N_1169);
nand U4452 (N_4452,N_129,N_2254);
or U4453 (N_4453,N_223,N_1570);
nor U4454 (N_4454,N_7,N_897);
and U4455 (N_4455,N_1954,N_2068);
or U4456 (N_4456,N_1702,N_1764);
and U4457 (N_4457,N_656,N_33);
nand U4458 (N_4458,N_63,N_1270);
nor U4459 (N_4459,N_1971,N_347);
nor U4460 (N_4460,N_2070,N_751);
nor U4461 (N_4461,N_1682,N_1566);
nor U4462 (N_4462,N_101,N_949);
nor U4463 (N_4463,N_560,N_1704);
or U4464 (N_4464,N_1561,N_1927);
nand U4465 (N_4465,N_1338,N_1516);
nand U4466 (N_4466,N_1019,N_768);
and U4467 (N_4467,N_2438,N_2128);
nor U4468 (N_4468,N_1944,N_1002);
and U4469 (N_4469,N_210,N_1407);
and U4470 (N_4470,N_455,N_1460);
and U4471 (N_4471,N_2437,N_2395);
nor U4472 (N_4472,N_370,N_1759);
nor U4473 (N_4473,N_507,N_1059);
nand U4474 (N_4474,N_1480,N_967);
and U4475 (N_4475,N_2308,N_30);
and U4476 (N_4476,N_380,N_1518);
nor U4477 (N_4477,N_1952,N_541);
or U4478 (N_4478,N_817,N_1849);
or U4479 (N_4479,N_705,N_1552);
and U4480 (N_4480,N_2482,N_2259);
nor U4481 (N_4481,N_1617,N_1978);
and U4482 (N_4482,N_2304,N_982);
nand U4483 (N_4483,N_560,N_1130);
nor U4484 (N_4484,N_1824,N_1366);
and U4485 (N_4485,N_2183,N_1999);
nor U4486 (N_4486,N_145,N_473);
nand U4487 (N_4487,N_2039,N_2488);
nor U4488 (N_4488,N_600,N_1164);
nand U4489 (N_4489,N_784,N_688);
or U4490 (N_4490,N_2348,N_443);
and U4491 (N_4491,N_1031,N_2353);
and U4492 (N_4492,N_1494,N_44);
or U4493 (N_4493,N_1663,N_2110);
nor U4494 (N_4494,N_2457,N_447);
and U4495 (N_4495,N_188,N_1463);
or U4496 (N_4496,N_2194,N_1970);
nand U4497 (N_4497,N_2414,N_987);
nor U4498 (N_4498,N_1767,N_1448);
or U4499 (N_4499,N_415,N_778);
nand U4500 (N_4500,N_918,N_1836);
and U4501 (N_4501,N_1525,N_1607);
nor U4502 (N_4502,N_613,N_2091);
nand U4503 (N_4503,N_2214,N_1161);
and U4504 (N_4504,N_113,N_1759);
or U4505 (N_4505,N_2127,N_51);
or U4506 (N_4506,N_2138,N_2477);
nand U4507 (N_4507,N_319,N_92);
nand U4508 (N_4508,N_1763,N_1219);
nand U4509 (N_4509,N_1449,N_1477);
nand U4510 (N_4510,N_981,N_369);
nor U4511 (N_4511,N_300,N_2087);
and U4512 (N_4512,N_1258,N_462);
nor U4513 (N_4513,N_1062,N_491);
and U4514 (N_4514,N_1095,N_1537);
and U4515 (N_4515,N_1720,N_1236);
nand U4516 (N_4516,N_210,N_981);
and U4517 (N_4517,N_203,N_2213);
nand U4518 (N_4518,N_433,N_2101);
nor U4519 (N_4519,N_2331,N_1881);
nand U4520 (N_4520,N_2278,N_1262);
or U4521 (N_4521,N_2080,N_2153);
nor U4522 (N_4522,N_1124,N_2030);
nor U4523 (N_4523,N_432,N_1271);
and U4524 (N_4524,N_1781,N_608);
and U4525 (N_4525,N_2302,N_2460);
and U4526 (N_4526,N_2215,N_2229);
nor U4527 (N_4527,N_2311,N_293);
nor U4528 (N_4528,N_2070,N_942);
and U4529 (N_4529,N_1464,N_2055);
nor U4530 (N_4530,N_278,N_2181);
or U4531 (N_4531,N_2176,N_2017);
or U4532 (N_4532,N_2418,N_984);
or U4533 (N_4533,N_2084,N_1998);
or U4534 (N_4534,N_348,N_913);
or U4535 (N_4535,N_2294,N_459);
nor U4536 (N_4536,N_598,N_807);
nor U4537 (N_4537,N_1474,N_115);
and U4538 (N_4538,N_729,N_349);
or U4539 (N_4539,N_990,N_1554);
and U4540 (N_4540,N_1139,N_1042);
or U4541 (N_4541,N_425,N_707);
nand U4542 (N_4542,N_300,N_481);
or U4543 (N_4543,N_2083,N_1022);
nand U4544 (N_4544,N_2326,N_111);
or U4545 (N_4545,N_51,N_2364);
or U4546 (N_4546,N_1424,N_1463);
and U4547 (N_4547,N_1493,N_1413);
nand U4548 (N_4548,N_688,N_1355);
nor U4549 (N_4549,N_1286,N_171);
nor U4550 (N_4550,N_740,N_2223);
xnor U4551 (N_4551,N_80,N_2352);
or U4552 (N_4552,N_231,N_2041);
or U4553 (N_4553,N_846,N_2489);
or U4554 (N_4554,N_1265,N_2385);
nor U4555 (N_4555,N_129,N_514);
and U4556 (N_4556,N_1489,N_781);
nand U4557 (N_4557,N_524,N_1852);
and U4558 (N_4558,N_1034,N_588);
or U4559 (N_4559,N_1952,N_642);
nand U4560 (N_4560,N_1694,N_2209);
nor U4561 (N_4561,N_413,N_2450);
or U4562 (N_4562,N_1416,N_878);
and U4563 (N_4563,N_474,N_7);
nor U4564 (N_4564,N_1641,N_520);
and U4565 (N_4565,N_879,N_2004);
or U4566 (N_4566,N_2147,N_402);
or U4567 (N_4567,N_1747,N_1247);
and U4568 (N_4568,N_650,N_1797);
and U4569 (N_4569,N_850,N_2094);
or U4570 (N_4570,N_1609,N_1388);
or U4571 (N_4571,N_2036,N_443);
and U4572 (N_4572,N_1338,N_501);
nor U4573 (N_4573,N_2157,N_1498);
or U4574 (N_4574,N_1727,N_1656);
or U4575 (N_4575,N_668,N_1306);
and U4576 (N_4576,N_1771,N_1356);
nand U4577 (N_4577,N_504,N_1102);
and U4578 (N_4578,N_365,N_1586);
nand U4579 (N_4579,N_2451,N_850);
or U4580 (N_4580,N_1770,N_1545);
nor U4581 (N_4581,N_1412,N_521);
and U4582 (N_4582,N_626,N_2154);
nand U4583 (N_4583,N_1465,N_1317);
and U4584 (N_4584,N_2146,N_2472);
nand U4585 (N_4585,N_1244,N_47);
nand U4586 (N_4586,N_1005,N_1531);
xnor U4587 (N_4587,N_1402,N_1468);
and U4588 (N_4588,N_2362,N_1155);
and U4589 (N_4589,N_709,N_163);
and U4590 (N_4590,N_982,N_1017);
xnor U4591 (N_4591,N_2416,N_1873);
nor U4592 (N_4592,N_1043,N_1765);
nor U4593 (N_4593,N_2280,N_1435);
and U4594 (N_4594,N_96,N_1812);
and U4595 (N_4595,N_1808,N_1558);
nor U4596 (N_4596,N_761,N_1632);
nand U4597 (N_4597,N_368,N_2258);
and U4598 (N_4598,N_1701,N_613);
and U4599 (N_4599,N_1831,N_2308);
nor U4600 (N_4600,N_2015,N_384);
or U4601 (N_4601,N_1311,N_483);
or U4602 (N_4602,N_2239,N_2095);
and U4603 (N_4603,N_2490,N_1941);
and U4604 (N_4604,N_1013,N_177);
and U4605 (N_4605,N_1841,N_435);
or U4606 (N_4606,N_1756,N_2118);
and U4607 (N_4607,N_1820,N_451);
and U4608 (N_4608,N_2146,N_910);
nand U4609 (N_4609,N_1064,N_1296);
or U4610 (N_4610,N_878,N_58);
nand U4611 (N_4611,N_1851,N_2307);
nand U4612 (N_4612,N_1922,N_938);
nor U4613 (N_4613,N_134,N_2113);
nor U4614 (N_4614,N_1146,N_1105);
or U4615 (N_4615,N_2290,N_2385);
nor U4616 (N_4616,N_1492,N_2287);
or U4617 (N_4617,N_89,N_2158);
nand U4618 (N_4618,N_1743,N_14);
nand U4619 (N_4619,N_900,N_223);
nor U4620 (N_4620,N_952,N_1857);
and U4621 (N_4621,N_1598,N_1115);
and U4622 (N_4622,N_1763,N_2120);
and U4623 (N_4623,N_2045,N_735);
nor U4624 (N_4624,N_1373,N_1423);
or U4625 (N_4625,N_1725,N_1688);
and U4626 (N_4626,N_448,N_483);
or U4627 (N_4627,N_564,N_1063);
nand U4628 (N_4628,N_1440,N_149);
nor U4629 (N_4629,N_579,N_1733);
and U4630 (N_4630,N_2385,N_1088);
or U4631 (N_4631,N_2382,N_805);
nor U4632 (N_4632,N_6,N_1462);
and U4633 (N_4633,N_1430,N_1617);
and U4634 (N_4634,N_1627,N_1546);
nand U4635 (N_4635,N_2470,N_109);
nand U4636 (N_4636,N_523,N_2445);
nand U4637 (N_4637,N_653,N_2098);
nor U4638 (N_4638,N_106,N_2023);
nand U4639 (N_4639,N_2163,N_1195);
nand U4640 (N_4640,N_2056,N_462);
and U4641 (N_4641,N_1094,N_482);
nor U4642 (N_4642,N_1204,N_1646);
nand U4643 (N_4643,N_701,N_2237);
nor U4644 (N_4644,N_1320,N_1142);
nor U4645 (N_4645,N_212,N_165);
nand U4646 (N_4646,N_104,N_567);
nand U4647 (N_4647,N_1873,N_1385);
and U4648 (N_4648,N_1600,N_1417);
or U4649 (N_4649,N_107,N_461);
nand U4650 (N_4650,N_1399,N_2160);
nand U4651 (N_4651,N_1794,N_186);
nand U4652 (N_4652,N_1760,N_1683);
and U4653 (N_4653,N_1714,N_506);
nor U4654 (N_4654,N_329,N_1857);
or U4655 (N_4655,N_1342,N_2218);
and U4656 (N_4656,N_2259,N_749);
nand U4657 (N_4657,N_1720,N_553);
nor U4658 (N_4658,N_2039,N_851);
or U4659 (N_4659,N_608,N_2163);
or U4660 (N_4660,N_2239,N_619);
or U4661 (N_4661,N_1407,N_558);
nand U4662 (N_4662,N_2112,N_446);
nor U4663 (N_4663,N_1944,N_1065);
and U4664 (N_4664,N_918,N_1869);
nand U4665 (N_4665,N_1997,N_2442);
and U4666 (N_4666,N_2426,N_2242);
xnor U4667 (N_4667,N_773,N_906);
and U4668 (N_4668,N_283,N_1085);
and U4669 (N_4669,N_1690,N_739);
nor U4670 (N_4670,N_1193,N_1050);
and U4671 (N_4671,N_1125,N_1590);
nor U4672 (N_4672,N_1185,N_734);
nand U4673 (N_4673,N_77,N_368);
and U4674 (N_4674,N_1992,N_2438);
and U4675 (N_4675,N_2407,N_1442);
and U4676 (N_4676,N_1084,N_1813);
nor U4677 (N_4677,N_560,N_166);
nor U4678 (N_4678,N_2499,N_1110);
or U4679 (N_4679,N_130,N_960);
and U4680 (N_4680,N_2365,N_163);
and U4681 (N_4681,N_735,N_972);
and U4682 (N_4682,N_2204,N_308);
nand U4683 (N_4683,N_1256,N_1410);
and U4684 (N_4684,N_770,N_586);
nand U4685 (N_4685,N_1110,N_1409);
and U4686 (N_4686,N_1760,N_1259);
or U4687 (N_4687,N_284,N_554);
nor U4688 (N_4688,N_1737,N_432);
and U4689 (N_4689,N_163,N_1013);
nor U4690 (N_4690,N_1323,N_990);
or U4691 (N_4691,N_2158,N_880);
nand U4692 (N_4692,N_654,N_819);
or U4693 (N_4693,N_2296,N_146);
or U4694 (N_4694,N_433,N_1499);
nand U4695 (N_4695,N_1170,N_1166);
and U4696 (N_4696,N_1940,N_206);
xor U4697 (N_4697,N_1602,N_650);
or U4698 (N_4698,N_1527,N_1777);
nor U4699 (N_4699,N_253,N_2269);
nand U4700 (N_4700,N_1722,N_2045);
nor U4701 (N_4701,N_1064,N_2205);
xnor U4702 (N_4702,N_1018,N_845);
nand U4703 (N_4703,N_1865,N_1845);
nor U4704 (N_4704,N_2085,N_328);
nand U4705 (N_4705,N_601,N_595);
or U4706 (N_4706,N_630,N_690);
nand U4707 (N_4707,N_15,N_1255);
or U4708 (N_4708,N_1198,N_1370);
and U4709 (N_4709,N_1596,N_445);
nor U4710 (N_4710,N_1395,N_2160);
nor U4711 (N_4711,N_272,N_2497);
or U4712 (N_4712,N_871,N_444);
nand U4713 (N_4713,N_2052,N_1759);
and U4714 (N_4714,N_1169,N_1033);
and U4715 (N_4715,N_1018,N_1504);
and U4716 (N_4716,N_1954,N_305);
or U4717 (N_4717,N_1440,N_549);
or U4718 (N_4718,N_228,N_799);
nor U4719 (N_4719,N_2019,N_2020);
and U4720 (N_4720,N_632,N_1345);
nand U4721 (N_4721,N_2005,N_499);
or U4722 (N_4722,N_2467,N_1620);
or U4723 (N_4723,N_712,N_2256);
xor U4724 (N_4724,N_1997,N_856);
and U4725 (N_4725,N_1743,N_1943);
nand U4726 (N_4726,N_243,N_48);
or U4727 (N_4727,N_1677,N_1789);
or U4728 (N_4728,N_840,N_332);
and U4729 (N_4729,N_689,N_405);
nor U4730 (N_4730,N_2254,N_531);
or U4731 (N_4731,N_1779,N_965);
nor U4732 (N_4732,N_1579,N_1158);
and U4733 (N_4733,N_2423,N_2447);
nand U4734 (N_4734,N_2156,N_920);
or U4735 (N_4735,N_1395,N_1114);
nand U4736 (N_4736,N_1003,N_1806);
or U4737 (N_4737,N_143,N_1983);
and U4738 (N_4738,N_590,N_1641);
nand U4739 (N_4739,N_1196,N_2352);
and U4740 (N_4740,N_2021,N_48);
nand U4741 (N_4741,N_1729,N_1813);
nand U4742 (N_4742,N_24,N_255);
nor U4743 (N_4743,N_2164,N_1426);
and U4744 (N_4744,N_1931,N_2362);
nand U4745 (N_4745,N_2436,N_1046);
and U4746 (N_4746,N_946,N_184);
nor U4747 (N_4747,N_1343,N_469);
or U4748 (N_4748,N_1218,N_1487);
nand U4749 (N_4749,N_1943,N_2346);
nand U4750 (N_4750,N_2172,N_2162);
nand U4751 (N_4751,N_356,N_1366);
and U4752 (N_4752,N_1233,N_1673);
nor U4753 (N_4753,N_2065,N_1834);
and U4754 (N_4754,N_1823,N_1216);
and U4755 (N_4755,N_66,N_958);
nor U4756 (N_4756,N_1315,N_690);
nand U4757 (N_4757,N_1736,N_1847);
nor U4758 (N_4758,N_890,N_453);
or U4759 (N_4759,N_826,N_862);
or U4760 (N_4760,N_451,N_1053);
or U4761 (N_4761,N_1483,N_2491);
and U4762 (N_4762,N_2230,N_2302);
or U4763 (N_4763,N_2244,N_340);
or U4764 (N_4764,N_333,N_233);
nor U4765 (N_4765,N_1011,N_475);
and U4766 (N_4766,N_1344,N_1123);
or U4767 (N_4767,N_694,N_12);
nor U4768 (N_4768,N_86,N_1932);
nor U4769 (N_4769,N_528,N_1618);
nor U4770 (N_4770,N_170,N_16);
nor U4771 (N_4771,N_2050,N_931);
or U4772 (N_4772,N_1165,N_375);
or U4773 (N_4773,N_996,N_548);
or U4774 (N_4774,N_1821,N_2267);
nand U4775 (N_4775,N_2430,N_1836);
nand U4776 (N_4776,N_1580,N_906);
nand U4777 (N_4777,N_1241,N_1125);
nand U4778 (N_4778,N_1271,N_1308);
and U4779 (N_4779,N_875,N_732);
or U4780 (N_4780,N_474,N_2194);
nor U4781 (N_4781,N_2206,N_1142);
nor U4782 (N_4782,N_2338,N_196);
nor U4783 (N_4783,N_2076,N_1148);
or U4784 (N_4784,N_338,N_1479);
xnor U4785 (N_4785,N_1355,N_1846);
nand U4786 (N_4786,N_432,N_916);
nor U4787 (N_4787,N_620,N_1544);
nor U4788 (N_4788,N_1424,N_2415);
nor U4789 (N_4789,N_1348,N_509);
or U4790 (N_4790,N_1694,N_2151);
nor U4791 (N_4791,N_564,N_1133);
nor U4792 (N_4792,N_493,N_104);
nand U4793 (N_4793,N_1735,N_1670);
nor U4794 (N_4794,N_344,N_1486);
or U4795 (N_4795,N_2221,N_2343);
or U4796 (N_4796,N_1116,N_2177);
or U4797 (N_4797,N_1645,N_707);
or U4798 (N_4798,N_2116,N_768);
nand U4799 (N_4799,N_534,N_97);
or U4800 (N_4800,N_1016,N_1432);
nor U4801 (N_4801,N_1115,N_972);
nand U4802 (N_4802,N_492,N_1731);
nor U4803 (N_4803,N_1700,N_382);
or U4804 (N_4804,N_1941,N_1710);
or U4805 (N_4805,N_1917,N_2436);
nand U4806 (N_4806,N_1866,N_2109);
xor U4807 (N_4807,N_493,N_710);
or U4808 (N_4808,N_883,N_1915);
nor U4809 (N_4809,N_601,N_1829);
nor U4810 (N_4810,N_693,N_672);
xnor U4811 (N_4811,N_347,N_785);
nor U4812 (N_4812,N_728,N_100);
nand U4813 (N_4813,N_836,N_2143);
or U4814 (N_4814,N_1344,N_646);
or U4815 (N_4815,N_1875,N_481);
and U4816 (N_4816,N_1232,N_905);
or U4817 (N_4817,N_1162,N_1209);
nand U4818 (N_4818,N_2439,N_641);
and U4819 (N_4819,N_1367,N_78);
or U4820 (N_4820,N_1459,N_195);
and U4821 (N_4821,N_1895,N_1752);
nor U4822 (N_4822,N_621,N_1259);
nand U4823 (N_4823,N_130,N_228);
xor U4824 (N_4824,N_1105,N_1006);
nand U4825 (N_4825,N_2357,N_1650);
and U4826 (N_4826,N_1123,N_1495);
nand U4827 (N_4827,N_339,N_903);
nor U4828 (N_4828,N_1301,N_2122);
nor U4829 (N_4829,N_1584,N_1287);
and U4830 (N_4830,N_1309,N_1415);
and U4831 (N_4831,N_38,N_233);
and U4832 (N_4832,N_1318,N_999);
or U4833 (N_4833,N_2209,N_1348);
and U4834 (N_4834,N_2475,N_1685);
and U4835 (N_4835,N_2196,N_96);
or U4836 (N_4836,N_1660,N_275);
nand U4837 (N_4837,N_1996,N_903);
or U4838 (N_4838,N_2003,N_2316);
or U4839 (N_4839,N_2317,N_484);
nor U4840 (N_4840,N_1251,N_2356);
nand U4841 (N_4841,N_526,N_461);
and U4842 (N_4842,N_577,N_1573);
nand U4843 (N_4843,N_32,N_1540);
or U4844 (N_4844,N_221,N_1302);
nand U4845 (N_4845,N_2258,N_2031);
or U4846 (N_4846,N_1722,N_782);
or U4847 (N_4847,N_217,N_1507);
nor U4848 (N_4848,N_1657,N_1464);
and U4849 (N_4849,N_743,N_309);
or U4850 (N_4850,N_2330,N_1277);
or U4851 (N_4851,N_318,N_2493);
nor U4852 (N_4852,N_1684,N_1750);
nor U4853 (N_4853,N_1991,N_2093);
nand U4854 (N_4854,N_1982,N_1993);
or U4855 (N_4855,N_659,N_612);
nor U4856 (N_4856,N_1565,N_491);
nor U4857 (N_4857,N_1499,N_1786);
or U4858 (N_4858,N_625,N_286);
nand U4859 (N_4859,N_1946,N_1695);
or U4860 (N_4860,N_430,N_1600);
nor U4861 (N_4861,N_957,N_2207);
nand U4862 (N_4862,N_650,N_1442);
or U4863 (N_4863,N_1087,N_1607);
and U4864 (N_4864,N_1500,N_2002);
or U4865 (N_4865,N_764,N_2406);
nand U4866 (N_4866,N_466,N_2142);
nor U4867 (N_4867,N_2140,N_54);
nand U4868 (N_4868,N_1574,N_609);
or U4869 (N_4869,N_1769,N_569);
nor U4870 (N_4870,N_1315,N_1714);
nand U4871 (N_4871,N_2347,N_1380);
or U4872 (N_4872,N_1629,N_1059);
nand U4873 (N_4873,N_1356,N_2235);
nor U4874 (N_4874,N_753,N_754);
and U4875 (N_4875,N_1924,N_1530);
and U4876 (N_4876,N_1482,N_976);
or U4877 (N_4877,N_1490,N_2168);
or U4878 (N_4878,N_2290,N_2262);
nand U4879 (N_4879,N_1071,N_2312);
nor U4880 (N_4880,N_1639,N_1176);
or U4881 (N_4881,N_2355,N_2222);
nand U4882 (N_4882,N_248,N_1049);
nor U4883 (N_4883,N_648,N_994);
nand U4884 (N_4884,N_2310,N_1525);
nor U4885 (N_4885,N_2457,N_2327);
or U4886 (N_4886,N_1097,N_1471);
nor U4887 (N_4887,N_1600,N_414);
nand U4888 (N_4888,N_1357,N_2188);
or U4889 (N_4889,N_255,N_1073);
nand U4890 (N_4890,N_1576,N_1065);
nor U4891 (N_4891,N_1321,N_2460);
or U4892 (N_4892,N_1047,N_1192);
or U4893 (N_4893,N_481,N_1030);
and U4894 (N_4894,N_1748,N_1607);
and U4895 (N_4895,N_2208,N_747);
nor U4896 (N_4896,N_1438,N_1216);
or U4897 (N_4897,N_1042,N_1214);
nand U4898 (N_4898,N_1865,N_560);
nand U4899 (N_4899,N_1158,N_23);
and U4900 (N_4900,N_1377,N_1244);
nor U4901 (N_4901,N_359,N_1267);
or U4902 (N_4902,N_33,N_870);
nand U4903 (N_4903,N_801,N_1853);
nor U4904 (N_4904,N_1705,N_2125);
xnor U4905 (N_4905,N_2446,N_369);
nor U4906 (N_4906,N_2373,N_2052);
or U4907 (N_4907,N_1096,N_1432);
nand U4908 (N_4908,N_1852,N_876);
and U4909 (N_4909,N_110,N_2490);
and U4910 (N_4910,N_217,N_2216);
or U4911 (N_4911,N_2016,N_939);
nor U4912 (N_4912,N_3,N_473);
nand U4913 (N_4913,N_1887,N_65);
nor U4914 (N_4914,N_906,N_86);
or U4915 (N_4915,N_386,N_1731);
or U4916 (N_4916,N_717,N_671);
nand U4917 (N_4917,N_2393,N_2221);
nand U4918 (N_4918,N_914,N_183);
nand U4919 (N_4919,N_821,N_1023);
nand U4920 (N_4920,N_365,N_753);
nand U4921 (N_4921,N_1204,N_2411);
and U4922 (N_4922,N_1378,N_1611);
nand U4923 (N_4923,N_2046,N_1372);
and U4924 (N_4924,N_651,N_694);
nor U4925 (N_4925,N_2421,N_1383);
or U4926 (N_4926,N_603,N_2106);
nor U4927 (N_4927,N_1681,N_878);
nor U4928 (N_4928,N_717,N_1991);
or U4929 (N_4929,N_1959,N_2025);
nor U4930 (N_4930,N_247,N_1697);
nand U4931 (N_4931,N_1479,N_158);
or U4932 (N_4932,N_1471,N_2183);
nor U4933 (N_4933,N_781,N_529);
or U4934 (N_4934,N_292,N_1883);
xor U4935 (N_4935,N_172,N_405);
nand U4936 (N_4936,N_1872,N_565);
or U4937 (N_4937,N_529,N_1606);
or U4938 (N_4938,N_1944,N_524);
nor U4939 (N_4939,N_2207,N_125);
and U4940 (N_4940,N_1828,N_1554);
nor U4941 (N_4941,N_207,N_2369);
nand U4942 (N_4942,N_1970,N_1528);
nor U4943 (N_4943,N_2119,N_69);
nor U4944 (N_4944,N_388,N_940);
or U4945 (N_4945,N_631,N_2421);
and U4946 (N_4946,N_1555,N_1696);
nor U4947 (N_4947,N_1395,N_1699);
and U4948 (N_4948,N_2463,N_2211);
and U4949 (N_4949,N_1959,N_2195);
nand U4950 (N_4950,N_2309,N_2480);
nor U4951 (N_4951,N_2446,N_244);
and U4952 (N_4952,N_1488,N_362);
nand U4953 (N_4953,N_2189,N_1090);
nor U4954 (N_4954,N_2102,N_25);
or U4955 (N_4955,N_565,N_128);
nor U4956 (N_4956,N_1204,N_375);
nand U4957 (N_4957,N_1716,N_681);
or U4958 (N_4958,N_1041,N_2477);
and U4959 (N_4959,N_108,N_2034);
nand U4960 (N_4960,N_1735,N_2408);
and U4961 (N_4961,N_1472,N_2250);
xnor U4962 (N_4962,N_719,N_215);
nor U4963 (N_4963,N_2225,N_2388);
or U4964 (N_4964,N_1312,N_1619);
or U4965 (N_4965,N_1750,N_1863);
or U4966 (N_4966,N_911,N_2305);
nand U4967 (N_4967,N_551,N_268);
and U4968 (N_4968,N_1613,N_990);
or U4969 (N_4969,N_457,N_1569);
nand U4970 (N_4970,N_2317,N_1348);
nand U4971 (N_4971,N_2032,N_1862);
nand U4972 (N_4972,N_1949,N_1095);
nor U4973 (N_4973,N_1213,N_239);
and U4974 (N_4974,N_1131,N_798);
nor U4975 (N_4975,N_2262,N_1067);
nor U4976 (N_4976,N_1917,N_1927);
nor U4977 (N_4977,N_1773,N_1378);
and U4978 (N_4978,N_723,N_1988);
or U4979 (N_4979,N_1509,N_326);
and U4980 (N_4980,N_364,N_1181);
nand U4981 (N_4981,N_2419,N_325);
and U4982 (N_4982,N_629,N_1889);
nand U4983 (N_4983,N_1052,N_498);
and U4984 (N_4984,N_591,N_212);
nand U4985 (N_4985,N_316,N_2231);
nor U4986 (N_4986,N_1872,N_2048);
nand U4987 (N_4987,N_1376,N_1703);
and U4988 (N_4988,N_62,N_320);
nand U4989 (N_4989,N_1608,N_1901);
and U4990 (N_4990,N_1669,N_1616);
nand U4991 (N_4991,N_1015,N_1409);
nor U4992 (N_4992,N_1301,N_786);
nor U4993 (N_4993,N_1550,N_1779);
and U4994 (N_4994,N_1665,N_1759);
and U4995 (N_4995,N_1410,N_927);
nor U4996 (N_4996,N_1317,N_960);
nor U4997 (N_4997,N_887,N_1601);
and U4998 (N_4998,N_40,N_283);
and U4999 (N_4999,N_674,N_228);
and U5000 (N_5000,N_4707,N_3333);
or U5001 (N_5001,N_3331,N_4068);
nand U5002 (N_5002,N_4118,N_4503);
nor U5003 (N_5003,N_3217,N_4005);
nor U5004 (N_5004,N_3542,N_4139);
nor U5005 (N_5005,N_4859,N_3341);
nand U5006 (N_5006,N_4288,N_4823);
and U5007 (N_5007,N_4750,N_3149);
nor U5008 (N_5008,N_3844,N_3252);
nand U5009 (N_5009,N_2815,N_3439);
and U5010 (N_5010,N_3609,N_2915);
nor U5011 (N_5011,N_3226,N_4210);
or U5012 (N_5012,N_2828,N_4484);
nor U5013 (N_5013,N_2698,N_2773);
and U5014 (N_5014,N_4390,N_2971);
and U5015 (N_5015,N_3288,N_3811);
and U5016 (N_5016,N_4405,N_4975);
nand U5017 (N_5017,N_4386,N_3781);
nand U5018 (N_5018,N_4836,N_3214);
and U5019 (N_5019,N_3045,N_3472);
and U5020 (N_5020,N_3236,N_3995);
or U5021 (N_5021,N_3962,N_2977);
and U5022 (N_5022,N_3353,N_4282);
nand U5023 (N_5023,N_2673,N_4896);
nand U5024 (N_5024,N_4154,N_3795);
and U5025 (N_5025,N_4211,N_3038);
nor U5026 (N_5026,N_4334,N_4170);
and U5027 (N_5027,N_3643,N_3603);
or U5028 (N_5028,N_2502,N_3167);
and U5029 (N_5029,N_4027,N_4119);
or U5030 (N_5030,N_4042,N_3782);
or U5031 (N_5031,N_2694,N_4374);
nand U5032 (N_5032,N_3227,N_3517);
or U5033 (N_5033,N_2941,N_3201);
nand U5034 (N_5034,N_3897,N_3507);
nand U5035 (N_5035,N_4554,N_4489);
nor U5036 (N_5036,N_3604,N_2604);
or U5037 (N_5037,N_3810,N_3522);
nand U5038 (N_5038,N_4192,N_3230);
nor U5039 (N_5039,N_4522,N_4654);
and U5040 (N_5040,N_3898,N_4592);
nor U5041 (N_5041,N_3835,N_4011);
nand U5042 (N_5042,N_4748,N_4081);
or U5043 (N_5043,N_4728,N_4495);
nand U5044 (N_5044,N_3303,N_4837);
and U5045 (N_5045,N_3481,N_4983);
and U5046 (N_5046,N_3723,N_4356);
nor U5047 (N_5047,N_3705,N_2758);
and U5048 (N_5048,N_3212,N_4642);
and U5049 (N_5049,N_3516,N_4796);
nand U5050 (N_5050,N_3524,N_3202);
and U5051 (N_5051,N_2998,N_3399);
and U5052 (N_5052,N_4772,N_4371);
nor U5053 (N_5053,N_2591,N_4057);
nand U5054 (N_5054,N_4219,N_3368);
nor U5055 (N_5055,N_3185,N_3686);
or U5056 (N_5056,N_3939,N_4150);
and U5057 (N_5057,N_3878,N_2609);
nor U5058 (N_5058,N_4074,N_4652);
nor U5059 (N_5059,N_4215,N_3678);
nor U5060 (N_5060,N_2830,N_3848);
nor U5061 (N_5061,N_3461,N_2857);
or U5062 (N_5062,N_4569,N_2532);
nor U5063 (N_5063,N_3042,N_4218);
or U5064 (N_5064,N_4603,N_3283);
nor U5065 (N_5065,N_3463,N_4263);
or U5066 (N_5066,N_3793,N_2631);
nor U5067 (N_5067,N_3944,N_2702);
and U5068 (N_5068,N_3390,N_4014);
or U5069 (N_5069,N_4292,N_3457);
or U5070 (N_5070,N_2798,N_4309);
nand U5071 (N_5071,N_4962,N_3145);
and U5072 (N_5072,N_4391,N_2782);
or U5073 (N_5073,N_3946,N_3605);
or U5074 (N_5074,N_4037,N_4467);
nor U5075 (N_5075,N_4621,N_3616);
or U5076 (N_5076,N_4440,N_4879);
nand U5077 (N_5077,N_4771,N_4166);
and U5078 (N_5078,N_3757,N_3111);
and U5079 (N_5079,N_4141,N_4075);
nand U5080 (N_5080,N_4528,N_3961);
nand U5081 (N_5081,N_3891,N_4559);
nor U5082 (N_5082,N_4945,N_2903);
nor U5083 (N_5083,N_2512,N_4612);
and U5084 (N_5084,N_3969,N_4903);
and U5085 (N_5085,N_3278,N_4913);
nor U5086 (N_5086,N_3363,N_4850);
nor U5087 (N_5087,N_3446,N_3486);
nor U5088 (N_5088,N_2564,N_4167);
nor U5089 (N_5089,N_3165,N_3398);
and U5090 (N_5090,N_2671,N_2685);
and U5091 (N_5091,N_3385,N_3137);
and U5092 (N_5092,N_4753,N_2660);
nand U5093 (N_5093,N_4846,N_2797);
nor U5094 (N_5094,N_4711,N_2722);
nand U5095 (N_5095,N_3578,N_2668);
and U5096 (N_5096,N_3139,N_4350);
or U5097 (N_5097,N_2736,N_3647);
and U5098 (N_5098,N_4110,N_4313);
or U5099 (N_5099,N_4449,N_4638);
and U5100 (N_5100,N_3450,N_2642);
nor U5101 (N_5101,N_3365,N_4636);
nor U5102 (N_5102,N_4957,N_3014);
or U5103 (N_5103,N_4464,N_2728);
and U5104 (N_5104,N_4687,N_4841);
nand U5105 (N_5105,N_4947,N_3364);
xor U5106 (N_5106,N_4804,N_3220);
or U5107 (N_5107,N_4583,N_3753);
nand U5108 (N_5108,N_4774,N_3340);
nor U5109 (N_5109,N_3631,N_2901);
or U5110 (N_5110,N_4257,N_3701);
nand U5111 (N_5111,N_2672,N_4000);
nor U5112 (N_5112,N_3970,N_3788);
nand U5113 (N_5113,N_2839,N_4778);
and U5114 (N_5114,N_3455,N_3071);
or U5115 (N_5115,N_3211,N_3965);
and U5116 (N_5116,N_2602,N_2827);
or U5117 (N_5117,N_3979,N_3142);
or U5118 (N_5118,N_3445,N_3180);
or U5119 (N_5119,N_2813,N_4286);
nand U5120 (N_5120,N_4819,N_3689);
and U5121 (N_5121,N_4889,N_3648);
or U5122 (N_5122,N_4053,N_3594);
and U5123 (N_5123,N_4199,N_4222);
or U5124 (N_5124,N_2619,N_3242);
and U5125 (N_5125,N_2536,N_3294);
or U5126 (N_5126,N_3460,N_3092);
nand U5127 (N_5127,N_3050,N_2877);
nor U5128 (N_5128,N_2554,N_2675);
or U5129 (N_5129,N_3987,N_4754);
nand U5130 (N_5130,N_3411,N_3200);
or U5131 (N_5131,N_2772,N_4546);
nand U5132 (N_5132,N_2973,N_4773);
or U5133 (N_5133,N_3598,N_3095);
or U5134 (N_5134,N_4744,N_2939);
nand U5135 (N_5135,N_3482,N_3816);
nand U5136 (N_5136,N_4404,N_3651);
and U5137 (N_5137,N_3478,N_3624);
nand U5138 (N_5138,N_2691,N_2885);
and U5139 (N_5139,N_4996,N_4157);
nor U5140 (N_5140,N_3090,N_3556);
nand U5141 (N_5141,N_4809,N_4646);
or U5142 (N_5142,N_4954,N_4409);
or U5143 (N_5143,N_2718,N_4240);
xnor U5144 (N_5144,N_3821,N_3727);
or U5145 (N_5145,N_4269,N_4106);
and U5146 (N_5146,N_2795,N_4377);
and U5147 (N_5147,N_3162,N_3641);
nor U5148 (N_5148,N_2820,N_3915);
and U5149 (N_5149,N_3527,N_2834);
nor U5150 (N_5150,N_3345,N_2683);
nand U5151 (N_5151,N_2754,N_3859);
nor U5152 (N_5152,N_3001,N_4358);
and U5153 (N_5153,N_3775,N_2542);
and U5154 (N_5154,N_3102,N_2819);
and U5155 (N_5155,N_3151,N_3058);
nand U5156 (N_5156,N_4426,N_3983);
nor U5157 (N_5157,N_3313,N_4320);
nor U5158 (N_5158,N_4419,N_2897);
nor U5159 (N_5159,N_3442,N_2909);
nor U5160 (N_5160,N_3925,N_3657);
or U5161 (N_5161,N_4331,N_2553);
or U5162 (N_5162,N_3825,N_3144);
nand U5163 (N_5163,N_3082,N_3739);
nand U5164 (N_5164,N_3218,N_2561);
nand U5165 (N_5165,N_2555,N_4822);
and U5166 (N_5166,N_3259,N_4010);
nor U5167 (N_5167,N_4738,N_3763);
and U5168 (N_5168,N_2812,N_3312);
or U5169 (N_5169,N_4985,N_4415);
or U5170 (N_5170,N_2509,N_2572);
or U5171 (N_5171,N_4740,N_2558);
and U5172 (N_5172,N_4630,N_2986);
nand U5173 (N_5173,N_3376,N_3510);
nor U5174 (N_5174,N_4930,N_4665);
and U5175 (N_5175,N_3459,N_4152);
nand U5176 (N_5176,N_2898,N_3555);
nor U5177 (N_5177,N_3026,N_4697);
nor U5178 (N_5178,N_4710,N_3113);
or U5179 (N_5179,N_4884,N_4732);
and U5180 (N_5180,N_4557,N_3491);
nand U5181 (N_5181,N_3266,N_4212);
or U5182 (N_5182,N_4452,N_3537);
nand U5183 (N_5183,N_3855,N_2521);
or U5184 (N_5184,N_4311,N_4741);
nand U5185 (N_5185,N_4626,N_3830);
and U5186 (N_5186,N_2988,N_2711);
and U5187 (N_5187,N_3468,N_4757);
nor U5188 (N_5188,N_4226,N_3749);
and U5189 (N_5189,N_3268,N_4022);
and U5190 (N_5190,N_3662,N_3762);
nand U5191 (N_5191,N_3140,N_3628);
or U5192 (N_5192,N_3130,N_3083);
or U5193 (N_5193,N_4712,N_4927);
nand U5194 (N_5194,N_3154,N_4049);
nand U5195 (N_5195,N_4287,N_3941);
or U5196 (N_5196,N_3543,N_2684);
nand U5197 (N_5197,N_3632,N_3447);
nand U5198 (N_5198,N_3564,N_2927);
and U5199 (N_5199,N_4656,N_4560);
nor U5200 (N_5200,N_4545,N_2992);
and U5201 (N_5201,N_4971,N_4101);
nor U5202 (N_5202,N_3208,N_4759);
or U5203 (N_5203,N_4250,N_3438);
nor U5204 (N_5204,N_4802,N_4629);
nand U5205 (N_5205,N_4297,N_2716);
and U5206 (N_5206,N_3231,N_3356);
and U5207 (N_5207,N_3237,N_2662);
and U5208 (N_5208,N_4535,N_4285);
and U5209 (N_5209,N_4907,N_2551);
or U5210 (N_5210,N_3867,N_3526);
and U5211 (N_5211,N_4003,N_4379);
and U5212 (N_5212,N_2507,N_4591);
or U5213 (N_5213,N_3173,N_4653);
and U5214 (N_5214,N_4742,N_4127);
nor U5215 (N_5215,N_3794,N_4004);
and U5216 (N_5216,N_4843,N_2814);
or U5217 (N_5217,N_3721,N_4031);
or U5218 (N_5218,N_2636,N_4949);
or U5219 (N_5219,N_2771,N_4082);
nor U5220 (N_5220,N_3694,N_4190);
or U5221 (N_5221,N_3136,N_4335);
nor U5222 (N_5222,N_4733,N_3204);
or U5223 (N_5223,N_4264,N_3474);
and U5224 (N_5224,N_4259,N_3471);
nand U5225 (N_5225,N_3467,N_2535);
or U5226 (N_5226,N_2779,N_3067);
or U5227 (N_5227,N_2862,N_4091);
or U5228 (N_5228,N_2818,N_4716);
or U5229 (N_5229,N_4100,N_3415);
and U5230 (N_5230,N_4186,N_3930);
nand U5231 (N_5231,N_2578,N_2981);
or U5232 (N_5232,N_4084,N_2732);
and U5233 (N_5233,N_4805,N_3016);
nor U5234 (N_5234,N_3298,N_4709);
or U5235 (N_5235,N_3518,N_4800);
and U5236 (N_5236,N_4487,N_2679);
nor U5237 (N_5237,N_4129,N_3325);
nor U5238 (N_5238,N_3973,N_4970);
nor U5239 (N_5239,N_2664,N_3697);
or U5240 (N_5240,N_3525,N_3942);
and U5241 (N_5241,N_4359,N_4046);
and U5242 (N_5242,N_4465,N_2737);
xor U5243 (N_5243,N_4238,N_3738);
and U5244 (N_5244,N_2518,N_4956);
nor U5245 (N_5245,N_3956,N_3704);
and U5246 (N_5246,N_3464,N_2968);
nor U5247 (N_5247,N_3258,N_2606);
nand U5248 (N_5248,N_3778,N_3311);
nand U5249 (N_5249,N_3671,N_3406);
or U5250 (N_5250,N_3361,N_4851);
and U5251 (N_5251,N_3837,N_3745);
and U5252 (N_5252,N_2517,N_4734);
nand U5253 (N_5253,N_3244,N_4811);
and U5254 (N_5254,N_3501,N_3017);
nand U5255 (N_5255,N_4013,N_3764);
nand U5256 (N_5256,N_3620,N_2822);
nor U5257 (N_5257,N_3346,N_4981);
or U5258 (N_5258,N_4087,N_3229);
nor U5259 (N_5259,N_4008,N_3735);
nor U5260 (N_5260,N_3125,N_3074);
nor U5261 (N_5261,N_4873,N_3172);
nand U5262 (N_5262,N_3819,N_3344);
or U5263 (N_5263,N_4516,N_4848);
or U5264 (N_5264,N_4727,N_3621);
and U5265 (N_5265,N_4389,N_3256);
or U5266 (N_5266,N_2719,N_3622);
or U5267 (N_5267,N_2928,N_3886);
or U5268 (N_5268,N_4904,N_3393);
xor U5269 (N_5269,N_3053,N_3748);
or U5270 (N_5270,N_3269,N_3724);
and U5271 (N_5271,N_4078,N_4015);
nand U5272 (N_5272,N_2610,N_4891);
and U5273 (N_5273,N_4149,N_3563);
nor U5274 (N_5274,N_4195,N_3077);
or U5275 (N_5275,N_3696,N_3339);
and U5276 (N_5276,N_4136,N_2816);
or U5277 (N_5277,N_3908,N_2868);
nor U5278 (N_5278,N_3008,N_4530);
nor U5279 (N_5279,N_4790,N_4617);
xor U5280 (N_5280,N_3126,N_4348);
and U5281 (N_5281,N_2787,N_4887);
nand U5282 (N_5282,N_3558,N_3655);
nor U5283 (N_5283,N_4911,N_3530);
or U5284 (N_5284,N_3998,N_4067);
nor U5285 (N_5285,N_4310,N_3098);
nand U5286 (N_5286,N_3384,N_2666);
nor U5287 (N_5287,N_4420,N_4402);
nand U5288 (N_5288,N_3840,N_2759);
nor U5289 (N_5289,N_2891,N_3660);
and U5290 (N_5290,N_4121,N_3533);
xor U5291 (N_5291,N_4436,N_3932);
nand U5292 (N_5292,N_3011,N_3146);
or U5293 (N_5293,N_4980,N_4797);
nand U5294 (N_5294,N_3550,N_4724);
or U5295 (N_5295,N_4604,N_4547);
nand U5296 (N_5296,N_2991,N_3466);
and U5297 (N_5297,N_4073,N_2661);
nand U5298 (N_5298,N_2692,N_3424);
nand U5299 (N_5299,N_3338,N_4302);
nor U5300 (N_5300,N_4095,N_4897);
and U5301 (N_5301,N_3366,N_4613);
nand U5302 (N_5302,N_4135,N_3685);
and U5303 (N_5303,N_4399,N_2665);
xor U5304 (N_5304,N_4381,N_4161);
nand U5305 (N_5305,N_3473,N_4993);
and U5306 (N_5306,N_4541,N_3304);
nor U5307 (N_5307,N_3565,N_3302);
or U5308 (N_5308,N_2714,N_4050);
or U5309 (N_5309,N_4729,N_2628);
or U5310 (N_5310,N_2693,N_4555);
nand U5311 (N_5311,N_3263,N_4360);
nand U5312 (N_5312,N_4673,N_2725);
and U5313 (N_5313,N_2888,N_3186);
or U5314 (N_5314,N_4023,N_4853);
nand U5315 (N_5315,N_4726,N_3693);
and U5316 (N_5316,N_2566,N_3037);
and U5317 (N_5317,N_3640,N_3433);
nand U5318 (N_5318,N_3034,N_3881);
or U5319 (N_5319,N_4434,N_4574);
nor U5320 (N_5320,N_4698,N_3907);
and U5321 (N_5321,N_2794,N_3726);
or U5322 (N_5322,N_2529,N_3076);
and U5323 (N_5323,N_4585,N_2763);
nand U5324 (N_5324,N_4179,N_4478);
or U5325 (N_5325,N_3465,N_4977);
and U5326 (N_5326,N_4885,N_2644);
nor U5327 (N_5327,N_3271,N_3926);
nor U5328 (N_5328,N_3275,N_3408);
and U5329 (N_5329,N_4628,N_3870);
nand U5330 (N_5330,N_4538,N_4725);
nand U5331 (N_5331,N_4433,N_2570);
nor U5332 (N_5332,N_4382,N_3319);
and U5333 (N_5333,N_3645,N_4364);
nor U5334 (N_5334,N_3423,N_3427);
or U5335 (N_5335,N_3536,N_3470);
or U5336 (N_5336,N_4755,N_3495);
or U5337 (N_5337,N_4156,N_3375);
and U5338 (N_5338,N_4443,N_4083);
and U5339 (N_5339,N_3358,N_4735);
nand U5340 (N_5340,N_4984,N_4342);
and U5341 (N_5341,N_2710,N_3695);
and U5342 (N_5342,N_4045,N_2634);
or U5343 (N_5343,N_2522,N_4283);
nor U5344 (N_5344,N_2639,N_4827);
or U5345 (N_5345,N_2588,N_4459);
or U5346 (N_5346,N_3255,N_4634);
or U5347 (N_5347,N_3857,N_2645);
or U5348 (N_5348,N_4942,N_3958);
and U5349 (N_5349,N_4163,N_3232);
and U5350 (N_5350,N_2520,N_4648);
nor U5351 (N_5351,N_4306,N_3751);
nor U5352 (N_5352,N_2584,N_3197);
nor U5353 (N_5353,N_2984,N_4806);
nor U5354 (N_5354,N_4052,N_3044);
and U5355 (N_5355,N_4563,N_4953);
and U5356 (N_5356,N_4810,N_2846);
and U5357 (N_5357,N_4312,N_4908);
nor U5358 (N_5358,N_4565,N_4507);
nand U5359 (N_5359,N_3822,N_3260);
nor U5360 (N_5360,N_3623,N_3119);
nand U5361 (N_5361,N_4245,N_2743);
and U5362 (N_5362,N_3206,N_3318);
nand U5363 (N_5363,N_3078,N_3086);
nand U5364 (N_5364,N_3910,N_4122);
nor U5365 (N_5365,N_3952,N_2844);
or U5366 (N_5366,N_4036,N_4808);
or U5367 (N_5367,N_3843,N_3216);
nor U5368 (N_5368,N_2937,N_4854);
nor U5369 (N_5369,N_4833,N_4609);
nor U5370 (N_5370,N_3354,N_3213);
nand U5371 (N_5371,N_4221,N_3625);
nand U5372 (N_5372,N_2617,N_4883);
nor U5373 (N_5373,N_3948,N_4357);
or U5374 (N_5374,N_3571,N_3971);
nand U5375 (N_5375,N_3093,N_3813);
or U5376 (N_5376,N_3006,N_2687);
nand U5377 (N_5377,N_3722,N_4517);
and U5378 (N_5378,N_3324,N_4303);
or U5379 (N_5379,N_4909,N_3383);
nand U5380 (N_5380,N_3513,N_4227);
or U5381 (N_5381,N_4279,N_4779);
nor U5382 (N_5382,N_3613,N_2859);
nor U5383 (N_5383,N_3959,N_4474);
or U5384 (N_5384,N_2576,N_3317);
and U5385 (N_5385,N_4147,N_4940);
nand U5386 (N_5386,N_3733,N_3496);
nor U5387 (N_5387,N_4544,N_4183);
or U5388 (N_5388,N_4088,N_3326);
and U5389 (N_5389,N_3322,N_3574);
nand U5390 (N_5390,N_3305,N_3182);
or U5391 (N_5391,N_4300,N_3039);
nor U5392 (N_5392,N_2573,N_4761);
or U5393 (N_5393,N_3316,N_3520);
or U5394 (N_5394,N_2921,N_2525);
or U5395 (N_5395,N_3417,N_2781);
and U5396 (N_5396,N_3426,N_3994);
nor U5397 (N_5397,N_4793,N_3619);
nand U5398 (N_5398,N_3777,N_4069);
nand U5399 (N_5399,N_3239,N_4328);
or U5400 (N_5400,N_3179,N_3335);
and U5401 (N_5401,N_4966,N_4339);
nor U5402 (N_5402,N_3360,N_2893);
nand U5403 (N_5403,N_2889,N_3947);
nor U5404 (N_5404,N_4995,N_3276);
nor U5405 (N_5405,N_2530,N_3847);
nand U5406 (N_5406,N_3924,N_3249);
and U5407 (N_5407,N_3688,N_2600);
and U5408 (N_5408,N_4830,N_3002);
or U5409 (N_5409,N_4989,N_4616);
nor U5410 (N_5410,N_2976,N_4463);
or U5411 (N_5411,N_3935,N_4316);
nand U5412 (N_5412,N_4214,N_3561);
or U5413 (N_5413,N_4644,N_3401);
nand U5414 (N_5414,N_3487,N_4886);
nor U5415 (N_5415,N_4573,N_4160);
and U5416 (N_5416,N_3416,N_3892);
nor U5417 (N_5417,N_2817,N_4182);
nand U5418 (N_5418,N_4025,N_4140);
nor U5419 (N_5419,N_3434,N_4699);
or U5420 (N_5420,N_3453,N_2966);
nor U5421 (N_5421,N_4817,N_3673);
or U5422 (N_5422,N_4718,N_2552);
and U5423 (N_5423,N_3989,N_2999);
nor U5424 (N_5424,N_4345,N_4441);
and U5425 (N_5425,N_4587,N_3035);
and U5426 (N_5426,N_3668,N_3754);
and U5427 (N_5427,N_2805,N_4184);
and U5428 (N_5428,N_3418,N_4553);
nand U5429 (N_5429,N_3786,N_2641);
nand U5430 (N_5430,N_4237,N_3192);
nand U5431 (N_5431,N_3658,N_2808);
nand U5432 (N_5432,N_3681,N_3676);
and U5433 (N_5433,N_3065,N_4632);
or U5434 (N_5434,N_3589,N_3707);
and U5435 (N_5435,N_2880,N_4066);
nor U5436 (N_5436,N_3388,N_4020);
nand U5437 (N_5437,N_3240,N_4143);
nand U5438 (N_5438,N_2824,N_3976);
or U5439 (N_5439,N_4667,N_2919);
or U5440 (N_5440,N_4151,N_4787);
nor U5441 (N_5441,N_2648,N_2592);
and U5442 (N_5442,N_4447,N_2646);
and U5443 (N_5443,N_4708,N_2733);
nand U5444 (N_5444,N_3797,N_3400);
nand U5445 (N_5445,N_3798,N_3854);
and U5446 (N_5446,N_3118,N_3927);
and U5447 (N_5447,N_4960,N_4691);
nand U5448 (N_5448,N_3858,N_4905);
nor U5449 (N_5449,N_3716,N_4874);
nand U5450 (N_5450,N_3068,N_3646);
and U5451 (N_5451,N_4562,N_4427);
and U5452 (N_5452,N_3123,N_4469);
nand U5453 (N_5453,N_3503,N_4398);
and U5454 (N_5454,N_3792,N_4839);
or U5455 (N_5455,N_3287,N_3320);
or U5456 (N_5456,N_2842,N_3802);
nor U5457 (N_5457,N_3051,N_4798);
and U5458 (N_5458,N_2930,N_2560);
or U5459 (N_5459,N_4207,N_3055);
nand U5460 (N_5460,N_2949,N_3024);
or U5461 (N_5461,N_4470,N_3337);
and U5462 (N_5462,N_4281,N_3277);
nand U5463 (N_5463,N_3549,N_4935);
nor U5464 (N_5464,N_2829,N_3048);
nor U5465 (N_5465,N_3394,N_4571);
nor U5466 (N_5466,N_3490,N_3099);
nand U5467 (N_5467,N_4177,N_4675);
or U5468 (N_5468,N_2938,N_3159);
or U5469 (N_5469,N_4035,N_3284);
or U5470 (N_5470,N_4365,N_3209);
nor U5471 (N_5471,N_2882,N_4992);
nand U5472 (N_5472,N_4533,N_2950);
or U5473 (N_5473,N_4900,N_3851);
and U5474 (N_5474,N_2583,N_4120);
nand U5475 (N_5475,N_4175,N_4070);
nor U5476 (N_5476,N_3022,N_4747);
or U5477 (N_5477,N_4669,N_4499);
nand U5478 (N_5478,N_3535,N_2659);
nor U5479 (N_5479,N_3634,N_3968);
or U5480 (N_5480,N_4138,N_4422);
nor U5481 (N_5481,N_4209,N_3814);
nand U5482 (N_5482,N_4006,N_2550);
nand U5483 (N_5483,N_4265,N_4987);
nand U5484 (N_5484,N_4397,N_3156);
and U5485 (N_5485,N_4230,N_2935);
and U5486 (N_5486,N_4700,N_4526);
or U5487 (N_5487,N_4875,N_4829);
and U5488 (N_5488,N_4137,N_3904);
nor U5489 (N_5489,N_4431,N_4531);
nand U5490 (N_5490,N_4527,N_2802);
nand U5491 (N_5491,N_4882,N_4291);
or U5492 (N_5492,N_3504,N_2845);
nand U5493 (N_5493,N_2653,N_3581);
or U5494 (N_5494,N_4668,N_4171);
and U5495 (N_5495,N_3766,N_3483);
or U5496 (N_5496,N_3462,N_4736);
and U5497 (N_5497,N_4028,N_4655);
nand U5498 (N_5498,N_3755,N_2537);
or U5499 (N_5499,N_3128,N_4169);
and U5500 (N_5500,N_4633,N_3062);
and U5501 (N_5501,N_2780,N_4089);
or U5502 (N_5502,N_3015,N_3018);
and U5503 (N_5503,N_3148,N_3860);
nor U5504 (N_5504,N_4588,N_3667);
nand U5505 (N_5505,N_3307,N_3991);
nor U5506 (N_5506,N_3692,N_2739);
or U5507 (N_5507,N_3272,N_3432);
and U5508 (N_5508,N_4155,N_2593);
nor U5509 (N_5509,N_3759,N_4417);
or U5510 (N_5510,N_2686,N_2669);
nor U5511 (N_5511,N_4248,N_2546);
and U5512 (N_5512,N_3253,N_4485);
or U5513 (N_5513,N_4657,N_3548);
nand U5514 (N_5514,N_2690,N_3920);
and U5515 (N_5515,N_4769,N_3141);
nand U5516 (N_5516,N_4739,N_2982);
nand U5517 (N_5517,N_3131,N_3043);
or U5518 (N_5518,N_2703,N_4615);
and U5519 (N_5519,N_2744,N_3984);
nand U5520 (N_5520,N_4094,N_4505);
nor U5521 (N_5521,N_4363,N_4564);
nand U5522 (N_5522,N_4959,N_4967);
nand U5523 (N_5523,N_4717,N_4205);
or U5524 (N_5524,N_3274,N_2740);
nand U5525 (N_5525,N_2916,N_3025);
and U5526 (N_5526,N_4719,N_4314);
or U5527 (N_5527,N_4509,N_4329);
nor U5528 (N_5528,N_4601,N_4520);
or U5529 (N_5529,N_4792,N_4099);
nor U5530 (N_5530,N_3444,N_2674);
and U5531 (N_5531,N_4702,N_3712);
nor U5532 (N_5532,N_3725,N_3404);
or U5533 (N_5533,N_2841,N_3552);
and U5534 (N_5534,N_4430,N_4387);
or U5535 (N_5535,N_3257,N_4494);
and U5536 (N_5536,N_4353,N_4918);
and U5537 (N_5537,N_2720,N_3291);
nand U5538 (N_5538,N_3582,N_4228);
nand U5539 (N_5539,N_2958,N_3484);
nand U5540 (N_5540,N_3347,N_3033);
and U5541 (N_5541,N_3590,N_4721);
nor U5542 (N_5542,N_4552,N_4033);
or U5543 (N_5543,N_4111,N_4385);
and U5544 (N_5544,N_4946,N_4939);
or U5545 (N_5545,N_3152,N_4361);
and U5546 (N_5546,N_3744,N_4519);
or U5547 (N_5547,N_3937,N_3732);
nor U5548 (N_5548,N_3396,N_3772);
nor U5549 (N_5549,N_2562,N_4685);
and U5550 (N_5550,N_4428,N_2515);
or U5551 (N_5551,N_3449,N_3081);
and U5552 (N_5552,N_3718,N_4868);
or U5553 (N_5553,N_2623,N_4450);
and U5554 (N_5554,N_4229,N_4115);
nor U5555 (N_5555,N_4176,N_3163);
nor U5556 (N_5556,N_4344,N_3817);
nand U5557 (N_5557,N_2647,N_4631);
nand U5558 (N_5558,N_4307,N_3703);
and U5559 (N_5559,N_4932,N_4479);
or U5560 (N_5560,N_4737,N_3349);
or U5561 (N_5561,N_3297,N_3183);
nor U5562 (N_5562,N_3719,N_2678);
nor U5563 (N_5563,N_4340,N_4758);
or U5564 (N_5564,N_3711,N_4117);
or U5565 (N_5565,N_3780,N_2980);
or U5566 (N_5566,N_2849,N_2920);
nand U5567 (N_5567,N_4187,N_3873);
nand U5568 (N_5568,N_3280,N_3760);
nand U5569 (N_5569,N_3012,N_2734);
or U5570 (N_5570,N_3729,N_3378);
nand U5571 (N_5571,N_4295,N_2832);
and U5572 (N_5572,N_3120,N_4937);
nand U5573 (N_5573,N_2757,N_3529);
or U5574 (N_5574,N_4369,N_4534);
and U5575 (N_5575,N_4408,N_4493);
nand U5576 (N_5576,N_3425,N_2954);
or U5577 (N_5577,N_3833,N_2590);
nand U5578 (N_5578,N_4392,N_4109);
and U5579 (N_5579,N_4341,N_2967);
nor U5580 (N_5580,N_4610,N_3429);
nand U5581 (N_5581,N_3084,N_2585);
and U5582 (N_5582,N_3007,N_3664);
xnor U5583 (N_5583,N_4595,N_3541);
or U5584 (N_5584,N_2985,N_3710);
and U5585 (N_5585,N_4506,N_4424);
and U5586 (N_5586,N_4326,N_3523);
and U5587 (N_5587,N_2848,N_2931);
nor U5588 (N_5588,N_4097,N_3502);
nor U5589 (N_5589,N_2775,N_3579);
or U5590 (N_5590,N_2946,N_3642);
nand U5591 (N_5591,N_4866,N_3829);
nor U5592 (N_5592,N_2975,N_3853);
nor U5593 (N_5593,N_2870,N_4188);
or U5594 (N_5594,N_3273,N_4130);
and U5595 (N_5595,N_4255,N_2911);
nand U5596 (N_5596,N_4203,N_3699);
or U5597 (N_5597,N_2777,N_2696);
and U5598 (N_5598,N_4777,N_2682);
or U5599 (N_5599,N_4007,N_4435);
nand U5600 (N_5600,N_3838,N_3586);
nor U5601 (N_5601,N_2622,N_4383);
and U5602 (N_5602,N_4123,N_3666);
nand U5603 (N_5603,N_4941,N_3734);
nand U5604 (N_5604,N_3403,N_3181);
nand U5605 (N_5605,N_4860,N_4041);
nor U5606 (N_5606,N_3412,N_2516);
and U5607 (N_5607,N_3852,N_4931);
nor U5608 (N_5608,N_4418,N_3567);
and U5609 (N_5609,N_3799,N_3607);
nand U5610 (N_5610,N_3557,N_4498);
nand U5611 (N_5611,N_3804,N_3477);
and U5612 (N_5612,N_2869,N_4062);
nand U5613 (N_5613,N_4556,N_3031);
nor U5614 (N_5614,N_3009,N_3189);
or U5615 (N_5615,N_3215,N_2705);
or U5616 (N_5616,N_4146,N_3355);
or U5617 (N_5617,N_4421,N_4680);
or U5618 (N_5618,N_2799,N_2633);
and U5619 (N_5619,N_4425,N_4396);
or U5620 (N_5620,N_4677,N_2603);
or U5621 (N_5621,N_2594,N_4597);
and U5622 (N_5622,N_2756,N_4400);
or U5623 (N_5623,N_4745,N_3769);
nand U5624 (N_5624,N_3949,N_2810);
nor U5625 (N_5625,N_3367,N_4521);
and U5626 (N_5626,N_4635,N_4423);
or U5627 (N_5627,N_3289,N_2534);
nor U5628 (N_5628,N_4325,N_4814);
nor U5629 (N_5629,N_3972,N_4902);
nand U5630 (N_5630,N_3221,N_2707);
nand U5631 (N_5631,N_4704,N_2618);
nor U5632 (N_5632,N_3414,N_4124);
nand U5633 (N_5633,N_3437,N_4262);
nor U5634 (N_5634,N_3115,N_3663);
nor U5635 (N_5635,N_3485,N_3789);
and U5636 (N_5636,N_2762,N_2786);
and U5637 (N_5637,N_3615,N_3992);
and U5638 (N_5638,N_3104,N_4780);
or U5639 (N_5639,N_2863,N_2879);
or U5640 (N_5640,N_4164,N_3234);
or U5641 (N_5641,N_3911,N_2883);
nand U5642 (N_5642,N_2676,N_3448);
and U5643 (N_5643,N_3514,N_4542);
nand U5644 (N_5644,N_4767,N_4686);
or U5645 (N_5645,N_3633,N_4304);
nand U5646 (N_5646,N_4267,N_4202);
and U5647 (N_5647,N_3841,N_2970);
and U5648 (N_5648,N_3545,N_3306);
and U5649 (N_5649,N_3559,N_3836);
or U5650 (N_5650,N_3177,N_4153);
or U5651 (N_5651,N_2587,N_3454);
nor U5652 (N_5652,N_4678,N_3175);
or U5653 (N_5653,N_4413,N_2783);
and U5654 (N_5654,N_4965,N_3982);
and U5655 (N_5655,N_4271,N_2789);
and U5656 (N_5656,N_4643,N_3912);
nand U5657 (N_5657,N_4454,N_3951);
and U5658 (N_5658,N_2785,N_4789);
nand U5659 (N_5659,N_4086,N_3877);
nand U5660 (N_5660,N_4162,N_4486);
and U5661 (N_5661,N_2574,N_4076);
and U5662 (N_5662,N_4690,N_3923);
and U5663 (N_5663,N_3166,N_2944);
or U5664 (N_5664,N_4990,N_2727);
nand U5665 (N_5665,N_3945,N_3301);
nor U5666 (N_5666,N_2729,N_2544);
nand U5667 (N_5667,N_4864,N_3964);
nor U5668 (N_5668,N_4722,N_3489);
and U5669 (N_5669,N_4622,N_4114);
nor U5670 (N_5670,N_3428,N_4579);
or U5671 (N_5671,N_3135,N_4844);
xnor U5672 (N_5672,N_3895,N_2549);
nor U5673 (N_5673,N_2917,N_2792);
or U5674 (N_5674,N_3413,N_3094);
and U5675 (N_5675,N_2922,N_2955);
nor U5676 (N_5676,N_3121,N_2663);
or U5677 (N_5677,N_2764,N_3379);
or U5678 (N_5678,N_2526,N_4071);
or U5679 (N_5679,N_3334,N_2580);
or U5680 (N_5680,N_3943,N_4093);
or U5681 (N_5681,N_2625,N_3861);
nor U5682 (N_5682,N_3874,N_3903);
nor U5683 (N_5683,N_2539,N_3776);
nand U5684 (N_5684,N_3713,N_4598);
or U5685 (N_5685,N_2960,N_4200);
and U5686 (N_5686,N_3295,N_3790);
nor U5687 (N_5687,N_3246,N_2627);
or U5688 (N_5688,N_4969,N_4445);
nand U5689 (N_5689,N_2508,N_4826);
nor U5690 (N_5690,N_2541,N_3381);
nor U5691 (N_5691,N_2831,N_2987);
and U5692 (N_5692,N_2996,N_2709);
nor U5693 (N_5693,N_2599,N_2708);
and U5694 (N_5694,N_3219,N_3824);
nor U5695 (N_5695,N_3611,N_2918);
and U5696 (N_5696,N_4232,N_4032);
or U5697 (N_5697,N_3100,N_3767);
or U5698 (N_5698,N_2867,N_4103);
nor U5699 (N_5699,N_3850,N_2905);
nor U5700 (N_5700,N_4372,N_4671);
or U5701 (N_5701,N_4529,N_4590);
and U5702 (N_5702,N_3988,N_4705);
and U5703 (N_5703,N_3885,N_3410);
or U5704 (N_5704,N_4784,N_4349);
nor U5705 (N_5705,N_3382,N_2567);
nor U5706 (N_5706,N_4395,N_4979);
or U5707 (N_5707,N_4549,N_2565);
nor U5708 (N_5708,N_2504,N_2910);
nor U5709 (N_5709,N_4749,N_4786);
nor U5710 (N_5710,N_4606,N_2978);
nand U5711 (N_5711,N_3612,N_4001);
nor U5712 (N_5712,N_4012,N_4038);
or U5713 (N_5713,N_2776,N_2531);
nand U5714 (N_5714,N_3057,N_4266);
or U5715 (N_5715,N_4842,N_3430);
nand U5716 (N_5716,N_2929,N_4246);
and U5717 (N_5717,N_2959,N_3352);
nand U5718 (N_5718,N_2855,N_4764);
nand U5719 (N_5719,N_3863,N_3940);
xnor U5720 (N_5720,N_3309,N_4943);
or U5721 (N_5721,N_3188,N_2962);
and U5722 (N_5722,N_3884,N_4414);
nor U5723 (N_5723,N_3540,N_4060);
nor U5724 (N_5724,N_4296,N_3362);
nand U5725 (N_5725,N_4788,N_3980);
or U5726 (N_5726,N_2895,N_2706);
nand U5727 (N_5727,N_4327,N_3019);
and U5728 (N_5728,N_4384,N_4504);
or U5729 (N_5729,N_4664,N_4224);
or U5730 (N_5730,N_4696,N_4694);
or U5731 (N_5731,N_4333,N_4714);
nor U5732 (N_5732,N_2865,N_3127);
and U5733 (N_5733,N_3110,N_2677);
or U5734 (N_5734,N_2899,N_3730);
or U5735 (N_5735,N_4444,N_4058);
or U5736 (N_5736,N_2796,N_2864);
or U5737 (N_5737,N_3199,N_4783);
nand U5738 (N_5738,N_4437,N_3158);
nand U5739 (N_5739,N_3521,N_2701);
or U5740 (N_5740,N_4775,N_4021);
or U5741 (N_5741,N_3900,N_3476);
xnor U5742 (N_5742,N_4756,N_3636);
and U5743 (N_5743,N_3265,N_3807);
or U5744 (N_5744,N_3882,N_3812);
nand U5745 (N_5745,N_4432,N_2924);
nor U5746 (N_5746,N_3512,N_4838);
nand U5747 (N_5747,N_4513,N_4950);
and U5748 (N_5748,N_3369,N_3061);
nand U5749 (N_5749,N_3653,N_3027);
and U5750 (N_5750,N_3004,N_4670);
and U5751 (N_5751,N_2932,N_4659);
nand U5752 (N_5752,N_3922,N_3405);
nor U5753 (N_5753,N_3876,N_3771);
nand U5754 (N_5754,N_4584,N_3103);
and U5755 (N_5755,N_4388,N_4986);
or U5756 (N_5756,N_4952,N_4540);
nand U5757 (N_5757,N_4193,N_4862);
or U5758 (N_5758,N_3828,N_2767);
nor U5759 (N_5759,N_3279,N_4496);
nand U5760 (N_5760,N_4178,N_4926);
nand U5761 (N_5761,N_4581,N_2638);
and U5762 (N_5762,N_3153,N_2774);
or U5763 (N_5763,N_4511,N_4551);
nand U5764 (N_5764,N_2934,N_4925);
nand U5765 (N_5765,N_2563,N_3440);
or U5766 (N_5766,N_4477,N_3750);
nand U5767 (N_5767,N_4048,N_4920);
or U5768 (N_5768,N_3389,N_3741);
or U5769 (N_5769,N_4145,N_2993);
nand U5770 (N_5770,N_4849,N_2712);
and U5771 (N_5771,N_4064,N_2747);
and U5772 (N_5772,N_3570,N_3546);
or U5773 (N_5773,N_2836,N_2942);
nand U5774 (N_5774,N_4799,N_3030);
and U5775 (N_5775,N_3469,N_2741);
nand U5776 (N_5776,N_3087,N_4801);
nand U5777 (N_5777,N_4040,N_2913);
and U5778 (N_5778,N_4856,N_4651);
or U5779 (N_5779,N_3372,N_4888);
nor U5780 (N_5780,N_3373,N_3282);
nor U5781 (N_5781,N_4834,N_4301);
xnor U5782 (N_5782,N_4252,N_2629);
nand U5783 (N_5783,N_3106,N_4321);
nor U5784 (N_5784,N_2607,N_4611);
and U5785 (N_5785,N_3665,N_3842);
or U5786 (N_5786,N_3190,N_4895);
xnor U5787 (N_5787,N_4092,N_3005);
and U5788 (N_5788,N_4890,N_4254);
and U5789 (N_5789,N_4869,N_4059);
and U5790 (N_5790,N_4490,N_4274);
nand U5791 (N_5791,N_3993,N_2995);
nor U5792 (N_5792,N_3241,N_4276);
and U5793 (N_5793,N_4198,N_4208);
or U5794 (N_5794,N_3672,N_4104);
or U5795 (N_5795,N_4508,N_3999);
and U5796 (N_5796,N_4679,N_4912);
nor U5797 (N_5797,N_3868,N_2688);
or U5798 (N_5798,N_4871,N_3108);
and U5799 (N_5799,N_3602,N_4994);
nor U5800 (N_5800,N_3117,N_4568);
nor U5801 (N_5801,N_2699,N_3056);
nor U5802 (N_5802,N_4855,N_3089);
or U5803 (N_5803,N_2871,N_4337);
nand U5804 (N_5804,N_4144,N_3953);
nand U5805 (N_5805,N_4770,N_3914);
nand U5806 (N_5806,N_2760,N_4180);
nand U5807 (N_5807,N_4236,N_4376);
and U5808 (N_5808,N_4457,N_4647);
and U5809 (N_5809,N_2878,N_2801);
nor U5810 (N_5810,N_3889,N_2731);
and U5811 (N_5811,N_4065,N_4821);
nor U5812 (N_5812,N_4963,N_3436);
nor U5813 (N_5813,N_2697,N_2596);
and U5814 (N_5814,N_2964,N_3905);
nand U5815 (N_5815,N_4116,N_2569);
or U5816 (N_5816,N_4991,N_3890);
and U5817 (N_5817,N_4277,N_4352);
nand U5818 (N_5818,N_4275,N_3592);
nand U5819 (N_5819,N_3917,N_4305);
and U5820 (N_5820,N_4936,N_2748);
nor U5821 (N_5821,N_4133,N_4401);
nand U5822 (N_5822,N_4523,N_2953);
and U5823 (N_5823,N_2577,N_4131);
nor U5824 (N_5824,N_3342,N_3330);
or U5825 (N_5825,N_3133,N_2904);
nor U5826 (N_5826,N_2614,N_4923);
nand U5827 (N_5827,N_2784,N_2853);
and U5828 (N_5828,N_4235,N_3032);
nand U5829 (N_5829,N_2652,N_4330);
nand U5830 (N_5830,N_2809,N_2689);
nand U5831 (N_5831,N_4047,N_2974);
or U5832 (N_5832,N_3974,N_2632);
nor U5833 (N_5833,N_2601,N_2543);
nand U5834 (N_5834,N_4867,N_3610);
nand U5835 (N_5835,N_3500,N_3452);
nor U5836 (N_5836,N_4148,N_4763);
nor U5837 (N_5837,N_4666,N_3114);
xnor U5838 (N_5838,N_3515,N_3680);
and U5839 (N_5839,N_4901,N_3332);
nand U5840 (N_5840,N_4492,N_3743);
and U5841 (N_5841,N_2626,N_2533);
nand U5842 (N_5842,N_4650,N_2527);
and U5843 (N_5843,N_2838,N_3562);
nand U5844 (N_5844,N_3419,N_3866);
nor U5845 (N_5845,N_3746,N_4054);
nor U5846 (N_5846,N_2506,N_3661);
nand U5847 (N_5847,N_4543,N_4410);
nor U5848 (N_5848,N_4475,N_3245);
nand U5849 (N_5849,N_3553,N_4407);
or U5850 (N_5850,N_4623,N_3787);
nand U5851 (N_5851,N_2874,N_4378);
nand U5852 (N_5852,N_4550,N_4857);
nand U5853 (N_5853,N_4766,N_3402);
or U5854 (N_5854,N_3264,N_4225);
or U5855 (N_5855,N_4009,N_2956);
nor U5856 (N_5856,N_3371,N_2961);
or U5857 (N_5857,N_4825,N_2713);
or U5858 (N_5858,N_4701,N_3737);
or U5859 (N_5859,N_3768,N_3551);
nor U5860 (N_5860,N_4958,N_4916);
and U5861 (N_5861,N_2548,N_3649);
and U5862 (N_5862,N_4730,N_4289);
nor U5863 (N_5863,N_3706,N_4416);
and U5864 (N_5864,N_2751,N_3285);
and U5865 (N_5865,N_2940,N_2788);
nand U5866 (N_5866,N_2902,N_4524);
nand U5867 (N_5867,N_3205,N_3899);
or U5868 (N_5868,N_3097,N_4355);
nor U5869 (N_5869,N_3687,N_3800);
or U5870 (N_5870,N_4290,N_4997);
nand U5871 (N_5871,N_2742,N_3534);
and U5872 (N_5872,N_3101,N_2519);
and U5873 (N_5873,N_3064,N_4688);
nand U5874 (N_5874,N_4865,N_3872);
and U5875 (N_5875,N_2650,N_4599);
nor U5876 (N_5876,N_3116,N_4512);
nor U5877 (N_5877,N_2914,N_4840);
nor U5878 (N_5878,N_3674,N_4938);
xnor U5879 (N_5879,N_4640,N_4863);
or U5880 (N_5880,N_2840,N_2948);
nor U5881 (N_5881,N_3519,N_4815);
or U5882 (N_5882,N_3629,N_3171);
and U5883 (N_5883,N_3323,N_4968);
nand U5884 (N_5884,N_3293,N_3528);
nor U5885 (N_5885,N_4765,N_4204);
or U5886 (N_5886,N_4582,N_4816);
nor U5887 (N_5887,N_3286,N_4572);
nand U5888 (N_5888,N_3576,N_3329);
nand U5889 (N_5889,N_3169,N_2825);
nor U5890 (N_5890,N_4315,N_3931);
nand U5891 (N_5891,N_2540,N_3587);
nor U5892 (N_5892,N_3879,N_4723);
or U5893 (N_5893,N_4620,N_4852);
and U5894 (N_5894,N_3174,N_3747);
and U5895 (N_5895,N_3784,N_4105);
or U5896 (N_5896,N_2851,N_4466);
and U5897 (N_5897,N_4596,N_3421);
nand U5898 (N_5898,N_2616,N_3235);
or U5899 (N_5899,N_4280,N_3107);
nand U5900 (N_5900,N_3773,N_4298);
nand U5901 (N_5901,N_4713,N_4446);
nand U5902 (N_5902,N_3985,N_4126);
and U5903 (N_5903,N_4681,N_2597);
and U5904 (N_5904,N_4558,N_2575);
nand U5905 (N_5905,N_2556,N_4593);
nor U5906 (N_5906,N_4090,N_2804);
nor U5907 (N_5907,N_2768,N_4605);
nand U5908 (N_5908,N_2876,N_4172);
or U5909 (N_5909,N_4343,N_4881);
nor U5910 (N_5910,N_3488,N_2791);
and U5911 (N_5911,N_4548,N_4168);
nand U5912 (N_5912,N_4539,N_3267);
or U5913 (N_5913,N_4270,N_3635);
nor U5914 (N_5914,N_2952,N_4063);
or U5915 (N_5915,N_4308,N_3690);
nor U5916 (N_5916,N_3990,N_4108);
nand U5917 (N_5917,N_2651,N_2852);
or U5918 (N_5918,N_4898,N_4928);
or U5919 (N_5919,N_3028,N_4017);
nor U5920 (N_5920,N_3717,N_3299);
or U5921 (N_5921,N_4256,N_4791);
and U5922 (N_5922,N_2538,N_4034);
nor U5923 (N_5923,N_4536,N_3374);
nand U5924 (N_5924,N_3088,N_4044);
or U5925 (N_5925,N_3222,N_2843);
or U5926 (N_5926,N_3679,N_3250);
and U5927 (N_5927,N_2680,N_4768);
nor U5928 (N_5928,N_3370,N_3596);
and U5929 (N_5929,N_3492,N_3963);
nor U5930 (N_5930,N_3731,N_4955);
and U5931 (N_5931,N_3498,N_4244);
and U5932 (N_5932,N_3864,N_4973);
nor U5933 (N_5933,N_4649,N_2621);
nand U5934 (N_5934,N_4812,N_2866);
nand U5935 (N_5935,N_3933,N_3950);
nor U5936 (N_5936,N_2500,N_4284);
or U5937 (N_5937,N_4016,N_3742);
nand U5938 (N_5938,N_3617,N_4861);
and U5939 (N_5939,N_3682,N_4368);
nor U5940 (N_5940,N_3584,N_2806);
and U5941 (N_5941,N_4072,N_3262);
nand U5942 (N_5942,N_3168,N_3203);
and U5943 (N_5943,N_3702,N_4429);
and U5944 (N_5944,N_2700,N_4442);
nor U5945 (N_5945,N_3310,N_3010);
nor U5946 (N_5946,N_3134,N_4061);
or U5947 (N_5947,N_3124,N_4501);
xnor U5948 (N_5948,N_4107,N_2847);
nor U5949 (N_5949,N_3547,N_3572);
nand U5950 (N_5950,N_3072,N_2667);
and U5951 (N_5951,N_3066,N_2730);
and U5952 (N_5952,N_4249,N_4951);
and U5953 (N_5953,N_3357,N_4319);
nor U5954 (N_5954,N_3435,N_4915);
nand U5955 (N_5955,N_2649,N_4518);
and U5956 (N_5956,N_3443,N_4600);
and U5957 (N_5957,N_2951,N_4056);
nand U5958 (N_5958,N_3109,N_4658);
nor U5959 (N_5959,N_3736,N_3573);
nand U5960 (N_5960,N_4231,N_4914);
and U5961 (N_5961,N_3779,N_3314);
nand U5962 (N_5962,N_4488,N_3296);
nor U5963 (N_5963,N_3575,N_3047);
nor U5964 (N_5964,N_2510,N_2835);
nor U5965 (N_5965,N_2887,N_4043);
or U5966 (N_5966,N_2800,N_2908);
and U5967 (N_5967,N_3997,N_3902);
nand U5968 (N_5968,N_3233,N_2559);
nor U5969 (N_5969,N_2643,N_3112);
or U5970 (N_5970,N_2715,N_4661);
nor U5971 (N_5971,N_4362,N_4336);
nor U5972 (N_5972,N_3913,N_2630);
nand U5973 (N_5973,N_3928,N_3013);
nor U5974 (N_5974,N_4835,N_2969);
and U5975 (N_5975,N_3261,N_3063);
or U5976 (N_5976,N_3938,N_2881);
and U5977 (N_5977,N_4858,N_4367);
or U5978 (N_5978,N_3327,N_4242);
or U5979 (N_5979,N_4934,N_4448);
nor U5980 (N_5980,N_4299,N_4972);
nor U5981 (N_5981,N_2807,N_2793);
and U5982 (N_5982,N_3281,N_4338);
nor U5983 (N_5983,N_3650,N_3627);
or U5984 (N_5984,N_2611,N_3506);
nor U5985 (N_5985,N_4917,N_4619);
and U5986 (N_5986,N_4332,N_3129);
nor U5987 (N_5987,N_2695,N_2595);
and U5988 (N_5988,N_3036,N_2613);
and U5989 (N_5989,N_3160,N_2620);
or U5990 (N_5990,N_2505,N_3409);
and U5991 (N_5991,N_4351,N_4174);
nor U5992 (N_5992,N_4234,N_3184);
nor U5993 (N_5993,N_2811,N_4406);
and U5994 (N_5994,N_4051,N_4999);
nand U5995 (N_5995,N_4039,N_3975);
and U5996 (N_5996,N_4468,N_3321);
nor U5997 (N_5997,N_3196,N_2860);
and U5998 (N_5998,N_2581,N_4085);
or U5999 (N_5999,N_2511,N_4683);
nand U6000 (N_6000,N_4618,N_4002);
nand U6001 (N_6001,N_4273,N_4831);
or U6002 (N_6002,N_2528,N_3883);
or U6003 (N_6003,N_3608,N_3637);
nor U6004 (N_6004,N_3023,N_4878);
or U6005 (N_6005,N_4580,N_4803);
or U6006 (N_6006,N_3887,N_3756);
nand U6007 (N_6007,N_3654,N_3977);
nor U6008 (N_6008,N_4899,N_4813);
or U6009 (N_6009,N_4055,N_4743);
and U6010 (N_6010,N_2557,N_3880);
nand U6011 (N_6011,N_4393,N_3194);
and U6012 (N_6012,N_2738,N_3380);
and U6013 (N_6013,N_3493,N_4514);
or U6014 (N_6014,N_2586,N_3343);
and U6015 (N_6015,N_2933,N_3052);
and U6016 (N_6016,N_4253,N_3967);
nand U6017 (N_6017,N_4323,N_2884);
nor U6018 (N_6018,N_3957,N_2726);
and U6019 (N_6019,N_3785,N_4480);
and U6020 (N_6020,N_3720,N_3511);
nor U6021 (N_6021,N_3906,N_2735);
nand U6022 (N_6022,N_3079,N_2826);
or U6023 (N_6023,N_4876,N_3187);
or U6024 (N_6024,N_3597,N_3041);
and U6025 (N_6025,N_3532,N_2655);
and U6026 (N_6026,N_3919,N_3300);
or U6027 (N_6027,N_3069,N_3803);
or U6028 (N_6028,N_3508,N_4196);
or U6029 (N_6029,N_3308,N_2723);
nand U6030 (N_6030,N_3138,N_2745);
and U6031 (N_6031,N_4578,N_3238);
and U6032 (N_6032,N_2890,N_4159);
nor U6033 (N_6033,N_3801,N_4471);
nand U6034 (N_6034,N_4201,N_4260);
or U6035 (N_6035,N_3080,N_3909);
or U6036 (N_6036,N_4019,N_4988);
nor U6037 (N_6037,N_3591,N_3808);
or U6038 (N_6038,N_4029,N_2605);
and U6039 (N_6039,N_2983,N_2925);
nand U6040 (N_6040,N_3805,N_4497);
and U6041 (N_6041,N_3585,N_4906);
nand U6042 (N_6042,N_4894,N_3936);
nand U6043 (N_6043,N_3865,N_4322);
and U6044 (N_6044,N_4026,N_4278);
nand U6045 (N_6045,N_4451,N_2778);
and U6046 (N_6046,N_4317,N_4241);
and U6047 (N_6047,N_4380,N_3839);
nor U6048 (N_6048,N_3630,N_2637);
nor U6049 (N_6049,N_4785,N_4347);
nor U6050 (N_6050,N_3155,N_4537);
nand U6051 (N_6051,N_4272,N_4872);
xnor U6052 (N_6052,N_3386,N_4460);
nand U6053 (N_6053,N_3105,N_4746);
nand U6054 (N_6054,N_3228,N_3669);
and U6055 (N_6055,N_4525,N_3774);
and U6056 (N_6056,N_4216,N_3207);
nor U6057 (N_6057,N_2752,N_2770);
nor U6058 (N_6058,N_2945,N_4870);
or U6059 (N_6059,N_2717,N_3251);
and U6060 (N_6060,N_3740,N_4403);
nand U6061 (N_6061,N_4239,N_2746);
and U6062 (N_6062,N_3600,N_4412);
nor U6063 (N_6063,N_4929,N_2579);
nand U6064 (N_6064,N_4820,N_4824);
and U6065 (N_6065,N_4191,N_4532);
or U6066 (N_6066,N_2656,N_2640);
xnor U6067 (N_6067,N_4324,N_4510);
nor U6068 (N_6068,N_4924,N_3350);
and U6069 (N_6069,N_3195,N_4692);
and U6070 (N_6070,N_3638,N_4194);
nand U6071 (N_6071,N_3918,N_2912);
nor U6072 (N_6072,N_4933,N_3765);
or U6073 (N_6073,N_4577,N_3652);
and U6074 (N_6074,N_3715,N_3888);
or U6075 (N_6075,N_2936,N_3176);
or U6076 (N_6076,N_2523,N_3040);
nand U6077 (N_6077,N_4624,N_2545);
nand U6078 (N_6078,N_2994,N_4411);
nor U6079 (N_6079,N_3796,N_3480);
and U6080 (N_6080,N_4370,N_4461);
nand U6081 (N_6081,N_2750,N_3351);
nand U6082 (N_6082,N_2907,N_3456);
nor U6083 (N_6083,N_3708,N_2501);
nor U6084 (N_6084,N_3392,N_3675);
nor U6085 (N_6085,N_3896,N_3986);
nor U6086 (N_6086,N_2972,N_4354);
or U6087 (N_6087,N_3003,N_4258);
nor U6088 (N_6088,N_4079,N_3191);
and U6089 (N_6089,N_3599,N_3588);
nand U6090 (N_6090,N_2582,N_2906);
or U6091 (N_6091,N_2753,N_3420);
nor U6092 (N_6092,N_2571,N_3916);
nand U6093 (N_6093,N_4181,N_3544);
nand U6094 (N_6094,N_4976,N_4080);
nand U6095 (N_6095,N_3070,N_3770);
or U6096 (N_6096,N_3831,N_4268);
and U6097 (N_6097,N_3451,N_4102);
or U6098 (N_6098,N_4567,N_3966);
or U6099 (N_6099,N_3820,N_3560);
nand U6100 (N_6100,N_2821,N_4481);
nor U6101 (N_6101,N_3431,N_4660);
nor U6102 (N_6102,N_4438,N_4462);
or U6103 (N_6103,N_3150,N_3315);
and U6104 (N_6104,N_3809,N_3210);
nor U6105 (N_6105,N_4394,N_3849);
and U6106 (N_6106,N_4500,N_4919);
nand U6107 (N_6107,N_4128,N_4776);
nand U6108 (N_6108,N_3397,N_3059);
nor U6109 (N_6109,N_3791,N_3761);
or U6110 (N_6110,N_2612,N_3714);
nor U6111 (N_6111,N_3247,N_3387);
nor U6112 (N_6112,N_3921,N_4828);
and U6113 (N_6113,N_4627,N_2524);
or U6114 (N_6114,N_4223,N_2681);
or U6115 (N_6115,N_3224,N_3458);
nand U6116 (N_6116,N_4158,N_3684);
and U6117 (N_6117,N_2886,N_2769);
or U6118 (N_6118,N_3554,N_3531);
and U6119 (N_6119,N_4575,N_3270);
nand U6120 (N_6120,N_4961,N_4456);
nand U6121 (N_6121,N_2873,N_2979);
nand U6122 (N_6122,N_2850,N_2654);
and U6123 (N_6123,N_2837,N_3292);
and U6124 (N_6124,N_4751,N_4561);
nor U6125 (N_6125,N_4672,N_4832);
and U6126 (N_6126,N_4220,N_4978);
or U6127 (N_6127,N_3060,N_4476);
nor U6128 (N_6128,N_3046,N_3170);
and U6129 (N_6129,N_4142,N_3815);
nand U6130 (N_6130,N_3096,N_3569);
and U6131 (N_6131,N_4847,N_3020);
or U6132 (N_6132,N_4782,N_4455);
nand U6133 (N_6133,N_3049,N_4173);
nand U6134 (N_6134,N_4112,N_3479);
and U6135 (N_6135,N_3075,N_2965);
and U6136 (N_6136,N_4645,N_4641);
xor U6137 (N_6137,N_3871,N_3254);
nand U6138 (N_6138,N_3132,N_3593);
nor U6139 (N_6139,N_2749,N_3021);
or U6140 (N_6140,N_3700,N_4693);
and U6141 (N_6141,N_3856,N_2861);
or U6142 (N_6142,N_3670,N_4373);
or U6143 (N_6143,N_3290,N_4794);
or U6144 (N_6144,N_4662,N_4637);
or U6145 (N_6145,N_4213,N_3639);
and U6146 (N_6146,N_2947,N_3538);
and U6147 (N_6147,N_2658,N_3580);
nor U6148 (N_6148,N_2598,N_3834);
nand U6149 (N_6149,N_3198,N_4570);
nor U6150 (N_6150,N_4720,N_4247);
and U6151 (N_6151,N_3996,N_4458);
or U6152 (N_6152,N_2990,N_2926);
and U6153 (N_6153,N_3243,N_4892);
or U6154 (N_6154,N_2963,N_2589);
or U6155 (N_6155,N_2608,N_3601);
nand U6156 (N_6156,N_2513,N_3806);
and U6157 (N_6157,N_4682,N_3223);
nor U6158 (N_6158,N_4251,N_3677);
and U6159 (N_6159,N_3348,N_2790);
nand U6160 (N_6160,N_3336,N_3614);
or U6161 (N_6161,N_2704,N_3606);
nor U6162 (N_6162,N_4132,N_3497);
and U6163 (N_6163,N_4944,N_4921);
nor U6164 (N_6164,N_3164,N_4217);
or U6165 (N_6165,N_2514,N_4261);
nor U6166 (N_6166,N_4795,N_3441);
nand U6167 (N_6167,N_3475,N_3509);
or U6168 (N_6168,N_4845,N_3085);
and U6169 (N_6169,N_4910,N_3143);
or U6170 (N_6170,N_4233,N_3029);
nor U6171 (N_6171,N_2615,N_2833);
nor U6172 (N_6172,N_3328,N_3539);
nor U6173 (N_6173,N_2755,N_3893);
nor U6174 (N_6174,N_3618,N_2875);
or U6175 (N_6175,N_4096,N_4243);
or U6176 (N_6176,N_3499,N_4974);
nand U6177 (N_6177,N_4453,N_3494);
nand U6178 (N_6178,N_2957,N_3955);
nand U6179 (N_6179,N_3626,N_2854);
nand U6180 (N_6180,N_4482,N_4502);
nand U6181 (N_6181,N_4030,N_3054);
and U6182 (N_6182,N_3193,N_3758);
nor U6183 (N_6183,N_3698,N_3073);
nand U6184 (N_6184,N_3377,N_3818);
or U6185 (N_6185,N_3823,N_3846);
or U6186 (N_6186,N_4472,N_3783);
nand U6187 (N_6187,N_3869,N_4674);
nand U6188 (N_6188,N_3728,N_4715);
or U6189 (N_6189,N_4602,N_4752);
nor U6190 (N_6190,N_4614,N_4293);
and U6191 (N_6191,N_3875,N_4589);
or U6192 (N_6192,N_4964,N_2997);
xor U6193 (N_6193,N_3568,N_4922);
and U6194 (N_6194,N_4689,N_4684);
or U6195 (N_6195,N_2923,N_4189);
or U6196 (N_6196,N_3752,N_4731);
nand U6197 (N_6197,N_2894,N_4375);
nand U6198 (N_6198,N_3901,N_3978);
nor U6199 (N_6199,N_2724,N_4781);
or U6200 (N_6200,N_3391,N_3359);
nor U6201 (N_6201,N_2766,N_2765);
nor U6202 (N_6202,N_4366,N_2823);
nor U6203 (N_6203,N_2568,N_3826);
nor U6204 (N_6204,N_3656,N_2900);
nor U6205 (N_6205,N_4948,N_4594);
nor U6206 (N_6206,N_3178,N_4893);
nand U6207 (N_6207,N_2547,N_4318);
and U6208 (N_6208,N_4608,N_2896);
nor U6209 (N_6209,N_4024,N_3395);
and U6210 (N_6210,N_3845,N_4880);
or U6211 (N_6211,N_3862,N_2803);
nor U6212 (N_6212,N_4165,N_2761);
and U6213 (N_6213,N_4586,N_4676);
and U6214 (N_6214,N_3583,N_4473);
and U6215 (N_6215,N_4491,N_4134);
and U6216 (N_6216,N_4113,N_3122);
and U6217 (N_6217,N_4515,N_3827);
nand U6218 (N_6218,N_4077,N_4760);
nand U6219 (N_6219,N_2721,N_4018);
nand U6220 (N_6220,N_3832,N_3659);
and U6221 (N_6221,N_3566,N_2503);
nand U6222 (N_6222,N_3147,N_3157);
and U6223 (N_6223,N_2670,N_4807);
and U6224 (N_6224,N_3225,N_4762);
and U6225 (N_6225,N_4982,N_2657);
or U6226 (N_6226,N_3248,N_4625);
nor U6227 (N_6227,N_4185,N_3422);
or U6228 (N_6228,N_3161,N_2624);
or U6229 (N_6229,N_2635,N_4663);
and U6230 (N_6230,N_3691,N_2872);
nor U6231 (N_6231,N_4294,N_4439);
or U6232 (N_6232,N_2892,N_4818);
and U6233 (N_6233,N_4998,N_4098);
and U6234 (N_6234,N_3644,N_3505);
nand U6235 (N_6235,N_4706,N_3981);
nand U6236 (N_6236,N_2856,N_4197);
nand U6237 (N_6237,N_3407,N_4607);
or U6238 (N_6238,N_2989,N_3709);
nand U6239 (N_6239,N_3934,N_3683);
and U6240 (N_6240,N_4206,N_3954);
nor U6241 (N_6241,N_4576,N_2943);
or U6242 (N_6242,N_3894,N_4695);
and U6243 (N_6243,N_4703,N_3929);
and U6244 (N_6244,N_4483,N_3595);
and U6245 (N_6245,N_4125,N_4639);
or U6246 (N_6246,N_4877,N_4566);
or U6247 (N_6247,N_2858,N_3960);
nor U6248 (N_6248,N_3577,N_3091);
and U6249 (N_6249,N_3000,N_4346);
xor U6250 (N_6250,N_4103,N_3374);
and U6251 (N_6251,N_2632,N_2717);
and U6252 (N_6252,N_4606,N_4031);
nor U6253 (N_6253,N_2928,N_4299);
or U6254 (N_6254,N_2840,N_4192);
and U6255 (N_6255,N_3088,N_4781);
and U6256 (N_6256,N_3031,N_2581);
nand U6257 (N_6257,N_4576,N_4615);
or U6258 (N_6258,N_3924,N_3501);
or U6259 (N_6259,N_3310,N_2755);
nor U6260 (N_6260,N_3924,N_3833);
and U6261 (N_6261,N_4245,N_4280);
or U6262 (N_6262,N_3472,N_2869);
or U6263 (N_6263,N_2567,N_3997);
or U6264 (N_6264,N_3177,N_4015);
nand U6265 (N_6265,N_3718,N_4635);
nand U6266 (N_6266,N_4731,N_2800);
nor U6267 (N_6267,N_3109,N_3775);
nor U6268 (N_6268,N_3855,N_2946);
and U6269 (N_6269,N_2502,N_3430);
nor U6270 (N_6270,N_2730,N_3027);
and U6271 (N_6271,N_3898,N_4352);
nor U6272 (N_6272,N_2820,N_4833);
and U6273 (N_6273,N_3827,N_2981);
or U6274 (N_6274,N_3561,N_4095);
and U6275 (N_6275,N_4549,N_4456);
or U6276 (N_6276,N_2868,N_4634);
nor U6277 (N_6277,N_3187,N_2703);
nand U6278 (N_6278,N_3715,N_2608);
nand U6279 (N_6279,N_3531,N_4774);
and U6280 (N_6280,N_3205,N_4500);
and U6281 (N_6281,N_3859,N_3779);
nand U6282 (N_6282,N_4010,N_4505);
nor U6283 (N_6283,N_3118,N_3062);
and U6284 (N_6284,N_4187,N_2983);
or U6285 (N_6285,N_3565,N_3923);
or U6286 (N_6286,N_3520,N_4937);
nor U6287 (N_6287,N_2750,N_3991);
nor U6288 (N_6288,N_2725,N_4212);
or U6289 (N_6289,N_4693,N_2916);
or U6290 (N_6290,N_3059,N_2693);
and U6291 (N_6291,N_3739,N_4302);
and U6292 (N_6292,N_4352,N_3539);
and U6293 (N_6293,N_3253,N_4588);
or U6294 (N_6294,N_4146,N_4359);
nor U6295 (N_6295,N_3159,N_4384);
nor U6296 (N_6296,N_3828,N_2977);
nand U6297 (N_6297,N_2779,N_3319);
nor U6298 (N_6298,N_3928,N_3075);
or U6299 (N_6299,N_3556,N_3405);
nand U6300 (N_6300,N_4277,N_4967);
nor U6301 (N_6301,N_4574,N_2685);
and U6302 (N_6302,N_3431,N_4564);
nand U6303 (N_6303,N_2750,N_4052);
or U6304 (N_6304,N_4095,N_3887);
or U6305 (N_6305,N_4222,N_4194);
or U6306 (N_6306,N_2836,N_2959);
nand U6307 (N_6307,N_3926,N_3586);
nand U6308 (N_6308,N_4358,N_2730);
nand U6309 (N_6309,N_2605,N_3983);
and U6310 (N_6310,N_4557,N_3387);
or U6311 (N_6311,N_4370,N_3117);
nor U6312 (N_6312,N_2588,N_3041);
and U6313 (N_6313,N_4181,N_4603);
nand U6314 (N_6314,N_4452,N_4465);
nand U6315 (N_6315,N_3209,N_2648);
nand U6316 (N_6316,N_2988,N_4002);
or U6317 (N_6317,N_4681,N_4405);
and U6318 (N_6318,N_4653,N_4399);
nand U6319 (N_6319,N_2612,N_4896);
nand U6320 (N_6320,N_4819,N_4712);
or U6321 (N_6321,N_2841,N_4318);
and U6322 (N_6322,N_4625,N_3041);
and U6323 (N_6323,N_4124,N_2553);
nand U6324 (N_6324,N_2953,N_4364);
or U6325 (N_6325,N_4857,N_4999);
xnor U6326 (N_6326,N_3814,N_2696);
nand U6327 (N_6327,N_4648,N_4103);
or U6328 (N_6328,N_3448,N_2814);
nand U6329 (N_6329,N_3487,N_2577);
nand U6330 (N_6330,N_3541,N_3417);
or U6331 (N_6331,N_4236,N_3861);
nand U6332 (N_6332,N_3766,N_4886);
nand U6333 (N_6333,N_4351,N_3004);
nor U6334 (N_6334,N_3925,N_3991);
nand U6335 (N_6335,N_2529,N_2583);
and U6336 (N_6336,N_4769,N_3785);
nor U6337 (N_6337,N_4652,N_3911);
nor U6338 (N_6338,N_4208,N_3856);
or U6339 (N_6339,N_4767,N_3345);
and U6340 (N_6340,N_4172,N_4747);
or U6341 (N_6341,N_3020,N_3408);
or U6342 (N_6342,N_2554,N_2609);
nand U6343 (N_6343,N_3731,N_3159);
nor U6344 (N_6344,N_4457,N_4371);
and U6345 (N_6345,N_4200,N_3636);
or U6346 (N_6346,N_3655,N_4677);
and U6347 (N_6347,N_4945,N_3546);
nand U6348 (N_6348,N_2617,N_2939);
or U6349 (N_6349,N_4033,N_3331);
or U6350 (N_6350,N_4643,N_2956);
nor U6351 (N_6351,N_2753,N_4505);
or U6352 (N_6352,N_3753,N_4655);
nor U6353 (N_6353,N_3236,N_2645);
and U6354 (N_6354,N_4542,N_4234);
or U6355 (N_6355,N_3386,N_3111);
or U6356 (N_6356,N_4380,N_2853);
nor U6357 (N_6357,N_4389,N_4567);
or U6358 (N_6358,N_2930,N_4090);
and U6359 (N_6359,N_2615,N_2611);
or U6360 (N_6360,N_4790,N_3033);
or U6361 (N_6361,N_4412,N_2760);
and U6362 (N_6362,N_3746,N_2713);
nand U6363 (N_6363,N_2836,N_4788);
or U6364 (N_6364,N_2812,N_4029);
xor U6365 (N_6365,N_2986,N_3087);
and U6366 (N_6366,N_3051,N_4702);
nand U6367 (N_6367,N_2666,N_4380);
or U6368 (N_6368,N_3418,N_3061);
or U6369 (N_6369,N_4149,N_3159);
nand U6370 (N_6370,N_4340,N_4635);
and U6371 (N_6371,N_4164,N_4329);
and U6372 (N_6372,N_2720,N_4439);
nor U6373 (N_6373,N_3490,N_3660);
nand U6374 (N_6374,N_4577,N_4898);
or U6375 (N_6375,N_4215,N_2789);
or U6376 (N_6376,N_4962,N_4545);
nand U6377 (N_6377,N_4457,N_4499);
nand U6378 (N_6378,N_3532,N_4037);
or U6379 (N_6379,N_3620,N_3440);
or U6380 (N_6380,N_2764,N_2699);
nand U6381 (N_6381,N_3703,N_4045);
and U6382 (N_6382,N_3800,N_3351);
nand U6383 (N_6383,N_4849,N_3544);
nand U6384 (N_6384,N_4041,N_3914);
nor U6385 (N_6385,N_2609,N_4047);
and U6386 (N_6386,N_2677,N_2696);
nor U6387 (N_6387,N_4763,N_4917);
and U6388 (N_6388,N_3485,N_3728);
or U6389 (N_6389,N_3364,N_3668);
nor U6390 (N_6390,N_2662,N_4009);
or U6391 (N_6391,N_3831,N_4545);
xnor U6392 (N_6392,N_4875,N_2711);
nand U6393 (N_6393,N_3966,N_2940);
or U6394 (N_6394,N_2714,N_3177);
nand U6395 (N_6395,N_3639,N_3791);
nand U6396 (N_6396,N_4891,N_3096);
nor U6397 (N_6397,N_2690,N_2976);
and U6398 (N_6398,N_2524,N_4602);
nor U6399 (N_6399,N_2792,N_2548);
or U6400 (N_6400,N_3049,N_3879);
and U6401 (N_6401,N_3720,N_4160);
and U6402 (N_6402,N_4131,N_2881);
and U6403 (N_6403,N_4979,N_4146);
nor U6404 (N_6404,N_3647,N_4618);
or U6405 (N_6405,N_4103,N_3249);
nor U6406 (N_6406,N_4256,N_3346);
and U6407 (N_6407,N_4147,N_4423);
nand U6408 (N_6408,N_3424,N_4791);
and U6409 (N_6409,N_4307,N_3977);
nand U6410 (N_6410,N_2559,N_3515);
nand U6411 (N_6411,N_4884,N_4310);
or U6412 (N_6412,N_3710,N_4038);
nand U6413 (N_6413,N_4235,N_4803);
nand U6414 (N_6414,N_4388,N_4693);
and U6415 (N_6415,N_2687,N_4782);
and U6416 (N_6416,N_4809,N_4396);
or U6417 (N_6417,N_3140,N_3168);
and U6418 (N_6418,N_3453,N_3396);
xor U6419 (N_6419,N_3493,N_3688);
nor U6420 (N_6420,N_2989,N_2861);
and U6421 (N_6421,N_4727,N_4582);
nor U6422 (N_6422,N_2895,N_4474);
nand U6423 (N_6423,N_4974,N_3808);
nand U6424 (N_6424,N_4276,N_4520);
and U6425 (N_6425,N_4905,N_3166);
nand U6426 (N_6426,N_3911,N_4076);
nand U6427 (N_6427,N_4349,N_3169);
or U6428 (N_6428,N_4181,N_4743);
nor U6429 (N_6429,N_4058,N_4858);
or U6430 (N_6430,N_3910,N_3044);
nand U6431 (N_6431,N_3622,N_3143);
nor U6432 (N_6432,N_3134,N_4640);
and U6433 (N_6433,N_4640,N_3847);
or U6434 (N_6434,N_3029,N_2948);
and U6435 (N_6435,N_3945,N_4357);
or U6436 (N_6436,N_3293,N_3394);
or U6437 (N_6437,N_2932,N_2559);
and U6438 (N_6438,N_4685,N_2568);
nor U6439 (N_6439,N_2979,N_4909);
and U6440 (N_6440,N_4843,N_4429);
and U6441 (N_6441,N_4500,N_3048);
nand U6442 (N_6442,N_2916,N_3129);
and U6443 (N_6443,N_3429,N_3077);
and U6444 (N_6444,N_2883,N_4348);
xor U6445 (N_6445,N_3194,N_3160);
or U6446 (N_6446,N_4312,N_3826);
and U6447 (N_6447,N_3258,N_2519);
xnor U6448 (N_6448,N_4716,N_2689);
nor U6449 (N_6449,N_2701,N_3874);
nor U6450 (N_6450,N_2563,N_3915);
nor U6451 (N_6451,N_3063,N_4854);
and U6452 (N_6452,N_3094,N_4931);
and U6453 (N_6453,N_4459,N_4783);
nand U6454 (N_6454,N_4037,N_2875);
or U6455 (N_6455,N_3812,N_3821);
or U6456 (N_6456,N_3353,N_4613);
nand U6457 (N_6457,N_2799,N_4881);
nor U6458 (N_6458,N_2902,N_3931);
nor U6459 (N_6459,N_4569,N_3309);
nand U6460 (N_6460,N_3264,N_4163);
xnor U6461 (N_6461,N_3356,N_3555);
and U6462 (N_6462,N_2716,N_3622);
and U6463 (N_6463,N_4639,N_4351);
and U6464 (N_6464,N_3744,N_3945);
nand U6465 (N_6465,N_3857,N_2755);
nand U6466 (N_6466,N_3861,N_4269);
nor U6467 (N_6467,N_2673,N_4891);
nor U6468 (N_6468,N_4144,N_2824);
nor U6469 (N_6469,N_2706,N_2847);
and U6470 (N_6470,N_3112,N_4843);
and U6471 (N_6471,N_3054,N_4464);
nand U6472 (N_6472,N_4602,N_3806);
nor U6473 (N_6473,N_4277,N_3953);
and U6474 (N_6474,N_3633,N_3483);
nor U6475 (N_6475,N_4433,N_4277);
nand U6476 (N_6476,N_4463,N_3026);
nor U6477 (N_6477,N_4151,N_3508);
and U6478 (N_6478,N_2822,N_4064);
or U6479 (N_6479,N_4360,N_3585);
nor U6480 (N_6480,N_3016,N_3030);
nand U6481 (N_6481,N_2778,N_2525);
nand U6482 (N_6482,N_4141,N_4754);
or U6483 (N_6483,N_2635,N_2746);
or U6484 (N_6484,N_2806,N_4007);
and U6485 (N_6485,N_2559,N_4698);
nand U6486 (N_6486,N_4097,N_3939);
or U6487 (N_6487,N_4826,N_4622);
or U6488 (N_6488,N_2749,N_4638);
or U6489 (N_6489,N_4017,N_3019);
nand U6490 (N_6490,N_3487,N_2867);
and U6491 (N_6491,N_3098,N_3021);
nor U6492 (N_6492,N_3607,N_3869);
nor U6493 (N_6493,N_3858,N_4466);
or U6494 (N_6494,N_3188,N_2864);
and U6495 (N_6495,N_3922,N_3317);
and U6496 (N_6496,N_4135,N_3418);
and U6497 (N_6497,N_3490,N_4544);
nand U6498 (N_6498,N_3273,N_3119);
or U6499 (N_6499,N_2625,N_4693);
nor U6500 (N_6500,N_3321,N_3748);
and U6501 (N_6501,N_4526,N_4575);
or U6502 (N_6502,N_3641,N_4026);
or U6503 (N_6503,N_2898,N_4775);
nand U6504 (N_6504,N_3239,N_4914);
nor U6505 (N_6505,N_3161,N_3654);
nand U6506 (N_6506,N_4003,N_2803);
nand U6507 (N_6507,N_4032,N_4123);
nand U6508 (N_6508,N_4550,N_3369);
or U6509 (N_6509,N_4845,N_4523);
or U6510 (N_6510,N_4543,N_3610);
and U6511 (N_6511,N_3176,N_2729);
and U6512 (N_6512,N_2791,N_3676);
and U6513 (N_6513,N_3825,N_2560);
nand U6514 (N_6514,N_4014,N_3612);
nand U6515 (N_6515,N_3909,N_2772);
nor U6516 (N_6516,N_3793,N_3405);
and U6517 (N_6517,N_4337,N_4499);
or U6518 (N_6518,N_4473,N_2857);
nor U6519 (N_6519,N_4856,N_3014);
or U6520 (N_6520,N_3883,N_4634);
nor U6521 (N_6521,N_4509,N_2971);
nor U6522 (N_6522,N_4012,N_4128);
nor U6523 (N_6523,N_2732,N_3186);
nor U6524 (N_6524,N_3391,N_3080);
nor U6525 (N_6525,N_3293,N_4944);
and U6526 (N_6526,N_3544,N_2980);
and U6527 (N_6527,N_4226,N_2575);
and U6528 (N_6528,N_3923,N_4488);
nor U6529 (N_6529,N_4483,N_3319);
nor U6530 (N_6530,N_3681,N_4017);
and U6531 (N_6531,N_3146,N_2590);
and U6532 (N_6532,N_4816,N_3688);
and U6533 (N_6533,N_4950,N_4693);
or U6534 (N_6534,N_3791,N_3952);
nor U6535 (N_6535,N_2962,N_2595);
nor U6536 (N_6536,N_4043,N_3057);
nor U6537 (N_6537,N_2841,N_3608);
and U6538 (N_6538,N_3819,N_4512);
or U6539 (N_6539,N_4288,N_3195);
nor U6540 (N_6540,N_4068,N_3607);
or U6541 (N_6541,N_4094,N_2864);
and U6542 (N_6542,N_3705,N_4053);
and U6543 (N_6543,N_4531,N_4329);
nand U6544 (N_6544,N_3968,N_2871);
and U6545 (N_6545,N_4708,N_4124);
or U6546 (N_6546,N_4902,N_3248);
or U6547 (N_6547,N_3625,N_3380);
nand U6548 (N_6548,N_4418,N_2734);
or U6549 (N_6549,N_2519,N_3796);
nand U6550 (N_6550,N_3810,N_3324);
and U6551 (N_6551,N_4035,N_3768);
nor U6552 (N_6552,N_4520,N_4448);
xor U6553 (N_6553,N_4480,N_3241);
and U6554 (N_6554,N_4601,N_2556);
xor U6555 (N_6555,N_3351,N_4749);
or U6556 (N_6556,N_4621,N_4428);
and U6557 (N_6557,N_3776,N_4913);
nand U6558 (N_6558,N_4722,N_4182);
and U6559 (N_6559,N_4883,N_3011);
nor U6560 (N_6560,N_4996,N_3656);
nor U6561 (N_6561,N_3619,N_3248);
or U6562 (N_6562,N_4004,N_4203);
and U6563 (N_6563,N_3291,N_3096);
nand U6564 (N_6564,N_3290,N_2611);
nor U6565 (N_6565,N_2966,N_3682);
and U6566 (N_6566,N_2750,N_2980);
nand U6567 (N_6567,N_4584,N_3541);
nor U6568 (N_6568,N_4851,N_3641);
and U6569 (N_6569,N_2957,N_4117);
and U6570 (N_6570,N_4156,N_3475);
nor U6571 (N_6571,N_2870,N_4032);
or U6572 (N_6572,N_3713,N_4909);
or U6573 (N_6573,N_3041,N_3676);
nor U6574 (N_6574,N_2941,N_4910);
nand U6575 (N_6575,N_4871,N_4809);
or U6576 (N_6576,N_2952,N_4734);
and U6577 (N_6577,N_4615,N_2921);
nor U6578 (N_6578,N_4369,N_2710);
nor U6579 (N_6579,N_2556,N_3255);
nand U6580 (N_6580,N_3764,N_4955);
and U6581 (N_6581,N_4988,N_2962);
or U6582 (N_6582,N_3608,N_4348);
and U6583 (N_6583,N_3182,N_3575);
nor U6584 (N_6584,N_2718,N_2832);
and U6585 (N_6585,N_2795,N_4660);
nand U6586 (N_6586,N_3309,N_4205);
or U6587 (N_6587,N_2681,N_3278);
nand U6588 (N_6588,N_4162,N_2785);
or U6589 (N_6589,N_2687,N_4213);
nor U6590 (N_6590,N_3836,N_2951);
or U6591 (N_6591,N_4901,N_4778);
or U6592 (N_6592,N_4039,N_3713);
nand U6593 (N_6593,N_3130,N_2604);
or U6594 (N_6594,N_4054,N_4709);
nor U6595 (N_6595,N_4166,N_4810);
and U6596 (N_6596,N_4857,N_4529);
or U6597 (N_6597,N_2657,N_2530);
xor U6598 (N_6598,N_2890,N_4470);
or U6599 (N_6599,N_4390,N_2950);
nor U6600 (N_6600,N_3495,N_3347);
nand U6601 (N_6601,N_2511,N_3308);
nand U6602 (N_6602,N_3389,N_2794);
and U6603 (N_6603,N_4741,N_4803);
or U6604 (N_6604,N_3744,N_2721);
and U6605 (N_6605,N_4831,N_2910);
and U6606 (N_6606,N_4045,N_4050);
nand U6607 (N_6607,N_3637,N_3421);
and U6608 (N_6608,N_4267,N_4887);
and U6609 (N_6609,N_4425,N_2500);
and U6610 (N_6610,N_3201,N_3175);
or U6611 (N_6611,N_2995,N_2730);
or U6612 (N_6612,N_4782,N_4319);
nor U6613 (N_6613,N_3245,N_3397);
nand U6614 (N_6614,N_3737,N_4291);
nand U6615 (N_6615,N_3653,N_4425);
or U6616 (N_6616,N_4402,N_3185);
nand U6617 (N_6617,N_3742,N_3003);
and U6618 (N_6618,N_3582,N_4674);
nand U6619 (N_6619,N_3538,N_3026);
and U6620 (N_6620,N_4616,N_4498);
and U6621 (N_6621,N_3993,N_3326);
or U6622 (N_6622,N_4194,N_4578);
and U6623 (N_6623,N_4834,N_2726);
and U6624 (N_6624,N_4237,N_3742);
nand U6625 (N_6625,N_3758,N_3062);
and U6626 (N_6626,N_2925,N_3917);
or U6627 (N_6627,N_4341,N_3047);
nand U6628 (N_6628,N_3599,N_4571);
nor U6629 (N_6629,N_2869,N_2885);
nor U6630 (N_6630,N_3843,N_2900);
nand U6631 (N_6631,N_3073,N_3027);
nor U6632 (N_6632,N_3905,N_2844);
and U6633 (N_6633,N_3565,N_4114);
nor U6634 (N_6634,N_3277,N_4471);
nand U6635 (N_6635,N_2826,N_4259);
nand U6636 (N_6636,N_4267,N_4816);
or U6637 (N_6637,N_3459,N_4071);
or U6638 (N_6638,N_3532,N_4758);
or U6639 (N_6639,N_4251,N_4052);
and U6640 (N_6640,N_4540,N_4159);
nor U6641 (N_6641,N_3357,N_3860);
nand U6642 (N_6642,N_4607,N_3868);
nor U6643 (N_6643,N_3844,N_4587);
or U6644 (N_6644,N_3909,N_3123);
nand U6645 (N_6645,N_3005,N_3688);
nor U6646 (N_6646,N_3992,N_3940);
nor U6647 (N_6647,N_3866,N_4658);
or U6648 (N_6648,N_4338,N_3897);
nand U6649 (N_6649,N_4756,N_2979);
and U6650 (N_6650,N_3030,N_3129);
and U6651 (N_6651,N_3045,N_3750);
and U6652 (N_6652,N_3127,N_4436);
nand U6653 (N_6653,N_4305,N_3318);
nor U6654 (N_6654,N_4671,N_4390);
or U6655 (N_6655,N_4082,N_3793);
nand U6656 (N_6656,N_3302,N_3039);
and U6657 (N_6657,N_3205,N_2592);
and U6658 (N_6658,N_3355,N_4602);
nor U6659 (N_6659,N_4328,N_3879);
nor U6660 (N_6660,N_3011,N_3109);
and U6661 (N_6661,N_3857,N_3501);
nand U6662 (N_6662,N_3341,N_4099);
or U6663 (N_6663,N_4702,N_4575);
and U6664 (N_6664,N_2995,N_4046);
nor U6665 (N_6665,N_3684,N_2991);
xor U6666 (N_6666,N_4582,N_3401);
and U6667 (N_6667,N_3609,N_3204);
nand U6668 (N_6668,N_4614,N_3572);
and U6669 (N_6669,N_3845,N_3480);
nor U6670 (N_6670,N_3797,N_3630);
nand U6671 (N_6671,N_3513,N_4563);
or U6672 (N_6672,N_4293,N_2784);
nand U6673 (N_6673,N_3045,N_2741);
or U6674 (N_6674,N_4004,N_4068);
nor U6675 (N_6675,N_4394,N_3677);
nor U6676 (N_6676,N_2995,N_4107);
nor U6677 (N_6677,N_2523,N_4286);
nand U6678 (N_6678,N_3884,N_3993);
nor U6679 (N_6679,N_3234,N_3983);
and U6680 (N_6680,N_4324,N_3629);
nand U6681 (N_6681,N_4665,N_4604);
or U6682 (N_6682,N_4481,N_2853);
or U6683 (N_6683,N_4981,N_3936);
nor U6684 (N_6684,N_3080,N_4919);
and U6685 (N_6685,N_3224,N_4561);
or U6686 (N_6686,N_4702,N_2936);
or U6687 (N_6687,N_4643,N_4912);
nand U6688 (N_6688,N_4528,N_2903);
and U6689 (N_6689,N_3153,N_2725);
and U6690 (N_6690,N_2587,N_2796);
or U6691 (N_6691,N_4415,N_4269);
nand U6692 (N_6692,N_3981,N_3919);
and U6693 (N_6693,N_4497,N_2937);
and U6694 (N_6694,N_4866,N_4858);
nand U6695 (N_6695,N_3622,N_3352);
nor U6696 (N_6696,N_4003,N_3845);
and U6697 (N_6697,N_4006,N_2754);
nand U6698 (N_6698,N_2691,N_4579);
and U6699 (N_6699,N_2534,N_2768);
or U6700 (N_6700,N_4141,N_4316);
nor U6701 (N_6701,N_2806,N_4742);
nor U6702 (N_6702,N_4651,N_4316);
or U6703 (N_6703,N_4036,N_3611);
or U6704 (N_6704,N_4466,N_4221);
and U6705 (N_6705,N_4842,N_3140);
nand U6706 (N_6706,N_4693,N_4561);
or U6707 (N_6707,N_2681,N_2550);
nor U6708 (N_6708,N_2908,N_3701);
nor U6709 (N_6709,N_2828,N_3327);
nand U6710 (N_6710,N_4053,N_4012);
nand U6711 (N_6711,N_3072,N_4901);
nor U6712 (N_6712,N_3514,N_3603);
nor U6713 (N_6713,N_4595,N_4138);
and U6714 (N_6714,N_3896,N_4144);
or U6715 (N_6715,N_2973,N_2575);
or U6716 (N_6716,N_4823,N_4564);
nand U6717 (N_6717,N_4391,N_2903);
or U6718 (N_6718,N_2899,N_3431);
or U6719 (N_6719,N_3807,N_2573);
and U6720 (N_6720,N_3659,N_3054);
or U6721 (N_6721,N_4069,N_3143);
nand U6722 (N_6722,N_4591,N_4184);
and U6723 (N_6723,N_3390,N_2722);
or U6724 (N_6724,N_3805,N_2780);
xor U6725 (N_6725,N_2529,N_3627);
nand U6726 (N_6726,N_4342,N_4848);
and U6727 (N_6727,N_4637,N_4914);
and U6728 (N_6728,N_3249,N_4346);
nor U6729 (N_6729,N_4980,N_4136);
nand U6730 (N_6730,N_3032,N_4638);
nand U6731 (N_6731,N_4912,N_3644);
nand U6732 (N_6732,N_2569,N_4645);
and U6733 (N_6733,N_2646,N_4223);
or U6734 (N_6734,N_3492,N_3758);
nand U6735 (N_6735,N_3622,N_4108);
nand U6736 (N_6736,N_2965,N_3924);
nand U6737 (N_6737,N_3921,N_3911);
and U6738 (N_6738,N_4823,N_3587);
nor U6739 (N_6739,N_3975,N_3249);
or U6740 (N_6740,N_3201,N_4483);
nor U6741 (N_6741,N_4290,N_3845);
or U6742 (N_6742,N_4643,N_4258);
or U6743 (N_6743,N_4732,N_3004);
or U6744 (N_6744,N_3346,N_3906);
or U6745 (N_6745,N_3741,N_2740);
nand U6746 (N_6746,N_4176,N_4667);
nand U6747 (N_6747,N_4149,N_3596);
xnor U6748 (N_6748,N_3710,N_4931);
and U6749 (N_6749,N_3860,N_4798);
nand U6750 (N_6750,N_3475,N_4974);
or U6751 (N_6751,N_2534,N_4884);
and U6752 (N_6752,N_4678,N_3127);
or U6753 (N_6753,N_4742,N_4832);
nand U6754 (N_6754,N_3999,N_3059);
nor U6755 (N_6755,N_3617,N_4993);
nor U6756 (N_6756,N_4120,N_4242);
and U6757 (N_6757,N_4040,N_2993);
nand U6758 (N_6758,N_4712,N_3235);
or U6759 (N_6759,N_3967,N_2543);
nor U6760 (N_6760,N_4887,N_2597);
and U6761 (N_6761,N_2778,N_3468);
and U6762 (N_6762,N_3732,N_3884);
nor U6763 (N_6763,N_4946,N_4328);
and U6764 (N_6764,N_4577,N_4989);
or U6765 (N_6765,N_4527,N_3299);
nor U6766 (N_6766,N_4263,N_2986);
and U6767 (N_6767,N_4366,N_3656);
and U6768 (N_6768,N_4413,N_4513);
xnor U6769 (N_6769,N_4990,N_4293);
nor U6770 (N_6770,N_4237,N_3867);
nand U6771 (N_6771,N_2851,N_3892);
or U6772 (N_6772,N_4104,N_4159);
nor U6773 (N_6773,N_2953,N_2742);
and U6774 (N_6774,N_4679,N_4360);
and U6775 (N_6775,N_4542,N_2695);
or U6776 (N_6776,N_2592,N_3206);
or U6777 (N_6777,N_3220,N_4510);
nand U6778 (N_6778,N_3178,N_4227);
nor U6779 (N_6779,N_4359,N_4231);
and U6780 (N_6780,N_3256,N_4849);
or U6781 (N_6781,N_3009,N_4651);
and U6782 (N_6782,N_4656,N_3084);
or U6783 (N_6783,N_3622,N_4801);
nand U6784 (N_6784,N_3549,N_4061);
or U6785 (N_6785,N_4633,N_3404);
and U6786 (N_6786,N_3690,N_3113);
nand U6787 (N_6787,N_3729,N_4306);
and U6788 (N_6788,N_3378,N_3283);
or U6789 (N_6789,N_3000,N_4887);
nand U6790 (N_6790,N_4788,N_3071);
and U6791 (N_6791,N_3888,N_3439);
nand U6792 (N_6792,N_3463,N_2625);
or U6793 (N_6793,N_3435,N_4336);
and U6794 (N_6794,N_4619,N_2859);
nor U6795 (N_6795,N_2643,N_3635);
nor U6796 (N_6796,N_2871,N_3751);
or U6797 (N_6797,N_3857,N_3138);
or U6798 (N_6798,N_4141,N_3942);
nand U6799 (N_6799,N_3460,N_3018);
nor U6800 (N_6800,N_4373,N_2962);
nor U6801 (N_6801,N_2547,N_3173);
nand U6802 (N_6802,N_2953,N_3302);
and U6803 (N_6803,N_3357,N_4527);
and U6804 (N_6804,N_4049,N_3012);
nor U6805 (N_6805,N_3059,N_4933);
nand U6806 (N_6806,N_3769,N_3869);
or U6807 (N_6807,N_3362,N_3490);
or U6808 (N_6808,N_4139,N_3345);
or U6809 (N_6809,N_2610,N_2922);
nand U6810 (N_6810,N_4891,N_3271);
and U6811 (N_6811,N_2646,N_4214);
nand U6812 (N_6812,N_4177,N_4312);
nand U6813 (N_6813,N_4397,N_3707);
or U6814 (N_6814,N_4230,N_3186);
and U6815 (N_6815,N_4552,N_3065);
and U6816 (N_6816,N_3091,N_4543);
nor U6817 (N_6817,N_2897,N_4739);
nor U6818 (N_6818,N_4331,N_3824);
nor U6819 (N_6819,N_4574,N_3586);
or U6820 (N_6820,N_4423,N_3848);
nand U6821 (N_6821,N_3318,N_4204);
nor U6822 (N_6822,N_3209,N_3126);
and U6823 (N_6823,N_4135,N_2952);
and U6824 (N_6824,N_2771,N_3859);
nand U6825 (N_6825,N_4294,N_4951);
and U6826 (N_6826,N_2965,N_3254);
nand U6827 (N_6827,N_2993,N_2581);
nor U6828 (N_6828,N_4235,N_2578);
or U6829 (N_6829,N_4634,N_3127);
and U6830 (N_6830,N_4393,N_3788);
and U6831 (N_6831,N_2804,N_3517);
nor U6832 (N_6832,N_2831,N_4468);
and U6833 (N_6833,N_4807,N_4636);
nor U6834 (N_6834,N_4857,N_2909);
or U6835 (N_6835,N_3326,N_4729);
nor U6836 (N_6836,N_3642,N_2566);
nand U6837 (N_6837,N_4164,N_2590);
nand U6838 (N_6838,N_4666,N_2773);
and U6839 (N_6839,N_4256,N_3506);
nor U6840 (N_6840,N_2977,N_3543);
or U6841 (N_6841,N_3347,N_3886);
nor U6842 (N_6842,N_3324,N_3961);
and U6843 (N_6843,N_4395,N_4079);
and U6844 (N_6844,N_3418,N_3112);
nor U6845 (N_6845,N_3791,N_4132);
nand U6846 (N_6846,N_2632,N_4255);
or U6847 (N_6847,N_3017,N_4997);
nor U6848 (N_6848,N_3904,N_4537);
nor U6849 (N_6849,N_4172,N_4263);
nand U6850 (N_6850,N_3462,N_3325);
nor U6851 (N_6851,N_2559,N_3949);
or U6852 (N_6852,N_3624,N_2924);
nor U6853 (N_6853,N_4091,N_3883);
and U6854 (N_6854,N_4825,N_2985);
nand U6855 (N_6855,N_3525,N_4650);
nand U6856 (N_6856,N_4100,N_2735);
or U6857 (N_6857,N_3631,N_3482);
nor U6858 (N_6858,N_3842,N_2900);
and U6859 (N_6859,N_3603,N_3207);
and U6860 (N_6860,N_4240,N_3603);
nand U6861 (N_6861,N_4768,N_3354);
nor U6862 (N_6862,N_4210,N_2865);
nand U6863 (N_6863,N_3890,N_4045);
nand U6864 (N_6864,N_4305,N_4777);
nor U6865 (N_6865,N_3940,N_4920);
and U6866 (N_6866,N_3921,N_2633);
nand U6867 (N_6867,N_4198,N_4171);
nand U6868 (N_6868,N_3272,N_2911);
nand U6869 (N_6869,N_3871,N_2947);
nand U6870 (N_6870,N_3886,N_4432);
nor U6871 (N_6871,N_3133,N_3572);
and U6872 (N_6872,N_3308,N_4700);
xor U6873 (N_6873,N_3462,N_3942);
and U6874 (N_6874,N_4818,N_4009);
or U6875 (N_6875,N_2898,N_4707);
and U6876 (N_6876,N_2795,N_4220);
nand U6877 (N_6877,N_2904,N_4254);
nand U6878 (N_6878,N_4512,N_3860);
nor U6879 (N_6879,N_4245,N_3634);
or U6880 (N_6880,N_3812,N_4599);
nor U6881 (N_6881,N_4647,N_3654);
and U6882 (N_6882,N_2534,N_4723);
or U6883 (N_6883,N_4157,N_2628);
nor U6884 (N_6884,N_4328,N_3735);
or U6885 (N_6885,N_3503,N_3480);
nand U6886 (N_6886,N_4837,N_3736);
xnor U6887 (N_6887,N_2944,N_4490);
nor U6888 (N_6888,N_3281,N_4545);
nand U6889 (N_6889,N_2567,N_3679);
nand U6890 (N_6890,N_4253,N_4245);
and U6891 (N_6891,N_3126,N_2722);
and U6892 (N_6892,N_3020,N_2968);
and U6893 (N_6893,N_3228,N_3385);
nor U6894 (N_6894,N_4878,N_3386);
or U6895 (N_6895,N_3285,N_2809);
nand U6896 (N_6896,N_3666,N_3037);
nand U6897 (N_6897,N_2977,N_3167);
nor U6898 (N_6898,N_3942,N_3859);
nor U6899 (N_6899,N_4600,N_3347);
nand U6900 (N_6900,N_2732,N_2801);
and U6901 (N_6901,N_4522,N_4642);
nor U6902 (N_6902,N_3244,N_2882);
or U6903 (N_6903,N_2507,N_3827);
and U6904 (N_6904,N_2653,N_3177);
and U6905 (N_6905,N_3803,N_4410);
or U6906 (N_6906,N_3462,N_3657);
nand U6907 (N_6907,N_4598,N_4426);
nand U6908 (N_6908,N_4636,N_2836);
nor U6909 (N_6909,N_3097,N_2788);
and U6910 (N_6910,N_4554,N_4229);
or U6911 (N_6911,N_3065,N_3149);
and U6912 (N_6912,N_4126,N_2980);
or U6913 (N_6913,N_3881,N_4523);
or U6914 (N_6914,N_4796,N_4757);
nor U6915 (N_6915,N_3121,N_4136);
nor U6916 (N_6916,N_4904,N_3607);
nor U6917 (N_6917,N_3783,N_3368);
or U6918 (N_6918,N_3439,N_3155);
or U6919 (N_6919,N_4511,N_3281);
nand U6920 (N_6920,N_4696,N_3081);
and U6921 (N_6921,N_4685,N_2864);
nor U6922 (N_6922,N_4992,N_3644);
nor U6923 (N_6923,N_4119,N_3547);
or U6924 (N_6924,N_2768,N_3949);
nand U6925 (N_6925,N_4488,N_4368);
or U6926 (N_6926,N_3596,N_3516);
nor U6927 (N_6927,N_4942,N_4504);
nand U6928 (N_6928,N_4023,N_3661);
nor U6929 (N_6929,N_3536,N_2915);
nor U6930 (N_6930,N_3559,N_4376);
or U6931 (N_6931,N_3366,N_4750);
and U6932 (N_6932,N_4805,N_4509);
or U6933 (N_6933,N_3119,N_3542);
nand U6934 (N_6934,N_3915,N_3047);
and U6935 (N_6935,N_4207,N_4376);
or U6936 (N_6936,N_4145,N_2810);
or U6937 (N_6937,N_4983,N_2624);
or U6938 (N_6938,N_4584,N_4805);
nor U6939 (N_6939,N_4847,N_3203);
nor U6940 (N_6940,N_4202,N_3203);
or U6941 (N_6941,N_3766,N_4719);
and U6942 (N_6942,N_4523,N_4613);
and U6943 (N_6943,N_4331,N_4367);
and U6944 (N_6944,N_3024,N_3139);
and U6945 (N_6945,N_4740,N_2985);
nand U6946 (N_6946,N_3487,N_4287);
nand U6947 (N_6947,N_4088,N_4159);
nor U6948 (N_6948,N_3480,N_4982);
nand U6949 (N_6949,N_2904,N_4427);
or U6950 (N_6950,N_4682,N_4463);
nor U6951 (N_6951,N_4545,N_2883);
nor U6952 (N_6952,N_4727,N_3839);
nor U6953 (N_6953,N_4320,N_2706);
and U6954 (N_6954,N_4161,N_4839);
and U6955 (N_6955,N_4585,N_3034);
and U6956 (N_6956,N_3865,N_4018);
and U6957 (N_6957,N_3825,N_4829);
or U6958 (N_6958,N_3520,N_4208);
or U6959 (N_6959,N_3431,N_4607);
nand U6960 (N_6960,N_4221,N_3531);
and U6961 (N_6961,N_3812,N_4744);
nand U6962 (N_6962,N_3641,N_4758);
nor U6963 (N_6963,N_4350,N_3259);
and U6964 (N_6964,N_4315,N_4357);
nand U6965 (N_6965,N_4401,N_3998);
nor U6966 (N_6966,N_3118,N_4227);
or U6967 (N_6967,N_2920,N_4754);
nor U6968 (N_6968,N_3658,N_4024);
nor U6969 (N_6969,N_3391,N_4781);
nor U6970 (N_6970,N_3759,N_4949);
and U6971 (N_6971,N_3633,N_4574);
and U6972 (N_6972,N_4003,N_4133);
or U6973 (N_6973,N_3909,N_3168);
or U6974 (N_6974,N_3398,N_4645);
nor U6975 (N_6975,N_3697,N_2724);
nor U6976 (N_6976,N_3785,N_2572);
or U6977 (N_6977,N_4701,N_4942);
nor U6978 (N_6978,N_4270,N_4163);
or U6979 (N_6979,N_3601,N_4499);
or U6980 (N_6980,N_2730,N_3861);
nor U6981 (N_6981,N_3477,N_4158);
and U6982 (N_6982,N_3234,N_2568);
and U6983 (N_6983,N_3300,N_2993);
nor U6984 (N_6984,N_4441,N_4767);
and U6985 (N_6985,N_4781,N_3485);
and U6986 (N_6986,N_4606,N_4738);
nor U6987 (N_6987,N_4042,N_2916);
nor U6988 (N_6988,N_3853,N_4629);
nor U6989 (N_6989,N_4511,N_4126);
and U6990 (N_6990,N_3819,N_3265);
nor U6991 (N_6991,N_3417,N_3274);
nand U6992 (N_6992,N_4096,N_2956);
nand U6993 (N_6993,N_3619,N_3943);
or U6994 (N_6994,N_4382,N_4015);
or U6995 (N_6995,N_3758,N_3903);
nor U6996 (N_6996,N_3388,N_4062);
and U6997 (N_6997,N_3856,N_4715);
nand U6998 (N_6998,N_2895,N_4013);
or U6999 (N_6999,N_2538,N_3454);
or U7000 (N_7000,N_4503,N_4094);
or U7001 (N_7001,N_3736,N_4293);
nor U7002 (N_7002,N_2557,N_3715);
or U7003 (N_7003,N_4067,N_2578);
and U7004 (N_7004,N_4104,N_3974);
or U7005 (N_7005,N_3170,N_3600);
nor U7006 (N_7006,N_2925,N_3852);
nand U7007 (N_7007,N_4224,N_3258);
and U7008 (N_7008,N_4273,N_3791);
and U7009 (N_7009,N_4943,N_2684);
or U7010 (N_7010,N_3594,N_3165);
and U7011 (N_7011,N_3355,N_3725);
nand U7012 (N_7012,N_3716,N_4396);
nor U7013 (N_7013,N_3221,N_4972);
nand U7014 (N_7014,N_4815,N_3461);
or U7015 (N_7015,N_4250,N_4309);
nand U7016 (N_7016,N_2875,N_4531);
nor U7017 (N_7017,N_4913,N_3629);
nor U7018 (N_7018,N_3544,N_2803);
nand U7019 (N_7019,N_4857,N_2955);
or U7020 (N_7020,N_3488,N_3026);
nand U7021 (N_7021,N_3362,N_4324);
and U7022 (N_7022,N_4170,N_3707);
and U7023 (N_7023,N_4494,N_3800);
nand U7024 (N_7024,N_2828,N_3046);
nor U7025 (N_7025,N_3781,N_4760);
nor U7026 (N_7026,N_3944,N_4064);
or U7027 (N_7027,N_4025,N_4052);
nor U7028 (N_7028,N_2740,N_4016);
or U7029 (N_7029,N_2560,N_2622);
or U7030 (N_7030,N_2931,N_3781);
nand U7031 (N_7031,N_2818,N_2724);
nand U7032 (N_7032,N_3331,N_4958);
and U7033 (N_7033,N_2892,N_3175);
nor U7034 (N_7034,N_2937,N_4739);
or U7035 (N_7035,N_3416,N_3492);
and U7036 (N_7036,N_3055,N_3217);
nor U7037 (N_7037,N_4480,N_4402);
nand U7038 (N_7038,N_3868,N_2799);
or U7039 (N_7039,N_3825,N_3038);
nor U7040 (N_7040,N_3101,N_4987);
or U7041 (N_7041,N_4787,N_4486);
nor U7042 (N_7042,N_4950,N_4689);
or U7043 (N_7043,N_3100,N_3955);
or U7044 (N_7044,N_2881,N_3107);
nand U7045 (N_7045,N_3051,N_3522);
nand U7046 (N_7046,N_2757,N_3467);
nor U7047 (N_7047,N_2890,N_3109);
nor U7048 (N_7048,N_4980,N_3772);
or U7049 (N_7049,N_4949,N_4979);
nor U7050 (N_7050,N_3246,N_3836);
and U7051 (N_7051,N_4362,N_4996);
or U7052 (N_7052,N_2681,N_4628);
nor U7053 (N_7053,N_4845,N_2947);
nor U7054 (N_7054,N_2892,N_2569);
or U7055 (N_7055,N_3264,N_4915);
nor U7056 (N_7056,N_3189,N_2853);
and U7057 (N_7057,N_2662,N_4448);
nor U7058 (N_7058,N_4166,N_4780);
and U7059 (N_7059,N_3058,N_2860);
nor U7060 (N_7060,N_3970,N_3790);
nand U7061 (N_7061,N_2618,N_3587);
or U7062 (N_7062,N_4300,N_4196);
nand U7063 (N_7063,N_3607,N_4058);
or U7064 (N_7064,N_3736,N_3878);
nor U7065 (N_7065,N_4313,N_4628);
nor U7066 (N_7066,N_4217,N_3651);
and U7067 (N_7067,N_4703,N_3942);
nand U7068 (N_7068,N_4509,N_3246);
nor U7069 (N_7069,N_4149,N_4175);
and U7070 (N_7070,N_4677,N_4420);
or U7071 (N_7071,N_4847,N_4634);
and U7072 (N_7072,N_3903,N_4497);
xor U7073 (N_7073,N_3627,N_4929);
nand U7074 (N_7074,N_3267,N_4713);
nand U7075 (N_7075,N_2679,N_4835);
and U7076 (N_7076,N_3183,N_2726);
nor U7077 (N_7077,N_2988,N_3347);
and U7078 (N_7078,N_4871,N_2732);
nor U7079 (N_7079,N_4618,N_3564);
and U7080 (N_7080,N_3312,N_4012);
or U7081 (N_7081,N_3004,N_2914);
nand U7082 (N_7082,N_2735,N_4130);
or U7083 (N_7083,N_3704,N_4655);
and U7084 (N_7084,N_3988,N_4676);
or U7085 (N_7085,N_3736,N_4563);
nor U7086 (N_7086,N_4866,N_4897);
nand U7087 (N_7087,N_4142,N_3062);
nand U7088 (N_7088,N_4675,N_3114);
nand U7089 (N_7089,N_3851,N_2798);
nor U7090 (N_7090,N_4830,N_3318);
nor U7091 (N_7091,N_3988,N_3380);
nand U7092 (N_7092,N_3871,N_2777);
and U7093 (N_7093,N_2551,N_3037);
and U7094 (N_7094,N_4247,N_2884);
or U7095 (N_7095,N_3726,N_4971);
nor U7096 (N_7096,N_4071,N_2540);
nand U7097 (N_7097,N_3870,N_2764);
or U7098 (N_7098,N_2842,N_3249);
nor U7099 (N_7099,N_2995,N_4718);
and U7100 (N_7100,N_3723,N_2507);
or U7101 (N_7101,N_4732,N_4404);
or U7102 (N_7102,N_4996,N_3696);
and U7103 (N_7103,N_3569,N_2585);
and U7104 (N_7104,N_4452,N_3713);
and U7105 (N_7105,N_4667,N_2559);
and U7106 (N_7106,N_4331,N_4395);
nor U7107 (N_7107,N_3269,N_4569);
and U7108 (N_7108,N_3136,N_4791);
nand U7109 (N_7109,N_4123,N_3677);
and U7110 (N_7110,N_4709,N_4932);
nand U7111 (N_7111,N_3023,N_4132);
nand U7112 (N_7112,N_4671,N_4724);
and U7113 (N_7113,N_2595,N_4532);
nand U7114 (N_7114,N_2929,N_2968);
and U7115 (N_7115,N_2688,N_4821);
nand U7116 (N_7116,N_4114,N_2863);
nor U7117 (N_7117,N_2523,N_3181);
nand U7118 (N_7118,N_2910,N_4686);
nor U7119 (N_7119,N_4922,N_3810);
and U7120 (N_7120,N_4593,N_3999);
nand U7121 (N_7121,N_4911,N_4971);
nor U7122 (N_7122,N_3754,N_2519);
or U7123 (N_7123,N_3942,N_3292);
or U7124 (N_7124,N_4106,N_3627);
nand U7125 (N_7125,N_3496,N_4760);
or U7126 (N_7126,N_4984,N_3725);
or U7127 (N_7127,N_3283,N_3359);
or U7128 (N_7128,N_3859,N_2566);
nand U7129 (N_7129,N_4180,N_3847);
nand U7130 (N_7130,N_4856,N_4649);
or U7131 (N_7131,N_3189,N_3055);
nand U7132 (N_7132,N_3207,N_2689);
or U7133 (N_7133,N_4121,N_3375);
xnor U7134 (N_7134,N_3813,N_4620);
and U7135 (N_7135,N_2969,N_2556);
nor U7136 (N_7136,N_3933,N_3096);
nor U7137 (N_7137,N_3217,N_3324);
nand U7138 (N_7138,N_3462,N_3876);
nor U7139 (N_7139,N_3517,N_4790);
or U7140 (N_7140,N_2669,N_3593);
or U7141 (N_7141,N_2883,N_3610);
and U7142 (N_7142,N_3779,N_4728);
nand U7143 (N_7143,N_3339,N_3028);
or U7144 (N_7144,N_2709,N_3639);
nor U7145 (N_7145,N_2624,N_4251);
or U7146 (N_7146,N_4470,N_4785);
nand U7147 (N_7147,N_4825,N_2652);
nand U7148 (N_7148,N_4099,N_3271);
and U7149 (N_7149,N_3010,N_2654);
xor U7150 (N_7150,N_2732,N_3091);
and U7151 (N_7151,N_3947,N_3640);
and U7152 (N_7152,N_4629,N_4433);
nor U7153 (N_7153,N_4272,N_4588);
nor U7154 (N_7154,N_2786,N_3975);
and U7155 (N_7155,N_4968,N_3048);
and U7156 (N_7156,N_3486,N_3089);
or U7157 (N_7157,N_3946,N_4244);
nor U7158 (N_7158,N_2734,N_3178);
nand U7159 (N_7159,N_3201,N_4398);
nor U7160 (N_7160,N_4565,N_3268);
nor U7161 (N_7161,N_3099,N_4470);
nand U7162 (N_7162,N_2955,N_4687);
nor U7163 (N_7163,N_4741,N_3273);
nor U7164 (N_7164,N_4787,N_4244);
nor U7165 (N_7165,N_2816,N_3298);
nand U7166 (N_7166,N_3565,N_3014);
nand U7167 (N_7167,N_4890,N_4112);
and U7168 (N_7168,N_3629,N_3689);
nand U7169 (N_7169,N_3018,N_3097);
nor U7170 (N_7170,N_2924,N_4214);
and U7171 (N_7171,N_4710,N_3607);
nand U7172 (N_7172,N_3460,N_3188);
and U7173 (N_7173,N_2903,N_3131);
nand U7174 (N_7174,N_4181,N_2538);
or U7175 (N_7175,N_4328,N_2562);
nand U7176 (N_7176,N_3625,N_2842);
nor U7177 (N_7177,N_4422,N_3785);
nor U7178 (N_7178,N_4835,N_2817);
and U7179 (N_7179,N_4504,N_4329);
and U7180 (N_7180,N_3213,N_3265);
nor U7181 (N_7181,N_2936,N_4947);
and U7182 (N_7182,N_4638,N_4492);
and U7183 (N_7183,N_4065,N_4856);
nand U7184 (N_7184,N_3665,N_2969);
nand U7185 (N_7185,N_4101,N_4825);
nand U7186 (N_7186,N_4195,N_3632);
nor U7187 (N_7187,N_4949,N_3905);
nor U7188 (N_7188,N_4252,N_4645);
nand U7189 (N_7189,N_4518,N_3984);
and U7190 (N_7190,N_3807,N_2528);
nor U7191 (N_7191,N_3913,N_4307);
nor U7192 (N_7192,N_3523,N_2536);
xor U7193 (N_7193,N_4527,N_4178);
and U7194 (N_7194,N_4206,N_4267);
or U7195 (N_7195,N_3230,N_3363);
nor U7196 (N_7196,N_4834,N_3137);
nand U7197 (N_7197,N_3727,N_3119);
nor U7198 (N_7198,N_3236,N_4396);
and U7199 (N_7199,N_3679,N_3808);
nand U7200 (N_7200,N_4006,N_2967);
nand U7201 (N_7201,N_3373,N_4858);
or U7202 (N_7202,N_3159,N_4907);
nor U7203 (N_7203,N_4499,N_4796);
and U7204 (N_7204,N_4482,N_3298);
or U7205 (N_7205,N_4709,N_3826);
and U7206 (N_7206,N_3648,N_3348);
nand U7207 (N_7207,N_3933,N_2608);
or U7208 (N_7208,N_3507,N_4557);
nor U7209 (N_7209,N_2831,N_4797);
nand U7210 (N_7210,N_3518,N_4308);
nand U7211 (N_7211,N_4176,N_3035);
nor U7212 (N_7212,N_4569,N_4484);
or U7213 (N_7213,N_4298,N_2764);
and U7214 (N_7214,N_3340,N_2528);
nor U7215 (N_7215,N_4794,N_3727);
or U7216 (N_7216,N_2543,N_4418);
nand U7217 (N_7217,N_4585,N_4399);
and U7218 (N_7218,N_4083,N_4231);
or U7219 (N_7219,N_4601,N_4348);
nor U7220 (N_7220,N_3072,N_4126);
xor U7221 (N_7221,N_3929,N_4227);
nand U7222 (N_7222,N_3801,N_4901);
nand U7223 (N_7223,N_2886,N_4075);
nand U7224 (N_7224,N_3339,N_2825);
nor U7225 (N_7225,N_4592,N_4636);
or U7226 (N_7226,N_2677,N_4184);
or U7227 (N_7227,N_2893,N_4279);
xor U7228 (N_7228,N_4714,N_2862);
or U7229 (N_7229,N_3773,N_3922);
xor U7230 (N_7230,N_4184,N_4606);
and U7231 (N_7231,N_3403,N_2509);
nand U7232 (N_7232,N_2829,N_2757);
or U7233 (N_7233,N_2982,N_3138);
and U7234 (N_7234,N_3521,N_4478);
nand U7235 (N_7235,N_2528,N_3067);
or U7236 (N_7236,N_2712,N_4532);
or U7237 (N_7237,N_4855,N_4474);
nand U7238 (N_7238,N_2969,N_3764);
nand U7239 (N_7239,N_3980,N_4620);
nand U7240 (N_7240,N_3329,N_3012);
nor U7241 (N_7241,N_2595,N_4754);
and U7242 (N_7242,N_3136,N_4873);
or U7243 (N_7243,N_3304,N_3177);
nor U7244 (N_7244,N_4081,N_3717);
or U7245 (N_7245,N_3673,N_4371);
or U7246 (N_7246,N_4745,N_4900);
and U7247 (N_7247,N_3327,N_3267);
nor U7248 (N_7248,N_4161,N_3601);
nand U7249 (N_7249,N_4175,N_4361);
nor U7250 (N_7250,N_4681,N_3751);
or U7251 (N_7251,N_4604,N_3039);
nand U7252 (N_7252,N_2504,N_4024);
nor U7253 (N_7253,N_4663,N_4510);
nor U7254 (N_7254,N_4666,N_2515);
nand U7255 (N_7255,N_2906,N_4115);
and U7256 (N_7256,N_4734,N_4604);
and U7257 (N_7257,N_4384,N_4764);
nand U7258 (N_7258,N_4324,N_4901);
and U7259 (N_7259,N_2854,N_3339);
and U7260 (N_7260,N_2789,N_4036);
nor U7261 (N_7261,N_2633,N_3351);
or U7262 (N_7262,N_3129,N_4037);
and U7263 (N_7263,N_4490,N_4130);
nand U7264 (N_7264,N_4076,N_2775);
nor U7265 (N_7265,N_4717,N_2525);
nor U7266 (N_7266,N_3802,N_3974);
or U7267 (N_7267,N_3353,N_4463);
or U7268 (N_7268,N_4382,N_4622);
or U7269 (N_7269,N_4135,N_4307);
nand U7270 (N_7270,N_4548,N_4977);
nand U7271 (N_7271,N_4437,N_2614);
nand U7272 (N_7272,N_4053,N_4794);
or U7273 (N_7273,N_4821,N_3151);
and U7274 (N_7274,N_4830,N_4228);
nor U7275 (N_7275,N_4106,N_3185);
nand U7276 (N_7276,N_2520,N_4530);
or U7277 (N_7277,N_2595,N_3748);
nor U7278 (N_7278,N_2761,N_4818);
or U7279 (N_7279,N_3929,N_3706);
nand U7280 (N_7280,N_3905,N_2668);
nand U7281 (N_7281,N_4960,N_4449);
nand U7282 (N_7282,N_3583,N_2900);
or U7283 (N_7283,N_4638,N_2520);
and U7284 (N_7284,N_4570,N_2555);
or U7285 (N_7285,N_2738,N_2989);
nor U7286 (N_7286,N_3476,N_2519);
nor U7287 (N_7287,N_2705,N_4271);
nor U7288 (N_7288,N_4019,N_3861);
or U7289 (N_7289,N_4001,N_4339);
and U7290 (N_7290,N_2620,N_3951);
nand U7291 (N_7291,N_3016,N_2688);
and U7292 (N_7292,N_4508,N_4027);
nor U7293 (N_7293,N_4710,N_4478);
nor U7294 (N_7294,N_2961,N_3520);
nor U7295 (N_7295,N_3692,N_3536);
xnor U7296 (N_7296,N_4065,N_4849);
or U7297 (N_7297,N_4015,N_3964);
and U7298 (N_7298,N_3341,N_3027);
nor U7299 (N_7299,N_4720,N_3546);
nand U7300 (N_7300,N_4846,N_4313);
and U7301 (N_7301,N_4174,N_4992);
and U7302 (N_7302,N_3558,N_3437);
nand U7303 (N_7303,N_2703,N_2981);
and U7304 (N_7304,N_2581,N_3849);
xor U7305 (N_7305,N_4973,N_4904);
nand U7306 (N_7306,N_4493,N_4562);
nor U7307 (N_7307,N_4885,N_3881);
and U7308 (N_7308,N_3208,N_3957);
xor U7309 (N_7309,N_3443,N_3368);
nor U7310 (N_7310,N_3261,N_3129);
nor U7311 (N_7311,N_3449,N_4463);
nand U7312 (N_7312,N_4509,N_2523);
or U7313 (N_7313,N_3118,N_3756);
and U7314 (N_7314,N_4833,N_4422);
xor U7315 (N_7315,N_4113,N_3908);
and U7316 (N_7316,N_4882,N_3757);
nand U7317 (N_7317,N_4807,N_3321);
nand U7318 (N_7318,N_4066,N_4261);
and U7319 (N_7319,N_4803,N_4072);
nand U7320 (N_7320,N_3467,N_3665);
and U7321 (N_7321,N_3257,N_3523);
or U7322 (N_7322,N_3891,N_2518);
nor U7323 (N_7323,N_4681,N_3558);
or U7324 (N_7324,N_2927,N_3292);
or U7325 (N_7325,N_4373,N_4335);
or U7326 (N_7326,N_4161,N_4694);
or U7327 (N_7327,N_3633,N_3052);
and U7328 (N_7328,N_4075,N_3541);
nand U7329 (N_7329,N_4016,N_4477);
and U7330 (N_7330,N_4561,N_3829);
nor U7331 (N_7331,N_4663,N_3235);
nor U7332 (N_7332,N_3410,N_2982);
nand U7333 (N_7333,N_4268,N_2910);
xnor U7334 (N_7334,N_2996,N_4958);
nor U7335 (N_7335,N_2765,N_2791);
and U7336 (N_7336,N_3599,N_4162);
or U7337 (N_7337,N_3736,N_3421);
nand U7338 (N_7338,N_4460,N_2867);
nand U7339 (N_7339,N_4217,N_4637);
nor U7340 (N_7340,N_4332,N_4204);
and U7341 (N_7341,N_3481,N_4718);
nor U7342 (N_7342,N_3699,N_4824);
and U7343 (N_7343,N_3367,N_2849);
or U7344 (N_7344,N_4918,N_3132);
and U7345 (N_7345,N_4543,N_4856);
and U7346 (N_7346,N_4162,N_4452);
nor U7347 (N_7347,N_4889,N_3616);
nand U7348 (N_7348,N_2570,N_4744);
nand U7349 (N_7349,N_3345,N_3102);
nor U7350 (N_7350,N_3298,N_4081);
nor U7351 (N_7351,N_4192,N_3002);
and U7352 (N_7352,N_4399,N_3417);
nand U7353 (N_7353,N_4272,N_4869);
and U7354 (N_7354,N_3628,N_3368);
and U7355 (N_7355,N_4189,N_4414);
or U7356 (N_7356,N_4892,N_4824);
or U7357 (N_7357,N_2752,N_3220);
and U7358 (N_7358,N_2955,N_2607);
or U7359 (N_7359,N_3466,N_2505);
nor U7360 (N_7360,N_3142,N_3977);
and U7361 (N_7361,N_2796,N_3784);
or U7362 (N_7362,N_2809,N_4046);
or U7363 (N_7363,N_3659,N_3376);
nand U7364 (N_7364,N_3397,N_3548);
and U7365 (N_7365,N_3284,N_3189);
nor U7366 (N_7366,N_4780,N_2724);
nand U7367 (N_7367,N_4284,N_3442);
and U7368 (N_7368,N_4277,N_3957);
or U7369 (N_7369,N_4442,N_3866);
or U7370 (N_7370,N_3756,N_4093);
nor U7371 (N_7371,N_4624,N_4446);
and U7372 (N_7372,N_3518,N_3487);
nor U7373 (N_7373,N_4020,N_2822);
nand U7374 (N_7374,N_3106,N_3019);
nand U7375 (N_7375,N_3764,N_4489);
xnor U7376 (N_7376,N_2959,N_3105);
or U7377 (N_7377,N_4507,N_3314);
nand U7378 (N_7378,N_2865,N_2775);
or U7379 (N_7379,N_3562,N_3623);
nor U7380 (N_7380,N_4654,N_4612);
nor U7381 (N_7381,N_3459,N_4517);
nor U7382 (N_7382,N_3800,N_2809);
nand U7383 (N_7383,N_4146,N_3353);
and U7384 (N_7384,N_4693,N_4499);
and U7385 (N_7385,N_3729,N_2971);
or U7386 (N_7386,N_2558,N_3019);
nor U7387 (N_7387,N_2504,N_4934);
or U7388 (N_7388,N_3797,N_3952);
nand U7389 (N_7389,N_4568,N_2896);
and U7390 (N_7390,N_2959,N_4978);
nor U7391 (N_7391,N_4504,N_4843);
and U7392 (N_7392,N_3668,N_3267);
or U7393 (N_7393,N_2613,N_4889);
or U7394 (N_7394,N_4119,N_4296);
nor U7395 (N_7395,N_4992,N_3836);
nor U7396 (N_7396,N_3441,N_4136);
nor U7397 (N_7397,N_4306,N_3105);
or U7398 (N_7398,N_4932,N_3704);
and U7399 (N_7399,N_3108,N_3105);
and U7400 (N_7400,N_3952,N_4036);
or U7401 (N_7401,N_3403,N_3708);
nand U7402 (N_7402,N_2698,N_2580);
nand U7403 (N_7403,N_4014,N_3386);
and U7404 (N_7404,N_3432,N_2733);
nor U7405 (N_7405,N_4444,N_4165);
nand U7406 (N_7406,N_2507,N_2926);
nor U7407 (N_7407,N_2865,N_3231);
nor U7408 (N_7408,N_3037,N_4689);
and U7409 (N_7409,N_4887,N_4382);
nor U7410 (N_7410,N_4110,N_4602);
nor U7411 (N_7411,N_3424,N_4296);
and U7412 (N_7412,N_4697,N_3194);
nor U7413 (N_7413,N_3558,N_2704);
or U7414 (N_7414,N_3089,N_4586);
nor U7415 (N_7415,N_3926,N_3201);
or U7416 (N_7416,N_3988,N_2766);
nand U7417 (N_7417,N_4239,N_4890);
nor U7418 (N_7418,N_4260,N_4725);
and U7419 (N_7419,N_3349,N_2973);
nand U7420 (N_7420,N_4343,N_3802);
nand U7421 (N_7421,N_3189,N_4258);
and U7422 (N_7422,N_2836,N_3134);
or U7423 (N_7423,N_3721,N_4122);
nand U7424 (N_7424,N_4095,N_4937);
or U7425 (N_7425,N_4285,N_4245);
nand U7426 (N_7426,N_3738,N_3208);
nor U7427 (N_7427,N_4978,N_2555);
nand U7428 (N_7428,N_3106,N_4929);
and U7429 (N_7429,N_4490,N_4527);
nand U7430 (N_7430,N_3337,N_3114);
nor U7431 (N_7431,N_3719,N_3238);
nor U7432 (N_7432,N_3097,N_4693);
or U7433 (N_7433,N_4852,N_2783);
nor U7434 (N_7434,N_3665,N_2500);
nand U7435 (N_7435,N_3135,N_4331);
or U7436 (N_7436,N_4884,N_2687);
and U7437 (N_7437,N_2538,N_3928);
xor U7438 (N_7438,N_4315,N_3554);
or U7439 (N_7439,N_4236,N_4847);
nand U7440 (N_7440,N_4801,N_3334);
nor U7441 (N_7441,N_3504,N_3213);
or U7442 (N_7442,N_3825,N_3011);
nand U7443 (N_7443,N_4314,N_3391);
and U7444 (N_7444,N_3880,N_3511);
and U7445 (N_7445,N_4446,N_3025);
nand U7446 (N_7446,N_3044,N_3747);
and U7447 (N_7447,N_4646,N_4721);
nand U7448 (N_7448,N_3900,N_4996);
xor U7449 (N_7449,N_4290,N_3790);
nor U7450 (N_7450,N_4753,N_2533);
nor U7451 (N_7451,N_2917,N_3990);
nand U7452 (N_7452,N_3823,N_4902);
or U7453 (N_7453,N_2550,N_3847);
nand U7454 (N_7454,N_4026,N_3664);
nor U7455 (N_7455,N_4450,N_3631);
or U7456 (N_7456,N_2592,N_2915);
nand U7457 (N_7457,N_3510,N_3267);
nand U7458 (N_7458,N_4823,N_3320);
nand U7459 (N_7459,N_3164,N_2671);
or U7460 (N_7460,N_4362,N_4663);
or U7461 (N_7461,N_3830,N_3883);
and U7462 (N_7462,N_4776,N_3556);
or U7463 (N_7463,N_3411,N_3313);
or U7464 (N_7464,N_4826,N_3924);
nand U7465 (N_7465,N_3800,N_4775);
nor U7466 (N_7466,N_3341,N_2746);
and U7467 (N_7467,N_4058,N_3498);
nand U7468 (N_7468,N_2597,N_3032);
or U7469 (N_7469,N_3627,N_4404);
nand U7470 (N_7470,N_3843,N_4849);
and U7471 (N_7471,N_4106,N_4485);
and U7472 (N_7472,N_4967,N_3744);
nor U7473 (N_7473,N_3105,N_3708);
nor U7474 (N_7474,N_3949,N_2727);
and U7475 (N_7475,N_2770,N_3828);
or U7476 (N_7476,N_3914,N_3654);
or U7477 (N_7477,N_3768,N_3688);
nand U7478 (N_7478,N_3176,N_3028);
nand U7479 (N_7479,N_2557,N_2771);
nand U7480 (N_7480,N_3248,N_4118);
and U7481 (N_7481,N_2958,N_4445);
or U7482 (N_7482,N_3247,N_4564);
nor U7483 (N_7483,N_4266,N_4023);
or U7484 (N_7484,N_3230,N_2692);
and U7485 (N_7485,N_4791,N_3984);
nand U7486 (N_7486,N_4470,N_2984);
and U7487 (N_7487,N_4228,N_3519);
or U7488 (N_7488,N_4666,N_3229);
nor U7489 (N_7489,N_4204,N_4441);
nand U7490 (N_7490,N_2807,N_4615);
nor U7491 (N_7491,N_3200,N_2597);
and U7492 (N_7492,N_4078,N_2657);
nand U7493 (N_7493,N_4158,N_4604);
nand U7494 (N_7494,N_3485,N_3219);
nand U7495 (N_7495,N_3115,N_4483);
nor U7496 (N_7496,N_2936,N_4150);
or U7497 (N_7497,N_3965,N_3830);
and U7498 (N_7498,N_3152,N_3405);
nor U7499 (N_7499,N_4593,N_3611);
or U7500 (N_7500,N_5133,N_5884);
nor U7501 (N_7501,N_6119,N_7004);
or U7502 (N_7502,N_5604,N_5638);
and U7503 (N_7503,N_5701,N_5451);
nor U7504 (N_7504,N_6317,N_5605);
or U7505 (N_7505,N_7247,N_7021);
or U7506 (N_7506,N_6356,N_5693);
nand U7507 (N_7507,N_6035,N_6655);
nor U7508 (N_7508,N_5428,N_5396);
nor U7509 (N_7509,N_6355,N_6742);
or U7510 (N_7510,N_7009,N_6756);
nand U7511 (N_7511,N_5808,N_6115);
and U7512 (N_7512,N_5768,N_5060);
or U7513 (N_7513,N_7163,N_5885);
or U7514 (N_7514,N_5826,N_7197);
nor U7515 (N_7515,N_7136,N_6582);
nor U7516 (N_7516,N_6164,N_6599);
or U7517 (N_7517,N_7262,N_5002);
or U7518 (N_7518,N_6306,N_7268);
nor U7519 (N_7519,N_7455,N_6628);
nand U7520 (N_7520,N_6762,N_6764);
or U7521 (N_7521,N_5890,N_7030);
nand U7522 (N_7522,N_6406,N_6022);
nor U7523 (N_7523,N_6825,N_7075);
or U7524 (N_7524,N_6382,N_7410);
or U7525 (N_7525,N_6358,N_6235);
nor U7526 (N_7526,N_6814,N_6052);
nand U7527 (N_7527,N_5508,N_6280);
and U7528 (N_7528,N_6697,N_6917);
and U7529 (N_7529,N_5365,N_5243);
and U7530 (N_7530,N_6156,N_7063);
or U7531 (N_7531,N_5104,N_6525);
or U7532 (N_7532,N_6696,N_6441);
nor U7533 (N_7533,N_6163,N_5953);
or U7534 (N_7534,N_6794,N_5470);
nand U7535 (N_7535,N_5718,N_6899);
or U7536 (N_7536,N_6617,N_7167);
nand U7537 (N_7537,N_6070,N_5902);
nor U7538 (N_7538,N_7064,N_5454);
and U7539 (N_7539,N_5027,N_5386);
or U7540 (N_7540,N_5651,N_6621);
nand U7541 (N_7541,N_5753,N_6836);
or U7542 (N_7542,N_6574,N_7202);
nand U7543 (N_7543,N_7470,N_5210);
nor U7544 (N_7544,N_6955,N_6593);
nor U7545 (N_7545,N_7036,N_6481);
nand U7546 (N_7546,N_7329,N_6694);
or U7547 (N_7547,N_5230,N_5769);
or U7548 (N_7548,N_5437,N_7111);
nor U7549 (N_7549,N_6568,N_5917);
nor U7550 (N_7550,N_6654,N_5945);
or U7551 (N_7551,N_6649,N_6321);
and U7552 (N_7552,N_6790,N_6201);
nand U7553 (N_7553,N_7284,N_5053);
or U7554 (N_7554,N_6660,N_6688);
or U7555 (N_7555,N_5786,N_6240);
and U7556 (N_7556,N_6592,N_7298);
or U7557 (N_7557,N_5240,N_6606);
nand U7558 (N_7558,N_6630,N_7311);
and U7559 (N_7559,N_6989,N_5985);
and U7560 (N_7560,N_5780,N_7142);
or U7561 (N_7561,N_5936,N_7144);
and U7562 (N_7562,N_5996,N_6904);
and U7563 (N_7563,N_7193,N_7319);
and U7564 (N_7564,N_5533,N_5477);
or U7565 (N_7565,N_6369,N_6155);
or U7566 (N_7566,N_5267,N_5789);
and U7567 (N_7567,N_6613,N_6906);
or U7568 (N_7568,N_5337,N_5379);
nand U7569 (N_7569,N_5655,N_7289);
and U7570 (N_7570,N_6449,N_5859);
and U7571 (N_7571,N_5233,N_7133);
nor U7572 (N_7572,N_5022,N_5727);
or U7573 (N_7573,N_7198,N_6859);
nor U7574 (N_7574,N_5755,N_6819);
nand U7575 (N_7575,N_5515,N_6512);
nand U7576 (N_7576,N_5375,N_6007);
nor U7577 (N_7577,N_5903,N_6982);
and U7578 (N_7578,N_5654,N_6934);
and U7579 (N_7579,N_6507,N_6735);
and U7580 (N_7580,N_6937,N_6784);
nand U7581 (N_7581,N_7043,N_6516);
nor U7582 (N_7582,N_5207,N_6097);
nor U7583 (N_7583,N_6184,N_7466);
nor U7584 (N_7584,N_6571,N_5648);
nor U7585 (N_7585,N_5328,N_7322);
and U7586 (N_7586,N_6996,N_5523);
or U7587 (N_7587,N_6653,N_7290);
nor U7588 (N_7588,N_7353,N_7074);
or U7589 (N_7589,N_7234,N_7086);
and U7590 (N_7590,N_6307,N_6731);
nor U7591 (N_7591,N_5425,N_6898);
and U7592 (N_7592,N_6840,N_7345);
nor U7593 (N_7593,N_5711,N_5958);
nand U7594 (N_7594,N_6259,N_6948);
and U7595 (N_7595,N_5620,N_6960);
and U7596 (N_7596,N_7259,N_6393);
and U7597 (N_7597,N_5181,N_5819);
and U7598 (N_7598,N_7215,N_6602);
or U7599 (N_7599,N_7393,N_6009);
nor U7600 (N_7600,N_6849,N_5406);
xnor U7601 (N_7601,N_6487,N_6206);
nand U7602 (N_7602,N_6505,N_7286);
and U7603 (N_7603,N_6277,N_5463);
and U7604 (N_7604,N_5736,N_6504);
or U7605 (N_7605,N_7467,N_6730);
and U7606 (N_7606,N_5992,N_7294);
nand U7607 (N_7607,N_7309,N_6792);
and U7608 (N_7608,N_5586,N_6074);
and U7609 (N_7609,N_6572,N_6413);
nor U7610 (N_7610,N_5626,N_6554);
or U7611 (N_7611,N_5566,N_7317);
or U7612 (N_7612,N_6919,N_6608);
nand U7613 (N_7613,N_7204,N_6539);
and U7614 (N_7614,N_6202,N_7464);
or U7615 (N_7615,N_5719,N_7090);
nor U7616 (N_7616,N_5969,N_5733);
nor U7617 (N_7617,N_7417,N_5762);
and U7618 (N_7618,N_6807,N_5290);
and U7619 (N_7619,N_5169,N_5025);
and U7620 (N_7620,N_6530,N_7060);
or U7621 (N_7621,N_5201,N_5632);
nand U7622 (N_7622,N_6935,N_5645);
or U7623 (N_7623,N_5547,N_6026);
and U7624 (N_7624,N_5834,N_6242);
and U7625 (N_7625,N_6652,N_7423);
and U7626 (N_7626,N_6172,N_7295);
and U7627 (N_7627,N_6800,N_5549);
or U7628 (N_7628,N_6222,N_7052);
nor U7629 (N_7629,N_7368,N_7229);
nand U7630 (N_7630,N_5561,N_6336);
nor U7631 (N_7631,N_6778,N_5976);
nor U7632 (N_7632,N_6152,N_5670);
nor U7633 (N_7633,N_6204,N_5756);
nand U7634 (N_7634,N_6331,N_7121);
nor U7635 (N_7635,N_7443,N_6651);
or U7636 (N_7636,N_5657,N_5828);
and U7637 (N_7637,N_5731,N_5042);
or U7638 (N_7638,N_5524,N_5007);
nand U7639 (N_7639,N_7428,N_6123);
nand U7640 (N_7640,N_5511,N_6057);
nor U7641 (N_7641,N_7475,N_5617);
nor U7642 (N_7642,N_6466,N_6815);
or U7643 (N_7643,N_6671,N_5000);
nand U7644 (N_7644,N_6169,N_5935);
nand U7645 (N_7645,N_5710,N_5125);
or U7646 (N_7646,N_7492,N_6526);
nor U7647 (N_7647,N_7025,N_7184);
nor U7648 (N_7648,N_6085,N_5389);
or U7649 (N_7649,N_7477,N_6011);
and U7650 (N_7650,N_7321,N_5841);
nor U7651 (N_7651,N_6001,N_5446);
or U7652 (N_7652,N_7178,N_6820);
nor U7653 (N_7653,N_7478,N_6460);
and U7654 (N_7654,N_7152,N_5244);
and U7655 (N_7655,N_6159,N_7331);
and U7656 (N_7656,N_6214,N_6179);
nand U7657 (N_7657,N_6839,N_6462);
or U7658 (N_7658,N_7489,N_5286);
or U7659 (N_7659,N_6886,N_6589);
and U7660 (N_7660,N_6618,N_6439);
nor U7661 (N_7661,N_5715,N_6863);
and U7662 (N_7662,N_7413,N_7397);
or U7663 (N_7663,N_5799,N_5732);
or U7664 (N_7664,N_7062,N_5362);
nand U7665 (N_7665,N_6028,N_5058);
nand U7666 (N_7666,N_5905,N_7399);
nor U7667 (N_7667,N_5581,N_6048);
and U7668 (N_7668,N_5616,N_6348);
nand U7669 (N_7669,N_7304,N_6707);
and U7670 (N_7670,N_5019,N_6344);
nor U7671 (N_7671,N_6146,N_6584);
nand U7672 (N_7672,N_5564,N_6230);
nor U7673 (N_7673,N_6614,N_6729);
nor U7674 (N_7674,N_5268,N_6434);
and U7675 (N_7675,N_6623,N_6997);
and U7676 (N_7676,N_5920,N_7186);
nor U7677 (N_7677,N_6973,N_6485);
or U7678 (N_7678,N_6737,N_6661);
nand U7679 (N_7679,N_5551,N_5763);
and U7680 (N_7680,N_6875,N_5873);
or U7681 (N_7681,N_6409,N_6289);
or U7682 (N_7682,N_7388,N_7446);
or U7683 (N_7683,N_5138,N_5330);
nand U7684 (N_7684,N_7491,N_6368);
nor U7685 (N_7685,N_5127,N_6698);
or U7686 (N_7686,N_5229,N_6263);
nor U7687 (N_7687,N_6767,N_5975);
nor U7688 (N_7688,N_5737,N_7211);
and U7689 (N_7689,N_5813,N_5827);
or U7690 (N_7690,N_7285,N_7291);
nand U7691 (N_7691,N_6685,N_5713);
nand U7692 (N_7692,N_5795,N_6797);
or U7693 (N_7693,N_6573,N_7131);
and U7694 (N_7694,N_6290,N_6776);
or U7695 (N_7695,N_7320,N_7155);
nand U7696 (N_7696,N_5539,N_6157);
and U7697 (N_7697,N_5583,N_5045);
nand U7698 (N_7698,N_5745,N_7409);
or U7699 (N_7699,N_7046,N_6012);
and U7700 (N_7700,N_6076,N_5948);
nand U7701 (N_7701,N_6940,N_6719);
nand U7702 (N_7702,N_7253,N_5298);
xnor U7703 (N_7703,N_6471,N_6780);
and U7704 (N_7704,N_6446,N_6639);
and U7705 (N_7705,N_6093,N_6284);
and U7706 (N_7706,N_5248,N_5754);
and U7707 (N_7707,N_7391,N_6394);
nand U7708 (N_7708,N_7348,N_7208);
and U7709 (N_7709,N_7244,N_5987);
nor U7710 (N_7710,N_6086,N_6850);
or U7711 (N_7711,N_6082,N_6665);
nand U7712 (N_7712,N_6787,N_5531);
and U7713 (N_7713,N_5923,N_7263);
and U7714 (N_7714,N_5792,N_6650);
nand U7715 (N_7715,N_7182,N_5692);
and U7716 (N_7716,N_7402,N_5944);
nor U7717 (N_7717,N_5722,N_5724);
and U7718 (N_7718,N_5874,N_6219);
or U7719 (N_7719,N_6761,N_5650);
or U7720 (N_7720,N_6854,N_6347);
or U7721 (N_7721,N_7306,N_5770);
and U7722 (N_7722,N_6956,N_7436);
or U7723 (N_7723,N_6842,N_7269);
nand U7724 (N_7724,N_5664,N_5788);
nand U7725 (N_7725,N_6153,N_7305);
nand U7726 (N_7726,N_5642,N_6049);
nor U7727 (N_7727,N_7481,N_5822);
and U7728 (N_7728,N_5590,N_6486);
or U7729 (N_7729,N_5319,N_5351);
and U7730 (N_7730,N_5610,N_5276);
nor U7731 (N_7731,N_6084,N_7378);
and U7732 (N_7732,N_6588,N_6817);
nor U7733 (N_7733,N_5155,N_7217);
nand U7734 (N_7734,N_5047,N_6978);
and U7735 (N_7735,N_6136,N_6553);
nand U7736 (N_7736,N_5546,N_5618);
nand U7737 (N_7737,N_5906,N_6773);
nor U7738 (N_7738,N_5501,N_6869);
nand U7739 (N_7739,N_7139,N_7112);
and U7740 (N_7740,N_5123,N_6490);
or U7741 (N_7741,N_6705,N_6432);
and U7742 (N_7742,N_5507,N_6522);
and U7743 (N_7743,N_5708,N_6734);
or U7744 (N_7744,N_5085,N_5333);
or U7745 (N_7745,N_6912,N_7314);
or U7746 (N_7746,N_7313,N_6519);
or U7747 (N_7747,N_5236,N_5823);
and U7748 (N_7748,N_5101,N_6351);
or U7749 (N_7749,N_5339,N_6689);
and U7750 (N_7750,N_5812,N_5052);
nor U7751 (N_7751,N_5177,N_7038);
or U7752 (N_7752,N_6081,N_6226);
nor U7753 (N_7753,N_7016,N_6619);
nor U7754 (N_7754,N_7199,N_5356);
nand U7755 (N_7755,N_6502,N_7071);
nand U7756 (N_7756,N_6562,N_6598);
nor U7757 (N_7757,N_5141,N_6291);
and U7758 (N_7758,N_6852,N_5416);
nand U7759 (N_7759,N_7218,N_6712);
and U7760 (N_7760,N_5439,N_7355);
and U7761 (N_7761,N_5432,N_7343);
and U7762 (N_7762,N_6129,N_6806);
nor U7763 (N_7763,N_6830,N_5904);
or U7764 (N_7764,N_5647,N_5496);
or U7765 (N_7765,N_5679,N_7376);
or U7766 (N_7766,N_7073,N_7001);
nand U7767 (N_7767,N_6835,N_5017);
xnor U7768 (N_7768,N_5352,N_5126);
and U7769 (N_7769,N_6957,N_5204);
nor U7770 (N_7770,N_7245,N_5311);
nor U7771 (N_7771,N_5185,N_5553);
xor U7772 (N_7772,N_5621,N_5166);
nor U7773 (N_7773,N_5223,N_6895);
or U7774 (N_7774,N_5237,N_5440);
nand U7775 (N_7775,N_6452,N_6103);
nor U7776 (N_7776,N_6386,N_7404);
nand U7777 (N_7777,N_6838,N_5609);
nand U7778 (N_7778,N_5306,N_6828);
or U7779 (N_7779,N_6110,N_5012);
or U7780 (N_7780,N_5594,N_7130);
and U7781 (N_7781,N_6322,N_6491);
or U7782 (N_7782,N_7473,N_5269);
and U7783 (N_7783,N_7371,N_6333);
and U7784 (N_7784,N_5039,N_5915);
or U7785 (N_7785,N_6569,N_7049);
xnor U7786 (N_7786,N_7354,N_7179);
nand U7787 (N_7787,N_6044,N_6175);
or U7788 (N_7788,N_6856,N_5433);
or U7789 (N_7789,N_6758,N_6751);
or U7790 (N_7790,N_5738,N_7087);
nand U7791 (N_7791,N_6664,N_7496);
or U7792 (N_7792,N_5317,N_6861);
and U7793 (N_7793,N_5111,N_7469);
and U7794 (N_7794,N_5238,N_6594);
nand U7795 (N_7795,N_6788,N_7141);
and U7796 (N_7796,N_6745,N_5213);
and U7797 (N_7797,N_5301,N_5212);
nor U7798 (N_7798,N_6190,N_6922);
nor U7799 (N_7799,N_5080,N_5649);
nor U7800 (N_7800,N_7093,N_7479);
and U7801 (N_7801,N_6565,N_5599);
nor U7802 (N_7802,N_5336,N_5790);
nand U7803 (N_7803,N_6804,N_6752);
nand U7804 (N_7804,N_5931,N_6677);
or U7805 (N_7805,N_5335,N_5965);
nor U7806 (N_7806,N_5993,N_5695);
nor U7807 (N_7807,N_6559,N_5461);
nand U7808 (N_7808,N_6943,N_7113);
and U7809 (N_7809,N_5982,N_5354);
or U7810 (N_7810,N_5807,N_6031);
nand U7811 (N_7811,N_5926,N_6073);
or U7812 (N_7812,N_5704,N_7497);
or U7813 (N_7813,N_6603,N_6892);
nor U7814 (N_7814,N_5305,N_7293);
and U7815 (N_7815,N_6278,N_5438);
and U7816 (N_7816,N_6120,N_5102);
and U7817 (N_7817,N_5054,N_5999);
and U7818 (N_7818,N_6902,N_7107);
and U7819 (N_7819,N_7084,N_5436);
nor U7820 (N_7820,N_5488,N_6400);
nor U7821 (N_7821,N_5146,N_5264);
nand U7822 (N_7822,N_6942,N_6475);
nor U7823 (N_7823,N_7239,N_5684);
nor U7824 (N_7824,N_7002,N_5625);
and U7825 (N_7825,N_6037,N_6670);
nor U7826 (N_7826,N_5259,N_5689);
and U7827 (N_7827,N_7027,N_5313);
and U7828 (N_7828,N_6888,N_6139);
nor U7829 (N_7829,N_7173,N_5830);
and U7830 (N_7830,N_6071,N_5459);
nand U7831 (N_7831,N_6265,N_6221);
and U7832 (N_7832,N_6102,N_7108);
nand U7833 (N_7833,N_5779,N_6450);
and U7834 (N_7834,N_6189,N_5287);
and U7835 (N_7835,N_7308,N_5500);
nand U7836 (N_7836,N_5803,N_6744);
and U7837 (N_7837,N_6959,N_5631);
or U7838 (N_7838,N_5653,N_5750);
nor U7839 (N_7839,N_6601,N_6061);
or U7840 (N_7840,N_5940,N_6312);
nand U7841 (N_7841,N_6018,N_6469);
or U7842 (N_7842,N_5815,N_7260);
nor U7843 (N_7843,N_6845,N_7273);
or U7844 (N_7844,N_5140,N_7254);
and U7845 (N_7845,N_6273,N_7316);
xnor U7846 (N_7846,N_6117,N_6437);
or U7847 (N_7847,N_5744,N_7424);
or U7848 (N_7848,N_6669,N_5797);
and U7849 (N_7849,N_6458,N_5189);
and U7850 (N_7850,N_7468,N_7080);
and U7851 (N_7851,N_5398,N_7408);
nor U7852 (N_7852,N_5748,N_5348);
or U7853 (N_7853,N_6045,N_5550);
nor U7854 (N_7854,N_5282,N_7437);
and U7855 (N_7855,N_7257,N_5124);
and U7856 (N_7856,N_6241,N_7120);
and U7857 (N_7857,N_5876,N_6233);
and U7858 (N_7858,N_5629,N_6950);
nand U7859 (N_7859,N_7126,N_7013);
nand U7860 (N_7860,N_6533,N_5573);
and U7861 (N_7861,N_5081,N_7041);
nand U7862 (N_7862,N_7281,N_5088);
nand U7863 (N_7863,N_5192,N_5558);
or U7864 (N_7864,N_6470,N_5014);
and U7865 (N_7865,N_5530,N_7237);
and U7866 (N_7866,N_5607,N_6676);
and U7867 (N_7867,N_6591,N_5005);
and U7868 (N_7868,N_6695,N_5899);
or U7869 (N_7869,N_5384,N_6821);
and U7870 (N_7870,N_6360,N_7207);
or U7871 (N_7871,N_5700,N_6337);
or U7872 (N_7872,N_7214,N_6126);
and U7873 (N_7873,N_5162,N_7008);
nand U7874 (N_7874,N_7159,N_7282);
or U7875 (N_7875,N_5209,N_6176);
and U7876 (N_7876,N_5656,N_6855);
nor U7877 (N_7877,N_5962,N_7264);
and U7878 (N_7878,N_7061,N_5278);
and U7879 (N_7879,N_5611,N_6443);
or U7880 (N_7880,N_5844,N_5382);
and U7881 (N_7881,N_6436,N_7056);
nand U7882 (N_7882,N_6447,N_6563);
nand U7883 (N_7883,N_5410,N_6638);
nor U7884 (N_7884,N_6124,N_6663);
or U7885 (N_7885,N_5893,N_6089);
or U7886 (N_7886,N_6033,N_5073);
or U7887 (N_7887,N_5293,N_5342);
nand U7888 (N_7888,N_5978,N_5911);
and U7889 (N_7889,N_7484,N_5036);
or U7890 (N_7890,N_6218,N_6193);
or U7891 (N_7891,N_5543,N_7267);
nand U7892 (N_7892,N_7082,N_6177);
and U7893 (N_7893,N_6112,N_6267);
and U7894 (N_7894,N_5652,N_7301);
and U7895 (N_7895,N_6472,N_6681);
and U7896 (N_7896,N_6182,N_7425);
or U7897 (N_7897,N_6805,N_6067);
or U7898 (N_7898,N_6027,N_5894);
or U7899 (N_7899,N_5215,N_5582);
nor U7900 (N_7900,N_5575,N_5570);
nand U7901 (N_7901,N_7377,N_6165);
nor U7902 (N_7902,N_6107,N_6923);
and U7903 (N_7903,N_5359,N_6596);
nand U7904 (N_7904,N_5746,N_7418);
nand U7905 (N_7905,N_5218,N_6298);
nor U7906 (N_7906,N_5688,N_6309);
and U7907 (N_7907,N_5691,N_5077);
or U7908 (N_7908,N_6227,N_5199);
and U7909 (N_7909,N_5071,N_5824);
and U7910 (N_7910,N_5775,N_7312);
nor U7911 (N_7911,N_5810,N_7138);
and U7912 (N_7912,N_6418,N_6738);
or U7913 (N_7913,N_5479,N_6520);
nor U7914 (N_7914,N_7325,N_6702);
nand U7915 (N_7915,N_5309,N_7185);
nor U7916 (N_7916,N_5341,N_7243);
or U7917 (N_7917,N_6144,N_5369);
nor U7918 (N_7918,N_5175,N_6812);
or U7919 (N_7919,N_5116,N_5499);
nand U7920 (N_7920,N_5989,N_5880);
nand U7921 (N_7921,N_6457,N_5951);
nand U7922 (N_7922,N_5697,N_5526);
nand U7923 (N_7923,N_5644,N_7300);
or U7924 (N_7924,N_5776,N_7297);
nand U7925 (N_7925,N_6397,N_6257);
or U7926 (N_7926,N_5947,N_6357);
nand U7927 (N_7927,N_5871,N_6476);
or U7928 (N_7928,N_5879,N_5661);
nand U7929 (N_7929,N_5514,N_5391);
nand U7930 (N_7930,N_6302,N_6166);
and U7931 (N_7931,N_5641,N_7118);
nand U7932 (N_7932,N_5933,N_7127);
nand U7933 (N_7933,N_7250,N_7122);
and U7934 (N_7934,N_5943,N_5430);
or U7935 (N_7935,N_5357,N_6410);
and U7936 (N_7936,N_6903,N_6867);
nor U7937 (N_7937,N_5971,N_7433);
nand U7938 (N_7938,N_5866,N_5739);
nand U7939 (N_7939,N_5404,N_5038);
or U7940 (N_7940,N_5308,N_7372);
nor U7941 (N_7941,N_7033,N_5453);
nand U7942 (N_7942,N_5318,N_5165);
nor U7943 (N_7943,N_5968,N_6316);
nand U7944 (N_7944,N_6170,N_6381);
and U7945 (N_7945,N_6104,N_7106);
nor U7946 (N_7946,N_5392,N_7438);
and U7947 (N_7947,N_6186,N_5628);
nor U7948 (N_7948,N_7369,N_6597);
nand U7949 (N_7949,N_5921,N_6438);
nor U7950 (N_7950,N_7176,N_5261);
or U7951 (N_7951,N_7145,N_6720);
nor U7952 (N_7952,N_6635,N_7441);
nor U7953 (N_7953,N_7089,N_7493);
or U7954 (N_7954,N_6249,N_5538);
nand U7955 (N_7955,N_6844,N_5100);
nand U7956 (N_7956,N_6367,N_5497);
nand U7957 (N_7957,N_6464,N_7482);
nor U7958 (N_7958,N_7092,N_5552);
or U7959 (N_7959,N_6423,N_5505);
nand U7960 (N_7960,N_5062,N_6180);
or U7961 (N_7961,N_6841,N_7488);
or U7962 (N_7962,N_5869,N_7318);
and U7963 (N_7963,N_5368,N_5272);
nor U7964 (N_7964,N_6557,N_7240);
and U7965 (N_7965,N_7209,N_5565);
and U7966 (N_7966,N_7006,N_5730);
and U7967 (N_7967,N_5990,N_5838);
nand U7968 (N_7968,N_6363,N_5672);
and U7969 (N_7969,N_6187,N_6640);
or U7970 (N_7970,N_6444,N_5856);
nand U7971 (N_7971,N_6748,N_6765);
nor U7972 (N_7972,N_5314,N_6154);
nand U7973 (N_7973,N_5250,N_5239);
and U7974 (N_7974,N_7037,N_7236);
or U7975 (N_7975,N_5984,N_6096);
nor U7976 (N_7976,N_6194,N_6105);
nor U7977 (N_7977,N_6605,N_6092);
nand U7978 (N_7978,N_5469,N_5134);
or U7979 (N_7979,N_7194,N_5429);
nor U7980 (N_7980,N_6951,N_5462);
or U7981 (N_7981,N_7005,N_5143);
nand U7982 (N_7982,N_6831,N_7485);
nor U7983 (N_7983,N_7261,N_6417);
and U7984 (N_7984,N_6142,N_5371);
nand U7985 (N_7985,N_7356,N_5145);
and U7986 (N_7986,N_6511,N_7200);
nand U7987 (N_7987,N_5928,N_5519);
or U7988 (N_7988,N_7022,N_6495);
nor U7989 (N_7989,N_7161,N_7249);
nor U7990 (N_7990,N_5271,N_7091);
or U7991 (N_7991,N_6286,N_6332);
or U7992 (N_7992,N_6723,N_6811);
nor U7993 (N_7993,N_7375,N_6134);
nand U7994 (N_7994,N_5242,N_5596);
or U7995 (N_7995,N_5850,N_6701);
or U7996 (N_7996,N_5414,N_6916);
nor U7997 (N_7997,N_5340,N_5296);
nor U7998 (N_7998,N_6258,N_6775);
or U7999 (N_7999,N_7123,N_6217);
and U8000 (N_8000,N_5279,N_6733);
and U8001 (N_8001,N_5343,N_5646);
nand U8002 (N_8002,N_5774,N_7232);
and U8003 (N_8003,N_6006,N_5316);
and U8004 (N_8004,N_5970,N_5929);
or U8005 (N_8005,N_6900,N_7109);
and U8006 (N_8006,N_5108,N_5484);
nand U8007 (N_8007,N_5481,N_5633);
or U8008 (N_8008,N_5562,N_5323);
or U8009 (N_8009,N_6576,N_6883);
or U8010 (N_8010,N_5709,N_5128);
or U8011 (N_8011,N_7432,N_6209);
and U8012 (N_8012,N_5798,N_5280);
or U8013 (N_8013,N_5941,N_6319);
or U8014 (N_8014,N_5387,N_5800);
or U8015 (N_8015,N_5498,N_7117);
or U8016 (N_8016,N_6891,N_5092);
nand U8017 (N_8017,N_6580,N_5112);
or U8018 (N_8018,N_5955,N_7116);
or U8019 (N_8019,N_6150,N_6497);
or U8020 (N_8020,N_6551,N_6931);
and U8021 (N_8021,N_7058,N_6188);
nor U8022 (N_8022,N_6459,N_6678);
or U8023 (N_8023,N_6637,N_7334);
nor U8024 (N_8024,N_5435,N_5887);
nor U8025 (N_8025,N_7252,N_7096);
and U8026 (N_8026,N_6160,N_6880);
nand U8027 (N_8027,N_6885,N_5716);
or U8028 (N_8028,N_7299,N_6445);
or U8029 (N_8029,N_6341,N_5897);
nor U8030 (N_8030,N_6645,N_6325);
nor U8031 (N_8031,N_6700,N_6518);
or U8032 (N_8032,N_5160,N_7374);
and U8033 (N_8033,N_6827,N_7153);
and U8034 (N_8034,N_7463,N_6636);
nor U8035 (N_8035,N_5835,N_6680);
or U8036 (N_8036,N_5480,N_5015);
nor U8037 (N_8037,N_5449,N_6149);
and U8038 (N_8038,N_5490,N_7280);
nand U8039 (N_8039,N_6025,N_6672);
nand U8040 (N_8040,N_6905,N_7448);
or U8041 (N_8041,N_7175,N_5096);
xor U8042 (N_8042,N_6373,N_5156);
nand U8043 (N_8043,N_6724,N_5378);
nor U8044 (N_8044,N_5934,N_5405);
nor U8045 (N_8045,N_5608,N_7054);
xnor U8046 (N_8046,N_7457,N_6711);
nor U8047 (N_8047,N_5513,N_7251);
or U8048 (N_8048,N_6162,N_5676);
or U8049 (N_8049,N_5374,N_6065);
nand U8050 (N_8050,N_6279,N_5956);
nor U8051 (N_8051,N_6690,N_6300);
nand U8052 (N_8052,N_6158,N_6809);
nand U8053 (N_8053,N_5872,N_5312);
or U8054 (N_8054,N_5458,N_5743);
nand U8055 (N_8055,N_5913,N_6857);
nor U8056 (N_8056,N_6879,N_6930);
and U8057 (N_8057,N_6294,N_6270);
nand U8058 (N_8058,N_6753,N_7419);
or U8059 (N_8059,N_5766,N_6709);
nor U8060 (N_8060,N_7406,N_7146);
and U8061 (N_8061,N_5004,N_5137);
and U8062 (N_8062,N_6543,N_7100);
nor U8063 (N_8063,N_5284,N_5603);
nor U8064 (N_8064,N_5532,N_7447);
nand U8065 (N_8065,N_6881,N_5606);
nor U8066 (N_8066,N_5257,N_6981);
or U8067 (N_8067,N_5548,N_5358);
and U8068 (N_8068,N_5380,N_5011);
nor U8069 (N_8069,N_6834,N_5057);
nor U8070 (N_8070,N_7101,N_6686);
or U8071 (N_8071,N_5959,N_7272);
nand U8072 (N_8072,N_5801,N_5662);
nor U8073 (N_8073,N_5867,N_5211);
or U8074 (N_8074,N_7328,N_7439);
nor U8075 (N_8075,N_5749,N_6499);
or U8076 (N_8076,N_6264,N_6313);
nand U8077 (N_8077,N_6781,N_6984);
or U8078 (N_8078,N_7405,N_5013);
nor U8079 (N_8079,N_6646,N_7019);
nor U8080 (N_8080,N_5778,N_6609);
or U8081 (N_8081,N_6320,N_7246);
and U8082 (N_8082,N_7422,N_5273);
nand U8083 (N_8083,N_6192,N_5781);
and U8084 (N_8084,N_5785,N_6684);
and U8085 (N_8085,N_6604,N_7366);
xor U8086 (N_8086,N_5855,N_5291);
or U8087 (N_8087,N_6200,N_6239);
or U8088 (N_8088,N_5690,N_6455);
or U8089 (N_8089,N_7047,N_5154);
or U8090 (N_8090,N_5050,N_6970);
nand U8091 (N_8091,N_6528,N_5878);
or U8092 (N_8092,N_6161,N_6372);
nand U8093 (N_8093,N_6889,N_6467);
and U8094 (N_8094,N_5241,N_5303);
and U8095 (N_8095,N_7370,N_7279);
nor U8096 (N_8096,N_6079,N_5266);
nand U8097 (N_8097,N_5474,N_5390);
nand U8098 (N_8098,N_6140,N_5373);
nor U8099 (N_8099,N_6283,N_6910);
nand U8100 (N_8100,N_6167,N_5512);
nor U8101 (N_8101,N_5916,N_5502);
or U8102 (N_8102,N_5861,N_5275);
nand U8103 (N_8103,N_6884,N_6039);
nand U8104 (N_8104,N_6442,N_5966);
nor U8105 (N_8105,N_5078,N_6577);
nand U8106 (N_8106,N_6928,N_6549);
and U8107 (N_8107,N_5703,N_6964);
and U8108 (N_8108,N_6483,N_7000);
nand U8109 (N_8109,N_5534,N_5227);
nand U8110 (N_8110,N_6435,N_5262);
nand U8111 (N_8111,N_6965,N_5270);
and U8112 (N_8112,N_5997,N_6275);
nand U8113 (N_8113,N_5252,N_5837);
or U8114 (N_8114,N_7213,N_5991);
nand U8115 (N_8115,N_6537,N_5584);
or U8116 (N_8116,N_5758,N_6412);
nor U8117 (N_8117,N_5814,N_7454);
nand U8118 (N_8118,N_5675,N_5402);
nor U8119 (N_8119,N_6101,N_6656);
nor U8120 (N_8120,N_6311,N_5721);
or U8121 (N_8121,N_6429,N_5193);
nand U8122 (N_8122,N_6030,N_6420);
and U8123 (N_8123,N_5326,N_5973);
nand U8124 (N_8124,N_6272,N_6371);
and U8125 (N_8125,N_5591,N_6925);
nand U8126 (N_8126,N_6095,N_6482);
nor U8127 (N_8127,N_7326,N_5152);
nor U8128 (N_8128,N_5946,N_5084);
and U8129 (N_8129,N_6293,N_5598);
and U8130 (N_8130,N_5344,N_6128);
or U8131 (N_8131,N_6967,N_6717);
nor U8132 (N_8132,N_6422,N_6749);
nand U8133 (N_8133,N_7114,N_5457);
and U8134 (N_8134,N_7160,N_6779);
nand U8135 (N_8135,N_6585,N_6269);
and U8136 (N_8136,N_5466,N_6419);
and U8137 (N_8137,N_7453,N_5195);
and U8138 (N_8138,N_5805,N_5274);
nor U8139 (N_8139,N_5419,N_5051);
nand U8140 (N_8140,N_6408,N_5467);
or U8141 (N_8141,N_5862,N_6514);
nor U8142 (N_8142,N_5952,N_6440);
nand U8143 (N_8143,N_5258,N_7296);
nor U8144 (N_8144,N_5334,N_6786);
nand U8145 (N_8145,N_7210,N_5967);
and U8146 (N_8146,N_5294,N_6380);
nand U8147 (N_8147,N_6496,N_6099);
nor U8148 (N_8148,N_7124,N_6247);
nor U8149 (N_8149,N_7225,N_5325);
nor U8150 (N_8150,N_5376,N_7099);
or U8151 (N_8151,N_6054,N_6404);
and U8152 (N_8152,N_5994,N_6143);
nand U8153 (N_8153,N_7076,N_7310);
nand U8154 (N_8154,N_5908,N_5136);
or U8155 (N_8155,N_5863,N_6532);
or U8156 (N_8156,N_6078,N_6586);
and U8157 (N_8157,N_6251,N_6759);
nor U8158 (N_8158,N_7292,N_5833);
nor U8159 (N_8159,N_6542,N_7201);
nor U8160 (N_8160,N_6350,N_6395);
nor U8161 (N_8161,N_7072,N_5151);
or U8162 (N_8162,N_6515,N_7346);
nor U8163 (N_8163,N_6816,N_5535);
or U8164 (N_8164,N_5698,N_6813);
and U8165 (N_8165,N_6231,N_5705);
nor U8166 (N_8166,N_5251,N_5483);
nand U8167 (N_8167,N_6043,N_5680);
or U8168 (N_8168,N_7499,N_5234);
nor U8169 (N_8169,N_6492,N_5782);
nand U8170 (N_8170,N_6237,N_5434);
nor U8171 (N_8171,N_5717,N_6979);
nor U8172 (N_8172,N_7498,N_6612);
nand U8173 (N_8173,N_7382,N_5347);
xnor U8174 (N_8174,N_7415,N_7035);
nand U8175 (N_8175,N_6521,N_5784);
and U8176 (N_8176,N_7042,N_6335);
nor U8177 (N_8177,N_5107,N_5949);
and U8178 (N_8178,N_5707,N_6168);
or U8179 (N_8179,N_5444,N_6454);
and U8180 (N_8180,N_5930,N_5728);
or U8181 (N_8181,N_5304,N_6060);
nor U8182 (N_8182,N_5074,N_5150);
nor U8183 (N_8183,N_7115,N_5568);
and U8184 (N_8184,N_7129,N_6587);
nand U8185 (N_8185,N_6484,N_5818);
and U8186 (N_8186,N_6971,N_6308);
or U8187 (N_8187,N_5578,N_5572);
nand U8188 (N_8188,N_5848,N_6864);
nand U8189 (N_8189,N_7387,N_5346);
nor U8190 (N_8190,N_6003,N_6824);
or U8191 (N_8191,N_7137,N_5542);
or U8192 (N_8192,N_5232,N_6962);
nand U8193 (N_8193,N_7458,N_5964);
nand U8194 (N_8194,N_6755,N_7449);
or U8195 (N_8195,N_6343,N_5910);
nand U8196 (N_8196,N_5179,N_5381);
nand U8197 (N_8197,N_7452,N_5714);
nor U8198 (N_8198,N_5510,N_7333);
or U8199 (N_8199,N_6013,N_6062);
or U8200 (N_8200,N_7020,N_6122);
nor U8201 (N_8201,N_6456,N_5300);
or U8202 (N_8202,N_5579,N_5909);
and U8203 (N_8203,N_5870,N_6523);
and U8204 (N_8204,N_6860,N_6947);
nand U8205 (N_8205,N_6610,N_6148);
or U8206 (N_8206,N_5367,N_6546);
nor U8207 (N_8207,N_6908,N_6529);
nand U8208 (N_8208,N_5178,N_7212);
nor U8209 (N_8209,N_6211,N_5541);
nand U8210 (N_8210,N_7143,N_6538);
or U8211 (N_8211,N_6216,N_5960);
nor U8212 (N_8212,N_7330,N_5377);
and U8213 (N_8213,N_6359,N_5026);
nor U8214 (N_8214,N_6246,N_7024);
and U8215 (N_8215,N_7238,N_6250);
and U8216 (N_8216,N_7222,N_5106);
and U8217 (N_8217,N_6741,N_6862);
and U8218 (N_8218,N_5517,N_6116);
or U8219 (N_8219,N_7003,N_6017);
nor U8220 (N_8220,N_6083,N_7032);
and U8221 (N_8221,N_5222,N_6262);
or U8222 (N_8222,N_5630,N_6352);
nand U8223 (N_8223,N_7337,N_6500);
nand U8224 (N_8224,N_6870,N_5288);
nor U8225 (N_8225,N_7386,N_6479);
or U8226 (N_8226,N_5361,N_6907);
and U8227 (N_8227,N_6561,N_6282);
nand U8228 (N_8228,N_5065,N_5687);
and U8229 (N_8229,N_5041,N_7363);
nand U8230 (N_8230,N_7332,N_5882);
nand U8231 (N_8231,N_5615,N_5401);
or U8232 (N_8232,N_5142,N_6223);
nor U8233 (N_8233,N_6135,N_5307);
or U8234 (N_8234,N_6991,N_6147);
nor U8235 (N_8235,N_5674,N_7360);
or U8236 (N_8236,N_6058,N_5849);
or U8237 (N_8237,N_6297,N_6229);
nand U8238 (N_8238,N_7394,N_6285);
or U8239 (N_8239,N_5099,N_6789);
nand U8240 (N_8240,N_6392,N_6590);
or U8241 (N_8241,N_5221,N_5158);
or U8242 (N_8242,N_7059,N_6354);
and U8243 (N_8243,N_5478,N_7351);
and U8244 (N_8244,N_5200,N_6975);
nor U8245 (N_8245,N_6036,N_6029);
and U8246 (N_8246,N_5253,N_6077);
nand U8247 (N_8247,N_7154,N_6005);
nor U8248 (N_8248,N_6772,N_7227);
and U8249 (N_8249,N_6252,N_5464);
and U8250 (N_8250,N_6622,N_6338);
or U8251 (N_8251,N_5220,N_6055);
and U8252 (N_8252,N_6673,N_6191);
and U8253 (N_8253,N_6056,N_7465);
nand U8254 (N_8254,N_5161,N_6624);
nand U8255 (N_8255,N_6266,N_6451);
nand U8256 (N_8256,N_5364,N_6301);
and U8257 (N_8257,N_5409,N_5528);
and U8258 (N_8258,N_5636,N_5190);
nand U8259 (N_8259,N_7057,N_5083);
nand U8260 (N_8260,N_6038,N_6244);
nor U8261 (N_8261,N_6958,N_5821);
and U8262 (N_8262,N_5349,N_6364);
nand U8263 (N_8263,N_5939,N_5009);
nor U8264 (N_8264,N_5246,N_5907);
nor U8265 (N_8265,N_6205,N_5619);
and U8266 (N_8266,N_6059,N_5113);
nor U8267 (N_8267,N_7339,N_7357);
or U8268 (N_8268,N_5048,N_6090);
or U8269 (N_8269,N_6388,N_6858);
or U8270 (N_8270,N_5660,N_6207);
nor U8271 (N_8271,N_5767,N_7034);
or U8272 (N_8272,N_6276,N_5665);
nor U8273 (N_8273,N_5901,N_6954);
or U8274 (N_8274,N_5972,N_6714);
or U8275 (N_8275,N_5327,N_7157);
nor U8276 (N_8276,N_6936,N_5094);
or U8277 (N_8277,N_7450,N_5345);
or U8278 (N_8278,N_5811,N_5896);
nor U8279 (N_8279,N_6345,N_5560);
nand U8280 (N_8280,N_6399,N_5168);
and U8281 (N_8281,N_5840,N_5747);
nor U8282 (N_8282,N_6977,N_5588);
nand U8283 (N_8283,N_5927,N_6401);
nor U8284 (N_8284,N_5635,N_6799);
or U8285 (N_8285,N_7283,N_5191);
nand U8286 (N_8286,N_5806,N_5033);
nand U8287 (N_8287,N_7461,N_7088);
or U8288 (N_8288,N_7189,N_6008);
nand U8289 (N_8289,N_7340,N_5892);
nand U8290 (N_8290,N_5148,N_5663);
nor U8291 (N_8291,N_6349,N_6100);
nor U8292 (N_8292,N_5460,N_5816);
nand U8293 (N_8293,N_5121,N_5938);
or U8294 (N_8294,N_5006,N_7358);
and U8295 (N_8295,N_6581,N_5465);
nor U8296 (N_8296,N_6334,N_7148);
or U8297 (N_8297,N_6010,N_6517);
nor U8298 (N_8298,N_7442,N_6774);
nor U8299 (N_8299,N_6939,N_5445);
and U8300 (N_8300,N_5576,N_7014);
or U8301 (N_8301,N_5046,N_7486);
xor U8302 (N_8302,N_5132,N_6489);
or U8303 (N_8303,N_6243,N_7070);
nand U8304 (N_8304,N_6387,N_5832);
and U8305 (N_8305,N_6127,N_5764);
or U8306 (N_8306,N_5765,N_5443);
and U8307 (N_8307,N_6238,N_6098);
and U8308 (N_8308,N_7097,N_5003);
nor U8309 (N_8309,N_5394,N_6727);
nand U8310 (N_8310,N_6051,N_6138);
or U8311 (N_8311,N_7172,N_6915);
nor U8312 (N_8312,N_6783,N_5089);
xor U8313 (N_8313,N_5895,N_5757);
nor U8314 (N_8314,N_5315,N_5563);
nand U8315 (N_8315,N_5858,N_5889);
nor U8316 (N_8316,N_5153,N_6949);
nand U8317 (N_8317,N_5164,N_6296);
nand U8318 (N_8318,N_7315,N_7383);
nand U8319 (N_8319,N_6498,N_5421);
or U8320 (N_8320,N_5412,N_6274);
nand U8321 (N_8321,N_6378,N_5998);
or U8322 (N_8322,N_7050,N_5556);
nor U8323 (N_8323,N_6132,N_6494);
or U8324 (N_8324,N_5536,N_6342);
nor U8325 (N_8325,N_5103,N_6739);
nor U8326 (N_8326,N_6236,N_6477);
and U8327 (N_8327,N_6428,N_7392);
or U8328 (N_8328,N_7169,N_6020);
nand U8329 (N_8329,N_5726,N_5370);
nand U8330 (N_8330,N_7053,N_5559);
nor U8331 (N_8331,N_6210,N_6798);
or U8332 (N_8332,N_6808,N_5117);
nand U8333 (N_8333,N_7205,N_5614);
or U8334 (N_8334,N_7132,N_7017);
or U8335 (N_8335,N_6268,N_5482);
or U8336 (N_8336,N_7451,N_6478);
nor U8337 (N_8337,N_7180,N_5804);
and U8338 (N_8338,N_5157,N_6421);
nor U8339 (N_8339,N_5400,N_5918);
and U8340 (N_8340,N_6882,N_6658);
xnor U8341 (N_8341,N_6353,N_6374);
nor U8342 (N_8342,N_6750,N_6503);
or U8343 (N_8343,N_5963,N_6575);
or U8344 (N_8344,N_7235,N_6691);
nand U8345 (N_8345,N_5110,N_6728);
or U8346 (N_8346,N_5912,N_7380);
or U8347 (N_8347,N_6224,N_5673);
and U8348 (N_8348,N_6746,N_6932);
nor U8349 (N_8349,N_5032,N_5571);
xor U8350 (N_8350,N_7171,N_6853);
nor U8351 (N_8351,N_7151,N_5643);
nor U8352 (N_8352,N_7379,N_6547);
nor U8353 (N_8353,N_5875,N_6938);
or U8354 (N_8354,N_5922,N_5115);
and U8355 (N_8355,N_5184,N_6550);
nor U8356 (N_8356,N_5217,N_6945);
nand U8357 (N_8357,N_6016,N_6473);
and U8358 (N_8358,N_6876,N_7216);
nor U8359 (N_8359,N_5522,N_7203);
nor U8360 (N_8360,N_5034,N_5403);
nor U8361 (N_8361,N_7162,N_5173);
or U8362 (N_8362,N_7230,N_7069);
or U8363 (N_8363,N_5456,N_5622);
nor U8364 (N_8364,N_6629,N_6463);
nand U8365 (N_8365,N_6641,N_7105);
nor U8366 (N_8366,N_7078,N_6185);
or U8367 (N_8367,N_5640,N_5281);
nor U8368 (N_8368,N_5087,N_7324);
nand U8369 (N_8369,N_6920,N_6901);
and U8370 (N_8370,N_6933,N_5677);
nor U8371 (N_8371,N_5197,N_5759);
or U8372 (N_8372,N_5491,N_5010);
or U8373 (N_8373,N_5950,N_5331);
and U8374 (N_8374,N_5426,N_6137);
or U8375 (N_8375,N_5056,N_7400);
and U8376 (N_8376,N_5729,N_6924);
or U8377 (N_8377,N_5600,N_5623);
nor U8378 (N_8378,N_6890,N_7103);
or U8379 (N_8379,N_6506,N_6556);
nand U8380 (N_8380,N_6040,N_6448);
nand U8381 (N_8381,N_6261,N_5415);
nor U8382 (N_8382,N_6715,N_5302);
and U8383 (N_8383,N_5397,N_5093);
or U8384 (N_8384,N_6877,N_6133);
xnor U8385 (N_8385,N_5068,N_5612);
nor U8386 (N_8386,N_7349,N_5455);
nand U8387 (N_8387,N_7010,N_7381);
nand U8388 (N_8388,N_5567,N_6770);
nor U8389 (N_8389,N_5320,N_5285);
or U8390 (N_8390,N_6315,N_6771);
or U8391 (N_8391,N_7287,N_5475);
and U8392 (N_8392,N_7416,N_6327);
nand U8393 (N_8393,N_7045,N_5760);
nand U8394 (N_8394,N_6366,N_5686);
or U8395 (N_8395,N_6987,N_6716);
nand U8396 (N_8396,N_7278,N_5144);
or U8397 (N_8397,N_5860,N_5411);
nor U8398 (N_8398,N_5372,N_6524);
nor U8399 (N_8399,N_5228,N_6848);
or U8400 (N_8400,N_5540,N_6330);
and U8401 (N_8401,N_5350,N_6024);
or U8402 (N_8402,N_5696,N_5289);
nor U8403 (N_8403,N_6763,N_6657);
and U8404 (N_8404,N_5487,N_6234);
and U8405 (N_8405,N_7040,N_5802);
or U8406 (N_8406,N_7174,N_6544);
and U8407 (N_8407,N_5035,N_6340);
nor U8408 (N_8408,N_7338,N_5506);
nor U8409 (N_8409,N_7140,N_6403);
nand U8410 (N_8410,N_6379,N_7066);
nand U8411 (N_8411,N_5544,N_6757);
nand U8412 (N_8412,N_5735,N_7471);
nand U8413 (N_8413,N_5883,N_6108);
nand U8414 (N_8414,N_6722,N_7026);
and U8415 (N_8415,N_5180,N_6736);
and U8416 (N_8416,N_6668,N_6540);
and U8417 (N_8417,N_6918,N_6832);
nand U8418 (N_8418,N_5118,N_6034);
or U8419 (N_8419,N_5321,N_6769);
xor U8420 (N_8420,N_5263,N_5592);
and U8421 (N_8421,N_5702,N_6248);
nor U8422 (N_8422,N_5843,N_5219);
nor U8423 (N_8423,N_6513,N_6199);
nand U8424 (N_8424,N_6893,N_7288);
or U8425 (N_8425,N_6963,N_6245);
nor U8426 (N_8426,N_6826,N_5366);
and U8427 (N_8427,N_5055,N_5914);
nand U8428 (N_8428,N_6570,N_5825);
or U8429 (N_8429,N_7226,N_5667);
nor U8430 (N_8430,N_6687,N_5898);
or U8431 (N_8431,N_7029,N_5075);
and U8432 (N_8432,N_5537,N_6872);
nand U8433 (N_8433,N_6303,N_6183);
nand U8434 (N_8434,N_5448,N_6130);
or U8435 (N_8435,N_6988,N_5723);
and U8436 (N_8436,N_7044,N_5545);
and U8437 (N_8437,N_6754,N_5120);
or U8438 (N_8438,N_6747,N_7081);
or U8439 (N_8439,N_6208,N_5363);
and U8440 (N_8440,N_5986,N_5008);
nor U8441 (N_8441,N_6019,N_6878);
and U8442 (N_8442,N_5595,N_7495);
or U8443 (N_8443,N_5783,N_7134);
and U8444 (N_8444,N_6843,N_5587);
nand U8445 (N_8445,N_6002,N_6914);
nand U8446 (N_8446,N_7427,N_7270);
or U8447 (N_8447,N_6431,N_7223);
and U8448 (N_8448,N_6326,N_7083);
or U8449 (N_8449,N_5016,N_6927);
nand U8450 (N_8450,N_5509,N_6385);
and U8451 (N_8451,N_6721,N_6545);
and U8452 (N_8452,N_6304,N_6699);
nor U8453 (N_8453,N_7196,N_7168);
and U8454 (N_8454,N_7384,N_6810);
and U8455 (N_8455,N_6064,N_5247);
nor U8456 (N_8456,N_6595,N_5174);
nand U8457 (N_8457,N_6548,N_6088);
or U8458 (N_8458,N_5525,N_6968);
or U8459 (N_8459,N_6430,N_6376);
nor U8460 (N_8460,N_6683,N_7335);
and U8461 (N_8461,N_5029,N_6894);
nor U8462 (N_8462,N_6871,N_5418);
nor U8463 (N_8463,N_5752,N_7079);
and U8464 (N_8464,N_6726,N_6634);
xor U8465 (N_8465,N_6708,N_7191);
and U8466 (N_8466,N_6583,N_6873);
or U8467 (N_8467,N_5399,N_6926);
nor U8468 (N_8468,N_5942,N_6941);
and U8469 (N_8469,N_5297,N_5044);
nor U8470 (N_8470,N_5720,N_6066);
or U8471 (N_8471,N_6607,N_5516);
or U8472 (N_8472,N_5864,N_7018);
nand U8473 (N_8473,N_7104,N_6468);
and U8474 (N_8474,N_5172,N_6391);
nand U8475 (N_8475,N_5706,N_6004);
or U8476 (N_8476,N_5063,N_6616);
nand U8477 (N_8477,N_6868,N_5961);
and U8478 (N_8478,N_6046,N_5932);
or U8479 (N_8479,N_6068,N_5877);
nor U8480 (N_8480,N_6053,N_7414);
nand U8481 (N_8481,N_6493,N_5079);
and U8482 (N_8482,N_5076,N_5476);
and U8483 (N_8483,N_6314,N_5473);
and U8484 (N_8484,N_5206,N_5468);
nand U8485 (N_8485,N_6921,N_5423);
and U8486 (N_8486,N_6536,N_7149);
nor U8487 (N_8487,N_5265,N_5853);
or U8488 (N_8488,N_5886,N_7007);
or U8489 (N_8489,N_5424,N_6626);
and U8490 (N_8490,N_6197,N_7177);
nand U8491 (N_8491,N_5751,N_5577);
or U8492 (N_8492,N_6405,N_5383);
or U8493 (N_8493,N_6801,N_5441);
and U8494 (N_8494,N_6600,N_7342);
and U8495 (N_8495,N_5624,N_6913);
nand U8496 (N_8496,N_7102,N_6390);
nor U8497 (N_8497,N_7255,N_7233);
or U8498 (N_8498,N_6042,N_7407);
or U8499 (N_8499,N_5122,N_6666);
or U8500 (N_8500,N_6995,N_5030);
or U8501 (N_8501,N_5322,N_6384);
nand U8502 (N_8502,N_5407,N_7095);
nor U8503 (N_8503,N_5683,N_6181);
nand U8504 (N_8504,N_5529,N_5235);
nor U8505 (N_8505,N_6414,N_5613);
nand U8506 (N_8506,N_6087,N_6647);
nand U8507 (N_8507,N_6212,N_5171);
and U8508 (N_8508,N_5831,N_5520);
nor U8509 (N_8509,N_6823,N_6865);
nor U8510 (N_8510,N_6310,N_6295);
xor U8511 (N_8511,N_6718,N_5527);
nand U8512 (N_8512,N_6072,N_5043);
or U8513 (N_8513,N_5049,N_5131);
or U8514 (N_8514,N_5408,N_5658);
and U8515 (N_8515,N_6822,N_5809);
or U8516 (N_8516,N_5925,N_5188);
nand U8517 (N_8517,N_5176,N_7430);
nand U8518 (N_8518,N_7031,N_5355);
nand U8519 (N_8519,N_6579,N_6323);
or U8520 (N_8520,N_6015,N_7462);
nor U8521 (N_8521,N_6174,N_6999);
and U8522 (N_8522,N_5974,N_5854);
and U8523 (N_8523,N_5037,N_5980);
nor U8524 (N_8524,N_7039,N_5427);
nand U8525 (N_8525,N_6141,N_7364);
nand U8526 (N_8526,N_5097,N_5836);
or U8527 (N_8527,N_5072,N_6080);
and U8528 (N_8528,N_6785,N_6847);
or U8529 (N_8529,N_7220,N_5888);
nand U8530 (N_8530,N_6171,N_6324);
or U8531 (N_8531,N_5597,N_7206);
nor U8532 (N_8532,N_5069,N_5881);
nor U8533 (N_8533,N_5119,N_6255);
and U8534 (N_8534,N_6837,N_6075);
and U8535 (N_8535,N_7373,N_5020);
and U8536 (N_8536,N_6782,N_7187);
nand U8537 (N_8537,N_6961,N_5114);
nor U8538 (N_8538,N_6662,N_5202);
or U8539 (N_8539,N_5791,N_6642);
or U8540 (N_8540,N_5442,N_7190);
and U8541 (N_8541,N_6228,N_5734);
or U8542 (N_8542,N_6887,N_7435);
and U8543 (N_8543,N_5794,N_5216);
nor U8544 (N_8544,N_6113,N_5666);
nor U8545 (N_8545,N_5554,N_6644);
nand U8546 (N_8546,N_6094,N_6510);
nor U8547 (N_8547,N_5332,N_6706);
and U8548 (N_8548,N_6407,N_6803);
nand U8549 (N_8549,N_6555,N_6791);
nor U8550 (N_8550,N_6389,N_6050);
and U8551 (N_8551,N_7156,N_7411);
nand U8552 (N_8552,N_6396,N_5741);
nor U8553 (N_8553,N_6632,N_6427);
or U8554 (N_8554,N_7028,N_7110);
nor U8555 (N_8555,N_6398,N_6534);
nor U8556 (N_8556,N_6986,N_7098);
nor U8557 (N_8557,N_6256,N_5761);
nor U8558 (N_8558,N_6552,N_5031);
nor U8559 (N_8559,N_6047,N_6564);
nand U8560 (N_8560,N_5957,N_5001);
nor U8561 (N_8561,N_5147,N_6213);
and U8562 (N_8562,N_7359,N_5385);
nor U8563 (N_8563,N_5845,N_5983);
or U8564 (N_8564,N_7274,N_6131);
and U8565 (N_8565,N_6659,N_5492);
and U8566 (N_8566,N_7385,N_7067);
nand U8567 (N_8567,N_5066,N_7483);
nand U8568 (N_8568,N_6766,N_5224);
or U8569 (N_8569,N_6710,N_5865);
and U8570 (N_8570,N_6225,N_5091);
and U8571 (N_8571,N_7361,N_5471);
nand U8572 (N_8572,N_5793,N_5329);
nand U8573 (N_8573,N_5388,N_5452);
and U8574 (N_8574,N_6109,N_6818);
or U8575 (N_8575,N_6287,N_6674);
nor U8576 (N_8576,N_6375,N_6023);
nor U8577 (N_8577,N_6909,N_7494);
nand U8578 (N_8578,N_6091,N_6994);
or U8579 (N_8579,N_7403,N_7221);
xor U8580 (N_8580,N_7183,N_6846);
and U8581 (N_8581,N_5671,N_6501);
or U8582 (N_8582,N_5249,N_6260);
and U8583 (N_8583,N_5900,N_6220);
and U8584 (N_8584,N_5712,N_5771);
nand U8585 (N_8585,N_5256,N_5260);
nor U8586 (N_8586,N_6535,N_5095);
nand U8587 (N_8587,N_6682,N_5194);
and U8588 (N_8588,N_5277,N_7228);
nor U8589 (N_8589,N_6725,N_5847);
nand U8590 (N_8590,N_5198,N_6474);
and U8591 (N_8591,N_5130,N_6679);
or U8592 (N_8592,N_5447,N_6866);
and U8593 (N_8593,N_5846,N_5283);
nor U8594 (N_8594,N_6281,N_6415);
nor U8595 (N_8595,N_7429,N_5979);
or U8596 (N_8596,N_5187,N_6362);
nor U8597 (N_8597,N_6196,N_6980);
nand U8598 (N_8598,N_7362,N_6111);
or U8599 (N_8599,N_6631,N_5393);
nor U8600 (N_8600,N_5725,N_5678);
nor U8601 (N_8601,N_5585,N_7150);
nor U8602 (N_8602,N_5518,N_5231);
nand U8603 (N_8603,N_6063,N_6069);
or U8604 (N_8604,N_6896,N_5170);
or U8605 (N_8605,N_6118,N_5954);
or U8606 (N_8606,N_6851,N_7474);
or U8607 (N_8607,N_5634,N_6667);
nor U8608 (N_8608,N_5486,N_6365);
nand U8609 (N_8609,N_7068,N_7085);
nor U8610 (N_8610,N_6426,N_6453);
or U8611 (N_8611,N_5601,N_7302);
nor U8612 (N_8612,N_7352,N_5018);
nor U8613 (N_8613,N_7303,N_5593);
or U8614 (N_8614,N_6985,N_6944);
and U8615 (N_8615,N_6178,N_7445);
or U8616 (N_8616,N_7224,N_7065);
nand U8617 (N_8617,N_6106,N_6625);
nor U8618 (N_8618,N_6508,N_6377);
xor U8619 (N_8619,N_5338,N_7051);
xor U8620 (N_8620,N_6339,N_5086);
nor U8621 (N_8621,N_5777,N_7365);
or U8622 (N_8622,N_5796,N_5574);
nand U8623 (N_8623,N_5852,N_5028);
nor U8624 (N_8624,N_6795,N_7265);
nor U8625 (N_8625,N_7055,N_5024);
and U8626 (N_8626,N_7119,N_7398);
nand U8627 (N_8627,N_6215,N_7164);
and U8628 (N_8628,N_5842,N_5135);
or U8629 (N_8629,N_6998,N_5295);
nand U8630 (N_8630,N_6952,N_6271);
nand U8631 (N_8631,N_5159,N_7444);
nor U8632 (N_8632,N_5205,N_6911);
and U8633 (N_8633,N_6558,N_5040);
nor U8634 (N_8634,N_5857,N_6969);
nand U8635 (N_8635,N_6946,N_6014);
nor U8636 (N_8636,N_5495,N_6874);
nor U8637 (N_8637,N_7307,N_6424);
nand U8638 (N_8638,N_6021,N_7166);
and U8639 (N_8639,N_6531,N_6703);
nor U8640 (N_8640,N_6361,N_7258);
or U8641 (N_8641,N_7094,N_7327);
nor U8642 (N_8642,N_5602,N_6743);
or U8643 (N_8643,N_5225,N_5694);
nand U8644 (N_8644,N_6254,N_7012);
or U8645 (N_8645,N_6620,N_7350);
nor U8646 (N_8646,N_6990,N_7135);
nand U8647 (N_8647,N_6329,N_5659);
and U8648 (N_8648,N_5839,N_6425);
nor U8649 (N_8649,N_7412,N_7011);
nand U8650 (N_8650,N_6768,N_7421);
nand U8651 (N_8651,N_6567,N_5167);
or U8652 (N_8652,N_5787,N_7367);
nor U8653 (N_8653,N_5981,N_7023);
nand U8654 (N_8654,N_6299,N_5292);
nor U8655 (N_8655,N_6675,N_7248);
nand U8656 (N_8656,N_5196,N_7170);
and U8657 (N_8657,N_6704,N_5557);
xnor U8658 (N_8658,N_6465,N_7195);
and U8659 (N_8659,N_7390,N_5489);
nand U8660 (N_8660,N_5109,N_5149);
nor U8661 (N_8661,N_7188,N_7276);
nor U8662 (N_8662,N_6692,N_5067);
or U8663 (N_8663,N_7395,N_6611);
and U8664 (N_8664,N_7219,N_5637);
or U8665 (N_8665,N_7277,N_5203);
and U8666 (N_8666,N_6488,N_5310);
nor U8667 (N_8667,N_6993,N_7336);
or U8668 (N_8668,N_7401,N_6693);
nand U8669 (N_8669,N_6627,N_6151);
nand U8670 (N_8670,N_7490,N_6643);
nor U8671 (N_8671,N_5504,N_7165);
nand U8672 (N_8672,N_6416,N_7480);
nor U8673 (N_8673,N_5829,N_6983);
and U8674 (N_8674,N_7181,N_5740);
nand U8675 (N_8675,N_5139,N_5061);
nor U8676 (N_8676,N_6288,N_5668);
nand U8677 (N_8677,N_7048,N_5163);
and U8678 (N_8678,N_5360,N_7241);
nand U8679 (N_8679,N_7158,N_6566);
nand U8680 (N_8680,N_7344,N_5977);
nand U8681 (N_8681,N_6328,N_6793);
nor U8682 (N_8682,N_5324,N_5988);
nand U8683 (N_8683,N_6173,N_7128);
and U8684 (N_8684,N_5098,N_7231);
nand U8685 (N_8685,N_5924,N_5919);
nor U8686 (N_8686,N_7271,N_5589);
nand U8687 (N_8687,N_7396,N_7472);
nor U8688 (N_8688,N_5699,N_5639);
nand U8689 (N_8689,N_5208,N_5214);
nand U8690 (N_8690,N_5472,N_6203);
nor U8691 (N_8691,N_7476,N_7242);
and U8692 (N_8692,N_5070,N_6976);
nor U8693 (N_8693,N_5627,N_5820);
and U8694 (N_8694,N_5420,N_6972);
and U8695 (N_8695,N_5580,N_5105);
nor U8696 (N_8696,N_5817,N_5450);
nor U8697 (N_8697,N_5431,N_7341);
nor U8698 (N_8698,N_6527,N_7434);
or U8699 (N_8699,N_5023,N_6777);
nor U8700 (N_8700,N_6305,N_5021);
or U8701 (N_8701,N_6346,N_5064);
nor U8702 (N_8702,N_6480,N_7347);
nor U8703 (N_8703,N_6833,N_7125);
nand U8704 (N_8704,N_7275,N_5254);
and U8705 (N_8705,N_5569,N_5555);
or U8706 (N_8706,N_5493,N_6402);
or U8707 (N_8707,N_6796,N_6732);
or U8708 (N_8708,N_6461,N_6615);
and U8709 (N_8709,N_7460,N_6992);
nor U8710 (N_8710,N_5183,N_6114);
and U8711 (N_8711,N_6145,N_5059);
nor U8712 (N_8712,N_6578,N_7389);
nand U8713 (N_8713,N_7487,N_5422);
nand U8714 (N_8714,N_7256,N_6760);
nand U8715 (N_8715,N_7440,N_6232);
or U8716 (N_8716,N_5685,N_5937);
and U8717 (N_8717,N_5773,N_5681);
and U8718 (N_8718,N_5682,N_7420);
nor U8719 (N_8719,N_6740,N_6195);
nand U8720 (N_8720,N_5395,N_7015);
nand U8721 (N_8721,N_7147,N_6292);
and U8722 (N_8722,N_6829,N_6713);
or U8723 (N_8723,N_6509,N_6560);
and U8724 (N_8724,N_6897,N_5417);
nor U8725 (N_8725,N_6198,N_6318);
nand U8726 (N_8726,N_5669,N_6541);
or U8727 (N_8727,N_5186,N_6966);
nand U8728 (N_8728,N_5090,N_6041);
nand U8729 (N_8729,N_7459,N_6433);
or U8730 (N_8730,N_5299,N_7426);
nand U8731 (N_8731,N_7323,N_5226);
or U8732 (N_8732,N_5521,N_6411);
nor U8733 (N_8733,N_6929,N_6633);
nor U8734 (N_8734,N_7077,N_7266);
and U8735 (N_8735,N_5868,N_6032);
or U8736 (N_8736,N_5503,N_7431);
nor U8737 (N_8737,N_6125,N_5851);
nand U8738 (N_8738,N_5772,N_5413);
or U8739 (N_8739,N_6253,N_5742);
or U8740 (N_8740,N_5485,N_6802);
and U8741 (N_8741,N_5245,N_7456);
and U8742 (N_8742,N_6974,N_6383);
nor U8743 (N_8743,N_5995,N_5891);
nor U8744 (N_8744,N_5255,N_5182);
and U8745 (N_8745,N_6953,N_6000);
nor U8746 (N_8746,N_6648,N_5494);
or U8747 (N_8747,N_5129,N_5082);
nor U8748 (N_8748,N_6121,N_5353);
or U8749 (N_8749,N_6370,N_7192);
nor U8750 (N_8750,N_7170,N_5593);
nor U8751 (N_8751,N_6975,N_5950);
nand U8752 (N_8752,N_5552,N_6616);
and U8753 (N_8753,N_7190,N_6812);
nor U8754 (N_8754,N_5408,N_7153);
or U8755 (N_8755,N_5712,N_5742);
or U8756 (N_8756,N_7371,N_5688);
nand U8757 (N_8757,N_6376,N_5714);
and U8758 (N_8758,N_6998,N_5523);
nor U8759 (N_8759,N_6275,N_6066);
nor U8760 (N_8760,N_7425,N_7129);
and U8761 (N_8761,N_5456,N_6956);
nand U8762 (N_8762,N_7408,N_6936);
nand U8763 (N_8763,N_5192,N_6953);
or U8764 (N_8764,N_7349,N_6177);
or U8765 (N_8765,N_7155,N_5679);
nor U8766 (N_8766,N_5832,N_5245);
nand U8767 (N_8767,N_5667,N_5938);
and U8768 (N_8768,N_6364,N_5422);
or U8769 (N_8769,N_6088,N_7034);
or U8770 (N_8770,N_5256,N_6149);
nand U8771 (N_8771,N_7118,N_5979);
and U8772 (N_8772,N_6851,N_5345);
or U8773 (N_8773,N_7036,N_6148);
and U8774 (N_8774,N_7085,N_6883);
nor U8775 (N_8775,N_6070,N_5172);
nor U8776 (N_8776,N_6716,N_6037);
nand U8777 (N_8777,N_6714,N_5024);
and U8778 (N_8778,N_5394,N_6890);
and U8779 (N_8779,N_7134,N_6635);
nor U8780 (N_8780,N_5671,N_5836);
and U8781 (N_8781,N_6661,N_7490);
nand U8782 (N_8782,N_7297,N_6860);
nor U8783 (N_8783,N_5864,N_6312);
or U8784 (N_8784,N_5548,N_5345);
and U8785 (N_8785,N_6974,N_6737);
nand U8786 (N_8786,N_6395,N_7084);
nand U8787 (N_8787,N_5695,N_5747);
nor U8788 (N_8788,N_5457,N_5084);
nand U8789 (N_8789,N_6223,N_7348);
nand U8790 (N_8790,N_5477,N_7319);
and U8791 (N_8791,N_6440,N_6124);
nand U8792 (N_8792,N_7254,N_6573);
nor U8793 (N_8793,N_6428,N_7086);
or U8794 (N_8794,N_7358,N_5503);
nor U8795 (N_8795,N_6693,N_6520);
nand U8796 (N_8796,N_6836,N_6113);
nand U8797 (N_8797,N_5355,N_5581);
and U8798 (N_8798,N_5470,N_7069);
nor U8799 (N_8799,N_6194,N_7227);
and U8800 (N_8800,N_6812,N_6230);
and U8801 (N_8801,N_7466,N_5522);
nor U8802 (N_8802,N_6764,N_5075);
nor U8803 (N_8803,N_5769,N_5744);
or U8804 (N_8804,N_7451,N_5643);
and U8805 (N_8805,N_5637,N_6503);
nor U8806 (N_8806,N_6274,N_5970);
and U8807 (N_8807,N_7082,N_6778);
nor U8808 (N_8808,N_5318,N_6801);
nand U8809 (N_8809,N_5340,N_5452);
nor U8810 (N_8810,N_5727,N_5852);
and U8811 (N_8811,N_6580,N_7270);
nand U8812 (N_8812,N_6499,N_5447);
nand U8813 (N_8813,N_6182,N_6197);
nor U8814 (N_8814,N_6115,N_6483);
or U8815 (N_8815,N_5696,N_6764);
xor U8816 (N_8816,N_6080,N_6062);
nor U8817 (N_8817,N_6412,N_7083);
nor U8818 (N_8818,N_5603,N_6353);
nor U8819 (N_8819,N_6262,N_5152);
or U8820 (N_8820,N_6316,N_5188);
nand U8821 (N_8821,N_5135,N_5136);
xnor U8822 (N_8822,N_7308,N_7083);
nor U8823 (N_8823,N_6414,N_5099);
or U8824 (N_8824,N_7390,N_7320);
nand U8825 (N_8825,N_6630,N_7138);
or U8826 (N_8826,N_6983,N_5302);
or U8827 (N_8827,N_5496,N_6084);
or U8828 (N_8828,N_6601,N_6184);
xnor U8829 (N_8829,N_6110,N_6921);
and U8830 (N_8830,N_6350,N_5226);
nor U8831 (N_8831,N_5906,N_6742);
and U8832 (N_8832,N_6836,N_5110);
or U8833 (N_8833,N_5845,N_6805);
nor U8834 (N_8834,N_5180,N_6894);
nor U8835 (N_8835,N_5009,N_7163);
nor U8836 (N_8836,N_7434,N_6095);
nand U8837 (N_8837,N_7418,N_5360);
nor U8838 (N_8838,N_7078,N_5801);
or U8839 (N_8839,N_5364,N_6085);
and U8840 (N_8840,N_7303,N_6598);
nand U8841 (N_8841,N_6785,N_6103);
nor U8842 (N_8842,N_5392,N_5527);
nor U8843 (N_8843,N_6716,N_7120);
or U8844 (N_8844,N_5313,N_6278);
nand U8845 (N_8845,N_7095,N_7251);
and U8846 (N_8846,N_5581,N_6529);
nand U8847 (N_8847,N_6669,N_6920);
nor U8848 (N_8848,N_6460,N_5210);
nand U8849 (N_8849,N_6710,N_5679);
or U8850 (N_8850,N_7447,N_5889);
or U8851 (N_8851,N_7149,N_7285);
nor U8852 (N_8852,N_7084,N_5586);
nand U8853 (N_8853,N_6144,N_6507);
nor U8854 (N_8854,N_5972,N_5849);
or U8855 (N_8855,N_5568,N_6224);
or U8856 (N_8856,N_5150,N_6723);
nor U8857 (N_8857,N_7184,N_6925);
nor U8858 (N_8858,N_7178,N_5153);
nor U8859 (N_8859,N_7355,N_7279);
nor U8860 (N_8860,N_7205,N_6347);
and U8861 (N_8861,N_5700,N_6619);
and U8862 (N_8862,N_5431,N_7120);
nand U8863 (N_8863,N_6776,N_7132);
or U8864 (N_8864,N_7475,N_6568);
nand U8865 (N_8865,N_6624,N_5597);
nand U8866 (N_8866,N_5366,N_6495);
or U8867 (N_8867,N_6590,N_5156);
and U8868 (N_8868,N_6250,N_6792);
or U8869 (N_8869,N_6038,N_6907);
and U8870 (N_8870,N_6100,N_5446);
and U8871 (N_8871,N_7418,N_5159);
and U8872 (N_8872,N_5727,N_6322);
nand U8873 (N_8873,N_5066,N_6778);
or U8874 (N_8874,N_5472,N_6903);
nor U8875 (N_8875,N_5431,N_6967);
or U8876 (N_8876,N_5152,N_6301);
nand U8877 (N_8877,N_7255,N_6799);
or U8878 (N_8878,N_6773,N_7099);
nand U8879 (N_8879,N_6869,N_7414);
nand U8880 (N_8880,N_6300,N_6040);
nor U8881 (N_8881,N_6911,N_5375);
nand U8882 (N_8882,N_5686,N_5468);
nor U8883 (N_8883,N_6529,N_6703);
or U8884 (N_8884,N_5354,N_5565);
nor U8885 (N_8885,N_6247,N_7087);
and U8886 (N_8886,N_6319,N_7082);
or U8887 (N_8887,N_5638,N_6740);
nor U8888 (N_8888,N_7497,N_6690);
and U8889 (N_8889,N_5388,N_6242);
and U8890 (N_8890,N_7430,N_5736);
or U8891 (N_8891,N_7492,N_5316);
and U8892 (N_8892,N_6173,N_5646);
and U8893 (N_8893,N_6518,N_6252);
or U8894 (N_8894,N_7293,N_7228);
nor U8895 (N_8895,N_7416,N_6194);
and U8896 (N_8896,N_7129,N_7011);
or U8897 (N_8897,N_6311,N_5197);
and U8898 (N_8898,N_6032,N_7447);
nand U8899 (N_8899,N_5623,N_5188);
and U8900 (N_8900,N_7303,N_5398);
nand U8901 (N_8901,N_7367,N_6928);
nor U8902 (N_8902,N_5937,N_5664);
nand U8903 (N_8903,N_7025,N_6695);
and U8904 (N_8904,N_6564,N_6844);
and U8905 (N_8905,N_5627,N_5440);
and U8906 (N_8906,N_6765,N_6421);
nand U8907 (N_8907,N_5040,N_7147);
and U8908 (N_8908,N_5360,N_7393);
nand U8909 (N_8909,N_5866,N_5359);
and U8910 (N_8910,N_7004,N_5975);
or U8911 (N_8911,N_7142,N_6347);
nand U8912 (N_8912,N_6444,N_6443);
nand U8913 (N_8913,N_6757,N_5390);
nor U8914 (N_8914,N_5478,N_5229);
nor U8915 (N_8915,N_6029,N_6021);
nand U8916 (N_8916,N_7268,N_7200);
and U8917 (N_8917,N_6942,N_5684);
nor U8918 (N_8918,N_6215,N_5130);
or U8919 (N_8919,N_7379,N_5237);
and U8920 (N_8920,N_6170,N_5706);
nor U8921 (N_8921,N_7067,N_7237);
or U8922 (N_8922,N_7155,N_7125);
or U8923 (N_8923,N_6969,N_6622);
nand U8924 (N_8924,N_5244,N_6564);
xor U8925 (N_8925,N_6001,N_6094);
nor U8926 (N_8926,N_5426,N_6755);
xor U8927 (N_8927,N_7143,N_6033);
and U8928 (N_8928,N_5149,N_6152);
or U8929 (N_8929,N_6431,N_5362);
nand U8930 (N_8930,N_5942,N_5358);
and U8931 (N_8931,N_5111,N_6635);
and U8932 (N_8932,N_5720,N_6961);
or U8933 (N_8933,N_5234,N_7253);
or U8934 (N_8934,N_6076,N_6860);
nand U8935 (N_8935,N_7428,N_5529);
nand U8936 (N_8936,N_7248,N_5719);
and U8937 (N_8937,N_5272,N_6341);
nor U8938 (N_8938,N_7116,N_6366);
nand U8939 (N_8939,N_7155,N_5222);
nand U8940 (N_8940,N_6813,N_6777);
nand U8941 (N_8941,N_5724,N_6952);
nand U8942 (N_8942,N_6882,N_7226);
nor U8943 (N_8943,N_6682,N_5226);
nor U8944 (N_8944,N_5093,N_5047);
or U8945 (N_8945,N_6438,N_5649);
nand U8946 (N_8946,N_5292,N_6072);
and U8947 (N_8947,N_5725,N_5360);
nor U8948 (N_8948,N_6103,N_6375);
or U8949 (N_8949,N_7248,N_5524);
or U8950 (N_8950,N_6269,N_6147);
nand U8951 (N_8951,N_6353,N_5802);
nand U8952 (N_8952,N_7439,N_6225);
and U8953 (N_8953,N_7388,N_5622);
nand U8954 (N_8954,N_7037,N_5806);
nand U8955 (N_8955,N_6296,N_7459);
nor U8956 (N_8956,N_5289,N_7218);
nand U8957 (N_8957,N_5056,N_6832);
nor U8958 (N_8958,N_5047,N_6715);
and U8959 (N_8959,N_6274,N_6824);
nand U8960 (N_8960,N_5220,N_6426);
or U8961 (N_8961,N_5909,N_5308);
and U8962 (N_8962,N_5786,N_5428);
or U8963 (N_8963,N_5547,N_6012);
and U8964 (N_8964,N_7007,N_5173);
and U8965 (N_8965,N_5171,N_7171);
nor U8966 (N_8966,N_6992,N_5461);
nor U8967 (N_8967,N_5516,N_7162);
and U8968 (N_8968,N_5062,N_5829);
nor U8969 (N_8969,N_7003,N_6862);
and U8970 (N_8970,N_6783,N_6997);
or U8971 (N_8971,N_5323,N_6222);
nor U8972 (N_8972,N_5035,N_5762);
nor U8973 (N_8973,N_7466,N_6200);
nand U8974 (N_8974,N_5337,N_6586);
or U8975 (N_8975,N_6029,N_5782);
or U8976 (N_8976,N_6281,N_5741);
and U8977 (N_8977,N_5725,N_5445);
or U8978 (N_8978,N_7450,N_5829);
or U8979 (N_8979,N_5829,N_6686);
or U8980 (N_8980,N_6577,N_7026);
nor U8981 (N_8981,N_7061,N_6434);
xor U8982 (N_8982,N_5087,N_5110);
nand U8983 (N_8983,N_5841,N_5430);
or U8984 (N_8984,N_6517,N_7432);
nand U8985 (N_8985,N_6134,N_6432);
nor U8986 (N_8986,N_6715,N_5598);
nand U8987 (N_8987,N_5219,N_6507);
nand U8988 (N_8988,N_5577,N_6413);
and U8989 (N_8989,N_7458,N_6228);
nand U8990 (N_8990,N_6701,N_7385);
and U8991 (N_8991,N_7382,N_6856);
nand U8992 (N_8992,N_6126,N_5157);
and U8993 (N_8993,N_5944,N_5892);
or U8994 (N_8994,N_5605,N_6214);
nor U8995 (N_8995,N_5960,N_7146);
nor U8996 (N_8996,N_5723,N_6794);
nand U8997 (N_8997,N_6303,N_6832);
or U8998 (N_8998,N_7436,N_6093);
or U8999 (N_8999,N_5559,N_6333);
nand U9000 (N_9000,N_6311,N_5810);
and U9001 (N_9001,N_5630,N_5792);
nand U9002 (N_9002,N_5468,N_5376);
nor U9003 (N_9003,N_6464,N_7163);
nor U9004 (N_9004,N_5638,N_7446);
and U9005 (N_9005,N_6281,N_6060);
nor U9006 (N_9006,N_7485,N_6136);
and U9007 (N_9007,N_7319,N_5019);
nand U9008 (N_9008,N_5338,N_5398);
and U9009 (N_9009,N_6811,N_6083);
nor U9010 (N_9010,N_6511,N_5199);
or U9011 (N_9011,N_6924,N_6944);
or U9012 (N_9012,N_7169,N_5648);
nand U9013 (N_9013,N_7246,N_5288);
nand U9014 (N_9014,N_6634,N_6395);
nand U9015 (N_9015,N_5427,N_7272);
or U9016 (N_9016,N_6109,N_6984);
nand U9017 (N_9017,N_5782,N_5023);
nor U9018 (N_9018,N_6144,N_6973);
or U9019 (N_9019,N_5424,N_7018);
and U9020 (N_9020,N_6410,N_7184);
nor U9021 (N_9021,N_7201,N_5549);
and U9022 (N_9022,N_6356,N_5316);
nand U9023 (N_9023,N_6896,N_7014);
and U9024 (N_9024,N_5256,N_7424);
and U9025 (N_9025,N_5533,N_6612);
nand U9026 (N_9026,N_5919,N_5279);
or U9027 (N_9027,N_6717,N_7097);
nor U9028 (N_9028,N_5525,N_5381);
and U9029 (N_9029,N_6597,N_5644);
nor U9030 (N_9030,N_6390,N_6471);
and U9031 (N_9031,N_7472,N_6865);
and U9032 (N_9032,N_5790,N_5183);
and U9033 (N_9033,N_5876,N_7246);
and U9034 (N_9034,N_7135,N_6568);
nand U9035 (N_9035,N_6915,N_6734);
and U9036 (N_9036,N_5796,N_7493);
nand U9037 (N_9037,N_5564,N_6189);
and U9038 (N_9038,N_5403,N_7197);
or U9039 (N_9039,N_6736,N_6953);
or U9040 (N_9040,N_5003,N_5772);
nor U9041 (N_9041,N_6033,N_5397);
nand U9042 (N_9042,N_5228,N_6720);
nand U9043 (N_9043,N_7066,N_5818);
nor U9044 (N_9044,N_6440,N_5453);
and U9045 (N_9045,N_5313,N_5924);
and U9046 (N_9046,N_5732,N_5323);
nand U9047 (N_9047,N_6862,N_6677);
and U9048 (N_9048,N_7438,N_5835);
nand U9049 (N_9049,N_5623,N_6385);
nand U9050 (N_9050,N_5549,N_5600);
nand U9051 (N_9051,N_5193,N_7114);
or U9052 (N_9052,N_6348,N_7256);
nand U9053 (N_9053,N_7445,N_6236);
nand U9054 (N_9054,N_6864,N_6901);
and U9055 (N_9055,N_6316,N_7373);
or U9056 (N_9056,N_6627,N_7291);
or U9057 (N_9057,N_5209,N_5606);
and U9058 (N_9058,N_6208,N_5186);
and U9059 (N_9059,N_5740,N_6680);
and U9060 (N_9060,N_5166,N_6429);
or U9061 (N_9061,N_6269,N_5576);
nor U9062 (N_9062,N_7450,N_6695);
and U9063 (N_9063,N_7286,N_6985);
nor U9064 (N_9064,N_5064,N_6082);
or U9065 (N_9065,N_6501,N_7067);
nand U9066 (N_9066,N_6955,N_6974);
and U9067 (N_9067,N_6020,N_6550);
and U9068 (N_9068,N_5377,N_6741);
and U9069 (N_9069,N_5984,N_5114);
and U9070 (N_9070,N_6115,N_5305);
nor U9071 (N_9071,N_5066,N_7312);
nand U9072 (N_9072,N_6058,N_7003);
and U9073 (N_9073,N_5144,N_7198);
nand U9074 (N_9074,N_6441,N_6388);
nor U9075 (N_9075,N_5231,N_5164);
nor U9076 (N_9076,N_6989,N_5649);
nor U9077 (N_9077,N_7394,N_5187);
or U9078 (N_9078,N_6331,N_7194);
or U9079 (N_9079,N_6416,N_7226);
nand U9080 (N_9080,N_5231,N_6068);
nor U9081 (N_9081,N_6751,N_5943);
nand U9082 (N_9082,N_6368,N_5703);
nor U9083 (N_9083,N_6185,N_6347);
and U9084 (N_9084,N_5820,N_6795);
nand U9085 (N_9085,N_5439,N_6341);
and U9086 (N_9086,N_7231,N_6272);
nand U9087 (N_9087,N_7440,N_5572);
nand U9088 (N_9088,N_6128,N_7011);
or U9089 (N_9089,N_7461,N_6123);
nand U9090 (N_9090,N_7246,N_7482);
or U9091 (N_9091,N_5042,N_6386);
and U9092 (N_9092,N_6381,N_5112);
or U9093 (N_9093,N_5611,N_6324);
nand U9094 (N_9094,N_5656,N_5085);
or U9095 (N_9095,N_6796,N_5535);
and U9096 (N_9096,N_5996,N_7222);
or U9097 (N_9097,N_6360,N_6943);
and U9098 (N_9098,N_6612,N_6686);
or U9099 (N_9099,N_6894,N_5879);
nand U9100 (N_9100,N_7456,N_7084);
and U9101 (N_9101,N_6718,N_6012);
nand U9102 (N_9102,N_5802,N_6893);
or U9103 (N_9103,N_6297,N_5116);
nand U9104 (N_9104,N_6892,N_7048);
nand U9105 (N_9105,N_6940,N_7009);
and U9106 (N_9106,N_5195,N_5470);
nor U9107 (N_9107,N_7499,N_5217);
nand U9108 (N_9108,N_6398,N_7342);
nand U9109 (N_9109,N_5718,N_7009);
or U9110 (N_9110,N_7071,N_5244);
or U9111 (N_9111,N_7418,N_6268);
xnor U9112 (N_9112,N_5957,N_5051);
and U9113 (N_9113,N_5437,N_5415);
nand U9114 (N_9114,N_5652,N_5567);
nor U9115 (N_9115,N_6455,N_7375);
nor U9116 (N_9116,N_6187,N_5150);
nand U9117 (N_9117,N_6891,N_6295);
or U9118 (N_9118,N_6177,N_6496);
nor U9119 (N_9119,N_5305,N_7376);
and U9120 (N_9120,N_5123,N_7100);
or U9121 (N_9121,N_5463,N_6558);
nor U9122 (N_9122,N_7059,N_6784);
or U9123 (N_9123,N_7085,N_5773);
and U9124 (N_9124,N_5574,N_6424);
nand U9125 (N_9125,N_7059,N_6590);
nand U9126 (N_9126,N_5386,N_5755);
nor U9127 (N_9127,N_6699,N_5005);
nor U9128 (N_9128,N_7151,N_5499);
and U9129 (N_9129,N_5997,N_5000);
nor U9130 (N_9130,N_7024,N_5766);
and U9131 (N_9131,N_6537,N_6429);
and U9132 (N_9132,N_6473,N_5770);
nand U9133 (N_9133,N_5434,N_5573);
nor U9134 (N_9134,N_5976,N_6084);
and U9135 (N_9135,N_6572,N_6635);
or U9136 (N_9136,N_5097,N_6393);
nand U9137 (N_9137,N_6423,N_7302);
or U9138 (N_9138,N_6541,N_5623);
nand U9139 (N_9139,N_7232,N_5122);
nor U9140 (N_9140,N_5983,N_6418);
nor U9141 (N_9141,N_7380,N_5900);
nor U9142 (N_9142,N_7197,N_6988);
nor U9143 (N_9143,N_5222,N_7496);
and U9144 (N_9144,N_6079,N_5885);
nor U9145 (N_9145,N_5349,N_6400);
and U9146 (N_9146,N_5144,N_5491);
and U9147 (N_9147,N_6243,N_7409);
or U9148 (N_9148,N_5102,N_5150);
or U9149 (N_9149,N_5834,N_5055);
nand U9150 (N_9150,N_5562,N_6998);
nand U9151 (N_9151,N_7488,N_6516);
or U9152 (N_9152,N_6405,N_7269);
and U9153 (N_9153,N_5964,N_7359);
nor U9154 (N_9154,N_5601,N_5015);
or U9155 (N_9155,N_7306,N_7352);
or U9156 (N_9156,N_6965,N_6659);
and U9157 (N_9157,N_5408,N_6287);
or U9158 (N_9158,N_6777,N_5039);
and U9159 (N_9159,N_6085,N_6327);
and U9160 (N_9160,N_7251,N_7394);
or U9161 (N_9161,N_6482,N_7342);
or U9162 (N_9162,N_6189,N_6144);
and U9163 (N_9163,N_5409,N_5238);
nor U9164 (N_9164,N_5612,N_5744);
nand U9165 (N_9165,N_6489,N_5608);
or U9166 (N_9166,N_6441,N_6307);
or U9167 (N_9167,N_5992,N_6224);
and U9168 (N_9168,N_6354,N_6637);
and U9169 (N_9169,N_5200,N_5448);
nor U9170 (N_9170,N_5705,N_5842);
nand U9171 (N_9171,N_5335,N_6434);
or U9172 (N_9172,N_6078,N_5065);
nor U9173 (N_9173,N_6295,N_7287);
nand U9174 (N_9174,N_6128,N_6051);
nand U9175 (N_9175,N_5248,N_7115);
nand U9176 (N_9176,N_6938,N_5926);
or U9177 (N_9177,N_5174,N_6219);
nand U9178 (N_9178,N_6298,N_7300);
and U9179 (N_9179,N_6095,N_5549);
or U9180 (N_9180,N_7133,N_7397);
nor U9181 (N_9181,N_5957,N_7186);
and U9182 (N_9182,N_6682,N_6745);
or U9183 (N_9183,N_6521,N_5569);
and U9184 (N_9184,N_5108,N_5408);
and U9185 (N_9185,N_6823,N_5014);
nand U9186 (N_9186,N_5539,N_7165);
and U9187 (N_9187,N_6813,N_5390);
or U9188 (N_9188,N_7362,N_6013);
nand U9189 (N_9189,N_6185,N_6188);
nand U9190 (N_9190,N_5109,N_6267);
nor U9191 (N_9191,N_5322,N_6947);
or U9192 (N_9192,N_6765,N_6574);
xnor U9193 (N_9193,N_7065,N_7103);
nand U9194 (N_9194,N_5526,N_5542);
and U9195 (N_9195,N_7178,N_5568);
and U9196 (N_9196,N_5546,N_5297);
nor U9197 (N_9197,N_6200,N_6927);
nor U9198 (N_9198,N_6812,N_6657);
nand U9199 (N_9199,N_7136,N_7057);
or U9200 (N_9200,N_7123,N_6155);
and U9201 (N_9201,N_6373,N_7352);
or U9202 (N_9202,N_5396,N_5135);
and U9203 (N_9203,N_6409,N_6223);
and U9204 (N_9204,N_5616,N_6387);
or U9205 (N_9205,N_7463,N_5483);
or U9206 (N_9206,N_5243,N_5263);
nand U9207 (N_9207,N_6617,N_5184);
and U9208 (N_9208,N_5044,N_7040);
or U9209 (N_9209,N_6756,N_6102);
nor U9210 (N_9210,N_6328,N_6029);
and U9211 (N_9211,N_6126,N_5894);
nand U9212 (N_9212,N_6247,N_5867);
nand U9213 (N_9213,N_6868,N_5975);
nor U9214 (N_9214,N_5931,N_5462);
and U9215 (N_9215,N_7036,N_7173);
or U9216 (N_9216,N_7481,N_7342);
nor U9217 (N_9217,N_7172,N_6272);
nand U9218 (N_9218,N_7418,N_6353);
nand U9219 (N_9219,N_6622,N_6082);
nor U9220 (N_9220,N_5749,N_6818);
xnor U9221 (N_9221,N_6753,N_5601);
and U9222 (N_9222,N_5482,N_5213);
nor U9223 (N_9223,N_7488,N_6882);
or U9224 (N_9224,N_5683,N_6723);
or U9225 (N_9225,N_5131,N_5595);
or U9226 (N_9226,N_5572,N_5996);
and U9227 (N_9227,N_7162,N_7235);
nand U9228 (N_9228,N_5008,N_6110);
nor U9229 (N_9229,N_5116,N_5217);
nand U9230 (N_9230,N_5289,N_6697);
xor U9231 (N_9231,N_6019,N_7099);
xor U9232 (N_9232,N_5875,N_7060);
or U9233 (N_9233,N_5059,N_5916);
nand U9234 (N_9234,N_5501,N_6678);
and U9235 (N_9235,N_5935,N_7240);
or U9236 (N_9236,N_6952,N_6653);
or U9237 (N_9237,N_5143,N_6146);
or U9238 (N_9238,N_7290,N_7247);
nand U9239 (N_9239,N_6716,N_6940);
or U9240 (N_9240,N_6030,N_6952);
nor U9241 (N_9241,N_6511,N_7058);
nor U9242 (N_9242,N_6346,N_5251);
nand U9243 (N_9243,N_5328,N_6549);
nand U9244 (N_9244,N_6083,N_6577);
or U9245 (N_9245,N_5128,N_6493);
nor U9246 (N_9246,N_5675,N_7039);
or U9247 (N_9247,N_5410,N_6301);
nand U9248 (N_9248,N_6911,N_5086);
and U9249 (N_9249,N_7216,N_6405);
or U9250 (N_9250,N_5092,N_5664);
and U9251 (N_9251,N_5868,N_5703);
and U9252 (N_9252,N_6390,N_6005);
and U9253 (N_9253,N_7366,N_6954);
nor U9254 (N_9254,N_5125,N_6589);
and U9255 (N_9255,N_6500,N_5375);
and U9256 (N_9256,N_7492,N_6496);
or U9257 (N_9257,N_6527,N_6184);
nand U9258 (N_9258,N_5150,N_7110);
nor U9259 (N_9259,N_5506,N_5817);
and U9260 (N_9260,N_6533,N_5044);
nor U9261 (N_9261,N_5257,N_5915);
or U9262 (N_9262,N_7274,N_5821);
nand U9263 (N_9263,N_7052,N_5179);
nand U9264 (N_9264,N_6477,N_7000);
nand U9265 (N_9265,N_6069,N_5106);
nor U9266 (N_9266,N_6480,N_5852);
and U9267 (N_9267,N_5286,N_5685);
xnor U9268 (N_9268,N_7173,N_5176);
and U9269 (N_9269,N_6655,N_5350);
nor U9270 (N_9270,N_5786,N_6217);
or U9271 (N_9271,N_5210,N_6811);
nor U9272 (N_9272,N_5606,N_6516);
and U9273 (N_9273,N_5466,N_5393);
nor U9274 (N_9274,N_5155,N_6741);
nand U9275 (N_9275,N_6234,N_5217);
nor U9276 (N_9276,N_7233,N_7006);
or U9277 (N_9277,N_5687,N_7435);
and U9278 (N_9278,N_5720,N_7409);
and U9279 (N_9279,N_6805,N_6142);
nand U9280 (N_9280,N_6259,N_7084);
and U9281 (N_9281,N_7160,N_7145);
or U9282 (N_9282,N_7091,N_5868);
and U9283 (N_9283,N_6000,N_6343);
and U9284 (N_9284,N_6890,N_7165);
or U9285 (N_9285,N_6044,N_6698);
nand U9286 (N_9286,N_7227,N_6115);
or U9287 (N_9287,N_5644,N_5537);
and U9288 (N_9288,N_6398,N_5139);
and U9289 (N_9289,N_7033,N_5044);
or U9290 (N_9290,N_5916,N_6585);
nor U9291 (N_9291,N_5218,N_6388);
and U9292 (N_9292,N_6033,N_5883);
nor U9293 (N_9293,N_6217,N_7355);
nand U9294 (N_9294,N_5062,N_7298);
or U9295 (N_9295,N_6810,N_5273);
and U9296 (N_9296,N_7117,N_5138);
and U9297 (N_9297,N_6633,N_7224);
or U9298 (N_9298,N_5711,N_6580);
or U9299 (N_9299,N_6264,N_7244);
and U9300 (N_9300,N_7259,N_5991);
nor U9301 (N_9301,N_5938,N_6345);
nor U9302 (N_9302,N_7345,N_6218);
nor U9303 (N_9303,N_5334,N_6750);
or U9304 (N_9304,N_5502,N_5115);
and U9305 (N_9305,N_6377,N_7420);
or U9306 (N_9306,N_7186,N_6065);
and U9307 (N_9307,N_5889,N_5433);
and U9308 (N_9308,N_5403,N_5816);
nand U9309 (N_9309,N_7159,N_6874);
or U9310 (N_9310,N_6194,N_5418);
and U9311 (N_9311,N_5097,N_5816);
and U9312 (N_9312,N_5871,N_6025);
and U9313 (N_9313,N_5094,N_5832);
and U9314 (N_9314,N_7418,N_6903);
and U9315 (N_9315,N_6097,N_7058);
xnor U9316 (N_9316,N_7104,N_5186);
and U9317 (N_9317,N_5184,N_6306);
nor U9318 (N_9318,N_6983,N_6540);
and U9319 (N_9319,N_5474,N_6079);
nor U9320 (N_9320,N_5254,N_6291);
or U9321 (N_9321,N_6775,N_6511);
or U9322 (N_9322,N_6454,N_6083);
nand U9323 (N_9323,N_6047,N_7460);
and U9324 (N_9324,N_6364,N_5362);
and U9325 (N_9325,N_6449,N_7248);
or U9326 (N_9326,N_7123,N_6688);
nor U9327 (N_9327,N_6591,N_6753);
nor U9328 (N_9328,N_5884,N_5770);
or U9329 (N_9329,N_5821,N_6575);
and U9330 (N_9330,N_5663,N_7147);
and U9331 (N_9331,N_6368,N_6737);
nor U9332 (N_9332,N_5832,N_5866);
nand U9333 (N_9333,N_6694,N_6871);
nand U9334 (N_9334,N_5060,N_5482);
or U9335 (N_9335,N_7056,N_5557);
or U9336 (N_9336,N_5170,N_7428);
nor U9337 (N_9337,N_7446,N_6760);
and U9338 (N_9338,N_7489,N_5725);
nand U9339 (N_9339,N_6548,N_6522);
and U9340 (N_9340,N_6765,N_6227);
nand U9341 (N_9341,N_5696,N_5522);
and U9342 (N_9342,N_5919,N_5477);
nor U9343 (N_9343,N_5518,N_6366);
and U9344 (N_9344,N_6319,N_5155);
or U9345 (N_9345,N_5835,N_5187);
nand U9346 (N_9346,N_6529,N_7096);
nor U9347 (N_9347,N_5660,N_7495);
and U9348 (N_9348,N_5744,N_6556);
or U9349 (N_9349,N_7026,N_6082);
nand U9350 (N_9350,N_5937,N_6031);
or U9351 (N_9351,N_7148,N_6033);
nand U9352 (N_9352,N_5832,N_6572);
and U9353 (N_9353,N_7037,N_7234);
nor U9354 (N_9354,N_5470,N_5078);
and U9355 (N_9355,N_5248,N_5869);
nor U9356 (N_9356,N_6093,N_6213);
and U9357 (N_9357,N_6198,N_5386);
or U9358 (N_9358,N_5384,N_6373);
and U9359 (N_9359,N_7094,N_7443);
nand U9360 (N_9360,N_5125,N_6286);
and U9361 (N_9361,N_7039,N_5007);
nand U9362 (N_9362,N_7182,N_6482);
xor U9363 (N_9363,N_5493,N_6451);
nand U9364 (N_9364,N_6265,N_5555);
or U9365 (N_9365,N_6491,N_5418);
nor U9366 (N_9366,N_7459,N_6757);
and U9367 (N_9367,N_6583,N_6571);
or U9368 (N_9368,N_5617,N_7386);
nor U9369 (N_9369,N_5309,N_5951);
nand U9370 (N_9370,N_5652,N_7007);
and U9371 (N_9371,N_7004,N_6404);
and U9372 (N_9372,N_5698,N_5170);
and U9373 (N_9373,N_7188,N_7404);
nor U9374 (N_9374,N_6390,N_7428);
or U9375 (N_9375,N_5165,N_7353);
and U9376 (N_9376,N_7201,N_6609);
nor U9377 (N_9377,N_6118,N_5370);
nand U9378 (N_9378,N_5935,N_6387);
nand U9379 (N_9379,N_6742,N_7151);
nand U9380 (N_9380,N_5438,N_7242);
nor U9381 (N_9381,N_5883,N_5958);
nand U9382 (N_9382,N_7154,N_6389);
or U9383 (N_9383,N_6554,N_6365);
nor U9384 (N_9384,N_5638,N_7007);
nand U9385 (N_9385,N_5460,N_5646);
or U9386 (N_9386,N_5812,N_5350);
nand U9387 (N_9387,N_6744,N_6863);
nand U9388 (N_9388,N_5285,N_5572);
nor U9389 (N_9389,N_6105,N_5507);
and U9390 (N_9390,N_7132,N_5766);
nand U9391 (N_9391,N_6270,N_5600);
and U9392 (N_9392,N_5112,N_7039);
nor U9393 (N_9393,N_5487,N_7279);
and U9394 (N_9394,N_5946,N_7383);
nor U9395 (N_9395,N_6173,N_6201);
nor U9396 (N_9396,N_7233,N_5262);
nand U9397 (N_9397,N_6688,N_7348);
nor U9398 (N_9398,N_7266,N_6977);
xor U9399 (N_9399,N_7335,N_6053);
nand U9400 (N_9400,N_5755,N_7003);
or U9401 (N_9401,N_6809,N_6440);
or U9402 (N_9402,N_6771,N_7186);
or U9403 (N_9403,N_6197,N_5462);
or U9404 (N_9404,N_5939,N_7032);
nand U9405 (N_9405,N_5098,N_7022);
nor U9406 (N_9406,N_7292,N_5189);
nor U9407 (N_9407,N_6509,N_7171);
or U9408 (N_9408,N_7491,N_5570);
nor U9409 (N_9409,N_7195,N_6424);
nand U9410 (N_9410,N_5355,N_6324);
or U9411 (N_9411,N_5000,N_6121);
nor U9412 (N_9412,N_6196,N_6695);
and U9413 (N_9413,N_6891,N_7428);
nor U9414 (N_9414,N_7364,N_6444);
nor U9415 (N_9415,N_5943,N_6620);
nand U9416 (N_9416,N_5895,N_7405);
nand U9417 (N_9417,N_5423,N_5920);
or U9418 (N_9418,N_6166,N_5937);
nand U9419 (N_9419,N_6761,N_5963);
nor U9420 (N_9420,N_5778,N_6875);
and U9421 (N_9421,N_6087,N_7020);
or U9422 (N_9422,N_6908,N_5926);
or U9423 (N_9423,N_5857,N_6824);
nor U9424 (N_9424,N_6976,N_6188);
and U9425 (N_9425,N_6410,N_6128);
nand U9426 (N_9426,N_6026,N_6886);
nor U9427 (N_9427,N_5397,N_7205);
and U9428 (N_9428,N_6237,N_6373);
nor U9429 (N_9429,N_7330,N_7488);
nand U9430 (N_9430,N_6879,N_7064);
nor U9431 (N_9431,N_6390,N_5246);
or U9432 (N_9432,N_6338,N_6545);
and U9433 (N_9433,N_5467,N_6743);
nand U9434 (N_9434,N_7040,N_7068);
and U9435 (N_9435,N_5324,N_6658);
or U9436 (N_9436,N_7025,N_6197);
or U9437 (N_9437,N_7359,N_7323);
and U9438 (N_9438,N_6254,N_5836);
or U9439 (N_9439,N_6516,N_6048);
or U9440 (N_9440,N_7313,N_7030);
nand U9441 (N_9441,N_7423,N_6493);
nor U9442 (N_9442,N_5739,N_6507);
and U9443 (N_9443,N_6610,N_6765);
nand U9444 (N_9444,N_6458,N_6592);
nand U9445 (N_9445,N_6634,N_6665);
or U9446 (N_9446,N_5458,N_5980);
or U9447 (N_9447,N_7011,N_6025);
nor U9448 (N_9448,N_5738,N_6745);
or U9449 (N_9449,N_6479,N_5038);
nor U9450 (N_9450,N_5317,N_7256);
nor U9451 (N_9451,N_7007,N_5781);
or U9452 (N_9452,N_5166,N_5324);
or U9453 (N_9453,N_5692,N_5219);
and U9454 (N_9454,N_7081,N_7209);
or U9455 (N_9455,N_7102,N_5205);
or U9456 (N_9456,N_6330,N_7384);
and U9457 (N_9457,N_5778,N_6305);
nand U9458 (N_9458,N_6323,N_5486);
nand U9459 (N_9459,N_7031,N_6348);
nand U9460 (N_9460,N_6746,N_5317);
and U9461 (N_9461,N_6169,N_6166);
or U9462 (N_9462,N_6344,N_7271);
and U9463 (N_9463,N_6341,N_7329);
or U9464 (N_9464,N_5317,N_5226);
nand U9465 (N_9465,N_5883,N_6560);
and U9466 (N_9466,N_6853,N_7214);
nand U9467 (N_9467,N_5642,N_5794);
and U9468 (N_9468,N_6034,N_5070);
and U9469 (N_9469,N_6158,N_5392);
or U9470 (N_9470,N_7158,N_7223);
nor U9471 (N_9471,N_6708,N_6901);
nand U9472 (N_9472,N_6296,N_6991);
or U9473 (N_9473,N_5889,N_7370);
nor U9474 (N_9474,N_6174,N_7206);
and U9475 (N_9475,N_5647,N_5770);
nand U9476 (N_9476,N_5779,N_7411);
and U9477 (N_9477,N_6220,N_6413);
or U9478 (N_9478,N_5305,N_7378);
or U9479 (N_9479,N_6271,N_6291);
or U9480 (N_9480,N_7368,N_7281);
and U9481 (N_9481,N_6346,N_5539);
or U9482 (N_9482,N_5779,N_5881);
nand U9483 (N_9483,N_7428,N_6807);
nor U9484 (N_9484,N_6461,N_6355);
and U9485 (N_9485,N_7150,N_7371);
or U9486 (N_9486,N_6836,N_7416);
xor U9487 (N_9487,N_5528,N_5275);
nand U9488 (N_9488,N_5766,N_6965);
nor U9489 (N_9489,N_7412,N_5073);
nor U9490 (N_9490,N_6997,N_5808);
or U9491 (N_9491,N_6456,N_5046);
and U9492 (N_9492,N_5449,N_6614);
nand U9493 (N_9493,N_6818,N_7144);
nand U9494 (N_9494,N_5389,N_5321);
nor U9495 (N_9495,N_6380,N_7499);
or U9496 (N_9496,N_6845,N_5273);
nand U9497 (N_9497,N_5743,N_6199);
xnor U9498 (N_9498,N_5985,N_6598);
or U9499 (N_9499,N_7166,N_5869);
and U9500 (N_9500,N_6257,N_5310);
and U9501 (N_9501,N_6016,N_6314);
nor U9502 (N_9502,N_5962,N_5580);
nand U9503 (N_9503,N_6296,N_6385);
nor U9504 (N_9504,N_6134,N_7117);
xor U9505 (N_9505,N_5368,N_7222);
nand U9506 (N_9506,N_6481,N_5912);
nor U9507 (N_9507,N_7434,N_6538);
nand U9508 (N_9508,N_5996,N_5603);
nor U9509 (N_9509,N_5777,N_6237);
and U9510 (N_9510,N_6965,N_5752);
and U9511 (N_9511,N_5988,N_5358);
and U9512 (N_9512,N_6516,N_6450);
and U9513 (N_9513,N_7072,N_6709);
nor U9514 (N_9514,N_6673,N_6541);
or U9515 (N_9515,N_5158,N_5164);
or U9516 (N_9516,N_6837,N_6673);
nand U9517 (N_9517,N_6315,N_6017);
nand U9518 (N_9518,N_7010,N_5780);
nor U9519 (N_9519,N_6857,N_5346);
nor U9520 (N_9520,N_6859,N_5414);
nor U9521 (N_9521,N_5120,N_6070);
and U9522 (N_9522,N_6386,N_7228);
nor U9523 (N_9523,N_7229,N_5627);
or U9524 (N_9524,N_6359,N_5611);
nand U9525 (N_9525,N_6368,N_5286);
or U9526 (N_9526,N_5198,N_5905);
or U9527 (N_9527,N_6455,N_7095);
and U9528 (N_9528,N_7286,N_6158);
nor U9529 (N_9529,N_6168,N_5636);
and U9530 (N_9530,N_6196,N_7377);
and U9531 (N_9531,N_7233,N_7045);
or U9532 (N_9532,N_5618,N_6549);
nor U9533 (N_9533,N_5051,N_5669);
nand U9534 (N_9534,N_6469,N_6804);
nor U9535 (N_9535,N_5474,N_6703);
nor U9536 (N_9536,N_6331,N_5145);
nor U9537 (N_9537,N_5990,N_5468);
and U9538 (N_9538,N_5994,N_7458);
or U9539 (N_9539,N_6080,N_5221);
and U9540 (N_9540,N_5776,N_7263);
nor U9541 (N_9541,N_7032,N_7349);
nand U9542 (N_9542,N_6855,N_6380);
or U9543 (N_9543,N_6485,N_5688);
nand U9544 (N_9544,N_7438,N_7228);
nand U9545 (N_9545,N_6321,N_7185);
or U9546 (N_9546,N_6362,N_7473);
nor U9547 (N_9547,N_5351,N_6265);
and U9548 (N_9548,N_7257,N_6885);
and U9549 (N_9549,N_6319,N_6927);
and U9550 (N_9550,N_6688,N_7147);
or U9551 (N_9551,N_7196,N_5328);
nor U9552 (N_9552,N_6687,N_6091);
nand U9553 (N_9553,N_5045,N_7120);
nand U9554 (N_9554,N_7367,N_5212);
nand U9555 (N_9555,N_7402,N_6768);
nand U9556 (N_9556,N_5861,N_5990);
or U9557 (N_9557,N_7195,N_6672);
nor U9558 (N_9558,N_6542,N_6813);
nor U9559 (N_9559,N_6996,N_5769);
and U9560 (N_9560,N_7293,N_5610);
and U9561 (N_9561,N_7291,N_6922);
nor U9562 (N_9562,N_6573,N_7079);
or U9563 (N_9563,N_5594,N_5792);
nor U9564 (N_9564,N_7208,N_7211);
nand U9565 (N_9565,N_6222,N_6513);
nand U9566 (N_9566,N_6690,N_5001);
nand U9567 (N_9567,N_5821,N_5615);
xor U9568 (N_9568,N_6468,N_6399);
and U9569 (N_9569,N_6407,N_5592);
or U9570 (N_9570,N_5871,N_5468);
or U9571 (N_9571,N_5588,N_7342);
nand U9572 (N_9572,N_6568,N_7163);
nor U9573 (N_9573,N_5664,N_6290);
or U9574 (N_9574,N_6519,N_5880);
nor U9575 (N_9575,N_7294,N_7183);
nand U9576 (N_9576,N_5318,N_7253);
nor U9577 (N_9577,N_6834,N_6507);
nor U9578 (N_9578,N_5794,N_5104);
nor U9579 (N_9579,N_6158,N_6744);
nor U9580 (N_9580,N_7374,N_7146);
nand U9581 (N_9581,N_5351,N_5075);
or U9582 (N_9582,N_5935,N_5657);
nor U9583 (N_9583,N_6546,N_6252);
and U9584 (N_9584,N_7477,N_6522);
and U9585 (N_9585,N_7054,N_7169);
and U9586 (N_9586,N_6331,N_7436);
and U9587 (N_9587,N_6611,N_5799);
nor U9588 (N_9588,N_6981,N_7155);
nor U9589 (N_9589,N_5633,N_5592);
nor U9590 (N_9590,N_7190,N_6278);
nand U9591 (N_9591,N_6199,N_6294);
nor U9592 (N_9592,N_6552,N_6481);
nand U9593 (N_9593,N_5855,N_7010);
nand U9594 (N_9594,N_5711,N_6108);
nand U9595 (N_9595,N_5262,N_6974);
nor U9596 (N_9596,N_6768,N_5951);
nor U9597 (N_9597,N_5082,N_5209);
and U9598 (N_9598,N_6204,N_6200);
or U9599 (N_9599,N_6860,N_5465);
nand U9600 (N_9600,N_5099,N_6052);
or U9601 (N_9601,N_6663,N_5093);
or U9602 (N_9602,N_6778,N_6877);
nor U9603 (N_9603,N_6480,N_6149);
or U9604 (N_9604,N_6918,N_5025);
or U9605 (N_9605,N_5202,N_5818);
nor U9606 (N_9606,N_5741,N_6180);
and U9607 (N_9607,N_5243,N_6452);
and U9608 (N_9608,N_6461,N_6645);
nor U9609 (N_9609,N_7398,N_6003);
nor U9610 (N_9610,N_5062,N_5853);
or U9611 (N_9611,N_5949,N_6373);
nor U9612 (N_9612,N_6701,N_6192);
nor U9613 (N_9613,N_6207,N_5360);
nand U9614 (N_9614,N_5875,N_6666);
nand U9615 (N_9615,N_6503,N_5850);
nand U9616 (N_9616,N_5366,N_5512);
and U9617 (N_9617,N_5899,N_5863);
nand U9618 (N_9618,N_7254,N_6322);
and U9619 (N_9619,N_5197,N_5003);
nand U9620 (N_9620,N_5341,N_6322);
and U9621 (N_9621,N_5702,N_7343);
nand U9622 (N_9622,N_5101,N_6558);
nand U9623 (N_9623,N_6904,N_7155);
nand U9624 (N_9624,N_6276,N_6173);
nand U9625 (N_9625,N_7475,N_5378);
nor U9626 (N_9626,N_6121,N_5682);
xor U9627 (N_9627,N_5132,N_6624);
nor U9628 (N_9628,N_7178,N_6974);
nand U9629 (N_9629,N_5552,N_6477);
nor U9630 (N_9630,N_6125,N_5800);
nand U9631 (N_9631,N_5737,N_7090);
nor U9632 (N_9632,N_5917,N_6934);
nand U9633 (N_9633,N_6200,N_5447);
or U9634 (N_9634,N_5582,N_5267);
and U9635 (N_9635,N_5911,N_5497);
and U9636 (N_9636,N_6448,N_5665);
nor U9637 (N_9637,N_6161,N_5558);
nand U9638 (N_9638,N_7349,N_5097);
nor U9639 (N_9639,N_5786,N_6390);
nor U9640 (N_9640,N_6571,N_6560);
or U9641 (N_9641,N_5766,N_7225);
and U9642 (N_9642,N_7366,N_6345);
or U9643 (N_9643,N_7456,N_6787);
nor U9644 (N_9644,N_6389,N_7067);
and U9645 (N_9645,N_7341,N_7446);
or U9646 (N_9646,N_6578,N_6646);
nor U9647 (N_9647,N_7390,N_6767);
nor U9648 (N_9648,N_7406,N_7069);
or U9649 (N_9649,N_6011,N_6392);
and U9650 (N_9650,N_5342,N_6544);
or U9651 (N_9651,N_7428,N_6433);
nand U9652 (N_9652,N_5396,N_5872);
nor U9653 (N_9653,N_5728,N_5085);
or U9654 (N_9654,N_6577,N_6036);
and U9655 (N_9655,N_5220,N_5295);
or U9656 (N_9656,N_7489,N_5217);
nand U9657 (N_9657,N_6437,N_6309);
nor U9658 (N_9658,N_6500,N_7449);
nand U9659 (N_9659,N_7404,N_5795);
or U9660 (N_9660,N_5514,N_5355);
xnor U9661 (N_9661,N_7157,N_5952);
or U9662 (N_9662,N_7159,N_7151);
nor U9663 (N_9663,N_6602,N_5511);
and U9664 (N_9664,N_5423,N_5791);
nand U9665 (N_9665,N_7347,N_5120);
nor U9666 (N_9666,N_6437,N_7376);
nor U9667 (N_9667,N_7463,N_5280);
nor U9668 (N_9668,N_5463,N_5803);
or U9669 (N_9669,N_6012,N_6657);
nand U9670 (N_9670,N_5997,N_5604);
nand U9671 (N_9671,N_5785,N_5535);
nand U9672 (N_9672,N_7370,N_7001);
and U9673 (N_9673,N_6817,N_6472);
nor U9674 (N_9674,N_7482,N_7258);
nor U9675 (N_9675,N_6218,N_6238);
nor U9676 (N_9676,N_7467,N_5167);
nor U9677 (N_9677,N_6804,N_7073);
nor U9678 (N_9678,N_7402,N_5038);
or U9679 (N_9679,N_6745,N_6994);
and U9680 (N_9680,N_6229,N_5029);
nor U9681 (N_9681,N_5531,N_6726);
nor U9682 (N_9682,N_6877,N_6714);
nor U9683 (N_9683,N_6040,N_7198);
or U9684 (N_9684,N_6917,N_5498);
and U9685 (N_9685,N_5555,N_6377);
and U9686 (N_9686,N_6706,N_5861);
nor U9687 (N_9687,N_7126,N_7187);
nand U9688 (N_9688,N_5776,N_5882);
nor U9689 (N_9689,N_5412,N_5336);
and U9690 (N_9690,N_5526,N_6012);
nor U9691 (N_9691,N_6046,N_5514);
or U9692 (N_9692,N_5666,N_6379);
and U9693 (N_9693,N_6658,N_6225);
nand U9694 (N_9694,N_6693,N_6716);
and U9695 (N_9695,N_5515,N_7158);
and U9696 (N_9696,N_6628,N_5190);
nor U9697 (N_9697,N_7052,N_6258);
nor U9698 (N_9698,N_6540,N_7074);
nand U9699 (N_9699,N_6810,N_6981);
xor U9700 (N_9700,N_5878,N_5932);
nor U9701 (N_9701,N_6086,N_5415);
and U9702 (N_9702,N_5840,N_5181);
nor U9703 (N_9703,N_6575,N_6260);
xor U9704 (N_9704,N_6000,N_6681);
and U9705 (N_9705,N_6964,N_7354);
or U9706 (N_9706,N_7418,N_6073);
nand U9707 (N_9707,N_5668,N_6486);
nand U9708 (N_9708,N_5469,N_5733);
nor U9709 (N_9709,N_5543,N_6809);
nor U9710 (N_9710,N_5549,N_6741);
nand U9711 (N_9711,N_6750,N_5284);
xnor U9712 (N_9712,N_6825,N_5769);
or U9713 (N_9713,N_6150,N_6867);
nor U9714 (N_9714,N_5770,N_5399);
and U9715 (N_9715,N_5846,N_7280);
and U9716 (N_9716,N_7489,N_5264);
and U9717 (N_9717,N_6010,N_5399);
nor U9718 (N_9718,N_5989,N_5043);
and U9719 (N_9719,N_7136,N_5788);
or U9720 (N_9720,N_6252,N_6584);
nor U9721 (N_9721,N_5978,N_5787);
or U9722 (N_9722,N_6838,N_7206);
nand U9723 (N_9723,N_6174,N_6056);
nor U9724 (N_9724,N_5200,N_5429);
nor U9725 (N_9725,N_7147,N_6439);
and U9726 (N_9726,N_6725,N_6825);
nand U9727 (N_9727,N_7432,N_7457);
and U9728 (N_9728,N_6058,N_5087);
nor U9729 (N_9729,N_6084,N_5665);
and U9730 (N_9730,N_5401,N_6475);
nor U9731 (N_9731,N_6766,N_5155);
and U9732 (N_9732,N_6064,N_5966);
or U9733 (N_9733,N_5560,N_7193);
nor U9734 (N_9734,N_6692,N_6259);
nor U9735 (N_9735,N_7215,N_7029);
or U9736 (N_9736,N_7107,N_7363);
or U9737 (N_9737,N_6383,N_6652);
or U9738 (N_9738,N_6422,N_5279);
and U9739 (N_9739,N_5681,N_6151);
nand U9740 (N_9740,N_5394,N_5997);
nand U9741 (N_9741,N_5540,N_5560);
or U9742 (N_9742,N_7079,N_5054);
nand U9743 (N_9743,N_6865,N_5231);
nand U9744 (N_9744,N_7214,N_5526);
nor U9745 (N_9745,N_5285,N_5972);
and U9746 (N_9746,N_5540,N_5763);
or U9747 (N_9747,N_5340,N_5779);
or U9748 (N_9748,N_6075,N_5813);
and U9749 (N_9749,N_7045,N_6331);
and U9750 (N_9750,N_6330,N_5434);
and U9751 (N_9751,N_6681,N_6383);
or U9752 (N_9752,N_7235,N_6697);
nand U9753 (N_9753,N_5186,N_6613);
nand U9754 (N_9754,N_6293,N_5893);
nand U9755 (N_9755,N_5076,N_6863);
or U9756 (N_9756,N_7232,N_5549);
or U9757 (N_9757,N_7009,N_5532);
nor U9758 (N_9758,N_7142,N_5465);
nand U9759 (N_9759,N_7368,N_6111);
nand U9760 (N_9760,N_5215,N_6270);
and U9761 (N_9761,N_5697,N_5705);
or U9762 (N_9762,N_5601,N_7131);
and U9763 (N_9763,N_6921,N_7012);
or U9764 (N_9764,N_6592,N_5285);
or U9765 (N_9765,N_7194,N_6764);
xor U9766 (N_9766,N_5801,N_6580);
nand U9767 (N_9767,N_5860,N_6237);
nor U9768 (N_9768,N_6194,N_7170);
nor U9769 (N_9769,N_5382,N_6983);
or U9770 (N_9770,N_6817,N_5673);
or U9771 (N_9771,N_6931,N_6985);
or U9772 (N_9772,N_5510,N_5043);
or U9773 (N_9773,N_6798,N_5702);
or U9774 (N_9774,N_6984,N_6731);
and U9775 (N_9775,N_6307,N_5093);
nand U9776 (N_9776,N_6016,N_5252);
nor U9777 (N_9777,N_6050,N_6763);
nand U9778 (N_9778,N_5943,N_6185);
or U9779 (N_9779,N_5313,N_7009);
nor U9780 (N_9780,N_5879,N_5476);
nand U9781 (N_9781,N_5588,N_7167);
and U9782 (N_9782,N_5621,N_6001);
nand U9783 (N_9783,N_6717,N_5744);
nand U9784 (N_9784,N_6055,N_6233);
nor U9785 (N_9785,N_5854,N_6665);
and U9786 (N_9786,N_7354,N_6984);
nand U9787 (N_9787,N_5810,N_6253);
nand U9788 (N_9788,N_5587,N_6033);
nand U9789 (N_9789,N_5880,N_6986);
or U9790 (N_9790,N_5239,N_5472);
or U9791 (N_9791,N_6351,N_6949);
nand U9792 (N_9792,N_6476,N_6743);
or U9793 (N_9793,N_5522,N_6702);
and U9794 (N_9794,N_6616,N_5716);
nor U9795 (N_9795,N_6323,N_6673);
or U9796 (N_9796,N_5962,N_6528);
nor U9797 (N_9797,N_7403,N_7133);
nor U9798 (N_9798,N_6642,N_6341);
and U9799 (N_9799,N_6131,N_6518);
and U9800 (N_9800,N_6400,N_6235);
or U9801 (N_9801,N_7004,N_5110);
and U9802 (N_9802,N_7326,N_5903);
nor U9803 (N_9803,N_5980,N_6096);
nand U9804 (N_9804,N_6248,N_5202);
nor U9805 (N_9805,N_6246,N_5942);
nor U9806 (N_9806,N_6647,N_6196);
and U9807 (N_9807,N_7190,N_6942);
and U9808 (N_9808,N_7369,N_7177);
or U9809 (N_9809,N_6348,N_5357);
and U9810 (N_9810,N_7317,N_7364);
nand U9811 (N_9811,N_7490,N_6198);
nor U9812 (N_9812,N_6202,N_7286);
nor U9813 (N_9813,N_5034,N_6216);
or U9814 (N_9814,N_5711,N_7232);
and U9815 (N_9815,N_6298,N_7381);
or U9816 (N_9816,N_7449,N_6345);
or U9817 (N_9817,N_6818,N_6445);
nor U9818 (N_9818,N_6548,N_6529);
and U9819 (N_9819,N_6293,N_5943);
nand U9820 (N_9820,N_6480,N_6470);
nor U9821 (N_9821,N_6209,N_7053);
nand U9822 (N_9822,N_6954,N_6914);
or U9823 (N_9823,N_7304,N_7341);
nor U9824 (N_9824,N_5037,N_7414);
nand U9825 (N_9825,N_7194,N_5532);
nor U9826 (N_9826,N_5126,N_5425);
and U9827 (N_9827,N_5119,N_5230);
or U9828 (N_9828,N_6819,N_6813);
nand U9829 (N_9829,N_6316,N_5876);
and U9830 (N_9830,N_5923,N_5850);
and U9831 (N_9831,N_6352,N_6591);
nor U9832 (N_9832,N_5124,N_5626);
nand U9833 (N_9833,N_7021,N_6856);
or U9834 (N_9834,N_6260,N_6741);
nor U9835 (N_9835,N_5584,N_6891);
nand U9836 (N_9836,N_5316,N_5954);
nand U9837 (N_9837,N_6367,N_6355);
or U9838 (N_9838,N_6273,N_7244);
and U9839 (N_9839,N_5164,N_6306);
or U9840 (N_9840,N_6232,N_6196);
nor U9841 (N_9841,N_6491,N_7172);
and U9842 (N_9842,N_7232,N_6281);
nand U9843 (N_9843,N_5381,N_6420);
and U9844 (N_9844,N_5713,N_7209);
nor U9845 (N_9845,N_5946,N_6288);
and U9846 (N_9846,N_6267,N_5721);
and U9847 (N_9847,N_6629,N_5556);
nor U9848 (N_9848,N_6539,N_5186);
nor U9849 (N_9849,N_6376,N_5295);
and U9850 (N_9850,N_5724,N_6421);
or U9851 (N_9851,N_5349,N_5275);
and U9852 (N_9852,N_5992,N_6718);
nor U9853 (N_9853,N_7265,N_6722);
or U9854 (N_9854,N_6850,N_5990);
nand U9855 (N_9855,N_6592,N_5640);
nand U9856 (N_9856,N_6931,N_5116);
nand U9857 (N_9857,N_5299,N_5937);
nand U9858 (N_9858,N_5455,N_6957);
and U9859 (N_9859,N_7121,N_5110);
nor U9860 (N_9860,N_5388,N_6828);
and U9861 (N_9861,N_5183,N_6614);
and U9862 (N_9862,N_6446,N_7187);
nor U9863 (N_9863,N_7190,N_6820);
and U9864 (N_9864,N_5545,N_5630);
and U9865 (N_9865,N_6533,N_5357);
nor U9866 (N_9866,N_6209,N_5986);
nor U9867 (N_9867,N_7205,N_6108);
and U9868 (N_9868,N_7036,N_6772);
and U9869 (N_9869,N_5797,N_5003);
or U9870 (N_9870,N_6935,N_6607);
xnor U9871 (N_9871,N_6595,N_5587);
nand U9872 (N_9872,N_6059,N_5163);
and U9873 (N_9873,N_5903,N_5394);
nor U9874 (N_9874,N_5939,N_6168);
nand U9875 (N_9875,N_7033,N_6036);
nor U9876 (N_9876,N_6996,N_6596);
nand U9877 (N_9877,N_5938,N_5669);
nor U9878 (N_9878,N_7462,N_6515);
and U9879 (N_9879,N_6756,N_5163);
nand U9880 (N_9880,N_7095,N_7176);
and U9881 (N_9881,N_6056,N_6177);
or U9882 (N_9882,N_5326,N_5224);
nor U9883 (N_9883,N_7169,N_5047);
and U9884 (N_9884,N_5436,N_5836);
or U9885 (N_9885,N_6216,N_7177);
or U9886 (N_9886,N_6790,N_6189);
nor U9887 (N_9887,N_6140,N_7269);
nand U9888 (N_9888,N_7307,N_5258);
nand U9889 (N_9889,N_6903,N_5543);
nor U9890 (N_9890,N_6199,N_7458);
nand U9891 (N_9891,N_6672,N_6334);
and U9892 (N_9892,N_6866,N_7267);
and U9893 (N_9893,N_5051,N_5039);
and U9894 (N_9894,N_6806,N_5000);
nand U9895 (N_9895,N_6416,N_5205);
or U9896 (N_9896,N_6513,N_6635);
nor U9897 (N_9897,N_6845,N_6571);
nand U9898 (N_9898,N_6352,N_5234);
and U9899 (N_9899,N_6092,N_5127);
and U9900 (N_9900,N_6159,N_5755);
nor U9901 (N_9901,N_7100,N_7208);
and U9902 (N_9902,N_7001,N_7480);
nor U9903 (N_9903,N_6550,N_6506);
nor U9904 (N_9904,N_5773,N_6912);
nand U9905 (N_9905,N_5293,N_5094);
or U9906 (N_9906,N_6193,N_5956);
and U9907 (N_9907,N_6355,N_5237);
nor U9908 (N_9908,N_6635,N_5650);
nor U9909 (N_9909,N_6106,N_7495);
and U9910 (N_9910,N_6508,N_5395);
nor U9911 (N_9911,N_5110,N_5835);
and U9912 (N_9912,N_6713,N_5369);
or U9913 (N_9913,N_7348,N_5924);
nand U9914 (N_9914,N_5852,N_7033);
xor U9915 (N_9915,N_6703,N_6663);
nand U9916 (N_9916,N_5926,N_7029);
nor U9917 (N_9917,N_6435,N_6680);
and U9918 (N_9918,N_5891,N_5332);
nand U9919 (N_9919,N_6344,N_6471);
and U9920 (N_9920,N_5808,N_5518);
or U9921 (N_9921,N_6093,N_5961);
or U9922 (N_9922,N_6039,N_6530);
nand U9923 (N_9923,N_6488,N_5957);
nor U9924 (N_9924,N_6414,N_6711);
nor U9925 (N_9925,N_6430,N_5493);
and U9926 (N_9926,N_6508,N_6178);
nor U9927 (N_9927,N_5504,N_6762);
nand U9928 (N_9928,N_6443,N_5494);
nand U9929 (N_9929,N_5975,N_7110);
nor U9930 (N_9930,N_5589,N_7290);
nor U9931 (N_9931,N_6319,N_5154);
and U9932 (N_9932,N_6463,N_6692);
and U9933 (N_9933,N_5931,N_5424);
and U9934 (N_9934,N_6341,N_5924);
and U9935 (N_9935,N_6634,N_6900);
nand U9936 (N_9936,N_7008,N_5547);
nor U9937 (N_9937,N_6656,N_7442);
nor U9938 (N_9938,N_5644,N_6615);
nor U9939 (N_9939,N_5320,N_5225);
nor U9940 (N_9940,N_5653,N_6207);
nand U9941 (N_9941,N_6797,N_5634);
nor U9942 (N_9942,N_5954,N_6379);
and U9943 (N_9943,N_5614,N_6143);
or U9944 (N_9944,N_5579,N_6700);
nand U9945 (N_9945,N_6548,N_5696);
nand U9946 (N_9946,N_5008,N_6899);
or U9947 (N_9947,N_6687,N_6217);
nand U9948 (N_9948,N_5488,N_6272);
nand U9949 (N_9949,N_5895,N_6417);
nor U9950 (N_9950,N_7206,N_7057);
nor U9951 (N_9951,N_5660,N_5709);
nor U9952 (N_9952,N_6819,N_5214);
or U9953 (N_9953,N_6052,N_5497);
and U9954 (N_9954,N_6953,N_7421);
or U9955 (N_9955,N_6627,N_5636);
or U9956 (N_9956,N_6670,N_5806);
or U9957 (N_9957,N_6898,N_5240);
nor U9958 (N_9958,N_6310,N_6355);
and U9959 (N_9959,N_6927,N_6031);
or U9960 (N_9960,N_5324,N_7008);
or U9961 (N_9961,N_7463,N_6663);
nor U9962 (N_9962,N_6235,N_5272);
or U9963 (N_9963,N_5051,N_6104);
nand U9964 (N_9964,N_5687,N_5551);
nor U9965 (N_9965,N_7151,N_6946);
or U9966 (N_9966,N_5534,N_5891);
and U9967 (N_9967,N_7325,N_7131);
or U9968 (N_9968,N_5070,N_5546);
and U9969 (N_9969,N_5362,N_6580);
nor U9970 (N_9970,N_6616,N_5868);
and U9971 (N_9971,N_5240,N_6333);
and U9972 (N_9972,N_6405,N_5192);
and U9973 (N_9973,N_7470,N_6455);
and U9974 (N_9974,N_6024,N_6842);
or U9975 (N_9975,N_6137,N_6860);
nand U9976 (N_9976,N_6573,N_6398);
nor U9977 (N_9977,N_5302,N_6934);
nor U9978 (N_9978,N_5407,N_6605);
and U9979 (N_9979,N_7376,N_5818);
or U9980 (N_9980,N_6585,N_6450);
nor U9981 (N_9981,N_6843,N_6823);
and U9982 (N_9982,N_5013,N_7238);
or U9983 (N_9983,N_6339,N_7099);
xor U9984 (N_9984,N_6407,N_6399);
nand U9985 (N_9985,N_6781,N_6149);
nand U9986 (N_9986,N_5986,N_7260);
or U9987 (N_9987,N_6193,N_6800);
nor U9988 (N_9988,N_7070,N_7406);
xor U9989 (N_9989,N_7421,N_5398);
or U9990 (N_9990,N_5150,N_6622);
and U9991 (N_9991,N_5456,N_7126);
nand U9992 (N_9992,N_5295,N_5678);
and U9993 (N_9993,N_7437,N_7074);
nor U9994 (N_9994,N_6588,N_5996);
xor U9995 (N_9995,N_5587,N_5246);
or U9996 (N_9996,N_5755,N_7214);
or U9997 (N_9997,N_6513,N_6702);
and U9998 (N_9998,N_6290,N_6805);
nand U9999 (N_9999,N_6749,N_7297);
or UO_0 (O_0,N_9591,N_9510);
nand UO_1 (O_1,N_8886,N_7981);
and UO_2 (O_2,N_9756,N_9008);
xnor UO_3 (O_3,N_8577,N_7849);
nor UO_4 (O_4,N_9328,N_9945);
and UO_5 (O_5,N_8617,N_8788);
or UO_6 (O_6,N_7684,N_8058);
and UO_7 (O_7,N_8094,N_9679);
or UO_8 (O_8,N_8305,N_7677);
or UO_9 (O_9,N_7843,N_8954);
nand UO_10 (O_10,N_9446,N_8380);
or UO_11 (O_11,N_9280,N_7708);
xor UO_12 (O_12,N_9727,N_9150);
nand UO_13 (O_13,N_8935,N_8665);
or UO_14 (O_14,N_8826,N_9893);
and UO_15 (O_15,N_9074,N_9031);
xor UO_16 (O_16,N_8450,N_8295);
xnor UO_17 (O_17,N_7940,N_9861);
and UO_18 (O_18,N_9780,N_8566);
nor UO_19 (O_19,N_8394,N_8492);
or UO_20 (O_20,N_9848,N_8174);
nor UO_21 (O_21,N_9115,N_8542);
nand UO_22 (O_22,N_8490,N_9991);
nand UO_23 (O_23,N_7837,N_9981);
nand UO_24 (O_24,N_8230,N_8589);
nand UO_25 (O_25,N_8554,N_9425);
and UO_26 (O_26,N_7530,N_8282);
nor UO_27 (O_27,N_8792,N_7746);
and UO_28 (O_28,N_9421,N_8606);
or UO_29 (O_29,N_9009,N_9605);
or UO_30 (O_30,N_8369,N_8103);
xnor UO_31 (O_31,N_8872,N_7789);
nor UO_32 (O_32,N_9768,N_9081);
nand UO_33 (O_33,N_8302,N_9118);
nand UO_34 (O_34,N_8914,N_7859);
or UO_35 (O_35,N_9391,N_8337);
nand UO_36 (O_36,N_8880,N_9284);
and UO_37 (O_37,N_8347,N_8791);
nor UO_38 (O_38,N_9672,N_7710);
and UO_39 (O_39,N_7962,N_7985);
or UO_40 (O_40,N_7871,N_7764);
and UO_41 (O_41,N_8100,N_8558);
nor UO_42 (O_42,N_7969,N_8258);
and UO_43 (O_43,N_8876,N_8698);
or UO_44 (O_44,N_8933,N_8359);
and UO_45 (O_45,N_9136,N_9970);
nor UO_46 (O_46,N_8655,N_9141);
nand UO_47 (O_47,N_9602,N_9289);
or UO_48 (O_48,N_9760,N_9046);
nand UO_49 (O_49,N_8390,N_9561);
nor UO_50 (O_50,N_8917,N_8565);
and UO_51 (O_51,N_9899,N_9573);
or UO_52 (O_52,N_8579,N_8470);
nand UO_53 (O_53,N_8304,N_7804);
nor UO_54 (O_54,N_9295,N_7755);
nor UO_55 (O_55,N_8653,N_8428);
nor UO_56 (O_56,N_7567,N_8136);
nand UO_57 (O_57,N_9469,N_9855);
nand UO_58 (O_58,N_8178,N_9127);
nor UO_59 (O_59,N_8027,N_9473);
and UO_60 (O_60,N_9846,N_7870);
and UO_61 (O_61,N_7572,N_9896);
or UO_62 (O_62,N_9942,N_8596);
and UO_63 (O_63,N_8766,N_7989);
and UO_64 (O_64,N_8623,N_9188);
nand UO_65 (O_65,N_9026,N_9546);
or UO_66 (O_66,N_8575,N_8603);
and UO_67 (O_67,N_8977,N_9729);
or UO_68 (O_68,N_8207,N_8229);
or UO_69 (O_69,N_8848,N_9116);
nand UO_70 (O_70,N_8402,N_9433);
nor UO_71 (O_71,N_7717,N_8355);
nand UO_72 (O_72,N_8619,N_8238);
nand UO_73 (O_73,N_7747,N_9211);
and UO_74 (O_74,N_9772,N_9304);
and UO_75 (O_75,N_7749,N_8348);
nor UO_76 (O_76,N_7992,N_9309);
nand UO_77 (O_77,N_7738,N_9025);
and UO_78 (O_78,N_8895,N_8367);
or UO_79 (O_79,N_9138,N_8076);
and UO_80 (O_80,N_7515,N_9769);
and UO_81 (O_81,N_9411,N_9373);
or UO_82 (O_82,N_9673,N_9283);
nor UO_83 (O_83,N_9778,N_8217);
and UO_84 (O_84,N_8869,N_8827);
or UO_85 (O_85,N_9944,N_9725);
and UO_86 (O_86,N_8863,N_8947);
nand UO_87 (O_87,N_7921,N_9441);
nand UO_88 (O_88,N_8731,N_9338);
or UO_89 (O_89,N_8971,N_8832);
or UO_90 (O_90,N_7922,N_8451);
nand UO_91 (O_91,N_8540,N_7792);
nand UO_92 (O_92,N_7598,N_8049);
nand UO_93 (O_93,N_9350,N_9869);
and UO_94 (O_94,N_8284,N_9627);
or UO_95 (O_95,N_7699,N_9832);
nand UO_96 (O_96,N_7984,N_9757);
nor UO_97 (O_97,N_8448,N_9206);
nand UO_98 (O_98,N_7865,N_8021);
or UO_99 (O_99,N_8545,N_7959);
nand UO_100 (O_100,N_8783,N_8530);
nor UO_101 (O_101,N_8400,N_7873);
and UO_102 (O_102,N_7835,N_9640);
and UO_103 (O_103,N_8997,N_9983);
nor UO_104 (O_104,N_8055,N_7787);
or UO_105 (O_105,N_9642,N_8440);
nand UO_106 (O_106,N_9424,N_9534);
or UO_107 (O_107,N_8148,N_7953);
or UO_108 (O_108,N_9496,N_7958);
nand UO_109 (O_109,N_8051,N_9487);
or UO_110 (O_110,N_7607,N_9464);
or UO_111 (O_111,N_8877,N_9887);
nor UO_112 (O_112,N_9108,N_8511);
or UO_113 (O_113,N_8068,N_7961);
nand UO_114 (O_114,N_8916,N_9785);
nor UO_115 (O_115,N_9299,N_7576);
nor UO_116 (O_116,N_9231,N_9964);
and UO_117 (O_117,N_8227,N_8059);
nor UO_118 (O_118,N_8852,N_9203);
nor UO_119 (O_119,N_7994,N_8910);
nor UO_120 (O_120,N_8250,N_9587);
or UO_121 (O_121,N_9799,N_9693);
nor UO_122 (O_122,N_7590,N_8855);
nand UO_123 (O_123,N_9315,N_8628);
or UO_124 (O_124,N_9875,N_8188);
nand UO_125 (O_125,N_9042,N_9916);
or UO_126 (O_126,N_7820,N_9296);
nor UO_127 (O_127,N_8341,N_9014);
nor UO_128 (O_128,N_8278,N_8667);
nand UO_129 (O_129,N_8761,N_9786);
nand UO_130 (O_130,N_9109,N_9213);
nand UO_131 (O_131,N_8981,N_9569);
and UO_132 (O_132,N_9824,N_8809);
nor UO_133 (O_133,N_7683,N_9683);
or UO_134 (O_134,N_8016,N_9761);
nand UO_135 (O_135,N_8210,N_8054);
nor UO_136 (O_136,N_7885,N_9645);
or UO_137 (O_137,N_8468,N_7838);
nand UO_138 (O_138,N_9189,N_8668);
nand UO_139 (O_139,N_9098,N_7650);
nand UO_140 (O_140,N_8953,N_9795);
and UO_141 (O_141,N_9200,N_9758);
and UO_142 (O_142,N_7601,N_7972);
nor UO_143 (O_143,N_9903,N_9531);
and UO_144 (O_144,N_9503,N_9142);
or UO_145 (O_145,N_9736,N_8241);
and UO_146 (O_146,N_9239,N_8275);
or UO_147 (O_147,N_8834,N_8097);
and UO_148 (O_148,N_9225,N_7848);
nor UO_149 (O_149,N_8962,N_8590);
nand UO_150 (O_150,N_9222,N_7739);
nand UO_151 (O_151,N_8677,N_7610);
nor UO_152 (O_152,N_9123,N_8563);
nor UO_153 (O_153,N_9608,N_8699);
or UO_154 (O_154,N_9449,N_9807);
and UO_155 (O_155,N_7622,N_9251);
nand UO_156 (O_156,N_9101,N_8967);
nand UO_157 (O_157,N_8138,N_7767);
and UO_158 (O_158,N_8621,N_9737);
nand UO_159 (O_159,N_9844,N_8700);
or UO_160 (O_160,N_7725,N_8899);
nand UO_161 (O_161,N_8568,N_9472);
and UO_162 (O_162,N_8972,N_7811);
nor UO_163 (O_163,N_9630,N_9963);
nand UO_164 (O_164,N_7704,N_7761);
nor UO_165 (O_165,N_8392,N_8356);
nand UO_166 (O_166,N_8649,N_7952);
or UO_167 (O_167,N_9180,N_9468);
nor UO_168 (O_168,N_9344,N_9484);
nand UO_169 (O_169,N_9417,N_9020);
and UO_170 (O_170,N_8990,N_9346);
nand UO_171 (O_171,N_8812,N_9985);
nand UO_172 (O_172,N_9860,N_8162);
nand UO_173 (O_173,N_8436,N_9245);
and UO_174 (O_174,N_8279,N_9360);
or UO_175 (O_175,N_9588,N_7971);
nand UO_176 (O_176,N_9646,N_7726);
or UO_177 (O_177,N_9670,N_7812);
and UO_178 (O_178,N_9518,N_9018);
or UO_179 (O_179,N_8332,N_9900);
nand UO_180 (O_180,N_8484,N_8574);
nand UO_181 (O_181,N_9380,N_9070);
or UO_182 (O_182,N_7654,N_8526);
and UO_183 (O_183,N_7852,N_8911);
nor UO_184 (O_184,N_7675,N_9183);
nor UO_185 (O_185,N_9764,N_8906);
nor UO_186 (O_186,N_9698,N_9389);
nor UO_187 (O_187,N_9481,N_7909);
nor UO_188 (O_188,N_9435,N_7617);
and UO_189 (O_189,N_7702,N_8544);
or UO_190 (O_190,N_9638,N_9146);
and UO_191 (O_191,N_9820,N_8339);
nor UO_192 (O_192,N_9652,N_8228);
and UO_193 (O_193,N_9864,N_7535);
and UO_194 (O_194,N_9741,N_8445);
and UO_195 (O_195,N_8312,N_8782);
or UO_196 (O_196,N_9654,N_8706);
or UO_197 (O_197,N_7892,N_8150);
and UO_198 (O_198,N_8888,N_8662);
nor UO_199 (O_199,N_9049,N_7942);
and UO_200 (O_200,N_7967,N_9447);
or UO_201 (O_201,N_9811,N_9984);
nand UO_202 (O_202,N_7529,N_8331);
or UO_203 (O_203,N_8318,N_7540);
or UO_204 (O_204,N_7554,N_9898);
or UO_205 (O_205,N_8363,N_9656);
and UO_206 (O_206,N_9462,N_8551);
or UO_207 (O_207,N_8104,N_8719);
nand UO_208 (O_208,N_7908,N_7730);
and UO_209 (O_209,N_9885,N_8158);
nand UO_210 (O_210,N_8401,N_9694);
or UO_211 (O_211,N_9514,N_9612);
or UO_212 (O_212,N_9374,N_9710);
and UO_213 (O_213,N_8319,N_7779);
nand UO_214 (O_214,N_8276,N_8062);
nor UO_215 (O_215,N_9437,N_9094);
and UO_216 (O_216,N_8893,N_9884);
nand UO_217 (O_217,N_8920,N_8815);
or UO_218 (O_218,N_8270,N_7839);
and UO_219 (O_219,N_7816,N_8516);
and UO_220 (O_220,N_9544,N_8583);
nor UO_221 (O_221,N_9133,N_7772);
nor UO_222 (O_222,N_8773,N_9524);
or UO_223 (O_223,N_8769,N_9621);
nor UO_224 (O_224,N_8539,N_8810);
nor UO_225 (O_225,N_9099,N_8465);
nor UO_226 (O_226,N_8758,N_8277);
nand UO_227 (O_227,N_7899,N_9474);
nand UO_228 (O_228,N_9781,N_8721);
or UO_229 (O_229,N_7603,N_8541);
and UO_230 (O_230,N_8446,N_9106);
and UO_231 (O_231,N_7823,N_8447);
and UO_232 (O_232,N_9738,N_8161);
nand UO_233 (O_233,N_9696,N_8976);
nor UO_234 (O_234,N_9798,N_9812);
nand UO_235 (O_235,N_8472,N_8930);
or UO_236 (O_236,N_7874,N_8065);
or UO_237 (O_237,N_9162,N_9614);
and UO_238 (O_238,N_9639,N_8866);
or UO_239 (O_239,N_8956,N_8125);
nor UO_240 (O_240,N_8842,N_7679);
or UO_241 (O_241,N_8416,N_7648);
or UO_242 (O_242,N_9731,N_9998);
nand UO_243 (O_243,N_9691,N_9671);
and UO_244 (O_244,N_9706,N_8555);
nor UO_245 (O_245,N_8582,N_9298);
nor UO_246 (O_246,N_9529,N_7932);
and UO_247 (O_247,N_9396,N_7748);
or UO_248 (O_248,N_9540,N_9692);
nor UO_249 (O_249,N_7732,N_8643);
or UO_250 (O_250,N_9782,N_8747);
nand UO_251 (O_251,N_7980,N_9332);
nand UO_252 (O_252,N_8708,N_9695);
nand UO_253 (O_253,N_9904,N_7933);
or UO_254 (O_254,N_8231,N_9689);
nor UO_255 (O_255,N_9556,N_8352);
nand UO_256 (O_256,N_8072,N_9072);
nor UO_257 (O_257,N_9443,N_9960);
nand UO_258 (O_258,N_9011,N_9385);
nand UO_259 (O_259,N_9023,N_7805);
and UO_260 (O_260,N_7623,N_9063);
nor UO_261 (O_261,N_9143,N_7813);
nor UO_262 (O_262,N_8715,N_7797);
nor UO_263 (O_263,N_9925,N_9132);
nor UO_264 (O_264,N_9300,N_8473);
nor UO_265 (O_265,N_7541,N_9651);
xnor UO_266 (O_266,N_9905,N_7580);
nand UO_267 (O_267,N_8638,N_8095);
nor UO_268 (O_268,N_8903,N_8743);
or UO_269 (O_269,N_9908,N_8265);
or UO_270 (O_270,N_8393,N_8196);
and UO_271 (O_271,N_9940,N_9618);
nand UO_272 (O_272,N_7819,N_9552);
nand UO_273 (O_273,N_7731,N_9831);
and UO_274 (O_274,N_7568,N_8042);
nand UO_275 (O_275,N_9452,N_9954);
or UO_276 (O_276,N_8673,N_8867);
nand UO_277 (O_277,N_9248,N_9575);
nand UO_278 (O_278,N_8133,N_8140);
and UO_279 (O_279,N_9230,N_7734);
nand UO_280 (O_280,N_7737,N_7524);
nand UO_281 (O_281,N_8285,N_9793);
and UO_282 (O_282,N_9148,N_9278);
nand UO_283 (O_283,N_8680,N_9705);
nand UO_284 (O_284,N_8248,N_7954);
nor UO_285 (O_285,N_9322,N_7509);
or UO_286 (O_286,N_7631,N_7864);
nor UO_287 (O_287,N_8588,N_9616);
nor UO_288 (O_288,N_9093,N_8198);
and UO_289 (O_289,N_7759,N_9595);
nor UO_290 (O_290,N_8658,N_9120);
and UO_291 (O_291,N_7740,N_7990);
and UO_292 (O_292,N_8159,N_9359);
or UO_293 (O_293,N_8324,N_9913);
and UO_294 (O_294,N_7894,N_8195);
nand UO_295 (O_295,N_8491,N_8508);
nor UO_296 (O_296,N_7685,N_9922);
nor UO_297 (O_297,N_8991,N_7707);
nand UO_298 (O_298,N_8115,N_7709);
nand UO_299 (O_299,N_9456,N_9323);
nor UO_300 (O_300,N_9247,N_8547);
and UO_301 (O_301,N_9862,N_7620);
nor UO_302 (O_302,N_9436,N_9947);
and UO_303 (O_303,N_8651,N_7914);
nor UO_304 (O_304,N_8129,N_9677);
or UO_305 (O_305,N_8950,N_9003);
and UO_306 (O_306,N_8108,N_7630);
and UO_307 (O_307,N_9131,N_8755);
and UO_308 (O_308,N_9301,N_9551);
nand UO_309 (O_309,N_7831,N_8892);
nor UO_310 (O_310,N_7766,N_7564);
nor UO_311 (O_311,N_9305,N_8414);
nor UO_312 (O_312,N_9220,N_8124);
or UO_313 (O_313,N_8366,N_9010);
or UO_314 (O_314,N_8625,N_8650);
and UO_315 (O_315,N_8796,N_9647);
nor UO_316 (O_316,N_8498,N_8439);
nor UO_317 (O_317,N_8695,N_7987);
nand UO_318 (O_318,N_7575,N_9229);
or UO_319 (O_319,N_8992,N_8461);
or UO_320 (O_320,N_8007,N_7505);
and UO_321 (O_321,N_9721,N_9157);
nand UO_322 (O_322,N_9166,N_9517);
or UO_323 (O_323,N_8800,N_8120);
nand UO_324 (O_324,N_9083,N_8028);
or UO_325 (O_325,N_8382,N_9815);
nand UO_326 (O_326,N_9366,N_9348);
and UO_327 (O_327,N_8806,N_9613);
or UO_328 (O_328,N_9177,N_9792);
and UO_329 (O_329,N_8531,N_9066);
nand UO_330 (O_330,N_9961,N_8252);
nand UO_331 (O_331,N_9990,N_9412);
nand UO_332 (O_332,N_9485,N_9941);
or UO_333 (O_333,N_8083,N_7521);
and UO_334 (O_334,N_7794,N_8576);
or UO_335 (O_335,N_7807,N_9075);
and UO_336 (O_336,N_9906,N_7999);
nand UO_337 (O_337,N_8580,N_9504);
nand UO_338 (O_338,N_9586,N_9833);
or UO_339 (O_339,N_8594,N_8626);
and UO_340 (O_340,N_8149,N_9653);
or UO_341 (O_341,N_7964,N_9851);
nor UO_342 (O_342,N_9314,N_8752);
or UO_343 (O_343,N_7851,N_8426);
nand UO_344 (O_344,N_9037,N_7532);
nor UO_345 (O_345,N_9372,N_7927);
and UO_346 (O_346,N_7676,N_9606);
nor UO_347 (O_347,N_7522,N_8040);
nor UO_348 (O_348,N_8281,N_7955);
nand UO_349 (O_349,N_9784,N_9221);
or UO_350 (O_350,N_9153,N_7960);
nor UO_351 (O_351,N_7700,N_8602);
nor UO_352 (O_352,N_9973,N_9949);
and UO_353 (O_353,N_8074,N_7713);
nor UO_354 (O_354,N_9926,N_9419);
nor UO_355 (O_355,N_9604,N_9628);
and UO_356 (O_356,N_9664,N_9726);
and UO_357 (O_357,N_9880,N_8884);
nor UO_358 (O_358,N_7667,N_7910);
nand UO_359 (O_359,N_9482,N_7784);
and UO_360 (O_360,N_8690,N_8767);
nand UO_361 (O_361,N_8894,N_8882);
and UO_362 (O_362,N_9865,N_9490);
nor UO_363 (O_363,N_8288,N_7586);
nor UO_364 (O_364,N_8734,N_8959);
nor UO_365 (O_365,N_8487,N_8194);
nand UO_366 (O_366,N_8182,N_8163);
nor UO_367 (O_367,N_7934,N_8837);
nand UO_368 (O_368,N_9173,N_9434);
or UO_369 (O_369,N_9246,N_8689);
nor UO_370 (O_370,N_8631,N_9713);
nand UO_371 (O_371,N_7658,N_7790);
or UO_372 (O_372,N_9717,N_8119);
and UO_373 (O_373,N_9345,N_7565);
or UO_374 (O_374,N_9467,N_9387);
or UO_375 (O_375,N_9545,N_7775);
nor UO_376 (O_376,N_9988,N_9825);
nand UO_377 (O_377,N_8504,N_9543);
or UO_378 (O_378,N_9102,N_7657);
or UO_379 (O_379,N_8020,N_8383);
nand UO_380 (O_380,N_9152,N_9835);
and UO_381 (O_381,N_7834,N_9410);
or UO_382 (O_382,N_9267,N_8750);
and UO_383 (O_383,N_8024,N_7822);
or UO_384 (O_384,N_9365,N_9596);
or UO_385 (O_385,N_8063,N_9006);
nor UO_386 (O_386,N_9353,N_8493);
and UO_387 (O_387,N_9069,N_7507);
nand UO_388 (O_388,N_7853,N_9261);
nor UO_389 (O_389,N_8984,N_7665);
and UO_390 (O_390,N_7881,N_8875);
and UO_391 (O_391,N_8881,N_9938);
and UO_392 (O_392,N_8050,N_8190);
nor UO_393 (O_393,N_9891,N_8529);
nand UO_394 (O_394,N_8396,N_7993);
nand UO_395 (O_395,N_9787,N_8897);
nand UO_396 (O_396,N_8514,N_9828);
or UO_397 (O_397,N_8441,N_9994);
or UO_398 (O_398,N_9956,N_8728);
nor UO_399 (O_399,N_9535,N_8840);
nor UO_400 (O_400,N_9740,N_8425);
nand UO_401 (O_401,N_8898,N_7946);
nor UO_402 (O_402,N_7979,N_7770);
nand UO_403 (O_403,N_9617,N_7893);
nand UO_404 (O_404,N_9107,N_8957);
nand UO_405 (O_405,N_9428,N_8586);
or UO_406 (O_406,N_9675,N_8116);
or UO_407 (O_407,N_9796,N_7600);
nand UO_408 (O_408,N_8543,N_7581);
or UO_409 (O_409,N_8336,N_9145);
nand UO_410 (O_410,N_7528,N_9933);
and UO_411 (O_411,N_8942,N_8458);
nand UO_412 (O_412,N_8137,N_9512);
nor UO_413 (O_413,N_8670,N_9397);
nand UO_414 (O_414,N_8527,N_9242);
or UO_415 (O_415,N_8176,N_9771);
nor UO_416 (O_416,N_9684,N_8372);
and UO_417 (O_417,N_8936,N_9803);
nor UO_418 (O_418,N_7588,N_8510);
or UO_419 (O_419,N_9147,N_7796);
nor UO_420 (O_420,N_9937,N_8034);
nand UO_421 (O_421,N_9499,N_8045);
and UO_422 (O_422,N_9732,N_9883);
nand UO_423 (O_423,N_9001,N_8488);
nor UO_424 (O_424,N_9746,N_9215);
nand UO_425 (O_425,N_9789,N_9182);
and UO_426 (O_426,N_8453,N_8033);
or UO_427 (O_427,N_8494,N_9021);
and UO_428 (O_428,N_9530,N_8298);
nor UO_429 (O_429,N_9742,N_7696);
and UO_430 (O_430,N_8406,N_8036);
xnor UO_431 (O_431,N_7947,N_9282);
and UO_432 (O_432,N_9307,N_9897);
nor UO_433 (O_433,N_7756,N_7693);
nor UO_434 (O_434,N_7956,N_8904);
nor UO_435 (O_435,N_9165,N_7597);
nand UO_436 (O_436,N_9273,N_9505);
nand UO_437 (O_437,N_8814,N_8139);
nand UO_438 (O_438,N_9407,N_8342);
or UO_439 (O_439,N_9598,N_7976);
or UO_440 (O_440,N_7688,N_9129);
or UO_441 (O_441,N_8532,N_9872);
or UO_442 (O_442,N_7968,N_8146);
nand UO_443 (O_443,N_8092,N_9939);
and UO_444 (O_444,N_9406,N_8986);
and UO_445 (O_445,N_9997,N_9124);
nor UO_446 (O_446,N_8693,N_7793);
and UO_447 (O_447,N_9414,N_9032);
nor UO_448 (O_448,N_8932,N_7841);
or UO_449 (O_449,N_8457,N_7558);
and UO_450 (O_450,N_9212,N_8128);
nand UO_451 (O_451,N_9583,N_9889);
nand UO_452 (O_452,N_9802,N_9678);
or UO_453 (O_453,N_9493,N_8987);
and UO_454 (O_454,N_7563,N_9558);
and UO_455 (O_455,N_9272,N_8317);
or UO_456 (O_456,N_9704,N_8310);
nor UO_457 (O_457,N_8171,N_8391);
or UO_458 (O_458,N_9376,N_9306);
nor UO_459 (O_459,N_8760,N_9680);
nand UO_460 (O_460,N_9868,N_8931);
or UO_461 (O_461,N_8014,N_8192);
nor UO_462 (O_462,N_9915,N_8325);
and UO_463 (O_463,N_9111,N_8927);
nor UO_464 (O_464,N_8887,N_9364);
nor UO_465 (O_465,N_8778,N_9119);
xnor UO_466 (O_466,N_9641,N_7795);
nor UO_467 (O_467,N_9114,N_9489);
nor UO_468 (O_468,N_8168,N_8569);
and UO_469 (O_469,N_7869,N_9056);
nor UO_470 (O_470,N_8320,N_9592);
nand UO_471 (O_471,N_8785,N_7846);
nand UO_472 (O_472,N_8422,N_7750);
and UO_473 (O_473,N_9405,N_8041);
nand UO_474 (O_474,N_8245,N_9228);
nor UO_475 (O_475,N_7856,N_9402);
and UO_476 (O_476,N_7924,N_8157);
nand UO_477 (O_477,N_8272,N_8787);
or UO_478 (O_478,N_9559,N_9666);
nor UO_479 (O_479,N_8013,N_8101);
and UO_480 (O_480,N_8587,N_8513);
or UO_481 (O_481,N_9470,N_9522);
nand UO_482 (O_482,N_9655,N_9912);
and UO_483 (O_483,N_7788,N_9565);
nor UO_484 (O_484,N_9058,N_8703);
and UO_485 (O_485,N_8219,N_7983);
or UO_486 (O_486,N_8346,N_7682);
or UO_487 (O_487,N_7608,N_9650);
and UO_488 (O_488,N_9574,N_7878);
or UO_489 (O_489,N_8521,N_9176);
nor UO_490 (O_490,N_8349,N_8296);
or UO_491 (O_491,N_8975,N_8857);
or UO_492 (O_492,N_8466,N_9386);
nor UO_493 (O_493,N_8813,N_7680);
nand UO_494 (O_494,N_7543,N_8710);
and UO_495 (O_495,N_9398,N_9699);
nand UO_496 (O_496,N_8824,N_8823);
or UO_497 (O_497,N_9399,N_8561);
nor UO_498 (O_498,N_8323,N_8454);
nor UO_499 (O_499,N_9975,N_9000);
nor UO_500 (O_500,N_7527,N_7917);
or UO_501 (O_501,N_9395,N_9682);
or UO_502 (O_502,N_7629,N_9777);
nand UO_503 (O_503,N_7723,N_8672);
nor UO_504 (O_504,N_9290,N_9202);
nand UO_505 (O_505,N_7826,N_8993);
and UO_506 (O_506,N_9810,N_9840);
and UO_507 (O_507,N_9330,N_9594);
xnor UO_508 (O_508,N_9708,N_9763);
or UO_509 (O_509,N_8633,N_9055);
or UO_510 (O_510,N_9814,N_9371);
and UO_511 (O_511,N_8057,N_9084);
nand UO_512 (O_512,N_7855,N_8641);
nand UO_513 (O_513,N_7579,N_8273);
or UO_514 (O_514,N_7647,N_8232);
and UO_515 (O_515,N_8333,N_8966);
nand UO_516 (O_516,N_9232,N_9553);
and UO_517 (O_517,N_8557,N_9920);
nor UO_518 (O_518,N_7988,N_9748);
nor UO_519 (O_519,N_9224,N_7808);
nor UO_520 (O_520,N_8535,N_7664);
or UO_521 (O_521,N_9509,N_9415);
and UO_522 (O_522,N_8839,N_9266);
nand UO_523 (O_523,N_8242,N_8327);
nor UO_524 (O_524,N_9836,N_7714);
nand UO_525 (O_525,N_9486,N_9064);
nand UO_526 (O_526,N_7890,N_7633);
nor UO_527 (O_527,N_8314,N_9770);
nand UO_528 (O_528,N_9800,N_8929);
nand UO_529 (O_529,N_9702,N_7503);
nand UO_530 (O_530,N_8682,N_7857);
or UO_531 (O_531,N_7780,N_8338);
and UO_532 (O_532,N_8481,N_8740);
nor UO_533 (O_533,N_7951,N_8556);
nor UO_534 (O_534,N_8365,N_7897);
or UO_535 (O_535,N_9513,N_8896);
and UO_536 (O_536,N_9537,N_8263);
nand UO_537 (O_537,N_9186,N_9174);
and UO_538 (O_538,N_9313,N_8830);
and UO_539 (O_539,N_8648,N_8343);
or UO_540 (O_540,N_8253,N_7926);
nand UO_541 (O_541,N_9845,N_9091);
or UO_542 (O_542,N_9674,N_9775);
nor UO_543 (O_543,N_8079,N_8674);
nand UO_544 (O_544,N_8502,N_7520);
or UO_545 (O_545,N_8417,N_7599);
and UO_546 (O_546,N_9035,N_7801);
nand UO_547 (O_547,N_7902,N_8524);
or UO_548 (O_548,N_9269,N_7642);
nor UO_549 (O_549,N_8746,N_8751);
nand UO_550 (O_550,N_9599,N_8404);
nor UO_551 (O_551,N_9325,N_7868);
nor UO_552 (O_552,N_7937,N_9762);
or UO_553 (O_553,N_8053,N_7830);
nand UO_554 (O_554,N_9542,N_8878);
nor UO_555 (O_555,N_8889,N_8452);
and UO_556 (O_556,N_8130,N_9714);
and UO_557 (O_557,N_8553,N_7814);
nand UO_558 (O_558,N_8890,N_7641);
and UO_559 (O_559,N_8560,N_9105);
nand UO_560 (O_560,N_8723,N_8089);
and UO_561 (O_561,N_7957,N_7587);
and UO_562 (O_562,N_8784,N_8608);
nand UO_563 (O_563,N_8326,N_8381);
nand UO_564 (O_564,N_8047,N_8085);
or UO_565 (O_565,N_9852,N_8435);
and UO_566 (O_566,N_7765,N_9377);
nor UO_567 (O_567,N_9571,N_8838);
or UO_568 (O_568,N_9209,N_9172);
nand UO_569 (O_569,N_8805,N_8449);
and UO_570 (O_570,N_9488,N_9375);
nor UO_571 (O_571,N_9525,N_8191);
nor UO_572 (O_572,N_8518,N_7975);
or UO_573 (O_573,N_8202,N_9155);
and UO_574 (O_574,N_9062,N_9404);
or UO_575 (O_575,N_9520,N_8147);
or UO_576 (O_576,N_7502,N_7534);
nand UO_577 (O_577,N_8803,N_8951);
nor UO_578 (O_578,N_9607,N_9707);
nor UO_579 (O_579,N_8604,N_7945);
or UO_580 (O_580,N_9027,N_8069);
nand UO_581 (O_581,N_9936,N_8850);
nor UO_582 (O_582,N_8358,N_8012);
nor UO_583 (O_583,N_9626,N_7690);
nand UO_584 (O_584,N_8073,N_8858);
or UO_585 (O_585,N_8483,N_7661);
and UO_586 (O_586,N_7546,N_7781);
nand UO_587 (O_587,N_9199,N_9079);
nand UO_588 (O_588,N_7694,N_9252);
or UO_589 (O_589,N_9663,N_8395);
nor UO_590 (O_590,N_9593,N_9311);
and UO_591 (O_591,N_8038,N_8614);
nor UO_592 (O_592,N_7655,N_8409);
nand UO_593 (O_593,N_9491,N_9050);
nand UO_594 (O_594,N_8434,N_8578);
and UO_595 (O_595,N_8635,N_9264);
nand UO_596 (O_596,N_9363,N_9629);
nand UO_597 (O_597,N_9051,N_9722);
nand UO_598 (O_598,N_8056,N_9805);
nand UO_599 (O_599,N_7901,N_7569);
or UO_600 (O_600,N_7836,N_9033);
or UO_601 (O_601,N_9057,N_7778);
or UO_602 (O_602,N_9801,N_9951);
nand UO_603 (O_603,N_8479,N_8663);
nand UO_604 (O_604,N_9847,N_8118);
or UO_605 (O_605,N_8988,N_9430);
and UO_606 (O_606,N_8572,N_7776);
and UO_607 (O_607,N_8462,N_8819);
and UO_608 (O_608,N_7653,N_7777);
nand UO_609 (O_609,N_7845,N_7619);
nor UO_610 (O_610,N_9210,N_7555);
nand UO_611 (O_611,N_8717,N_8093);
nor UO_612 (O_612,N_7919,N_9818);
nand UO_613 (O_613,N_8251,N_9268);
or UO_614 (O_614,N_7718,N_7741);
nand UO_615 (O_615,N_9223,N_9019);
nor UO_616 (O_616,N_9347,N_8066);
nand UO_617 (O_617,N_8738,N_8718);
and UO_618 (O_618,N_9910,N_8201);
xnor UO_619 (O_619,N_9822,N_7743);
nor UO_620 (O_620,N_8921,N_7666);
nand UO_621 (O_621,N_7640,N_8291);
and UO_622 (O_622,N_9190,N_7525);
nand UO_623 (O_623,N_9369,N_7621);
nand UO_624 (O_624,N_9358,N_8968);
and UO_625 (O_625,N_7783,N_9902);
or UO_626 (O_626,N_7512,N_9877);
or UO_627 (O_627,N_7785,N_9539);
nand UO_628 (O_628,N_7553,N_7757);
nand UO_629 (O_629,N_7504,N_8601);
xnor UO_630 (O_630,N_8442,N_7637);
nor UO_631 (O_631,N_7516,N_9611);
nor UO_632 (O_632,N_9361,N_9349);
and UO_633 (O_633,N_9584,N_8864);
or UO_634 (O_634,N_9039,N_9863);
nor UO_635 (O_635,N_9334,N_9751);
nor UO_636 (O_636,N_8088,N_9041);
nor UO_637 (O_637,N_7900,N_7977);
or UO_638 (O_638,N_7501,N_9843);
nor UO_639 (O_639,N_9337,N_9012);
nor UO_640 (O_640,N_9492,N_7923);
and UO_641 (O_641,N_8705,N_7651);
or UO_642 (O_642,N_9275,N_9408);
nor UO_643 (O_643,N_8862,N_7941);
or UO_644 (O_644,N_8172,N_9909);
nor UO_645 (O_645,N_9002,N_8820);
nor UO_646 (O_646,N_8167,N_9128);
or UO_647 (O_647,N_8595,N_8497);
and UO_648 (O_648,N_8776,N_8011);
and UO_649 (O_649,N_8683,N_8567);
nand UO_650 (O_650,N_9590,N_7809);
and UO_651 (O_651,N_8259,N_8505);
and UO_652 (O_652,N_9187,N_8405);
or UO_653 (O_653,N_8353,N_8109);
nand UO_654 (O_654,N_8046,N_8193);
or UO_655 (O_655,N_8902,N_9163);
and UO_656 (O_656,N_9343,N_9716);
and UO_657 (O_657,N_9427,N_8536);
nand UO_658 (O_658,N_8794,N_9719);
nor UO_659 (O_659,N_9959,N_7966);
and UO_660 (O_660,N_8306,N_9029);
or UO_661 (O_661,N_8105,N_8702);
nor UO_662 (O_662,N_9867,N_7905);
and UO_663 (O_663,N_9685,N_7719);
or UO_664 (O_664,N_7500,N_9088);
and UO_665 (O_665,N_8692,N_8132);
and UO_666 (O_666,N_9515,N_9533);
and UO_667 (O_667,N_8712,N_7896);
and UO_668 (O_668,N_9658,N_9297);
or UO_669 (O_669,N_9243,N_9048);
or UO_670 (O_670,N_9160,N_7549);
nor UO_671 (O_671,N_8883,N_7545);
and UO_672 (O_672,N_9995,N_7884);
or UO_673 (O_673,N_9977,N_8924);
and UO_674 (O_674,N_7913,N_7824);
or UO_675 (O_675,N_8610,N_9161);
nand UO_676 (O_676,N_9576,N_8996);
nor UO_677 (O_677,N_8963,N_7891);
nor UO_678 (O_678,N_9316,N_8311);
and UO_679 (O_679,N_8160,N_9390);
nor UO_680 (O_680,N_9310,N_8225);
and UO_681 (O_681,N_9103,N_8022);
nor UO_682 (O_682,N_9755,N_7907);
and UO_683 (O_683,N_7763,N_9958);
xor UO_684 (O_684,N_8745,N_7948);
and UO_685 (O_685,N_9071,N_9917);
or UO_686 (O_686,N_8865,N_7701);
and UO_687 (O_687,N_9422,N_8937);
or UO_688 (O_688,N_9204,N_8922);
nand UO_689 (O_689,N_8500,N_7506);
or UO_690 (O_690,N_9989,N_7578);
or UO_691 (O_691,N_8691,N_7963);
and UO_692 (O_692,N_8600,N_7526);
nand UO_693 (O_693,N_8843,N_9319);
and UO_694 (O_694,N_9874,N_9089);
nand UO_695 (O_695,N_7827,N_7887);
nand UO_696 (O_696,N_7513,N_9393);
nand UO_697 (O_697,N_8570,N_9955);
or UO_698 (O_698,N_9850,N_9620);
and UO_699 (O_699,N_7903,N_9317);
or UO_700 (O_700,N_8283,N_9842);
nor UO_701 (O_701,N_9164,N_8666);
and UO_702 (O_702,N_7875,N_8039);
nor UO_703 (O_703,N_9734,N_7791);
nand UO_704 (O_704,N_8552,N_8015);
or UO_705 (O_705,N_8111,N_8629);
nand UO_706 (O_706,N_8037,N_9550);
nand UO_707 (O_707,N_8913,N_8205);
nor UO_708 (O_708,N_8995,N_7715);
nor UO_709 (O_709,N_8714,N_7645);
nor UO_710 (O_710,N_9700,N_8008);
or UO_711 (O_711,N_7753,N_8874);
nor UO_712 (O_712,N_9078,N_9191);
or UO_713 (O_713,N_8236,N_9004);
nand UO_714 (O_714,N_7867,N_9834);
and UO_715 (O_715,N_7998,N_7612);
and UO_716 (O_716,N_9506,N_8926);
and UO_717 (O_717,N_9420,N_9724);
nor UO_718 (O_718,N_8009,N_7930);
or UO_719 (O_719,N_7721,N_8707);
nand UO_720 (O_720,N_7911,N_7678);
and UO_721 (O_721,N_8846,N_7832);
or UO_722 (O_722,N_8763,N_8742);
or UO_723 (O_723,N_9712,N_9097);
and UO_724 (O_724,N_9015,N_9632);
or UO_725 (O_725,N_7806,N_8155);
nor UO_726 (O_726,N_8460,N_8153);
and UO_727 (O_727,N_9028,N_7544);
nor UO_728 (O_728,N_9987,N_8989);
and UO_729 (O_729,N_8098,N_8301);
or UO_730 (O_730,N_8969,N_7754);
nor UO_731 (O_731,N_8455,N_9808);
nand UO_732 (O_732,N_8661,N_8934);
nor UO_733 (O_733,N_8928,N_8135);
nor UO_734 (O_734,N_9362,N_9381);
nand UO_735 (O_735,N_8960,N_8925);
or UO_736 (O_736,N_9779,N_7720);
and UO_737 (O_737,N_7644,N_9331);
or UO_738 (O_738,N_8528,N_8102);
and UO_739 (O_739,N_9439,N_8660);
and UO_740 (O_740,N_9125,N_7605);
nand UO_741 (O_741,N_8423,N_8585);
nand UO_742 (O_742,N_9541,N_8271);
or UO_743 (O_743,N_9036,N_8308);
nor UO_744 (O_744,N_9701,N_8260);
nor UO_745 (O_745,N_9379,N_8211);
nand UO_746 (O_746,N_9681,N_7895);
or UO_747 (O_747,N_7523,N_8156);
and UO_748 (O_748,N_8816,N_7872);
xor UO_749 (O_749,N_9856,N_9999);
nand UO_750 (O_750,N_8912,N_9827);
nand UO_751 (O_751,N_7613,N_9329);
nor UO_752 (O_752,N_9752,N_7925);
nor UO_753 (O_753,N_9455,N_9554);
nor UO_754 (O_754,N_8938,N_8744);
nor UO_755 (O_755,N_9619,N_9355);
and UO_756 (O_756,N_9285,N_9214);
and UO_757 (O_757,N_8389,N_8117);
nand UO_758 (O_758,N_7880,N_7508);
nand UO_759 (O_759,N_8257,N_9580);
and UO_760 (O_760,N_9333,N_9293);
nor UO_761 (O_761,N_8152,N_8851);
nand UO_762 (O_762,N_8321,N_8052);
nor UO_763 (O_763,N_8123,N_7689);
or UO_764 (O_764,N_7821,N_9871);
and UO_765 (O_765,N_8078,N_9356);
nand UO_766 (O_766,N_9876,N_7638);
or UO_767 (O_767,N_8330,N_7639);
nand UO_768 (O_768,N_8412,N_8371);
nor UO_769 (O_769,N_8607,N_8573);
nand UO_770 (O_770,N_8685,N_9817);
nand UO_771 (O_771,N_8274,N_9813);
or UO_772 (O_772,N_9723,N_8645);
and UO_773 (O_773,N_9783,N_9277);
nor UO_774 (O_774,N_9788,N_8090);
and UO_775 (O_775,N_9260,N_9532);
nor UO_776 (O_776,N_9388,N_9624);
and UO_777 (O_777,N_9054,N_8185);
or UO_778 (O_778,N_9965,N_9235);
and UO_779 (O_779,N_9837,N_9643);
and UO_780 (O_780,N_7712,N_8727);
nor UO_781 (O_781,N_9341,N_9982);
nor UO_782 (O_782,N_7609,N_8939);
or UO_783 (O_783,N_8980,N_8733);
or UO_784 (O_784,N_9578,N_8944);
and UO_785 (O_785,N_7810,N_8375);
nor UO_786 (O_786,N_8833,N_9450);
nand UO_787 (O_787,N_8430,N_8143);
or UO_788 (O_788,N_7752,N_8949);
nor UO_789 (O_789,N_9637,N_9024);
or UO_790 (O_790,N_9819,N_8154);
and UO_791 (O_791,N_8164,N_7577);
nor UO_792 (O_792,N_8467,N_9766);
and UO_793 (O_793,N_9384,N_9463);
or UO_794 (O_794,N_9858,N_9657);
nor UO_795 (O_795,N_9631,N_9809);
nor UO_796 (O_796,N_9413,N_9197);
nand UO_797 (O_797,N_8808,N_9254);
xnor UO_798 (O_798,N_8520,N_7912);
nand UO_799 (O_799,N_9043,N_7660);
nor UO_800 (O_800,N_7627,N_7518);
nor UO_801 (O_801,N_7519,N_8373);
or UO_802 (O_802,N_9237,N_8480);
or UO_803 (O_803,N_8303,N_9914);
nand UO_804 (O_804,N_9950,N_9005);
nand UO_805 (O_805,N_9357,N_7997);
or UO_806 (O_806,N_8943,N_9320);
nand UO_807 (O_807,N_7888,N_9193);
nor UO_808 (O_808,N_9194,N_9442);
or UO_809 (O_809,N_9882,N_9841);
or UO_810 (O_810,N_8286,N_8550);
xor UO_811 (O_811,N_8031,N_8795);
nor UO_812 (O_812,N_9418,N_8444);
nand UO_813 (O_813,N_7582,N_8345);
and UO_814 (O_814,N_7674,N_8907);
or UO_815 (O_815,N_8329,N_8671);
and UO_816 (O_816,N_7510,N_8035);
nand UO_817 (O_817,N_9676,N_8189);
nor UO_818 (O_818,N_9548,N_9564);
nor UO_819 (O_819,N_7920,N_7589);
nand UO_820 (O_820,N_9797,N_7995);
nand UO_821 (O_821,N_8534,N_9423);
nand UO_822 (O_822,N_9502,N_8106);
or UO_823 (O_823,N_8010,N_9547);
nand UO_824 (O_824,N_9073,N_7594);
and UO_825 (O_825,N_7557,N_7840);
nand UO_826 (O_826,N_7928,N_7671);
nor UO_827 (O_827,N_8519,N_8598);
or UO_828 (O_828,N_7842,N_8611);
or UO_829 (O_829,N_8915,N_8485);
nor UO_830 (O_830,N_7786,N_9555);
nand UO_831 (O_831,N_8584,N_7705);
or UO_832 (O_832,N_8591,N_9953);
nand UO_833 (O_833,N_8780,N_9255);
nor UO_834 (O_834,N_8096,N_9971);
nor UO_835 (O_835,N_7659,N_7986);
nor UO_836 (O_836,N_8187,N_9928);
nand UO_837 (O_837,N_8781,N_9401);
and UO_838 (O_838,N_8340,N_8676);
xor UO_839 (O_839,N_7592,N_9244);
or UO_840 (O_840,N_7548,N_9471);
nand UO_841 (O_841,N_7833,N_9403);
nor UO_842 (O_842,N_8026,N_9536);
nor UO_843 (O_843,N_9718,N_8474);
and UO_844 (O_844,N_9625,N_8091);
and UO_845 (O_845,N_9735,N_9816);
and UO_846 (O_846,N_8184,N_9562);
or UO_847 (O_847,N_8268,N_9567);
nor UO_848 (O_848,N_8000,N_7550);
and UO_849 (O_849,N_8017,N_9894);
nor UO_850 (O_850,N_7531,N_9234);
nor UO_851 (O_851,N_8630,N_8764);
or UO_852 (O_852,N_9986,N_9233);
or UO_853 (O_853,N_7818,N_8644);
xor UO_854 (O_854,N_8398,N_9067);
and UO_855 (O_855,N_8537,N_9258);
or UO_856 (O_856,N_8110,N_8822);
and UO_857 (O_857,N_8978,N_8679);
or UO_858 (O_858,N_8974,N_8646);
nor UO_859 (O_859,N_7828,N_9154);
or UO_860 (O_860,N_8686,N_9560);
and UO_861 (O_861,N_7760,N_9292);
and UO_862 (O_862,N_8517,N_8459);
and UO_863 (O_863,N_9185,N_9687);
and UO_864 (O_864,N_9321,N_8141);
or UO_865 (O_865,N_8793,N_8233);
or UO_866 (O_866,N_8798,N_7614);
and UO_867 (O_867,N_9516,N_7799);
or UO_868 (O_868,N_8082,N_7606);
nand UO_869 (O_869,N_8859,N_8994);
or UO_870 (O_870,N_9171,N_9167);
and UO_871 (O_871,N_8985,N_7602);
nand UO_872 (O_872,N_8269,N_7991);
or UO_873 (O_873,N_9259,N_9168);
and UO_874 (O_874,N_8564,N_8818);
nand UO_875 (O_875,N_8335,N_8144);
and UO_876 (O_876,N_8624,N_9216);
and UO_877 (O_877,N_8503,N_9523);
xor UO_878 (O_878,N_7906,N_8239);
or UO_879 (O_879,N_8941,N_7566);
nor UO_880 (O_880,N_9218,N_8387);
or UO_881 (O_881,N_9886,N_9743);
nand UO_882 (O_882,N_9568,N_8515);
nor UO_883 (O_883,N_9597,N_7915);
or UO_884 (O_884,N_9993,N_9276);
and UO_885 (O_885,N_9857,N_7798);
and UO_886 (O_886,N_7585,N_9175);
or UO_887 (O_887,N_9339,N_8735);
and UO_888 (O_888,N_9750,N_7538);
nor UO_889 (O_889,N_8165,N_9668);
nor UO_890 (O_890,N_9966,N_8255);
and UO_891 (O_891,N_9829,N_7965);
nand UO_892 (O_892,N_8512,N_9458);
or UO_893 (O_893,N_8362,N_7724);
nor UO_894 (O_894,N_8486,N_8077);
or UO_895 (O_895,N_9192,N_9662);
nand UO_896 (O_896,N_8243,N_7771);
nand UO_897 (O_897,N_7672,N_9431);
nand UO_898 (O_898,N_9461,N_7698);
nand UO_899 (O_899,N_8770,N_9526);
nand UO_900 (O_900,N_9178,N_8070);
and UO_901 (O_901,N_8309,N_8919);
and UO_902 (O_902,N_8214,N_9096);
and UO_903 (O_903,N_8249,N_9140);
nor UO_904 (O_904,N_7670,N_8946);
or UO_905 (O_905,N_7673,N_7898);
nor UO_906 (O_906,N_7636,N_8126);
or UO_907 (O_907,N_8828,N_8107);
nand UO_908 (O_908,N_7773,N_8821);
or UO_909 (O_909,N_9034,N_9948);
or UO_910 (O_910,N_7931,N_7596);
and UO_911 (O_911,N_8908,N_8262);
and UO_912 (O_912,N_7584,N_7728);
nand UO_913 (O_913,N_7692,N_8216);
nand UO_914 (O_914,N_8525,N_8765);
and UO_915 (O_915,N_9538,N_7829);
nand UO_916 (O_916,N_8754,N_9478);
or UO_917 (O_917,N_8533,N_7879);
and UO_918 (O_918,N_8546,N_9040);
or UO_919 (O_919,N_9279,N_7552);
nor UO_920 (O_920,N_8246,N_7883);
nor UO_921 (O_921,N_9007,N_8790);
nor UO_922 (O_922,N_8060,N_7517);
nor UO_923 (O_923,N_9017,N_8006);
nand UO_924 (O_924,N_7542,N_9265);
nand UO_925 (O_925,N_8099,N_8918);
nor UO_926 (O_926,N_9370,N_9151);
nand UO_927 (O_927,N_8370,N_9879);
or UO_928 (O_928,N_8801,N_7570);
and UO_929 (O_929,N_9207,N_9169);
or UO_930 (O_930,N_8799,N_7681);
nor UO_931 (O_931,N_8344,N_9753);
or UO_932 (O_932,N_8261,N_8112);
and UO_933 (O_933,N_8064,N_8802);
and UO_934 (O_934,N_8664,N_9804);
nand UO_935 (O_935,N_8004,N_8177);
nand UO_936 (O_936,N_8209,N_7618);
nor UO_937 (O_937,N_9144,N_8087);
or UO_938 (O_938,N_8197,N_9774);
xnor UO_939 (O_939,N_7669,N_7803);
or UO_940 (O_940,N_9733,N_9870);
or UO_941 (O_941,N_8701,N_8749);
and UO_942 (O_942,N_7583,N_9274);
or UO_943 (O_943,N_9340,N_9968);
and UO_944 (O_944,N_9623,N_8203);
nor UO_945 (O_945,N_8220,N_8443);
or UO_946 (O_946,N_9440,N_8200);
nand UO_947 (O_947,N_9929,N_8871);
and UO_948 (O_948,N_8181,N_8499);
or UO_949 (O_949,N_7970,N_7882);
or UO_950 (O_950,N_9217,N_7716);
nand UO_951 (O_951,N_9342,N_7974);
and UO_952 (O_952,N_7939,N_7800);
nand UO_953 (O_953,N_8361,N_9901);
nor UO_954 (O_954,N_9946,N_9895);
or UO_955 (O_955,N_8234,N_9747);
and UO_956 (O_956,N_8322,N_9511);
or UO_957 (O_957,N_9378,N_7744);
or UO_958 (O_958,N_8657,N_7850);
and UO_959 (O_959,N_8433,N_9838);
nor UO_960 (O_960,N_9495,N_8432);
and UO_961 (O_961,N_7573,N_7904);
and UO_962 (O_962,N_8581,N_9249);
nor UO_963 (O_963,N_9294,N_9519);
nor UO_964 (O_964,N_9444,N_8067);
nor UO_965 (O_965,N_9291,N_8071);
or UO_966 (O_966,N_8973,N_8377);
nand UO_967 (O_967,N_8613,N_8030);
and UO_968 (O_968,N_8961,N_9773);
or UO_969 (O_969,N_8386,N_8399);
or UO_970 (O_970,N_9767,N_9582);
nand UO_971 (O_971,N_7634,N_9601);
nor UO_972 (O_972,N_8797,N_8979);
nor UO_973 (O_973,N_7782,N_9610);
nand UO_974 (O_974,N_8221,N_9649);
or UO_975 (O_975,N_8420,N_9749);
and UO_976 (O_976,N_9137,N_8169);
nand UO_977 (O_977,N_9923,N_8983);
nand UO_978 (O_978,N_9709,N_8048);
nor UO_979 (O_979,N_8244,N_8771);
or UO_980 (O_980,N_9432,N_8873);
nor UO_981 (O_981,N_8522,N_9992);
xnor UO_982 (O_982,N_8456,N_9060);
nand UO_983 (O_983,N_8772,N_9241);
and UO_984 (O_984,N_9930,N_7862);
nand UO_985 (O_985,N_7982,N_8142);
nor UO_986 (O_986,N_9892,N_8835);
nand UO_987 (O_987,N_8175,N_8923);
and UO_988 (O_988,N_8825,N_8418);
nand UO_989 (O_989,N_9931,N_9281);
or UO_990 (O_990,N_9659,N_8247);
nand UO_991 (O_991,N_9198,N_8437);
nand UO_992 (O_992,N_8868,N_9669);
and UO_993 (O_993,N_9633,N_9907);
or UO_994 (O_994,N_9978,N_9240);
nor UO_995 (O_995,N_7943,N_9979);
nor UO_996 (O_996,N_9648,N_8955);
nand UO_997 (O_997,N_7643,N_9263);
nand UO_998 (O_998,N_9918,N_9383);
or UO_999 (O_999,N_8654,N_8208);
or UO_1000 (O_1000,N_9728,N_8627);
nor UO_1001 (O_1001,N_8179,N_9126);
and UO_1002 (O_1002,N_8509,N_9476);
and UO_1003 (O_1003,N_9826,N_8885);
and UO_1004 (O_1004,N_9609,N_9911);
or UO_1005 (O_1005,N_9924,N_9980);
nor UO_1006 (O_1006,N_9501,N_9589);
nand UO_1007 (O_1007,N_9149,N_8424);
nand UO_1008 (O_1008,N_8044,N_7938);
nand UO_1009 (O_1009,N_7537,N_8075);
nor UO_1010 (O_1010,N_9745,N_9416);
and UO_1011 (O_1011,N_8061,N_9932);
nand UO_1012 (O_1012,N_8756,N_9303);
nor UO_1013 (O_1013,N_7847,N_9849);
nand UO_1014 (O_1014,N_8496,N_7646);
nor UO_1015 (O_1015,N_8410,N_8762);
and UO_1016 (O_1016,N_8266,N_9100);
nand UO_1017 (O_1017,N_9943,N_8084);
and UO_1018 (O_1018,N_8403,N_7536);
nor UO_1019 (O_1019,N_8965,N_9622);
nor UO_1020 (O_1020,N_9065,N_7978);
or UO_1021 (O_1021,N_9113,N_8145);
and UO_1022 (O_1022,N_7817,N_7662);
or UO_1023 (O_1023,N_8180,N_8759);
or UO_1024 (O_1024,N_8495,N_8438);
nor UO_1025 (O_1025,N_7615,N_7936);
or UO_1026 (O_1026,N_7727,N_8299);
nand UO_1027 (O_1027,N_9448,N_8722);
nand UO_1028 (O_1028,N_9156,N_7539);
or UO_1029 (O_1029,N_8637,N_7758);
nand UO_1030 (O_1030,N_9454,N_8019);
or UO_1031 (O_1031,N_9238,N_9270);
nor UO_1032 (O_1032,N_9368,N_8003);
or UO_1033 (O_1033,N_9480,N_9287);
and UO_1034 (O_1034,N_7769,N_7935);
nand UO_1035 (O_1035,N_9759,N_8562);
nand UO_1036 (O_1036,N_8720,N_8292);
nand UO_1037 (O_1037,N_9354,N_8829);
nor UO_1038 (O_1038,N_9697,N_8647);
nand UO_1039 (O_1039,N_8616,N_8388);
or UO_1040 (O_1040,N_9092,N_8622);
nor UO_1041 (O_1041,N_9460,N_9082);
and UO_1042 (O_1042,N_8215,N_9112);
and UO_1043 (O_1043,N_9227,N_9076);
and UO_1044 (O_1044,N_8226,N_8632);
or UO_1045 (O_1045,N_9507,N_9130);
or UO_1046 (O_1046,N_7562,N_8477);
or UO_1047 (O_1047,N_8909,N_9392);
nand UO_1048 (O_1048,N_8652,N_8753);
or UO_1049 (O_1049,N_9045,N_7626);
and UO_1050 (O_1050,N_8287,N_9286);
nor UO_1051 (O_1051,N_8948,N_8804);
nand UO_1052 (O_1052,N_7722,N_7514);
or UO_1053 (O_1053,N_9549,N_8854);
and UO_1054 (O_1054,N_7625,N_8134);
nand UO_1055 (O_1055,N_8360,N_8121);
or UO_1056 (O_1056,N_8656,N_8029);
or UO_1057 (O_1057,N_9429,N_8489);
nand UO_1058 (O_1058,N_7825,N_9821);
nor UO_1059 (O_1059,N_8669,N_8639);
nor UO_1060 (O_1060,N_9475,N_8293);
nor UO_1061 (O_1061,N_8620,N_7996);
or UO_1062 (O_1062,N_8538,N_8901);
or UO_1063 (O_1063,N_7628,N_9158);
and UO_1064 (O_1064,N_7877,N_7591);
nand UO_1065 (O_1065,N_9479,N_8853);
and UO_1066 (O_1066,N_8634,N_7649);
nor UO_1067 (O_1067,N_8844,N_8334);
nor UO_1068 (O_1068,N_9324,N_9967);
nor UO_1069 (O_1069,N_7691,N_9205);
or UO_1070 (O_1070,N_8970,N_8599);
nand UO_1071 (O_1071,N_9690,N_9711);
nand UO_1072 (O_1072,N_8789,N_8411);
nor UO_1073 (O_1073,N_8845,N_8675);
and UO_1074 (O_1074,N_8475,N_8732);
nor UO_1075 (O_1075,N_8471,N_9059);
nand UO_1076 (O_1076,N_8289,N_8964);
and UO_1077 (O_1077,N_8429,N_8748);
nor UO_1078 (O_1078,N_8300,N_7559);
and UO_1079 (O_1079,N_9077,N_9790);
nor UO_1080 (O_1080,N_7635,N_7802);
nor UO_1081 (O_1081,N_9888,N_7944);
nand UO_1082 (O_1082,N_9335,N_9665);
and UO_1083 (O_1083,N_9196,N_9134);
nand UO_1084 (O_1084,N_8113,N_8636);
or UO_1085 (O_1085,N_9720,N_8523);
nor UO_1086 (O_1086,N_7560,N_8640);
and UO_1087 (O_1087,N_7686,N_9201);
or UO_1088 (O_1088,N_8618,N_8615);
nor UO_1089 (O_1089,N_8999,N_8357);
nor UO_1090 (O_1090,N_8592,N_8774);
or UO_1091 (O_1091,N_7745,N_9257);
and UO_1092 (O_1092,N_9179,N_7854);
nand UO_1093 (O_1093,N_8836,N_9934);
nor UO_1094 (O_1094,N_9409,N_9853);
nor UO_1095 (O_1095,N_8354,N_9952);
and UO_1096 (O_1096,N_8131,N_8807);
and UO_1097 (O_1097,N_9117,N_9776);
or UO_1098 (O_1098,N_9085,N_8478);
nand UO_1099 (O_1099,N_8612,N_8025);
nor UO_1100 (O_1100,N_9457,N_7687);
nand UO_1101 (O_1101,N_9873,N_7733);
nand UO_1102 (O_1102,N_8431,N_9581);
or UO_1103 (O_1103,N_8730,N_8757);
nand UO_1104 (O_1104,N_9139,N_8240);
nand UO_1105 (O_1105,N_8397,N_8697);
xnor UO_1106 (O_1106,N_9053,N_9660);
nor UO_1107 (O_1107,N_9047,N_9351);
nand UO_1108 (O_1108,N_7876,N_8775);
nand UO_1109 (O_1109,N_7742,N_9854);
or UO_1110 (O_1110,N_8737,N_9688);
nor UO_1111 (O_1111,N_7697,N_9095);
nor UO_1112 (O_1112,N_9030,N_8237);
nand UO_1113 (O_1113,N_9579,N_9090);
nor UO_1114 (O_1114,N_8709,N_8469);
or UO_1115 (O_1115,N_8415,N_9256);
and UO_1116 (O_1116,N_9110,N_9208);
nand UO_1117 (O_1117,N_8297,N_8847);
or UO_1118 (O_1118,N_9016,N_8413);
or UO_1119 (O_1119,N_8952,N_8817);
and UO_1120 (O_1120,N_8364,N_8741);
or UO_1121 (O_1121,N_9730,N_9823);
nor UO_1122 (O_1122,N_8023,N_8768);
and UO_1123 (O_1123,N_7866,N_9382);
nor UO_1124 (O_1124,N_9226,N_7695);
or UO_1125 (O_1125,N_7762,N_9557);
and UO_1126 (O_1126,N_7595,N_7858);
or UO_1127 (O_1127,N_8605,N_8313);
nand UO_1128 (O_1128,N_9236,N_9974);
nand UO_1129 (O_1129,N_8694,N_8235);
nand UO_1130 (O_1130,N_9013,N_8549);
or UO_1131 (O_1131,N_9919,N_9068);
nand UO_1132 (O_1132,N_8958,N_8482);
nor UO_1133 (O_1133,N_8593,N_9477);
or UO_1134 (O_1134,N_8368,N_8571);
nor UO_1135 (O_1135,N_8427,N_9308);
nand UO_1136 (O_1136,N_8739,N_9302);
nor UO_1137 (O_1137,N_7973,N_9754);
and UO_1138 (O_1138,N_8032,N_9600);
nand UO_1139 (O_1139,N_9326,N_9635);
nor UO_1140 (O_1140,N_9585,N_7751);
and UO_1141 (O_1141,N_9563,N_7863);
nand UO_1142 (O_1142,N_8724,N_9715);
and UO_1143 (O_1143,N_8900,N_8290);
nor UO_1144 (O_1144,N_9253,N_7656);
xnor UO_1145 (O_1145,N_8704,N_8385);
nor UO_1146 (O_1146,N_7706,N_8548);
and UO_1147 (O_1147,N_9661,N_8716);
and UO_1148 (O_1148,N_7593,N_8002);
nor UO_1149 (O_1149,N_7889,N_8280);
and UO_1150 (O_1150,N_8005,N_8407);
or UO_1151 (O_1151,N_9806,N_7950);
nor UO_1152 (O_1152,N_9336,N_8696);
or UO_1153 (O_1153,N_8870,N_9830);
and UO_1154 (O_1154,N_8212,N_9445);
xor UO_1155 (O_1155,N_7768,N_7916);
nor UO_1156 (O_1156,N_9367,N_8982);
and UO_1157 (O_1157,N_9318,N_8294);
nand UO_1158 (O_1158,N_8127,N_7929);
nand UO_1159 (O_1159,N_9394,N_9794);
nor UO_1160 (O_1160,N_7624,N_9459);
nor UO_1161 (O_1161,N_7561,N_9976);
nor UO_1162 (O_1162,N_8186,N_7886);
nor UO_1163 (O_1163,N_9453,N_9765);
or UO_1164 (O_1164,N_9644,N_8384);
and UO_1165 (O_1165,N_9570,N_9500);
nor UO_1166 (O_1166,N_8223,N_9312);
nor UO_1167 (O_1167,N_8378,N_8506);
nand UO_1168 (O_1168,N_8860,N_8811);
and UO_1169 (O_1169,N_9038,N_7736);
or UO_1170 (O_1170,N_9703,N_7632);
xor UO_1171 (O_1171,N_9250,N_8849);
nor UO_1172 (O_1172,N_8779,N_8081);
nand UO_1173 (O_1173,N_8351,N_9497);
nor UO_1174 (O_1174,N_9603,N_9667);
nor UO_1175 (O_1175,N_7551,N_9686);
or UO_1176 (O_1176,N_8507,N_9566);
nor UO_1177 (O_1177,N_8307,N_9996);
nor UO_1178 (O_1178,N_9508,N_9438);
and UO_1179 (O_1179,N_9170,N_7574);
or UO_1180 (O_1180,N_7861,N_9327);
nand UO_1181 (O_1181,N_8328,N_7652);
nand UO_1182 (O_1182,N_9498,N_8998);
nor UO_1183 (O_1183,N_8419,N_9577);
or UO_1184 (O_1184,N_8711,N_9878);
nor UO_1185 (O_1185,N_9061,N_7774);
or UO_1186 (O_1186,N_9521,N_8018);
nor UO_1187 (O_1187,N_8642,N_7571);
or UO_1188 (O_1188,N_9271,N_7604);
nand UO_1189 (O_1189,N_7663,N_8905);
nor UO_1190 (O_1190,N_8421,N_8464);
and UO_1191 (O_1191,N_9195,N_8856);
or UO_1192 (O_1192,N_9866,N_7735);
nor UO_1193 (O_1193,N_9839,N_9466);
or UO_1194 (O_1194,N_9104,N_8713);
and UO_1195 (O_1195,N_9859,N_8206);
or UO_1196 (O_1196,N_8678,N_8879);
nor UO_1197 (O_1197,N_9426,N_8681);
nor UO_1198 (O_1198,N_8945,N_8408);
and UO_1199 (O_1199,N_8183,N_8831);
and UO_1200 (O_1200,N_9288,N_8841);
nand UO_1201 (O_1201,N_9086,N_9572);
nor UO_1202 (O_1202,N_8122,N_8264);
or UO_1203 (O_1203,N_9080,N_9219);
nor UO_1204 (O_1204,N_9122,N_8199);
nand UO_1205 (O_1205,N_7533,N_8609);
or UO_1206 (O_1206,N_8688,N_8213);
and UO_1207 (O_1207,N_9615,N_8218);
nand UO_1208 (O_1208,N_8043,N_8086);
and UO_1209 (O_1209,N_9465,N_9634);
nand UO_1210 (O_1210,N_8376,N_8463);
and UO_1211 (O_1211,N_9962,N_8736);
nand UO_1212 (O_1212,N_8001,N_8725);
and UO_1213 (O_1213,N_7616,N_7556);
nand UO_1214 (O_1214,N_8204,N_7511);
nand UO_1215 (O_1215,N_9181,N_8224);
or UO_1216 (O_1216,N_7918,N_7668);
nand UO_1217 (O_1217,N_7703,N_8316);
and UO_1218 (O_1218,N_7860,N_8597);
nand UO_1219 (O_1219,N_9957,N_9135);
or UO_1220 (O_1220,N_8559,N_9400);
nor UO_1221 (O_1221,N_8222,N_9352);
or UO_1222 (O_1222,N_8080,N_7949);
or UO_1223 (O_1223,N_9121,N_8891);
nand UO_1224 (O_1224,N_9087,N_8476);
or UO_1225 (O_1225,N_8786,N_9052);
and UO_1226 (O_1226,N_8501,N_9739);
and UO_1227 (O_1227,N_8379,N_8173);
nand UO_1228 (O_1228,N_9636,N_8777);
and UO_1229 (O_1229,N_8659,N_9262);
nand UO_1230 (O_1230,N_9969,N_9184);
nor UO_1231 (O_1231,N_9881,N_8684);
nor UO_1232 (O_1232,N_9972,N_8256);
and UO_1233 (O_1233,N_7815,N_7711);
and UO_1234 (O_1234,N_9159,N_8350);
and UO_1235 (O_1235,N_8374,N_8687);
and UO_1236 (O_1236,N_8254,N_8166);
and UO_1237 (O_1237,N_8940,N_7547);
and UO_1238 (O_1238,N_9044,N_8726);
or UO_1239 (O_1239,N_9451,N_7844);
or UO_1240 (O_1240,N_9921,N_9483);
and UO_1241 (O_1241,N_8267,N_9528);
nor UO_1242 (O_1242,N_9927,N_9494);
nor UO_1243 (O_1243,N_7611,N_8861);
nor UO_1244 (O_1244,N_9890,N_9791);
nor UO_1245 (O_1245,N_8114,N_9935);
and UO_1246 (O_1246,N_9022,N_7729);
or UO_1247 (O_1247,N_9744,N_8729);
nand UO_1248 (O_1248,N_8151,N_9527);
nand UO_1249 (O_1249,N_8170,N_8315);
nand UO_1250 (O_1250,N_9264,N_7501);
nor UO_1251 (O_1251,N_7654,N_8103);
nor UO_1252 (O_1252,N_9980,N_9225);
or UO_1253 (O_1253,N_9329,N_9855);
or UO_1254 (O_1254,N_8729,N_7924);
nand UO_1255 (O_1255,N_8367,N_7884);
or UO_1256 (O_1256,N_9307,N_9518);
and UO_1257 (O_1257,N_8814,N_8220);
nor UO_1258 (O_1258,N_9511,N_9629);
or UO_1259 (O_1259,N_9356,N_9196);
and UO_1260 (O_1260,N_8290,N_8593);
and UO_1261 (O_1261,N_9178,N_9601);
nor UO_1262 (O_1262,N_9467,N_8301);
or UO_1263 (O_1263,N_9768,N_9534);
and UO_1264 (O_1264,N_7949,N_9511);
or UO_1265 (O_1265,N_9671,N_8688);
or UO_1266 (O_1266,N_8575,N_8261);
or UO_1267 (O_1267,N_7512,N_8473);
or UO_1268 (O_1268,N_8241,N_9377);
or UO_1269 (O_1269,N_8778,N_9533);
nand UO_1270 (O_1270,N_8479,N_8171);
nor UO_1271 (O_1271,N_8105,N_9324);
or UO_1272 (O_1272,N_9342,N_9445);
and UO_1273 (O_1273,N_8391,N_8610);
nand UO_1274 (O_1274,N_9656,N_7757);
nor UO_1275 (O_1275,N_9160,N_9568);
nand UO_1276 (O_1276,N_9244,N_8261);
nand UO_1277 (O_1277,N_9142,N_7887);
nand UO_1278 (O_1278,N_8336,N_9941);
nand UO_1279 (O_1279,N_9346,N_9957);
nor UO_1280 (O_1280,N_9236,N_8347);
nand UO_1281 (O_1281,N_9802,N_9783);
nor UO_1282 (O_1282,N_9446,N_9921);
nand UO_1283 (O_1283,N_9518,N_8781);
nor UO_1284 (O_1284,N_9283,N_8962);
and UO_1285 (O_1285,N_8397,N_8885);
nor UO_1286 (O_1286,N_8876,N_8858);
and UO_1287 (O_1287,N_7639,N_9979);
nor UO_1288 (O_1288,N_7909,N_9696);
and UO_1289 (O_1289,N_9851,N_8811);
nor UO_1290 (O_1290,N_8041,N_9229);
nand UO_1291 (O_1291,N_8371,N_9570);
and UO_1292 (O_1292,N_8774,N_8741);
and UO_1293 (O_1293,N_7780,N_8390);
and UO_1294 (O_1294,N_9751,N_9967);
nor UO_1295 (O_1295,N_8321,N_8490);
or UO_1296 (O_1296,N_7854,N_8340);
or UO_1297 (O_1297,N_9027,N_8391);
nor UO_1298 (O_1298,N_8079,N_9852);
nand UO_1299 (O_1299,N_9158,N_9001);
or UO_1300 (O_1300,N_9777,N_8227);
nor UO_1301 (O_1301,N_9307,N_8709);
or UO_1302 (O_1302,N_8544,N_9208);
nand UO_1303 (O_1303,N_8825,N_7639);
nor UO_1304 (O_1304,N_7504,N_9448);
nor UO_1305 (O_1305,N_9649,N_8583);
nor UO_1306 (O_1306,N_8406,N_8117);
nand UO_1307 (O_1307,N_8767,N_8778);
or UO_1308 (O_1308,N_9874,N_8289);
nor UO_1309 (O_1309,N_9374,N_9005);
or UO_1310 (O_1310,N_8524,N_7986);
nand UO_1311 (O_1311,N_8632,N_7664);
or UO_1312 (O_1312,N_7502,N_8976);
or UO_1313 (O_1313,N_8978,N_8645);
nand UO_1314 (O_1314,N_9962,N_7693);
and UO_1315 (O_1315,N_9946,N_7942);
and UO_1316 (O_1316,N_9619,N_9688);
or UO_1317 (O_1317,N_8161,N_7521);
nand UO_1318 (O_1318,N_8626,N_8834);
and UO_1319 (O_1319,N_7513,N_7920);
nand UO_1320 (O_1320,N_7952,N_8369);
nand UO_1321 (O_1321,N_7820,N_7728);
nand UO_1322 (O_1322,N_8230,N_7759);
nand UO_1323 (O_1323,N_7874,N_8733);
or UO_1324 (O_1324,N_8715,N_8943);
and UO_1325 (O_1325,N_8010,N_9621);
or UO_1326 (O_1326,N_8151,N_8353);
nand UO_1327 (O_1327,N_9026,N_7821);
nor UO_1328 (O_1328,N_9747,N_9908);
and UO_1329 (O_1329,N_8187,N_7951);
and UO_1330 (O_1330,N_8761,N_8740);
or UO_1331 (O_1331,N_9473,N_9311);
and UO_1332 (O_1332,N_9878,N_9567);
nand UO_1333 (O_1333,N_8341,N_7779);
nor UO_1334 (O_1334,N_8188,N_8570);
nand UO_1335 (O_1335,N_9966,N_9381);
nand UO_1336 (O_1336,N_8213,N_7890);
nand UO_1337 (O_1337,N_7598,N_7859);
and UO_1338 (O_1338,N_8114,N_8465);
and UO_1339 (O_1339,N_9711,N_9469);
and UO_1340 (O_1340,N_8072,N_7820);
and UO_1341 (O_1341,N_9847,N_9044);
xnor UO_1342 (O_1342,N_7691,N_9370);
and UO_1343 (O_1343,N_8246,N_9261);
or UO_1344 (O_1344,N_9298,N_9547);
or UO_1345 (O_1345,N_9950,N_7788);
nand UO_1346 (O_1346,N_9720,N_9879);
nor UO_1347 (O_1347,N_8164,N_8181);
nor UO_1348 (O_1348,N_8631,N_8779);
nand UO_1349 (O_1349,N_8932,N_7792);
or UO_1350 (O_1350,N_8837,N_9902);
and UO_1351 (O_1351,N_9324,N_8097);
and UO_1352 (O_1352,N_8712,N_8569);
and UO_1353 (O_1353,N_8607,N_7904);
nor UO_1354 (O_1354,N_8929,N_9022);
nor UO_1355 (O_1355,N_8920,N_8239);
nand UO_1356 (O_1356,N_9380,N_9775);
nor UO_1357 (O_1357,N_8755,N_7750);
or UO_1358 (O_1358,N_8755,N_7941);
and UO_1359 (O_1359,N_8748,N_8308);
nor UO_1360 (O_1360,N_7658,N_9906);
nor UO_1361 (O_1361,N_8629,N_8895);
or UO_1362 (O_1362,N_8774,N_7936);
nor UO_1363 (O_1363,N_7953,N_9592);
nand UO_1364 (O_1364,N_8292,N_9043);
nand UO_1365 (O_1365,N_9391,N_9584);
nor UO_1366 (O_1366,N_8769,N_8276);
nor UO_1367 (O_1367,N_7547,N_7975);
nor UO_1368 (O_1368,N_7901,N_8232);
or UO_1369 (O_1369,N_7557,N_8955);
nand UO_1370 (O_1370,N_8986,N_9636);
or UO_1371 (O_1371,N_7995,N_9106);
and UO_1372 (O_1372,N_8600,N_9650);
nand UO_1373 (O_1373,N_9750,N_8183);
nand UO_1374 (O_1374,N_9787,N_8596);
and UO_1375 (O_1375,N_9300,N_9303);
or UO_1376 (O_1376,N_8292,N_8471);
or UO_1377 (O_1377,N_9413,N_8216);
nand UO_1378 (O_1378,N_7700,N_8902);
and UO_1379 (O_1379,N_9888,N_7667);
or UO_1380 (O_1380,N_9635,N_7715);
nor UO_1381 (O_1381,N_7517,N_9288);
nand UO_1382 (O_1382,N_8376,N_9878);
and UO_1383 (O_1383,N_8506,N_9800);
nor UO_1384 (O_1384,N_7635,N_9054);
nor UO_1385 (O_1385,N_7804,N_8733);
nor UO_1386 (O_1386,N_9576,N_8893);
nand UO_1387 (O_1387,N_8924,N_9582);
or UO_1388 (O_1388,N_8531,N_8618);
nor UO_1389 (O_1389,N_8600,N_9604);
or UO_1390 (O_1390,N_9517,N_7756);
nand UO_1391 (O_1391,N_9682,N_8704);
or UO_1392 (O_1392,N_8693,N_9163);
or UO_1393 (O_1393,N_8058,N_8385);
nand UO_1394 (O_1394,N_8532,N_7752);
nand UO_1395 (O_1395,N_8501,N_8091);
and UO_1396 (O_1396,N_8045,N_9930);
nand UO_1397 (O_1397,N_8819,N_9530);
and UO_1398 (O_1398,N_8335,N_8503);
nor UO_1399 (O_1399,N_9957,N_9549);
and UO_1400 (O_1400,N_8808,N_8049);
nand UO_1401 (O_1401,N_9077,N_7616);
and UO_1402 (O_1402,N_7953,N_7817);
nand UO_1403 (O_1403,N_7776,N_8845);
and UO_1404 (O_1404,N_7660,N_8733);
nor UO_1405 (O_1405,N_7728,N_8093);
nand UO_1406 (O_1406,N_8368,N_7815);
nand UO_1407 (O_1407,N_7905,N_7533);
nand UO_1408 (O_1408,N_9943,N_9549);
and UO_1409 (O_1409,N_9435,N_8105);
or UO_1410 (O_1410,N_8362,N_9155);
or UO_1411 (O_1411,N_8435,N_9279);
nor UO_1412 (O_1412,N_9937,N_7919);
nor UO_1413 (O_1413,N_9755,N_8474);
nand UO_1414 (O_1414,N_8241,N_8076);
and UO_1415 (O_1415,N_9484,N_9524);
or UO_1416 (O_1416,N_9606,N_9564);
nor UO_1417 (O_1417,N_9807,N_9100);
nand UO_1418 (O_1418,N_8184,N_8819);
nand UO_1419 (O_1419,N_7914,N_9681);
xnor UO_1420 (O_1420,N_9098,N_8597);
or UO_1421 (O_1421,N_8105,N_7868);
and UO_1422 (O_1422,N_9089,N_9401);
or UO_1423 (O_1423,N_8053,N_9418);
or UO_1424 (O_1424,N_8079,N_7966);
nand UO_1425 (O_1425,N_9519,N_8010);
nand UO_1426 (O_1426,N_8812,N_9321);
or UO_1427 (O_1427,N_7939,N_8283);
nor UO_1428 (O_1428,N_8200,N_9887);
nor UO_1429 (O_1429,N_9703,N_8548);
nor UO_1430 (O_1430,N_9247,N_9858);
and UO_1431 (O_1431,N_9435,N_8527);
nand UO_1432 (O_1432,N_7673,N_8420);
and UO_1433 (O_1433,N_9267,N_8182);
and UO_1434 (O_1434,N_7645,N_7612);
nand UO_1435 (O_1435,N_8323,N_9558);
nor UO_1436 (O_1436,N_8899,N_9976);
and UO_1437 (O_1437,N_9319,N_8653);
nor UO_1438 (O_1438,N_9548,N_8413);
nand UO_1439 (O_1439,N_8694,N_8495);
nor UO_1440 (O_1440,N_9175,N_9984);
and UO_1441 (O_1441,N_8682,N_7913);
nor UO_1442 (O_1442,N_8213,N_8820);
or UO_1443 (O_1443,N_8466,N_9286);
and UO_1444 (O_1444,N_9348,N_9351);
or UO_1445 (O_1445,N_8263,N_7976);
nand UO_1446 (O_1446,N_9750,N_9123);
or UO_1447 (O_1447,N_8589,N_7979);
nor UO_1448 (O_1448,N_7849,N_9348);
and UO_1449 (O_1449,N_8958,N_9033);
nor UO_1450 (O_1450,N_8274,N_9361);
and UO_1451 (O_1451,N_8306,N_9753);
nor UO_1452 (O_1452,N_9209,N_9911);
and UO_1453 (O_1453,N_9732,N_7803);
nand UO_1454 (O_1454,N_9316,N_7839);
or UO_1455 (O_1455,N_9033,N_9168);
and UO_1456 (O_1456,N_7989,N_7551);
and UO_1457 (O_1457,N_8510,N_9448);
nor UO_1458 (O_1458,N_7814,N_7654);
and UO_1459 (O_1459,N_9583,N_8998);
and UO_1460 (O_1460,N_8051,N_9989);
or UO_1461 (O_1461,N_7559,N_8152);
nand UO_1462 (O_1462,N_9064,N_9701);
nor UO_1463 (O_1463,N_8239,N_9328);
and UO_1464 (O_1464,N_7747,N_8225);
nand UO_1465 (O_1465,N_9386,N_8750);
or UO_1466 (O_1466,N_9030,N_9397);
or UO_1467 (O_1467,N_8985,N_9299);
nand UO_1468 (O_1468,N_7866,N_7667);
nand UO_1469 (O_1469,N_8989,N_8943);
nand UO_1470 (O_1470,N_7658,N_9700);
and UO_1471 (O_1471,N_9048,N_7711);
or UO_1472 (O_1472,N_8694,N_7768);
xnor UO_1473 (O_1473,N_8993,N_9195);
nand UO_1474 (O_1474,N_8579,N_8323);
nor UO_1475 (O_1475,N_9121,N_9271);
and UO_1476 (O_1476,N_9347,N_8371);
or UO_1477 (O_1477,N_7533,N_8824);
and UO_1478 (O_1478,N_7988,N_9512);
nand UO_1479 (O_1479,N_9863,N_9423);
nand UO_1480 (O_1480,N_8281,N_9857);
nor UO_1481 (O_1481,N_7829,N_8756);
nor UO_1482 (O_1482,N_8207,N_8162);
and UO_1483 (O_1483,N_9841,N_9600);
or UO_1484 (O_1484,N_8330,N_9965);
nand UO_1485 (O_1485,N_8242,N_8345);
or UO_1486 (O_1486,N_8489,N_8410);
and UO_1487 (O_1487,N_9438,N_9172);
nor UO_1488 (O_1488,N_9147,N_8164);
nor UO_1489 (O_1489,N_9389,N_8410);
and UO_1490 (O_1490,N_8468,N_7540);
or UO_1491 (O_1491,N_8020,N_8348);
or UO_1492 (O_1492,N_7903,N_8888);
or UO_1493 (O_1493,N_9705,N_8445);
or UO_1494 (O_1494,N_9785,N_9374);
nand UO_1495 (O_1495,N_9148,N_9865);
nor UO_1496 (O_1496,N_8112,N_9332);
and UO_1497 (O_1497,N_8923,N_9483);
nand UO_1498 (O_1498,N_9828,N_9980);
nand UO_1499 (O_1499,N_9325,N_9041);
endmodule